`include "common.h"

module chip_6502(
  input eclk, ereset,
  output ab0,
  output ab1,
  output ab2,
  output ab3,
  output ab4,
  output ab5,
  output ab6,
  output ab7,
  output ab8,
  output ab9,
  output ab10,
  output ab11,
  output ab12,
  output ab13,
  output ab14,
  output ab15,
  input db0_i,
  output db0_o,
  output db0_t,
  input db1_i,
  output db1_o,
  output db1_t,
  input db2_i,
  output db2_o,
  output db2_t,
  input db3_i,
  output db3_o,
  output db3_t,
  input db4_i,
  output db4_o,
  output db4_t,
  input db5_i,
  output db5_o,
  output db5_t,
  input db6_i,
  output db6_o,
  output db6_t,
  input db7_i,
  output db7_o,
  output db7_t,
  input res,
  output rw,
  output sync,
  input so,
  input clk0,
  output clk1out,
  output clk2out,
  input rdy,
  input nmi,
  input irq
);

  wire signed [`W-1:0] DBNeg_i0;
  wire signed [`W-1:0] DBNeg_i1;
  wire signed [`W-1:0] DBNeg_i2;
  wire signed [`W-1:0] DBNeg_i3;
  wire signed [`W-1:0] DBNeg_v;
  wire signed [`W-1:0] n344_i0;
  wire signed [`W-1:0] n344_i1;
  wire signed [`W-1:0] n344_i2;
  wire signed [`W-1:0] n344_i3;
  wire signed [`W-1:0] n344_i4;
  wire signed [`W-1:0] n344_v;
  wire signed [`W-1:0] n345_i0;
  wire signed [`W-1:0] n345_i1;
  wire signed [`W-1:0] n345_i2;
  wire signed [`W-1:0] n345_i3;
  wire signed [`W-1:0] n345_v;
  wire signed [`W-1:0] n347_i0;
  wire signed [`W-1:0] n347_i1;
  wire signed [`W-1:0] n347_i2;
  wire signed [`W-1:0] n347_i3;
  wire signed [`W-1:0] n347_i4;
  wire signed [`W-1:0] n347_v;
  wire signed [`W-1:0] n340_i0;
  wire signed [`W-1:0] n340_i1;
  wire signed [`W-1:0] n340_i2;
  wire signed [`W-1:0] n340_v;
  wire signed [`W-1:0] op_T4_i0;
  wire signed [`W-1:0] op_T4_i1;
  wire signed [`W-1:0] op_T4_i2;
  wire signed [`W-1:0] op_T4_v;
  wire signed [`W-1:0] x_op_T3_ind_y_i0;
  wire signed [`W-1:0] x_op_T3_ind_y_i1;
  wire signed [`W-1:0] x_op_T3_ind_y_i2;
  wire signed [`W-1:0] x_op_T3_ind_y_v;
  wire signed [`W-1:0] p3_i0;
  wire signed [`W-1:0] p3_i1;
  wire signed [`W-1:0] p3_v;
  wire signed [`W-1:0] ab13_i0;
  wire signed [`W-1:0] ab13_i1;
  wire signed [`W-1:0] ab13_i2;
  wire signed [`W-1:0] ab13_v;
  wire signed [`W-1:0] n298_i0;
  wire signed [`W-1:0] n298_i1;
  wire signed [`W-1:0] n298_i2;
  wire signed [`W-1:0] n298_v;
  wire signed [`W-1:0] n299_i0;
  wire signed [`W-1:0] n299_i1;
  wire signed [`W-1:0] n299_i2;
  wire signed [`W-1:0] n299_v;
  wire signed [`W-1:0] n296_i0;
  wire signed [`W-1:0] n296_i1;
  wire signed [`W-1:0] n296_i2;
  wire signed [`W-1:0] n296_i3;
  wire signed [`W-1:0] n296_i4;
  wire signed [`W-1:0] n296_i5;
  wire signed [`W-1:0] n296_v;
  wire signed [`W-1:0] n297_i0;
  wire signed [`W-1:0] n297_i1;
  wire signed [`W-1:0] n297_i2;
  wire signed [`W-1:0] n297_v;
  wire signed [`W-1:0] pipeUNK20_i0;
  wire signed [`W-1:0] pipeUNK20_i1;
  wire signed [`W-1:0] pipeUNK20_v;
  wire signed [`W-1:0] __AxB1__C01_i0;
  wire signed [`W-1:0] __AxB1__C01_i1;
  wire signed [`W-1:0] __AxB1__C01_i2;
  wire signed [`W-1:0] __AxB1__C01_v;
  wire signed [`W-1:0] pch1_i0;
  wire signed [`W-1:0] pch1_i1;
  wire signed [`W-1:0] pch1_i2;
  wire signed [`W-1:0] pch1_v;
  wire signed [`W-1:0] n293_i0;
  wire signed [`W-1:0] n293_i1;
  wire signed [`W-1:0] n293_i2;
  wire signed [`W-1:0] n293_i3;
  wire signed [`W-1:0] n293_i4;
  wire signed [`W-1:0] n293_v;
  wire signed [`W-1:0] n597_i0;
  wire signed [`W-1:0] n597_i1;
  wire signed [`W-1:0] n597_v;
  wire signed [`W-1:0] n291_i0;
  wire signed [`W-1:0] n291_i1;
  wire signed [`W-1:0] n291_i2;
  wire signed [`W-1:0] n291_i3;
  wire signed [`W-1:0] n291_v;
  wire signed [`W-1:0] n270_i0;
  wire signed [`W-1:0] n270_i1;
  wire signed [`W-1:0] n270_i2;
  wire signed [`W-1:0] n270_i3;
  wire signed [`W-1:0] n270_i4;
  wire signed [`W-1:0] n270_i5;
  wire signed [`W-1:0] n270_i6;
  wire signed [`W-1:0] n270_v;
  wire signed [`W-1:0] op_T0_jsr_i0;
  wire signed [`W-1:0] op_T0_jsr_i1;
  wire signed [`W-1:0] op_T0_jsr_i2;
  wire signed [`W-1:0] op_T0_jsr_i3;
  wire signed [`W-1:0] op_T0_jsr_v;
  wire signed [`W-1:0] n272_i0;
  wire signed [`W-1:0] n272_i1;
  wire signed [`W-1:0] n272_i2;
  wire signed [`W-1:0] n272_i3;
  wire signed [`W-1:0] n272_v;
  wire signed [`W-1:0] op_T2_abs_access_i0;
  wire signed [`W-1:0] op_T2_abs_access_i1;
  wire signed [`W-1:0] op_T2_abs_access_i2;
  wire signed [`W-1:0] op_T2_abs_access_i3;
  wire signed [`W-1:0] op_T2_abs_access_i4;
  wire signed [`W-1:0] op_T2_abs_access_v;
  wire signed [`W-1:0] __AxBxC_3_i0;
  wire signed [`W-1:0] __AxBxC_3_i1;
  wire signed [`W-1:0] __AxBxC_3_i2;
  wire signed [`W-1:0] __AxBxC_3_v;
  wire signed [`W-1:0] n275_i0;
  wire signed [`W-1:0] n275_i1;
  wire signed [`W-1:0] n275_i2;
  wire signed [`W-1:0] n275_v;
  wire signed [`W-1:0] notalu2_i0;
  wire signed [`W-1:0] notalu2_i1;
  wire signed [`W-1:0] notalu2_v;
  wire signed [`W-1:0] n277_i0;
  wire signed [`W-1:0] n277_i1;
  wire signed [`W-1:0] n277_i2;
  wire signed [`W-1:0] n277_i3;
  wire signed [`W-1:0] n277_i4;
  wire signed [`W-1:0] n277_i5;
  wire signed [`W-1:0] n277_v;
  wire signed [`W-1:0] n278_i0;
  wire signed [`W-1:0] n278_i1;
  wire signed [`W-1:0] n278_i2;
  wire signed [`W-1:0] n278_v;
  wire signed [`W-1:0] n279_i0;
  wire signed [`W-1:0] n279_i1;
  wire signed [`W-1:0] n279_i2;
  wire signed [`W-1:0] n279_v;
  wire signed [`W-1:0] n108_i0;
  wire signed [`W-1:0] n108_i1;
  wire signed [`W-1:0] n108_i2;
  wire signed [`W-1:0] n108_v;
  wire signed [`W-1:0] n109_i0;
  wire signed [`W-1:0] n109_i1;
  wire signed [`W-1:0] n109_i2;
  wire signed [`W-1:0] n109_v;
  wire signed [`W-1:0] n102_i0;
  wire signed [`W-1:0] n102_i1;
  wire signed [`W-1:0] n102_i2;
  wire signed [`W-1:0] n102_v;
  wire signed [`W-1:0] irq_i0;
  wire signed [`W-1:0] irq_i1;
  wire signed [`W-1:0] irq_v;
  wire signed [`W-1:0] n101_i0;
  wire signed [`W-1:0] n101_i1;
  wire signed [`W-1:0] n101_v;
  wire signed [`W-1:0] _ABL1_i0;
  wire signed [`W-1:0] _ABL1_i1;
  wire signed [`W-1:0] _ABL1_i2;
  wire signed [`W-1:0] _ABL1_v;
  wire signed [`W-1:0] n104_i0;
  wire signed [`W-1:0] n104_i1;
  wire signed [`W-1:0] n104_i2;
  wire signed [`W-1:0] n104_v;
  wire signed [`W-1:0] n105_i0;
  wire signed [`W-1:0] n105_i1;
  wire signed [`W-1:0] n105_i2;
  wire signed [`W-1:0] n105_i3;
  wire signed [`W-1:0] n105_v;
  wire signed [`W-1:0] pipeUNK04_i0;
  wire signed [`W-1:0] pipeUNK04_i1;
  wire signed [`W-1:0] pipeUNK04_v;
  wire signed [`W-1:0] x1_i0;
  wire signed [`W-1:0] x1_i1;
  wire signed [`W-1:0] x1_i2;
  wire signed [`W-1:0] x1_v;
  wire signed [`W-1:0] n91_i0;
  wire signed [`W-1:0] n91_i1;
  wire signed [`W-1:0] n91_i2;
  wire signed [`W-1:0] n91_i3;
  wire signed [`W-1:0] n91_v;
  wire signed [`W-1:0] n90_i0;
  wire signed [`W-1:0] n90_i1;
  wire signed [`W-1:0] n90_i2;
  wire signed [`W-1:0] n90_i3;
  wire signed [`W-1:0] n90_i4;
  wire signed [`W-1:0] n90_v;
  wire signed [`W-1:0] n93_i0;
  wire signed [`W-1:0] n93_i1;
  wire signed [`W-1:0] n93_i2;
  wire signed [`W-1:0] n93_v;
  wire signed [`W-1:0] _ABH3_i0;
  wire signed [`W-1:0] _ABH3_i1;
  wire signed [`W-1:0] _ABH3_i2;
  wire signed [`W-1:0] _ABH3_v;
  wire signed [`W-1:0] n95_i0;
  wire signed [`W-1:0] n95_i1;
  wire signed [`W-1:0] n95_v;
  wire signed [`W-1:0] n94_i0;
  wire signed [`W-1:0] n94_i1;
  wire signed [`W-1:0] n94_v;
  wire signed [`W-1:0] dor0_i0;
  wire signed [`W-1:0] dor0_i1;
  wire signed [`W-1:0] dor0_i2;
  wire signed [`W-1:0] dor0_i3;
  wire signed [`W-1:0] dor0_i4;
  wire signed [`W-1:0] dor0_v;
  wire signed [`W-1:0] alub3_i0;
  wire signed [`W-1:0] alub3_i1;
  wire signed [`W-1:0] alub3_i2;
  wire signed [`W-1:0] alub3_i3;
  wire signed [`W-1:0] alub3_i4;
  wire signed [`W-1:0] alub3_v;
  wire signed [`W-1:0] op_T0_eor_i0;
  wire signed [`W-1:0] op_T0_eor_i1;
  wire signed [`W-1:0] op_T0_eor_i2;
  wire signed [`W-1:0] op_T0_eor_v;
  wire signed [`W-1:0] pd0_clearIR_i0;
  wire signed [`W-1:0] pd0_clearIR_i1;
  wire signed [`W-1:0] pd0_clearIR_i2;
  wire signed [`W-1:0] pd0_clearIR_i3;
  wire signed [`W-1:0] pd0_clearIR_i4;
  wire signed [`W-1:0] pd0_clearIR_v;
  wire signed [`W-1:0] n1621_i0;
  wire signed [`W-1:0] n1621_i1;
  wire signed [`W-1:0] n1621_i2;
  wire signed [`W-1:0] n1621_v;
  wire signed [`W-1:0] n1620_i0;
  wire signed [`W-1:0] n1620_i1;
  wire signed [`W-1:0] n1620_i2;
  wire signed [`W-1:0] n1620_v;
  wire signed [`W-1:0] alua6_i0;
  wire signed [`W-1:0] alua6_i1;
  wire signed [`W-1:0] alua6_i2;
  wire signed [`W-1:0] alua6_i3;
  wire signed [`W-1:0] alua6_v;
  wire signed [`W-1:0] ir1_i0;
  wire signed [`W-1:0] ir1_i1;
  wire signed [`W-1:0] ir1_i2;
  wire signed [`W-1:0] ir1_i3;
  wire signed [`W-1:0] ir1_v;
  wire signed [`W-1:0] n1625_i0;
  wire signed [`W-1:0] n1625_i1;
  wire signed [`W-1:0] n1625_v;
  wire signed [`W-1:0] n1624_i0;
  wire signed [`W-1:0] n1624_i1;
  wire signed [`W-1:0] n1624_v;
  wire signed [`W-1:0] n1629_i0;
  wire signed [`W-1:0] n1629_i1;
  wire signed [`W-1:0] n1629_i2;
  wire signed [`W-1:0] n1629_v;
  wire signed [`W-1:0] aluanandb0_i0;
  wire signed [`W-1:0] aluanandb0_i1;
  wire signed [`W-1:0] aluanandb0_i2;
  wire signed [`W-1:0] aluanandb0_i3;
  wire signed [`W-1:0] aluanandb0_i4;
  wire signed [`W-1:0] aluanandb0_i5;
  wire signed [`W-1:0] aluanandb0_v;
  wire signed [`W-1:0] n559_i0;
  wire signed [`W-1:0] n559_i1;
  wire signed [`W-1:0] n559_v;
  wire signed [`W-1:0] _AxB_0__C0in_i0;
  wire signed [`W-1:0] _AxB_0__C0in_i1;
  wire signed [`W-1:0] _AxB_0__C0in_i2;
  wire signed [`W-1:0] _AxB_0__C0in_v;
  wire signed [`W-1:0] pipe_T0_i0;
  wire signed [`W-1:0] pipe_T0_i1;
  wire signed [`W-1:0] pipe_T0_i2;
  wire signed [`W-1:0] pipe_T0_v;
  wire signed [`W-1:0] n556_i0;
  wire signed [`W-1:0] n556_i1;
  wire signed [`W-1:0] n556_i2;
  wire signed [`W-1:0] n556_v;
  wire signed [`W-1:0] n551_i0;
  wire signed [`W-1:0] n551_i1;
  wire signed [`W-1:0] n551_i2;
  wire signed [`W-1:0] n551_v;
  wire signed [`W-1:0] n550_i0;
  wire signed [`W-1:0] n550_i1;
  wire signed [`W-1:0] n550_i2;
  wire signed [`W-1:0] n550_v;
  wire signed [`W-1:0] n553_i0;
  wire signed [`W-1:0] n553_i1;
  wire signed [`W-1:0] n553_i2;
  wire signed [`W-1:0] n553_v;
  wire signed [`W-1:0] op_T0_php_pha_i0;
  wire signed [`W-1:0] op_T0_php_pha_i1;
  wire signed [`W-1:0] op_T0_php_pha_i2;
  wire signed [`W-1:0] op_T0_php_pha_v;
  wire signed [`W-1:0] n1199_i0;
  wire signed [`W-1:0] n1199_i1;
  wire signed [`W-1:0] n1199_i2;
  wire signed [`W-1:0] n1199_v;
  wire signed [`W-1:0] n1191_i0;
  wire signed [`W-1:0] n1191_i1;
  wire signed [`W-1:0] n1191_i2;
  wire signed [`W-1:0] n1191_v;
  wire signed [`W-1:0] n1190_i0;
  wire signed [`W-1:0] n1190_i1;
  wire signed [`W-1:0] n1190_i2;
  wire signed [`W-1:0] n1190_v;
  wire signed [`W-1:0] n_0_ADL2_i0;
  wire signed [`W-1:0] n_0_ADL2_i1;
  wire signed [`W-1:0] n_0_ADL2_i2;
  wire signed [`W-1:0] n_0_ADL2_v;
  wire signed [`W-1:0] n1192_i0;
  wire signed [`W-1:0] n1192_i1;
  wire signed [`W-1:0] n1192_i2;
  wire signed [`W-1:0] n1192_v;
  wire signed [`W-1:0] n1195_i0;
  wire signed [`W-1:0] n1195_i1;
  wire signed [`W-1:0] n1195_i2;
  wire signed [`W-1:0] n1195_i3;
  wire signed [`W-1:0] n1195_v;
  wire signed [`W-1:0] n1194_i0;
  wire signed [`W-1:0] n1194_i1;
  wire signed [`W-1:0] n1194_i2;
  wire signed [`W-1:0] n1194_i3;
  wire signed [`W-1:0] n1194_v;
  wire signed [`W-1:0] __AxBxC_6_i0;
  wire signed [`W-1:0] __AxBxC_6_i1;
  wire signed [`W-1:0] __AxBxC_6_i2;
  wire signed [`W-1:0] __AxBxC_6_v;
  wire signed [`W-1:0] op_SUMS_i0;
  wire signed [`W-1:0] op_SUMS_i1;
  wire signed [`W-1:0] op_SUMS_i2;
  wire signed [`W-1:0] op_SUMS_v;
  wire signed [`W-1:0] n1177_i0;
  wire signed [`W-1:0] n1177_i1;
  wire signed [`W-1:0] n1177_v;
  wire signed [`W-1:0] pipeUNK21_i0;
  wire signed [`W-1:0] pipeUNK21_i1;
  wire signed [`W-1:0] pipeUNK21_v;
  wire signed [`W-1:0] n1175_i0;
  wire signed [`W-1:0] n1175_i1;
  wire signed [`W-1:0] n1175_i2;
  wire signed [`W-1:0] n1175_i3;
  wire signed [`W-1:0] n1175_v;
  wire signed [`W-1:0] _op_branch_bit7_i0;
  wire signed [`W-1:0] _op_branch_bit7_i1;
  wire signed [`W-1:0] _op_branch_bit7_i2;
  wire signed [`W-1:0] _op_branch_bit7_i3;
  wire signed [`W-1:0] _op_branch_bit7_i4;
  wire signed [`W-1:0] _op_branch_bit7_v;
  wire signed [`W-1:0] x_op_T0_tya_i0;
  wire signed [`W-1:0] x_op_T0_tya_i1;
  wire signed [`W-1:0] x_op_T0_tya_i2;
  wire signed [`W-1:0] x_op_T0_tya_v;
  wire signed [`W-1:0] clk0_i0;
  wire signed [`W-1:0] clk0_i1;
  wire signed [`W-1:0] clk0_i2;
  wire signed [`W-1:0] clk0_v;
  wire signed [`W-1:0] n1170_i0;
  wire signed [`W-1:0] n1170_i1;
  wire signed [`W-1:0] n1170_i2;
  wire signed [`W-1:0] n1170_v;
  wire signed [`W-1:0] n1179_i0;
  wire signed [`W-1:0] n1179_i1;
  wire signed [`W-1:0] n1179_i2;
  wire signed [`W-1:0] n1179_v;
  wire signed [`W-1:0] n1178_i0;
  wire signed [`W-1:0] n1178_i1;
  wire signed [`W-1:0] n1178_i2;
  wire signed [`W-1:0] n1178_v;
  wire signed [`W-1:0] n510_i0;
  wire signed [`W-1:0] n510_i1;
  wire signed [`W-1:0] n510_i2;
  wire signed [`W-1:0] n510_v;
  wire signed [`W-1:0] n513_i0;
  wire signed [`W-1:0] n513_i1;
  wire signed [`W-1:0] n513_i2;
  wire signed [`W-1:0] n513_v;
  wire signed [`W-1:0] C01_i0;
  wire signed [`W-1:0] C01_i1;
  wire signed [`W-1:0] C01_i2;
  wire signed [`W-1:0] C01_i3;
  wire signed [`W-1:0] C01_v;
  wire signed [`W-1:0] notidl3_i0;
  wire signed [`W-1:0] notidl3_i1;
  wire signed [`W-1:0] notidl3_v;
  wire signed [`W-1:0] sb2_i0;
  wire signed [`W-1:0] sb2_i1;
  wire signed [`W-1:0] sb2_i2;
  wire signed [`W-1:0] sb2_i3;
  wire signed [`W-1:0] sb2_i4;
  wire signed [`W-1:0] sb2_i5;
  wire signed [`W-1:0] sb2_i6;
  wire signed [`W-1:0] sb2_i7;
  wire signed [`W-1:0] sb2_i8;
  wire signed [`W-1:0] sb2_i9;
  wire signed [`W-1:0] sb2_i10;
  wire signed [`W-1:0] sb2_i11;
  wire signed [`W-1:0] sb2_i12;
  wire signed [`W-1:0] sb2_v;
  wire signed [`W-1:0] n512_i0;
  wire signed [`W-1:0] n512_i1;
  wire signed [`W-1:0] n512_v;
  wire signed [`W-1:0] n1281_i0;
  wire signed [`W-1:0] n1281_i1;
  wire signed [`W-1:0] n1281_i2;
  wire signed [`W-1:0] n1281_v;
  wire signed [`W-1:0] pipeUNK12_i0;
  wire signed [`W-1:0] pipeUNK12_i1;
  wire signed [`W-1:0] pipeUNK12_v;
  wire signed [`W-1:0] adl1_i0;
  wire signed [`W-1:0] adl1_i1;
  wire signed [`W-1:0] adl1_i2;
  wire signed [`W-1:0] adl1_i3;
  wire signed [`W-1:0] adl1_i4;
  wire signed [`W-1:0] adl1_i5;
  wire signed [`W-1:0] adl1_i6;
  wire signed [`W-1:0] adl1_i7;
  wire signed [`W-1:0] adl1_i8;
  wire signed [`W-1:0] adl1_v;
  wire signed [`W-1:0] n515_i0;
  wire signed [`W-1:0] n515_i1;
  wire signed [`W-1:0] n515_i2;
  wire signed [`W-1:0] n515_v;
  wire signed [`W-1:0] fetch_i0;
  wire signed [`W-1:0] fetch_i1;
  wire signed [`W-1:0] fetch_i2;
  wire signed [`W-1:0] fetch_i3;
  wire signed [`W-1:0] fetch_i4;
  wire signed [`W-1:0] fetch_i5;
  wire signed [`W-1:0] fetch_i6;
  wire signed [`W-1:0] fetch_i7;
  wire signed [`W-1:0] fetch_i8;
  wire signed [`W-1:0] fetch_i9;
  wire signed [`W-1:0] fetch_i10;
  wire signed [`W-1:0] fetch_v;
  wire signed [`W-1:0] n1289_i0;
  wire signed [`W-1:0] n1289_i1;
  wire signed [`W-1:0] n1289_i2;
  wire signed [`W-1:0] n1289_v;
  wire signed [`W-1:0] notdor2_i0;
  wire signed [`W-1:0] notdor2_i1;
  wire signed [`W-1:0] notdor2_v;
  wire signed [`W-1:0] n1579_i0;
  wire signed [`W-1:0] n1579_i1;
  wire signed [`W-1:0] n1579_v;
  wire signed [`W-1:0] n1578_i0;
  wire signed [`W-1:0] n1578_i1;
  wire signed [`W-1:0] n1578_i2;
  wire signed [`W-1:0] n1578_v;
  wire signed [`W-1:0] n689_i0;
  wire signed [`W-1:0] n689_i1;
  wire signed [`W-1:0] n689_i2;
  wire signed [`W-1:0] n689_v;
  wire signed [`W-1:0] sb7_i0;
  wire signed [`W-1:0] sb7_i1;
  wire signed [`W-1:0] sb7_i2;
  wire signed [`W-1:0] sb7_i3;
  wire signed [`W-1:0] sb7_i4;
  wire signed [`W-1:0] sb7_i5;
  wire signed [`W-1:0] sb7_i6;
  wire signed [`W-1:0] sb7_i7;
  wire signed [`W-1:0] sb7_i8;
  wire signed [`W-1:0] sb7_i9;
  wire signed [`W-1:0] sb7_i10;
  wire signed [`W-1:0] sb7_i11;
  wire signed [`W-1:0] sb7_i12;
  wire signed [`W-1:0] sb7_v;
  wire signed [`W-1:0] pipeUNK28_i0;
  wire signed [`W-1:0] pipeUNK28_i1;
  wire signed [`W-1:0] pipeUNK28_v;
  wire signed [`W-1:0] Pout0_i0;
  wire signed [`W-1:0] Pout0_i1;
  wire signed [`W-1:0] Pout0_i2;
  wire signed [`W-1:0] Pout0_v;
  wire signed [`W-1:0] n1570_i0;
  wire signed [`W-1:0] n1570_i1;
  wire signed [`W-1:0] n1570_v;
  wire signed [`W-1:0] n681_i0;
  wire signed [`W-1:0] n681_i1;
  wire signed [`W-1:0] n681_i2;
  wire signed [`W-1:0] n681_i3;
  wire signed [`W-1:0] n681_i4;
  wire signed [`W-1:0] n681_i5;
  wire signed [`W-1:0] n681_i6;
  wire signed [`W-1:0] n681_v;
  wire signed [`W-1:0] ir3_i0;
  wire signed [`W-1:0] ir3_i1;
  wire signed [`W-1:0] ir3_i2;
  wire signed [`W-1:0] ir3_i3;
  wire signed [`W-1:0] ir3_i4;
  wire signed [`W-1:0] ir3_i5;
  wire signed [`W-1:0] ir3_i6;
  wire signed [`W-1:0] ir3_i7;
  wire signed [`W-1:0] ir3_i8;
  wire signed [`W-1:0] ir3_i9;
  wire signed [`W-1:0] ir3_i10;
  wire signed [`W-1:0] ir3_i11;
  wire signed [`W-1:0] ir3_i12;
  wire signed [`W-1:0] ir3_i13;
  wire signed [`W-1:0] ir3_i14;
  wire signed [`W-1:0] ir3_i15;
  wire signed [`W-1:0] ir3_i16;
  wire signed [`W-1:0] ir3_i17;
  wire signed [`W-1:0] ir3_i18;
  wire signed [`W-1:0] ir3_i19;
  wire signed [`W-1:0] ir3_i20;
  wire signed [`W-1:0] ir3_i21;
  wire signed [`W-1:0] ir3_i22;
  wire signed [`W-1:0] ir3_i23;
  wire signed [`W-1:0] ir3_i24;
  wire signed [`W-1:0] ir3_i25;
  wire signed [`W-1:0] ir3_i26;
  wire signed [`W-1:0] ir3_i27;
  wire signed [`W-1:0] ir3_i28;
  wire signed [`W-1:0] ir3_i29;
  wire signed [`W-1:0] ir3_i30;
  wire signed [`W-1:0] ir3_i31;
  wire signed [`W-1:0] ir3_i32;
  wire signed [`W-1:0] ir3_i33;
  wire signed [`W-1:0] ir3_i34;
  wire signed [`W-1:0] ir3_i35;
  wire signed [`W-1:0] ir3_i36;
  wire signed [`W-1:0] ir3_i37;
  wire signed [`W-1:0] ir3_i38;
  wire signed [`W-1:0] ir3_i39;
  wire signed [`W-1:0] ir3_i40;
  wire signed [`W-1:0] ir3_i41;
  wire signed [`W-1:0] ir3_v;
  wire signed [`W-1:0] n1575_i0;
  wire signed [`W-1:0] n1575_i1;
  wire signed [`W-1:0] n1575_i2;
  wire signed [`W-1:0] n1575_i3;
  wire signed [`W-1:0] n1575_v;
  wire signed [`W-1:0] op_T0_tsx_i0;
  wire signed [`W-1:0] op_T0_tsx_i1;
  wire signed [`W-1:0] op_T0_tsx_i2;
  wire signed [`W-1:0] op_T0_tsx_v;
  wire signed [`W-1:0] n458_i0;
  wire signed [`W-1:0] n458_i1;
  wire signed [`W-1:0] n458_i2;
  wire signed [`W-1:0] n458_v;
  wire signed [`W-1:0] pcl5_i0;
  wire signed [`W-1:0] pcl5_i1;
  wire signed [`W-1:0] pcl5_i2;
  wire signed [`W-1:0] pcl5_v;
  wire signed [`W-1:0] n621_i0;
  wire signed [`W-1:0] n621_i1;
  wire signed [`W-1:0] n621_v;
  wire signed [`W-1:0] notdor4_i0;
  wire signed [`W-1:0] notdor4_i1;
  wire signed [`W-1:0] notdor4_v;
  wire signed [`W-1:0] n1224_i0;
  wire signed [`W-1:0] n1224_i1;
  wire signed [`W-1:0] n1224_i2;
  wire signed [`W-1:0] n1224_v;
  wire signed [`W-1:0] p1_i0;
  wire signed [`W-1:0] p1_i1;
  wire signed [`W-1:0] p1_v;
  wire signed [`W-1:0] n1222_i0;
  wire signed [`W-1:0] n1222_i1;
  wire signed [`W-1:0] n1222_i2;
  wire signed [`W-1:0] n1222_v;
  wire signed [`W-1:0] n1221_i0;
  wire signed [`W-1:0] n1221_i1;
  wire signed [`W-1:0] n1221_v;
  wire signed [`W-1:0] n624_i0;
  wire signed [`W-1:0] n624_i1;
  wire signed [`W-1:0] n624_i2;
  wire signed [`W-1:0] n624_v;
  wire signed [`W-1:0] n1371_i0;
  wire signed [`W-1:0] n1371_i1;
  wire signed [`W-1:0] n1371_i2;
  wire signed [`W-1:0] n1371_v;
  wire signed [`W-1:0] Pout7_i0;
  wire signed [`W-1:0] Pout7_i1;
  wire signed [`W-1:0] Pout7_i2;
  wire signed [`W-1:0] Pout7_v;
  wire signed [`W-1:0] n404_i0;
  wire signed [`W-1:0] n404_i1;
  wire signed [`W-1:0] n404_i2;
  wire signed [`W-1:0] n404_i3;
  wire signed [`W-1:0] n404_i4;
  wire signed [`W-1:0] n404_v;
  wire signed [`W-1:0] n1375_i0;
  wire signed [`W-1:0] n1375_i1;
  wire signed [`W-1:0] n1375_i2;
  wire signed [`W-1:0] n1375_v;
  wire signed [`W-1:0] n1374_i0;
  wire signed [`W-1:0] n1374_i1;
  wire signed [`W-1:0] n1374_i2;
  wire signed [`W-1:0] n1374_i3;
  wire signed [`W-1:0] n1374_v;
  wire signed [`W-1:0] alu0_i0;
  wire signed [`W-1:0] alu0_i1;
  wire signed [`W-1:0] alu0_i2;
  wire signed [`W-1:0] alu0_i3;
  wire signed [`W-1:0] alu0_v;
  wire signed [`W-1:0] ab1_i0;
  wire signed [`W-1:0] ab1_i1;
  wire signed [`W-1:0] ab1_i2;
  wire signed [`W-1:0] ab1_v;
  wire signed [`W-1:0] n1379_i0;
  wire signed [`W-1:0] n1379_i1;
  wire signed [`W-1:0] n1379_i2;
  wire signed [`W-1:0] n1379_v;
  wire signed [`W-1:0] n409_i0;
  wire signed [`W-1:0] n409_i1;
  wire signed [`W-1:0] n409_i2;
  wire signed [`W-1:0] n409_i3;
  wire signed [`W-1:0] n409_v;
  wire signed [`W-1:0] n408_i0;
  wire signed [`W-1:0] n408_i1;
  wire signed [`W-1:0] n408_v;
  wire signed [`W-1:0] n453_i0;
  wire signed [`W-1:0] n453_i1;
  wire signed [`W-1:0] n453_i2;
  wire signed [`W-1:0] n453_i3;
  wire signed [`W-1:0] n453_v;
  wire signed [`W-1:0] n1344_i0;
  wire signed [`W-1:0] n1344_i1;
  wire signed [`W-1:0] n1344_i2;
  wire signed [`W-1:0] n1344_i3;
  wire signed [`W-1:0] n1344_i4;
  wire signed [`W-1:0] n1344_v;
  wire signed [`W-1:0] n1345_i0;
  wire signed [`W-1:0] n1345_i1;
  wire signed [`W-1:0] n1345_i2;
  wire signed [`W-1:0] n1345_i3;
  wire signed [`W-1:0] n1345_i4;
  wire signed [`W-1:0] n1345_v;
  wire signed [`W-1:0] n1346_i0;
  wire signed [`W-1:0] n1346_i1;
  wire signed [`W-1:0] n1346_i2;
  wire signed [`W-1:0] n1346_i3;
  wire signed [`W-1:0] n1346_v;
  wire signed [`W-1:0] n1347_i0;
  wire signed [`W-1:0] n1347_i1;
  wire signed [`W-1:0] n1347_i2;
  wire signed [`W-1:0] n1347_v;
  wire signed [`W-1:0] n1245_i0;
  wire signed [`W-1:0] n1245_i1;
  wire signed [`W-1:0] n1245_i2;
  wire signed [`W-1:0] n1245_v;
  wire signed [`W-1:0] dpc36_IPC_i0;
  wire signed [`W-1:0] dpc36_IPC_i1;
  wire signed [`W-1:0] dpc36_IPC_i2;
  wire signed [`W-1:0] dpc36_IPC_i3;
  wire signed [`W-1:0] dpc36_IPC_i4;
  wire signed [`W-1:0] dpc36_IPC_v;
  wire signed [`W-1:0] n378_i0;
  wire signed [`W-1:0] n378_i1;
  wire signed [`W-1:0] n378_i2;
  wire signed [`W-1:0] n378_i3;
  wire signed [`W-1:0] n378_v;
  wire signed [`W-1:0] __AxBxC_0_i0;
  wire signed [`W-1:0] __AxBxC_0_i1;
  wire signed [`W-1:0] __AxBxC_0_i2;
  wire signed [`W-1:0] __AxBxC_0_v;
  wire signed [`W-1:0] op_T5_brk_i0;
  wire signed [`W-1:0] op_T5_brk_i1;
  wire signed [`W-1:0] op_T5_brk_i2;
  wire signed [`W-1:0] op_T5_brk_i3;
  wire signed [`W-1:0] op_T5_brk_v;
  wire signed [`W-1:0] n373_i0;
  wire signed [`W-1:0] n373_i1;
  wire signed [`W-1:0] n373_i2;
  wire signed [`W-1:0] n373_v;
  wire signed [`W-1:0] n372_i0;
  wire signed [`W-1:0] n372_i1;
  wire signed [`W-1:0] n372_i2;
  wire signed [`W-1:0] n372_v;
  wire signed [`W-1:0] n374_i0;
  wire signed [`W-1:0] n374_i1;
  wire signed [`W-1:0] n374_i2;
  wire signed [`W-1:0] n374_v;
  wire signed [`W-1:0] pcl6_i0;
  wire signed [`W-1:0] pcl6_i1;
  wire signed [`W-1:0] pcl6_i2;
  wire signed [`W-1:0] pcl6_v;
  wire signed [`W-1:0] abl1_i0;
  wire signed [`W-1:0] abl1_i1;
  wire signed [`W-1:0] abl1_i2;
  wire signed [`W-1:0] abl1_i3;
  wire signed [`W-1:0] abl1_i4;
  wire signed [`W-1:0] abl1_v;
  wire signed [`W-1:0] n393_i0;
  wire signed [`W-1:0] n393_i1;
  wire signed [`W-1:0] n393_v;
  wire signed [`W-1:0] n392_i0;
  wire signed [`W-1:0] n392_i1;
  wire signed [`W-1:0] n392_i2;
  wire signed [`W-1:0] n392_i3;
  wire signed [`W-1:0] n392_v;
  wire signed [`W-1:0] idl7_i0;
  wire signed [`W-1:0] idl7_i1;
  wire signed [`W-1:0] idl7_i2;
  wire signed [`W-1:0] idl7_v;
  wire signed [`W-1:0] n390_i0;
  wire signed [`W-1:0] n390_i1;
  wire signed [`W-1:0] n390_i2;
  wire signed [`W-1:0] n390_v;
  wire signed [`W-1:0] n397_i0;
  wire signed [`W-1:0] n397_i1;
  wire signed [`W-1:0] n397_i2;
  wire signed [`W-1:0] n397_v;
  wire signed [`W-1:0] n396_i0;
  wire signed [`W-1:0] n396_i1;
  wire signed [`W-1:0] n396_i2;
  wire signed [`W-1:0] n396_v;
  wire signed [`W-1:0] notalu0_i0;
  wire signed [`W-1:0] notalu0_i1;
  wire signed [`W-1:0] notalu0_v;
  wire signed [`W-1:0] ab11_i0;
  wire signed [`W-1:0] ab11_i1;
  wire signed [`W-1:0] ab11_i2;
  wire signed [`W-1:0] ab11_v;
  wire signed [`W-1:0] n398_i0;
  wire signed [`W-1:0] n398_i1;
  wire signed [`W-1:0] n398_v;
  wire signed [`W-1:0] notir6_i0;
  wire signed [`W-1:0] notir6_i1;
  wire signed [`W-1:0] notir6_i2;
  wire signed [`W-1:0] notir6_i3;
  wire signed [`W-1:0] notir6_i4;
  wire signed [`W-1:0] notir6_i5;
  wire signed [`W-1:0] notir6_i6;
  wire signed [`W-1:0] notir6_i7;
  wire signed [`W-1:0] notir6_i8;
  wire signed [`W-1:0] notir6_i9;
  wire signed [`W-1:0] notir6_i10;
  wire signed [`W-1:0] notir6_i11;
  wire signed [`W-1:0] notir6_i12;
  wire signed [`W-1:0] notir6_i13;
  wire signed [`W-1:0] notir6_i14;
  wire signed [`W-1:0] notir6_i15;
  wire signed [`W-1:0] notir6_i16;
  wire signed [`W-1:0] notir6_i17;
  wire signed [`W-1:0] notir6_i18;
  wire signed [`W-1:0] notir6_i19;
  wire signed [`W-1:0] notir6_i20;
  wire signed [`W-1:0] notir6_i21;
  wire signed [`W-1:0] notir6_i22;
  wire signed [`W-1:0] notir6_i23;
  wire signed [`W-1:0] notir6_i24;
  wire signed [`W-1:0] notir6_i25;
  wire signed [`W-1:0] notir6_i26;
  wire signed [`W-1:0] notir6_i27;
  wire signed [`W-1:0] notir6_i28;
  wire signed [`W-1:0] notir6_i29;
  wire signed [`W-1:0] notir6_i30;
  wire signed [`W-1:0] notir6_i31;
  wire signed [`W-1:0] notir6_i32;
  wire signed [`W-1:0] notir6_i33;
  wire signed [`W-1:0] notir6_i34;
  wire signed [`W-1:0] notir6_i35;
  wire signed [`W-1:0] notir6_i36;
  wire signed [`W-1:0] notir6_i37;
  wire signed [`W-1:0] notir6_i38;
  wire signed [`W-1:0] notir6_i39;
  wire signed [`W-1:0] notir6_v;
  wire signed [`W-1:0] op_shift_right_i0;
  wire signed [`W-1:0] op_shift_right_i1;
  wire signed [`W-1:0] op_shift_right_i2;
  wire signed [`W-1:0] op_shift_right_v;
  wire signed [`W-1:0] op_T0_txs_i0;
  wire signed [`W-1:0] op_T0_txs_i1;
  wire signed [`W-1:0] op_T0_txs_i2;
  wire signed [`W-1:0] op_T0_txs_i3;
  wire signed [`W-1:0] op_T0_txs_v;
  wire signed [`W-1:0] op_ror_i0;
  wire signed [`W-1:0] op_ror_i1;
  wire signed [`W-1:0] op_ror_i2;
  wire signed [`W-1:0] op_ror_v;
  wire signed [`W-1:0] dpc33_PCHDB_i0;
  wire signed [`W-1:0] dpc33_PCHDB_i1;
  wire signed [`W-1:0] dpc33_PCHDB_i2;
  wire signed [`W-1:0] dpc33_PCHDB_i3;
  wire signed [`W-1:0] dpc33_PCHDB_i4;
  wire signed [`W-1:0] dpc33_PCHDB_i5;
  wire signed [`W-1:0] dpc33_PCHDB_i6;
  wire signed [`W-1:0] dpc33_PCHDB_i7;
  wire signed [`W-1:0] dpc33_PCHDB_i8;
  wire signed [`W-1:0] dpc33_PCHDB_i9;
  wire signed [`W-1:0] dpc33_PCHDB_v;
  wire signed [`W-1:0] n241_i0;
  wire signed [`W-1:0] n241_i1;
  wire signed [`W-1:0] n241_i2;
  wire signed [`W-1:0] n241_i3;
  wire signed [`W-1:0] n241_v;
  wire signed [`W-1:0] idl5_i0;
  wire signed [`W-1:0] idl5_i1;
  wire signed [`W-1:0] idl5_i2;
  wire signed [`W-1:0] idl5_v;
  wire signed [`W-1:0] n243_i0;
  wire signed [`W-1:0] n243_i1;
  wire signed [`W-1:0] n243_i2;
  wire signed [`W-1:0] n243_v;
  wire signed [`W-1:0] n242_i0;
  wire signed [`W-1:0] n242_i1;
  wire signed [`W-1:0] n242_i2;
  wire signed [`W-1:0] n242_i3;
  wire signed [`W-1:0] n242_v;
  wire signed [`W-1:0] n249_i0;
  wire signed [`W-1:0] n249_i1;
  wire signed [`W-1:0] n249_i2;
  wire signed [`W-1:0] n249_i3;
  wire signed [`W-1:0] n249_v;
  wire signed [`W-1:0] notRdy0_i0;
  wire signed [`W-1:0] notRdy0_i1;
  wire signed [`W-1:0] notRdy0_i2;
  wire signed [`W-1:0] notRdy0_i3;
  wire signed [`W-1:0] notRdy0_i4;
  wire signed [`W-1:0] notRdy0_i5;
  wire signed [`W-1:0] notRdy0_i6;
  wire signed [`W-1:0] notRdy0_i7;
  wire signed [`W-1:0] notRdy0_i8;
  wire signed [`W-1:0] notRdy0_i9;
  wire signed [`W-1:0] notRdy0_i10;
  wire signed [`W-1:0] notRdy0_i11;
  wire signed [`W-1:0] notRdy0_i12;
  wire signed [`W-1:0] notRdy0_i13;
  wire signed [`W-1:0] notRdy0_i14;
  wire signed [`W-1:0] notRdy0_i15;
  wire signed [`W-1:0] notRdy0_i16;
  wire signed [`W-1:0] notRdy0_i17;
  wire signed [`W-1:0] notRdy0_i18;
  wire signed [`W-1:0] notRdy0_i19;
  wire signed [`W-1:0] notRdy0_i20;
  wire signed [`W-1:0] notRdy0_i21;
  wire signed [`W-1:0] notRdy0_i22;
  wire signed [`W-1:0] notRdy0_i23;
  wire signed [`W-1:0] notRdy0_i24;
  wire signed [`W-1:0] notRdy0_i25;
  wire signed [`W-1:0] notRdy0_i26;
  wire signed [`W-1:0] notRdy0_i27;
  wire signed [`W-1:0] notRdy0_i28;
  wire signed [`W-1:0] notRdy0_i29;
  wire signed [`W-1:0] notRdy0_i30;
  wire signed [`W-1:0] notRdy0_i31;
  wire signed [`W-1:0] notRdy0_i32;
  wire signed [`W-1:0] notRdy0_i33;
  wire signed [`W-1:0] notRdy0_i34;
  wire signed [`W-1:0] notRdy0_i35;
  wire signed [`W-1:0] notRdy0_i36;
  wire signed [`W-1:0] notRdy0_v;
  wire signed [`W-1:0] op_T0_txa_i0;
  wire signed [`W-1:0] op_T0_txa_i1;
  wire signed [`W-1:0] op_T0_txa_i2;
  wire signed [`W-1:0] op_T0_txa_v;
  wire signed [`W-1:0] abl7_i0;
  wire signed [`W-1:0] abl7_i1;
  wire signed [`W-1:0] abl7_i2;
  wire signed [`W-1:0] abl7_i3;
  wire signed [`W-1:0] abl7_i4;
  wire signed [`W-1:0] abl7_v;
  wire signed [`W-1:0] n177_i0;
  wire signed [`W-1:0] n177_i1;
  wire signed [`W-1:0] n177_i2;
  wire signed [`W-1:0] n177_v;
  wire signed [`W-1:0] n176_i0;
  wire signed [`W-1:0] n176_i1;
  wire signed [`W-1:0] n176_i2;
  wire signed [`W-1:0] n176_v;
  wire signed [`W-1:0] db5_i0;
  wire signed [`W-1:0] db5_i1;
  wire signed [`W-1:0] db5_i2;
  wire signed [`W-1:0] db5_i3;
  wire signed [`W-1:0] db5_i4;
  wire signed [`W-1:0] db5_v;
  wire signed [`W-1:0] _AxB_6__C56_i0;
  wire signed [`W-1:0] _AxB_6__C56_i1;
  wire signed [`W-1:0] _AxB_6__C56_i2;
  wire signed [`W-1:0] _AxB_6__C56_v;
  wire signed [`W-1:0] n172_i0;
  wire signed [`W-1:0] n172_i1;
  wire signed [`W-1:0] n172_i2;
  wire signed [`W-1:0] n172_i3;
  wire signed [`W-1:0] n172_v;
  wire signed [`W-1:0] n171_i0;
  wire signed [`W-1:0] n171_i1;
  wire signed [`W-1:0] n171_i2;
  wire signed [`W-1:0] n171_i3;
  wire signed [`W-1:0] n171_v;
  wire signed [`W-1:0] pipeVectorA1_i0;
  wire signed [`W-1:0] pipeVectorA1_i1;
  wire signed [`W-1:0] pipeVectorA1_v;
  wire signed [`W-1:0] abl2_i0;
  wire signed [`W-1:0] abl2_i1;
  wire signed [`W-1:0] abl2_i2;
  wire signed [`W-1:0] abl2_i3;
  wire signed [`W-1:0] abl2_i4;
  wire signed [`W-1:0] abl2_v;
  wire signed [`W-1:0] n1500_i0;
  wire signed [`W-1:0] n1500_i1;
  wire signed [`W-1:0] n1500_i2;
  wire signed [`W-1:0] n1500_v;
  wire signed [`W-1:0] pcl2_i0;
  wire signed [`W-1:0] pcl2_i1;
  wire signed [`W-1:0] pcl2_i2;
  wire signed [`W-1:0] pcl2_v;
  wire signed [`W-1:0] n652_i0;
  wire signed [`W-1:0] n652_i1;
  wire signed [`W-1:0] n652_i2;
  wire signed [`W-1:0] n652_i3;
  wire signed [`W-1:0] n652_i4;
  wire signed [`W-1:0] n652_v;
  wire signed [`W-1:0] n1507_i0;
  wire signed [`W-1:0] n1507_i1;
  wire signed [`W-1:0] n1507_i2;
  wire signed [`W-1:0] n1507_v;
  wire signed [`W-1:0] op_T0_and_i0;
  wire signed [`W-1:0] op_T0_and_i1;
  wire signed [`W-1:0] op_T0_and_i2;
  wire signed [`W-1:0] op_T0_and_v;
  wire signed [`W-1:0] n1505_i0;
  wire signed [`W-1:0] n1505_i1;
  wire signed [`W-1:0] n1505_v;
  wire signed [`W-1:0] n1364_i0;
  wire signed [`W-1:0] n1364_i1;
  wire signed [`W-1:0] n1364_i2;
  wire signed [`W-1:0] n1364_i3;
  wire signed [`W-1:0] n1364_v;
  wire signed [`W-1:0] n659_i0;
  wire signed [`W-1:0] n659_i1;
  wire signed [`W-1:0] n659_i2;
  wire signed [`W-1:0] n659_i3;
  wire signed [`W-1:0] n659_v;
  wire signed [`W-1:0] n1115_i0;
  wire signed [`W-1:0] n1115_i1;
  wire signed [`W-1:0] n1115_i2;
  wire signed [`W-1:0] n1115_v;
  wire signed [`W-1:0] n1618_i0;
  wire signed [`W-1:0] n1618_i1;
  wire signed [`W-1:0] n1618_i2;
  wire signed [`W-1:0] n1618_i3;
  wire signed [`W-1:0] n1618_i4;
  wire signed [`W-1:0] n1618_v;
  wire signed [`W-1:0] n1619_i0;
  wire signed [`W-1:0] n1619_i1;
  wire signed [`W-1:0] n1619_i2;
  wire signed [`W-1:0] n1619_v;
  wire signed [`W-1:0] n1614_i0;
  wire signed [`W-1:0] n1614_i1;
  wire signed [`W-1:0] n1614_i2;
  wire signed [`W-1:0] n1614_v;
  wire signed [`W-1:0] op_T4_rts_i0;
  wire signed [`W-1:0] op_T4_rts_i1;
  wire signed [`W-1:0] op_T4_rts_i2;
  wire signed [`W-1:0] op_T4_rts_v;
  wire signed [`W-1:0] n1613_i0;
  wire signed [`W-1:0] n1613_i1;
  wire signed [`W-1:0] n1613_i2;
  wire signed [`W-1:0] n1613_i3;
  wire signed [`W-1:0] n1613_v;
  wire signed [`W-1:0] n1610_i0;
  wire signed [`W-1:0] n1610_i1;
  wire signed [`W-1:0] n1610_i2;
  wire signed [`W-1:0] n1610_v;
  wire signed [`W-1:0] pcl7_i0;
  wire signed [`W-1:0] pcl7_i1;
  wire signed [`W-1:0] pcl7_i2;
  wire signed [`W-1:0] pcl7_v;
  wire signed [`W-1:0] op_T0_clc_sec_i0;
  wire signed [`W-1:0] op_T0_clc_sec_i1;
  wire signed [`W-1:0] op_T0_clc_sec_i2;
  wire signed [`W-1:0] op_T0_clc_sec_v;
  wire signed [`W-1:0] alua4_i0;
  wire signed [`W-1:0] alua4_i1;
  wire signed [`W-1:0] alua4_i2;
  wire signed [`W-1:0] alua4_i3;
  wire signed [`W-1:0] alua4_v;
  wire signed [`W-1:0] abh4_i0;
  wire signed [`W-1:0] abh4_i1;
  wire signed [`W-1:0] abh4_i2;
  wire signed [`W-1:0] abh4_i3;
  wire signed [`W-1:0] abh4_i4;
  wire signed [`W-1:0] abh4_v;
  wire signed [`W-1:0] n1140_i0;
  wire signed [`W-1:0] n1140_i1;
  wire signed [`W-1:0] n1140_i2;
  wire signed [`W-1:0] n1140_v;
  wire signed [`W-1:0] n1141_i0;
  wire signed [`W-1:0] n1141_i1;
  wire signed [`W-1:0] n1141_i2;
  wire signed [`W-1:0] n1141_v;
  wire signed [`W-1:0] alucout_i0;
  wire signed [`W-1:0] alucout_i1;
  wire signed [`W-1:0] alucout_i2;
  wire signed [`W-1:0] alucout_i3;
  wire signed [`W-1:0] alucout_v;
  wire signed [`W-1:0] n1147_i0;
  wire signed [`W-1:0] n1147_i1;
  wire signed [`W-1:0] n1147_i2;
  wire signed [`W-1:0] n1147_i3;
  wire signed [`W-1:0] n1147_v;
  wire signed [`W-1:0] DA_C45_i0;
  wire signed [`W-1:0] DA_C45_i1;
  wire signed [`W-1:0] DA_C45_i2;
  wire signed [`W-1:0] DA_C45_i3;
  wire signed [`W-1:0] DA_C45_v;
  wire signed [`W-1:0] n1145_i0;
  wire signed [`W-1:0] n1145_i1;
  wire signed [`W-1:0] n1145_i2;
  wire signed [`W-1:0] n1145_v;
  wire signed [`W-1:0] y1_i0;
  wire signed [`W-1:0] y1_i1;
  wire signed [`W-1:0] y1_i2;
  wire signed [`W-1:0] y1_v;
  wire signed [`W-1:0] n1149_i0;
  wire signed [`W-1:0] n1149_i1;
  wire signed [`W-1:0] n1149_v;
  wire signed [`W-1:0] n692_i0;
  wire signed [`W-1:0] n692_i1;
  wire signed [`W-1:0] n692_i2;
  wire signed [`W-1:0] n692_i3;
  wire signed [`W-1:0] n692_v;
  wire signed [`W-1:0] BRtaken_i0;
  wire signed [`W-1:0] BRtaken_i1;
  wire signed [`W-1:0] BRtaken_i2;
  wire signed [`W-1:0] BRtaken_i3;
  wire signed [`W-1:0] BRtaken_v;
  wire signed [`W-1:0] op_asl_rol_i0;
  wire signed [`W-1:0] op_asl_rol_i1;
  wire signed [`W-1:0] op_asl_rol_i2;
  wire signed [`W-1:0] op_asl_rol_i3;
  wire signed [`W-1:0] op_asl_rol_v;
  wire signed [`W-1:0] n696_i0;
  wire signed [`W-1:0] n696_i1;
  wire signed [`W-1:0] n696_i2;
  wire signed [`W-1:0] n696_v;
  wire signed [`W-1:0] notalu1_i0;
  wire signed [`W-1:0] notalu1_i1;
  wire signed [`W-1:0] notalu1_v;
  wire signed [`W-1:0] n694_i0;
  wire signed [`W-1:0] n694_i1;
  wire signed [`W-1:0] n694_i2;
  wire signed [`W-1:0] n694_i3;
  wire signed [`W-1:0] n694_i4;
  wire signed [`W-1:0] n694_v;
  wire signed [`W-1:0] n1541_i0;
  wire signed [`W-1:0] n1541_i1;
  wire signed [`W-1:0] n1541_i2;
  wire signed [`W-1:0] n1541_i3;
  wire signed [`W-1:0] n1541_v;
  wire signed [`W-1:0] n698_i0;
  wire signed [`W-1:0] n698_i1;
  wire signed [`W-1:0] n698_v;
  wire signed [`W-1:0] _DA_ADD2_i0;
  wire signed [`W-1:0] _DA_ADD2_i1;
  wire signed [`W-1:0] _DA_ADD2_i2;
  wire signed [`W-1:0] _DA_ADD2_i3;
  wire signed [`W-1:0] _DA_ADD2_v;
  wire signed [`W-1:0] n1548_i0;
  wire signed [`W-1:0] n1548_i1;
  wire signed [`W-1:0] n1548_i2;
  wire signed [`W-1:0] n1548_v;
  wire signed [`W-1:0] n1549_i0;
  wire signed [`W-1:0] n1549_i1;
  wire signed [`W-1:0] n1549_i2;
  wire signed [`W-1:0] n1549_v;
  wire signed [`W-1:0] n543_i0;
  wire signed [`W-1:0] n543_i1;
  wire signed [`W-1:0] n543_i2;
  wire signed [`W-1:0] n543_i3;
  wire signed [`W-1:0] n543_v;
  wire signed [`W-1:0] pd4_clearIR_i0;
  wire signed [`W-1:0] pd4_clearIR_i1;
  wire signed [`W-1:0] pd4_clearIR_i2;
  wire signed [`W-1:0] pd4_clearIR_i3;
  wire signed [`W-1:0] pd4_clearIR_i4;
  wire signed [`W-1:0] pd4_clearIR_i5;
  wire signed [`W-1:0] pd4_clearIR_v;
  wire signed [`W-1:0] n541_i0;
  wire signed [`W-1:0] n541_i1;
  wire signed [`W-1:0] n541_i2;
  wire signed [`W-1:0] n541_v;
  wire signed [`W-1:0] op_shift_i0;
  wire signed [`W-1:0] op_shift_i1;
  wire signed [`W-1:0] op_shift_i2;
  wire signed [`W-1:0] op_shift_v;
  wire signed [`W-1:0] n544_i0;
  wire signed [`W-1:0] n544_i1;
  wire signed [`W-1:0] n544_i2;
  wire signed [`W-1:0] n544_v;
  wire signed [`W-1:0] n548_i0;
  wire signed [`W-1:0] n548_i1;
  wire signed [`W-1:0] n548_i2;
  wire signed [`W-1:0] n548_v;
  wire signed [`W-1:0] dpc11_SBADD_i0;
  wire signed [`W-1:0] dpc11_SBADD_i1;
  wire signed [`W-1:0] dpc11_SBADD_i2;
  wire signed [`W-1:0] dpc11_SBADD_i3;
  wire signed [`W-1:0] dpc11_SBADD_i4;
  wire signed [`W-1:0] dpc11_SBADD_i5;
  wire signed [`W-1:0] dpc11_SBADD_i6;
  wire signed [`W-1:0] dpc11_SBADD_i7;
  wire signed [`W-1:0] dpc11_SBADD_i8;
  wire signed [`W-1:0] dpc11_SBADD_i9;
  wire signed [`W-1:0] dpc11_SBADD_v;
  wire signed [`W-1:0] n761_i0;
  wire signed [`W-1:0] n761_i1;
  wire signed [`W-1:0] n761_i2;
  wire signed [`W-1:0] n761_i3;
  wire signed [`W-1:0] n761_i4;
  wire signed [`W-1:0] n761_i5;
  wire signed [`W-1:0] n761_v;
  wire signed [`W-1:0] dpc40_ADLPCL_i0;
  wire signed [`W-1:0] dpc40_ADLPCL_i1;
  wire signed [`W-1:0] dpc40_ADLPCL_i2;
  wire signed [`W-1:0] dpc40_ADLPCL_i3;
  wire signed [`W-1:0] dpc40_ADLPCL_i4;
  wire signed [`W-1:0] dpc40_ADLPCL_i5;
  wire signed [`W-1:0] dpc40_ADLPCL_i6;
  wire signed [`W-1:0] dpc40_ADLPCL_i7;
  wire signed [`W-1:0] dpc40_ADLPCL_i8;
  wire signed [`W-1:0] dpc40_ADLPCL_i9;
  wire signed [`W-1:0] dpc40_ADLPCL_v;
  wire signed [`W-1:0] n415_i0;
  wire signed [`W-1:0] n415_i1;
  wire signed [`W-1:0] n415_v;
  wire signed [`W-1:0] n417_i0;
  wire signed [`W-1:0] n417_i1;
  wire signed [`W-1:0] n417_i2;
  wire signed [`W-1:0] n417_v;
  wire signed [`W-1:0] n1389_i0;
  wire signed [`W-1:0] n1389_i1;
  wire signed [`W-1:0] n1389_i2;
  wire signed [`W-1:0] n1389_i3;
  wire signed [`W-1:0] n1389_i4;
  wire signed [`W-1:0] n1389_v;
  wire signed [`W-1:0] notalucout_i0;
  wire signed [`W-1:0] notalucout_i1;
  wire signed [`W-1:0] notalucout_i2;
  wire signed [`W-1:0] notalucout_i3;
  wire signed [`W-1:0] notalucout_v;
  wire signed [`W-1:0] adl0_i0;
  wire signed [`W-1:0] adl0_i1;
  wire signed [`W-1:0] adl0_i2;
  wire signed [`W-1:0] adl0_i3;
  wire signed [`W-1:0] adl0_i4;
  wire signed [`W-1:0] adl0_i5;
  wire signed [`W-1:0] adl0_i6;
  wire signed [`W-1:0] adl0_i7;
  wire signed [`W-1:0] adl0_i8;
  wire signed [`W-1:0] adl0_v;
  wire signed [`W-1:0] ir2_i0;
  wire signed [`W-1:0] ir2_i1;
  wire signed [`W-1:0] ir2_i2;
  wire signed [`W-1:0] ir2_i3;
  wire signed [`W-1:0] ir2_i4;
  wire signed [`W-1:0] ir2_i5;
  wire signed [`W-1:0] ir2_i6;
  wire signed [`W-1:0] ir2_i7;
  wire signed [`W-1:0] ir2_i8;
  wire signed [`W-1:0] ir2_i9;
  wire signed [`W-1:0] ir2_i10;
  wire signed [`W-1:0] ir2_i11;
  wire signed [`W-1:0] ir2_i12;
  wire signed [`W-1:0] ir2_i13;
  wire signed [`W-1:0] ir2_i14;
  wire signed [`W-1:0] ir2_i15;
  wire signed [`W-1:0] ir2_i16;
  wire signed [`W-1:0] ir2_i17;
  wire signed [`W-1:0] ir2_i18;
  wire signed [`W-1:0] ir2_i19;
  wire signed [`W-1:0] ir2_i20;
  wire signed [`W-1:0] ir2_i21;
  wire signed [`W-1:0] ir2_i22;
  wire signed [`W-1:0] ir2_i23;
  wire signed [`W-1:0] ir2_i24;
  wire signed [`W-1:0] ir2_i25;
  wire signed [`W-1:0] ir2_i26;
  wire signed [`W-1:0] ir2_i27;
  wire signed [`W-1:0] ir2_i28;
  wire signed [`W-1:0] ir2_i29;
  wire signed [`W-1:0] ir2_i30;
  wire signed [`W-1:0] ir2_i31;
  wire signed [`W-1:0] ir2_i32;
  wire signed [`W-1:0] ir2_i33;
  wire signed [`W-1:0] ir2_i34;
  wire signed [`W-1:0] ir2_i35;
  wire signed [`W-1:0] ir2_i36;
  wire signed [`W-1:0] ir2_i37;
  wire signed [`W-1:0] ir2_i38;
  wire signed [`W-1:0] ir2_i39;
  wire signed [`W-1:0] ir2_i40;
  wire signed [`W-1:0] ir2_i41;
  wire signed [`W-1:0] ir2_i42;
  wire signed [`W-1:0] ir2_i43;
  wire signed [`W-1:0] ir2_i44;
  wire signed [`W-1:0] ir2_i45;
  wire signed [`W-1:0] ir2_i46;
  wire signed [`W-1:0] ir2_i47;
  wire signed [`W-1:0] ir2_i48;
  wire signed [`W-1:0] ir2_i49;
  wire signed [`W-1:0] ir2_i50;
  wire signed [`W-1:0] ir2_i51;
  wire signed [`W-1:0] ir2_i52;
  wire signed [`W-1:0] ir2_i53;
  wire signed [`W-1:0] ir2_i54;
  wire signed [`W-1:0] ir2_i55;
  wire signed [`W-1:0] ir2_i56;
  wire signed [`W-1:0] ir2_i57;
  wire signed [`W-1:0] ir2_i58;
  wire signed [`W-1:0] ir2_i59;
  wire signed [`W-1:0] ir2_i60;
  wire signed [`W-1:0] ir2_i61;
  wire signed [`W-1:0] ir2_i62;
  wire signed [`W-1:0] ir2_i63;
  wire signed [`W-1:0] ir2_i64;
  wire signed [`W-1:0] ir2_i65;
  wire signed [`W-1:0] ir2_i66;
  wire signed [`W-1:0] ir2_i67;
  wire signed [`W-1:0] ir2_i68;
  wire signed [`W-1:0] ir2_i69;
  wire signed [`W-1:0] ir2_i70;
  wire signed [`W-1:0] ir2_i71;
  wire signed [`W-1:0] ir2_i72;
  wire signed [`W-1:0] ir2_v;
  wire signed [`W-1:0] op_T5_mem_ind_idx_i0;
  wire signed [`W-1:0] op_T5_mem_ind_idx_i1;
  wire signed [`W-1:0] op_T5_mem_ind_idx_i2;
  wire signed [`W-1:0] op_T5_mem_ind_idx_v;
  wire signed [`W-1:0] n1386_i0;
  wire signed [`W-1:0] n1386_i1;
  wire signed [`W-1:0] n1386_i2;
  wire signed [`W-1:0] n1386_v;
  wire signed [`W-1:0] n1387_i0;
  wire signed [`W-1:0] n1387_i1;
  wire signed [`W-1:0] n1387_i2;
  wire signed [`W-1:0] n1387_i3;
  wire signed [`W-1:0] n1387_v;
  wire signed [`W-1:0] n1380_i0;
  wire signed [`W-1:0] n1380_i1;
  wire signed [`W-1:0] n1380_i2;
  wire signed [`W-1:0] n1380_i3;
  wire signed [`W-1:0] n1380_v;
  wire signed [`W-1:0] op_T3_jmp_i0;
  wire signed [`W-1:0] op_T3_jmp_i1;
  wire signed [`W-1:0] op_T3_jmp_i2;
  wire signed [`W-1:0] op_T3_jmp_v;
  wire signed [`W-1:0] brk_done_i0;
  wire signed [`W-1:0] brk_done_i1;
  wire signed [`W-1:0] brk_done_i2;
  wire signed [`W-1:0] brk_done_i3;
  wire signed [`W-1:0] brk_done_i4;
  wire signed [`W-1:0] brk_done_i5;
  wire signed [`W-1:0] brk_done_i6;
  wire signed [`W-1:0] brk_done_i7;
  wire signed [`W-1:0] brk_done_i8;
  wire signed [`W-1:0] brk_done_v;
  wire signed [`W-1:0] n1383_i0;
  wire signed [`W-1:0] n1383_i1;
  wire signed [`W-1:0] n1383_i2;
  wire signed [`W-1:0] n1383_v;
  wire signed [`W-1:0] n368_i0;
  wire signed [`W-1:0] n368_i1;
  wire signed [`W-1:0] n368_i2;
  wire signed [`W-1:0] n368_v;
  wire signed [`W-1:0] pd4_i0;
  wire signed [`W-1:0] pd4_i1;
  wire signed [`W-1:0] pd4_v;
  wire signed [`W-1:0] n366_i0;
  wire signed [`W-1:0] n366_i1;
  wire signed [`W-1:0] n366_i2;
  wire signed [`W-1:0] n366_v;
  wire signed [`W-1:0] _ABL4_i0;
  wire signed [`W-1:0] _ABL4_i1;
  wire signed [`W-1:0] _ABL4_i2;
  wire signed [`W-1:0] _ABL4_v;
  wire signed [`W-1:0] PD_0xx0xx0x_i0;
  wire signed [`W-1:0] PD_0xx0xx0x_i1;
  wire signed [`W-1:0] PD_0xx0xx0x_i2;
  wire signed [`W-1:0] PD_0xx0xx0x_v;
  wire signed [`W-1:0] dpc14_SRS_i0;
  wire signed [`W-1:0] dpc14_SRS_i1;
  wire signed [`W-1:0] dpc14_SRS_i2;
  wire signed [`W-1:0] dpc14_SRS_i3;
  wire signed [`W-1:0] dpc14_SRS_i4;
  wire signed [`W-1:0] dpc14_SRS_i5;
  wire signed [`W-1:0] dpc14_SRS_i6;
  wire signed [`W-1:0] dpc14_SRS_i7;
  wire signed [`W-1:0] dpc14_SRS_i8;
  wire signed [`W-1:0] dpc14_SRS_i9;
  wire signed [`W-1:0] dpc14_SRS_v;
  wire signed [`W-1:0] n360_i0;
  wire signed [`W-1:0] n360_i1;
  wire signed [`W-1:0] n360_v;
  wire signed [`W-1:0] pd1_i0;
  wire signed [`W-1:0] pd1_i1;
  wire signed [`W-1:0] pd1_v;
  wire signed [`W-1:0] n381_i0;
  wire signed [`W-1:0] n381_i1;
  wire signed [`W-1:0] n381_i2;
  wire signed [`W-1:0] n381_i3;
  wire signed [`W-1:0] n381_v;
  wire signed [`W-1:0] op_T0_iny_dey_i0;
  wire signed [`W-1:0] op_T0_iny_dey_i1;
  wire signed [`W-1:0] op_T0_iny_dey_i2;
  wire signed [`W-1:0] op_T0_iny_dey_v;
  wire signed [`W-1:0] n383_i0;
  wire signed [`W-1:0] n383_i1;
  wire signed [`W-1:0] n383_i2;
  wire signed [`W-1:0] n383_i3;
  wire signed [`W-1:0] n383_v;
  wire signed [`W-1:0] n384_i0;
  wire signed [`W-1:0] n384_i1;
  wire signed [`W-1:0] n384_i2;
  wire signed [`W-1:0] n384_i3;
  wire signed [`W-1:0] n384_v;
  wire signed [`W-1:0] n385_i0;
  wire signed [`W-1:0] n385_i1;
  wire signed [`W-1:0] n385_i2;
  wire signed [`W-1:0] n385_v;
  wire signed [`W-1:0] n386_i0;
  wire signed [`W-1:0] n386_i1;
  wire signed [`W-1:0] n386_i2;
  wire signed [`W-1:0] n386_i3;
  wire signed [`W-1:0] n386_v;
  wire signed [`W-1:0] n388_i0;
  wire signed [`W-1:0] n388_i1;
  wire signed [`W-1:0] n388_i2;
  wire signed [`W-1:0] n388_v;
  wire signed [`W-1:0] n389_i0;
  wire signed [`W-1:0] n389_i1;
  wire signed [`W-1:0] n389_i2;
  wire signed [`W-1:0] n389_i3;
  wire signed [`W-1:0] n389_i4;
  wire signed [`W-1:0] n389_v;
  wire signed [`W-1:0] op_T2_idx_x_xy_i0;
  wire signed [`W-1:0] op_T2_idx_x_xy_i1;
  wire signed [`W-1:0] op_T2_idx_x_xy_i2;
  wire signed [`W-1:0] op_T2_idx_x_xy_i3;
  wire signed [`W-1:0] op_T2_idx_x_xy_v;
  wire signed [`W-1:0] op_jsr_i0;
  wire signed [`W-1:0] op_jsr_i1;
  wire signed [`W-1:0] op_jsr_i2;
  wire signed [`W-1:0] op_jsr_v;
  wire signed [`W-1:0] _op_set_C_i0;
  wire signed [`W-1:0] _op_set_C_i1;
  wire signed [`W-1:0] _op_set_C_i2;
  wire signed [`W-1:0] _op_set_C_v;
  wire signed [`W-1:0] n253_i0;
  wire signed [`W-1:0] n253_i1;
  wire signed [`W-1:0] n253_i2;
  wire signed [`W-1:0] n253_i3;
  wire signed [`W-1:0] n253_v;
  wire signed [`W-1:0] notaluoutmux1_i0;
  wire signed [`W-1:0] notaluoutmux1_i1;
  wire signed [`W-1:0] notaluoutmux1_i2;
  wire signed [`W-1:0] notaluoutmux1_i3;
  wire signed [`W-1:0] notaluoutmux1_i4;
  wire signed [`W-1:0] notaluoutmux1_i5;
  wire signed [`W-1:0] notaluoutmux1_v;
  wire signed [`W-1:0] n251_i0;
  wire signed [`W-1:0] n251_i1;
  wire signed [`W-1:0] n251_i2;
  wire signed [`W-1:0] n251_i3;
  wire signed [`W-1:0] n251_v;
  wire signed [`W-1:0] n256_i0;
  wire signed [`W-1:0] n256_i1;
  wire signed [`W-1:0] n256_i2;
  wire signed [`W-1:0] n256_v;
  wire signed [`W-1:0] op_T0_tya_i0;
  wire signed [`W-1:0] op_T0_tya_i1;
  wire signed [`W-1:0] op_T0_tya_i2;
  wire signed [`W-1:0] op_T0_tya_v;
  wire signed [`W-1:0] n254_i0;
  wire signed [`W-1:0] n254_i1;
  wire signed [`W-1:0] n254_i2;
  wire signed [`W-1:0] n254_v;
  wire signed [`W-1:0] n255_i0;
  wire signed [`W-1:0] n255_i1;
  wire signed [`W-1:0] n255_i2;
  wire signed [`W-1:0] n255_v;
  wire signed [`W-1:0] n168_i0;
  wire signed [`W-1:0] n168_i1;
  wire signed [`W-1:0] n168_i2;
  wire signed [`W-1:0] n168_v;
  wire signed [`W-1:0] n169_i0;
  wire signed [`W-1:0] n169_i1;
  wire signed [`W-1:0] n169_i2;
  wire signed [`W-1:0] n169_v;
  wire signed [`W-1:0] DC78_phi2_i0;
  wire signed [`W-1:0] DC78_phi2_i1;
  wire signed [`W-1:0] DC78_phi2_v;
  wire signed [`W-1:0] sb5_i0;
  wire signed [`W-1:0] sb5_i1;
  wire signed [`W-1:0] sb5_i2;
  wire signed [`W-1:0] sb5_i3;
  wire signed [`W-1:0] sb5_i4;
  wire signed [`W-1:0] sb5_i5;
  wire signed [`W-1:0] sb5_i6;
  wire signed [`W-1:0] sb5_i7;
  wire signed [`W-1:0] sb5_i8;
  wire signed [`W-1:0] sb5_i9;
  wire signed [`W-1:0] sb5_i10;
  wire signed [`W-1:0] sb5_i11;
  wire signed [`W-1:0] sb5_i12;
  wire signed [`W-1:0] sb5_v;
  wire signed [`W-1:0] op_T0_tax_i0;
  wire signed [`W-1:0] op_T0_tax_i1;
  wire signed [`W-1:0] op_T0_tax_i2;
  wire signed [`W-1:0] op_T0_tax_v;
  wire signed [`W-1:0] n160_i0;
  wire signed [`W-1:0] n160_i1;
  wire signed [`W-1:0] n160_i2;
  wire signed [`W-1:0] n160_v;
  wire signed [`W-1:0] n161_i0;
  wire signed [`W-1:0] n161_i1;
  wire signed [`W-1:0] n161_i2;
  wire signed [`W-1:0] n161_i3;
  wire signed [`W-1:0] n161_v;
  wire signed [`W-1:0] a3_i0;
  wire signed [`W-1:0] a3_i1;
  wire signed [`W-1:0] a3_i2;
  wire signed [`W-1:0] a3_v;
  wire signed [`W-1:0] n163_i0;
  wire signed [`W-1:0] n163_i1;
  wire signed [`W-1:0] n163_i2;
  wire signed [`W-1:0] n163_i3;
  wire signed [`W-1:0] n163_v;
  wire signed [`W-1:0] n1090_i0;
  wire signed [`W-1:0] n1090_i1;
  wire signed [`W-1:0] n1090_i2;
  wire signed [`W-1:0] n1090_v;
  wire signed [`W-1:0] dasb6_i0;
  wire signed [`W-1:0] dasb6_i1;
  wire signed [`W-1:0] dasb6_i2;
  wire signed [`W-1:0] dasb6_v;
  wire signed [`W-1:0] n1093_i0;
  wire signed [`W-1:0] n1093_i1;
  wire signed [`W-1:0] n1093_i2;
  wire signed [`W-1:0] n1093_v;
  wire signed [`W-1:0] s5_i0;
  wire signed [`W-1:0] s5_i1;
  wire signed [`W-1:0] s5_i2;
  wire signed [`W-1:0] s5_v;
  wire signed [`W-1:0] n1099_i0;
  wire signed [`W-1:0] n1099_i1;
  wire signed [`W-1:0] n1099_i2;
  wire signed [`W-1:0] n1099_v;
  wire signed [`W-1:0] n1609_i0;
  wire signed [`W-1:0] n1609_i1;
  wire signed [`W-1:0] n1609_i2;
  wire signed [`W-1:0] n1609_v;
  wire signed [`W-1:0] n1608_i0;
  wire signed [`W-1:0] n1608_i1;
  wire signed [`W-1:0] n1608_i2;
  wire signed [`W-1:0] n1608_v;
  wire signed [`W-1:0] op_sty_cpy_mem_i0;
  wire signed [`W-1:0] op_sty_cpy_mem_i1;
  wire signed [`W-1:0] op_sty_cpy_mem_i2;
  wire signed [`W-1:0] op_sty_cpy_mem_i3;
  wire signed [`W-1:0] op_sty_cpy_mem_v;
  wire signed [`W-1:0] n1600_i0;
  wire signed [`W-1:0] n1600_i1;
  wire signed [`W-1:0] n1600_i2;
  wire signed [`W-1:0] n1600_v;
  wire signed [`W-1:0] nots4_i0;
  wire signed [`W-1:0] nots4_i1;
  wire signed [`W-1:0] nots4_v;
  wire signed [`W-1:0] n1602_i0;
  wire signed [`W-1:0] n1602_i1;
  wire signed [`W-1:0] n1602_v;
  wire signed [`W-1:0] n1605_i0;
  wire signed [`W-1:0] n1605_i1;
  wire signed [`W-1:0] n1605_i2;
  wire signed [`W-1:0] n1605_i3;
  wire signed [`W-1:0] n1605_v;
  wire signed [`W-1:0] pipeUNK14_i0;
  wire signed [`W-1:0] pipeUNK14_i1;
  wire signed [`W-1:0] pipeUNK14_v;
  wire signed [`W-1:0] n1606_i0;
  wire signed [`W-1:0] n1606_i1;
  wire signed [`W-1:0] n1606_v;
  wire signed [`W-1:0] pd1_clearIR_i0;
  wire signed [`W-1:0] pd1_clearIR_i1;
  wire signed [`W-1:0] pd1_clearIR_i2;
  wire signed [`W-1:0] pd1_clearIR_i3;
  wire signed [`W-1:0] pd1_clearIR_v;
  wire signed [`W-1:0] alurawcout_i0;
  wire signed [`W-1:0] alurawcout_i1;
  wire signed [`W-1:0] alurawcout_i2;
  wire signed [`W-1:0] alurawcout_v;
  wire signed [`W-1:0] n803_i0;
  wire signed [`W-1:0] n803_i1;
  wire signed [`W-1:0] n803_i2;
  wire signed [`W-1:0] n803_v;
  wire signed [`W-1:0] dpc0_YSB_i0;
  wire signed [`W-1:0] dpc0_YSB_i1;
  wire signed [`W-1:0] dpc0_YSB_i2;
  wire signed [`W-1:0] dpc0_YSB_i3;
  wire signed [`W-1:0] dpc0_YSB_i4;
  wire signed [`W-1:0] dpc0_YSB_i5;
  wire signed [`W-1:0] dpc0_YSB_i6;
  wire signed [`W-1:0] dpc0_YSB_i7;
  wire signed [`W-1:0] dpc0_YSB_i8;
  wire signed [`W-1:0] dpc0_YSB_i9;
  wire signed [`W-1:0] dpc0_YSB_v;
  wire signed [`W-1:0] n800_i0;
  wire signed [`W-1:0] n800_i1;
  wire signed [`W-1:0] n800_i2;
  wire signed [`W-1:0] n800_v;
  wire signed [`W-1:0] n807_i0;
  wire signed [`W-1:0] n807_i1;
  wire signed [`W-1:0] n807_i2;
  wire signed [`W-1:0] n807_v;
  wire signed [`W-1:0] n806_v;
  wire signed [`W-1:0] n805_i0;
  wire signed [`W-1:0] n805_i1;
  wire signed [`W-1:0] n805_v;
  wire signed [`W-1:0] op_T4_brk_jsr_i0;
  wire signed [`W-1:0] op_T4_brk_jsr_i1;
  wire signed [`W-1:0] op_T4_brk_jsr_i2;
  wire signed [`W-1:0] op_T4_brk_jsr_v;
  wire signed [`W-1:0] n1159_i0;
  wire signed [`W-1:0] n1159_i1;
  wire signed [`W-1:0] n1159_i2;
  wire signed [`W-1:0] n1159_v;
  wire signed [`W-1:0] x_op_T__adc_sbc_i0;
  wire signed [`W-1:0] x_op_T__adc_sbc_i1;
  wire signed [`W-1:0] x_op_T__adc_sbc_i2;
  wire signed [`W-1:0] x_op_T__adc_sbc_i3;
  wire signed [`W-1:0] x_op_T__adc_sbc_v;
  wire signed [`W-1:0] n1154_i0;
  wire signed [`W-1:0] n1154_i1;
  wire signed [`W-1:0] n1154_i2;
  wire signed [`W-1:0] n1154_v;
  wire signed [`W-1:0] n1157_i0;
  wire signed [`W-1:0] n1157_i1;
  wire signed [`W-1:0] n1157_i2;
  wire signed [`W-1:0] n1157_v;
  wire signed [`W-1:0] rw_i0;
  wire signed [`W-1:0] rw_i1;
  wire signed [`W-1:0] rw_i2;
  wire signed [`W-1:0] rw_v;
  wire signed [`W-1:0] sb1_i0;
  wire signed [`W-1:0] sb1_i1;
  wire signed [`W-1:0] sb1_i2;
  wire signed [`W-1:0] sb1_i3;
  wire signed [`W-1:0] sb1_i4;
  wire signed [`W-1:0] sb1_i5;
  wire signed [`W-1:0] sb1_i6;
  wire signed [`W-1:0] sb1_i7;
  wire signed [`W-1:0] sb1_i8;
  wire signed [`W-1:0] sb1_i9;
  wire signed [`W-1:0] sb1_i10;
  wire signed [`W-1:0] sb1_i11;
  wire signed [`W-1:0] sb1_i12;
  wire signed [`W-1:0] sb1_v;
  wire signed [`W-1:0] n1153_i0;
  wire signed [`W-1:0] n1153_i1;
  wire signed [`W-1:0] n1153_i2;
  wire signed [`W-1:0] n1153_i3;
  wire signed [`W-1:0] n1153_v;
  wire signed [`W-1:0] n1152_i0;
  wire signed [`W-1:0] n1152_i1;
  wire signed [`W-1:0] n1152_i2;
  wire signed [`W-1:0] n1152_v;
  wire signed [`W-1:0] dpc13_ORS_i0;
  wire signed [`W-1:0] dpc13_ORS_i1;
  wire signed [`W-1:0] dpc13_ORS_i2;
  wire signed [`W-1:0] dpc13_ORS_i3;
  wire signed [`W-1:0] dpc13_ORS_i4;
  wire signed [`W-1:0] dpc13_ORS_i5;
  wire signed [`W-1:0] dpc13_ORS_i6;
  wire signed [`W-1:0] dpc13_ORS_i7;
  wire signed [`W-1:0] dpc13_ORS_i8;
  wire signed [`W-1:0] dpc13_ORS_i9;
  wire signed [`W-1:0] dpc13_ORS_v;
  wire signed [`W-1:0] pch6_i0;
  wire signed [`W-1:0] pch6_i1;
  wire signed [`W-1:0] pch6_i2;
  wire signed [`W-1:0] pch6_v;
  wire signed [`W-1:0] p2_i0;
  wire signed [`W-1:0] p2_i1;
  wire signed [`W-1:0] p2_v;
  wire signed [`W-1:0] n1552_i0;
  wire signed [`W-1:0] n1552_i1;
  wire signed [`W-1:0] n1552_i2;
  wire signed [`W-1:0] n1552_v;
  wire signed [`W-1:0] op_T3_abs_idx_i0;
  wire signed [`W-1:0] op_T3_abs_idx_i1;
  wire signed [`W-1:0] op_T3_abs_idx_i2;
  wire signed [`W-1:0] op_T3_abs_idx_v;
  wire signed [`W-1:0] op_brk_rti_i0;
  wire signed [`W-1:0] op_brk_rti_i1;
  wire signed [`W-1:0] op_brk_rti_i2;
  wire signed [`W-1:0] op_brk_rti_v;
  wire signed [`W-1:0] pipeUNK34_i0;
  wire signed [`W-1:0] pipeUNK34_i1;
  wire signed [`W-1:0] pipeUNK34_v;
  wire signed [`W-1:0] n50_i0;
  wire signed [`W-1:0] n50_i1;
  wire signed [`W-1:0] n50_v;
  wire signed [`W-1:0] op_lsr_ror_dec_inc_i0;
  wire signed [`W-1:0] op_lsr_ror_dec_inc_i1;
  wire signed [`W-1:0] op_lsr_ror_dec_inc_i2;
  wire signed [`W-1:0] op_lsr_ror_dec_inc_v;
  wire signed [`W-1:0] adh1_i0;
  wire signed [`W-1:0] adh1_i1;
  wire signed [`W-1:0] adh1_i2;
  wire signed [`W-1:0] adh1_i3;
  wire signed [`W-1:0] adh1_i4;
  wire signed [`W-1:0] adh1_i5;
  wire signed [`W-1:0] adh1_i6;
  wire signed [`W-1:0] adh1_v;
  wire signed [`W-1:0] pipeT_SYNC_i0;
  wire signed [`W-1:0] pipeT_SYNC_i1;
  wire signed [`W-1:0] pipeT_SYNC_v;
  wire signed [`W-1:0] pclp7_i0;
  wire signed [`W-1:0] pclp7_i1;
  wire signed [`W-1:0] pclp7_v;
  wire signed [`W-1:0] pchp7_i0;
  wire signed [`W-1:0] pchp7_i1;
  wire signed [`W-1:0] pchp7_i2;
  wire signed [`W-1:0] pchp7_v;
  wire signed [`W-1:0] dpc23_SBAC_i0;
  wire signed [`W-1:0] dpc23_SBAC_i1;
  wire signed [`W-1:0] dpc23_SBAC_i2;
  wire signed [`W-1:0] dpc23_SBAC_i3;
  wire signed [`W-1:0] dpc23_SBAC_i4;
  wire signed [`W-1:0] dpc23_SBAC_i5;
  wire signed [`W-1:0] dpc23_SBAC_i6;
  wire signed [`W-1:0] dpc23_SBAC_i7;
  wire signed [`W-1:0] dpc23_SBAC_i8;
  wire signed [`W-1:0] dpc23_SBAC_i9;
  wire signed [`W-1:0] dpc23_SBAC_v;
  wire signed [`W-1:0] n533_i0;
  wire signed [`W-1:0] n533_i1;
  wire signed [`W-1:0] n533_i2;
  wire signed [`W-1:0] n533_v;
  wire signed [`W-1:0] __AxBxC_7_i0;
  wire signed [`W-1:0] __AxBxC_7_i1;
  wire signed [`W-1:0] __AxBxC_7_i2;
  wire signed [`W-1:0] __AxBxC_7_v;
  wire signed [`W-1:0] n531_i0;
  wire signed [`W-1:0] n531_i1;
  wire signed [`W-1:0] n531_i2;
  wire signed [`W-1:0] n531_i3;
  wire signed [`W-1:0] n531_v;
  wire signed [`W-1:0] dasb0_i0;
  wire signed [`W-1:0] dasb0_i1;
  wire signed [`W-1:0] dasb0_i2;
  wire signed [`W-1:0] dasb0_i3;
  wire signed [`W-1:0] dasb0_i4;
  wire signed [`W-1:0] dasb0_i5;
  wire signed [`W-1:0] dasb0_i6;
  wire signed [`W-1:0] dasb0_i7;
  wire signed [`W-1:0] dasb0_i8;
  wire signed [`W-1:0] dasb0_i9;
  wire signed [`W-1:0] dasb0_i10;
  wire signed [`W-1:0] dasb0_i11;
  wire signed [`W-1:0] dasb0_i12;
  wire signed [`W-1:0] dasb0_v;
  wire signed [`W-1:0] sync_i0;
  wire signed [`W-1:0] sync_i1;
  wire signed [`W-1:0] sync_i2;
  wire signed [`W-1:0] sync_v;
  wire signed [`W-1:0] n538_i0;
  wire signed [`W-1:0] n538_i1;
  wire signed [`W-1:0] n538_i2;
  wire signed [`W-1:0] n538_v;
  wire signed [`W-1:0] _ABH7_i0;
  wire signed [`W-1:0] _ABH7_i1;
  wire signed [`W-1:0] _ABH7_i2;
  wire signed [`W-1:0] _ABH7_v;
  wire signed [`W-1:0] n428_i0;
  wire signed [`W-1:0] n428_i1;
  wire signed [`W-1:0] n428_i2;
  wire signed [`W-1:0] n428_v;
  wire signed [`W-1:0] n1399_i0;
  wire signed [`W-1:0] n1399_i1;
  wire signed [`W-1:0] n1399_i2;
  wire signed [`W-1:0] n1399_i3;
  wire signed [`W-1:0] n1399_v;
  wire signed [`W-1:0] n1398_i0;
  wire signed [`W-1:0] n1398_i1;
  wire signed [`W-1:0] n1398_i2;
  wire signed [`W-1:0] n1398_i3;
  wire signed [`W-1:0] n1398_i4;
  wire signed [`W-1:0] n1398_i5;
  wire signed [`W-1:0] n1398_v;
  wire signed [`W-1:0] op_T0_shift_a_i0;
  wire signed [`W-1:0] op_T0_shift_a_i1;
  wire signed [`W-1:0] op_T0_shift_a_i2;
  wire signed [`W-1:0] op_T0_shift_a_i3;
  wire signed [`W-1:0] op_T0_shift_a_v;
  wire signed [`W-1:0] n1395_i0;
  wire signed [`W-1:0] n1395_i1;
  wire signed [`W-1:0] n1395_v;
  wire signed [`W-1:0] notir5_i0;
  wire signed [`W-1:0] notir5_i1;
  wire signed [`W-1:0] notir5_i2;
  wire signed [`W-1:0] notir5_i3;
  wire signed [`W-1:0] notir5_i4;
  wire signed [`W-1:0] notir5_i5;
  wire signed [`W-1:0] notir5_i6;
  wire signed [`W-1:0] notir5_i7;
  wire signed [`W-1:0] notir5_i8;
  wire signed [`W-1:0] notir5_i9;
  wire signed [`W-1:0] notir5_i10;
  wire signed [`W-1:0] notir5_i11;
  wire signed [`W-1:0] notir5_i12;
  wire signed [`W-1:0] notir5_i13;
  wire signed [`W-1:0] notir5_i14;
  wire signed [`W-1:0] notir5_i15;
  wire signed [`W-1:0] notir5_i16;
  wire signed [`W-1:0] notir5_i17;
  wire signed [`W-1:0] notir5_i18;
  wire signed [`W-1:0] notir5_i19;
  wire signed [`W-1:0] notir5_i20;
  wire signed [`W-1:0] notir5_i21;
  wire signed [`W-1:0] notir5_i22;
  wire signed [`W-1:0] notir5_i23;
  wire signed [`W-1:0] notir5_i24;
  wire signed [`W-1:0] notir5_i25;
  wire signed [`W-1:0] notir5_i26;
  wire signed [`W-1:0] notir5_i27;
  wire signed [`W-1:0] notir5_i28;
  wire signed [`W-1:0] notir5_i29;
  wire signed [`W-1:0] notir5_i30;
  wire signed [`W-1:0] notir5_i31;
  wire signed [`W-1:0] notir5_i32;
  wire signed [`W-1:0] notir5_i33;
  wire signed [`W-1:0] notir5_i34;
  wire signed [`W-1:0] notir5_i35;
  wire signed [`W-1:0] notir5_i36;
  wire signed [`W-1:0] notir5_i37;
  wire signed [`W-1:0] notir5_v;
  wire signed [`W-1:0] db4_i0;
  wire signed [`W-1:0] db4_i1;
  wire signed [`W-1:0] db4_i2;
  wire signed [`W-1:0] db4_i3;
  wire signed [`W-1:0] db4_i4;
  wire signed [`W-1:0] db4_v;
  wire signed [`W-1:0] n1392_i0;
  wire signed [`W-1:0] n1392_i1;
  wire signed [`W-1:0] n1392_i2;
  wire signed [`W-1:0] n1392_i3;
  wire signed [`W-1:0] n1392_v;
  wire signed [`W-1:0] _C56_i0;
  wire signed [`W-1:0] _C56_i1;
  wire signed [`W-1:0] _C56_i2;
  wire signed [`W-1:0] _C56_i3;
  wire signed [`W-1:0] _C56_v;
  wire signed [`W-1:0] alua5_i0;
  wire signed [`W-1:0] alua5_i1;
  wire signed [`W-1:0] alua5_i2;
  wire signed [`W-1:0] alua5_i3;
  wire signed [`W-1:0] alua5_v;
  wire signed [`W-1:0] _TWOCYCLE_i0;
  wire signed [`W-1:0] _TWOCYCLE_i1;
  wire signed [`W-1:0] _TWOCYCLE_i2;
  wire signed [`W-1:0] _TWOCYCLE_v;
  wire signed [`W-1:0] n853_i0;
  wire signed [`W-1:0] n853_i1;
  wire signed [`W-1:0] n853_i2;
  wire signed [`W-1:0] n853_i3;
  wire signed [`W-1:0] n853_v;
  wire signed [`W-1:0] pipeUNK26_i0;
  wire signed [`W-1:0] pipeUNK26_i1;
  wire signed [`W-1:0] pipeUNK26_v;
  wire signed [`W-1:0] dpc28_0ADH0_i0;
  wire signed [`W-1:0] dpc28_0ADH0_i1;
  wire signed [`W-1:0] dpc28_0ADH0_i2;
  wire signed [`W-1:0] dpc28_0ADH0_v;
  wire signed [`W-1:0] n228_i0;
  wire signed [`W-1:0] n228_i1;
  wire signed [`W-1:0] n228_i2;
  wire signed [`W-1:0] n228_v;
  wire signed [`W-1:0] n227_i0;
  wire signed [`W-1:0] n227_i1;
  wire signed [`W-1:0] n227_i2;
  wire signed [`W-1:0] n227_v;
  wire signed [`W-1:0] n226_i0;
  wire signed [`W-1:0] n226_i1;
  wire signed [`W-1:0] n226_v;
  wire signed [`W-1:0] n225_i0;
  wire signed [`W-1:0] n225_i1;
  wire signed [`W-1:0] n225_i2;
  wire signed [`W-1:0] n225_v;
  wire signed [`W-1:0] n224_i0;
  wire signed [`W-1:0] n224_i1;
  wire signed [`W-1:0] n224_i2;
  wire signed [`W-1:0] n224_i3;
  wire signed [`W-1:0] n224_v;
  wire signed [`W-1:0] n223_i0;
  wire signed [`W-1:0] n223_i1;
  wire signed [`W-1:0] n223_v;
  wire signed [`W-1:0] notdor0_i0;
  wire signed [`W-1:0] notdor0_i1;
  wire signed [`W-1:0] notdor0_v;
  wire signed [`W-1:0] n221_i0;
  wire signed [`W-1:0] n221_i1;
  wire signed [`W-1:0] n221_i2;
  wire signed [`W-1:0] n221_v;
  wire signed [`W-1:0] n220_i0;
  wire signed [`W-1:0] n220_i1;
  wire signed [`W-1:0] n220_i2;
  wire signed [`W-1:0] n220_i3;
  wire signed [`W-1:0] n220_v;
  wire signed [`W-1:0] pipeUNK39_i0;
  wire signed [`W-1:0] pipeUNK39_i1;
  wire signed [`W-1:0] pipeUNK39_v;
  wire signed [`W-1:0] _ABL0_i0;
  wire signed [`W-1:0] _ABL0_i1;
  wire signed [`W-1:0] _ABL0_i2;
  wire signed [`W-1:0] _ABL0_v;
  wire signed [`W-1:0] n152_i0;
  wire signed [`W-1:0] n152_i1;
  wire signed [`W-1:0] n152_i2;
  wire signed [`W-1:0] n152_v;
  wire signed [`W-1:0] aluanorb1_i0;
  wire signed [`W-1:0] aluanorb1_i1;
  wire signed [`W-1:0] aluanorb1_i2;
  wire signed [`W-1:0] aluanorb1_i3;
  wire signed [`W-1:0] aluanorb1_i4;
  wire signed [`W-1:0] aluanorb1_v;
  wire signed [`W-1:0] n154_i0;
  wire signed [`W-1:0] n154_i1;
  wire signed [`W-1:0] n154_i2;
  wire signed [`W-1:0] n154_i3;
  wire signed [`W-1:0] n154_v;
  wire signed [`W-1:0] op_T2_stack_access_i0;
  wire signed [`W-1:0] op_T2_stack_access_i1;
  wire signed [`W-1:0] op_T2_stack_access_i2;
  wire signed [`W-1:0] op_T2_stack_access_v;
  wire signed [`W-1:0] clock2_i0;
  wire signed [`W-1:0] clock2_i1;
  wire signed [`W-1:0] clock2_i2;
  wire signed [`W-1:0] clock2_i3;
  wire signed [`W-1:0] clock2_i4;
  wire signed [`W-1:0] clock2_i5;
  wire signed [`W-1:0] clock2_i6;
  wire signed [`W-1:0] clock2_i7;
  wire signed [`W-1:0] clock2_i8;
  wire signed [`W-1:0] clock2_i9;
  wire signed [`W-1:0] clock2_i10;
  wire signed [`W-1:0] clock2_i11;
  wire signed [`W-1:0] clock2_i12;
  wire signed [`W-1:0] clock2_i13;
  wire signed [`W-1:0] clock2_v;
  wire signed [`W-1:0] res_i0;
  wire signed [`W-1:0] res_i1;
  wire signed [`W-1:0] res_v;
  wire signed [`W-1:0] notdor7_i0;
  wire signed [`W-1:0] notdor7_i1;
  wire signed [`W-1:0] notdor7_v;
  wire signed [`W-1:0] n1293_i0;
  wire signed [`W-1:0] n1293_i1;
  wire signed [`W-1:0] n1293_i2;
  wire signed [`W-1:0] n1293_v;
  wire signed [`W-1:0] n1256_i0;
  wire signed [`W-1:0] n1256_i1;
  wire signed [`W-1:0] n1256_i2;
  wire signed [`W-1:0] n1256_v;
  wire signed [`W-1:0] t4_i0;
  wire signed [`W-1:0] t4_i1;
  wire signed [`W-1:0] t4_i2;
  wire signed [`W-1:0] t4_i3;
  wire signed [`W-1:0] t4_i4;
  wire signed [`W-1:0] t4_i5;
  wire signed [`W-1:0] t4_i6;
  wire signed [`W-1:0] t4_i7;
  wire signed [`W-1:0] t4_i8;
  wire signed [`W-1:0] t4_i9;
  wire signed [`W-1:0] t4_i10;
  wire signed [`W-1:0] t4_i11;
  wire signed [`W-1:0] t4_i12;
  wire signed [`W-1:0] t4_i13;
  wire signed [`W-1:0] t4_v;
  wire signed [`W-1:0] __AxB_0_i0;
  wire signed [`W-1:0] __AxB_0_i1;
  wire signed [`W-1:0] __AxB_0_i2;
  wire signed [`W-1:0] __AxB_0_i3;
  wire signed [`W-1:0] __AxB_0_i4;
  wire signed [`W-1:0] __AxB_0_v;
  wire signed [`W-1:0] n1526_i0;
  wire signed [`W-1:0] n1526_i1;
  wire signed [`W-1:0] n1526_i2;
  wire signed [`W-1:0] n1526_v;
  wire signed [`W-1:0] n818_i0;
  wire signed [`W-1:0] n818_i1;
  wire signed [`W-1:0] n818_i2;
  wire signed [`W-1:0] n818_i3;
  wire signed [`W-1:0] n818_v;
  wire signed [`W-1:0] n819_i0;
  wire signed [`W-1:0] n819_i1;
  wire signed [`W-1:0] n819_i2;
  wire signed [`W-1:0] n819_i3;
  wire signed [`W-1:0] n819_v;
  wire signed [`W-1:0] n1255_i0;
  wire signed [`W-1:0] n1255_i1;
  wire signed [`W-1:0] n1255_i2;
  wire signed [`W-1:0] n1255_v;
  wire signed [`W-1:0] n810_i0;
  wire signed [`W-1:0] n810_i1;
  wire signed [`W-1:0] n810_i2;
  wire signed [`W-1:0] n810_v;
  wire signed [`W-1:0] n811_i0;
  wire signed [`W-1:0] n811_i1;
  wire signed [`W-1:0] n811_i2;
  wire signed [`W-1:0] n811_i3;
  wire signed [`W-1:0] n811_i4;
  wire signed [`W-1:0] n811_v;
  wire signed [`W-1:0] n812_i0;
  wire signed [`W-1:0] n812_i1;
  wire signed [`W-1:0] n812_i2;
  wire signed [`W-1:0] n812_v;
  wire signed [`W-1:0] n813_i0;
  wire signed [`W-1:0] n813_i1;
  wire signed [`W-1:0] n813_i2;
  wire signed [`W-1:0] n813_v;
  wire signed [`W-1:0] n815_i0;
  wire signed [`W-1:0] n815_i1;
  wire signed [`W-1:0] n815_i2;
  wire signed [`W-1:0] n815_v;
  wire signed [`W-1:0] __AxB5__C45_i0;
  wire signed [`W-1:0] __AxB5__C45_i1;
  wire signed [`W-1:0] __AxB5__C45_i2;
  wire signed [`W-1:0] __AxB5__C45_v;
  wire signed [`W-1:0] abl3_i0;
  wire signed [`W-1:0] abl3_i1;
  wire signed [`W-1:0] abl3_i2;
  wire signed [`W-1:0] abl3_i3;
  wire signed [`W-1:0] abl3_i4;
  wire signed [`W-1:0] abl3_v;
  wire signed [`W-1:0] n1251_i0;
  wire signed [`W-1:0] n1251_i1;
  wire signed [`W-1:0] n1251_i2;
  wire signed [`W-1:0] n1251_i3;
  wire signed [`W-1:0] n1251_v;
  wire signed [`W-1:0] notalu4_i0;
  wire signed [`W-1:0] notalu4_i1;
  wire signed [`W-1:0] notalu4_v;
  wire signed [`W-1:0] n1491_i0;
  wire signed [`W-1:0] n1491_i1;
  wire signed [`W-1:0] n1491_i2;
  wire signed [`W-1:0] n1491_i3;
  wire signed [`W-1:0] n1491_v;
  wire signed [`W-1:0] n1492_i0;
  wire signed [`W-1:0] n1492_i1;
  wire signed [`W-1:0] n1492_i2;
  wire signed [`W-1:0] n1492_i3;
  wire signed [`W-1:0] n1492_v;
  wire signed [`W-1:0] ab7_i0;
  wire signed [`W-1:0] ab7_i1;
  wire signed [`W-1:0] ab7_i2;
  wire signed [`W-1:0] ab7_v;
  wire signed [`W-1:0] dasb7_i0;
  wire signed [`W-1:0] dasb7_i1;
  wire signed [`W-1:0] dasb7_i2;
  wire signed [`W-1:0] dasb7_v;
  wire signed [`W-1:0] n1495_i0;
  wire signed [`W-1:0] n1495_i1;
  wire signed [`W-1:0] n1495_i2;
  wire signed [`W-1:0] n1495_v;
  wire signed [`W-1:0] n1496_i0;
  wire signed [`W-1:0] n1496_i1;
  wire signed [`W-1:0] n1496_i2;
  wire signed [`W-1:0] n1496_i3;
  wire signed [`W-1:0] n1496_i4;
  wire signed [`W-1:0] n1496_v;
  wire signed [`W-1:0] n1497_i0;
  wire signed [`W-1:0] n1497_i1;
  wire signed [`W-1:0] n1497_i2;
  wire signed [`W-1:0] n1497_v;
  wire signed [`W-1:0] n1499_i0;
  wire signed [`W-1:0] n1499_i1;
  wire signed [`W-1:0] n1499_i2;
  wire signed [`W-1:0] n1499_i3;
  wire signed [`W-1:0] n1499_v;
  wire signed [`W-1:0] n423_i0;
  wire signed [`W-1:0] n423_i1;
  wire signed [`W-1:0] n423_i2;
  wire signed [`W-1:0] n423_v;
  wire signed [`W-1:0] dpc4_SSB_i0;
  wire signed [`W-1:0] dpc4_SSB_i1;
  wire signed [`W-1:0] dpc4_SSB_i2;
  wire signed [`W-1:0] dpc4_SSB_i3;
  wire signed [`W-1:0] dpc4_SSB_i4;
  wire signed [`W-1:0] dpc4_SSB_i5;
  wire signed [`W-1:0] dpc4_SSB_i6;
  wire signed [`W-1:0] dpc4_SSB_i7;
  wire signed [`W-1:0] dpc4_SSB_i8;
  wire signed [`W-1:0] dpc4_SSB_i9;
  wire signed [`W-1:0] dpc4_SSB_v;
  wire signed [`W-1:0] s4_i0;
  wire signed [`W-1:0] s4_i1;
  wire signed [`W-1:0] s4_i2;
  wire signed [`W-1:0] s4_v;
  wire signed [`W-1:0] dpc34_PCLC_i0;
  wire signed [`W-1:0] dpc34_PCLC_i1;
  wire signed [`W-1:0] dpc34_PCLC_i2;
  wire signed [`W-1:0] dpc34_PCLC_i3;
  wire signed [`W-1:0] dpc34_PCLC_i4;
  wire signed [`W-1:0] dpc34_PCLC_v;
  wire signed [`W-1:0] n1705_i0;
  wire signed [`W-1:0] n1705_i1;
  wire signed [`W-1:0] n1705_i2;
  wire signed [`W-1:0] n1705_v;
  wire signed [`W-1:0] n1708_i0;
  wire signed [`W-1:0] n1708_i1;
  wire signed [`W-1:0] n1708_i2;
  wire signed [`W-1:0] n1708_i3;
  wire signed [`W-1:0] n1708_i4;
  wire signed [`W-1:0] n1708_v;
  wire signed [`W-1:0] n1709_i0;
  wire signed [`W-1:0] n1709_i1;
  wire signed [`W-1:0] n1709_i2;
  wire signed [`W-1:0] n1709_i3;
  wire signed [`W-1:0] n1709_v;
  wire signed [`W-1:0] n424_i0;
  wire signed [`W-1:0] n424_i1;
  wire signed [`W-1:0] n424_i2;
  wire signed [`W-1:0] n424_v;
  wire signed [`W-1:0] n1391_i0;
  wire signed [`W-1:0] n1391_i1;
  wire signed [`W-1:0] n1391_i2;
  wire signed [`W-1:0] n1391_v;
  wire signed [`W-1:0] _ABH5_i0;
  wire signed [`W-1:0] _ABH5_i1;
  wire signed [`W-1:0] _ABH5_i2;
  wire signed [`W-1:0] _ABH5_v;
  wire signed [`W-1:0] n1129_i0;
  wire signed [`W-1:0] n1129_i1;
  wire signed [`W-1:0] n1129_i2;
  wire signed [`W-1:0] n1129_i3;
  wire signed [`W-1:0] n1129_v;
  wire signed [`W-1:0] n1120_i0;
  wire signed [`W-1:0] n1120_i1;
  wire signed [`W-1:0] n1120_i2;
  wire signed [`W-1:0] n1120_v;
  wire signed [`W-1:0] n1121_i0;
  wire signed [`W-1:0] n1121_i1;
  wire signed [`W-1:0] n1121_v;
  wire signed [`W-1:0] _C12_i0;
  wire signed [`W-1:0] _C12_i1;
  wire signed [`W-1:0] _C12_i2;
  wire signed [`W-1:0] _C12_i3;
  wire signed [`W-1:0] _C12_v;
  wire signed [`W-1:0] notalu7_i0;
  wire signed [`W-1:0] notalu7_i1;
  wire signed [`W-1:0] notalu7_v;
  wire signed [`W-1:0] n1124_i0;
  wire signed [`W-1:0] n1124_i1;
  wire signed [`W-1:0] n1124_v;
  wire signed [`W-1:0] notir3_i0;
  wire signed [`W-1:0] notir3_i1;
  wire signed [`W-1:0] notir3_i2;
  wire signed [`W-1:0] notir3_i3;
  wire signed [`W-1:0] notir3_i4;
  wire signed [`W-1:0] notir3_i5;
  wire signed [`W-1:0] notir3_i6;
  wire signed [`W-1:0] notir3_i7;
  wire signed [`W-1:0] notir3_i8;
  wire signed [`W-1:0] notir3_i9;
  wire signed [`W-1:0] notir3_i10;
  wire signed [`W-1:0] notir3_i11;
  wire signed [`W-1:0] notir3_i12;
  wire signed [`W-1:0] notir3_i13;
  wire signed [`W-1:0] notir3_i14;
  wire signed [`W-1:0] notir3_i15;
  wire signed [`W-1:0] notir3_i16;
  wire signed [`W-1:0] notir3_i17;
  wire signed [`W-1:0] notir3_i18;
  wire signed [`W-1:0] notir3_i19;
  wire signed [`W-1:0] notir3_i20;
  wire signed [`W-1:0] notir3_i21;
  wire signed [`W-1:0] notir3_i22;
  wire signed [`W-1:0] notir3_i23;
  wire signed [`W-1:0] notir3_i24;
  wire signed [`W-1:0] notir3_i25;
  wire signed [`W-1:0] notir3_i26;
  wire signed [`W-1:0] notir3_i27;
  wire signed [`W-1:0] notir3_i28;
  wire signed [`W-1:0] notir3_i29;
  wire signed [`W-1:0] notir3_i30;
  wire signed [`W-1:0] notir3_i31;
  wire signed [`W-1:0] notir3_i32;
  wire signed [`W-1:0] notir3_i33;
  wire signed [`W-1:0] notir3_i34;
  wire signed [`W-1:0] notir3_i35;
  wire signed [`W-1:0] notir3_i36;
  wire signed [`W-1:0] notir3_i37;
  wire signed [`W-1:0] notir3_i38;
  wire signed [`W-1:0] notir3_i39;
  wire signed [`W-1:0] notir3_i40;
  wire signed [`W-1:0] notir3_i41;
  wire signed [`W-1:0] notir3_i42;
  wire signed [`W-1:0] notir3_i43;
  wire signed [`W-1:0] notir3_i44;
  wire signed [`W-1:0] notir3_i45;
  wire signed [`W-1:0] notir3_i46;
  wire signed [`W-1:0] notir3_i47;
  wire signed [`W-1:0] notir3_i48;
  wire signed [`W-1:0] notir3_i49;
  wire signed [`W-1:0] notir3_i50;
  wire signed [`W-1:0] notir3_i51;
  wire signed [`W-1:0] notir3_v;
  wire signed [`W-1:0] n1126_i0;
  wire signed [`W-1:0] n1126_i1;
  wire signed [`W-1:0] n1126_v;
  wire signed [`W-1:0] n525_i0;
  wire signed [`W-1:0] n525_i1;
  wire signed [`W-1:0] n525_i2;
  wire signed [`W-1:0] n525_i3;
  wire signed [`W-1:0] n525_v;
  wire signed [`W-1:0] n526_i0;
  wire signed [`W-1:0] n526_i1;
  wire signed [`W-1:0] n526_v;
  wire signed [`W-1:0] notdor1_i0;
  wire signed [`W-1:0] notdor1_i1;
  wire signed [`W-1:0] notdor1_v;
  wire signed [`W-1:0] n520_i0;
  wire signed [`W-1:0] n520_i1;
  wire signed [`W-1:0] n520_i2;
  wire signed [`W-1:0] n520_v;
  wire signed [`W-1:0] n521_i0;
  wire signed [`W-1:0] n521_i1;
  wire signed [`W-1:0] n521_v;
  wire signed [`W-1:0] op_ORS_i0;
  wire signed [`W-1:0] op_ORS_i1;
  wire signed [`W-1:0] op_ORS_i2;
  wire signed [`W-1:0] op_ORS_i3;
  wire signed [`W-1:0] op_ORS_v;
  wire signed [`W-1:0] n523_i0;
  wire signed [`W-1:0] n523_i1;
  wire signed [`W-1:0] n523_i2;
  wire signed [`W-1:0] n523_i3;
  wire signed [`W-1:0] n523_i4;
  wire signed [`W-1:0] n523_v;
  wire signed [`W-1:0] n1014_i0;
  wire signed [`W-1:0] n1014_i1;
  wire signed [`W-1:0] n1014_i2;
  wire signed [`W-1:0] n1014_i3;
  wire signed [`W-1:0] n1014_v;
  wire signed [`W-1:0] dpc21_ADDADL_i0;
  wire signed [`W-1:0] dpc21_ADDADL_i1;
  wire signed [`W-1:0] dpc21_ADDADL_i2;
  wire signed [`W-1:0] dpc21_ADDADL_i3;
  wire signed [`W-1:0] dpc21_ADDADL_i4;
  wire signed [`W-1:0] dpc21_ADDADL_i5;
  wire signed [`W-1:0] dpc21_ADDADL_i6;
  wire signed [`W-1:0] dpc21_ADDADL_i7;
  wire signed [`W-1:0] dpc21_ADDADL_i8;
  wire signed [`W-1:0] dpc21_ADDADL_i9;
  wire signed [`W-1:0] dpc21_ADDADL_v;
  wire signed [`W-1:0] n1016_i0;
  wire signed [`W-1:0] n1016_i1;
  wire signed [`W-1:0] n1016_i2;
  wire signed [`W-1:0] n1016_v;
  wire signed [`W-1:0] n1017_i0;
  wire signed [`W-1:0] n1017_i1;
  wire signed [`W-1:0] n1017_i2;
  wire signed [`W-1:0] n1017_v;
  wire signed [`W-1:0] n1010_i0;
  wire signed [`W-1:0] n1010_i1;
  wire signed [`W-1:0] n1010_i2;
  wire signed [`W-1:0] n1010_i3;
  wire signed [`W-1:0] n1010_v;
  wire signed [`W-1:0] pipeUNK11_i0;
  wire signed [`W-1:0] pipeUNK11_i1;
  wire signed [`W-1:0] pipeUNK11_v;
  wire signed [`W-1:0] a1_i0;
  wire signed [`W-1:0] a1_i1;
  wire signed [`W-1:0] a1_i2;
  wire signed [`W-1:0] a1_v;
  wire signed [`W-1:0] dpc32_PCHADH_i0;
  wire signed [`W-1:0] dpc32_PCHADH_i1;
  wire signed [`W-1:0] dpc32_PCHADH_i2;
  wire signed [`W-1:0] dpc32_PCHADH_i3;
  wire signed [`W-1:0] dpc32_PCHADH_i4;
  wire signed [`W-1:0] dpc32_PCHADH_i5;
  wire signed [`W-1:0] dpc32_PCHADH_i6;
  wire signed [`W-1:0] dpc32_PCHADH_i7;
  wire signed [`W-1:0] dpc32_PCHADH_i8;
  wire signed [`W-1:0] dpc32_PCHADH_i9;
  wire signed [`W-1:0] dpc32_PCHADH_v;
  wire signed [`W-1:0] A_B5_i0;
  wire signed [`W-1:0] A_B5_i1;
  wire signed [`W-1:0] A_B5_i2;
  wire signed [`W-1:0] A_B5_v;
  wire signed [`W-1:0] ab12_i0;
  wire signed [`W-1:0] ab12_i1;
  wire signed [`W-1:0] ab12_i2;
  wire signed [`W-1:0] ab12_v;
  wire signed [`W-1:0] n1230_i0;
  wire signed [`W-1:0] n1230_i1;
  wire signed [`W-1:0] n1230_i2;
  wire signed [`W-1:0] n1230_i3;
  wire signed [`W-1:0] n1230_v;
  wire signed [`W-1:0] n1231_i0;
  wire signed [`W-1:0] n1231_i1;
  wire signed [`W-1:0] n1231_i2;
  wire signed [`W-1:0] n1231_v;
  wire signed [`W-1:0] abl4_i0;
  wire signed [`W-1:0] abl4_i1;
  wire signed [`W-1:0] abl4_i2;
  wire signed [`W-1:0] abl4_i3;
  wire signed [`W-1:0] abl4_i4;
  wire signed [`W-1:0] abl4_v;
  wire signed [`W-1:0] op_T0_cpy_iny_i0;
  wire signed [`W-1:0] op_T0_cpy_iny_i1;
  wire signed [`W-1:0] op_T0_cpy_iny_i2;
  wire signed [`W-1:0] op_T0_cpy_iny_v;
  wire signed [`W-1:0] n1238_i0;
  wire signed [`W-1:0] n1238_i1;
  wire signed [`W-1:0] n1238_i2;
  wire signed [`W-1:0] n1238_v;
  wire signed [`W-1:0] op_T2_branch_i0;
  wire signed [`W-1:0] op_T2_branch_i1;
  wire signed [`W-1:0] op_T2_branch_i2;
  wire signed [`W-1:0] op_T2_branch_v;
  wire signed [`W-1:0] dpc38_PCLADL_i0;
  wire signed [`W-1:0] dpc38_PCLADL_i1;
  wire signed [`W-1:0] dpc38_PCLADL_i2;
  wire signed [`W-1:0] dpc38_PCLADL_i3;
  wire signed [`W-1:0] dpc38_PCLADL_i4;
  wire signed [`W-1:0] dpc38_PCLADL_i5;
  wire signed [`W-1:0] dpc38_PCLADL_i6;
  wire signed [`W-1:0] dpc38_PCLADL_i7;
  wire signed [`W-1:0] dpc38_PCLADL_i8;
  wire signed [`W-1:0] dpc38_PCLADL_i9;
  wire signed [`W-1:0] dpc38_PCLADL_v;
  wire signed [`W-1:0] Pout3_i0;
  wire signed [`W-1:0] Pout3_i1;
  wire signed [`W-1:0] Pout3_i2;
  wire signed [`W-1:0] Pout3_i3;
  wire signed [`W-1:0] Pout3_i4;
  wire signed [`W-1:0] Pout3_v;
  wire signed [`W-1:0] n436_i0;
  wire signed [`W-1:0] n436_i1;
  wire signed [`W-1:0] n436_i2;
  wire signed [`W-1:0] n436_i3;
  wire signed [`W-1:0] n436_v;
  wire signed [`W-1:0] dpc10_ADLADD_i0;
  wire signed [`W-1:0] dpc10_ADLADD_i1;
  wire signed [`W-1:0] dpc10_ADLADD_i2;
  wire signed [`W-1:0] dpc10_ADLADD_i3;
  wire signed [`W-1:0] dpc10_ADLADD_i4;
  wire signed [`W-1:0] dpc10_ADLADD_i5;
  wire signed [`W-1:0] dpc10_ADLADD_i6;
  wire signed [`W-1:0] dpc10_ADLADD_i7;
  wire signed [`W-1:0] dpc10_ADLADD_i8;
  wire signed [`W-1:0] dpc10_ADLADD_i9;
  wire signed [`W-1:0] dpc10_ADLADD_v;
  wire signed [`W-1:0] op_rmw_i0;
  wire signed [`W-1:0] op_rmw_i1;
  wire signed [`W-1:0] op_rmw_i2;
  wire signed [`W-1:0] op_rmw_v;
  wire signed [`W-1:0] ab4_i0;
  wire signed [`W-1:0] ab4_i1;
  wire signed [`W-1:0] ab4_i2;
  wire signed [`W-1:0] ab4_v;
  wire signed [`W-1:0] n432_i0;
  wire signed [`W-1:0] n432_i1;
  wire signed [`W-1:0] n432_i2;
  wire signed [`W-1:0] n432_i3;
  wire signed [`W-1:0] n432_v;
  wire signed [`W-1:0] n430_i0;
  wire signed [`W-1:0] n430_i1;
  wire signed [`W-1:0] n430_i2;
  wire signed [`W-1:0] n430_i3;
  wire signed [`W-1:0] n430_i4;
  wire signed [`W-1:0] n430_v;
  wire signed [`W-1:0] n238_i0;
  wire signed [`W-1:0] n238_i1;
  wire signed [`W-1:0] n238_i2;
  wire signed [`W-1:0] n238_v;
  wire signed [`W-1:0] abl5_i0;
  wire signed [`W-1:0] abl5_i1;
  wire signed [`W-1:0] abl5_i2;
  wire signed [`W-1:0] abl5_i3;
  wire signed [`W-1:0] abl5_i4;
  wire signed [`W-1:0] abl5_v;
  wire signed [`W-1:0] alub6_i0;
  wire signed [`W-1:0] alub6_i1;
  wire signed [`W-1:0] alub6_i2;
  wire signed [`W-1:0] alub6_i3;
  wire signed [`W-1:0] alub6_i4;
  wire signed [`W-1:0] alub6_v;
  wire signed [`W-1:0] n236_i0;
  wire signed [`W-1:0] n236_i1;
  wire signed [`W-1:0] n236_i2;
  wire signed [`W-1:0] n236_i3;
  wire signed [`W-1:0] n236_i4;
  wire signed [`W-1:0] n236_i5;
  wire signed [`W-1:0] n236_i6;
  wire signed [`W-1:0] n236_i7;
  wire signed [`W-1:0] n236_v;
  wire signed [`W-1:0] ab8_i0;
  wire signed [`W-1:0] ab8_i1;
  wire signed [`W-1:0] ab8_i2;
  wire signed [`W-1:0] ab8_v;
  wire signed [`W-1:0] n231_i0;
  wire signed [`W-1:0] n231_i1;
  wire signed [`W-1:0] n231_i2;
  wire signed [`W-1:0] n231_v;
  wire signed [`W-1:0] n232_i0;
  wire signed [`W-1:0] n232_i1;
  wire signed [`W-1:0] n232_i2;
  wire signed [`W-1:0] n232_i3;
  wire signed [`W-1:0] n232_i4;
  wire signed [`W-1:0] n232_v;
  wire signed [`W-1:0] n233_i0;
  wire signed [`W-1:0] n233_i1;
  wire signed [`W-1:0] n233_i2;
  wire signed [`W-1:0] n233_v;
  wire signed [`W-1:0] x2_i0;
  wire signed [`W-1:0] x2_i1;
  wire signed [`W-1:0] x2_i2;
  wire signed [`W-1:0] x2_v;
  wire signed [`W-1:0] n146_i0;
  wire signed [`W-1:0] n146_i1;
  wire signed [`W-1:0] n146_i2;
  wire signed [`W-1:0] n146_i3;
  wire signed [`W-1:0] n146_i4;
  wire signed [`W-1:0] n146_v;
  wire signed [`W-1:0] n147_i0;
  wire signed [`W-1:0] n147_i1;
  wire signed [`W-1:0] n147_i2;
  wire signed [`W-1:0] n147_v;
  wire signed [`W-1:0] op_sta_cmp_i0;
  wire signed [`W-1:0] op_sta_cmp_i1;
  wire signed [`W-1:0] op_sta_cmp_i2;
  wire signed [`W-1:0] op_sta_cmp_v;
  wire signed [`W-1:0] C45_i0;
  wire signed [`W-1:0] C45_i1;
  wire signed [`W-1:0] C45_i2;
  wire signed [`W-1:0] C45_i3;
  wire signed [`W-1:0] C45_v;
  wire signed [`W-1:0] aluanorb0_i0;
  wire signed [`W-1:0] aluanorb0_i1;
  wire signed [`W-1:0] aluanorb0_i2;
  wire signed [`W-1:0] aluanorb0_i3;
  wire signed [`W-1:0] aluanorb0_i4;
  wire signed [`W-1:0] aluanorb0_i5;
  wire signed [`W-1:0] aluanorb0_v;
  wire signed [`W-1:0] dpc27_SBADH_i0;
  wire signed [`W-1:0] dpc27_SBADH_i1;
  wire signed [`W-1:0] dpc27_SBADH_i2;
  wire signed [`W-1:0] dpc27_SBADH_i3;
  wire signed [`W-1:0] dpc27_SBADH_i4;
  wire signed [`W-1:0] dpc27_SBADH_i5;
  wire signed [`W-1:0] dpc27_SBADH_i6;
  wire signed [`W-1:0] dpc27_SBADH_i7;
  wire signed [`W-1:0] dpc27_SBADH_i8;
  wire signed [`W-1:0] dpc27_SBADH_i9;
  wire signed [`W-1:0] dpc27_SBADH_v;
  wire signed [`W-1:0] n141_i0;
  wire signed [`W-1:0] n141_i1;
  wire signed [`W-1:0] n141_i2;
  wire signed [`W-1:0] n141_i3;
  wire signed [`W-1:0] n141_i4;
  wire signed [`W-1:0] n141_v;
  wire signed [`W-1:0] ab9_i0;
  wire signed [`W-1:0] ab9_i1;
  wire signed [`W-1:0] ab9_i2;
  wire signed [`W-1:0] ab9_v;
  wire signed [`W-1:0] n149_i0;
  wire signed [`W-1:0] n149_i1;
  wire signed [`W-1:0] n149_i2;
  wire signed [`W-1:0] n149_i3;
  wire signed [`W-1:0] n149_v;
  wire signed [`W-1:0] aluvout_i0;
  wire signed [`W-1:0] aluvout_i1;
  wire signed [`W-1:0] aluvout_i2;
  wire signed [`W-1:0] aluvout_v;
  wire signed [`W-1:0] n933_i0;
  wire signed [`W-1:0] n933_i1;
  wire signed [`W-1:0] n933_i2;
  wire signed [`W-1:0] n933_v;
  wire signed [`W-1:0] op_T2_php_pha_i0;
  wire signed [`W-1:0] op_T2_php_pha_i1;
  wire signed [`W-1:0] op_T2_php_pha_i2;
  wire signed [`W-1:0] op_T2_php_pha_i3;
  wire signed [`W-1:0] op_T2_php_pha_v;
  wire signed [`W-1:0] n931_i0;
  wire signed [`W-1:0] n931_i1;
  wire signed [`W-1:0] n931_i2;
  wire signed [`W-1:0] n931_v;
  wire signed [`W-1:0] n930_i0;
  wire signed [`W-1:0] n930_i1;
  wire signed [`W-1:0] n930_i2;
  wire signed [`W-1:0] n930_v;
  wire signed [`W-1:0] n937_i0;
  wire signed [`W-1:0] n937_i1;
  wire signed [`W-1:0] n937_i2;
  wire signed [`W-1:0] n937_i3;
  wire signed [`W-1:0] n937_i4;
  wire signed [`W-1:0] n937_v;
  wire signed [`W-1:0] n936_i0;
  wire signed [`W-1:0] n936_i1;
  wire signed [`W-1:0] n936_i2;
  wire signed [`W-1:0] n936_i3;
  wire signed [`W-1:0] n936_i4;
  wire signed [`W-1:0] n936_i5;
  wire signed [`W-1:0] n936_v;
  wire signed [`W-1:0] n935_i0;
  wire signed [`W-1:0] n935_i1;
  wire signed [`W-1:0] n935_i2;
  wire signed [`W-1:0] n935_v;
  wire signed [`W-1:0] op_SRS_i0;
  wire signed [`W-1:0] op_SRS_i1;
  wire signed [`W-1:0] op_SRS_i2;
  wire signed [`W-1:0] op_SRS_i3;
  wire signed [`W-1:0] op_SRS_i4;
  wire signed [`W-1:0] op_SRS_i5;
  wire signed [`W-1:0] op_SRS_i6;
  wire signed [`W-1:0] op_SRS_v;
  wire signed [`W-1:0] pd5_i0;
  wire signed [`W-1:0] pd5_i1;
  wire signed [`W-1:0] pd5_v;
  wire signed [`W-1:0] nots3_i0;
  wire signed [`W-1:0] nots3_i1;
  wire signed [`W-1:0] nots3_v;
  wire signed [`W-1:0] _ABL3_i0;
  wire signed [`W-1:0] _ABL3_i1;
  wire signed [`W-1:0] _ABL3_i2;
  wire signed [`W-1:0] _ABL3_v;
  wire signed [`W-1:0] n824_i0;
  wire signed [`W-1:0] n824_i1;
  wire signed [`W-1:0] n824_i2;
  wire signed [`W-1:0] n824_i3;
  wire signed [`W-1:0] n824_i4;
  wire signed [`W-1:0] n824_v;
  wire signed [`W-1:0] D1x1_i0;
  wire signed [`W-1:0] D1x1_i1;
  wire signed [`W-1:0] D1x1_i2;
  wire signed [`W-1:0] D1x1_i3;
  wire signed [`W-1:0] D1x1_i4;
  wire signed [`W-1:0] D1x1_v;
  wire signed [`W-1:0] n826_i0;
  wire signed [`W-1:0] n826_i1;
  wire signed [`W-1:0] n826_i2;
  wire signed [`W-1:0] n826_v;
  wire signed [`W-1:0] ADH_ABH_i0;
  wire signed [`W-1:0] ADH_ABH_i1;
  wire signed [`W-1:0] ADH_ABH_i2;
  wire signed [`W-1:0] ADH_ABH_i3;
  wire signed [`W-1:0] ADH_ABH_i4;
  wire signed [`W-1:0] ADH_ABH_i5;
  wire signed [`W-1:0] ADH_ABH_i6;
  wire signed [`W-1:0] ADH_ABH_i7;
  wire signed [`W-1:0] ADH_ABH_i8;
  wire signed [`W-1:0] ADH_ABH_i9;
  wire signed [`W-1:0] ADH_ABH_v;
  wire signed [`W-1:0] pchp4_i0;
  wire signed [`W-1:0] pchp4_i1;
  wire signed [`W-1:0] pchp4_v;
  wire signed [`W-1:0] notdor3_i0;
  wire signed [`W-1:0] notdor3_i1;
  wire signed [`W-1:0] notdor3_v;
  wire signed [`W-1:0] op_T__adc_sbc_i0;
  wire signed [`W-1:0] op_T__adc_sbc_i1;
  wire signed [`W-1:0] op_T__adc_sbc_i2;
  wire signed [`W-1:0] op_T__adc_sbc_v;
  wire signed [`W-1:0] op_T__iny_dey_i0;
  wire signed [`W-1:0] op_T__iny_dey_i1;
  wire signed [`W-1:0] op_T__iny_dey_i2;
  wire signed [`W-1:0] op_T__iny_dey_v;
  wire signed [`W-1:0] VEC1_i0;
  wire signed [`W-1:0] VEC1_i1;
  wire signed [`W-1:0] VEC1_i2;
  wire signed [`W-1:0] VEC1_i3;
  wire signed [`W-1:0] VEC1_i4;
  wire signed [`W-1:0] VEC1_v;
  wire signed [`W-1:0] op_T3_plp_pla_i0;
  wire signed [`W-1:0] op_T3_plp_pla_i1;
  wire signed [`W-1:0] op_T3_plp_pla_i2;
  wire signed [`W-1:0] op_T3_plp_pla_v;
  wire signed [`W-1:0] n1486_i0;
  wire signed [`W-1:0] n1486_i1;
  wire signed [`W-1:0] n1486_i2;
  wire signed [`W-1:0] n1486_v;
  wire signed [`W-1:0] notidl2_i0;
  wire signed [`W-1:0] notidl2_i1;
  wire signed [`W-1:0] notidl2_v;
  wire signed [`W-1:0] n1484_i0;
  wire signed [`W-1:0] n1484_i1;
  wire signed [`W-1:0] n1484_i2;
  wire signed [`W-1:0] n1484_v;
  wire signed [`W-1:0] n1488_i0;
  wire signed [`W-1:0] n1488_i1;
  wire signed [`W-1:0] n1488_i2;
  wire signed [`W-1:0] n1488_i3;
  wire signed [`W-1:0] n1488_v;
  wire signed [`W-1:0] n797_i0;
  wire signed [`W-1:0] n797_i1;
  wire signed [`W-1:0] n797_i2;
  wire signed [`W-1:0] n797_v;
  wire signed [`W-1:0] n796_i0;
  wire signed [`W-1:0] n796_i1;
  wire signed [`W-1:0] n796_v;
  wire signed [`W-1:0] n795_i0;
  wire signed [`W-1:0] n795_i1;
  wire signed [`W-1:0] n795_i2;
  wire signed [`W-1:0] n795_v;
  wire signed [`W-1:0] n794_i0;
  wire signed [`W-1:0] n794_i1;
  wire signed [`W-1:0] n794_i2;
  wire signed [`W-1:0] n794_v;
  wire signed [`W-1:0] n1717_i0;
  wire signed [`W-1:0] n1717_i1;
  wire signed [`W-1:0] n1717_i2;
  wire signed [`W-1:0] n1717_v;
  wire signed [`W-1:0] n1716_i0;
  wire signed [`W-1:0] n1716_i1;
  wire signed [`W-1:0] n1716_i2;
  wire signed [`W-1:0] n1716_v;
  wire signed [`W-1:0] op_push_pull_i0;
  wire signed [`W-1:0] op_push_pull_i1;
  wire signed [`W-1:0] op_push_pull_i2;
  wire signed [`W-1:0] op_push_pull_i3;
  wire signed [`W-1:0] op_push_pull_v;
  wire signed [`W-1:0] n790_i0;
  wire signed [`W-1:0] n790_i1;
  wire signed [`W-1:0] n790_i2;
  wire signed [`W-1:0] n790_i3;
  wire signed [`W-1:0] n790_i4;
  wire signed [`W-1:0] n790_v;
  wire signed [`W-1:0] n1719_i0;
  wire signed [`W-1:0] n1719_i1;
  wire signed [`W-1:0] n1719_i2;
  wire signed [`W-1:0] n1719_v;
  wire signed [`W-1:0] n1718_i0;
  wire signed [`W-1:0] n1718_i1;
  wire signed [`W-1:0] n1718_i2;
  wire signed [`W-1:0] n1718_v;
  wire signed [`W-1:0] n799_i0;
  wire signed [`W-1:0] n799_i1;
  wire signed [`W-1:0] n799_v;
  wire signed [`W-1:0] n798_i0;
  wire signed [`W-1:0] n798_i1;
  wire signed [`W-1:0] n798_i2;
  wire signed [`W-1:0] n798_v;
  wire signed [`W-1:0] n1270_i0;
  wire signed [`W-1:0] n1270_i1;
  wire signed [`W-1:0] n1270_i2;
  wire signed [`W-1:0] n1270_i3;
  wire signed [`W-1:0] n1270_v;
  wire signed [`W-1:0] n1271_i0;
  wire signed [`W-1:0] n1271_i1;
  wire signed [`W-1:0] n1271_i2;
  wire signed [`W-1:0] n1271_v;
  wire signed [`W-1:0] n610_i0;
  wire signed [`W-1:0] n610_i1;
  wire signed [`W-1:0] n610_v;
  wire signed [`W-1:0] pcl0_i0;
  wire signed [`W-1:0] pcl0_i1;
  wire signed [`W-1:0] pcl0_i2;
  wire signed [`W-1:0] pcl0_v;
  wire signed [`W-1:0] n1138_i0;
  wire signed [`W-1:0] n1138_i1;
  wire signed [`W-1:0] n1138_i2;
  wire signed [`W-1:0] n1138_v;
  wire signed [`W-1:0] n1133_i0;
  wire signed [`W-1:0] n1133_i1;
  wire signed [`W-1:0] n1133_i2;
  wire signed [`W-1:0] n1133_v;
  wire signed [`W-1:0] n1132_i0;
  wire signed [`W-1:0] n1132_i1;
  wire signed [`W-1:0] n1132_v;
  wire signed [`W-1:0] pipe_WR_phi2_i0;
  wire signed [`W-1:0] pipe_WR_phi2_i1;
  wire signed [`W-1:0] pipe_WR_phi2_v;
  wire signed [`W-1:0] n1130_i0;
  wire signed [`W-1:0] n1130_i1;
  wire signed [`W-1:0] n1130_i2;
  wire signed [`W-1:0] n1130_i3;
  wire signed [`W-1:0] n1130_v;
  wire signed [`W-1:0] n1137_i0;
  wire signed [`W-1:0] n1137_i1;
  wire signed [`W-1:0] n1137_i2;
  wire signed [`W-1:0] n1137_v;
  wire signed [`W-1:0] a6_i0;
  wire signed [`W-1:0] a6_i1;
  wire signed [`W-1:0] a6_i2;
  wire signed [`W-1:0] a6_v;
  wire signed [`W-1:0] n1135_i0;
  wire signed [`W-1:0] n1135_i1;
  wire signed [`W-1:0] n1135_i2;
  wire signed [`W-1:0] n1135_i3;
  wire signed [`W-1:0] n1135_v;
  wire signed [`W-1:0] _VEC_i0;
  wire signed [`W-1:0] _VEC_i1;
  wire signed [`W-1:0] _VEC_i2;
  wire signed [`W-1:0] _VEC_i3;
  wire signed [`W-1:0] _VEC_i4;
  wire signed [`W-1:0] _VEC_v;
  wire signed [`W-1:0] n1276_i0;
  wire signed [`W-1:0] n1276_i1;
  wire signed [`W-1:0] n1276_v;
  wire signed [`W-1:0] n1277_i0;
  wire signed [`W-1:0] n1277_i1;
  wire signed [`W-1:0] n1277_i2;
  wire signed [`W-1:0] n1277_i3;
  wire signed [`W-1:0] n1277_v;
  wire signed [`W-1:0] n519_i0;
  wire signed [`W-1:0] n519_i1;
  wire signed [`W-1:0] n519_i2;
  wire signed [`W-1:0] n519_i3;
  wire signed [`W-1:0] n519_i4;
  wire signed [`W-1:0] n519_v;
  wire signed [`W-1:0] n518_i0;
  wire signed [`W-1:0] n518_i1;
  wire signed [`W-1:0] n518_i2;
  wire signed [`W-1:0] n518_i3;
  wire signed [`W-1:0] n518_v;
  wire signed [`W-1:0] dasb1_i0;
  wire signed [`W-1:0] dasb1_i1;
  wire signed [`W-1:0] dasb1_i2;
  wire signed [`W-1:0] dasb1_v;
  wire signed [`W-1:0] pipeUNK29_i0;
  wire signed [`W-1:0] pipeUNK29_i1;
  wire signed [`W-1:0] pipeUNK29_i2;
  wire signed [`W-1:0] pipeUNK29_v;
  wire signed [`W-1:0] n1007_i0;
  wire signed [`W-1:0] n1007_i1;
  wire signed [`W-1:0] n1007_i2;
  wire signed [`W-1:0] n1007_v;
  wire signed [`W-1:0] op_implied_i0;
  wire signed [`W-1:0] op_implied_i1;
  wire signed [`W-1:0] op_implied_i2;
  wire signed [`W-1:0] op_implied_v;
  wire signed [`W-1:0] db0_i0;
  wire signed [`W-1:0] db0_i1;
  wire signed [`W-1:0] db0_i2;
  wire signed [`W-1:0] db0_i3;
  wire signed [`W-1:0] db0_i4;
  wire signed [`W-1:0] db0_v;
  wire signed [`W-1:0] _C23_i0;
  wire signed [`W-1:0] _C23_i1;
  wire signed [`W-1:0] _C23_i2;
  wire signed [`W-1:0] _C23_i3;
  wire signed [`W-1:0] _C23_v;
  wire signed [`W-1:0] n1002_i0;
  wire signed [`W-1:0] n1002_i1;
  wire signed [`W-1:0] n1002_i2;
  wire signed [`W-1:0] n1002_i3;
  wire signed [`W-1:0] n1002_i4;
  wire signed [`W-1:0] n1002_i5;
  wire signed [`W-1:0] n1002_v;
  wire signed [`W-1:0] op_store_i0;
  wire signed [`W-1:0] op_store_i1;
  wire signed [`W-1:0] op_store_i2;
  wire signed [`W-1:0] op_store_v;
  wire signed [`W-1:0] pclp0_i0;
  wire signed [`W-1:0] pclp0_i1;
  wire signed [`W-1:0] pclp0_i2;
  wire signed [`W-1:0] pclp0_v;
  wire signed [`W-1:0] op_T0_plp_i0;
  wire signed [`W-1:0] op_T0_plp_i1;
  wire signed [`W-1:0] op_T0_plp_i2;
  wire signed [`W-1:0] op_T0_plp_v;
  wire signed [`W-1:0] n1225_i0;
  wire signed [`W-1:0] n1225_i1;
  wire signed [`W-1:0] n1225_i2;
  wire signed [`W-1:0] n1225_i3;
  wire signed [`W-1:0] n1225_i4;
  wire signed [`W-1:0] n1225_v;
  wire signed [`W-1:0] n620_i0;
  wire signed [`W-1:0] n620_i1;
  wire signed [`W-1:0] n620_i2;
  wire signed [`W-1:0] n620_i3;
  wire signed [`W-1:0] n620_v;
  wire signed [`W-1:0] n1223_i0;
  wire signed [`W-1:0] n1223_i1;
  wire signed [`W-1:0] n1223_i2;
  wire signed [`W-1:0] n1223_i3;
  wire signed [`W-1:0] n1223_v;
  wire signed [`W-1:0] n626_i0;
  wire signed [`W-1:0] n626_i1;
  wire signed [`W-1:0] n626_i2;
  wire signed [`W-1:0] n626_v;
  wire signed [`W-1:0] n625_i0;
  wire signed [`W-1:0] n625_i1;
  wire signed [`W-1:0] n625_i2;
  wire signed [`W-1:0] n625_i3;
  wire signed [`W-1:0] n625_v;
  wire signed [`W-1:0] AxB5_i0;
  wire signed [`W-1:0] AxB5_i1;
  wire signed [`W-1:0] AxB5_i2;
  wire signed [`W-1:0] AxB5_i3;
  wire signed [`W-1:0] AxB5_i4;
  wire signed [`W-1:0] AxB5_i5;
  wire signed [`W-1:0] AxB5_v;
  wire signed [`W-1:0] n629_i0;
  wire signed [`W-1:0] n629_i1;
  wire signed [`W-1:0] n629_i2;
  wire signed [`W-1:0] n629_v;
  wire signed [`W-1:0] n628_i0;
  wire signed [`W-1:0] n628_i1;
  wire signed [`W-1:0] n628_i2;
  wire signed [`W-1:0] n628_i3;
  wire signed [`W-1:0] n628_v;
  wire signed [`W-1:0] n1229_i0;
  wire signed [`W-1:0] n1229_i1;
  wire signed [`W-1:0] n1229_i2;
  wire signed [`W-1:0] n1229_v;
  wire signed [`W-1:0] op_ANDS_i0;
  wire signed [`W-1:0] op_ANDS_i1;
  wire signed [`W-1:0] op_ANDS_i2;
  wire signed [`W-1:0] op_ANDS_i3;
  wire signed [`W-1:0] op_ANDS_i4;
  wire signed [`W-1:0] op_ANDS_i5;
  wire signed [`W-1:0] op_ANDS_i6;
  wire signed [`W-1:0] op_ANDS_v;
  wire signed [`W-1:0] alub7_i0;
  wire signed [`W-1:0] alub7_i1;
  wire signed [`W-1:0] alub7_i2;
  wire signed [`W-1:0] alub7_i3;
  wire signed [`W-1:0] alub7_i4;
  wire signed [`W-1:0] alub7_v;
  wire signed [`W-1:0] n1286_i0;
  wire signed [`W-1:0] n1286_i1;
  wire signed [`W-1:0] n1286_i2;
  wire signed [`W-1:0] n1286_v;
  wire signed [`W-1:0] n11_i0;
  wire signed [`W-1:0] n11_i1;
  wire signed [`W-1:0] n11_i2;
  wire signed [`W-1:0] n11_v;
  wire signed [`W-1:0] n10_i0;
  wire signed [`W-1:0] n10_i1;
  wire signed [`W-1:0] n10_i2;
  wire signed [`W-1:0] n10_v;
  wire signed [`W-1:0] adh6_i0;
  wire signed [`W-1:0] adh6_i1;
  wire signed [`W-1:0] adh6_i2;
  wire signed [`W-1:0] adh6_i3;
  wire signed [`W-1:0] adh6_i4;
  wire signed [`W-1:0] adh6_i5;
  wire signed [`W-1:0] adh6_i6;
  wire signed [`W-1:0] adh6_v;
  wire signed [`W-1:0] n15_i0;
  wire signed [`W-1:0] n15_i1;
  wire signed [`W-1:0] n15_v;
  wire signed [`W-1:0] n14_i0;
  wire signed [`W-1:0] n14_i1;
  wire signed [`W-1:0] n14_i2;
  wire signed [`W-1:0] n14_v;
  wire signed [`W-1:0] n17_i0;
  wire signed [`W-1:0] n17_i1;
  wire signed [`W-1:0] n17_i2;
  wire signed [`W-1:0] n17_i3;
  wire signed [`W-1:0] n17_i4;
  wire signed [`W-1:0] n17_v;
  wire signed [`W-1:0] n16_i0;
  wire signed [`W-1:0] n16_i1;
  wire signed [`W-1:0] n16_i2;
  wire signed [`W-1:0] n16_i3;
  wire signed [`W-1:0] n16_i4;
  wire signed [`W-1:0] n16_i5;
  wire signed [`W-1:0] n16_v;
  wire signed [`W-1:0] n19_i0;
  wire signed [`W-1:0] n19_i1;
  wire signed [`W-1:0] n19_i2;
  wire signed [`W-1:0] n19_v;
  wire signed [`W-1:0] n18_i0;
  wire signed [`W-1:0] n18_i1;
  wire signed [`W-1:0] n18_v;
  wire signed [`W-1:0] n688_i0;
  wire signed [`W-1:0] n688_i1;
  wire signed [`W-1:0] n688_v;
  wire signed [`W-1:0] n201_i0;
  wire signed [`W-1:0] n201_i1;
  wire signed [`W-1:0] n201_i2;
  wire signed [`W-1:0] n201_i3;
  wire signed [`W-1:0] n201_v;
  wire signed [`W-1:0] n200_i0;
  wire signed [`W-1:0] n200_i1;
  wire signed [`W-1:0] n200_i2;
  wire signed [`W-1:0] n200_i3;
  wire signed [`W-1:0] n200_i4;
  wire signed [`W-1:0] n200_v;
  wire signed [`W-1:0] dpc29_0ADH17_i0;
  wire signed [`W-1:0] dpc29_0ADH17_i1;
  wire signed [`W-1:0] dpc29_0ADH17_i2;
  wire signed [`W-1:0] dpc29_0ADH17_i3;
  wire signed [`W-1:0] dpc29_0ADH17_i4;
  wire signed [`W-1:0] dpc29_0ADH17_i5;
  wire signed [`W-1:0] dpc29_0ADH17_i6;
  wire signed [`W-1:0] dpc29_0ADH17_i7;
  wire signed [`W-1:0] dpc29_0ADH17_i8;
  wire signed [`W-1:0] dpc29_0ADH17_v;
  wire signed [`W-1:0] pch7_i0;
  wire signed [`W-1:0] pch7_i1;
  wire signed [`W-1:0] pch7_i2;
  wire signed [`W-1:0] pch7_v;
  wire signed [`W-1:0] op_T2_ADL_ADD_i0;
  wire signed [`W-1:0] op_T2_ADL_ADD_i1;
  wire signed [`W-1:0] op_T2_ADL_ADD_i2;
  wire signed [`W-1:0] op_T2_ADL_ADD_v;
  wire signed [`W-1:0] n207_i0;
  wire signed [`W-1:0] n207_i1;
  wire signed [`W-1:0] n207_i2;
  wire signed [`W-1:0] n207_v;
  wire signed [`W-1:0] n206_i0;
  wire signed [`W-1:0] n206_i1;
  wire signed [`W-1:0] n206_i2;
  wire signed [`W-1:0] n206_i3;
  wire signed [`W-1:0] n206_i4;
  wire signed [`W-1:0] n206_i5;
  wire signed [`W-1:0] n206_v;
  wire signed [`W-1:0] n209_i0;
  wire signed [`W-1:0] n209_i1;
  wire signed [`W-1:0] n209_i2;
  wire signed [`W-1:0] n209_i3;
  wire signed [`W-1:0] n209_i4;
  wire signed [`W-1:0] n209_v;
  wire signed [`W-1:0] n208_i0;
  wire signed [`W-1:0] n208_i1;
  wire signed [`W-1:0] n208_i2;
  wire signed [`W-1:0] n208_i3;
  wire signed [`W-1:0] n208_i4;
  wire signed [`W-1:0] n208_v;
  wire signed [`W-1:0] n1573_i0;
  wire signed [`W-1:0] n1573_i1;
  wire signed [`W-1:0] n1573_i2;
  wire signed [`W-1:0] n1573_v;
  wire signed [`W-1:0] adl3_i0;
  wire signed [`W-1:0] adl3_i1;
  wire signed [`W-1:0] adl3_i2;
  wire signed [`W-1:0] adl3_i3;
  wire signed [`W-1:0] adl3_i4;
  wire signed [`W-1:0] adl3_i5;
  wire signed [`W-1:0] adl3_i6;
  wire signed [`W-1:0] adl3_i7;
  wire signed [`W-1:0] adl3_v;
  wire signed [`W-1:0] _C45_i0;
  wire signed [`W-1:0] _C45_i1;
  wire signed [`W-1:0] _C45_i2;
  wire signed [`W-1:0] _C45_i3;
  wire signed [`W-1:0] _C45_i4;
  wire signed [`W-1:0] _C45_v;
  wire signed [`W-1:0] n_0_ADL1_i0;
  wire signed [`W-1:0] n_0_ADL1_i1;
  wire signed [`W-1:0] n_0_ADL1_i2;
  wire signed [`W-1:0] n_0_ADL1_v;
  wire signed [`W-1:0] pipeUNK15_i0;
  wire signed [`W-1:0] pipeUNK15_i1;
  wire signed [`W-1:0] pipeUNK15_v;
  wire signed [`W-1:0] n680_i0;
  wire signed [`W-1:0] n680_i1;
  wire signed [`W-1:0] n680_v;
  wire signed [`W-1:0] pipedpc28_i0;
  wire signed [`W-1:0] pipedpc28_i1;
  wire signed [`W-1:0] pipedpc28_v;
  wire signed [`W-1:0] n1574_i0;
  wire signed [`W-1:0] n1574_i1;
  wire signed [`W-1:0] n1574_v;
  wire signed [`W-1:0] n928_i0;
  wire signed [`W-1:0] n928_i1;
  wire signed [`W-1:0] n928_i2;
  wire signed [`W-1:0] n928_v;
  wire signed [`W-1:0] n929_i0;
  wire signed [`W-1:0] n929_i1;
  wire signed [`W-1:0] n929_i2;
  wire signed [`W-1:0] n929_i3;
  wire signed [`W-1:0] n929_i4;
  wire signed [`W-1:0] n929_v;
  wire signed [`W-1:0] n920_i0;
  wire signed [`W-1:0] n920_i1;
  wire signed [`W-1:0] n920_i2;
  wire signed [`W-1:0] n920_v;
  wire signed [`W-1:0] dpc17_SUMS_i0;
  wire signed [`W-1:0] dpc17_SUMS_i1;
  wire signed [`W-1:0] dpc17_SUMS_i2;
  wire signed [`W-1:0] dpc17_SUMS_i3;
  wire signed [`W-1:0] dpc17_SUMS_i4;
  wire signed [`W-1:0] dpc17_SUMS_i5;
  wire signed [`W-1:0] dpc17_SUMS_i6;
  wire signed [`W-1:0] dpc17_SUMS_i7;
  wire signed [`W-1:0] dpc17_SUMS_i8;
  wire signed [`W-1:0] dpc17_SUMS_i9;
  wire signed [`W-1:0] dpc17_SUMS_v;
  wire signed [`W-1:0] n923_i0;
  wire signed [`W-1:0] n923_i1;
  wire signed [`W-1:0] n923_i2;
  wire signed [`W-1:0] n923_i3;
  wire signed [`W-1:0] n923_i4;
  wire signed [`W-1:0] n923_v;
  wire signed [`W-1:0] _op_store_i0;
  wire signed [`W-1:0] _op_store_i1;
  wire signed [`W-1:0] _op_store_i2;
  wire signed [`W-1:0] _op_store_i3;
  wire signed [`W-1:0] _op_store_v;
  wire signed [`W-1:0] C1x5Reset_i0;
  wire signed [`W-1:0] C1x5Reset_i1;
  wire signed [`W-1:0] C1x5Reset_i2;
  wire signed [`W-1:0] C1x5Reset_i3;
  wire signed [`W-1:0] C1x5Reset_i4;
  wire signed [`W-1:0] C1x5Reset_i5;
  wire signed [`W-1:0] C1x5Reset_v;
  wire signed [`W-1:0] n927_i0;
  wire signed [`W-1:0] n927_i1;
  wire signed [`W-1:0] n927_i2;
  wire signed [`W-1:0] n927_v;
  wire signed [`W-1:0] pipeUNK19_i0;
  wire signed [`W-1:0] pipeUNK19_i1;
  wire signed [`W-1:0] pipeUNK19_v;
  wire signed [`W-1:0] idb6_i0;
  wire signed [`W-1:0] idb6_i1;
  wire signed [`W-1:0] idb6_i2;
  wire signed [`W-1:0] idb6_i3;
  wire signed [`W-1:0] idb6_i4;
  wire signed [`W-1:0] idb6_i5;
  wire signed [`W-1:0] idb6_i6;
  wire signed [`W-1:0] idb6_i7;
  wire signed [`W-1:0] idb6_i8;
  wire signed [`W-1:0] idb6_i9;
  wire signed [`W-1:0] idb6_i10;
  wire signed [`W-1:0] idb6_i11;
  wire signed [`W-1:0] idb6_v;
  wire signed [`W-1:0] n830_i0;
  wire signed [`W-1:0] n830_i1;
  wire signed [`W-1:0] n830_i2;
  wire signed [`W-1:0] n830_i3;
  wire signed [`W-1:0] n830_v;
  wire signed [`W-1:0] n831_i0;
  wire signed [`W-1:0] n831_i1;
  wire signed [`W-1:0] n831_i2;
  wire signed [`W-1:0] n831_i3;
  wire signed [`W-1:0] n831_i4;
  wire signed [`W-1:0] n831_v;
  wire signed [`W-1:0] n837_i0;
  wire signed [`W-1:0] n837_i1;
  wire signed [`W-1:0] n837_i2;
  wire signed [`W-1:0] n837_v;
  wire signed [`W-1:0] n834_i0;
  wire signed [`W-1:0] n834_i1;
  wire signed [`W-1:0] n834_i2;
  wire signed [`W-1:0] n834_i3;
  wire signed [`W-1:0] n834_i4;
  wire signed [`W-1:0] n834_v;
  wire signed [`W-1:0] n838_i0;
  wire signed [`W-1:0] n838_i1;
  wire signed [`W-1:0] n838_i2;
  wire signed [`W-1:0] n838_v;
  wire signed [`W-1:0] n839_i0;
  wire signed [`W-1:0] n839_i1;
  wire signed [`W-1:0] n839_i2;
  wire signed [`W-1:0] n839_v;
  wire signed [`W-1:0] n3_i0;
  wire signed [`W-1:0] n3_i1;
  wire signed [`W-1:0] n3_i2;
  wire signed [`W-1:0] n3_i3;
  wire signed [`W-1:0] n3_i4;
  wire signed [`W-1:0] n3_v;
  wire signed [`W-1:0] op_T5_rti_i0;
  wire signed [`W-1:0] op_T5_rti_i1;
  wire signed [`W-1:0] op_T5_rti_i2;
  wire signed [`W-1:0] op_T5_rti_i3;
  wire signed [`W-1:0] op_T5_rti_v;
  wire signed [`W-1:0] n785_i0;
  wire signed [`W-1:0] n785_i1;
  wire signed [`W-1:0] n785_v;
  wire signed [`W-1:0] op_T__dex_i0;
  wire signed [`W-1:0] op_T__dex_i1;
  wire signed [`W-1:0] op_T__dex_i2;
  wire signed [`W-1:0] op_T__dex_v;
  wire signed [`W-1:0] op_T0_sbc_i0;
  wire signed [`W-1:0] op_T0_sbc_i1;
  wire signed [`W-1:0] op_T0_sbc_i2;
  wire signed [`W-1:0] op_T0_sbc_i3;
  wire signed [`W-1:0] op_T0_sbc_i4;
  wire signed [`W-1:0] op_T0_sbc_v;
  wire signed [`W-1:0] pchp0_i0;
  wire signed [`W-1:0] pchp0_i1;
  wire signed [`W-1:0] pchp0_v;
  wire signed [`W-1:0] n781_i0;
  wire signed [`W-1:0] n781_i1;
  wire signed [`W-1:0] n781_i2;
  wire signed [`W-1:0] n781_i3;
  wire signed [`W-1:0] n781_i4;
  wire signed [`W-1:0] n781_i5;
  wire signed [`W-1:0] n781_i6;
  wire signed [`W-1:0] n781_i7;
  wire signed [`W-1:0] n781_i8;
  wire signed [`W-1:0] n781_v;
  wire signed [`W-1:0] n782_i0;
  wire signed [`W-1:0] n782_i1;
  wire signed [`W-1:0] n782_i2;
  wire signed [`W-1:0] n782_v;
  wire signed [`W-1:0] n783_i0;
  wire signed [`W-1:0] n783_i1;
  wire signed [`W-1:0] n783_i2;
  wire signed [`W-1:0] n783_i3;
  wire signed [`W-1:0] n783_i4;
  wire signed [`W-1:0] n783_v;
  wire signed [`W-1:0] n1724_i0;
  wire signed [`W-1:0] n1724_i1;
  wire signed [`W-1:0] n1724_i2;
  wire signed [`W-1:0] n1724_i3;
  wire signed [`W-1:0] n1724_v;
  wire signed [`W-1:0] op_T2_i0;
  wire signed [`W-1:0] op_T2_i1;
  wire signed [`W-1:0] op_T2_i2;
  wire signed [`W-1:0] op_T2_v;
  wire signed [`W-1:0] n789_i0;
  wire signed [`W-1:0] n789_i1;
  wire signed [`W-1:0] n789_i2;
  wire signed [`W-1:0] n789_v;
  wire signed [`W-1:0] n1720_i0;
  wire signed [`W-1:0] n1720_i1;
  wire signed [`W-1:0] n1720_i2;
  wire signed [`W-1:0] n1720_i3;
  wire signed [`W-1:0] n1720_v;
  wire signed [`W-1:0] op_branch_done_i0;
  wire signed [`W-1:0] op_branch_done_i1;
  wire signed [`W-1:0] op_branch_done_i2;
  wire signed [`W-1:0] op_branch_done_i3;
  wire signed [`W-1:0] op_branch_done_v;
  wire signed [`W-1:0] op_T3_ind_y_i0;
  wire signed [`W-1:0] op_T3_ind_y_i1;
  wire signed [`W-1:0] op_T3_ind_y_i2;
  wire signed [`W-1:0] op_T3_ind_y_v;
  wire signed [`W-1:0] n61_i0;
  wire signed [`W-1:0] n61_i1;
  wire signed [`W-1:0] n61_i2;
  wire signed [`W-1:0] n61_i3;
  wire signed [`W-1:0] n61_v;
  wire signed [`W-1:0] n62_i0;
  wire signed [`W-1:0] n62_i1;
  wire signed [`W-1:0] n62_i2;
  wire signed [`W-1:0] n62_v;
  wire signed [`W-1:0] dor7_i0;
  wire signed [`W-1:0] dor7_i1;
  wire signed [`W-1:0] dor7_i2;
  wire signed [`W-1:0] dor7_i3;
  wire signed [`W-1:0] dor7_i4;
  wire signed [`W-1:0] dor7_v;
  wire signed [`W-1:0] y0_i0;
  wire signed [`W-1:0] y0_i1;
  wire signed [`W-1:0] y0_i2;
  wire signed [`W-1:0] y0_v;
  wire signed [`W-1:0] _AxB_4__C34_i0;
  wire signed [`W-1:0] _AxB_4__C34_i1;
  wire signed [`W-1:0] _AxB_4__C34_i2;
  wire signed [`W-1:0] _AxB_4__C34_v;
  wire signed [`W-1:0] n66_i0;
  wire signed [`W-1:0] n66_i1;
  wire signed [`W-1:0] n66_i2;
  wire signed [`W-1:0] n66_i3;
  wire signed [`W-1:0] n66_v;
  wire signed [`W-1:0] Reset0_i0;
  wire signed [`W-1:0] Reset0_i1;
  wire signed [`W-1:0] Reset0_i2;
  wire signed [`W-1:0] Reset0_i3;
  wire signed [`W-1:0] Reset0_i4;
  wire signed [`W-1:0] Reset0_i5;
  wire signed [`W-1:0] Reset0_v;
  wire signed [`W-1:0] notalu6_i0;
  wire signed [`W-1:0] notalu6_i1;
  wire signed [`W-1:0] notalu6_v;
  wire signed [`W-1:0] n69_i0;
  wire signed [`W-1:0] n69_i1;
  wire signed [`W-1:0] n69_v;
  wire signed [`W-1:0] adh0_i0;
  wire signed [`W-1:0] adh0_i1;
  wire signed [`W-1:0] adh0_i2;
  wire signed [`W-1:0] adh0_i3;
  wire signed [`W-1:0] adh0_i4;
  wire signed [`W-1:0] adh0_i5;
  wire signed [`W-1:0] adh0_i6;
  wire signed [`W-1:0] adh0_v;
  wire signed [`W-1:0] n1588_i0;
  wire signed [`W-1:0] n1588_i1;
  wire signed [`W-1:0] n1588_i2;
  wire signed [`W-1:0] n1588_v;
  wire signed [`W-1:0] op_T4_jmp_i0;
  wire signed [`W-1:0] op_T4_jmp_i1;
  wire signed [`W-1:0] op_T4_jmp_i2;
  wire signed [`W-1:0] op_T4_jmp_i3;
  wire signed [`W-1:0] op_T4_jmp_v;
  wire signed [`W-1:0] op_T2_stack_i0;
  wire signed [`W-1:0] op_T2_stack_i1;
  wire signed [`W-1:0] op_T2_stack_i2;
  wire signed [`W-1:0] op_T2_stack_i3;
  wire signed [`W-1:0] op_T2_stack_v;
  wire signed [`W-1:0] n1580_i0;
  wire signed [`W-1:0] n1580_i1;
  wire signed [`W-1:0] n1580_i2;
  wire signed [`W-1:0] n1580_i3;
  wire signed [`W-1:0] n1580_v;
  wire signed [`W-1:0] n1581_i0;
  wire signed [`W-1:0] n1581_i1;
  wire signed [`W-1:0] n1581_v;
  wire signed [`W-1:0] n1586_i0;
  wire signed [`W-1:0] n1586_i1;
  wire signed [`W-1:0] n1586_i2;
  wire signed [`W-1:0] n1586_v;
  wire signed [`W-1:0] pipeT4out_i0;
  wire signed [`W-1:0] pipeT4out_i1;
  wire signed [`W-1:0] pipeT4out_i2;
  wire signed [`W-1:0] pipeT4out_v;
  wire signed [`W-1:0] n1585_i0;
  wire signed [`W-1:0] n1585_i1;
  wire signed [`W-1:0] n1585_i2;
  wire signed [`W-1:0] n1585_v;
  wire signed [`W-1:0] n1038_i0;
  wire signed [`W-1:0] n1038_i1;
  wire signed [`W-1:0] n1038_i2;
  wire signed [`W-1:0] n1038_v;
  wire signed [`W-1:0] DC34_i0;
  wire signed [`W-1:0] DC34_i1;
  wire signed [`W-1:0] DC34_i2;
  wire signed [`W-1:0] DC34_v;
  wire signed [`W-1:0] n509_i0;
  wire signed [`W-1:0] n509_i1;
  wire signed [`W-1:0] n509_v;
  wire signed [`W-1:0] NMIP_i0;
  wire signed [`W-1:0] NMIP_i1;
  wire signed [`W-1:0] NMIP_i2;
  wire signed [`W-1:0] NMIP_i3;
  wire signed [`W-1:0] NMIP_v;
  wire signed [`W-1:0] op_T0_ora_i0;
  wire signed [`W-1:0] op_T0_ora_i1;
  wire signed [`W-1:0] op_T0_ora_i2;
  wire signed [`W-1:0] op_T0_ora_v;
  wire signed [`W-1:0] op_T3_stack_bit_jmp_i0;
  wire signed [`W-1:0] op_T3_stack_bit_jmp_i1;
  wire signed [`W-1:0] op_T3_stack_bit_jmp_i2;
  wire signed [`W-1:0] op_T3_stack_bit_jmp_v;
  wire signed [`W-1:0] pch2_i0;
  wire signed [`W-1:0] pch2_i1;
  wire signed [`W-1:0] pch2_i2;
  wire signed [`W-1:0] pch2_v;
  wire signed [`W-1:0] n1037_i0;
  wire signed [`W-1:0] n1037_i1;
  wire signed [`W-1:0] n1037_i2;
  wire signed [`W-1:0] n1037_v;
  wire signed [`W-1:0] C56_i0;
  wire signed [`W-1:0] C56_i1;
  wire signed [`W-1:0] C56_i2;
  wire signed [`W-1:0] C56_i3;
  wire signed [`W-1:0] C56_v;
  wire signed [`W-1:0] n402_i0;
  wire signed [`W-1:0] n402_i1;
  wire signed [`W-1:0] n402_v;
  wire signed [`W-1:0] n630_i0;
  wire signed [`W-1:0] n630_i1;
  wire signed [`W-1:0] n630_i2;
  wire signed [`W-1:0] n630_i3;
  wire signed [`W-1:0] n630_v;
  wire signed [`W-1:0] n631_i0;
  wire signed [`W-1:0] n631_i1;
  wire signed [`W-1:0] n631_i2;
  wire signed [`W-1:0] n631_i3;
  wire signed [`W-1:0] n631_v;
  wire signed [`W-1:0] op_T5_ind_x_i0;
  wire signed [`W-1:0] op_T5_ind_x_i1;
  wire signed [`W-1:0] op_T5_ind_x_i2;
  wire signed [`W-1:0] op_T5_ind_x_i3;
  wire signed [`W-1:0] op_T5_ind_x_v;
  wire signed [`W-1:0] n1211_i0;
  wire signed [`W-1:0] n1211_i1;
  wire signed [`W-1:0] n1211_i2;
  wire signed [`W-1:0] n1211_i3;
  wire signed [`W-1:0] n1211_i4;
  wire signed [`W-1:0] n1211_v;
  wire signed [`W-1:0] n634_i0;
  wire signed [`W-1:0] n634_i1;
  wire signed [`W-1:0] n634_i2;
  wire signed [`W-1:0] n634_v;
  wire signed [`W-1:0] __AxB7__C67_i0;
  wire signed [`W-1:0] __AxB7__C67_i1;
  wire signed [`W-1:0] __AxB7__C67_i2;
  wire signed [`W-1:0] __AxB7__C67_v;
  wire signed [`W-1:0] n1214_i0;
  wire signed [`W-1:0] n1214_i1;
  wire signed [`W-1:0] n1214_i2;
  wire signed [`W-1:0] n1214_v;
  wire signed [`W-1:0] n637_i0;
  wire signed [`W-1:0] n637_i1;
  wire signed [`W-1:0] n637_i2;
  wire signed [`W-1:0] n637_v;
  wire signed [`W-1:0] n638_i0;
  wire signed [`W-1:0] n638_i1;
  wire signed [`W-1:0] n638_i2;
  wire signed [`W-1:0] n638_v;
  wire signed [`W-1:0] ADL_ABL_i0;
  wire signed [`W-1:0] ADL_ABL_i1;
  wire signed [`W-1:0] ADL_ABL_i2;
  wire signed [`W-1:0] ADL_ABL_i3;
  wire signed [`W-1:0] ADL_ABL_i4;
  wire signed [`W-1:0] ADL_ABL_i5;
  wire signed [`W-1:0] ADL_ABL_i6;
  wire signed [`W-1:0] ADL_ABL_i7;
  wire signed [`W-1:0] ADL_ABL_i8;
  wire signed [`W-1:0] ADL_ABL_i9;
  wire signed [`W-1:0] ADL_ABL_v;
  wire signed [`W-1:0] n1218_i0;
  wire signed [`W-1:0] n1218_i1;
  wire signed [`W-1:0] n1218_i2;
  wire signed [`W-1:0] n1218_v;
  wire signed [`W-1:0] n1376_i0;
  wire signed [`W-1:0] n1376_i1;
  wire signed [`W-1:0] n1376_i2;
  wire signed [`W-1:0] n1376_v;
  wire signed [`W-1:0] n465_i0;
  wire signed [`W-1:0] n465_i1;
  wire signed [`W-1:0] n465_i2;
  wire signed [`W-1:0] n465_v;
  wire signed [`W-1:0] n1107_i0;
  wire signed [`W-1:0] n1107_i1;
  wire signed [`W-1:0] n1107_i2;
  wire signed [`W-1:0] n1107_v;
  wire signed [`W-1:0] pipeUNK42_i0;
  wire signed [`W-1:0] pipeUNK42_i1;
  wire signed [`W-1:0] pipeUNK42_v;
  wire signed [`W-1:0] n1105_i0;
  wire signed [`W-1:0] n1105_i1;
  wire signed [`W-1:0] n1105_i2;
  wire signed [`W-1:0] n1105_v;
  wire signed [`W-1:0] n1450_i0;
  wire signed [`W-1:0] n1450_i1;
  wire signed [`W-1:0] n1450_v;
  wire signed [`W-1:0] n1452_i0;
  wire signed [`W-1:0] n1452_i1;
  wire signed [`W-1:0] n1452_v;
  wire signed [`W-1:0] dor5_i0;
  wire signed [`W-1:0] dor5_i1;
  wire signed [`W-1:0] dor5_i2;
  wire signed [`W-1:0] dor5_i3;
  wire signed [`W-1:0] dor5_i4;
  wire signed [`W-1:0] dor5_v;
  wire signed [`W-1:0] n1458_i0;
  wire signed [`W-1:0] n1458_i1;
  wire signed [`W-1:0] n1458_i2;
  wire signed [`W-1:0] n1458_i3;
  wire signed [`W-1:0] n1458_i4;
  wire signed [`W-1:0] n1458_v;
  wire signed [`W-1:0] __AxB_6_i0;
  wire signed [`W-1:0] __AxB_6_i1;
  wire signed [`W-1:0] __AxB_6_i2;
  wire signed [`W-1:0] __AxB_6_i3;
  wire signed [`W-1:0] __AxB_6_i4;
  wire signed [`W-1:0] __AxB_6_i5;
  wire signed [`W-1:0] __AxB_6_i6;
  wire signed [`W-1:0] __AxB_6_v;
  wire signed [`W-1:0] idb0_i0;
  wire signed [`W-1:0] idb0_i1;
  wire signed [`W-1:0] idb0_i2;
  wire signed [`W-1:0] idb0_i3;
  wire signed [`W-1:0] idb0_i4;
  wire signed [`W-1:0] idb0_i5;
  wire signed [`W-1:0] idb0_i6;
  wire signed [`W-1:0] idb0_i7;
  wire signed [`W-1:0] idb0_i8;
  wire signed [`W-1:0] idb0_i9;
  wire signed [`W-1:0] idb0_i10;
  wire signed [`W-1:0] idb0_i11;
  wire signed [`W-1:0] idb0_v;
  wire signed [`W-1:0] n1109_i0;
  wire signed [`W-1:0] n1109_i1;
  wire signed [`W-1:0] n1109_i2;
  wire signed [`W-1:0] n1109_i3;
  wire signed [`W-1:0] n1109_i4;
  wire signed [`W-1:0] n1109_v;
  wire signed [`W-1:0] n1722_i0;
  wire signed [`W-1:0] n1722_i1;
  wire signed [`W-1:0] n1722_i2;
  wire signed [`W-1:0] n1722_i3;
  wire signed [`W-1:0] n1722_i4;
  wire signed [`W-1:0] n1722_v;
  wire signed [`W-1:0] DA_AB2_i0;
  wire signed [`W-1:0] DA_AB2_i1;
  wire signed [`W-1:0] DA_AB2_i2;
  wire signed [`W-1:0] DA_AB2_i3;
  wire signed [`W-1:0] DA_AB2_v;
  wire signed [`W-1:0] n_0_ADL0_i0;
  wire signed [`W-1:0] n_0_ADL0_i1;
  wire signed [`W-1:0] n_0_ADL0_i2;
  wire signed [`W-1:0] n_0_ADL0_i3;
  wire signed [`W-1:0] n_0_ADL0_v;
  wire signed [`W-1:0] dpc19_ADDSB7_i0;
  wire signed [`W-1:0] dpc19_ADDSB7_i1;
  wire signed [`W-1:0] dpc19_ADDSB7_i2;
  wire signed [`W-1:0] dpc19_ADDSB7_v;
  wire signed [`W-1:0] pipeUNK10_i0;
  wire signed [`W-1:0] pipeUNK10_i1;
  wire signed [`W-1:0] pipeUNK10_v;
  wire signed [`W-1:0] n212_i0;
  wire signed [`W-1:0] n212_i1;
  wire signed [`W-1:0] n212_i2;
  wire signed [`W-1:0] n212_v;
  wire signed [`W-1:0] n213_i0;
  wire signed [`W-1:0] n213_i1;
  wire signed [`W-1:0] n213_i2;
  wire signed [`W-1:0] n213_v;
  wire signed [`W-1:0] n210_i0;
  wire signed [`W-1:0] n210_i1;
  wire signed [`W-1:0] n210_i2;
  wire signed [`W-1:0] n210_i3;
  wire signed [`W-1:0] n210_v;
  wire signed [`W-1:0] ab3_i0;
  wire signed [`W-1:0] ab3_i1;
  wire signed [`W-1:0] ab3_i2;
  wire signed [`W-1:0] ab3_v;
  wire signed [`W-1:0] n218_i0;
  wire signed [`W-1:0] n218_i1;
  wire signed [`W-1:0] n218_i2;
  wire signed [`W-1:0] n218_v;
  wire signed [`W-1:0] op_T2_mem_zp_i0;
  wire signed [`W-1:0] op_T2_mem_zp_i1;
  wire signed [`W-1:0] op_T2_mem_zp_i2;
  wire signed [`W-1:0] op_T2_mem_zp_v;
  wire signed [`W-1:0] op_T0_tay_i0;
  wire signed [`W-1:0] op_T0_tay_i1;
  wire signed [`W-1:0] op_T0_tay_i2;
  wire signed [`W-1:0] op_T0_tay_v;
  wire signed [`W-1:0] n919_i0;
  wire signed [`W-1:0] n919_i1;
  wire signed [`W-1:0] n919_i2;
  wire signed [`W-1:0] n919_i3;
  wire signed [`W-1:0] n919_i4;
  wire signed [`W-1:0] n919_v;
  wire signed [`W-1:0] n918_i0;
  wire signed [`W-1:0] n918_i1;
  wire signed [`W-1:0] n918_i2;
  wire signed [`W-1:0] n918_v;
  wire signed [`W-1:0] n917_i0;
  wire signed [`W-1:0] n917_i1;
  wire signed [`W-1:0] n917_i2;
  wire signed [`W-1:0] n917_v;
  wire signed [`W-1:0] n916_i0;
  wire signed [`W-1:0] n916_i1;
  wire signed [`W-1:0] n916_i2;
  wire signed [`W-1:0] n916_i3;
  wire signed [`W-1:0] n916_v;
  wire signed [`W-1:0] alucin_i0;
  wire signed [`W-1:0] alucin_i1;
  wire signed [`W-1:0] alucin_i2;
  wire signed [`W-1:0] alucin_v;
  wire signed [`W-1:0] n913_i0;
  wire signed [`W-1:0] n913_i1;
  wire signed [`W-1:0] n913_i2;
  wire signed [`W-1:0] n913_v;
  wire signed [`W-1:0] n847_i0;
  wire signed [`W-1:0] n847_i1;
  wire signed [`W-1:0] n847_i2;
  wire signed [`W-1:0] n847_v;
  wire signed [`W-1:0] n846_i0;
  wire signed [`W-1:0] n846_i1;
  wire signed [`W-1:0] n846_i2;
  wire signed [`W-1:0] n846_i3;
  wire signed [`W-1:0] n846_v;
  wire signed [`W-1:0] n845_i0;
  wire signed [`W-1:0] n845_i1;
  wire signed [`W-1:0] n845_i2;
  wire signed [`W-1:0] n845_v;
  wire signed [`W-1:0] n844_i0;
  wire signed [`W-1:0] n844_i1;
  wire signed [`W-1:0] n844_i2;
  wire signed [`W-1:0] n844_i3;
  wire signed [`W-1:0] n844_v;
  wire signed [`W-1:0] y7_i0;
  wire signed [`W-1:0] y7_i1;
  wire signed [`W-1:0] y7_i2;
  wire signed [`W-1:0] y7_v;
  wire signed [`W-1:0] n842_i0;
  wire signed [`W-1:0] n842_i1;
  wire signed [`W-1:0] n842_i2;
  wire signed [`W-1:0] n842_i3;
  wire signed [`W-1:0] n842_v;
  wire signed [`W-1:0] aluanandb1_i0;
  wire signed [`W-1:0] aluanandb1_i1;
  wire signed [`W-1:0] aluanandb1_i2;
  wire signed [`W-1:0] aluanandb1_i3;
  wire signed [`W-1:0] aluanandb1_i4;
  wire signed [`W-1:0] aluanandb1_v;
  wire signed [`W-1:0] _op_branch_bit6_i0;
  wire signed [`W-1:0] _op_branch_bit6_i1;
  wire signed [`W-1:0] _op_branch_bit6_i2;
  wire signed [`W-1:0] _op_branch_bit6_i3;
  wire signed [`W-1:0] _op_branch_bit6_i4;
  wire signed [`W-1:0] _op_branch_bit6_v;
  wire signed [`W-1:0] n849_i0;
  wire signed [`W-1:0] n849_i1;
  wire signed [`W-1:0] n849_i2;
  wire signed [`W-1:0] n849_v;
  wire signed [`W-1:0] pipeUNK33_i0;
  wire signed [`W-1:0] pipeUNK33_i1;
  wire signed [`W-1:0] pipeUNK33_v;
  wire signed [`W-1:0] n663_i0;
  wire signed [`W-1:0] n663_i1;
  wire signed [`W-1:0] n663_v;
  wire signed [`W-1:0] pd3_clearIR_i0;
  wire signed [`W-1:0] pd3_clearIR_i1;
  wire signed [`W-1:0] pd3_clearIR_i2;
  wire signed [`W-1:0] pd3_clearIR_i3;
  wire signed [`W-1:0] pd3_clearIR_v;
  wire signed [`W-1:0] n662_i0;
  wire signed [`W-1:0] n662_i1;
  wire signed [`W-1:0] n662_i2;
  wire signed [`W-1:0] n662_v;
  wire signed [`W-1:0] n1039_i0;
  wire signed [`W-1:0] n1039_i1;
  wire signed [`W-1:0] n1039_i2;
  wire signed [`W-1:0] n1039_v;
  wire signed [`W-1:0] n753_i0;
  wire signed [`W-1:0] n753_i1;
  wire signed [`W-1:0] n753_i2;
  wire signed [`W-1:0] n753_i3;
  wire signed [`W-1:0] n753_v;
  wire signed [`W-1:0] nots2_i0;
  wire signed [`W-1:0] nots2_i1;
  wire signed [`W-1:0] nots2_v;
  wire signed [`W-1:0] pchp6_i0;
  wire signed [`W-1:0] pchp6_i1;
  wire signed [`W-1:0] pchp6_v;
  wire signed [`W-1:0] op_T2_php_i0;
  wire signed [`W-1:0] op_T2_php_i1;
  wire signed [`W-1:0] op_T2_php_i2;
  wire signed [`W-1:0] op_T2_php_v;
  wire signed [`W-1:0] n757_i0;
  wire signed [`W-1:0] n757_i1;
  wire signed [`W-1:0] n757_i2;
  wire signed [`W-1:0] n757_v;
  wire signed [`W-1:0] n756_i0;
  wire signed [`W-1:0] n756_i1;
  wire signed [`W-1:0] n756_v;
  wire signed [`W-1:0] n755_i0;
  wire signed [`W-1:0] n755_i1;
  wire signed [`W-1:0] n755_i2;
  wire signed [`W-1:0] n755_i3;
  wire signed [`W-1:0] n755_v;
  wire signed [`W-1:0] n754_i0;
  wire signed [`W-1:0] n754_i1;
  wire signed [`W-1:0] n754_i2;
  wire signed [`W-1:0] n754_i3;
  wire signed [`W-1:0] n754_v;
  wire signed [`W-1:0] n759_i0;
  wire signed [`W-1:0] n759_i1;
  wire signed [`W-1:0] n759_v;
  wire signed [`W-1:0] pd0_i0;
  wire signed [`W-1:0] pd0_i1;
  wire signed [`W-1:0] pd0_v;
  wire signed [`W-1:0] n1595_i0;
  wire signed [`W-1:0] n1595_i1;
  wire signed [`W-1:0] n1595_i2;
  wire signed [`W-1:0] n1595_v;
  wire signed [`W-1:0] n506_i0;
  wire signed [`W-1:0] n506_i1;
  wire signed [`W-1:0] n506_i2;
  wire signed [`W-1:0] n506_i3;
  wire signed [`W-1:0] n506_v;
  wire signed [`W-1:0] idl0_i0;
  wire signed [`W-1:0] idl0_i1;
  wire signed [`W-1:0] idl0_i2;
  wire signed [`W-1:0] idl0_v;
  wire signed [`W-1:0] n1596_i0;
  wire signed [`W-1:0] n1596_i1;
  wire signed [`W-1:0] n1596_i2;
  wire signed [`W-1:0] n1596_i3;
  wire signed [`W-1:0] n1596_v;
  wire signed [`W-1:0] db6_i0;
  wire signed [`W-1:0] db6_i1;
  wire signed [`W-1:0] db6_i2;
  wire signed [`W-1:0] db6_i3;
  wire signed [`W-1:0] db6_i4;
  wire signed [`W-1:0] db6_v;
  wire signed [`W-1:0] n1593_i0;
  wire signed [`W-1:0] n1593_i1;
  wire signed [`W-1:0] n1593_i2;
  wire signed [`W-1:0] n1593_i3;
  wire signed [`W-1:0] n1593_v;
  wire signed [`W-1:0] n1033_i0;
  wire signed [`W-1:0] n1033_i1;
  wire signed [`W-1:0] n1033_i2;
  wire signed [`W-1:0] n1033_v;
  wire signed [`W-1:0] n1599_i0;
  wire signed [`W-1:0] n1599_i1;
  wire signed [`W-1:0] n1599_i2;
  wire signed [`W-1:0] n1599_i3;
  wire signed [`W-1:0] n1599_v;
  wire signed [`W-1:0] n1025_i0;
  wire signed [`W-1:0] n1025_i1;
  wire signed [`W-1:0] n1025_i2;
  wire signed [`W-1:0] n1025_v;
  wire signed [`W-1:0] n1024_i0;
  wire signed [`W-1:0] n1024_i1;
  wire signed [`W-1:0] n1024_i2;
  wire signed [`W-1:0] n1024_i3;
  wire signed [`W-1:0] n1024_v;
  wire signed [`W-1:0] n1027_i0;
  wire signed [`W-1:0] n1027_i1;
  wire signed [`W-1:0] n1027_v;
  wire signed [`W-1:0] C12_i0;
  wire signed [`W-1:0] C12_i1;
  wire signed [`W-1:0] C12_i2;
  wire signed [`W-1:0] C12_i3;
  wire signed [`W-1:0] C12_v;
  wire signed [`W-1:0] aluaorb1_i0;
  wire signed [`W-1:0] aluaorb1_i1;
  wire signed [`W-1:0] aluaorb1_i2;
  wire signed [`W-1:0] aluaorb1_v;
  wire signed [`W-1:0] n1020_i0;
  wire signed [`W-1:0] n1020_i1;
  wire signed [`W-1:0] n1020_v;
  wire signed [`W-1:0] C23_i0;
  wire signed [`W-1:0] C23_i1;
  wire signed [`W-1:0] C23_i2;
  wire signed [`W-1:0] C23_i3;
  wire signed [`W-1:0] C23_v;
  wire signed [`W-1:0] pcl1_i0;
  wire signed [`W-1:0] pcl1_i1;
  wire signed [`W-1:0] pcl1_i2;
  wire signed [`W-1:0] pcl1_v;
  wire signed [`W-1:0] pipephi2Reset0x_i0;
  wire signed [`W-1:0] pipephi2Reset0x_i1;
  wire signed [`W-1:0] pipephi2Reset0x_v;
  wire signed [`W-1:0] nots6_i0;
  wire signed [`W-1:0] nots6_i1;
  wire signed [`W-1:0] nots6_v;
  wire signed [`W-1:0] n1028_i0;
  wire signed [`W-1:0] n1028_i1;
  wire signed [`W-1:0] n1028_i2;
  wire signed [`W-1:0] n1028_v;
  wire signed [`W-1:0] n503_i0;
  wire signed [`W-1:0] n503_i1;
  wire signed [`W-1:0] n503_i2;
  wire signed [`W-1:0] n503_v;
  wire signed [`W-1:0] n1034_i0;
  wire signed [`W-1:0] n1034_i1;
  wire signed [`W-1:0] n1034_i2;
  wire signed [`W-1:0] n1034_i3;
  wire signed [`W-1:0] n1034_v;
  wire signed [`W-1:0] n501_i0;
  wire signed [`W-1:0] n501_i1;
  wire signed [`W-1:0] n501_i2;
  wire signed [`W-1:0] n501_v;
  wire signed [`W-1:0] s6_i0;
  wire signed [`W-1:0] s6_i1;
  wire signed [`W-1:0] s6_i2;
  wire signed [`W-1:0] s6_v;
  wire signed [`W-1:0] op_T3_mem_abs_i0;
  wire signed [`W-1:0] op_T3_mem_abs_i1;
  wire signed [`W-1:0] op_T3_mem_abs_i2;
  wire signed [`W-1:0] op_T3_mem_abs_v;
  wire signed [`W-1:0] alu4_i0;
  wire signed [`W-1:0] alu4_i1;
  wire signed [`W-1:0] alu4_i2;
  wire signed [`W-1:0] alu4_i3;
  wire signed [`W-1:0] alu4_v;
  wire signed [`W-1:0] nots5_i0;
  wire signed [`W-1:0] nots5_i1;
  wire signed [`W-1:0] nots5_v;
  wire signed [`W-1:0] n600_i0;
  wire signed [`W-1:0] n600_i1;
  wire signed [`W-1:0] n600_i2;
  wire signed [`W-1:0] n600_i3;
  wire signed [`W-1:0] n600_i4;
  wire signed [`W-1:0] n600_v;
  wire signed [`W-1:0] n603_i0;
  wire signed [`W-1:0] n603_i1;
  wire signed [`W-1:0] n603_i2;
  wire signed [`W-1:0] n603_v;
  wire signed [`W-1:0] n1213_i0;
  wire signed [`W-1:0] n1213_i1;
  wire signed [`W-1:0] n1213_i2;
  wire signed [`W-1:0] n1213_v;
  wire signed [`W-1:0] n1205_i0;
  wire signed [`W-1:0] n1205_i1;
  wire signed [`W-1:0] n1205_i2;
  wire signed [`W-1:0] n1205_i3;
  wire signed [`W-1:0] n1205_v;
  wire signed [`W-1:0] op_T2_ind_y_i0;
  wire signed [`W-1:0] op_T2_ind_y_i1;
  wire signed [`W-1:0] op_T2_ind_y_i2;
  wire signed [`W-1:0] op_T2_ind_y_v;
  wire signed [`W-1:0] n1206_i0;
  wire signed [`W-1:0] n1206_i1;
  wire signed [`W-1:0] n1206_i2;
  wire signed [`W-1:0] n1206_i3;
  wire signed [`W-1:0] n1206_i4;
  wire signed [`W-1:0] n1206_v;
  wire signed [`W-1:0] n609_i0;
  wire signed [`W-1:0] n609_i1;
  wire signed [`W-1:0] n609_i2;
  wire signed [`W-1:0] n609_i3;
  wire signed [`W-1:0] n609_i4;
  wire signed [`W-1:0] n609_v;
  wire signed [`W-1:0] n608_i0;
  wire signed [`W-1:0] n608_i1;
  wire signed [`W-1:0] n608_i2;
  wire signed [`W-1:0] n608_v;
  wire signed [`W-1:0] n1202_i0;
  wire signed [`W-1:0] n1202_i1;
  wire signed [`W-1:0] n1202_i2;
  wire signed [`W-1:0] n1202_i3;
  wire signed [`W-1:0] n1202_v;
  wire signed [`W-1:0] n1560_i0;
  wire signed [`W-1:0] n1560_i1;
  wire signed [`W-1:0] n1560_i2;
  wire signed [`W-1:0] n1560_v;
  wire signed [`W-1:0] x0_i0;
  wire signed [`W-1:0] x0_i1;
  wire signed [`W-1:0] x0_i2;
  wire signed [`W-1:0] x0_v;
  wire signed [`W-1:0] n635_i0;
  wire signed [`W-1:0] n635_i1;
  wire signed [`W-1:0] n635_i2;
  wire signed [`W-1:0] n635_i3;
  wire signed [`W-1:0] n635_v;
  wire signed [`W-1:0] n636_i0;
  wire signed [`W-1:0] n636_i1;
  wire signed [`W-1:0] n636_i2;
  wire signed [`W-1:0] n636_v;
  wire signed [`W-1:0] n1215_i0;
  wire signed [`W-1:0] n1215_i1;
  wire signed [`W-1:0] n1215_i2;
  wire signed [`W-1:0] n1215_i3;
  wire signed [`W-1:0] n1215_v;
  wire signed [`W-1:0] n1447_i0;
  wire signed [`W-1:0] n1447_i1;
  wire signed [`W-1:0] n1447_v;
  wire signed [`W-1:0] n1446_i0;
  wire signed [`W-1:0] n1446_i1;
  wire signed [`W-1:0] n1446_i2;
  wire signed [`W-1:0] n1446_v;
  wire signed [`W-1:0] ir4_i0;
  wire signed [`W-1:0] ir4_i1;
  wire signed [`W-1:0] ir4_i2;
  wire signed [`W-1:0] ir4_i3;
  wire signed [`W-1:0] ir4_i4;
  wire signed [`W-1:0] ir4_i5;
  wire signed [`W-1:0] ir4_i6;
  wire signed [`W-1:0] ir4_i7;
  wire signed [`W-1:0] ir4_i8;
  wire signed [`W-1:0] ir4_i9;
  wire signed [`W-1:0] ir4_i10;
  wire signed [`W-1:0] ir4_i11;
  wire signed [`W-1:0] ir4_i12;
  wire signed [`W-1:0] ir4_i13;
  wire signed [`W-1:0] ir4_i14;
  wire signed [`W-1:0] ir4_i15;
  wire signed [`W-1:0] ir4_i16;
  wire signed [`W-1:0] ir4_i17;
  wire signed [`W-1:0] ir4_i18;
  wire signed [`W-1:0] ir4_i19;
  wire signed [`W-1:0] ir4_i20;
  wire signed [`W-1:0] ir4_i21;
  wire signed [`W-1:0] ir4_i22;
  wire signed [`W-1:0] ir4_i23;
  wire signed [`W-1:0] ir4_i24;
  wire signed [`W-1:0] ir4_i25;
  wire signed [`W-1:0] ir4_i26;
  wire signed [`W-1:0] ir4_i27;
  wire signed [`W-1:0] ir4_i28;
  wire signed [`W-1:0] ir4_i29;
  wire signed [`W-1:0] ir4_i30;
  wire signed [`W-1:0] ir4_i31;
  wire signed [`W-1:0] ir4_i32;
  wire signed [`W-1:0] ir4_i33;
  wire signed [`W-1:0] ir4_i34;
  wire signed [`W-1:0] ir4_i35;
  wire signed [`W-1:0] ir4_i36;
  wire signed [`W-1:0] ir4_i37;
  wire signed [`W-1:0] ir4_i38;
  wire signed [`W-1:0] ir4_i39;
  wire signed [`W-1:0] ir4_i40;
  wire signed [`W-1:0] ir4_i41;
  wire signed [`W-1:0] ir4_i42;
  wire signed [`W-1:0] ir4_i43;
  wire signed [`W-1:0] ir4_i44;
  wire signed [`W-1:0] ir4_i45;
  wire signed [`W-1:0] ir4_i46;
  wire signed [`W-1:0] ir4_i47;
  wire signed [`W-1:0] ir4_i48;
  wire signed [`W-1:0] ir4_i49;
  wire signed [`W-1:0] ir4_i50;
  wire signed [`W-1:0] ir4_i51;
  wire signed [`W-1:0] ir4_i52;
  wire signed [`W-1:0] ir4_i53;
  wire signed [`W-1:0] ir4_i54;
  wire signed [`W-1:0] ir4_i55;
  wire signed [`W-1:0] ir4_i56;
  wire signed [`W-1:0] ir4_i57;
  wire signed [`W-1:0] ir4_i58;
  wire signed [`W-1:0] ir4_i59;
  wire signed [`W-1:0] ir4_i60;
  wire signed [`W-1:0] ir4_i61;
  wire signed [`W-1:0] ir4_i62;
  wire signed [`W-1:0] ir4_i63;
  wire signed [`W-1:0] ir4_i64;
  wire signed [`W-1:0] ir4_i65;
  wire signed [`W-1:0] ir4_i66;
  wire signed [`W-1:0] ir4_i67;
  wire signed [`W-1:0] ir4_i68;
  wire signed [`W-1:0] ir4_i69;
  wire signed [`W-1:0] ir4_i70;
  wire signed [`W-1:0] ir4_v;
  wire signed [`W-1:0] ab10_i0;
  wire signed [`W-1:0] ab10_i1;
  wire signed [`W-1:0] ab10_i2;
  wire signed [`W-1:0] ab10_v;
  wire signed [`W-1:0] pipeUNK13_i0;
  wire signed [`W-1:0] pipeUNK13_i1;
  wire signed [`W-1:0] pipeUNK13_v;
  wire signed [`W-1:0] n1117_i0;
  wire signed [`W-1:0] n1117_i1;
  wire signed [`W-1:0] n1117_i2;
  wire signed [`W-1:0] n1117_v;
  wire signed [`W-1:0] idl6_i0;
  wire signed [`W-1:0] idl6_i1;
  wire signed [`W-1:0] idl6_i2;
  wire signed [`W-1:0] idl6_v;
  wire signed [`W-1:0] Pout4_i0;
  wire signed [`W-1:0] Pout4_i1;
  wire signed [`W-1:0] Pout4_i2;
  wire signed [`W-1:0] Pout4_v;
  wire signed [`W-1:0] n1449_i0;
  wire signed [`W-1:0] n1449_i1;
  wire signed [`W-1:0] n1449_i2;
  wire signed [`W-1:0] n1449_v;
  wire signed [`W-1:0] n1448_i0;
  wire signed [`W-1:0] n1448_i1;
  wire signed [`W-1:0] n1448_i2;
  wire signed [`W-1:0] n1448_v;
  wire signed [`W-1:0] n1219_i0;
  wire signed [`W-1:0] n1219_i1;
  wire signed [`W-1:0] n1219_i2;
  wire signed [`W-1:0] n1219_v;
  wire signed [`W-1:0] x_op_T4_ind_y_i0;
  wire signed [`W-1:0] x_op_T4_ind_y_i1;
  wire signed [`W-1:0] x_op_T4_ind_y_i2;
  wire signed [`W-1:0] x_op_T4_ind_y_i3;
  wire signed [`W-1:0] x_op_T4_ind_y_v;
  wire signed [`W-1:0] n460_i0;
  wire signed [`W-1:0] n460_i1;
  wire signed [`W-1:0] n460_v;
  wire signed [`W-1:0] abh7_i0;
  wire signed [`W-1:0] abh7_i1;
  wire signed [`W-1:0] abh7_i2;
  wire signed [`W-1:0] abh7_i3;
  wire signed [`W-1:0] abh7_i4;
  wire signed [`W-1:0] abh7_v;
  wire signed [`W-1:0] n488_i0;
  wire signed [`W-1:0] n488_i1;
  wire signed [`W-1:0] n488_i2;
  wire signed [`W-1:0] n488_i3;
  wire signed [`W-1:0] n488_i4;
  wire signed [`W-1:0] n488_v;
  wire signed [`W-1:0] op_T2_brk_i0;
  wire signed [`W-1:0] op_T2_brk_i1;
  wire signed [`W-1:0] op_T2_brk_i2;
  wire signed [`W-1:0] op_T2_brk_v;
  wire signed [`W-1:0] __AxBxC_5_i0;
  wire signed [`W-1:0] __AxBxC_5_i1;
  wire signed [`W-1:0] __AxBxC_5_i2;
  wire signed [`W-1:0] __AxBxC_5_v;
  wire signed [`W-1:0] n485_i0;
  wire signed [`W-1:0] n485_i1;
  wire signed [`W-1:0] n485_i2;
  wire signed [`W-1:0] n485_v;
  wire signed [`W-1:0] n484_i0;
  wire signed [`W-1:0] n484_i1;
  wire signed [`W-1:0] n484_i2;
  wire signed [`W-1:0] n484_v;
  wire signed [`W-1:0] adh5_i0;
  wire signed [`W-1:0] adh5_i1;
  wire signed [`W-1:0] adh5_i2;
  wire signed [`W-1:0] adh5_i3;
  wire signed [`W-1:0] adh5_i4;
  wire signed [`W-1:0] adh5_i5;
  wire signed [`W-1:0] adh5_i6;
  wire signed [`W-1:0] adh5_v;
  wire signed [`W-1:0] n481_i0;
  wire signed [`W-1:0] n481_i1;
  wire signed [`W-1:0] n481_i2;
  wire signed [`W-1:0] n481_i3;
  wire signed [`W-1:0] n481_i4;
  wire signed [`W-1:0] n481_v;
  wire signed [`W-1:0] n480_i0;
  wire signed [`W-1:0] n480_i1;
  wire signed [`W-1:0] n480_i2;
  wire signed [`W-1:0] n480_v;
  wire signed [`W-1:0] pipeUNK09_i0;
  wire signed [`W-1:0] pipeUNK09_i1;
  wire signed [`W-1:0] pipeUNK09_i2;
  wire signed [`W-1:0] pipeUNK09_i3;
  wire signed [`W-1:0] pipeUNK09_v;
  wire signed [`W-1:0] n198_i0;
  wire signed [`W-1:0] n198_i1;
  wire signed [`W-1:0] n198_i2;
  wire signed [`W-1:0] n198_i3;
  wire signed [`W-1:0] n198_v;
  wire signed [`W-1:0] ab15_i0;
  wire signed [`W-1:0] ab15_i1;
  wire signed [`W-1:0] ab15_i2;
  wire signed [`W-1:0] ab15_v;
  wire signed [`W-1:0] notir0_i0;
  wire signed [`W-1:0] notir0_i1;
  wire signed [`W-1:0] notir0_i2;
  wire signed [`W-1:0] notir0_i3;
  wire signed [`W-1:0] notir0_i4;
  wire signed [`W-1:0] notir0_i5;
  wire signed [`W-1:0] notir0_i6;
  wire signed [`W-1:0] notir0_i7;
  wire signed [`W-1:0] notir0_i8;
  wire signed [`W-1:0] notir0_i9;
  wire signed [`W-1:0] notir0_i10;
  wire signed [`W-1:0] notir0_i11;
  wire signed [`W-1:0] notir0_i12;
  wire signed [`W-1:0] notir0_i13;
  wire signed [`W-1:0] notir0_i14;
  wire signed [`W-1:0] notir0_i15;
  wire signed [`W-1:0] notir0_i16;
  wire signed [`W-1:0] notir0_i17;
  wire signed [`W-1:0] notir0_i18;
  wire signed [`W-1:0] notir0_i19;
  wire signed [`W-1:0] notir0_i20;
  wire signed [`W-1:0] notir0_i21;
  wire signed [`W-1:0] notir0_i22;
  wire signed [`W-1:0] notir0_i23;
  wire signed [`W-1:0] notir0_i24;
  wire signed [`W-1:0] notir0_i25;
  wire signed [`W-1:0] notir0_i26;
  wire signed [`W-1:0] notir0_i27;
  wire signed [`W-1:0] notir0_i28;
  wire signed [`W-1:0] notir0_v;
  wire signed [`W-1:0] pipeUNK37_i0;
  wire signed [`W-1:0] pipeUNK37_i1;
  wire signed [`W-1:0] pipeUNK37_v;
  wire signed [`W-1:0] n196_i0;
  wire signed [`W-1:0] n196_i1;
  wire signed [`W-1:0] n196_i2;
  wire signed [`W-1:0] n196_v;
  wire signed [`W-1:0] n191_i0;
  wire signed [`W-1:0] n191_i1;
  wire signed [`W-1:0] n191_i2;
  wire signed [`W-1:0] n191_v;
  wire signed [`W-1:0] n190_i0;
  wire signed [`W-1:0] n190_i1;
  wire signed [`W-1:0] n190_v;
  wire signed [`W-1:0] _AxB_2__C12_i0;
  wire signed [`W-1:0] _AxB_2__C12_i1;
  wire signed [`W-1:0] _AxB_2__C12_i2;
  wire signed [`W-1:0] _AxB_2__C12_v;
  wire signed [`W-1:0] n192_i0;
  wire signed [`W-1:0] n192_i1;
  wire signed [`W-1:0] n192_i2;
  wire signed [`W-1:0] n192_i3;
  wire signed [`W-1:0] n192_i4;
  wire signed [`W-1:0] n192_v;
  wire signed [`W-1:0] n1106_i0;
  wire signed [`W-1:0] n1106_i1;
  wire signed [`W-1:0] n1106_i2;
  wire signed [`W-1:0] n1106_v;
  wire signed [`W-1:0] n1455_i0;
  wire signed [`W-1:0] n1455_i1;
  wire signed [`W-1:0] n1455_i2;
  wire signed [`W-1:0] n1455_i3;
  wire signed [`W-1:0] n1455_v;
  wire signed [`W-1:0] n1274_i0;
  wire signed [`W-1:0] n1274_i1;
  wire signed [`W-1:0] n1274_v;
  wire signed [`W-1:0] n1457_i0;
  wire signed [`W-1:0] n1457_i1;
  wire signed [`W-1:0] n1457_i2;
  wire signed [`W-1:0] n1457_v;
  wire signed [`W-1:0] pclp1_i0;
  wire signed [`W-1:0] pclp1_i1;
  wire signed [`W-1:0] pclp1_v;
  wire signed [`W-1:0] n1100_i0;
  wire signed [`W-1:0] n1100_i1;
  wire signed [`W-1:0] n1100_i2;
  wire signed [`W-1:0] n1100_i3;
  wire signed [`W-1:0] n1100_v;
  wire signed [`W-1:0] n1101_i0;
  wire signed [`W-1:0] n1101_i1;
  wire signed [`W-1:0] n1101_i2;
  wire signed [`W-1:0] n1101_v;
  wire signed [`W-1:0] n902_i0;
  wire signed [`W-1:0] n902_i1;
  wire signed [`W-1:0] n902_i2;
  wire signed [`W-1:0] n902_v;
  wire signed [`W-1:0] pcl4_i0;
  wire signed [`W-1:0] pcl4_i1;
  wire signed [`W-1:0] pcl4_i2;
  wire signed [`W-1:0] pcl4_v;
  wire signed [`W-1:0] _DA_ADD1_i0;
  wire signed [`W-1:0] _DA_ADD1_i1;
  wire signed [`W-1:0] _DA_ADD1_i2;
  wire signed [`W-1:0] _DA_ADD1_i3;
  wire signed [`W-1:0] _DA_ADD1_i4;
  wire signed [`W-1:0] _DA_ADD1_i5;
  wire signed [`W-1:0] _DA_ADD1_v;
  wire signed [`W-1:0] n906_i0;
  wire signed [`W-1:0] n906_i1;
  wire signed [`W-1:0] n906_i2;
  wire signed [`W-1:0] n906_i3;
  wire signed [`W-1:0] n906_v;
  wire signed [`W-1:0] _ABH1_i0;
  wire signed [`W-1:0] _ABH1_i1;
  wire signed [`W-1:0] _ABH1_i2;
  wire signed [`W-1:0] _ABH1_v;
  wire signed [`W-1:0] op_T3_mem_zp_idx_i0;
  wire signed [`W-1:0] op_T3_mem_zp_idx_i1;
  wire signed [`W-1:0] op_T3_mem_zp_idx_i2;
  wire signed [`W-1:0] op_T3_mem_zp_idx_v;
  wire signed [`W-1:0] n905_i0;
  wire signed [`W-1:0] n905_i1;
  wire signed [`W-1:0] n905_i2;
  wire signed [`W-1:0] n905_v;
  wire signed [`W-1:0] n420_i0;
  wire signed [`W-1:0] n420_i1;
  wire signed [`W-1:0] n420_i2;
  wire signed [`W-1:0] n420_v;
  wire signed [`W-1:0] t5_i0;
  wire signed [`W-1:0] t5_i1;
  wire signed [`W-1:0] t5_i2;
  wire signed [`W-1:0] t5_i3;
  wire signed [`W-1:0] t5_i4;
  wire signed [`W-1:0] t5_i5;
  wire signed [`W-1:0] t5_i6;
  wire signed [`W-1:0] t5_i7;
  wire signed [`W-1:0] t5_i8;
  wire signed [`W-1:0] t5_i9;
  wire signed [`W-1:0] t5_i10;
  wire signed [`W-1:0] t5_v;
  wire signed [`W-1:0] n854_i0;
  wire signed [`W-1:0] n854_i1;
  wire signed [`W-1:0] n854_i2;
  wire signed [`W-1:0] n854_i3;
  wire signed [`W-1:0] n854_v;
  wire signed [`W-1:0] n855_i0;
  wire signed [`W-1:0] n855_i1;
  wire signed [`W-1:0] n855_i2;
  wire signed [`W-1:0] n855_v;
  wire signed [`W-1:0] op_rti_rts_i0;
  wire signed [`W-1:0] op_rti_rts_i1;
  wire signed [`W-1:0] op_rti_rts_i2;
  wire signed [`W-1:0] op_rti_rts_i3;
  wire signed [`W-1:0] op_rti_rts_i4;
  wire signed [`W-1:0] op_rti_rts_v;
  wire signed [`W-1:0] n850_i0;
  wire signed [`W-1:0] n850_i1;
  wire signed [`W-1:0] n850_i2;
  wire signed [`W-1:0] n850_i3;
  wire signed [`W-1:0] n850_v;
  wire signed [`W-1:0] abh3_i0;
  wire signed [`W-1:0] abh3_i1;
  wire signed [`W-1:0] abh3_i2;
  wire signed [`W-1:0] abh3_i3;
  wire signed [`W-1:0] abh3_i4;
  wire signed [`W-1:0] abh3_v;
  wire signed [`W-1:0] n852_i0;
  wire signed [`W-1:0] n852_i1;
  wire signed [`W-1:0] n852_i2;
  wire signed [`W-1:0] n852_i3;
  wire signed [`W-1:0] n852_v;
  wire signed [`W-1:0] op_T5_rts_i0;
  wire signed [`W-1:0] op_T5_rts_i1;
  wire signed [`W-1:0] op_T5_rts_i2;
  wire signed [`W-1:0] op_T5_rts_i3;
  wire signed [`W-1:0] op_T5_rts_i4;
  wire signed [`W-1:0] op_T5_rts_i5;
  wire signed [`W-1:0] op_T5_rts_v;
  wire signed [`W-1:0] a5_i0;
  wire signed [`W-1:0] a5_i1;
  wire signed [`W-1:0] a5_i2;
  wire signed [`W-1:0] a5_v;
  wire signed [`W-1:0] dpc9_DBADD_i0;
  wire signed [`W-1:0] dpc9_DBADD_i1;
  wire signed [`W-1:0] dpc9_DBADD_i2;
  wire signed [`W-1:0] dpc9_DBADD_i3;
  wire signed [`W-1:0] dpc9_DBADD_i4;
  wire signed [`W-1:0] dpc9_DBADD_i5;
  wire signed [`W-1:0] dpc9_DBADD_i6;
  wire signed [`W-1:0] dpc9_DBADD_i7;
  wire signed [`W-1:0] dpc9_DBADD_i8;
  wire signed [`W-1:0] dpc9_DBADD_i9;
  wire signed [`W-1:0] dpc9_DBADD_v;
  wire signed [`W-1:0] n6_i0;
  wire signed [`W-1:0] n6_i1;
  wire signed [`W-1:0] n6_i2;
  wire signed [`W-1:0] n6_i3;
  wire signed [`W-1:0] n6_v;
  wire signed [`W-1:0] AxB1_i0;
  wire signed [`W-1:0] AxB1_i1;
  wire signed [`W-1:0] AxB1_i2;
  wire signed [`W-1:0] AxB1_i3;
  wire signed [`W-1:0] AxB1_i4;
  wire signed [`W-1:0] AxB1_i5;
  wire signed [`W-1:0] AxB1_v;
  wire signed [`W-1:0] n611_i0;
  wire signed [`W-1:0] n611_i1;
  wire signed [`W-1:0] n611_i2;
  wire signed [`W-1:0] n611_i3;
  wire signed [`W-1:0] n611_v;
  wire signed [`W-1:0] n740_i0;
  wire signed [`W-1:0] n740_i1;
  wire signed [`W-1:0] n740_i2;
  wire signed [`W-1:0] n740_i3;
  wire signed [`W-1:0] n740_i4;
  wire signed [`W-1:0] n740_i5;
  wire signed [`W-1:0] n740_v;
  wire signed [`W-1:0] dpc31_PCHPCH_i0;
  wire signed [`W-1:0] dpc31_PCHPCH_i1;
  wire signed [`W-1:0] dpc31_PCHPCH_i2;
  wire signed [`W-1:0] dpc31_PCHPCH_i3;
  wire signed [`W-1:0] dpc31_PCHPCH_i4;
  wire signed [`W-1:0] dpc31_PCHPCH_i5;
  wire signed [`W-1:0] dpc31_PCHPCH_i6;
  wire signed [`W-1:0] dpc31_PCHPCH_i7;
  wire signed [`W-1:0] dpc31_PCHPCH_i8;
  wire signed [`W-1:0] dpc31_PCHPCH_i9;
  wire signed [`W-1:0] dpc31_PCHPCH_v;
  wire signed [`W-1:0] n743_i0;
  wire signed [`W-1:0] n743_i1;
  wire signed [`W-1:0] n743_i2;
  wire signed [`W-1:0] n743_i3;
  wire signed [`W-1:0] n743_i4;
  wire signed [`W-1:0] n743_v;
  wire signed [`W-1:0] DBZ_i0;
  wire signed [`W-1:0] DBZ_i1;
  wire signed [`W-1:0] DBZ_i2;
  wire signed [`W-1:0] DBZ_v;
  wire signed [`W-1:0] n745_i0;
  wire signed [`W-1:0] n745_i1;
  wire signed [`W-1:0] n745_v;
  wire signed [`W-1:0] dor1_i0;
  wire signed [`W-1:0] dor1_i1;
  wire signed [`W-1:0] dor1_i2;
  wire signed [`W-1:0] dor1_i3;
  wire signed [`W-1:0] dor1_i4;
  wire signed [`W-1:0] dor1_v;
  wire signed [`W-1:0] n747_i0;
  wire signed [`W-1:0] n747_i1;
  wire signed [`W-1:0] n747_i2;
  wire signed [`W-1:0] n747_i3;
  wire signed [`W-1:0] n747_v;
  wire signed [`W-1:0] n748_i0;
  wire signed [`W-1:0] n748_i1;
  wire signed [`W-1:0] n748_i2;
  wire signed [`W-1:0] n748_i3;
  wire signed [`W-1:0] n748_v;
  wire signed [`W-1:0] n617_i0;
  wire signed [`W-1:0] n617_i1;
  wire signed [`W-1:0] n617_i2;
  wire signed [`W-1:0] n617_i3;
  wire signed [`W-1:0] n617_v;
  wire signed [`W-1:0] x_op_push_pull_i0;
  wire signed [`W-1:0] x_op_push_pull_i1;
  wire signed [`W-1:0] x_op_push_pull_i2;
  wire signed [`W-1:0] x_op_push_pull_v;
  wire signed [`W-1:0] pipeUNK16_i0;
  wire signed [`W-1:0] pipeUNK16_i1;
  wire signed [`W-1:0] pipeUNK16_v;
  wire signed [`W-1:0] x_op_jmp_i0;
  wire signed [`W-1:0] x_op_jmp_i1;
  wire signed [`W-1:0] x_op_jmp_i2;
  wire signed [`W-1:0] x_op_jmp_i3;
  wire signed [`W-1:0] x_op_jmp_v;
  wire signed [`W-1:0] n1054_i0;
  wire signed [`W-1:0] n1054_i1;
  wire signed [`W-1:0] n1054_i2;
  wire signed [`W-1:0] n1054_v;
  wire signed [`W-1:0] n1055_i0;
  wire signed [`W-1:0] n1055_i1;
  wire signed [`W-1:0] n1055_i2;
  wire signed [`W-1:0] n1055_v;
  wire signed [`W-1:0] n1056_i0;
  wire signed [`W-1:0] n1056_i1;
  wire signed [`W-1:0] n1056_i2;
  wire signed [`W-1:0] n1056_v;
  wire signed [`W-1:0] op_T2_abs_i0;
  wire signed [`W-1:0] op_T2_abs_i1;
  wire signed [`W-1:0] op_T2_abs_i2;
  wire signed [`W-1:0] op_T2_abs_v;
  wire signed [`W-1:0] n1059_i0;
  wire signed [`W-1:0] n1059_v;
  wire signed [`W-1:0] n1696_i0;
  wire signed [`W-1:0] n1696_i1;
  wire signed [`W-1:0] n1696_i2;
  wire signed [`W-1:0] n1696_v;
  wire signed [`W-1:0] n1697_i0;
  wire signed [`W-1:0] n1697_i1;
  wire signed [`W-1:0] n1697_i2;
  wire signed [`W-1:0] n1697_v;
  wire signed [`W-1:0] n1694_i0;
  wire signed [`W-1:0] n1694_i1;
  wire signed [`W-1:0] n1694_i2;
  wire signed [`W-1:0] n1694_i3;
  wire signed [`W-1:0] n1694_v;
  wire signed [`W-1:0] n1693_i0;
  wire signed [`W-1:0] n1693_i1;
  wire signed [`W-1:0] n1693_v;
  wire signed [`W-1:0] pd7_i0;
  wire signed [`W-1:0] pd7_i1;
  wire signed [`W-1:0] pd7_v;
  wire signed [`W-1:0] n1691_i0;
  wire signed [`W-1:0] n1691_i1;
  wire signed [`W-1:0] n1691_i2;
  wire signed [`W-1:0] n1691_i3;
  wire signed [`W-1:0] n1691_i4;
  wire signed [`W-1:0] n1691_i5;
  wire signed [`W-1:0] n1691_i6;
  wire signed [`W-1:0] n1691_v;
  wire signed [`W-1:0] dpc24_ACSB_i0;
  wire signed [`W-1:0] dpc24_ACSB_i1;
  wire signed [`W-1:0] dpc24_ACSB_i2;
  wire signed [`W-1:0] dpc24_ACSB_i3;
  wire signed [`W-1:0] dpc24_ACSB_i4;
  wire signed [`W-1:0] dpc24_ACSB_i5;
  wire signed [`W-1:0] dpc24_ACSB_i6;
  wire signed [`W-1:0] dpc24_ACSB_i7;
  wire signed [`W-1:0] dpc24_ACSB_i8;
  wire signed [`W-1:0] dpc24_ACSB_i9;
  wire signed [`W-1:0] dpc24_ACSB_v;
  wire signed [`W-1:0] n1699_i0;
  wire signed [`W-1:0] n1699_i1;
  wire signed [`W-1:0] n1699_v;
  wire signed [`W-1:0] n618_i0;
  wire signed [`W-1:0] n618_i1;
  wire signed [`W-1:0] n618_i2;
  wire signed [`W-1:0] n618_i3;
  wire signed [`W-1:0] n618_i4;
  wire signed [`W-1:0] n618_v;
  wire signed [`W-1:0] n612_i0;
  wire signed [`W-1:0] n612_i1;
  wire signed [`W-1:0] n612_i2;
  wire signed [`W-1:0] n612_v;
  wire signed [`W-1:0] n613_i0;
  wire signed [`W-1:0] n613_i1;
  wire signed [`W-1:0] n613_i2;
  wire signed [`W-1:0] n613_i3;
  wire signed [`W-1:0] n613_v;
  wire signed [`W-1:0] n1272_i0;
  wire signed [`W-1:0] n1272_i1;
  wire signed [`W-1:0] n1272_v;
  wire signed [`W-1:0] op_T0_i0;
  wire signed [`W-1:0] op_T0_i1;
  wire signed [`W-1:0] op_T0_i2;
  wire signed [`W-1:0] op_T0_v;
  wire signed [`W-1:0] n616_i0;
  wire signed [`W-1:0] n616_i1;
  wire signed [`W-1:0] n616_i2;
  wire signed [`W-1:0] n616_i3;
  wire signed [`W-1:0] n616_v;
  wire signed [`W-1:0] n1275_i0;
  wire signed [`W-1:0] n1275_i1;
  wire signed [`W-1:0] n1275_i2;
  wire signed [`W-1:0] n1275_v;
  wire signed [`W-1:0] pipeUNK31_i0;
  wire signed [`W-1:0] pipeUNK31_i1;
  wire signed [`W-1:0] pipeUNK31_v;
  wire signed [`W-1:0] y5_i0;
  wire signed [`W-1:0] y5_i1;
  wire signed [`W-1:0] y5_i2;
  wire signed [`W-1:0] y5_v;
  wire signed [`W-1:0] n1472_i0;
  wire signed [`W-1:0] n1472_i1;
  wire signed [`W-1:0] n1472_v;
  wire signed [`W-1:0] idb2_i0;
  wire signed [`W-1:0] idb2_i1;
  wire signed [`W-1:0] idb2_i2;
  wire signed [`W-1:0] idb2_i3;
  wire signed [`W-1:0] idb2_i4;
  wire signed [`W-1:0] idb2_i5;
  wire signed [`W-1:0] idb2_i6;
  wire signed [`W-1:0] idb2_i7;
  wire signed [`W-1:0] idb2_i8;
  wire signed [`W-1:0] idb2_i9;
  wire signed [`W-1:0] idb2_i10;
  wire signed [`W-1:0] idb2_i11;
  wire signed [`W-1:0] idb2_v;
  wire signed [`W-1:0] n1471_i0;
  wire signed [`W-1:0] n1471_i1;
  wire signed [`W-1:0] n1471_i2;
  wire signed [`W-1:0] n1471_v;
  wire signed [`W-1:0] x_op_T0_bit_i0;
  wire signed [`W-1:0] x_op_T0_bit_i1;
  wire signed [`W-1:0] x_op_T0_bit_i2;
  wire signed [`W-1:0] x_op_T0_bit_v;
  wire signed [`W-1:0] n1477_i0;
  wire signed [`W-1:0] n1477_i1;
  wire signed [`W-1:0] n1477_v;
  wire signed [`W-1:0] n1474_i0;
  wire signed [`W-1:0] n1474_i1;
  wire signed [`W-1:0] n1474_i2;
  wire signed [`W-1:0] n1474_v;
  wire signed [`W-1:0] dasb3_i0;
  wire signed [`W-1:0] dasb3_i1;
  wire signed [`W-1:0] dasb3_i2;
  wire signed [`W-1:0] dasb3_v;
  wire signed [`W-1:0] op_T0_brk_rti_i0;
  wire signed [`W-1:0] op_T0_brk_rti_i1;
  wire signed [`W-1:0] op_T0_brk_rti_i2;
  wire signed [`W-1:0] op_T0_brk_rti_v;
  wire signed [`W-1:0] n1479_i0;
  wire signed [`W-1:0] n1479_i1;
  wire signed [`W-1:0] n1479_i2;
  wire signed [`W-1:0] n1479_v;
  wire signed [`W-1:0] n1304_i0;
  wire signed [`W-1:0] n1304_i1;
  wire signed [`W-1:0] n1304_i2;
  wire signed [`W-1:0] n1304_v;
  wire signed [`W-1:0] n1305_i0;
  wire signed [`W-1:0] n1305_i1;
  wire signed [`W-1:0] n1305_i2;
  wire signed [`W-1:0] n1305_v;
  wire signed [`W-1:0] idl4_i0;
  wire signed [`W-1:0] idl4_i1;
  wire signed [`W-1:0] idl4_i2;
  wire signed [`W-1:0] idl4_v;
  wire signed [`W-1:0] _ABL6_i0;
  wire signed [`W-1:0] _ABL6_i1;
  wire signed [`W-1:0] _ABL6_i2;
  wire signed [`W-1:0] _ABL6_v;
  wire signed [`W-1:0] n1300_i0;
  wire signed [`W-1:0] n1300_i1;
  wire signed [`W-1:0] n1300_i2;
  wire signed [`W-1:0] n1300_v;
  wire signed [`W-1:0] n1301_i0;
  wire signed [`W-1:0] n1301_i1;
  wire signed [`W-1:0] n1301_i2;
  wire signed [`W-1:0] n1301_i3;
  wire signed [`W-1:0] n1301_i4;
  wire signed [`W-1:0] n1301_v;
  wire signed [`W-1:0] idb3_i0;
  wire signed [`W-1:0] idb3_i1;
  wire signed [`W-1:0] idb3_i2;
  wire signed [`W-1:0] idb3_i3;
  wire signed [`W-1:0] idb3_i4;
  wire signed [`W-1:0] idb3_i5;
  wire signed [`W-1:0] idb3_i6;
  wire signed [`W-1:0] idb3_i7;
  wire signed [`W-1:0] idb3_i8;
  wire signed [`W-1:0] idb3_i9;
  wire signed [`W-1:0] idb3_i10;
  wire signed [`W-1:0] idb3_i11;
  wire signed [`W-1:0] idb3_v;
  wire signed [`W-1:0] n1303_i0;
  wire signed [`W-1:0] n1303_i1;
  wire signed [`W-1:0] n1303_i2;
  wire signed [`W-1:0] n1303_v;
  wire signed [`W-1:0] notaluvout_i0;
  wire signed [`W-1:0] notaluvout_i1;
  wire signed [`W-1:0] notaluvout_i2;
  wire signed [`W-1:0] notaluvout_v;
  wire signed [`W-1:0] n1309_i0;
  wire signed [`W-1:0] n1309_i1;
  wire signed [`W-1:0] n1309_i2;
  wire signed [`W-1:0] n1309_v;
  wire signed [`W-1:0] notidl5_i0;
  wire signed [`W-1:0] notidl5_i1;
  wire signed [`W-1:0] notidl5_v;
  wire signed [`W-1:0] n499_i0;
  wire signed [`W-1:0] n499_i1;
  wire signed [`W-1:0] n499_i2;
  wire signed [`W-1:0] n499_i3;
  wire signed [`W-1:0] n499_v;
  wire signed [`W-1:0] n494_i0;
  wire signed [`W-1:0] n494_i1;
  wire signed [`W-1:0] n494_i2;
  wire signed [`W-1:0] n494_v;
  wire signed [`W-1:0] notalu3_i0;
  wire signed [`W-1:0] notalu3_i1;
  wire signed [`W-1:0] notalu3_v;
  wire signed [`W-1:0] n496_i0;
  wire signed [`W-1:0] n496_i1;
  wire signed [`W-1:0] n496_i2;
  wire signed [`W-1:0] n496_v;
  wire signed [`W-1:0] n490_i0;
  wire signed [`W-1:0] n490_i1;
  wire signed [`W-1:0] n490_i2;
  wire signed [`W-1:0] n490_v;
  wire signed [`W-1:0] n491_i0;
  wire signed [`W-1:0] n491_i1;
  wire signed [`W-1:0] n491_i2;
  wire signed [`W-1:0] n491_v;
  wire signed [`W-1:0] op_T4_ind_y_i0;
  wire signed [`W-1:0] op_T4_ind_y_i1;
  wire signed [`W-1:0] op_T4_ind_y_i2;
  wire signed [`W-1:0] op_T4_ind_y_v;
  wire signed [`W-1:0] idb7_i0;
  wire signed [`W-1:0] idb7_i1;
  wire signed [`W-1:0] idb7_i2;
  wire signed [`W-1:0] idb7_i3;
  wire signed [`W-1:0] idb7_i4;
  wire signed [`W-1:0] idb7_i5;
  wire signed [`W-1:0] idb7_i6;
  wire signed [`W-1:0] idb7_i7;
  wire signed [`W-1:0] idb7_i8;
  wire signed [`W-1:0] idb7_i9;
  wire signed [`W-1:0] idb7_i10;
  wire signed [`W-1:0] idb7_i11;
  wire signed [`W-1:0] idb7_v;
  wire signed [`W-1:0] n24_i0;
  wire signed [`W-1:0] n24_i1;
  wire signed [`W-1:0] n24_v;
  wire signed [`W-1:0] n25_i0;
  wire signed [`W-1:0] n25_i1;
  wire signed [`W-1:0] n25_i2;
  wire signed [`W-1:0] n25_v;
  wire signed [`W-1:0] notir4_i0;
  wire signed [`W-1:0] notir4_i1;
  wire signed [`W-1:0] notir4_i2;
  wire signed [`W-1:0] notir4_i3;
  wire signed [`W-1:0] notir4_i4;
  wire signed [`W-1:0] notir4_i5;
  wire signed [`W-1:0] notir4_i6;
  wire signed [`W-1:0] notir4_i7;
  wire signed [`W-1:0] notir4_i8;
  wire signed [`W-1:0] notir4_i9;
  wire signed [`W-1:0] notir4_i10;
  wire signed [`W-1:0] notir4_i11;
  wire signed [`W-1:0] notir4_i12;
  wire signed [`W-1:0] notir4_i13;
  wire signed [`W-1:0] notir4_i14;
  wire signed [`W-1:0] notir4_i15;
  wire signed [`W-1:0] notir4_i16;
  wire signed [`W-1:0] notir4_i17;
  wire signed [`W-1:0] notir4_i18;
  wire signed [`W-1:0] notir4_i19;
  wire signed [`W-1:0] notir4_i20;
  wire signed [`W-1:0] notir4_i21;
  wire signed [`W-1:0] notir4_i22;
  wire signed [`W-1:0] notir4_i23;
  wire signed [`W-1:0] notir4_i24;
  wire signed [`W-1:0] notir4_i25;
  wire signed [`W-1:0] notir4_i26;
  wire signed [`W-1:0] notir4_v;
  wire signed [`W-1:0] n27_i0;
  wire signed [`W-1:0] n27_i1;
  wire signed [`W-1:0] n27_i2;
  wire signed [`W-1:0] n27_i3;
  wire signed [`W-1:0] n27_i4;
  wire signed [`W-1:0] n27_v;
  wire signed [`W-1:0] n20_i0;
  wire signed [`W-1:0] n20_i1;
  wire signed [`W-1:0] n20_i2;
  wire signed [`W-1:0] n20_v;
  wire signed [`W-1:0] n21_i0;
  wire signed [`W-1:0] n21_i1;
  wire signed [`W-1:0] n21_i2;
  wire signed [`W-1:0] n21_i3;
  wire signed [`W-1:0] n21_v;
  wire signed [`W-1:0] __AxBxC_2_i0;
  wire signed [`W-1:0] __AxBxC_2_i1;
  wire signed [`W-1:0] __AxBxC_2_i2;
  wire signed [`W-1:0] __AxBxC_2_v;
  wire signed [`W-1:0] n23_i0;
  wire signed [`W-1:0] n23_i1;
  wire signed [`W-1:0] n23_i2;
  wire signed [`W-1:0] n23_i3;
  wire signed [`W-1:0] n23_v;
  wire signed [`W-1:0] _ABL7_i0;
  wire signed [`W-1:0] _ABL7_i1;
  wire signed [`W-1:0] _ABL7_i2;
  wire signed [`W-1:0] _ABL7_v;
  wire signed [`W-1:0] n29_i0;
  wire signed [`W-1:0] n29_i1;
  wire signed [`W-1:0] n29_i2;
  wire signed [`W-1:0] n29_v;
  wire signed [`W-1:0] n7_i0;
  wire signed [`W-1:0] n7_i1;
  wire signed [`W-1:0] n7_i2;
  wire signed [`W-1:0] n7_v;
  wire signed [`W-1:0] n410_i0;
  wire signed [`W-1:0] n410_i1;
  wire signed [`W-1:0] n410_i2;
  wire signed [`W-1:0] n410_i3;
  wire signed [`W-1:0] n410_i4;
  wire signed [`W-1:0] n410_v;
  wire signed [`W-1:0] n590_i0;
  wire signed [`W-1:0] n590_i1;
  wire signed [`W-1:0] n590_v;
  wire signed [`W-1:0] n1085_i0;
  wire signed [`W-1:0] n1085_i1;
  wire signed [`W-1:0] n1085_i2;
  wire signed [`W-1:0] n1085_v;
  wire signed [`W-1:0] _C67_i0;
  wire signed [`W-1:0] _C67_i1;
  wire signed [`W-1:0] _C67_i2;
  wire signed [`W-1:0] _C67_i3;
  wire signed [`W-1:0] _C67_v;
  wire signed [`W-1:0] n1083_i0;
  wire signed [`W-1:0] n1083_i1;
  wire signed [`W-1:0] n1083_i2;
  wire signed [`W-1:0] n1083_i3;
  wire signed [`W-1:0] n1083_i4;
  wire signed [`W-1:0] n1083_v;
  wire signed [`W-1:0] op_T0_jmp_i0;
  wire signed [`W-1:0] op_T0_jmp_i1;
  wire signed [`W-1:0] op_T0_jmp_i2;
  wire signed [`W-1:0] op_T0_jmp_v;
  wire signed [`W-1:0] alub0_i0;
  wire signed [`W-1:0] alub0_i1;
  wire signed [`W-1:0] alub0_i2;
  wire signed [`W-1:0] alub0_i3;
  wire signed [`W-1:0] alub0_i4;
  wire signed [`W-1:0] alub0_v;
  wire signed [`W-1:0] n976_i0;
  wire signed [`W-1:0] n976_i1;
  wire signed [`W-1:0] n976_i2;
  wire signed [`W-1:0] n976_i3;
  wire signed [`W-1:0] n976_i4;
  wire signed [`W-1:0] n976_v;
  wire signed [`W-1:0] n975_i0;
  wire signed [`W-1:0] n975_i1;
  wire signed [`W-1:0] n975_i2;
  wire signed [`W-1:0] n975_v;
  wire signed [`W-1:0] pipeUNK02_i0;
  wire signed [`W-1:0] pipeUNK02_i1;
  wire signed [`W-1:0] pipeUNK02_v;
  wire signed [`W-1:0] n973_i0;
  wire signed [`W-1:0] n973_i1;
  wire signed [`W-1:0] n973_i2;
  wire signed [`W-1:0] n973_v;
  wire signed [`W-1:0] t2_i0;
  wire signed [`W-1:0] t2_i1;
  wire signed [`W-1:0] t2_i2;
  wire signed [`W-1:0] t2_i3;
  wire signed [`W-1:0] t2_i4;
  wire signed [`W-1:0] t2_i5;
  wire signed [`W-1:0] t2_i6;
  wire signed [`W-1:0] t2_i7;
  wire signed [`W-1:0] t2_i8;
  wire signed [`W-1:0] t2_i9;
  wire signed [`W-1:0] t2_i10;
  wire signed [`W-1:0] t2_i11;
  wire signed [`W-1:0] t2_i12;
  wire signed [`W-1:0] t2_i13;
  wire signed [`W-1:0] t2_i14;
  wire signed [`W-1:0] t2_i15;
  wire signed [`W-1:0] t2_i16;
  wire signed [`W-1:0] t2_i17;
  wire signed [`W-1:0] t2_i18;
  wire signed [`W-1:0] t2_i19;
  wire signed [`W-1:0] t2_i20;
  wire signed [`W-1:0] t2_i21;
  wire signed [`W-1:0] t2_v;
  wire signed [`W-1:0] pipeUNK23_i0;
  wire signed [`W-1:0] pipeUNK23_i1;
  wire signed [`W-1:0] pipeUNK23_v;
  wire signed [`W-1:0] n979_i0;
  wire signed [`W-1:0] n979_i1;
  wire signed [`W-1:0] n979_i2;
  wire signed [`W-1:0] n979_v;
  wire signed [`W-1:0] a2_i0;
  wire signed [`W-1:0] a2_i1;
  wire signed [`W-1:0] a2_i2;
  wire signed [`W-1:0] a2_v;
  wire signed [`W-1:0] n182_i0;
  wire signed [`W-1:0] n182_i1;
  wire signed [`W-1:0] n182_i2;
  wire signed [`W-1:0] n182_i3;
  wire signed [`W-1:0] n182_i4;
  wire signed [`W-1:0] n182_v;
  wire signed [`W-1:0] s1_i0;
  wire signed [`W-1:0] s1_i1;
  wire signed [`W-1:0] s1_i2;
  wire signed [`W-1:0] s1_v;
  wire signed [`W-1:0] n180_i0;
  wire signed [`W-1:0] n180_i1;
  wire signed [`W-1:0] n180_i2;
  wire signed [`W-1:0] n180_v;
  wire signed [`W-1:0] nots7_i0;
  wire signed [`W-1:0] nots7_i1;
  wire signed [`W-1:0] nots7_v;
  wire signed [`W-1:0] notRnWprepad_i0;
  wire signed [`W-1:0] notRnWprepad_i1;
  wire signed [`W-1:0] notRnWprepad_i2;
  wire signed [`W-1:0] notRnWprepad_i3;
  wire signed [`W-1:0] notRnWprepad_i4;
  wire signed [`W-1:0] notRnWprepad_v;
  wire signed [`W-1:0] n184_i0;
  wire signed [`W-1:0] n184_i1;
  wire signed [`W-1:0] n184_i2;
  wire signed [`W-1:0] n184_v;
  wire signed [`W-1:0] n188_i0;
  wire signed [`W-1:0] n188_i1;
  wire signed [`W-1:0] n188_i2;
  wire signed [`W-1:0] n188_i3;
  wire signed [`W-1:0] n188_v;
  wire signed [`W-1:0] n1464_i0;
  wire signed [`W-1:0] n1464_i1;
  wire signed [`W-1:0] n1464_i2;
  wire signed [`W-1:0] n1464_v;
  wire signed [`W-1:0] n869_i0;
  wire signed [`W-1:0] n869_i1;
  wire signed [`W-1:0] n869_i2;
  wire signed [`W-1:0] n869_i3;
  wire signed [`W-1:0] n869_v;
  wire signed [`W-1:0] pclp3_i0;
  wire signed [`W-1:0] pclp3_i1;
  wire signed [`W-1:0] pclp3_v;
  wire signed [`W-1:0] n861_i0;
  wire signed [`W-1:0] n861_i1;
  wire signed [`W-1:0] n861_i2;
  wire signed [`W-1:0] n861_v;
  wire signed [`W-1:0] __AxB3__C23_i0;
  wire signed [`W-1:0] __AxB3__C23_i1;
  wire signed [`W-1:0] __AxB3__C23_i2;
  wire signed [`W-1:0] __AxB3__C23_v;
  wire signed [`W-1:0] dpc43_DL_DB_i0;
  wire signed [`W-1:0] dpc43_DL_DB_i1;
  wire signed [`W-1:0] dpc43_DL_DB_i2;
  wire signed [`W-1:0] dpc43_DL_DB_i3;
  wire signed [`W-1:0] dpc43_DL_DB_i4;
  wire signed [`W-1:0] dpc43_DL_DB_i5;
  wire signed [`W-1:0] dpc43_DL_DB_i6;
  wire signed [`W-1:0] dpc43_DL_DB_i7;
  wire signed [`W-1:0] dpc43_DL_DB_i8;
  wire signed [`W-1:0] dpc43_DL_DB_i9;
  wire signed [`W-1:0] dpc43_DL_DB_v;
  wire signed [`W-1:0] n862_i0;
  wire signed [`W-1:0] n862_i1;
  wire signed [`W-1:0] n862_i2;
  wire signed [`W-1:0] n862_i3;
  wire signed [`W-1:0] n862_i4;
  wire signed [`W-1:0] n862_i5;
  wire signed [`W-1:0] n862_i6;
  wire signed [`W-1:0] n862_i7;
  wire signed [`W-1:0] n862_i8;
  wire signed [`W-1:0] n862_i9;
  wire signed [`W-1:0] n862_v;
  wire signed [`W-1:0] n865_i0;
  wire signed [`W-1:0] n865_i1;
  wire signed [`W-1:0] n865_v;
  wire signed [`W-1:0] n867_i0;
  wire signed [`W-1:0] n867_i1;
  wire signed [`W-1:0] n867_i2;
  wire signed [`W-1:0] n867_v;
  wire signed [`W-1:0] n866_i0;
  wire signed [`W-1:0] n866_v;
  wire signed [`W-1:0] n883_i0;
  wire signed [`W-1:0] n883_i1;
  wire signed [`W-1:0] n883_i2;
  wire signed [`W-1:0] n883_v;
  wire signed [`W-1:0] n882_i0;
  wire signed [`W-1:0] n882_i1;
  wire signed [`W-1:0] n882_i2;
  wire signed [`W-1:0] n882_v;
  wire signed [`W-1:0] n880_i0;
  wire signed [`W-1:0] n880_i1;
  wire signed [`W-1:0] n880_i2;
  wire signed [`W-1:0] n880_v;
  wire signed [`W-1:0] ab6_i0;
  wire signed [`W-1:0] ab6_i1;
  wire signed [`W-1:0] ab6_i2;
  wire signed [`W-1:0] ab6_v;
  wire signed [`W-1:0] n885_i0;
  wire signed [`W-1:0] n885_i1;
  wire signed [`W-1:0] n885_i2;
  wire signed [`W-1:0] n885_v;
  wire signed [`W-1:0] n884_i0;
  wire signed [`W-1:0] n884_i1;
  wire signed [`W-1:0] n884_i2;
  wire signed [`W-1:0] n884_v;
  wire signed [`W-1:0] n889_i0;
  wire signed [`W-1:0] n889_i1;
  wire signed [`W-1:0] n889_i2;
  wire signed [`W-1:0] n889_v;
  wire signed [`W-1:0] n888_i0;
  wire signed [`W-1:0] n888_i1;
  wire signed [`W-1:0] n888_i2;
  wire signed [`W-1:0] n888_v;
  wire signed [`W-1:0] abh5_i0;
  wire signed [`W-1:0] abh5_i1;
  wire signed [`W-1:0] abh5_i2;
  wire signed [`W-1:0] abh5_i3;
  wire signed [`W-1:0] abh5_i4;
  wire signed [`W-1:0] abh5_v;
  wire signed [`W-1:0] n774_i0;
  wire signed [`W-1:0] n774_i1;
  wire signed [`W-1:0] n774_i2;
  wire signed [`W-1:0] n774_v;
  wire signed [`W-1:0] x7_i0;
  wire signed [`W-1:0] x7_i1;
  wire signed [`W-1:0] x7_i2;
  wire signed [`W-1:0] x7_v;
  wire signed [`W-1:0] op_T5_jsr_i0;
  wire signed [`W-1:0] op_T5_jsr_i1;
  wire signed [`W-1:0] op_T5_jsr_i2;
  wire signed [`W-1:0] op_T5_jsr_v;
  wire signed [`W-1:0] n771_i0;
  wire signed [`W-1:0] n771_i1;
  wire signed [`W-1:0] n771_i2;
  wire signed [`W-1:0] n771_i3;
  wire signed [`W-1:0] n771_i4;
  wire signed [`W-1:0] n771_v;
  wire signed [`W-1:0] n770_i0;
  wire signed [`W-1:0] n770_i1;
  wire signed [`W-1:0] n770_i2;
  wire signed [`W-1:0] n770_i3;
  wire signed [`W-1:0] n770_v;
  wire signed [`W-1:0] n773_i0;
  wire signed [`W-1:0] n773_i1;
  wire signed [`W-1:0] n773_i2;
  wire signed [`W-1:0] n773_v;
  wire signed [`W-1:0] n772_i0;
  wire signed [`W-1:0] n772_i1;
  wire signed [`W-1:0] n772_i2;
  wire signed [`W-1:0] n772_i3;
  wire signed [`W-1:0] n772_v;
  wire signed [`W-1:0] n779_i0;
  wire signed [`W-1:0] n779_i1;
  wire signed [`W-1:0] n779_i2;
  wire signed [`W-1:0] n779_i3;
  wire signed [`W-1:0] n779_v;
  wire signed [`W-1:0] ONEBYTE_i0;
  wire signed [`W-1:0] ONEBYTE_i1;
  wire signed [`W-1:0] ONEBYTE_i2;
  wire signed [`W-1:0] ONEBYTE_v;
  wire signed [`W-1:0] n419_i0;
  wire signed [`W-1:0] n419_i1;
  wire signed [`W-1:0] n419_i2;
  wire signed [`W-1:0] n419_v;
  wire signed [`W-1:0] Pout6_i0;
  wire signed [`W-1:0] Pout6_i1;
  wire signed [`W-1:0] Pout6_i2;
  wire signed [`W-1:0] Pout6_v;
  wire signed [`W-1:0] op_T0_dex_i0;
  wire signed [`W-1:0] op_T0_dex_i1;
  wire signed [`W-1:0] op_T0_dex_i2;
  wire signed [`W-1:0] op_T0_dex_v;
  wire signed [`W-1:0] n75_i0;
  wire signed [`W-1:0] n75_i1;
  wire signed [`W-1:0] n75_i2;
  wire signed [`W-1:0] n75_v;
  wire signed [`W-1:0] pipeUNK27_i0;
  wire signed [`W-1:0] pipeUNK27_i1;
  wire signed [`W-1:0] pipeUNK27_v;
  wire signed [`W-1:0] n72_i0;
  wire signed [`W-1:0] n72_i1;
  wire signed [`W-1:0] n72_i2;
  wire signed [`W-1:0] n72_i3;
  wire signed [`W-1:0] n72_i4;
  wire signed [`W-1:0] n72_v;
  wire signed [`W-1:0] n71_i0;
  wire signed [`W-1:0] n71_i1;
  wire signed [`W-1:0] n71_i2;
  wire signed [`W-1:0] n71_v;
  wire signed [`W-1:0] n70_i0;
  wire signed [`W-1:0] n70_i1;
  wire signed [`W-1:0] n70_i2;
  wire signed [`W-1:0] n70_v;
  wire signed [`W-1:0] n79_i0;
  wire signed [`W-1:0] n79_i1;
  wire signed [`W-1:0] n79_i2;
  wire signed [`W-1:0] n79_v;
  wire signed [`W-1:0] C34_i0;
  wire signed [`W-1:0] C34_i1;
  wire signed [`W-1:0] C34_i2;
  wire signed [`W-1:0] C34_i3;
  wire signed [`W-1:0] C34_i4;
  wire signed [`W-1:0] C34_i5;
  wire signed [`W-1:0] C34_v;
  wire signed [`W-1:0] n1043_i0;
  wire signed [`W-1:0] n1043_i1;
  wire signed [`W-1:0] n1043_i2;
  wire signed [`W-1:0] n1043_v;
  wire signed [`W-1:0] H1x1_i0;
  wire signed [`W-1:0] H1x1_i1;
  wire signed [`W-1:0] H1x1_i2;
  wire signed [`W-1:0] H1x1_i3;
  wire signed [`W-1:0] H1x1_i4;
  wire signed [`W-1:0] H1x1_i5;
  wire signed [`W-1:0] H1x1_i6;
  wire signed [`W-1:0] H1x1_i7;
  wire signed [`W-1:0] H1x1_i8;
  wire signed [`W-1:0] H1x1_v;
  wire signed [`W-1:0] n1041_i0;
  wire signed [`W-1:0] n1041_i1;
  wire signed [`W-1:0] n1041_i2;
  wire signed [`W-1:0] n1041_v;
  wire signed [`W-1:0] n1047_i0;
  wire signed [`W-1:0] n1047_i1;
  wire signed [`W-1:0] n1047_i2;
  wire signed [`W-1:0] n1047_v;
  wire signed [`W-1:0] n1046_i0;
  wire signed [`W-1:0] n1046_i1;
  wire signed [`W-1:0] n1046_i2;
  wire signed [`W-1:0] n1046_v;
  wire signed [`W-1:0] n1045_i0;
  wire signed [`W-1:0] n1045_i1;
  wire signed [`W-1:0] n1045_i2;
  wire signed [`W-1:0] n1045_i3;
  wire signed [`W-1:0] n1045_i4;
  wire signed [`W-1:0] n1045_v;
  wire signed [`W-1:0] n1044_i0;
  wire signed [`W-1:0] n1044_i1;
  wire signed [`W-1:0] n1044_i2;
  wire signed [`W-1:0] n1044_v;
  wire signed [`W-1:0] n1049_i0;
  wire signed [`W-1:0] n1049_i1;
  wire signed [`W-1:0] n1049_v;
  wire signed [`W-1:0] _op_branch_done_i0;
  wire signed [`W-1:0] _op_branch_done_i1;
  wire signed [`W-1:0] _op_branch_done_i2;
  wire signed [`W-1:0] _op_branch_done_v;
  wire signed [`W-1:0] alua3_i0;
  wire signed [`W-1:0] alua3_i1;
  wire signed [`W-1:0] alua3_i2;
  wire signed [`W-1:0] alua3_i3;
  wire signed [`W-1:0] alua3_v;
  wire signed [`W-1:0] n1683_i0;
  wire signed [`W-1:0] n1683_i1;
  wire signed [`W-1:0] n1683_v;
  wire signed [`W-1:0] n1682_i0;
  wire signed [`W-1:0] n1682_i1;
  wire signed [`W-1:0] n1682_i2;
  wire signed [`W-1:0] n1682_v;
  wire signed [`W-1:0] n1684_i0;
  wire signed [`W-1:0] n1684_i1;
  wire signed [`W-1:0] n1684_i2;
  wire signed [`W-1:0] n1684_v;
  wire signed [`W-1:0] n1687_i0;
  wire signed [`W-1:0] n1687_i1;
  wire signed [`W-1:0] n1687_i2;
  wire signed [`W-1:0] n1687_v;
  wire signed [`W-1:0] op_EORS_i0;
  wire signed [`W-1:0] op_EORS_i1;
  wire signed [`W-1:0] op_EORS_i2;
  wire signed [`W-1:0] op_EORS_i3;
  wire signed [`W-1:0] op_EORS_v;
  wire signed [`W-1:0] n1688_i0;
  wire signed [`W-1:0] n1688_i1;
  wire signed [`W-1:0] n1688_i2;
  wire signed [`W-1:0] n1688_v;
  wire signed [`W-1:0] n1269_i0;
  wire signed [`W-1:0] n1269_i1;
  wire signed [`W-1:0] n1269_i2;
  wire signed [`W-1:0] n1269_v;
  wire signed [`W-1:0] _DBZ_i0;
  wire signed [`W-1:0] _DBZ_i1;
  wire signed [`W-1:0] _DBZ_i2;
  wire signed [`W-1:0] _DBZ_v;
  wire signed [`W-1:0] n669_i0;
  wire signed [`W-1:0] n669_i1;
  wire signed [`W-1:0] n669_i2;
  wire signed [`W-1:0] n669_v;
  wire signed [`W-1:0] _ABH4_i0;
  wire signed [`W-1:0] _ABH4_i1;
  wire signed [`W-1:0] _ABH4_i2;
  wire signed [`W-1:0] _ABH4_v;
  wire signed [`W-1:0] pd5_clearIR_i0;
  wire signed [`W-1:0] pd5_clearIR_i1;
  wire signed [`W-1:0] pd5_clearIR_i2;
  wire signed [`W-1:0] pd5_clearIR_v;
  wire signed [`W-1:0] n1262_i0;
  wire signed [`W-1:0] n1262_i1;
  wire signed [`W-1:0] n1262_i2;
  wire signed [`W-1:0] n1262_i3;
  wire signed [`W-1:0] n1262_v;
  wire signed [`W-1:0] op_T0_ldy_mem_i0;
  wire signed [`W-1:0] op_T0_ldy_mem_i1;
  wire signed [`W-1:0] op_T0_ldy_mem_i2;
  wire signed [`W-1:0] op_T0_ldy_mem_v;
  wire signed [`W-1:0] n664_i0;
  wire signed [`W-1:0] n664_i1;
  wire signed [`W-1:0] n664_i2;
  wire signed [`W-1:0] n664_v;
  wire signed [`W-1:0] n1267_i0;
  wire signed [`W-1:0] n1267_i1;
  wire signed [`W-1:0] n1267_i2;
  wire signed [`W-1:0] n1267_v;
  wire signed [`W-1:0] notdor5_i0;
  wire signed [`W-1:0] notdor5_i1;
  wire signed [`W-1:0] notdor5_v;
  wire signed [`W-1:0] op_T3_branch_i0;
  wire signed [`W-1:0] op_T3_branch_i1;
  wire signed [`W-1:0] op_T3_branch_i2;
  wire signed [`W-1:0] op_T3_branch_i3;
  wire signed [`W-1:0] op_T3_branch_v;
  wire signed [`W-1:0] clk2out_i0;
  wire signed [`W-1:0] clk2out_i1;
  wire signed [`W-1:0] clk2out_i2;
  wire signed [`W-1:0] clk2out_v;
  wire signed [`W-1:0] n1469_i0;
  wire signed [`W-1:0] n1469_i1;
  wire signed [`W-1:0] n1469_i2;
  wire signed [`W-1:0] n1469_v;
  wire signed [`W-1:0] dpc5_SADL_i0;
  wire signed [`W-1:0] dpc5_SADL_i1;
  wire signed [`W-1:0] dpc5_SADL_i2;
  wire signed [`W-1:0] dpc5_SADL_i3;
  wire signed [`W-1:0] dpc5_SADL_i4;
  wire signed [`W-1:0] dpc5_SADL_i5;
  wire signed [`W-1:0] dpc5_SADL_i6;
  wire signed [`W-1:0] dpc5_SADL_i7;
  wire signed [`W-1:0] dpc5_SADL_i8;
  wire signed [`W-1:0] dpc5_SADL_i9;
  wire signed [`W-1:0] dpc5_SADL_v;
  wire signed [`W-1:0] VEC0_i0;
  wire signed [`W-1:0] VEC0_i1;
  wire signed [`W-1:0] VEC0_i2;
  wire signed [`W-1:0] VEC0_i3;
  wire signed [`W-1:0] VEC0_i4;
  wire signed [`W-1:0] VEC0_v;
  wire signed [`W-1:0] n1018_i0;
  wire signed [`W-1:0] n1018_i1;
  wire signed [`W-1:0] n1018_i2;
  wire signed [`W-1:0] n1018_v;
  wire signed [`W-1:0] n1467_i0;
  wire signed [`W-1:0] n1467_i1;
  wire signed [`W-1:0] n1467_i2;
  wire signed [`W-1:0] n1467_v;
  wire signed [`W-1:0] op_rol_ror_i0;
  wire signed [`W-1:0] op_rol_ror_i1;
  wire signed [`W-1:0] op_rol_ror_i2;
  wire signed [`W-1:0] op_rol_ror_v;
  wire signed [`W-1:0] pd6_clearIR_i0;
  wire signed [`W-1:0] pd6_clearIR_i1;
  wire signed [`W-1:0] pd6_clearIR_i2;
  wire signed [`W-1:0] pd6_clearIR_v;
  wire signed [`W-1:0] n1463_i0;
  wire signed [`W-1:0] n1463_i1;
  wire signed [`W-1:0] n1463_i2;
  wire signed [`W-1:0] n1463_i3;
  wire signed [`W-1:0] n1463_v;
  wire signed [`W-1:0] PD_xxxx10x0_i0;
  wire signed [`W-1:0] PD_xxxx10x0_i1;
  wire signed [`W-1:0] PD_xxxx10x0_i2;
  wire signed [`W-1:0] PD_xxxx10x0_i3;
  wire signed [`W-1:0] PD_xxxx10x0_v;
  wire signed [`W-1:0] n1316_i0;
  wire signed [`W-1:0] n1316_i1;
  wire signed [`W-1:0] n1316_i2;
  wire signed [`W-1:0] n1316_i3;
  wire signed [`W-1:0] n1316_i4;
  wire signed [`W-1:0] n1316_v;
  wire signed [`W-1:0] n1315_i0;
  wire signed [`W-1:0] n1315_i1;
  wire signed [`W-1:0] n1315_i2;
  wire signed [`W-1:0] n1315_i3;
  wire signed [`W-1:0] n1315_v;
  wire signed [`W-1:0] C67_i0;
  wire signed [`W-1:0] C67_i1;
  wire signed [`W-1:0] C67_i2;
  wire signed [`W-1:0] C67_i3;
  wire signed [`W-1:0] C67_i4;
  wire signed [`W-1:0] C67_i5;
  wire signed [`W-1:0] C67_v;
  wire signed [`W-1:0] A_B3_i0;
  wire signed [`W-1:0] A_B3_i1;
  wire signed [`W-1:0] A_B3_i2;
  wire signed [`W-1:0] A_B3_v;
  wire signed [`W-1:0] n1312_i0;
  wire signed [`W-1:0] n1312_i1;
  wire signed [`W-1:0] n1312_i2;
  wire signed [`W-1:0] n1312_v;
  wire signed [`W-1:0] op_T4_rti_i0;
  wire signed [`W-1:0] op_T4_rti_i1;
  wire signed [`W-1:0] op_T4_rti_i2;
  wire signed [`W-1:0] op_T4_rti_v;
  wire signed [`W-1:0] n1319_i0;
  wire signed [`W-1:0] n1319_i1;
  wire signed [`W-1:0] n1319_i2;
  wire signed [`W-1:0] n1319_v;
  wire signed [`W-1:0] n1318_i0;
  wire signed [`W-1:0] n1318_i1;
  wire signed [`W-1:0] n1318_i2;
  wire signed [`W-1:0] n1318_i3;
  wire signed [`W-1:0] n1318_i4;
  wire signed [`W-1:0] n1318_i5;
  wire signed [`W-1:0] n1318_v;
  wire signed [`W-1:0] xx_op_T5_jsr_i0;
  wire signed [`W-1:0] xx_op_T5_jsr_i1;
  wire signed [`W-1:0] xx_op_T5_jsr_i2;
  wire signed [`W-1:0] xx_op_T5_jsr_v;
  wire signed [`W-1:0] idl3_i0;
  wire signed [`W-1:0] idl3_i1;
  wire signed [`W-1:0] idl3_i2;
  wire signed [`W-1:0] idl3_v;
  wire signed [`W-1:0] notidl7_i0;
  wire signed [`W-1:0] notidl7_i1;
  wire signed [`W-1:0] notidl7_v;
  wire signed [`W-1:0] n319_i0;
  wire signed [`W-1:0] n319_i1;
  wire signed [`W-1:0] n319_i2;
  wire signed [`W-1:0] n319_v;
  wire signed [`W-1:0] n318_i0;
  wire signed [`W-1:0] n318_i1;
  wire signed [`W-1:0] n318_i2;
  wire signed [`W-1:0] n318_i3;
  wire signed [`W-1:0] n318_i4;
  wire signed [`W-1:0] n318_v;
  wire signed [`W-1:0] n312_i0;
  wire signed [`W-1:0] n312_i1;
  wire signed [`W-1:0] n312_i2;
  wire signed [`W-1:0] n312_i3;
  wire signed [`W-1:0] n312_v;
  wire signed [`W-1:0] n311_i0;
  wire signed [`W-1:0] n311_i1;
  wire signed [`W-1:0] n311_i2;
  wire signed [`W-1:0] n311_i3;
  wire signed [`W-1:0] n311_v;
  wire signed [`W-1:0] n310_i0;
  wire signed [`W-1:0] n310_i1;
  wire signed [`W-1:0] n310_i2;
  wire signed [`W-1:0] n310_v;
  wire signed [`W-1:0] n317_i0;
  wire signed [`W-1:0] n317_i1;
  wire signed [`W-1:0] n317_i2;
  wire signed [`W-1:0] n317_v;
  wire signed [`W-1:0] adh3_i0;
  wire signed [`W-1:0] adh3_i1;
  wire signed [`W-1:0] adh3_i2;
  wire signed [`W-1:0] adh3_i3;
  wire signed [`W-1:0] adh3_i4;
  wire signed [`W-1:0] adh3_i5;
  wire signed [`W-1:0] adh3_i6;
  wire signed [`W-1:0] adh3_v;
  wire signed [`W-1:0] alu5_i0;
  wire signed [`W-1:0] alu5_i1;
  wire signed [`W-1:0] alu5_i2;
  wire signed [`W-1:0] alu5_i3;
  wire signed [`W-1:0] alu5_i4;
  wire signed [`W-1:0] alu5_v;
  wire signed [`W-1:0] n1335_i0;
  wire signed [`W-1:0] n1335_i1;
  wire signed [`W-1:0] n1335_i2;
  wire signed [`W-1:0] n1335_v;
  wire signed [`W-1:0] dpc35_PCHC_i0;
  wire signed [`W-1:0] dpc35_PCHC_i1;
  wire signed [`W-1:0] dpc35_PCHC_i2;
  wire signed [`W-1:0] dpc35_PCHC_i3;
  wire signed [`W-1:0] dpc35_PCHC_v;
  wire signed [`W-1:0] n441_i0;
  wire signed [`W-1:0] n441_i1;
  wire signed [`W-1:0] n441_i2;
  wire signed [`W-1:0] n441_v;
  wire signed [`W-1:0] n440_i0;
  wire signed [`W-1:0] n440_i1;
  wire signed [`W-1:0] n440_i2;
  wire signed [`W-1:0] n440_i3;
  wire signed [`W-1:0] n440_i4;
  wire signed [`W-1:0] n440_i5;
  wire signed [`W-1:0] n440_i6;
  wire signed [`W-1:0] n440_i7;
  wire signed [`W-1:0] n440_i8;
  wire signed [`W-1:0] n440_i9;
  wire signed [`W-1:0] n440_i10;
  wire signed [`W-1:0] n440_v;
  wire signed [`W-1:0] dpc26_ACDB_i0;
  wire signed [`W-1:0] dpc26_ACDB_i1;
  wire signed [`W-1:0] dpc26_ACDB_i2;
  wire signed [`W-1:0] dpc26_ACDB_i3;
  wire signed [`W-1:0] dpc26_ACDB_i4;
  wire signed [`W-1:0] dpc26_ACDB_i5;
  wire signed [`W-1:0] dpc26_ACDB_i6;
  wire signed [`W-1:0] dpc26_ACDB_i7;
  wire signed [`W-1:0] dpc26_ACDB_i8;
  wire signed [`W-1:0] dpc26_ACDB_i9;
  wire signed [`W-1:0] dpc26_ACDB_v;
  wire signed [`W-1:0] n1333_i0;
  wire signed [`W-1:0] n1333_i1;
  wire signed [`W-1:0] n1333_v;
  wire signed [`W-1:0] dor3_i0;
  wire signed [`W-1:0] dor3_i1;
  wire signed [`W-1:0] dor3_i2;
  wire signed [`W-1:0] dor3_i3;
  wire signed [`W-1:0] dor3_i4;
  wire signed [`W-1:0] dor3_v;
  wire signed [`W-1:0] n632_i0;
  wire signed [`W-1:0] n632_i1;
  wire signed [`W-1:0] n632_i2;
  wire signed [`W-1:0] n632_v;
  wire signed [`W-1:0] n1521_i0;
  wire signed [`W-1:0] n1521_i1;
  wire signed [`W-1:0] n1521_i2;
  wire signed [`W-1:0] n1521_v;
  wire signed [`W-1:0] n633_i0;
  wire signed [`W-1:0] n633_v;
  wire signed [`W-1:0] n964_i0;
  wire signed [`W-1:0] n964_i1;
  wire signed [`W-1:0] n964_i2;
  wire signed [`W-1:0] n964_i3;
  wire signed [`W-1:0] n964_v;
  wire signed [`W-1:0] __AxBxC_1_i0;
  wire signed [`W-1:0] __AxBxC_1_i1;
  wire signed [`W-1:0] __AxBxC_1_i2;
  wire signed [`W-1:0] __AxBxC_1_v;
  wire signed [`W-1:0] n966_i0;
  wire signed [`W-1:0] n966_i1;
  wire signed [`W-1:0] n966_i2;
  wire signed [`W-1:0] n966_i3;
  wire signed [`W-1:0] n966_v;
  wire signed [`W-1:0] nnT2BR_i0;
  wire signed [`W-1:0] nnT2BR_i1;
  wire signed [`W-1:0] nnT2BR_i2;
  wire signed [`W-1:0] nnT2BR_i3;
  wire signed [`W-1:0] nnT2BR_i4;
  wire signed [`W-1:0] nnT2BR_i5;
  wire signed [`W-1:0] nnT2BR_i6;
  wire signed [`W-1:0] nnT2BR_i7;
  wire signed [`W-1:0] nnT2BR_i8;
  wire signed [`W-1:0] nnT2BR_i9;
  wire signed [`W-1:0] nnT2BR_i10;
  wire signed [`W-1:0] nnT2BR_v;
  wire signed [`W-1:0] pipeUNK32_i0;
  wire signed [`W-1:0] pipeUNK32_i1;
  wire signed [`W-1:0] pipeUNK32_v;
  wire signed [`W-1:0] n961_i0;
  wire signed [`W-1:0] n961_i1;
  wire signed [`W-1:0] n961_i2;
  wire signed [`W-1:0] n961_v;
  wire signed [`W-1:0] n962_i0;
  wire signed [`W-1:0] n962_i1;
  wire signed [`W-1:0] n962_i2;
  wire signed [`W-1:0] n962_v;
  wire signed [`W-1:0] n963_i0;
  wire signed [`W-1:0] n963_i1;
  wire signed [`W-1:0] n963_i2;
  wire signed [`W-1:0] n963_v;
  wire signed [`W-1:0] n968_i0;
  wire signed [`W-1:0] n968_i1;
  wire signed [`W-1:0] n968_v;
  wire signed [`W-1:0] n969_i0;
  wire signed [`W-1:0] n969_i1;
  wire signed [`W-1:0] n969_i2;
  wire signed [`W-1:0] n969_v;
  wire signed [`W-1:0] n400_i0;
  wire signed [`W-1:0] n400_i1;
  wire signed [`W-1:0] n400_i2;
  wire signed [`W-1:0] n400_i3;
  wire signed [`W-1:0] n400_v;
  wire signed [`W-1:0] AxB7_i0;
  wire signed [`W-1:0] AxB7_i1;
  wire signed [`W-1:0] AxB7_i2;
  wire signed [`W-1:0] AxB7_i3;
  wire signed [`W-1:0] AxB7_i4;
  wire signed [`W-1:0] AxB7_i5;
  wire signed [`W-1:0] AxB7_v;
  wire signed [`W-1:0] n878_i0;
  wire signed [`W-1:0] n878_i1;
  wire signed [`W-1:0] n878_v;
  wire signed [`W-1:0] n1240_i0;
  wire signed [`W-1:0] n1240_i1;
  wire signed [`W-1:0] n1240_i2;
  wire signed [`W-1:0] n1240_v;
  wire signed [`W-1:0] n876_i0;
  wire signed [`W-1:0] n876_i1;
  wire signed [`W-1:0] n876_i2;
  wire signed [`W-1:0] n876_v;
  wire signed [`W-1:0] n877_i0;
  wire signed [`W-1:0] n877_i1;
  wire signed [`W-1:0] n877_i2;
  wire signed [`W-1:0] n877_v;
  wire signed [`W-1:0] dpc6_SBS_i0;
  wire signed [`W-1:0] dpc6_SBS_i1;
  wire signed [`W-1:0] dpc6_SBS_i2;
  wire signed [`W-1:0] dpc6_SBS_i3;
  wire signed [`W-1:0] dpc6_SBS_i4;
  wire signed [`W-1:0] dpc6_SBS_i5;
  wire signed [`W-1:0] dpc6_SBS_i6;
  wire signed [`W-1:0] dpc6_SBS_i7;
  wire signed [`W-1:0] dpc6_SBS_i8;
  wire signed [`W-1:0] dpc6_SBS_i9;
  wire signed [`W-1:0] dpc6_SBS_v;
  wire signed [`W-1:0] n875_i0;
  wire signed [`W-1:0] n875_i1;
  wire signed [`W-1:0] n875_i2;
  wire signed [`W-1:0] n875_v;
  wire signed [`W-1:0] alu1_i0;
  wire signed [`W-1:0] alu1_i1;
  wire signed [`W-1:0] alu1_i2;
  wire signed [`W-1:0] alu1_i3;
  wire signed [`W-1:0] alu1_i4;
  wire signed [`W-1:0] alu1_v;
  wire signed [`W-1:0] op_T__ora_and_eor_adc_i0;
  wire signed [`W-1:0] op_T__ora_and_eor_adc_i1;
  wire signed [`W-1:0] op_T__ora_and_eor_adc_i2;
  wire signed [`W-1:0] op_T__ora_and_eor_adc_v;
  wire signed [`W-1:0] idl1_i0;
  wire signed [`W-1:0] idl1_i1;
  wire signed [`W-1:0] idl1_i2;
  wire signed [`W-1:0] idl1_v;
  wire signed [`W-1:0] n871_i0;
  wire signed [`W-1:0] n871_i1;
  wire signed [`W-1:0] n871_i2;
  wire signed [`W-1:0] n871_i3;
  wire signed [`W-1:0] n871_v;
  wire signed [`W-1:0] adl2_i0;
  wire signed [`W-1:0] adl2_i1;
  wire signed [`W-1:0] adl2_i2;
  wire signed [`W-1:0] adl2_i3;
  wire signed [`W-1:0] adl2_i4;
  wire signed [`W-1:0] adl2_i5;
  wire signed [`W-1:0] adl2_i6;
  wire signed [`W-1:0] adl2_i7;
  wire signed [`W-1:0] adl2_i8;
  wire signed [`W-1:0] adl2_v;
  wire signed [`W-1:0] n9_i0;
  wire signed [`W-1:0] n9_v;
  wire signed [`W-1:0] n1533_i0;
  wire signed [`W-1:0] n1533_i1;
  wire signed [`W-1:0] n1533_i2;
  wire signed [`W-1:0] n1533_v;
  wire signed [`W-1:0] n644_i0;
  wire signed [`W-1:0] n644_i1;
  wire signed [`W-1:0] n644_v;
  wire signed [`W-1:0] n890_i0;
  wire signed [`W-1:0] n890_i1;
  wire signed [`W-1:0] n890_i2;
  wire signed [`W-1:0] n890_v;
  wire signed [`W-1:0] idb4_i0;
  wire signed [`W-1:0] idb4_i1;
  wire signed [`W-1:0] idb4_i2;
  wire signed [`W-1:0] idb4_i3;
  wire signed [`W-1:0] idb4_i4;
  wire signed [`W-1:0] idb4_i5;
  wire signed [`W-1:0] idb4_i6;
  wire signed [`W-1:0] idb4_i7;
  wire signed [`W-1:0] idb4_i8;
  wire signed [`W-1:0] idb4_i9;
  wire signed [`W-1:0] idb4_i10;
  wire signed [`W-1:0] idb4_v;
  wire signed [`W-1:0] notalu5_i0;
  wire signed [`W-1:0] notalu5_i1;
  wire signed [`W-1:0] notalu5_v;
  wire signed [`W-1:0] pd3_i0;
  wire signed [`W-1:0] pd3_i1;
  wire signed [`W-1:0] pd3_v;
  wire signed [`W-1:0] n1247_i0;
  wire signed [`W-1:0] n1247_i1;
  wire signed [`W-1:0] n1247_i2;
  wire signed [`W-1:0] n1247_i3;
  wire signed [`W-1:0] n1247_i4;
  wire signed [`W-1:0] n1247_i5;
  wire signed [`W-1:0] n1247_i6;
  wire signed [`W-1:0] n1247_i7;
  wire signed [`W-1:0] n1247_i8;
  wire signed [`W-1:0] n1247_i9;
  wire signed [`W-1:0] n1247_i10;
  wire signed [`W-1:0] n1247_i11;
  wire signed [`W-1:0] n1247_i12;
  wire signed [`W-1:0] n1247_i13;
  wire signed [`W-1:0] n1247_i14;
  wire signed [`W-1:0] n1247_i15;
  wire signed [`W-1:0] n1247_i16;
  wire signed [`W-1:0] n1247_i17;
  wire signed [`W-1:0] n1247_i18;
  wire signed [`W-1:0] n1247_i19;
  wire signed [`W-1:0] n1247_v;
  wire signed [`W-1:0] n896_i0;
  wire signed [`W-1:0] n896_i1;
  wire signed [`W-1:0] n896_i2;
  wire signed [`W-1:0] n896_v;
  wire signed [`W-1:0] n897_i0;
  wire signed [`W-1:0] n897_i1;
  wire signed [`W-1:0] n897_v;
  wire signed [`W-1:0] dpc39_PCLPCL_i0;
  wire signed [`W-1:0] dpc39_PCLPCL_i1;
  wire signed [`W-1:0] dpc39_PCLPCL_i2;
  wire signed [`W-1:0] dpc39_PCLPCL_i3;
  wire signed [`W-1:0] dpc39_PCLPCL_i4;
  wire signed [`W-1:0] dpc39_PCLPCL_i5;
  wire signed [`W-1:0] dpc39_PCLPCL_i6;
  wire signed [`W-1:0] dpc39_PCLPCL_i7;
  wire signed [`W-1:0] dpc39_PCLPCL_i8;
  wire signed [`W-1:0] dpc39_PCLPCL_i9;
  wire signed [`W-1:0] dpc39_PCLPCL_v;
  wire signed [`W-1:0] pipeUNK18_i0;
  wire signed [`W-1:0] pipeUNK18_i1;
  wire signed [`W-1:0] pipeUNK18_v;
  wire signed [`W-1:0] pipeUNK01_i0;
  wire signed [`W-1:0] pipeUNK01_i1;
  wire signed [`W-1:0] pipeUNK01_v;
  wire signed [`W-1:0] n641_i0;
  wire signed [`W-1:0] n641_i1;
  wire signed [`W-1:0] n641_i2;
  wire signed [`W-1:0] n641_i3;
  wire signed [`W-1:0] n641_v;
  wire signed [`W-1:0] _ABH2_i0;
  wire signed [`W-1:0] _ABH2_i1;
  wire signed [`W-1:0] _ABH2_i2;
  wire signed [`W-1:0] _ABH2_v;
  wire signed [`W-1:0] n769_i0;
  wire signed [`W-1:0] n769_i1;
  wire signed [`W-1:0] n769_i2;
  wire signed [`W-1:0] n769_i3;
  wire signed [`W-1:0] n769_v;
  wire signed [`W-1:0] n762_i0;
  wire signed [`W-1:0] n762_i1;
  wire signed [`W-1:0] n762_i2;
  wire signed [`W-1:0] n762_v;
  wire signed [`W-1:0] n763_i0;
  wire signed [`W-1:0] n763_i1;
  wire signed [`W-1:0] n763_i2;
  wire signed [`W-1:0] n763_v;
  wire signed [`W-1:0] n760_i0;
  wire signed [`W-1:0] n760_i1;
  wire signed [`W-1:0] n760_v;
  wire signed [`W-1:0] clock1_i0;
  wire signed [`W-1:0] clock1_i1;
  wire signed [`W-1:0] clock1_i2;
  wire signed [`W-1:0] clock1_i3;
  wire signed [`W-1:0] clock1_i4;
  wire signed [`W-1:0] clock1_i5;
  wire signed [`W-1:0] clock1_i6;
  wire signed [`W-1:0] clock1_i7;
  wire signed [`W-1:0] clock1_i8;
  wire signed [`W-1:0] clock1_i9;
  wire signed [`W-1:0] clock1_i10;
  wire signed [`W-1:0] clock1_i11;
  wire signed [`W-1:0] clock1_i12;
  wire signed [`W-1:0] clock1_i13;
  wire signed [`W-1:0] clock1_i14;
  wire signed [`W-1:0] clock1_i15;
  wire signed [`W-1:0] clock1_i16;
  wire signed [`W-1:0] clock1_i17;
  wire signed [`W-1:0] clock1_i18;
  wire signed [`W-1:0] clock1_i19;
  wire signed [`W-1:0] clock1_i20;
  wire signed [`W-1:0] clock1_i21;
  wire signed [`W-1:0] clock1_i22;
  wire signed [`W-1:0] clock1_i23;
  wire signed [`W-1:0] clock1_i24;
  wire signed [`W-1:0] clock1_i25;
  wire signed [`W-1:0] clock1_i26;
  wire signed [`W-1:0] clock1_i27;
  wire signed [`W-1:0] clock1_i28;
  wire signed [`W-1:0] clock1_i29;
  wire signed [`W-1:0] clock1_i30;
  wire signed [`W-1:0] clock1_i31;
  wire signed [`W-1:0] clock1_i32;
  wire signed [`W-1:0] clock1_i33;
  wire signed [`W-1:0] clock1_i34;
  wire signed [`W-1:0] clock1_i35;
  wire signed [`W-1:0] clock1_i36;
  wire signed [`W-1:0] clock1_i37;
  wire signed [`W-1:0] clock1_i38;
  wire signed [`W-1:0] clock1_i39;
  wire signed [`W-1:0] clock1_i40;
  wire signed [`W-1:0] clock1_v;
  wire signed [`W-1:0] n767_i0;
  wire signed [`W-1:0] n767_i1;
  wire signed [`W-1:0] n767_i2;
  wire signed [`W-1:0] n767_i3;
  wire signed [`W-1:0] n767_v;
  wire signed [`W-1:0] op_jmp_i0;
  wire signed [`W-1:0] op_jmp_i1;
  wire signed [`W-1:0] op_jmp_i2;
  wire signed [`W-1:0] op_jmp_v;
  wire signed [`W-1:0] alu7_i0;
  wire signed [`W-1:0] alu7_i1;
  wire signed [`W-1:0] alu7_i2;
  wire signed [`W-1:0] alu7_i3;
  wire signed [`W-1:0] alu7_v;
  wire signed [`W-1:0] pipeUNK17_i0;
  wire signed [`W-1:0] pipeUNK17_i1;
  wire signed [`W-1:0] pipeUNK17_v;
  wire signed [`W-1:0] pclp2_i0;
  wire signed [`W-1:0] pclp2_i1;
  wire signed [`W-1:0] pclp2_i2;
  wire signed [`W-1:0] pclp2_v;
  wire signed [`W-1:0] n1076_i0;
  wire signed [`W-1:0] n1076_i1;
  wire signed [`W-1:0] n1076_i2;
  wire signed [`W-1:0] n1076_v;
  wire signed [`W-1:0] clearIR_i0;
  wire signed [`W-1:0] clearIR_i1;
  wire signed [`W-1:0] clearIR_i2;
  wire signed [`W-1:0] clearIR_i3;
  wire signed [`W-1:0] clearIR_i4;
  wire signed [`W-1:0] clearIR_i5;
  wire signed [`W-1:0] clearIR_i6;
  wire signed [`W-1:0] clearIR_i7;
  wire signed [`W-1:0] clearIR_i8;
  wire signed [`W-1:0] clearIR_i9;
  wire signed [`W-1:0] clearIR_v;
  wire signed [`W-1:0] op_T0_shift_right_a_i0;
  wire signed [`W-1:0] op_T0_shift_right_a_i1;
  wire signed [`W-1:0] op_T0_shift_right_a_i2;
  wire signed [`W-1:0] op_T0_shift_right_a_v;
  wire signed [`W-1:0] n1075_i0;
  wire signed [`W-1:0] n1075_i1;
  wire signed [`W-1:0] n1075_i2;
  wire signed [`W-1:0] n1075_v;
  wire signed [`W-1:0] n1072_i0;
  wire signed [`W-1:0] n1072_i1;
  wire signed [`W-1:0] n1072_i2;
  wire signed [`W-1:0] n1072_v;
  wire signed [`W-1:0] n1073_i0;
  wire signed [`W-1:0] n1073_i1;
  wire signed [`W-1:0] n1073_i2;
  wire signed [`W-1:0] n1073_v;
  wire signed [`W-1:0] n1070_i0;
  wire signed [`W-1:0] n1070_i1;
  wire signed [`W-1:0] n1070_i2;
  wire signed [`W-1:0] n1070_i3;
  wire signed [`W-1:0] n1070_i4;
  wire signed [`W-1:0] n1070_v;
  wire signed [`W-1:0] n1071_i0;
  wire signed [`W-1:0] n1071_i1;
  wire signed [`W-1:0] n1071_i2;
  wire signed [`W-1:0] n1071_i3;
  wire signed [`W-1:0] n1071_i4;
  wire signed [`W-1:0] n1071_i5;
  wire signed [`W-1:0] n1071_v;
  wire signed [`W-1:0] alub5_i0;
  wire signed [`W-1:0] alub5_i1;
  wire signed [`W-1:0] alub5_i2;
  wire signed [`W-1:0] alub5_i3;
  wire signed [`W-1:0] alub5_i4;
  wire signed [`W-1:0] alub5_v;
  wire signed [`W-1:0] n1679_i0;
  wire signed [`W-1:0] n1679_i1;
  wire signed [`W-1:0] n1679_v;
  wire signed [`W-1:0] n1674_i0;
  wire signed [`W-1:0] n1674_i1;
  wire signed [`W-1:0] n1674_v;
  wire signed [`W-1:0] n1675_i0;
  wire signed [`W-1:0] n1675_i1;
  wire signed [`W-1:0] n1675_i2;
  wire signed [`W-1:0] n1675_v;
  wire signed [`W-1:0] n1676_i0;
  wire signed [`W-1:0] n1676_i1;
  wire signed [`W-1:0] n1676_i2;
  wire signed [`W-1:0] n1676_i3;
  wire signed [`W-1:0] n1676_v;
  wire signed [`W-1:0] n1677_i0;
  wire signed [`W-1:0] n1677_i1;
  wire signed [`W-1:0] n1677_i2;
  wire signed [`W-1:0] n1677_i3;
  wire signed [`W-1:0] n1677_v;
  wire signed [`W-1:0] pch0_i0;
  wire signed [`W-1:0] pch0_i1;
  wire signed [`W-1:0] pch0_i2;
  wire signed [`W-1:0] pch0_v;
  wire signed [`W-1:0] pd2_clearIR_i0;
  wire signed [`W-1:0] pd2_clearIR_i1;
  wire signed [`W-1:0] pd2_clearIR_i2;
  wire signed [`W-1:0] pd2_clearIR_i3;
  wire signed [`W-1:0] pd2_clearIR_i4;
  wire signed [`W-1:0] pd2_clearIR_i5;
  wire signed [`W-1:0] pd2_clearIR_v;
  wire signed [`W-1:0] so_i0;
  wire signed [`W-1:0] so_i1;
  wire signed [`W-1:0] so_i2;
  wire signed [`W-1:0] so_v;
  wire signed [`W-1:0] n1673_i0;
  wire signed [`W-1:0] n1673_i1;
  wire signed [`W-1:0] n1673_v;
  wire signed [`W-1:0] n1094_i0;
  wire signed [`W-1:0] n1094_i1;
  wire signed [`W-1:0] n1094_i2;
  wire signed [`W-1:0] n1094_v;
  wire signed [`W-1:0] n1095_i0;
  wire signed [`W-1:0] n1095_i1;
  wire signed [`W-1:0] n1095_i2;
  wire signed [`W-1:0] n1095_i3;
  wire signed [`W-1:0] n1095_v;
  wire signed [`W-1:0] abl0_i0;
  wire signed [`W-1:0] abl0_i1;
  wire signed [`W-1:0] abl0_i2;
  wire signed [`W-1:0] abl0_i3;
  wire signed [`W-1:0] abl0_i4;
  wire signed [`W-1:0] abl0_v;
  wire signed [`W-1:0] n1097_i0;
  wire signed [`W-1:0] n1097_i1;
  wire signed [`W-1:0] n1097_i2;
  wire signed [`W-1:0] n1097_v;
  wire signed [`W-1:0] n678_i0;
  wire signed [`W-1:0] n678_i1;
  wire signed [`W-1:0] n678_i2;
  wire signed [`W-1:0] n678_i3;
  wire signed [`W-1:0] n678_v;
  wire signed [`W-1:0] n1091_i0;
  wire signed [`W-1:0] n1091_i1;
  wire signed [`W-1:0] n1091_i2;
  wire signed [`W-1:0] n1091_v;
  wire signed [`W-1:0] n642_i0;
  wire signed [`W-1:0] n642_i1;
  wire signed [`W-1:0] n642_i2;
  wire signed [`W-1:0] n642_i3;
  wire signed [`W-1:0] n642_v;
  wire signed [`W-1:0] n674_i0;
  wire signed [`W-1:0] n674_i1;
  wire signed [`W-1:0] n674_i2;
  wire signed [`W-1:0] n674_v;
  wire signed [`W-1:0] n675_i0;
  wire signed [`W-1:0] n675_i1;
  wire signed [`W-1:0] n675_v;
  wire signed [`W-1:0] n676_i0;
  wire signed [`W-1:0] n676_i1;
  wire signed [`W-1:0] n676_i2;
  wire signed [`W-1:0] n676_i3;
  wire signed [`W-1:0] n676_v;
  wire signed [`W-1:0] op_T3_abs_idx_ind_i0;
  wire signed [`W-1:0] op_T3_abs_idx_ind_i1;
  wire signed [`W-1:0] op_T3_abs_idx_ind_i2;
  wire signed [`W-1:0] op_T3_abs_idx_ind_v;
  wire signed [`W-1:0] n670_i0;
  wire signed [`W-1:0] n670_i1;
  wire signed [`W-1:0] n670_i2;
  wire signed [`W-1:0] n670_i3;
  wire signed [`W-1:0] n670_v;
  wire signed [`W-1:0] n671_i0;
  wire signed [`W-1:0] n671_i1;
  wire signed [`W-1:0] n671_v;
  wire signed [`W-1:0] ab14_i0;
  wire signed [`W-1:0] ab14_i1;
  wire signed [`W-1:0] ab14_i2;
  wire signed [`W-1:0] ab14_v;
  wire signed [`W-1:0] n673_i0;
  wire signed [`W-1:0] n673_i1;
  wire signed [`W-1:0] n673_i2;
  wire signed [`W-1:0] n673_v;
  wire signed [`W-1:0] notdor6_i0;
  wire signed [`W-1:0] notdor6_i1;
  wire signed [`W-1:0] notdor6_v;
  wire signed [`W-1:0] op_T0_cld_sed_i0;
  wire signed [`W-1:0] op_T0_cld_sed_i1;
  wire signed [`W-1:0] op_T0_cld_sed_i2;
  wire signed [`W-1:0] op_T0_cld_sed_v;
  wire signed [`W-1:0] pd7_clearIR_i0;
  wire signed [`W-1:0] pd7_clearIR_i1;
  wire signed [`W-1:0] pd7_clearIR_i2;
  wire signed [`W-1:0] pd7_clearIR_i3;
  wire signed [`W-1:0] pd7_clearIR_v;
  wire signed [`W-1:0] n1411_i0;
  wire signed [`W-1:0] n1411_i1;
  wire signed [`W-1:0] n1411_v;
  wire signed [`W-1:0] n1412_i0;
  wire signed [`W-1:0] n1412_i1;
  wire signed [`W-1:0] n1412_i2;
  wire signed [`W-1:0] n1412_v;
  wire signed [`W-1:0] n1413_i0;
  wire signed [`W-1:0] n1413_i1;
  wire signed [`W-1:0] n1413_i2;
  wire signed [`W-1:0] n1413_v;
  wire signed [`W-1:0] alu3_i0;
  wire signed [`W-1:0] alu3_i1;
  wire signed [`W-1:0] alu3_i2;
  wire signed [`W-1:0] alu3_i3;
  wire signed [`W-1:0] alu3_v;
  wire signed [`W-1:0] dor6_i0;
  wire signed [`W-1:0] dor6_i1;
  wire signed [`W-1:0] dor6_i2;
  wire signed [`W-1:0] dor6_i3;
  wire signed [`W-1:0] dor6_i4;
  wire signed [`W-1:0] dor6_v;
  wire signed [`W-1:0] n1416_i0;
  wire signed [`W-1:0] n1416_i1;
  wire signed [`W-1:0] n1416_i2;
  wire signed [`W-1:0] n1416_v;
  wire signed [`W-1:0] n1417_i0;
  wire signed [`W-1:0] n1417_i1;
  wire signed [`W-1:0] n1417_i2;
  wire signed [`W-1:0] n1417_v;
  wire signed [`W-1:0] n1323_i0;
  wire signed [`W-1:0] n1323_i1;
  wire signed [`W-1:0] n1323_i2;
  wire signed [`W-1:0] n1323_v;
  wire signed [`W-1:0] notir7_i0;
  wire signed [`W-1:0] notir7_i1;
  wire signed [`W-1:0] notir7_i2;
  wire signed [`W-1:0] notir7_i3;
  wire signed [`W-1:0] notir7_i4;
  wire signed [`W-1:0] notir7_i5;
  wire signed [`W-1:0] notir7_i6;
  wire signed [`W-1:0] notir7_i7;
  wire signed [`W-1:0] notir7_i8;
  wire signed [`W-1:0] notir7_i9;
  wire signed [`W-1:0] notir7_i10;
  wire signed [`W-1:0] notir7_i11;
  wire signed [`W-1:0] notir7_i12;
  wire signed [`W-1:0] notir7_i13;
  wire signed [`W-1:0] notir7_i14;
  wire signed [`W-1:0] notir7_i15;
  wire signed [`W-1:0] notir7_i16;
  wire signed [`W-1:0] notir7_i17;
  wire signed [`W-1:0] notir7_i18;
  wire signed [`W-1:0] notir7_i19;
  wire signed [`W-1:0] notir7_i20;
  wire signed [`W-1:0] notir7_i21;
  wire signed [`W-1:0] notir7_i22;
  wire signed [`W-1:0] notir7_i23;
  wire signed [`W-1:0] notir7_i24;
  wire signed [`W-1:0] notir7_i25;
  wire signed [`W-1:0] notir7_i26;
  wire signed [`W-1:0] notir7_i27;
  wire signed [`W-1:0] notir7_i28;
  wire signed [`W-1:0] notir7_i29;
  wire signed [`W-1:0] notir7_i30;
  wire signed [`W-1:0] notir7_i31;
  wire signed [`W-1:0] notir7_i32;
  wire signed [`W-1:0] notir7_i33;
  wire signed [`W-1:0] notir7_i34;
  wire signed [`W-1:0] notir7_i35;
  wire signed [`W-1:0] notir7_v;
  wire signed [`W-1:0] s3_i0;
  wire signed [`W-1:0] s3_i1;
  wire signed [`W-1:0] s3_i2;
  wire signed [`W-1:0] s3_v;
  wire signed [`W-1:0] pclp5_i0;
  wire signed [`W-1:0] pclp5_i1;
  wire signed [`W-1:0] pclp5_v;
  wire signed [`W-1:0] _C78_i0;
  wire signed [`W-1:0] _C78_i1;
  wire signed [`W-1:0] _C78_i2;
  wire signed [`W-1:0] _C78_v;
  wire signed [`W-1:0] op_T__shift_a_i0;
  wire signed [`W-1:0] op_T__shift_a_i1;
  wire signed [`W-1:0] op_T__shift_a_i2;
  wire signed [`W-1:0] op_T__shift_a_v;
  wire signed [`W-1:0] n1325_i0;
  wire signed [`W-1:0] n1325_i1;
  wire signed [`W-1:0] n1325_i2;
  wire signed [`W-1:0] n1325_v;
  wire signed [`W-1:0] ir7_i0;
  wire signed [`W-1:0] ir7_i1;
  wire signed [`W-1:0] ir7_i2;
  wire signed [`W-1:0] ir7_i3;
  wire signed [`W-1:0] ir7_i4;
  wire signed [`W-1:0] ir7_i5;
  wire signed [`W-1:0] ir7_i6;
  wire signed [`W-1:0] ir7_i7;
  wire signed [`W-1:0] ir7_i8;
  wire signed [`W-1:0] ir7_i9;
  wire signed [`W-1:0] ir7_i10;
  wire signed [`W-1:0] ir7_i11;
  wire signed [`W-1:0] ir7_i12;
  wire signed [`W-1:0] ir7_i13;
  wire signed [`W-1:0] ir7_i14;
  wire signed [`W-1:0] ir7_i15;
  wire signed [`W-1:0] ir7_i16;
  wire signed [`W-1:0] ir7_i17;
  wire signed [`W-1:0] ir7_i18;
  wire signed [`W-1:0] ir7_i19;
  wire signed [`W-1:0] ir7_i20;
  wire signed [`W-1:0] ir7_i21;
  wire signed [`W-1:0] ir7_i22;
  wire signed [`W-1:0] ir7_i23;
  wire signed [`W-1:0] ir7_i24;
  wire signed [`W-1:0] ir7_i25;
  wire signed [`W-1:0] ir7_i26;
  wire signed [`W-1:0] ir7_i27;
  wire signed [`W-1:0] ir7_i28;
  wire signed [`W-1:0] ir7_i29;
  wire signed [`W-1:0] ir7_i30;
  wire signed [`W-1:0] ir7_i31;
  wire signed [`W-1:0] ir7_i32;
  wire signed [`W-1:0] ir7_i33;
  wire signed [`W-1:0] ir7_i34;
  wire signed [`W-1:0] ir7_i35;
  wire signed [`W-1:0] ir7_i36;
  wire signed [`W-1:0] ir7_i37;
  wire signed [`W-1:0] ir7_i38;
  wire signed [`W-1:0] ir7_i39;
  wire signed [`W-1:0] ir7_i40;
  wire signed [`W-1:0] ir7_i41;
  wire signed [`W-1:0] ir7_i42;
  wire signed [`W-1:0] ir7_i43;
  wire signed [`W-1:0] ir7_i44;
  wire signed [`W-1:0] ir7_i45;
  wire signed [`W-1:0] ir7_i46;
  wire signed [`W-1:0] ir7_i47;
  wire signed [`W-1:0] ir7_i48;
  wire signed [`W-1:0] ir7_i49;
  wire signed [`W-1:0] ir7_i50;
  wire signed [`W-1:0] ir7_i51;
  wire signed [`W-1:0] ir7_i52;
  wire signed [`W-1:0] ir7_i53;
  wire signed [`W-1:0] ir7_i54;
  wire signed [`W-1:0] ir7_i55;
  wire signed [`W-1:0] ir7_i56;
  wire signed [`W-1:0] ir7_i57;
  wire signed [`W-1:0] ir7_i58;
  wire signed [`W-1:0] ir7_i59;
  wire signed [`W-1:0] ir7_i60;
  wire signed [`W-1:0] ir7_v;
  wire signed [`W-1:0] ir5_i0;
  wire signed [`W-1:0] ir5_i1;
  wire signed [`W-1:0] ir5_i2;
  wire signed [`W-1:0] ir5_i3;
  wire signed [`W-1:0] ir5_i4;
  wire signed [`W-1:0] ir5_i5;
  wire signed [`W-1:0] ir5_i6;
  wire signed [`W-1:0] ir5_i7;
  wire signed [`W-1:0] ir5_i8;
  wire signed [`W-1:0] ir5_i9;
  wire signed [`W-1:0] ir5_i10;
  wire signed [`W-1:0] ir5_i11;
  wire signed [`W-1:0] ir5_i12;
  wire signed [`W-1:0] ir5_i13;
  wire signed [`W-1:0] ir5_i14;
  wire signed [`W-1:0] ir5_i15;
  wire signed [`W-1:0] ir5_i16;
  wire signed [`W-1:0] ir5_i17;
  wire signed [`W-1:0] ir5_i18;
  wire signed [`W-1:0] ir5_i19;
  wire signed [`W-1:0] ir5_i20;
  wire signed [`W-1:0] ir5_i21;
  wire signed [`W-1:0] ir5_i22;
  wire signed [`W-1:0] ir5_i23;
  wire signed [`W-1:0] ir5_i24;
  wire signed [`W-1:0] ir5_i25;
  wire signed [`W-1:0] ir5_i26;
  wire signed [`W-1:0] ir5_i27;
  wire signed [`W-1:0] ir5_i28;
  wire signed [`W-1:0] ir5_i29;
  wire signed [`W-1:0] ir5_i30;
  wire signed [`W-1:0] ir5_i31;
  wire signed [`W-1:0] ir5_i32;
  wire signed [`W-1:0] ir5_i33;
  wire signed [`W-1:0] ir5_v;
  wire signed [`W-1:0] n5_i0;
  wire signed [`W-1:0] n5_i1;
  wire signed [`W-1:0] n5_i2;
  wire signed [`W-1:0] n5_v;
  wire signed [`W-1:0] n647_i0;
  wire signed [`W-1:0] n647_i1;
  wire signed [`W-1:0] n647_i2;
  wire signed [`W-1:0] n647_i3;
  wire signed [`W-1:0] n647_i4;
  wire signed [`W-1:0] n647_i5;
  wire signed [`W-1:0] n647_v;
  wire signed [`W-1:0] op_T2_ind_i0;
  wire signed [`W-1:0] op_T2_ind_i1;
  wire signed [`W-1:0] op_T2_ind_i2;
  wire signed [`W-1:0] op_T2_ind_v;
  wire signed [`W-1:0] n1257_i0;
  wire signed [`W-1:0] n1257_i1;
  wire signed [`W-1:0] n1257_i2;
  wire signed [`W-1:0] n1257_i3;
  wire signed [`W-1:0] n1257_i4;
  wire signed [`W-1:0] n1257_v;
  wire signed [`W-1:0] n1254_i0;
  wire signed [`W-1:0] n1254_i1;
  wire signed [`W-1:0] n1254_i2;
  wire signed [`W-1:0] n1254_i3;
  wire signed [`W-1:0] n1254_v;
  wire signed [`W-1:0] n1527_i0;
  wire signed [`W-1:0] n1527_i1;
  wire signed [`W-1:0] n1527_v;
  wire signed [`W-1:0] op_plp_pla_i0;
  wire signed [`W-1:0] op_plp_pla_i1;
  wire signed [`W-1:0] op_plp_pla_i2;
  wire signed [`W-1:0] op_plp_pla_v;
  wire signed [`W-1:0] n1253_i0;
  wire signed [`W-1:0] n1253_i1;
  wire signed [`W-1:0] n1253_i2;
  wire signed [`W-1:0] n1253_i3;
  wire signed [`W-1:0] n1253_i4;
  wire signed [`W-1:0] n1253_v;
  wire signed [`W-1:0] alua7_i0;
  wire signed [`W-1:0] alua7_i1;
  wire signed [`W-1:0] alua7_i2;
  wire signed [`W-1:0] alua7_i3;
  wire signed [`W-1:0] alua7_v;
  wire signed [`W-1:0] n1523_i0;
  wire signed [`W-1:0] n1523_i1;
  wire signed [`W-1:0] n1523_i2;
  wire signed [`W-1:0] n1523_i3;
  wire signed [`W-1:0] n1523_v;
  wire signed [`W-1:0] n1528_i0;
  wire signed [`W-1:0] n1528_i1;
  wire signed [`W-1:0] n1528_v;
  wire signed [`W-1:0] n1529_i0;
  wire signed [`W-1:0] n1529_i1;
  wire signed [`W-1:0] n1529_v;
  wire signed [`W-1:0] n1258_i0;
  wire signed [`W-1:0] n1258_i1;
  wire signed [`W-1:0] n1258_i2;
  wire signed [`W-1:0] n1258_i3;
  wire signed [`W-1:0] n1258_i4;
  wire signed [`W-1:0] n1258_i5;
  wire signed [`W-1:0] n1258_i6;
  wire signed [`W-1:0] n1258_i7;
  wire signed [`W-1:0] n1258_v;
  wire signed [`W-1:0] op_T4_ind_x_i0;
  wire signed [`W-1:0] op_T4_ind_x_i1;
  wire signed [`W-1:0] op_T4_ind_x_i2;
  wire signed [`W-1:0] op_T4_ind_x_i3;
  wire signed [`W-1:0] op_T4_ind_x_v;
  wire signed [`W-1:0] __AxB_4_i0;
  wire signed [`W-1:0] __AxB_4_i1;
  wire signed [`W-1:0] __AxB_4_i2;
  wire signed [`W-1:0] __AxB_4_i3;
  wire signed [`W-1:0] __AxB_4_i4;
  wire signed [`W-1:0] __AxB_4_v;
  wire signed [`W-1:0] op_T2_jmp_abs_i0;
  wire signed [`W-1:0] op_T2_jmp_abs_i1;
  wire signed [`W-1:0] op_T2_jmp_abs_i2;
  wire signed [`W-1:0] op_T2_jmp_abs_v;
  wire signed [`W-1:0] n300_i0;
  wire signed [`W-1:0] n300_i1;
  wire signed [`W-1:0] n300_i2;
  wire signed [`W-1:0] n300_v;
  wire signed [`W-1:0] op_T__cmp_i0;
  wire signed [`W-1:0] op_T__cmp_i1;
  wire signed [`W-1:0] op_T__cmp_i2;
  wire signed [`W-1:0] op_T__cmp_v;
  wire signed [`W-1:0] PD_xxx010x1_i0;
  wire signed [`W-1:0] PD_xxx010x1_i1;
  wire signed [`W-1:0] PD_xxx010x1_i2;
  wire signed [`W-1:0] PD_xxx010x1_v;
  wire signed [`W-1:0] op_T0_bit_i0;
  wire signed [`W-1:0] op_T0_bit_i1;
  wire signed [`W-1:0] op_T0_bit_i2;
  wire signed [`W-1:0] op_T0_bit_v;
  wire signed [`W-1:0] n304_i0;
  wire signed [`W-1:0] n304_i1;
  wire signed [`W-1:0] n304_i2;
  wire signed [`W-1:0] n304_i3;
  wire signed [`W-1:0] n304_i4;
  wire signed [`W-1:0] n304_i5;
  wire signed [`W-1:0] n304_v;
  wire signed [`W-1:0] y3_i0;
  wire signed [`W-1:0] y3_i1;
  wire signed [`W-1:0] y3_i2;
  wire signed [`W-1:0] y3_v;
  wire signed [`W-1:0] n306_i0;
  wire signed [`W-1:0] n306_i1;
  wire signed [`W-1:0] n306_i2;
  wire signed [`W-1:0] n306_v;
  wire signed [`W-1:0] n307_i0;
  wire signed [`W-1:0] n307_i1;
  wire signed [`W-1:0] n307_i2;
  wire signed [`W-1:0] n307_v;
  wire signed [`W-1:0] n473_i0;
  wire signed [`W-1:0] n473_i1;
  wire signed [`W-1:0] n473_i2;
  wire signed [`W-1:0] n473_v;
  wire signed [`W-1:0] DA_C01_i0;
  wire signed [`W-1:0] DA_C01_i1;
  wire signed [`W-1:0] DA_C01_i2;
  wire signed [`W-1:0] DA_C01_i3;
  wire signed [`W-1:0] DA_C01_v;
  wire signed [`W-1:0] n959_i0;
  wire signed [`W-1:0] n959_i1;
  wire signed [`W-1:0] n959_i2;
  wire signed [`W-1:0] n959_i3;
  wire signed [`W-1:0] n959_v;
  wire signed [`W-1:0] n958_i0;
  wire signed [`W-1:0] n958_i1;
  wire signed [`W-1:0] n958_i2;
  wire signed [`W-1:0] n958_i3;
  wire signed [`W-1:0] n958_v;
  wire signed [`W-1:0] n951_i0;
  wire signed [`W-1:0] n951_i1;
  wire signed [`W-1:0] n951_i2;
  wire signed [`W-1:0] n951_i3;
  wire signed [`W-1:0] n951_v;
  wire signed [`W-1:0] op_T__cpx_cpy_abs_i0;
  wire signed [`W-1:0] op_T__cpx_cpy_abs_i1;
  wire signed [`W-1:0] op_T__cpx_cpy_abs_i2;
  wire signed [`W-1:0] op_T__cpx_cpy_abs_v;
  wire signed [`W-1:0] n953_i0;
  wire signed [`W-1:0] n953_i1;
  wire signed [`W-1:0] n953_i2;
  wire signed [`W-1:0] n953_v;
  wire signed [`W-1:0] n952_i0;
  wire signed [`W-1:0] n952_i1;
  wire signed [`W-1:0] n952_i2;
  wire signed [`W-1:0] n952_i3;
  wire signed [`W-1:0] n952_v;
  wire signed [`W-1:0] pd2_i0;
  wire signed [`W-1:0] pd2_i1;
  wire signed [`W-1:0] pd2_v;
  wire signed [`W-1:0] n954_i0;
  wire signed [`W-1:0] n954_i1;
  wire signed [`W-1:0] n954_i2;
  wire signed [`W-1:0] n954_i3;
  wire signed [`W-1:0] n954_i4;
  wire signed [`W-1:0] n954_v;
  wire signed [`W-1:0] notaluoutmux0_i0;
  wire signed [`W-1:0] notaluoutmux0_i1;
  wire signed [`W-1:0] notaluoutmux0_i2;
  wire signed [`W-1:0] notaluoutmux0_i3;
  wire signed [`W-1:0] notaluoutmux0_i4;
  wire signed [`W-1:0] notaluoutmux0_i5;
  wire signed [`W-1:0] notaluoutmux0_v;
  wire signed [`W-1:0] n956_i0;
  wire signed [`W-1:0] n956_i1;
  wire signed [`W-1:0] n956_i2;
  wire signed [`W-1:0] n956_v;
  wire signed [`W-1:0] n507_i0;
  wire signed [`W-1:0] n507_i1;
  wire signed [`W-1:0] n507_i2;
  wire signed [`W-1:0] n507_i3;
  wire signed [`W-1:0] n507_v;
  wire signed [`W-1:0] dpc2_XSB_i0;
  wire signed [`W-1:0] dpc2_XSB_i1;
  wire signed [`W-1:0] dpc2_XSB_i2;
  wire signed [`W-1:0] dpc2_XSB_i3;
  wire signed [`W-1:0] dpc2_XSB_i4;
  wire signed [`W-1:0] dpc2_XSB_i5;
  wire signed [`W-1:0] dpc2_XSB_i6;
  wire signed [`W-1:0] dpc2_XSB_i7;
  wire signed [`W-1:0] dpc2_XSB_i8;
  wire signed [`W-1:0] dpc2_XSB_i9;
  wire signed [`W-1:0] dpc2_XSB_v;
  wire signed [`W-1:0] n666_i0;
  wire signed [`W-1:0] n666_i1;
  wire signed [`W-1:0] n666_v;
  wire signed [`W-1:0] n504_i0;
  wire signed [`W-1:0] n504_i1;
  wire signed [`W-1:0] n504_i2;
  wire signed [`W-1:0] n504_v;
  wire signed [`W-1:0] n1260_i0;
  wire signed [`W-1:0] n1260_i1;
  wire signed [`W-1:0] n1260_i2;
  wire signed [`W-1:0] n1260_i3;
  wire signed [`W-1:0] n1260_v;
  wire signed [`W-1:0] n719_i0;
  wire signed [`W-1:0] n719_i1;
  wire signed [`W-1:0] n719_i2;
  wire signed [`W-1:0] n719_i3;
  wire signed [`W-1:0] n719_v;
  wire signed [`W-1:0] n718_i0;
  wire signed [`W-1:0] n718_i1;
  wire signed [`W-1:0] n718_i2;
  wire signed [`W-1:0] n718_v;
  wire signed [`W-1:0] n717_i0;
  wire signed [`W-1:0] n717_i1;
  wire signed [`W-1:0] n717_i2;
  wire signed [`W-1:0] n717_i3;
  wire signed [`W-1:0] n717_v;
  wire signed [`W-1:0] n715_i0;
  wire signed [`W-1:0] n715_i1;
  wire signed [`W-1:0] n715_i2;
  wire signed [`W-1:0] n715_i3;
  wire signed [`W-1:0] n715_v;
  wire signed [`W-1:0] n714_i0;
  wire signed [`W-1:0] n714_i1;
  wire signed [`W-1:0] n714_i2;
  wire signed [`W-1:0] n714_v;
  wire signed [`W-1:0] abh1_i0;
  wire signed [`W-1:0] abh1_i1;
  wire signed [`W-1:0] abh1_i2;
  wire signed [`W-1:0] abh1_i3;
  wire signed [`W-1:0] abh1_i4;
  wire signed [`W-1:0] abh1_v;
  wire signed [`W-1:0] op_T2_jsr_i0;
  wire signed [`W-1:0] op_T2_jsr_i1;
  wire signed [`W-1:0] op_T2_jsr_i2;
  wire signed [`W-1:0] op_T2_jsr_i3;
  wire signed [`W-1:0] op_T2_jsr_i4;
  wire signed [`W-1:0] op_T2_jsr_v;
  wire signed [`W-1:0] cp1_i0;
  wire signed [`W-1:0] cp1_i1;
  wire signed [`W-1:0] cp1_i2;
  wire signed [`W-1:0] cp1_i3;
  wire signed [`W-1:0] cp1_i4;
  wire signed [`W-1:0] cp1_i5;
  wire signed [`W-1:0] cp1_i6;
  wire signed [`W-1:0] cp1_i7;
  wire signed [`W-1:0] cp1_i8;
  wire signed [`W-1:0] cp1_i9;
  wire signed [`W-1:0] cp1_i10;
  wire signed [`W-1:0] cp1_i11;
  wire signed [`W-1:0] cp1_i12;
  wire signed [`W-1:0] cp1_i13;
  wire signed [`W-1:0] cp1_i14;
  wire signed [`W-1:0] cp1_i15;
  wire signed [`W-1:0] cp1_i16;
  wire signed [`W-1:0] cp1_i17;
  wire signed [`W-1:0] cp1_i18;
  wire signed [`W-1:0] cp1_i19;
  wire signed [`W-1:0] cp1_i20;
  wire signed [`W-1:0] cp1_i21;
  wire signed [`W-1:0] cp1_i22;
  wire signed [`W-1:0] cp1_i23;
  wire signed [`W-1:0] cp1_i24;
  wire signed [`W-1:0] cp1_i25;
  wire signed [`W-1:0] cp1_i26;
  wire signed [`W-1:0] cp1_i27;
  wire signed [`W-1:0] cp1_i28;
  wire signed [`W-1:0] cp1_i29;
  wire signed [`W-1:0] cp1_i30;
  wire signed [`W-1:0] cp1_i31;
  wire signed [`W-1:0] cp1_i32;
  wire signed [`W-1:0] cp1_i33;
  wire signed [`W-1:0] cp1_i34;
  wire signed [`W-1:0] cp1_i35;
  wire signed [`W-1:0] cp1_i36;
  wire signed [`W-1:0] cp1_i37;
  wire signed [`W-1:0] cp1_i38;
  wire signed [`W-1:0] cp1_i39;
  wire signed [`W-1:0] cp1_i40;
  wire signed [`W-1:0] cp1_i41;
  wire signed [`W-1:0] cp1_i42;
  wire signed [`W-1:0] cp1_i43;
  wire signed [`W-1:0] cp1_i44;
  wire signed [`W-1:0] cp1_i45;
  wire signed [`W-1:0] cp1_i46;
  wire signed [`W-1:0] cp1_i47;
  wire signed [`W-1:0] cp1_i48;
  wire signed [`W-1:0] cp1_i49;
  wire signed [`W-1:0] cp1_i50;
  wire signed [`W-1:0] cp1_i51;
  wire signed [`W-1:0] cp1_i52;
  wire signed [`W-1:0] cp1_i53;
  wire signed [`W-1:0] cp1_i54;
  wire signed [`W-1:0] cp1_i55;
  wire signed [`W-1:0] cp1_i56;
  wire signed [`W-1:0] cp1_i57;
  wire signed [`W-1:0] cp1_i58;
  wire signed [`W-1:0] cp1_i59;
  wire signed [`W-1:0] cp1_i60;
  wire signed [`W-1:0] cp1_i61;
  wire signed [`W-1:0] cp1_i62;
  wire signed [`W-1:0] cp1_i63;
  wire signed [`W-1:0] cp1_i64;
  wire signed [`W-1:0] cp1_i65;
  wire signed [`W-1:0] cp1_i66;
  wire signed [`W-1:0] cp1_i67;
  wire signed [`W-1:0] cp1_i68;
  wire signed [`W-1:0] cp1_i69;
  wire signed [`W-1:0] cp1_i70;
  wire signed [`W-1:0] cp1_i71;
  wire signed [`W-1:0] cp1_i72;
  wire signed [`W-1:0] cp1_i73;
  wire signed [`W-1:0] cp1_i74;
  wire signed [`W-1:0] cp1_i75;
  wire signed [`W-1:0] cp1_i76;
  wire signed [`W-1:0] cp1_i77;
  wire signed [`W-1:0] cp1_i78;
  wire signed [`W-1:0] cp1_i79;
  wire signed [`W-1:0] cp1_i80;
  wire signed [`W-1:0] cp1_i81;
  wire signed [`W-1:0] cp1_i82;
  wire signed [`W-1:0] cp1_i83;
  wire signed [`W-1:0] cp1_i84;
  wire signed [`W-1:0] cp1_i85;
  wire signed [`W-1:0] cp1_i86;
  wire signed [`W-1:0] cp1_i87;
  wire signed [`W-1:0] cp1_i88;
  wire signed [`W-1:0] cp1_i89;
  wire signed [`W-1:0] cp1_i90;
  wire signed [`W-1:0] cp1_i91;
  wire signed [`W-1:0] cp1_i92;
  wire signed [`W-1:0] cp1_i93;
  wire signed [`W-1:0] cp1_i94;
  wire signed [`W-1:0] cp1_i95;
  wire signed [`W-1:0] cp1_i96;
  wire signed [`W-1:0] cp1_i97;
  wire signed [`W-1:0] cp1_i98;
  wire signed [`W-1:0] cp1_i99;
  wire signed [`W-1:0] cp1_i100;
  wire signed [`W-1:0] cp1_i101;
  wire signed [`W-1:0] cp1_i102;
  wire signed [`W-1:0] cp1_i103;
  wire signed [`W-1:0] cp1_v;
  wire signed [`W-1:0] n1265_i0;
  wire signed [`W-1:0] n1265_i1;
  wire signed [`W-1:0] n1265_i2;
  wire signed [`W-1:0] n1265_i3;
  wire signed [`W-1:0] n1265_v;
  wire signed [`W-1:0] n1069_i0;
  wire signed [`W-1:0] n1069_i1;
  wire signed [`W-1:0] n1069_i2;
  wire signed [`W-1:0] n1069_v;
  wire signed [`W-1:0] dpc8_nDBADD_i0;
  wire signed [`W-1:0] dpc8_nDBADD_i1;
  wire signed [`W-1:0] dpc8_nDBADD_i2;
  wire signed [`W-1:0] dpc8_nDBADD_i3;
  wire signed [`W-1:0] dpc8_nDBADD_i4;
  wire signed [`W-1:0] dpc8_nDBADD_i5;
  wire signed [`W-1:0] dpc8_nDBADD_i6;
  wire signed [`W-1:0] dpc8_nDBADD_i7;
  wire signed [`W-1:0] dpc8_nDBADD_i8;
  wire signed [`W-1:0] dpc8_nDBADD_i9;
  wire signed [`W-1:0] dpc8_nDBADD_v;
  wire signed [`W-1:0] n1061_i0;
  wire signed [`W-1:0] n1061_i1;
  wire signed [`W-1:0] n1061_v;
  wire signed [`W-1:0] dpc25_SBDB_i0;
  wire signed [`W-1:0] dpc25_SBDB_i1;
  wire signed [`W-1:0] dpc25_SBDB_i2;
  wire signed [`W-1:0] dpc25_SBDB_i3;
  wire signed [`W-1:0] dpc25_SBDB_i4;
  wire signed [`W-1:0] dpc25_SBDB_i5;
  wire signed [`W-1:0] dpc25_SBDB_i6;
  wire signed [`W-1:0] dpc25_SBDB_i7;
  wire signed [`W-1:0] dpc25_SBDB_i8;
  wire signed [`W-1:0] dpc25_SBDB_i9;
  wire signed [`W-1:0] dpc25_SBDB_v;
  wire signed [`W-1:0] n1063_i0;
  wire signed [`W-1:0] n1063_i1;
  wire signed [`W-1:0] n1063_i2;
  wire signed [`W-1:0] n1063_i3;
  wire signed [`W-1:0] n1063_i4;
  wire signed [`W-1:0] n1063_i5;
  wire signed [`W-1:0] n1063_v;
  wire signed [`W-1:0] _ABH0_i0;
  wire signed [`W-1:0] _ABH0_i1;
  wire signed [`W-1:0] _ABH0_i2;
  wire signed [`W-1:0] _ABH0_v;
  wire signed [`W-1:0] n1065_i0;
  wire signed [`W-1:0] n1065_i1;
  wire signed [`W-1:0] n1065_i2;
  wire signed [`W-1:0] n1065_v;
  wire signed [`W-1:0] nots1_i0;
  wire signed [`W-1:0] nots1_i1;
  wire signed [`W-1:0] nots1_v;
  wire signed [`W-1:0] n1067_i0;
  wire signed [`W-1:0] n1067_i1;
  wire signed [`W-1:0] n1067_i2;
  wire signed [`W-1:0] n1067_v;
  wire signed [`W-1:0] idl2_i0;
  wire signed [`W-1:0] idl2_i1;
  wire signed [`W-1:0] idl2_i2;
  wire signed [`W-1:0] idl2_v;
  wire signed [`W-1:0] pd6_i0;
  wire signed [`W-1:0] pd6_i1;
  wire signed [`W-1:0] pd6_v;
  wire signed [`W-1:0] n1668_i0;
  wire signed [`W-1:0] n1668_i1;
  wire signed [`W-1:0] n1668_i2;
  wire signed [`W-1:0] n1668_v;
  wire signed [`W-1:0] dpc16_EORS_i0;
  wire signed [`W-1:0] dpc16_EORS_i1;
  wire signed [`W-1:0] dpc16_EORS_i2;
  wire signed [`W-1:0] dpc16_EORS_i3;
  wire signed [`W-1:0] dpc16_EORS_i4;
  wire signed [`W-1:0] dpc16_EORS_i5;
  wire signed [`W-1:0] dpc16_EORS_i6;
  wire signed [`W-1:0] dpc16_EORS_i7;
  wire signed [`W-1:0] dpc16_EORS_i8;
  wire signed [`W-1:0] dpc16_EORS_i9;
  wire signed [`W-1:0] dpc16_EORS_v;
  wire signed [`W-1:0] op_T__asl_rol_a_i0;
  wire signed [`W-1:0] op_T__asl_rol_a_i1;
  wire signed [`W-1:0] op_T__asl_rol_a_i2;
  wire signed [`W-1:0] op_T__asl_rol_a_v;
  wire signed [`W-1:0] op_T__inx_i0;
  wire signed [`W-1:0] op_T__inx_i1;
  wire signed [`W-1:0] op_T__inx_i2;
  wire signed [`W-1:0] op_T__inx_v;
  wire signed [`W-1:0] n1662_i0;
  wire signed [`W-1:0] n1662_i1;
  wire signed [`W-1:0] n1662_i2;
  wire signed [`W-1:0] n1662_i3;
  wire signed [`W-1:0] n1662_v;
  wire signed [`W-1:0] n1661_i0;
  wire signed [`W-1:0] n1661_i1;
  wire signed [`W-1:0] n1661_i2;
  wire signed [`W-1:0] n1661_i3;
  wire signed [`W-1:0] n1661_v;
  wire signed [`W-1:0] n1660_i0;
  wire signed [`W-1:0] n1660_i1;
  wire signed [`W-1:0] n1660_i2;
  wire signed [`W-1:0] n1660_i3;
  wire signed [`W-1:0] n1660_v;
  wire signed [`W-1:0] n1087_i0;
  wire signed [`W-1:0] n1087_i1;
  wire signed [`W-1:0] n1087_i2;
  wire signed [`W-1:0] n1087_v;
  wire signed [`W-1:0] op_T2_pha_i0;
  wire signed [`W-1:0] op_T2_pha_i1;
  wire signed [`W-1:0] op_T2_pha_i2;
  wire signed [`W-1:0] op_T2_pha_v;
  wire signed [`W-1:0] n593_i0;
  wire signed [`W-1:0] n593_i1;
  wire signed [`W-1:0] n593_i2;
  wire signed [`W-1:0] n593_v;
  wire signed [`W-1:0] n1084_i0;
  wire signed [`W-1:0] n1084_i1;
  wire signed [`W-1:0] n1084_i2;
  wire signed [`W-1:0] n1084_i3;
  wire signed [`W-1:0] n1084_i4;
  wire signed [`W-1:0] n1084_v;
  wire signed [`W-1:0] n595_i0;
  wire signed [`W-1:0] n595_i1;
  wire signed [`W-1:0] n595_i2;
  wire signed [`W-1:0] n595_i3;
  wire signed [`W-1:0] n595_v;
  wire signed [`W-1:0] n1082_i0;
  wire signed [`W-1:0] n1082_i1;
  wire signed [`W-1:0] n1082_i2;
  wire signed [`W-1:0] n1082_v;
  wire signed [`W-1:0] n1081_i0;
  wire signed [`W-1:0] n1081_i1;
  wire signed [`W-1:0] n1081_i2;
  wire signed [`W-1:0] n1081_i3;
  wire signed [`W-1:0] n1081_v;
  wire signed [`W-1:0] n599_i0;
  wire signed [`W-1:0] n599_i1;
  wire signed [`W-1:0] n599_v;
  wire signed [`W-1:0] n598_i0;
  wire signed [`W-1:0] n598_i1;
  wire signed [`W-1:0] n598_v;
  wire signed [`W-1:0] n1089_i0;
  wire signed [`W-1:0] n1089_i1;
  wire signed [`W-1:0] n1089_i2;
  wire signed [`W-1:0] n1089_v;
  wire signed [`W-1:0] dor4_i0;
  wire signed [`W-1:0] dor4_i1;
  wire signed [`W-1:0] dor4_i2;
  wire signed [`W-1:0] dor4_i3;
  wire signed [`W-1:0] dor4_i4;
  wire signed [`W-1:0] dor4_v;
  wire signed [`W-1:0] n1409_i0;
  wire signed [`W-1:0] n1409_i1;
  wire signed [`W-1:0] n1409_v;
  wire signed [`W-1:0] n1408_i0;
  wire signed [`W-1:0] n1408_i1;
  wire signed [`W-1:0] n1408_i2;
  wire signed [`W-1:0] n1408_v;
  wire signed [`W-1:0] s0_i0;
  wire signed [`W-1:0] s0_i1;
  wire signed [`W-1:0] s0_i2;
  wire signed [`W-1:0] s0_v;
  wire signed [`W-1:0] n1402_i0;
  wire signed [`W-1:0] n1402_i1;
  wire signed [`W-1:0] n1402_i2;
  wire signed [`W-1:0] n1402_v;
  wire signed [`W-1:0] n1401_i0;
  wire signed [`W-1:0] n1401_i1;
  wire signed [`W-1:0] n1401_i2;
  wire signed [`W-1:0] n1401_v;
  wire signed [`W-1:0] n1400_i0;
  wire signed [`W-1:0] n1400_i1;
  wire signed [`W-1:0] n1400_i2;
  wire signed [`W-1:0] n1400_v;
  wire signed [`W-1:0] dasb4_i0;
  wire signed [`W-1:0] dasb4_i1;
  wire signed [`W-1:0] dasb4_i2;
  wire signed [`W-1:0] dasb4_i3;
  wire signed [`W-1:0] dasb4_i4;
  wire signed [`W-1:0] dasb4_i5;
  wire signed [`W-1:0] dasb4_i6;
  wire signed [`W-1:0] dasb4_i7;
  wire signed [`W-1:0] dasb4_i8;
  wire signed [`W-1:0] dasb4_i9;
  wire signed [`W-1:0] dasb4_i10;
  wire signed [`W-1:0] dasb4_i11;
  wire signed [`W-1:0] dasb4_i12;
  wire signed [`W-1:0] dasb4_v;
  wire signed [`W-1:0] n1404_i0;
  wire signed [`W-1:0] n1404_i1;
  wire signed [`W-1:0] n1404_v;
  wire signed [`W-1:0] pipephi2Reset0_i0;
  wire signed [`W-1:0] pipephi2Reset0_i1;
  wire signed [`W-1:0] pipephi2Reset0_v;
  wire signed [`W-1:0] x6_i0;
  wire signed [`W-1:0] x6_i1;
  wire signed [`W-1:0] x6_i2;
  wire signed [`W-1:0] x6_v;
  wire signed [`W-1:0] n1339_i0;
  wire signed [`W-1:0] n1339_i1;
  wire signed [`W-1:0] n1339_i2;
  wire signed [`W-1:0] n1339_v;
  wire signed [`W-1:0] n1338_i0;
  wire signed [`W-1:0] n1338_i1;
  wire signed [`W-1:0] n1338_v;
  wire signed [`W-1:0] aluaorb0_i0;
  wire signed [`W-1:0] aluaorb0_i1;
  wire signed [`W-1:0] aluaorb0_i2;
  wire signed [`W-1:0] aluaorb0_v;
  wire signed [`W-1:0] pipeUNK06_i0;
  wire signed [`W-1:0] pipeUNK06_i1;
  wire signed [`W-1:0] pipeUNK06_i2;
  wire signed [`W-1:0] pipeUNK06_v;
  wire signed [`W-1:0] n442_i0;
  wire signed [`W-1:0] n442_i1;
  wire signed [`W-1:0] n442_i2;
  wire signed [`W-1:0] n442_v;
  wire signed [`W-1:0] op_T0_cpx_cpy_inx_iny_i0;
  wire signed [`W-1:0] op_T0_cpx_cpy_inx_iny_i1;
  wire signed [`W-1:0] op_T0_cpx_cpy_inx_iny_i2;
  wire signed [`W-1:0] op_T0_cpx_cpy_inx_iny_v;
  wire signed [`W-1:0] sb6_i0;
  wire signed [`W-1:0] sb6_i1;
  wire signed [`W-1:0] sb6_i2;
  wire signed [`W-1:0] sb6_i3;
  wire signed [`W-1:0] sb6_i4;
  wire signed [`W-1:0] sb6_i5;
  wire signed [`W-1:0] sb6_i6;
  wire signed [`W-1:0] sb6_i7;
  wire signed [`W-1:0] sb6_i8;
  wire signed [`W-1:0] sb6_i9;
  wire signed [`W-1:0] sb6_i10;
  wire signed [`W-1:0] sb6_i11;
  wire signed [`W-1:0] sb6_i12;
  wire signed [`W-1:0] sb6_v;
  wire signed [`W-1:0] x_op_T3_abs_idx_i0;
  wire signed [`W-1:0] x_op_T3_abs_idx_i1;
  wire signed [`W-1:0] x_op_T3_abs_idx_i2;
  wire signed [`W-1:0] x_op_T3_abs_idx_v;
  wire signed [`W-1:0] op_T5_rti_rts_i0;
  wire signed [`W-1:0] op_T5_rti_rts_i1;
  wire signed [`W-1:0] op_T5_rti_rts_i2;
  wire signed [`W-1:0] op_T5_rti_rts_v;
  wire signed [`W-1:0] n445_i0;
  wire signed [`W-1:0] n445_i1;
  wire signed [`W-1:0] n445_i2;
  wire signed [`W-1:0] n445_i3;
  wire signed [`W-1:0] n445_i4;
  wire signed [`W-1:0] n445_v;
  wire signed [`W-1:0] alua2_i0;
  wire signed [`W-1:0] alua2_i1;
  wire signed [`W-1:0] alua2_i2;
  wire signed [`W-1:0] alua2_i3;
  wire signed [`W-1:0] alua2_v;
  wire signed [`W-1:0] n1545_i0;
  wire signed [`W-1:0] n1545_i1;
  wire signed [`W-1:0] n1545_i2;
  wire signed [`W-1:0] n1545_v;
  wire signed [`W-1:0] n1542_i0;
  wire signed [`W-1:0] n1542_i1;
  wire signed [`W-1:0] n1542_i2;
  wire signed [`W-1:0] n1542_i3;
  wire signed [`W-1:0] n1542_i4;
  wire signed [`W-1:0] n1542_v;
  wire signed [`W-1:0] x_op_T0_txa_i0;
  wire signed [`W-1:0] x_op_T0_txa_i1;
  wire signed [`W-1:0] x_op_T0_txa_i2;
  wire signed [`W-1:0] x_op_T0_txa_v;
  wire signed [`W-1:0] pclp4_i0;
  wire signed [`W-1:0] pclp4_i1;
  wire signed [`W-1:0] pclp4_i2;
  wire signed [`W-1:0] pclp4_v;
  wire signed [`W-1:0] n38_i0;
  wire signed [`W-1:0] n38_i1;
  wire signed [`W-1:0] n38_i2;
  wire signed [`W-1:0] n38_v;
  wire signed [`W-1:0] op_from_x_i0;
  wire signed [`W-1:0] op_from_x_i1;
  wire signed [`W-1:0] op_from_x_i2;
  wire signed [`W-1:0] op_from_x_i3;
  wire signed [`W-1:0] op_from_x_v;
  wire signed [`W-1:0] pchp5_i0;
  wire signed [`W-1:0] pchp5_i1;
  wire signed [`W-1:0] pchp5_i2;
  wire signed [`W-1:0] pchp5_v;
  wire signed [`W-1:0] p0_i0;
  wire signed [`W-1:0] p0_i1;
  wire signed [`W-1:0] p0_v;
  wire signed [`W-1:0] n31_i0;
  wire signed [`W-1:0] n31_i1;
  wire signed [`W-1:0] n31_i2;
  wire signed [`W-1:0] n31_i3;
  wire signed [`W-1:0] n31_i4;
  wire signed [`W-1:0] n31_i5;
  wire signed [`W-1:0] n31_i6;
  wire signed [`W-1:0] n31_v;
  wire signed [`W-1:0] n695_i0;
  wire signed [`W-1:0] n695_i1;
  wire signed [`W-1:0] n695_i2;
  wire signed [`W-1:0] n695_v;
  wire signed [`W-1:0] n37_i0;
  wire signed [`W-1:0] n37_i1;
  wire signed [`W-1:0] n37_i2;
  wire signed [`W-1:0] n37_v;
  wire signed [`W-1:0] n36_i0;
  wire signed [`W-1:0] n36_i1;
  wire signed [`W-1:0] n36_i2;
  wire signed [`W-1:0] n36_i3;
  wire signed [`W-1:0] n36_v;
  wire signed [`W-1:0] n35_i0;
  wire signed [`W-1:0] n35_i1;
  wire signed [`W-1:0] n35_i2;
  wire signed [`W-1:0] n35_i3;
  wire signed [`W-1:0] n35_v;
  wire signed [`W-1:0] n34_i0;
  wire signed [`W-1:0] n34_i1;
  wire signed [`W-1:0] n34_i2;
  wire signed [`W-1:0] n34_v;
  wire signed [`W-1:0] notidl6_i0;
  wire signed [`W-1:0] notidl6_i1;
  wire signed [`W-1:0] notidl6_v;
  wire signed [`W-1:0] AxB3_i0;
  wire signed [`W-1:0] AxB3_i1;
  wire signed [`W-1:0] AxB3_i2;
  wire signed [`W-1:0] AxB3_i3;
  wire signed [`W-1:0] AxB3_i4;
  wire signed [`W-1:0] AxB3_i5;
  wire signed [`W-1:0] AxB3_v;
  wire signed [`W-1:0] n643_i0;
  wire signed [`W-1:0] n643_i1;
  wire signed [`W-1:0] n643_i2;
  wire signed [`W-1:0] n643_v;
  wire signed [`W-1:0] n1534_i0;
  wire signed [`W-1:0] n1534_i1;
  wire signed [`W-1:0] n1534_i2;
  wire signed [`W-1:0] n1534_i3;
  wire signed [`W-1:0] n1534_v;
  wire signed [`W-1:0] n645_i0;
  wire signed [`W-1:0] n645_i1;
  wire signed [`W-1:0] n645_i2;
  wire signed [`W-1:0] n645_i3;
  wire signed [`W-1:0] n645_v;
  wire signed [`W-1:0] n1244_i0;
  wire signed [`W-1:0] n1244_i1;
  wire signed [`W-1:0] n1244_i2;
  wire signed [`W-1:0] n1244_v;
  wire signed [`W-1:0] n1531_i0;
  wire signed [`W-1:0] n1531_i1;
  wire signed [`W-1:0] n1531_i2;
  wire signed [`W-1:0] n1531_i3;
  wire signed [`W-1:0] n1531_v;
  wire signed [`W-1:0] n646_i0;
  wire signed [`W-1:0] n646_i1;
  wire signed [`W-1:0] n646_i2;
  wire signed [`W-1:0] n646_i3;
  wire signed [`W-1:0] n646_i4;
  wire signed [`W-1:0] n646_i5;
  wire signed [`W-1:0] n646_i6;
  wire signed [`W-1:0] n646_i7;
  wire signed [`W-1:0] n646_i8;
  wire signed [`W-1:0] n646_v;
  wire signed [`W-1:0] n649_i0;
  wire signed [`W-1:0] n649_i1;
  wire signed [`W-1:0] n649_i2;
  wire signed [`W-1:0] n649_i3;
  wire signed [`W-1:0] n649_i4;
  wire signed [`W-1:0] n649_v;
  wire signed [`W-1:0] alua1_i0;
  wire signed [`W-1:0] alua1_i1;
  wire signed [`W-1:0] alua1_i2;
  wire signed [`W-1:0] alua1_i3;
  wire signed [`W-1:0] alua1_v;
  wire signed [`W-1:0] adh7_i0;
  wire signed [`W-1:0] adh7_i1;
  wire signed [`W-1:0] adh7_i2;
  wire signed [`W-1:0] adh7_i3;
  wire signed [`W-1:0] adh7_i4;
  wire signed [`W-1:0] adh7_i5;
  wire signed [`W-1:0] adh7_i6;
  wire signed [`W-1:0] adh7_v;
  wire signed [`W-1:0] n339_i0;
  wire signed [`W-1:0] n339_i1;
  wire signed [`W-1:0] n339_v;
  wire signed [`W-1:0] pipeUNK08_i0;
  wire signed [`W-1:0] pipeUNK08_i1;
  wire signed [`W-1:0] pipeUNK08_v;
  wire signed [`W-1:0] n335_i0;
  wire signed [`W-1:0] n335_i1;
  wire signed [`W-1:0] n335_i2;
  wire signed [`W-1:0] n335_i3;
  wire signed [`W-1:0] n335_i4;
  wire signed [`W-1:0] n335_i5;
  wire signed [`W-1:0] n335_i6;
  wire signed [`W-1:0] n335_i7;
  wire signed [`W-1:0] n335_v;
  wire signed [`W-1:0] n334_i0;
  wire signed [`W-1:0] n334_i1;
  wire signed [`W-1:0] n334_i2;
  wire signed [`W-1:0] n334_i3;
  wire signed [`W-1:0] n334_i4;
  wire signed [`W-1:0] n334_v;
  wire signed [`W-1:0] ir6_i0;
  wire signed [`W-1:0] ir6_i1;
  wire signed [`W-1:0] ir6_i2;
  wire signed [`W-1:0] ir6_i3;
  wire signed [`W-1:0] ir6_i4;
  wire signed [`W-1:0] ir6_i5;
  wire signed [`W-1:0] ir6_i6;
  wire signed [`W-1:0] ir6_i7;
  wire signed [`W-1:0] ir6_i8;
  wire signed [`W-1:0] ir6_i9;
  wire signed [`W-1:0] ir6_i10;
  wire signed [`W-1:0] ir6_i11;
  wire signed [`W-1:0] ir6_i12;
  wire signed [`W-1:0] ir6_i13;
  wire signed [`W-1:0] ir6_i14;
  wire signed [`W-1:0] ir6_i15;
  wire signed [`W-1:0] ir6_i16;
  wire signed [`W-1:0] ir6_i17;
  wire signed [`W-1:0] ir6_i18;
  wire signed [`W-1:0] ir6_i19;
  wire signed [`W-1:0] ir6_i20;
  wire signed [`W-1:0] ir6_i21;
  wire signed [`W-1:0] ir6_i22;
  wire signed [`W-1:0] ir6_i23;
  wire signed [`W-1:0] ir6_i24;
  wire signed [`W-1:0] ir6_i25;
  wire signed [`W-1:0] ir6_i26;
  wire signed [`W-1:0] ir6_i27;
  wire signed [`W-1:0] ir6_i28;
  wire signed [`W-1:0] ir6_i29;
  wire signed [`W-1:0] ir6_i30;
  wire signed [`W-1:0] ir6_i31;
  wire signed [`W-1:0] ir6_i32;
  wire signed [`W-1:0] ir6_i33;
  wire signed [`W-1:0] ir6_i34;
  wire signed [`W-1:0] ir6_i35;
  wire signed [`W-1:0] ir6_i36;
  wire signed [`W-1:0] ir6_i37;
  wire signed [`W-1:0] ir6_i38;
  wire signed [`W-1:0] ir6_i39;
  wire signed [`W-1:0] ir6_i40;
  wire signed [`W-1:0] ir6_i41;
  wire signed [`W-1:0] ir6_i42;
  wire signed [`W-1:0] ir6_i43;
  wire signed [`W-1:0] ir6_v;
  wire signed [`W-1:0] n336_i0;
  wire signed [`W-1:0] n336_i1;
  wire signed [`W-1:0] n336_i2;
  wire signed [`W-1:0] n336_i3;
  wire signed [`W-1:0] n336_i4;
  wire signed [`W-1:0] n336_i5;
  wire signed [`W-1:0] n336_i6;
  wire signed [`W-1:0] n336_v;
  wire signed [`W-1:0] alu6_i0;
  wire signed [`W-1:0] alu6_i1;
  wire signed [`W-1:0] alu6_i2;
  wire signed [`W-1:0] alu6_i3;
  wire signed [`W-1:0] alu6_i4;
  wire signed [`W-1:0] alu6_v;
  wire signed [`W-1:0] n330_i0;
  wire signed [`W-1:0] n330_i1;
  wire signed [`W-1:0] n330_i2;
  wire signed [`W-1:0] n330_i3;
  wire signed [`W-1:0] n330_v;
  wire signed [`W-1:0] DC78_i0;
  wire signed [`W-1:0] DC78_i1;
  wire signed [`W-1:0] DC78_i2;
  wire signed [`W-1:0] DC78_v;
  wire signed [`W-1:0] n332_i0;
  wire signed [`W-1:0] n332_i1;
  wire signed [`W-1:0] n332_i2;
  wire signed [`W-1:0] n332_i3;
  wire signed [`W-1:0] n332_i4;
  wire signed [`W-1:0] n332_v;
  wire signed [`W-1:0] n1026_i0;
  wire signed [`W-1:0] n1026_i1;
  wire signed [`W-1:0] n1026_i2;
  wire signed [`W-1:0] n1026_i3;
  wire signed [`W-1:0] n1026_v;
  wire signed [`W-1:0] n8_i0;
  wire signed [`W-1:0] n8_i1;
  wire signed [`W-1:0] n8_i2;
  wire signed [`W-1:0] n8_i3;
  wire signed [`W-1:0] n8_i4;
  wire signed [`W-1:0] n8_v;
  wire signed [`W-1:0] n1462_i0;
  wire signed [`W-1:0] n1462_i1;
  wire signed [`W-1:0] n1462_i2;
  wire signed [`W-1:0] n1462_v;
  wire signed [`W-1:0] INTG_i0;
  wire signed [`W-1:0] INTG_i1;
  wire signed [`W-1:0] INTG_i2;
  wire signed [`W-1:0] INTG_i3;
  wire signed [`W-1:0] INTG_v;
  wire signed [`W-1:0] pch4_i0;
  wire signed [`W-1:0] pch4_i1;
  wire signed [`W-1:0] pch4_i2;
  wire signed [`W-1:0] pch4_v;
  wire signed [`W-1:0] n946_i0;
  wire signed [`W-1:0] n946_i1;
  wire signed [`W-1:0] n946_i2;
  wire signed [`W-1:0] n946_v;
  wire signed [`W-1:0] n947_i0;
  wire signed [`W-1:0] n947_i1;
  wire signed [`W-1:0] n947_i2;
  wire signed [`W-1:0] n947_v;
  wire signed [`W-1:0] n944_i0;
  wire signed [`W-1:0] n944_i1;
  wire signed [`W-1:0] n944_i2;
  wire signed [`W-1:0] n944_v;
  wire signed [`W-1:0] db2_i0;
  wire signed [`W-1:0] db2_i1;
  wire signed [`W-1:0] db2_i2;
  wire signed [`W-1:0] db2_i3;
  wire signed [`W-1:0] db2_i4;
  wire signed [`W-1:0] db2_v;
  wire signed [`W-1:0] cclk_i0;
  wire signed [`W-1:0] cclk_i1;
  wire signed [`W-1:0] cclk_i2;
  wire signed [`W-1:0] cclk_i3;
  wire signed [`W-1:0] cclk_i4;
  wire signed [`W-1:0] cclk_i5;
  wire signed [`W-1:0] cclk_i6;
  wire signed [`W-1:0] cclk_i7;
  wire signed [`W-1:0] cclk_i8;
  wire signed [`W-1:0] cclk_i9;
  wire signed [`W-1:0] cclk_i10;
  wire signed [`W-1:0] cclk_i11;
  wire signed [`W-1:0] cclk_i12;
  wire signed [`W-1:0] cclk_i13;
  wire signed [`W-1:0] cclk_i14;
  wire signed [`W-1:0] cclk_i15;
  wire signed [`W-1:0] cclk_i16;
  wire signed [`W-1:0] cclk_i17;
  wire signed [`W-1:0] cclk_i18;
  wire signed [`W-1:0] cclk_i19;
  wire signed [`W-1:0] cclk_i20;
  wire signed [`W-1:0] cclk_i21;
  wire signed [`W-1:0] cclk_i22;
  wire signed [`W-1:0] cclk_i23;
  wire signed [`W-1:0] cclk_i24;
  wire signed [`W-1:0] cclk_i25;
  wire signed [`W-1:0] cclk_i26;
  wire signed [`W-1:0] cclk_i27;
  wire signed [`W-1:0] cclk_i28;
  wire signed [`W-1:0] cclk_i29;
  wire signed [`W-1:0] cclk_i30;
  wire signed [`W-1:0] cclk_i31;
  wire signed [`W-1:0] cclk_i32;
  wire signed [`W-1:0] cclk_i33;
  wire signed [`W-1:0] cclk_i34;
  wire signed [`W-1:0] cclk_i35;
  wire signed [`W-1:0] cclk_i36;
  wire signed [`W-1:0] cclk_i37;
  wire signed [`W-1:0] cclk_i38;
  wire signed [`W-1:0] cclk_i39;
  wire signed [`W-1:0] cclk_i40;
  wire signed [`W-1:0] cclk_i41;
  wire signed [`W-1:0] cclk_i42;
  wire signed [`W-1:0] cclk_i43;
  wire signed [`W-1:0] cclk_i44;
  wire signed [`W-1:0] cclk_i45;
  wire signed [`W-1:0] cclk_i46;
  wire signed [`W-1:0] cclk_i47;
  wire signed [`W-1:0] cclk_i48;
  wire signed [`W-1:0] cclk_i49;
  wire signed [`W-1:0] cclk_i50;
  wire signed [`W-1:0] cclk_i51;
  wire signed [`W-1:0] cclk_i52;
  wire signed [`W-1:0] cclk_i53;
  wire signed [`W-1:0] cclk_i54;
  wire signed [`W-1:0] cclk_i55;
  wire signed [`W-1:0] cclk_i56;
  wire signed [`W-1:0] cclk_i57;
  wire signed [`W-1:0] cclk_i58;
  wire signed [`W-1:0] cclk_i59;
  wire signed [`W-1:0] cclk_i60;
  wire signed [`W-1:0] cclk_i61;
  wire signed [`W-1:0] cclk_i62;
  wire signed [`W-1:0] cclk_i63;
  wire signed [`W-1:0] cclk_i64;
  wire signed [`W-1:0] cclk_i65;
  wire signed [`W-1:0] cclk_i66;
  wire signed [`W-1:0] cclk_i67;
  wire signed [`W-1:0] cclk_i68;
  wire signed [`W-1:0] cclk_i69;
  wire signed [`W-1:0] cclk_i70;
  wire signed [`W-1:0] cclk_i71;
  wire signed [`W-1:0] cclk_i72;
  wire signed [`W-1:0] cclk_i73;
  wire signed [`W-1:0] cclk_i74;
  wire signed [`W-1:0] cclk_i75;
  wire signed [`W-1:0] cclk_i76;
  wire signed [`W-1:0] cclk_i77;
  wire signed [`W-1:0] cclk_i78;
  wire signed [`W-1:0] cclk_i79;
  wire signed [`W-1:0] cclk_i80;
  wire signed [`W-1:0] cclk_i81;
  wire signed [`W-1:0] cclk_i82;
  wire signed [`W-1:0] cclk_i83;
  wire signed [`W-1:0] cclk_i84;
  wire signed [`W-1:0] cclk_i85;
  wire signed [`W-1:0] cclk_i86;
  wire signed [`W-1:0] cclk_i87;
  wire signed [`W-1:0] cclk_i88;
  wire signed [`W-1:0] cclk_i89;
  wire signed [`W-1:0] cclk_i90;
  wire signed [`W-1:0] cclk_i91;
  wire signed [`W-1:0] cclk_i92;
  wire signed [`W-1:0] cclk_i93;
  wire signed [`W-1:0] cclk_i94;
  wire signed [`W-1:0] cclk_i95;
  wire signed [`W-1:0] cclk_i96;
  wire signed [`W-1:0] cclk_i97;
  wire signed [`W-1:0] cclk_i98;
  wire signed [`W-1:0] cclk_i99;
  wire signed [`W-1:0] cclk_i100;
  wire signed [`W-1:0] cclk_i101;
  wire signed [`W-1:0] cclk_i102;
  wire signed [`W-1:0] cclk_i103;
  wire signed [`W-1:0] cclk_i104;
  wire signed [`W-1:0] cclk_i105;
  wire signed [`W-1:0] cclk_i106;
  wire signed [`W-1:0] cclk_i107;
  wire signed [`W-1:0] cclk_i108;
  wire signed [`W-1:0] cclk_i109;
  wire signed [`W-1:0] cclk_i110;
  wire signed [`W-1:0] cclk_i111;
  wire signed [`W-1:0] cclk_i112;
  wire signed [`W-1:0] cclk_i113;
  wire signed [`W-1:0] cclk_i114;
  wire signed [`W-1:0] cclk_i115;
  wire signed [`W-1:0] cclk_i116;
  wire signed [`W-1:0] cclk_i117;
  wire signed [`W-1:0] cclk_i118;
  wire signed [`W-1:0] cclk_i119;
  wire signed [`W-1:0] cclk_i120;
  wire signed [`W-1:0] cclk_i121;
  wire signed [`W-1:0] cclk_i122;
  wire signed [`W-1:0] cclk_i123;
  wire signed [`W-1:0] cclk_i124;
  wire signed [`W-1:0] cclk_i125;
  wire signed [`W-1:0] cclk_i126;
  wire signed [`W-1:0] cclk_i127;
  wire signed [`W-1:0] cclk_i128;
  wire signed [`W-1:0] cclk_i129;
  wire signed [`W-1:0] cclk_i130;
  wire signed [`W-1:0] cclk_i131;
  wire signed [`W-1:0] cclk_i132;
  wire signed [`W-1:0] cclk_i133;
  wire signed [`W-1:0] cclk_i134;
  wire signed [`W-1:0] cclk_i135;
  wire signed [`W-1:0] cclk_i136;
  wire signed [`W-1:0] cclk_i137;
  wire signed [`W-1:0] cclk_i138;
  wire signed [`W-1:0] cclk_i139;
  wire signed [`W-1:0] cclk_i140;
  wire signed [`W-1:0] cclk_i141;
  wire signed [`W-1:0] cclk_i142;
  wire signed [`W-1:0] cclk_i143;
  wire signed [`W-1:0] cclk_i144;
  wire signed [`W-1:0] cclk_i145;
  wire signed [`W-1:0] cclk_i146;
  wire signed [`W-1:0] cclk_i147;
  wire signed [`W-1:0] cclk_i148;
  wire signed [`W-1:0] cclk_i149;
  wire signed [`W-1:0] cclk_i150;
  wire signed [`W-1:0] cclk_i151;
  wire signed [`W-1:0] cclk_i152;
  wire signed [`W-1:0] cclk_i153;
  wire signed [`W-1:0] cclk_i154;
  wire signed [`W-1:0] cclk_i155;
  wire signed [`W-1:0] cclk_i156;
  wire signed [`W-1:0] cclk_i157;
  wire signed [`W-1:0] cclk_i158;
  wire signed [`W-1:0] cclk_i159;
  wire signed [`W-1:0] cclk_i160;
  wire signed [`W-1:0] cclk_i161;
  wire signed [`W-1:0] cclk_i162;
  wire signed [`W-1:0] cclk_i163;
  wire signed [`W-1:0] cclk_i164;
  wire signed [`W-1:0] cclk_i165;
  wire signed [`W-1:0] cclk_i166;
  wire signed [`W-1:0] cclk_i167;
  wire signed [`W-1:0] cclk_i168;
  wire signed [`W-1:0] cclk_i169;
  wire signed [`W-1:0] cclk_i170;
  wire signed [`W-1:0] cclk_i171;
  wire signed [`W-1:0] cclk_i172;
  wire signed [`W-1:0] cclk_i173;
  wire signed [`W-1:0] cclk_i174;
  wire signed [`W-1:0] cclk_i175;
  wire signed [`W-1:0] cclk_i176;
  wire signed [`W-1:0] cclk_i177;
  wire signed [`W-1:0] cclk_i178;
  wire signed [`W-1:0] cclk_i179;
  wire signed [`W-1:0] cclk_i180;
  wire signed [`W-1:0] cclk_i181;
  wire signed [`W-1:0] cclk_i182;
  wire signed [`W-1:0] cclk_i183;
  wire signed [`W-1:0] cclk_i184;
  wire signed [`W-1:0] cclk_i185;
  wire signed [`W-1:0] cclk_i186;
  wire signed [`W-1:0] cclk_i187;
  wire signed [`W-1:0] cclk_i188;
  wire signed [`W-1:0] cclk_i189;
  wire signed [`W-1:0] cclk_i190;
  wire signed [`W-1:0] cclk_i191;
  wire signed [`W-1:0] cclk_i192;
  wire signed [`W-1:0] cclk_i193;
  wire signed [`W-1:0] cclk_i194;
  wire signed [`W-1:0] cclk_i195;
  wire signed [`W-1:0] cclk_i196;
  wire signed [`W-1:0] cclk_i197;
  wire signed [`W-1:0] cclk_i198;
  wire signed [`W-1:0] cclk_i199;
  wire signed [`W-1:0] cclk_i200;
  wire signed [`W-1:0] cclk_i201;
  wire signed [`W-1:0] cclk_i202;
  wire signed [`W-1:0] cclk_i203;
  wire signed [`W-1:0] cclk_i204;
  wire signed [`W-1:0] cclk_i205;
  wire signed [`W-1:0] cclk_i206;
  wire signed [`W-1:0] cclk_i207;
  wire signed [`W-1:0] cclk_i208;
  wire signed [`W-1:0] cclk_i209;
  wire signed [`W-1:0] cclk_i210;
  wire signed [`W-1:0] cclk_i211;
  wire signed [`W-1:0] cclk_i212;
  wire signed [`W-1:0] cclk_i213;
  wire signed [`W-1:0] cclk_i214;
  wire signed [`W-1:0] cclk_i215;
  wire signed [`W-1:0] cclk_i216;
  wire signed [`W-1:0] cclk_i217;
  wire signed [`W-1:0] cclk_i218;
  wire signed [`W-1:0] cclk_i219;
  wire signed [`W-1:0] cclk_i220;
  wire signed [`W-1:0] cclk_i221;
  wire signed [`W-1:0] cclk_i222;
  wire signed [`W-1:0] cclk_i223;
  wire signed [`W-1:0] cclk_i224;
  wire signed [`W-1:0] cclk_i225;
  wire signed [`W-1:0] cclk_i226;
  wire signed [`W-1:0] cclk_i227;
  wire signed [`W-1:0] cclk_i228;
  wire signed [`W-1:0] cclk_i229;
  wire signed [`W-1:0] cclk_i230;
  wire signed [`W-1:0] cclk_i231;
  wire signed [`W-1:0] cclk_i232;
  wire signed [`W-1:0] cclk_i233;
  wire signed [`W-1:0] cclk_i234;
  wire signed [`W-1:0] cclk_i235;
  wire signed [`W-1:0] cclk_i236;
  wire signed [`W-1:0] cclk_i237;
  wire signed [`W-1:0] cclk_i238;
  wire signed [`W-1:0] cclk_i239;
  wire signed [`W-1:0] cclk_i240;
  wire signed [`W-1:0] cclk_i241;
  wire signed [`W-1:0] cclk_i242;
  wire signed [`W-1:0] cclk_i243;
  wire signed [`W-1:0] cclk_i244;
  wire signed [`W-1:0] cclk_i245;
  wire signed [`W-1:0] cclk_i246;
  wire signed [`W-1:0] cclk_i247;
  wire signed [`W-1:0] cclk_i248;
  wire signed [`W-1:0] cclk_i249;
  wire signed [`W-1:0] cclk_i250;
  wire signed [`W-1:0] cclk_i251;
  wire signed [`W-1:0] cclk_i252;
  wire signed [`W-1:0] cclk_i253;
  wire signed [`W-1:0] cclk_i254;
  wire signed [`W-1:0] cclk_i255;
  wire signed [`W-1:0] cclk_i256;
  wire signed [`W-1:0] cclk_i257;
  wire signed [`W-1:0] cclk_i258;
  wire signed [`W-1:0] cclk_i259;
  wire signed [`W-1:0] cclk_i260;
  wire signed [`W-1:0] cclk_i261;
  wire signed [`W-1:0] cclk_i262;
  wire signed [`W-1:0] cclk_i263;
  wire signed [`W-1:0] cclk_i264;
  wire signed [`W-1:0] cclk_i265;
  wire signed [`W-1:0] cclk_i266;
  wire signed [`W-1:0] cclk_i267;
  wire signed [`W-1:0] cclk_i268;
  wire signed [`W-1:0] cclk_i269;
  wire signed [`W-1:0] cclk_i270;
  wire signed [`W-1:0] cclk_i271;
  wire signed [`W-1:0] cclk_i272;
  wire signed [`W-1:0] cclk_i273;
  wire signed [`W-1:0] cclk_i274;
  wire signed [`W-1:0] cclk_v;
  wire signed [`W-1:0] pipeT5out_i0;
  wire signed [`W-1:0] pipeT5out_i1;
  wire signed [`W-1:0] pipeT5out_v;
  wire signed [`W-1:0] n133_i0;
  wire signed [`W-1:0] n133_i1;
  wire signed [`W-1:0] n133_i2;
  wire signed [`W-1:0] n133_i3;
  wire signed [`W-1:0] n133_v;
  wire signed [`W-1:0] n132_i0;
  wire signed [`W-1:0] n132_i1;
  wire signed [`W-1:0] n132_i2;
  wire signed [`W-1:0] n132_v;
  wire signed [`W-1:0] op_T0_pla_i0;
  wire signed [`W-1:0] op_T0_pla_i1;
  wire signed [`W-1:0] op_T0_pla_i2;
  wire signed [`W-1:0] op_T0_pla_v;
  wire signed [`W-1:0] n130_i0;
  wire signed [`W-1:0] n130_i1;
  wire signed [`W-1:0] n130_i2;
  wire signed [`W-1:0] n130_v;
  wire signed [`W-1:0] n135_i0;
  wire signed [`W-1:0] n135_i1;
  wire signed [`W-1:0] n135_i2;
  wire signed [`W-1:0] n135_v;
  wire signed [`W-1:0] n134_i0;
  wire signed [`W-1:0] n134_i1;
  wire signed [`W-1:0] n134_i2;
  wire signed [`W-1:0] n134_i3;
  wire signed [`W-1:0] n134_v;
  wire signed [`W-1:0] n139_i0;
  wire signed [`W-1:0] n139_i1;
  wire signed [`W-1:0] n139_i2;
  wire signed [`W-1:0] n139_v;
  wire signed [`W-1:0] n138_i0;
  wire signed [`W-1:0] n138_i1;
  wire signed [`W-1:0] n138_i2;
  wire signed [`W-1:0] n138_i3;
  wire signed [`W-1:0] n138_v;
  wire signed [`W-1:0] n708_i0;
  wire signed [`W-1:0] n708_i1;
  wire signed [`W-1:0] n708_i2;
  wire signed [`W-1:0] n708_v;
  wire signed [`W-1:0] n709_i0;
  wire signed [`W-1:0] n709_i1;
  wire signed [`W-1:0] n709_i2;
  wire signed [`W-1:0] n709_v;
  wire signed [`W-1:0] alub2_i0;
  wire signed [`W-1:0] alub2_i1;
  wire signed [`W-1:0] alub2_i2;
  wire signed [`W-1:0] alub2_i3;
  wire signed [`W-1:0] alub2_i4;
  wire signed [`W-1:0] alub2_v;
  wire signed [`W-1:0] pipeT3out_i0;
  wire signed [`W-1:0] pipeT3out_i1;
  wire signed [`W-1:0] pipeT3out_i2;
  wire signed [`W-1:0] pipeT3out_v;
  wire signed [`W-1:0] _ABL2_i0;
  wire signed [`W-1:0] _ABL2_i1;
  wire signed [`W-1:0] _ABL2_i2;
  wire signed [`W-1:0] _ABL2_v;
  wire signed [`W-1:0] n700_i0;
  wire signed [`W-1:0] n700_i1;
  wire signed [`W-1:0] n700_i2;
  wire signed [`W-1:0] n700_i3;
  wire signed [`W-1:0] n700_v;
  wire signed [`W-1:0] __AxB_2_i0;
  wire signed [`W-1:0] __AxB_2_i1;
  wire signed [`W-1:0] __AxB_2_i2;
  wire signed [`W-1:0] __AxB_2_i3;
  wire signed [`W-1:0] __AxB_2_i4;
  wire signed [`W-1:0] __AxB_2_v;
  wire signed [`W-1:0] notir1_i0;
  wire signed [`W-1:0] notir1_i1;
  wire signed [`W-1:0] notir1_i2;
  wire signed [`W-1:0] notir1_i3;
  wire signed [`W-1:0] notir1_i4;
  wire signed [`W-1:0] notir1_i5;
  wire signed [`W-1:0] notir1_i6;
  wire signed [`W-1:0] notir1_i7;
  wire signed [`W-1:0] notir1_i8;
  wire signed [`W-1:0] notir1_i9;
  wire signed [`W-1:0] notir1_i10;
  wire signed [`W-1:0] notir1_i11;
  wire signed [`W-1:0] notir1_i12;
  wire signed [`W-1:0] notir1_i13;
  wire signed [`W-1:0] notir1_i14;
  wire signed [`W-1:0] notir1_i15;
  wire signed [`W-1:0] notir1_i16;
  wire signed [`W-1:0] notir1_i17;
  wire signed [`W-1:0] notir1_i18;
  wire signed [`W-1:0] notir1_i19;
  wire signed [`W-1:0] notir1_i20;
  wire signed [`W-1:0] notir1_i21;
  wire signed [`W-1:0] notir1_i22;
  wire signed [`W-1:0] notir1_i23;
  wire signed [`W-1:0] notir1_v;
  wire signed [`W-1:0] n88_i0;
  wire signed [`W-1:0] n88_i1;
  wire signed [`W-1:0] n88_v;
  wire signed [`W-1:0] rdy_i0;
  wire signed [`W-1:0] rdy_i1;
  wire signed [`W-1:0] rdy_i2;
  wire signed [`W-1:0] rdy_v;
  wire signed [`W-1:0] db1_i0;
  wire signed [`W-1:0] db1_i1;
  wire signed [`W-1:0] db1_i2;
  wire signed [`W-1:0] db1_i3;
  wire signed [`W-1:0] db1_i4;
  wire signed [`W-1:0] db1_v;
  wire signed [`W-1:0] n83_i0;
  wire signed [`W-1:0] n83_i1;
  wire signed [`W-1:0] n83_i2;
  wire signed [`W-1:0] n83_i3;
  wire signed [`W-1:0] n83_v;
  wire signed [`W-1:0] n80_i0;
  wire signed [`W-1:0] n80_i1;
  wire signed [`W-1:0] n80_i2;
  wire signed [`W-1:0] n80_v;
  wire signed [`W-1:0] s2_i0;
  wire signed [`W-1:0] s2_i1;
  wire signed [`W-1:0] s2_i2;
  wire signed [`W-1:0] s2_v;
  wire signed [`W-1:0] n86_i0;
  wire signed [`W-1:0] n86_i1;
  wire signed [`W-1:0] n86_i2;
  wire signed [`W-1:0] n86_i3;
  wire signed [`W-1:0] n86_v;
  wire signed [`W-1:0] n87_i0;
  wire signed [`W-1:0] n87_i1;
  wire signed [`W-1:0] n87_i2;
  wire signed [`W-1:0] n87_i3;
  wire signed [`W-1:0] n87_v;
  wire signed [`W-1:0] op_T2_ind_x_i0;
  wire signed [`W-1:0] op_T2_ind_x_i1;
  wire signed [`W-1:0] op_T2_ind_x_i2;
  wire signed [`W-1:0] op_T2_ind_x_v;
  wire signed [`W-1:0] x4_i0;
  wire signed [`W-1:0] x4_i1;
  wire signed [`W-1:0] x4_i2;
  wire signed [`W-1:0] x4_v;
  wire signed [`W-1:0] op_T0_cpx_inx_i0;
  wire signed [`W-1:0] op_T0_cpx_inx_i1;
  wire signed [`W-1:0] op_T0_cpx_inx_i2;
  wire signed [`W-1:0] op_T0_cpx_inx_v;
  wire signed [`W-1:0] pipeUNK30_i0;
  wire signed [`W-1:0] pipeUNK30_i1;
  wire signed [`W-1:0] pipeUNK30_v;
  wire signed [`W-1:0] a7_i0;
  wire signed [`W-1:0] a7_i1;
  wire signed [`W-1:0] a7_i2;
  wire signed [`W-1:0] a7_v;
  wire signed [`W-1:0] n1650_i0;
  wire signed [`W-1:0] n1650_i1;
  wire signed [`W-1:0] n1650_i2;
  wire signed [`W-1:0] n1650_v;
  wire signed [`W-1:0] adh2_i0;
  wire signed [`W-1:0] adh2_i1;
  wire signed [`W-1:0] adh2_i2;
  wire signed [`W-1:0] adh2_i3;
  wire signed [`W-1:0] adh2_i4;
  wire signed [`W-1:0] adh2_i5;
  wire signed [`W-1:0] adh2_i6;
  wire signed [`W-1:0] adh2_v;
  wire signed [`W-1:0] n1657_i0;
  wire signed [`W-1:0] n1657_i1;
  wire signed [`W-1:0] n1657_i2;
  wire signed [`W-1:0] n1657_v;
  wire signed [`W-1:0] n1654_i0;
  wire signed [`W-1:0] n1654_i1;
  wire signed [`W-1:0] n1654_i2;
  wire signed [`W-1:0] n1654_i3;
  wire signed [`W-1:0] n1654_i4;
  wire signed [`W-1:0] n1654_v;
  wire signed [`W-1:0] n1655_i0;
  wire signed [`W-1:0] n1655_i1;
  wire signed [`W-1:0] n1655_i2;
  wire signed [`W-1:0] n1655_v;
  wire signed [`W-1:0] n586_i0;
  wire signed [`W-1:0] n586_i1;
  wire signed [`W-1:0] n586_i2;
  wire signed [`W-1:0] n586_v;
  wire signed [`W-1:0] n587_i0;
  wire signed [`W-1:0] n587_i1;
  wire signed [`W-1:0] n587_i2;
  wire signed [`W-1:0] n587_v;
  wire signed [`W-1:0] pch3_i0;
  wire signed [`W-1:0] pch3_i1;
  wire signed [`W-1:0] pch3_i2;
  wire signed [`W-1:0] pch3_v;
  wire signed [`W-1:0] n582_i0;
  wire signed [`W-1:0] n582_i1;
  wire signed [`W-1:0] n582_i2;
  wire signed [`W-1:0] n582_i3;
  wire signed [`W-1:0] n582_v;
  wire signed [`W-1:0] n583_i0;
  wire signed [`W-1:0] n583_i1;
  wire signed [`W-1:0] n583_i2;
  wire signed [`W-1:0] n583_v;
  wire signed [`W-1:0] n581_i0;
  wire signed [`W-1:0] n581_i1;
  wire signed [`W-1:0] n581_v;
  wire signed [`W-1:0] n588_i0;
  wire signed [`W-1:0] n588_i1;
  wire signed [`W-1:0] n588_i2;
  wire signed [`W-1:0] n588_v;
  wire signed [`W-1:0] x5_i0;
  wire signed [`W-1:0] x5_i1;
  wire signed [`W-1:0] x5_i2;
  wire signed [`W-1:0] x5_v;
  wire signed [`W-1:0] pipeUNK03_i0;
  wire signed [`W-1:0] pipeUNK03_i1;
  wire signed [`W-1:0] pipeUNK03_i2;
  wire signed [`W-1:0] pipeUNK03_v;
  wire signed [`W-1:0] adl4_i0;
  wire signed [`W-1:0] adl4_i1;
  wire signed [`W-1:0] adl4_i2;
  wire signed [`W-1:0] adl4_i3;
  wire signed [`W-1:0] adl4_i4;
  wire signed [`W-1:0] adl4_i5;
  wire signed [`W-1:0] adl4_i6;
  wire signed [`W-1:0] adl4_i7;
  wire signed [`W-1:0] adl4_v;
  wire signed [`W-1:0] n1434_i0;
  wire signed [`W-1:0] n1434_i1;
  wire signed [`W-1:0] n1434_i2;
  wire signed [`W-1:0] n1434_v;
  wire signed [`W-1:0] s7_i0;
  wire signed [`W-1:0] s7_i1;
  wire signed [`W-1:0] s7_i2;
  wire signed [`W-1:0] s7_v;
  wire signed [`W-1:0] alub1_i0;
  wire signed [`W-1:0] alub1_i1;
  wire signed [`W-1:0] alub1_i2;
  wire signed [`W-1:0] alub1_i3;
  wire signed [`W-1:0] alub1_i4;
  wire signed [`W-1:0] alub1_v;
  wire signed [`W-1:0] n1433_i0;
  wire signed [`W-1:0] n1433_i1;
  wire signed [`W-1:0] n1433_i2;
  wire signed [`W-1:0] n1433_v;
  wire signed [`W-1:0] x_op_T3_plp_pla_i0;
  wire signed [`W-1:0] x_op_T3_plp_pla_i1;
  wire signed [`W-1:0] x_op_T3_plp_pla_i2;
  wire signed [`W-1:0] x_op_T3_plp_pla_v;
  wire signed [`W-1:0] pipe_VEC_i0;
  wire signed [`W-1:0] pipe_VEC_i1;
  wire signed [`W-1:0] pipe_VEC_v;
  wire signed [`W-1:0] nots0_i0;
  wire signed [`W-1:0] nots0_i1;
  wire signed [`W-1:0] nots0_v;
  wire signed [`W-1:0] pipeUNK41_i0;
  wire signed [`W-1:0] pipeUNK41_i1;
  wire signed [`W-1:0] pipeUNK41_v;
  wire signed [`W-1:0] n1439_i0;
  wire signed [`W-1:0] n1439_i1;
  wire signed [`W-1:0] n1439_i2;
  wire signed [`W-1:0] n1439_v;
  wire signed [`W-1:0] db7_i0;
  wire signed [`W-1:0] db7_i1;
  wire signed [`W-1:0] db7_i2;
  wire signed [`W-1:0] db7_i3;
  wire signed [`W-1:0] db7_i4;
  wire signed [`W-1:0] db7_v;
  wire signed [`W-1:0] n459_i0;
  wire signed [`W-1:0] n459_i1;
  wire signed [`W-1:0] n459_v;
  wire signed [`W-1:0] dasb2_i0;
  wire signed [`W-1:0] dasb2_i1;
  wire signed [`W-1:0] dasb2_i2;
  wire signed [`W-1:0] dasb2_v;
  wire signed [`W-1:0] n1341_i0;
  wire signed [`W-1:0] n1341_i1;
  wire signed [`W-1:0] n1341_v;
  wire signed [`W-1:0] op_T0_acc_i0;
  wire signed [`W-1:0] op_T0_acc_i1;
  wire signed [`W-1:0] op_T0_acc_i2;
  wire signed [`W-1:0] op_T0_acc_v;
  wire signed [`W-1:0] n1343_i0;
  wire signed [`W-1:0] n1343_i1;
  wire signed [`W-1:0] n1343_i2;
  wire signed [`W-1:0] n1343_v;
  wire signed [`W-1:0] pipeUNK40_i0;
  wire signed [`W-1:0] pipeUNK40_i1;
  wire signed [`W-1:0] pipeUNK40_v;
  wire signed [`W-1:0] n457_i0;
  wire signed [`W-1:0] n457_i1;
  wire signed [`W-1:0] n457_i2;
  wire signed [`W-1:0] n457_v;
  wire signed [`W-1:0] n1377_i0;
  wire signed [`W-1:0] n1377_i1;
  wire signed [`W-1:0] n1377_i2;
  wire signed [`W-1:0] n1377_v;
  wire signed [`W-1:0] idb5_i0;
  wire signed [`W-1:0] idb5_i1;
  wire signed [`W-1:0] idb5_i2;
  wire signed [`W-1:0] idb5_i3;
  wire signed [`W-1:0] idb5_i4;
  wire signed [`W-1:0] idb5_i5;
  wire signed [`W-1:0] idb5_i6;
  wire signed [`W-1:0] idb5_i7;
  wire signed [`W-1:0] idb5_i8;
  wire signed [`W-1:0] idb5_i9;
  wire signed [`W-1:0] idb5_v;
  wire signed [`W-1:0] dpc7_SS_i0;
  wire signed [`W-1:0] dpc7_SS_i1;
  wire signed [`W-1:0] dpc7_SS_i2;
  wire signed [`W-1:0] dpc7_SS_i3;
  wire signed [`W-1:0] dpc7_SS_i4;
  wire signed [`W-1:0] dpc7_SS_i5;
  wire signed [`W-1:0] dpc7_SS_i6;
  wire signed [`W-1:0] dpc7_SS_i7;
  wire signed [`W-1:0] dpc7_SS_i8;
  wire signed [`W-1:0] dpc7_SS_i9;
  wire signed [`W-1:0] dpc7_SS_v;
  wire signed [`W-1:0] n1501_i0;
  wire signed [`W-1:0] n1501_i1;
  wire signed [`W-1:0] n1501_i2;
  wire signed [`W-1:0] n1501_v;
  wire signed [`W-1:0] _C01_i0;
  wire signed [`W-1:0] _C01_i1;
  wire signed [`W-1:0] _C01_i2;
  wire signed [`W-1:0] _C01_i3;
  wire signed [`W-1:0] _C01_v;
  wire signed [`W-1:0] n653_i0;
  wire signed [`W-1:0] n653_i1;
  wire signed [`W-1:0] n653_v;
  wire signed [`W-1:0] db3_i0;
  wire signed [`W-1:0] db3_i1;
  wire signed [`W-1:0] db3_i2;
  wire signed [`W-1:0] db3_i3;
  wire signed [`W-1:0] db3_i4;
  wire signed [`W-1:0] db3_v;
  wire signed [`W-1:0] __AxBxC_4_i0;
  wire signed [`W-1:0] __AxBxC_4_i1;
  wire signed [`W-1:0] __AxBxC_4_i2;
  wire signed [`W-1:0] __AxBxC_4_v;
  wire signed [`W-1:0] n1509_i0;
  wire signed [`W-1:0] n1509_i1;
  wire signed [`W-1:0] n1509_v;
  wire signed [`W-1:0] n658_i0;
  wire signed [`W-1:0] n658_i1;
  wire signed [`W-1:0] n658_i2;
  wire signed [`W-1:0] n658_i3;
  wire signed [`W-1:0] n658_v;
  wire signed [`W-1:0] DA_AxB2_i0;
  wire signed [`W-1:0] DA_AxB2_i1;
  wire signed [`W-1:0] DA_AxB2_i2;
  wire signed [`W-1:0] DA_AxB2_v;
  wire signed [`W-1:0] n55_i0;
  wire signed [`W-1:0] n55_i1;
  wire signed [`W-1:0] n55_v;
  wire signed [`W-1:0] n322_i0;
  wire signed [`W-1:0] n322_i1;
  wire signed [`W-1:0] n322_i2;
  wire signed [`W-1:0] n322_v;
  wire signed [`W-1:0] n323_i0;
  wire signed [`W-1:0] n323_i1;
  wire signed [`W-1:0] n323_v;
  wire signed [`W-1:0] n320_i0;
  wire signed [`W-1:0] n320_i1;
  wire signed [`W-1:0] n320_i2;
  wire signed [`W-1:0] n320_i3;
  wire signed [`W-1:0] n320_v;
  wire signed [`W-1:0] n321_i0;
  wire signed [`W-1:0] n321_i1;
  wire signed [`W-1:0] n321_i2;
  wire signed [`W-1:0] n321_i3;
  wire signed [`W-1:0] n321_v;
  wire signed [`W-1:0] n326_i0;
  wire signed [`W-1:0] n326_i1;
  wire signed [`W-1:0] n326_i2;
  wire signed [`W-1:0] n326_i3;
  wire signed [`W-1:0] n326_i4;
  wire signed [`W-1:0] n326_v;
  wire signed [`W-1:0] n327_i0;
  wire signed [`W-1:0] n327_i1;
  wire signed [`W-1:0] n327_i2;
  wire signed [`W-1:0] n327_v;
  wire signed [`W-1:0] op_inc_nop_i0;
  wire signed [`W-1:0] op_inc_nop_i1;
  wire signed [`W-1:0] op_inc_nop_i2;
  wire signed [`W-1:0] op_inc_nop_v;
  wire signed [`W-1:0] dpc1_SBY_i0;
  wire signed [`W-1:0] dpc1_SBY_i1;
  wire signed [`W-1:0] dpc1_SBY_i2;
  wire signed [`W-1:0] dpc1_SBY_i3;
  wire signed [`W-1:0] dpc1_SBY_i4;
  wire signed [`W-1:0] dpc1_SBY_i5;
  wire signed [`W-1:0] dpc1_SBY_i6;
  wire signed [`W-1:0] dpc1_SBY_i7;
  wire signed [`W-1:0] dpc1_SBY_i8;
  wire signed [`W-1:0] dpc1_SBY_i9;
  wire signed [`W-1:0] dpc1_SBY_v;
  wire signed [`W-1:0] ir0_i0;
  wire signed [`W-1:0] ir0_i1;
  wire signed [`W-1:0] ir0_i2;
  wire signed [`W-1:0] ir0_i3;
  wire signed [`W-1:0] ir0_i4;
  wire signed [`W-1:0] ir0_v;
  wire signed [`W-1:0] n329_i0;
  wire signed [`W-1:0] n329_i1;
  wire signed [`W-1:0] n329_i2;
  wire signed [`W-1:0] n329_i3;
  wire signed [`W-1:0] n329_v;
  wire signed [`W-1:0] ab2_i0;
  wire signed [`W-1:0] ab2_i1;
  wire signed [`W-1:0] ab2_i2;
  wire signed [`W-1:0] ab2_v;
  wire signed [`W-1:0] n1594_i0;
  wire signed [`W-1:0] n1594_i1;
  wire signed [`W-1:0] n1594_i2;
  wire signed [`W-1:0] n1594_v;
  wire signed [`W-1:0] n1592_i0;
  wire signed [`W-1:0] n1592_i1;
  wire signed [`W-1:0] n1592_i2;
  wire signed [`W-1:0] n1592_i3;
  wire signed [`W-1:0] n1592_i4;
  wire signed [`W-1:0] n1592_v;
  wire signed [`W-1:0] n995_i0;
  wire signed [`W-1:0] n995_i1;
  wire signed [`W-1:0] n995_i2;
  wire signed [`W-1:0] n995_v;
  wire signed [`W-1:0] n994_i0;
  wire signed [`W-1:0] n994_i1;
  wire signed [`W-1:0] n994_i2;
  wire signed [`W-1:0] n994_i3;
  wire signed [`W-1:0] n994_v;
  wire signed [`W-1:0] abh6_i0;
  wire signed [`W-1:0] abh6_i1;
  wire signed [`W-1:0] abh6_i2;
  wire signed [`W-1:0] abh6_i3;
  wire signed [`W-1:0] abh6_i4;
  wire signed [`W-1:0] abh6_v;
  wire signed [`W-1:0] irline3_i0;
  wire signed [`W-1:0] irline3_i1;
  wire signed [`W-1:0] irline3_i2;
  wire signed [`W-1:0] irline3_i3;
  wire signed [`W-1:0] irline3_i4;
  wire signed [`W-1:0] irline3_i5;
  wire signed [`W-1:0] irline3_i6;
  wire signed [`W-1:0] irline3_i7;
  wire signed [`W-1:0] irline3_i8;
  wire signed [`W-1:0] irline3_i9;
  wire signed [`W-1:0] irline3_i10;
  wire signed [`W-1:0] irline3_i11;
  wire signed [`W-1:0] irline3_i12;
  wire signed [`W-1:0] irline3_i13;
  wire signed [`W-1:0] irline3_i14;
  wire signed [`W-1:0] irline3_i15;
  wire signed [`W-1:0] irline3_i16;
  wire signed [`W-1:0] irline3_i17;
  wire signed [`W-1:0] irline3_i18;
  wire signed [`W-1:0] irline3_i19;
  wire signed [`W-1:0] irline3_i20;
  wire signed [`W-1:0] irline3_i21;
  wire signed [`W-1:0] irline3_i22;
  wire signed [`W-1:0] irline3_i23;
  wire signed [`W-1:0] irline3_i24;
  wire signed [`W-1:0] irline3_i25;
  wire signed [`W-1:0] irline3_i26;
  wire signed [`W-1:0] irline3_i27;
  wire signed [`W-1:0] irline3_i28;
  wire signed [`W-1:0] irline3_i29;
  wire signed [`W-1:0] irline3_i30;
  wire signed [`W-1:0] irline3_i31;
  wire signed [`W-1:0] irline3_i32;
  wire signed [`W-1:0] irline3_i33;
  wire signed [`W-1:0] irline3_i34;
  wire signed [`W-1:0] irline3_i35;
  wire signed [`W-1:0] irline3_i36;
  wire signed [`W-1:0] irline3_i37;
  wire signed [`W-1:0] irline3_i38;
  wire signed [`W-1:0] irline3_i39;
  wire signed [`W-1:0] irline3_i40;
  wire signed [`W-1:0] irline3_i41;
  wire signed [`W-1:0] irline3_i42;
  wire signed [`W-1:0] irline3_i43;
  wire signed [`W-1:0] irline3_i44;
  wire signed [`W-1:0] irline3_i45;
  wire signed [`W-1:0] irline3_i46;
  wire signed [`W-1:0] irline3_i47;
  wire signed [`W-1:0] irline3_i48;
  wire signed [`W-1:0] irline3_i49;
  wire signed [`W-1:0] irline3_i50;
  wire signed [`W-1:0] irline3_i51;
  wire signed [`W-1:0] irline3_i52;
  wire signed [`W-1:0] irline3_i53;
  wire signed [`W-1:0] irline3_i54;
  wire signed [`W-1:0] irline3_i55;
  wire signed [`W-1:0] irline3_i56;
  wire signed [`W-1:0] irline3_i57;
  wire signed [`W-1:0] irline3_i58;
  wire signed [`W-1:0] irline3_i59;
  wire signed [`W-1:0] irline3_i60;
  wire signed [`W-1:0] irline3_i61;
  wire signed [`W-1:0] irline3_i62;
  wire signed [`W-1:0] irline3_i63;
  wire signed [`W-1:0] irline3_i64;
  wire signed [`W-1:0] irline3_v;
  wire signed [`W-1:0] idb1_i0;
  wire signed [`W-1:0] idb1_i1;
  wire signed [`W-1:0] idb1_i2;
  wire signed [`W-1:0] idb1_i3;
  wire signed [`W-1:0] idb1_i4;
  wire signed [`W-1:0] idb1_i5;
  wire signed [`W-1:0] idb1_i6;
  wire signed [`W-1:0] idb1_i7;
  wire signed [`W-1:0] idb1_i8;
  wire signed [`W-1:0] idb1_i9;
  wire signed [`W-1:0] idb1_i10;
  wire signed [`W-1:0] idb1_i11;
  wire signed [`W-1:0] idb1_v;
  wire signed [`W-1:0] n990_i0;
  wire signed [`W-1:0] n990_i1;
  wire signed [`W-1:0] n990_i2;
  wire signed [`W-1:0] n990_i3;
  wire signed [`W-1:0] n990_v;
  wire signed [`W-1:0] n993_i0;
  wire signed [`W-1:0] n993_i1;
  wire signed [`W-1:0] n993_v;
  wire signed [`W-1:0] n992_i0;
  wire signed [`W-1:0] n992_i1;
  wire signed [`W-1:0] n992_i2;
  wire signed [`W-1:0] n992_v;
  wire signed [`W-1:0] n999_i0;
  wire signed [`W-1:0] n999_i1;
  wire signed [`W-1:0] n999_i2;
  wire signed [`W-1:0] n999_i3;
  wire signed [`W-1:0] n999_v;
  wire signed [`W-1:0] n998_i0;
  wire signed [`W-1:0] n998_i1;
  wire signed [`W-1:0] n998_i2;
  wire signed [`W-1:0] n998_i3;
  wire signed [`W-1:0] n998_i4;
  wire signed [`W-1:0] n998_v;
  wire signed [`W-1:0] op_T3_i0;
  wire signed [`W-1:0] op_T3_i1;
  wire signed [`W-1:0] op_T3_i2;
  wire signed [`W-1:0] op_T3_v;
  wire signed [`W-1:0] adl6_i0;
  wire signed [`W-1:0] adl6_i1;
  wire signed [`W-1:0] adl6_i2;
  wire signed [`W-1:0] adl6_i3;
  wire signed [`W-1:0] adl6_i4;
  wire signed [`W-1:0] adl6_i5;
  wire signed [`W-1:0] adl6_i6;
  wire signed [`W-1:0] adl6_i7;
  wire signed [`W-1:0] adl6_v;
  wire signed [`W-1:0] n122_i0;
  wire signed [`W-1:0] n122_i1;
  wire signed [`W-1:0] n122_i2;
  wire signed [`W-1:0] n122_v;
  wire signed [`W-1:0] n123_i0;
  wire signed [`W-1:0] n123_i1;
  wire signed [`W-1:0] n123_i2;
  wire signed [`W-1:0] n123_v;
  wire signed [`W-1:0] pchp3_i0;
  wire signed [`W-1:0] pchp3_i1;
  wire signed [`W-1:0] pchp3_i2;
  wire signed [`W-1:0] pchp3_v;
  wire signed [`W-1:0] PD_n_0xx0xx0x_i0;
  wire signed [`W-1:0] PD_n_0xx0xx0x_i1;
  wire signed [`W-1:0] PD_n_0xx0xx0x_i2;
  wire signed [`W-1:0] PD_n_0xx0xx0x_v;
  wire signed [`W-1:0] n126_i0;
  wire signed [`W-1:0] n126_i1;
  wire signed [`W-1:0] n126_v;
  wire signed [`W-1:0] n127_i0;
  wire signed [`W-1:0] n127_i1;
  wire signed [`W-1:0] n127_i2;
  wire signed [`W-1:0] n127_i3;
  wire signed [`W-1:0] n127_v;
  wire signed [`W-1:0] n128_i0;
  wire signed [`W-1:0] n128_i1;
  wire signed [`W-1:0] n128_i2;
  wire signed [`W-1:0] n128_v;
  wire signed [`W-1:0] dpc20_ADDSB06_i0;
  wire signed [`W-1:0] dpc20_ADDSB06_i1;
  wire signed [`W-1:0] dpc20_ADDSB06_i2;
  wire signed [`W-1:0] dpc20_ADDSB06_i3;
  wire signed [`W-1:0] dpc20_ADDSB06_i4;
  wire signed [`W-1:0] dpc20_ADDSB06_i5;
  wire signed [`W-1:0] dpc20_ADDSB06_i6;
  wire signed [`W-1:0] dpc20_ADDSB06_i7;
  wire signed [`W-1:0] dpc20_ADDSB06_i8;
  wire signed [`W-1:0] dpc20_ADDSB06_v;
  wire signed [`W-1:0] alub4_i0;
  wire signed [`W-1:0] alub4_i1;
  wire signed [`W-1:0] alub4_i2;
  wire signed [`W-1:0] alub4_i3;
  wire signed [`W-1:0] alub4_i4;
  wire signed [`W-1:0] alub4_v;
  wire signed [`W-1:0] n1647_i0;
  wire signed [`W-1:0] n1647_i1;
  wire signed [`W-1:0] n1647_i2;
  wire signed [`W-1:0] n1647_i3;
  wire signed [`W-1:0] n1647_i4;
  wire signed [`W-1:0] n1647_v;
  wire signed [`W-1:0] op_T__bit_i0;
  wire signed [`W-1:0] op_T__bit_i1;
  wire signed [`W-1:0] op_T__bit_i2;
  wire signed [`W-1:0] op_T__bit_i3;
  wire signed [`W-1:0] op_T__bit_v;
  wire signed [`W-1:0] n1641_i0;
  wire signed [`W-1:0] n1641_i1;
  wire signed [`W-1:0] n1641_i2;
  wire signed [`W-1:0] n1641_v;
  wire signed [`W-1:0] n1640_i0;
  wire signed [`W-1:0] n1640_i1;
  wire signed [`W-1:0] n1640_i2;
  wire signed [`W-1:0] n1640_v;
  wire signed [`W-1:0] n1643_i0;
  wire signed [`W-1:0] n1643_i1;
  wire signed [`W-1:0] n1643_i2;
  wire signed [`W-1:0] n1643_i3;
  wire signed [`W-1:0] n1643_i4;
  wire signed [`W-1:0] n1643_v;
  wire signed [`W-1:0] n1642_i0;
  wire signed [`W-1:0] n1642_i1;
  wire signed [`W-1:0] n1642_i2;
  wire signed [`W-1:0] n1642_v;
  wire signed [`W-1:0] n1649_i0;
  wire signed [`W-1:0] n1649_i1;
  wire signed [`W-1:0] n1649_i2;
  wire signed [`W-1:0] n1649_i3;
  wire signed [`W-1:0] n1649_v;
  wire signed [`W-1:0] x3_i0;
  wire signed [`W-1:0] x3_i1;
  wire signed [`W-1:0] x3_i2;
  wire signed [`W-1:0] x3_v;
  wire signed [`W-1:0] n1252_i0;
  wire signed [`W-1:0] n1252_i1;
  wire signed [`W-1:0] n1252_v;
  wire signed [`W-1:0] op_T3_jsr_i0;
  wire signed [`W-1:0] op_T3_jsr_i1;
  wire signed [`W-1:0] op_T3_jsr_i2;
  wire signed [`W-1:0] op_T3_jsr_v;
  wire signed [`W-1:0] n578_i0;
  wire signed [`W-1:0] n578_i1;
  wire signed [`W-1:0] n578_i2;
  wire signed [`W-1:0] n578_i3;
  wire signed [`W-1:0] n578_v;
  wire signed [`W-1:0] n604_i0;
  wire signed [`W-1:0] n604_i1;
  wire signed [`W-1:0] n604_i2;
  wire signed [`W-1:0] n604_i3;
  wire signed [`W-1:0] n604_i4;
  wire signed [`W-1:0] n604_v;
  wire signed [`W-1:0] y2_i0;
  wire signed [`W-1:0] y2_i1;
  wire signed [`W-1:0] y2_i2;
  wire signed [`W-1:0] y2_v;
  wire signed [`W-1:0] n572_i0;
  wire signed [`W-1:0] n572_i1;
  wire signed [`W-1:0] n572_i2;
  wire signed [`W-1:0] n572_i3;
  wire signed [`W-1:0] n572_v;
  wire signed [`W-1:0] n571_i0;
  wire signed [`W-1:0] n571_i1;
  wire signed [`W-1:0] n571_i2;
  wire signed [`W-1:0] n571_v;
  wire signed [`W-1:0] n570_i0;
  wire signed [`W-1:0] n570_i1;
  wire signed [`W-1:0] n570_i2;
  wire signed [`W-1:0] n570_v;
  wire signed [`W-1:0] notidl1_i0;
  wire signed [`W-1:0] notidl1_i1;
  wire signed [`W-1:0] notidl1_v;
  wire signed [`W-1:0] op_T0_adc_sbc_i0;
  wire signed [`W-1:0] op_T0_adc_sbc_i1;
  wire signed [`W-1:0] op_T0_adc_sbc_i2;
  wire signed [`W-1:0] op_T0_adc_sbc_i3;
  wire signed [`W-1:0] op_T0_adc_sbc_v;
  wire signed [`W-1:0] dpc15_ANDS_i0;
  wire signed [`W-1:0] dpc15_ANDS_i1;
  wire signed [`W-1:0] dpc15_ANDS_i2;
  wire signed [`W-1:0] dpc15_ANDS_i3;
  wire signed [`W-1:0] dpc15_ANDS_i4;
  wire signed [`W-1:0] dpc15_ANDS_i5;
  wire signed [`W-1:0] dpc15_ANDS_i6;
  wire signed [`W-1:0] dpc15_ANDS_i7;
  wire signed [`W-1:0] dpc15_ANDS_i8;
  wire signed [`W-1:0] dpc15_ANDS_i9;
  wire signed [`W-1:0] dpc15_ANDS_v;
  wire signed [`W-1:0] n1209_i0;
  wire signed [`W-1:0] n1209_i1;
  wire signed [`W-1:0] n1209_i2;
  wire signed [`W-1:0] n1209_v;
  wire signed [`W-1:0] Pout2_i0;
  wire signed [`W-1:0] Pout2_i1;
  wire signed [`W-1:0] Pout2_i2;
  wire signed [`W-1:0] Pout2_v;
  wire signed [`W-1:0] op_T0_lda_i0;
  wire signed [`W-1:0] op_T0_lda_i1;
  wire signed [`W-1:0] op_T0_lda_i2;
  wire signed [`W-1:0] op_T0_lda_i3;
  wire signed [`W-1:0] op_T0_lda_v;
  wire signed [`W-1:0] n1423_i0;
  wire signed [`W-1:0] n1423_i1;
  wire signed [`W-1:0] n1423_i2;
  wire signed [`W-1:0] n1423_i3;
  wire signed [`W-1:0] n1423_v;
  wire signed [`W-1:0] _C34_i0;
  wire signed [`W-1:0] _C34_i1;
  wire signed [`W-1:0] _C34_i2;
  wire signed [`W-1:0] _C34_i3;
  wire signed [`W-1:0] _C34_v;
  wire signed [`W-1:0] n1424_i0;
  wire signed [`W-1:0] n1424_i1;
  wire signed [`W-1:0] n1424_i2;
  wire signed [`W-1:0] n1424_i3;
  wire signed [`W-1:0] n1424_v;
  wire signed [`W-1:0] n1427_i0;
  wire signed [`W-1:0] n1427_i1;
  wire signed [`W-1:0] n1427_i2;
  wire signed [`W-1:0] n1427_v;
  wire signed [`W-1:0] abh0_i0;
  wire signed [`W-1:0] abh0_i1;
  wire signed [`W-1:0] abh0_i2;
  wire signed [`W-1:0] abh0_i3;
  wire signed [`W-1:0] abh0_i4;
  wire signed [`W-1:0] abh0_v;
  wire signed [`W-1:0] op_T3_ind_x_i0;
  wire signed [`W-1:0] op_T3_ind_x_i1;
  wire signed [`W-1:0] op_T3_ind_x_i2;
  wire signed [`W-1:0] op_T3_ind_x_i3;
  wire signed [`W-1:0] op_T3_ind_x_v;
  wire signed [`W-1:0] n602_i0;
  wire signed [`W-1:0] n602_i1;
  wire signed [`W-1:0] n602_i2;
  wire signed [`W-1:0] n602_v;
  wire signed [`W-1:0] pclp6_i0;
  wire signed [`W-1:0] pclp6_i1;
  wire signed [`W-1:0] pclp6_i2;
  wire signed [`W-1:0] pclp6_v;
  wire signed [`W-1:0] n730_i0;
  wire signed [`W-1:0] n730_i1;
  wire signed [`W-1:0] n730_i2;
  wire signed [`W-1:0] n730_v;
  wire signed [`W-1:0] n733_i0;
  wire signed [`W-1:0] n733_i1;
  wire signed [`W-1:0] n733_i2;
  wire signed [`W-1:0] n733_i3;
  wire signed [`W-1:0] n733_v;
  wire signed [`W-1:0] n732_i0;
  wire signed [`W-1:0] n732_i1;
  wire signed [`W-1:0] n732_i2;
  wire signed [`W-1:0] n732_i3;
  wire signed [`W-1:0] n732_v;
  wire signed [`W-1:0] n735_i0;
  wire signed [`W-1:0] n735_i1;
  wire signed [`W-1:0] n735_i2;
  wire signed [`W-1:0] n735_v;
  wire signed [`W-1:0] a0_i0;
  wire signed [`W-1:0] a0_i1;
  wire signed [`W-1:0] a0_i2;
  wire signed [`W-1:0] a0_v;
  wire signed [`W-1:0] ab5_i0;
  wire signed [`W-1:0] ab5_i1;
  wire signed [`W-1:0] ab5_i2;
  wire signed [`W-1:0] ab5_v;
  wire signed [`W-1:0] n739_i0;
  wire signed [`W-1:0] n739_i1;
  wire signed [`W-1:0] n739_i2;
  wire signed [`W-1:0] n739_i3;
  wire signed [`W-1:0] n739_v;
  wire signed [`W-1:0] pcl3_i0;
  wire signed [`W-1:0] pcl3_i1;
  wire signed [`W-1:0] pcl3_i2;
  wire signed [`W-1:0] pcl3_v;
  wire signed [`W-1:0] n1358_i0;
  wire signed [`W-1:0] n1358_i1;
  wire signed [`W-1:0] n1358_i2;
  wire signed [`W-1:0] n1358_i3;
  wire signed [`W-1:0] n1358_v;
  wire signed [`W-1:0] n469_i0;
  wire signed [`W-1:0] n469_i1;
  wire signed [`W-1:0] n469_v;
  wire signed [`W-1:0] n468_i0;
  wire signed [`W-1:0] n468_i1;
  wire signed [`W-1:0] n468_i2;
  wire signed [`W-1:0] n468_v;
  wire signed [`W-1:0] _WR_i0;
  wire signed [`W-1:0] _WR_i1;
  wire signed [`W-1:0] _WR_i2;
  wire signed [`W-1:0] _WR_v;
  wire signed [`W-1:0] n467_i0;
  wire signed [`W-1:0] n467_i1;
  wire signed [`W-1:0] n467_i2;
  wire signed [`W-1:0] n467_i3;
  wire signed [`W-1:0] n467_v;
  wire signed [`W-1:0] n466_i0;
  wire signed [`W-1:0] n466_i1;
  wire signed [`W-1:0] n466_i2;
  wire signed [`W-1:0] n466_i3;
  wire signed [`W-1:0] n466_v;
  wire signed [`W-1:0] n1357_i0;
  wire signed [`W-1:0] n1357_i1;
  wire signed [`W-1:0] n1357_i2;
  wire signed [`W-1:0] n1357_i3;
  wire signed [`W-1:0] n1357_i4;
  wire signed [`W-1:0] n1357_i5;
  wire signed [`W-1:0] n1357_v;
  wire signed [`W-1:0] n1356_i0;
  wire signed [`W-1:0] n1356_i1;
  wire signed [`W-1:0] n1356_i2;
  wire signed [`W-1:0] n1356_v;
  wire signed [`W-1:0] op_T0_cmp_i0;
  wire signed [`W-1:0] op_T0_cmp_i1;
  wire signed [`W-1:0] op_T0_cmp_i2;
  wire signed [`W-1:0] op_T0_cmp_v;
  wire signed [`W-1:0] n462_i0;
  wire signed [`W-1:0] n462_i1;
  wire signed [`W-1:0] n462_i2;
  wire signed [`W-1:0] n462_i3;
  wire signed [`W-1:0] n462_v;
  wire signed [`W-1:0] n1519_i0;
  wire signed [`W-1:0] n1519_i1;
  wire signed [`W-1:0] n1519_i2;
  wire signed [`W-1:0] n1519_v;
  wire signed [`W-1:0] n1518_i0;
  wire signed [`W-1:0] n1518_i1;
  wire signed [`W-1:0] n1518_i2;
  wire signed [`W-1:0] n1518_v;
  wire signed [`W-1:0] n1517_i0;
  wire signed [`W-1:0] n1517_i1;
  wire signed [`W-1:0] n1517_i2;
  wire signed [`W-1:0] n1517_v;
  wire signed [`W-1:0] notidl4_i0;
  wire signed [`W-1:0] notidl4_i1;
  wire signed [`W-1:0] notidl4_v;
  wire signed [`W-1:0] n1511_i0;
  wire signed [`W-1:0] n1511_i1;
  wire signed [`W-1:0] n1511_i2;
  wire signed [`W-1:0] n1511_v;
  wire signed [`W-1:0] _ABL5_i0;
  wire signed [`W-1:0] _ABL5_i1;
  wire signed [`W-1:0] _ABL5_i2;
  wire signed [`W-1:0] _ABL5_v;
  wire signed [`W-1:0] op_T2_abs_y_i0;
  wire signed [`W-1:0] op_T2_abs_y_i1;
  wire signed [`W-1:0] op_T2_abs_y_i2;
  wire signed [`W-1:0] op_T2_abs_y_v;
  wire signed [`W-1:0] pipeVectorA0_i0;
  wire signed [`W-1:0] pipeVectorA0_i1;
  wire signed [`W-1:0] pipeVectorA0_v;
  wire signed [`W-1:0] n355_i0;
  wire signed [`W-1:0] n355_i1;
  wire signed [`W-1:0] n355_i2;
  wire signed [`W-1:0] n355_i3;
  wire signed [`W-1:0] n355_v;
  wire signed [`W-1:0] op_T4_abs_idx_i0;
  wire signed [`W-1:0] op_T4_abs_idx_i1;
  wire signed [`W-1:0] op_T4_abs_idx_i2;
  wire signed [`W-1:0] op_T4_abs_idx_v;
  wire signed [`W-1:0] RnWstretched_i0;
  wire signed [`W-1:0] RnWstretched_i1;
  wire signed [`W-1:0] RnWstretched_i2;
  wire signed [`W-1:0] RnWstretched_i3;
  wire signed [`W-1:0] RnWstretched_i4;
  wire signed [`W-1:0] RnWstretched_i5;
  wire signed [`W-1:0] RnWstretched_i6;
  wire signed [`W-1:0] RnWstretched_i7;
  wire signed [`W-1:0] RnWstretched_i8;
  wire signed [`W-1:0] RnWstretched_i9;
  wire signed [`W-1:0] RnWstretched_i10;
  wire signed [`W-1:0] RnWstretched_i11;
  wire signed [`W-1:0] RnWstretched_i12;
  wire signed [`W-1:0] RnWstretched_i13;
  wire signed [`W-1:0] RnWstretched_i14;
  wire signed [`W-1:0] RnWstretched_i15;
  wire signed [`W-1:0] RnWstretched_i16;
  wire signed [`W-1:0] RnWstretched_i17;
  wire signed [`W-1:0] RnWstretched_i18;
  wire signed [`W-1:0] RnWstretched_i19;
  wire signed [`W-1:0] RnWstretched_i20;
  wire signed [`W-1:0] RnWstretched_i21;
  wire signed [`W-1:0] RnWstretched_i22;
  wire signed [`W-1:0] RnWstretched_i23;
  wire signed [`W-1:0] RnWstretched_i24;
  wire signed [`W-1:0] RnWstretched_i25;
  wire signed [`W-1:0] RnWstretched_v;
  wire signed [`W-1:0] op_T4_brk_i0;
  wire signed [`W-1:0] op_T4_brk_i1;
  wire signed [`W-1:0] op_T4_brk_i2;
  wire signed [`W-1:0] op_T4_brk_i3;
  wire signed [`W-1:0] op_T4_brk_v;
  wire signed [`W-1:0] n351_i0;
  wire signed [`W-1:0] n351_i1;
  wire signed [`W-1:0] n351_i2;
  wire signed [`W-1:0] n351_v;
  wire signed [`W-1:0] n350_i0;
  wire signed [`W-1:0] n350_i1;
  wire signed [`W-1:0] n350_i2;
  wire signed [`W-1:0] n350_i3;
  wire signed [`W-1:0] n350_i4;
  wire signed [`W-1:0] n350_v;
  wire signed [`W-1:0] n359_i0;
  wire signed [`W-1:0] n359_i1;
  wire signed [`W-1:0] n359_i2;
  wire signed [`W-1:0] n359_i3;
  wire signed [`W-1:0] n359_v;
  wire signed [`W-1:0] n358_i0;
  wire signed [`W-1:0] n358_i1;
  wire signed [`W-1:0] n358_i2;
  wire signed [`W-1:0] n358_i3;
  wire signed [`W-1:0] n358_i4;
  wire signed [`W-1:0] n358_v;
  wire signed [`W-1:0] n1111_i0;
  wire signed [`W-1:0] n1111_i1;
  wire signed [`W-1:0] n1111_i2;
  wire signed [`W-1:0] n1111_i3;
  wire signed [`W-1:0] n1111_v;
  wire signed [`W-1:0] n1110_i0;
  wire signed [`W-1:0] n1110_i1;
  wire signed [`W-1:0] n1110_i2;
  wire signed [`W-1:0] n1110_i3;
  wire signed [`W-1:0] n1110_v;
  wire signed [`W-1:0] n1113_i0;
  wire signed [`W-1:0] n1113_i1;
  wire signed [`W-1:0] n1113_v;
  wire signed [`W-1:0] _ABH6_i0;
  wire signed [`W-1:0] _ABH6_i1;
  wire signed [`W-1:0] _ABH6_i2;
  wire signed [`W-1:0] _ABH6_v;
  wire signed [`W-1:0] n288_i0;
  wire signed [`W-1:0] n288_i1;
  wire signed [`W-1:0] n288_i2;
  wire signed [`W-1:0] n288_i3;
  wire signed [`W-1:0] n288_v;
  wire signed [`W-1:0] Pout1_i0;
  wire signed [`W-1:0] Pout1_i1;
  wire signed [`W-1:0] Pout1_i2;
  wire signed [`W-1:0] Pout1_v;
  wire signed [`W-1:0] op_T4_mem_abs_idx_i0;
  wire signed [`W-1:0] op_T4_mem_abs_idx_i1;
  wire signed [`W-1:0] op_T4_mem_abs_idx_i2;
  wire signed [`W-1:0] op_T4_mem_abs_idx_v;
  wire signed [`W-1:0] n280_i0;
  wire signed [`W-1:0] n280_i1;
  wire signed [`W-1:0] n280_i2;
  wire signed [`W-1:0] n280_i3;
  wire signed [`W-1:0] n280_i4;
  wire signed [`W-1:0] n280_v;
  wire signed [`W-1:0] dpc37_PCLDB_i0;
  wire signed [`W-1:0] dpc37_PCLDB_i1;
  wire signed [`W-1:0] dpc37_PCLDB_i2;
  wire signed [`W-1:0] dpc37_PCLDB_i3;
  wire signed [`W-1:0] dpc37_PCLDB_i4;
  wire signed [`W-1:0] dpc37_PCLDB_i5;
  wire signed [`W-1:0] dpc37_PCLDB_i6;
  wire signed [`W-1:0] dpc37_PCLDB_i7;
  wire signed [`W-1:0] dpc37_PCLDB_i8;
  wire signed [`W-1:0] dpc37_PCLDB_i9;
  wire signed [`W-1:0] dpc37_PCLDB_v;
  wire signed [`W-1:0] n282_i0;
  wire signed [`W-1:0] n282_i1;
  wire signed [`W-1:0] n282_i2;
  wire signed [`W-1:0] n282_v;
  wire signed [`W-1:0] op_T2_zp_zp_idx_i0;
  wire signed [`W-1:0] op_T2_zp_zp_idx_i1;
  wire signed [`W-1:0] op_T2_zp_zp_idx_i2;
  wire signed [`W-1:0] op_T2_zp_zp_idx_v;
  wire signed [`W-1:0] n284_i0;
  wire signed [`W-1:0] n284_i1;
  wire signed [`W-1:0] n284_i2;
  wire signed [`W-1:0] n284_v;
  wire signed [`W-1:0] abh2_i0;
  wire signed [`W-1:0] abh2_i1;
  wire signed [`W-1:0] abh2_i2;
  wire signed [`W-1:0] abh2_i3;
  wire signed [`W-1:0] abh2_i4;
  wire signed [`W-1:0] abh2_v;
  wire signed [`W-1:0] op_T0_tay_ldy_not_idx_i0;
  wire signed [`W-1:0] op_T0_tay_ldy_not_idx_i1;
  wire signed [`W-1:0] op_T0_tay_ldy_not_idx_i2;
  wire signed [`W-1:0] op_T0_tay_ldy_not_idx_v;
  wire signed [`W-1:0] n1441_i0;
  wire signed [`W-1:0] n1441_i1;
  wire signed [`W-1:0] n1441_i2;
  wire signed [`W-1:0] n1441_v;
  wire signed [`W-1:0] n1440_i0;
  wire signed [`W-1:0] n1440_i1;
  wire signed [`W-1:0] n1440_i2;
  wire signed [`W-1:0] n1440_v;
  wire signed [`W-1:0] dasb5_i0;
  wire signed [`W-1:0] dasb5_i1;
  wire signed [`W-1:0] dasb5_i2;
  wire signed [`W-1:0] dasb5_v;
  wire signed [`W-1:0] n262_i0;
  wire signed [`W-1:0] n262_i1;
  wire signed [`W-1:0] n262_i2;
  wire signed [`W-1:0] n262_v;
  wire signed [`W-1:0] n261_i0;
  wire signed [`W-1:0] n261_i1;
  wire signed [`W-1:0] n261_i2;
  wire signed [`W-1:0] n261_v;
  wire signed [`W-1:0] n260_i0;
  wire signed [`W-1:0] n260_i1;
  wire signed [`W-1:0] n260_i2;
  wire signed [`W-1:0] n260_v;
  wire signed [`W-1:0] n267_i0;
  wire signed [`W-1:0] n267_i1;
  wire signed [`W-1:0] n267_i2;
  wire signed [`W-1:0] n267_v;
  wire signed [`W-1:0] n266_i0;
  wire signed [`W-1:0] n266_i1;
  wire signed [`W-1:0] n266_v;
  wire signed [`W-1:0] n265_i0;
  wire signed [`W-1:0] n265_i1;
  wire signed [`W-1:0] n265_v;
  wire signed [`W-1:0] n264_i0;
  wire signed [`W-1:0] n264_i1;
  wire signed [`W-1:0] n264_i2;
  wire signed [`W-1:0] n264_i3;
  wire signed [`W-1:0] n264_i4;
  wire signed [`W-1:0] n264_i5;
  wire signed [`W-1:0] n264_v;
  wire signed [`W-1:0] n269_i0;
  wire signed [`W-1:0] n269_i1;
  wire signed [`W-1:0] n269_i2;
  wire signed [`W-1:0] n269_v;
  wire signed [`W-1:0] ab0_i0;
  wire signed [`W-1:0] ab0_i1;
  wire signed [`W-1:0] ab0_i2;
  wire signed [`W-1:0] ab0_v;
  wire signed [`W-1:0] op_xy_i0;
  wire signed [`W-1:0] op_xy_i1;
  wire signed [`W-1:0] op_xy_i2;
  wire signed [`W-1:0] op_xy_i3;
  wire signed [`W-1:0] op_xy_v;
  wire signed [`W-1:0] n1291_i0;
  wire signed [`W-1:0] n1291_i1;
  wire signed [`W-1:0] n1291_v;
  wire signed [`W-1:0] n1296_i0;
  wire signed [`W-1:0] n1296_i1;
  wire signed [`W-1:0] n1296_i2;
  wire signed [`W-1:0] n1296_v;
  wire signed [`W-1:0] n1565_i0;
  wire signed [`W-1:0] n1565_i1;
  wire signed [`W-1:0] n1565_v;
  wire signed [`W-1:0] PD_1xx000x0_i0;
  wire signed [`W-1:0] PD_1xx000x0_i1;
  wire signed [`W-1:0] PD_1xx000x0_i2;
  wire signed [`W-1:0] PD_1xx000x0_v;
  wire signed [`W-1:0] n1295_i0;
  wire signed [`W-1:0] n1295_i1;
  wire signed [`W-1:0] n1295_i2;
  wire signed [`W-1:0] n1295_i3;
  wire signed [`W-1:0] n1295_v;
  wire signed [`W-1:0] n988_i0;
  wire signed [`W-1:0] n988_i1;
  wire signed [`W-1:0] n988_i2;
  wire signed [`W-1:0] n988_i3;
  wire signed [`W-1:0] n988_v;
  wire signed [`W-1:0] y4_i0;
  wire signed [`W-1:0] y4_i1;
  wire signed [`W-1:0] y4_i2;
  wire signed [`W-1:0] y4_v;
  wire signed [`W-1:0] n982_i0;
  wire signed [`W-1:0] n982_i1;
  wire signed [`W-1:0] n982_v;
  wire signed [`W-1:0] n983_i0;
  wire signed [`W-1:0] n983_i1;
  wire signed [`W-1:0] n983_i2;
  wire signed [`W-1:0] n983_v;
  wire signed [`W-1:0] n980_i0;
  wire signed [`W-1:0] n980_i1;
  wire signed [`W-1:0] n980_i2;
  wire signed [`W-1:0] n980_v;
  wire signed [`W-1:0] n981_i0;
  wire signed [`W-1:0] n981_i1;
  wire signed [`W-1:0] n981_i2;
  wire signed [`W-1:0] n981_v;
  wire signed [`W-1:0] n986_i0;
  wire signed [`W-1:0] n986_i1;
  wire signed [`W-1:0] n986_i2;
  wire signed [`W-1:0] n986_v;
  wire signed [`W-1:0] n987_i0;
  wire signed [`W-1:0] n987_i1;
  wire signed [`W-1:0] n987_i2;
  wire signed [`W-1:0] n987_v;
  wire signed [`W-1:0] dpc12_0ADD_i0;
  wire signed [`W-1:0] dpc12_0ADD_i1;
  wire signed [`W-1:0] dpc12_0ADD_i2;
  wire signed [`W-1:0] dpc12_0ADD_i3;
  wire signed [`W-1:0] dpc12_0ADD_i4;
  wire signed [`W-1:0] dpc12_0ADD_i5;
  wire signed [`W-1:0] dpc12_0ADD_i6;
  wire signed [`W-1:0] dpc12_0ADD_i7;
  wire signed [`W-1:0] dpc12_0ADD_i8;
  wire signed [`W-1:0] dpc12_0ADD_i9;
  wire signed [`W-1:0] dpc12_0ADD_v;
  wire signed [`W-1:0] op_T0_ldx_tax_tsx_i0;
  wire signed [`W-1:0] op_T0_ldx_tax_tsx_i1;
  wire signed [`W-1:0] op_T0_ldx_tax_tsx_i2;
  wire signed [`W-1:0] op_T0_ldx_tax_tsx_v;
  wire signed [`W-1:0] y6_i0;
  wire signed [`W-1:0] y6_i1;
  wire signed [`W-1:0] y6_i2;
  wire signed [`W-1:0] y6_v;
  wire signed [`W-1:0] pchp2_i0;
  wire signed [`W-1:0] pchp2_i1;
  wire signed [`W-1:0] pchp2_v;
  wire signed [`W-1:0] A_B7_i0;
  wire signed [`W-1:0] A_B7_i1;
  wire signed [`W-1:0] A_B7_i2;
  wire signed [`W-1:0] A_B7_v;
  wire signed [`W-1:0] notidl0_i0;
  wire signed [`W-1:0] notidl0_i1;
  wire signed [`W-1:0] notidl0_v;
  wire signed [`W-1:0] n111_i0;
  wire signed [`W-1:0] n111_i1;
  wire signed [`W-1:0] n111_i2;
  wire signed [`W-1:0] n111_v;
  wire signed [`W-1:0] n110_i0;
  wire signed [`W-1:0] n110_i1;
  wire signed [`W-1:0] n110_i2;
  wire signed [`W-1:0] n110_v;
  wire signed [`W-1:0] pchp1_i0;
  wire signed [`W-1:0] pchp1_i1;
  wire signed [`W-1:0] pchp1_i2;
  wire signed [`W-1:0] pchp1_v;
  wire signed [`W-1:0] n119_i0;
  wire signed [`W-1:0] n119_i1;
  wire signed [`W-1:0] n119_i2;
  wire signed [`W-1:0] n119_v;
  wire signed [`W-1:0] n118_i0;
  wire signed [`W-1:0] n118_i1;
  wire signed [`W-1:0] n118_i2;
  wire signed [`W-1:0] n118_v;
  wire signed [`W-1:0] _DBE_i0;
  wire signed [`W-1:0] _DBE_i1;
  wire signed [`W-1:0] _DBE_i2;
  wire signed [`W-1:0] _DBE_v;
  wire signed [`W-1:0] adl5_i0;
  wire signed [`W-1:0] adl5_i1;
  wire signed [`W-1:0] adl5_i2;
  wire signed [`W-1:0] adl5_i3;
  wire signed [`W-1:0] adl5_i4;
  wire signed [`W-1:0] adl5_i5;
  wire signed [`W-1:0] adl5_i6;
  wire signed [`W-1:0] adl5_i7;
  wire signed [`W-1:0] adl5_v;
  wire signed [`W-1:0] n1631_i0;
  wire signed [`W-1:0] n1631_i1;
  wire signed [`W-1:0] n1631_i2;
  wire signed [`W-1:0] n1631_v;
  wire signed [`W-1:0] n1632_i0;
  wire signed [`W-1:0] n1632_i1;
  wire signed [`W-1:0] n1632_i2;
  wire signed [`W-1:0] n1632_i3;
  wire signed [`W-1:0] n1632_i4;
  wire signed [`W-1:0] n1632_v;
  wire signed [`W-1:0] n1633_i0;
  wire signed [`W-1:0] n1633_i1;
  wire signed [`W-1:0] n1633_i2;
  wire signed [`W-1:0] n1633_v;
  wire signed [`W-1:0] dor2_i0;
  wire signed [`W-1:0] dor2_i1;
  wire signed [`W-1:0] dor2_i2;
  wire signed [`W-1:0] dor2_i3;
  wire signed [`W-1:0] dor2_i4;
  wire signed [`W-1:0] dor2_v;
  wire signed [`W-1:0] n1635_i0;
  wire signed [`W-1:0] n1635_i1;
  wire signed [`W-1:0] n1635_i2;
  wire signed [`W-1:0] n1635_v;
  wire signed [`W-1:0] alu2_i0;
  wire signed [`W-1:0] alu2_i1;
  wire signed [`W-1:0] alu2_i2;
  wire signed [`W-1:0] alu2_i3;
  wire signed [`W-1:0] alu2_i4;
  wire signed [`W-1:0] alu2_v;
  wire signed [`W-1:0] n1638_i0;
  wire signed [`W-1:0] n1638_i1;
  wire signed [`W-1:0] n1638_i2;
  wire signed [`W-1:0] n1638_v;
  wire signed [`W-1:0] n1639_i0;
  wire signed [`W-1:0] n1639_i1;
  wire signed [`W-1:0] n1639_i2;
  wire signed [`W-1:0] n1639_v;
  wire signed [`W-1:0] n568_i0;
  wire signed [`W-1:0] n568_i1;
  wire signed [`W-1:0] n568_i2;
  wire signed [`W-1:0] n568_v;
  wire signed [`W-1:0] C78_phi2_i0;
  wire signed [`W-1:0] C78_phi2_i1;
  wire signed [`W-1:0] C78_phi2_v;
  wire signed [`W-1:0] pipeUNK22_i0;
  wire signed [`W-1:0] pipeUNK22_i1;
  wire signed [`W-1:0] pipeUNK22_v;
  wire signed [`W-1:0] n562_i0;
  wire signed [`W-1:0] n562_i1;
  wire signed [`W-1:0] n562_v;
  wire signed [`W-1:0] n564_i0;
  wire signed [`W-1:0] n564_i1;
  wire signed [`W-1:0] n564_i2;
  wire signed [`W-1:0] n564_i3;
  wire signed [`W-1:0] n564_v;
  wire signed [`W-1:0] n565_i0;
  wire signed [`W-1:0] n565_i1;
  wire signed [`W-1:0] n565_i2;
  wire signed [`W-1:0] n565_v;
  wire signed [`W-1:0] n566_i0;
  wire signed [`W-1:0] n566_i1;
  wire signed [`W-1:0] n566_i2;
  wire signed [`W-1:0] n566_v;
  wire signed [`W-1:0] n567_i0;
  wire signed [`W-1:0] n567_i1;
  wire signed [`W-1:0] n567_i2;
  wire signed [`W-1:0] n567_i3;
  wire signed [`W-1:0] n567_i4;
  wire signed [`W-1:0] n567_v;
  wire signed [`W-1:0] sb3_i0;
  wire signed [`W-1:0] sb3_i1;
  wire signed [`W-1:0] sb3_i2;
  wire signed [`W-1:0] sb3_i3;
  wire signed [`W-1:0] sb3_i4;
  wire signed [`W-1:0] sb3_i5;
  wire signed [`W-1:0] sb3_i6;
  wire signed [`W-1:0] sb3_i7;
  wire signed [`W-1:0] sb3_i8;
  wire signed [`W-1:0] sb3_i9;
  wire signed [`W-1:0] sb3_i10;
  wire signed [`W-1:0] sb3_i11;
  wire signed [`W-1:0] sb3_i12;
  wire signed [`W-1:0] sb3_v;
  wire signed [`W-1:0] dpc3_SBX_i0;
  wire signed [`W-1:0] dpc3_SBX_i1;
  wire signed [`W-1:0] dpc3_SBX_i2;
  wire signed [`W-1:0] dpc3_SBX_i3;
  wire signed [`W-1:0] dpc3_SBX_i4;
  wire signed [`W-1:0] dpc3_SBX_i5;
  wire signed [`W-1:0] dpc3_SBX_i6;
  wire signed [`W-1:0] dpc3_SBX_i7;
  wire signed [`W-1:0] dpc3_SBX_i8;
  wire signed [`W-1:0] dpc3_SBX_i9;
  wire signed [`W-1:0] dpc3_SBX_v;
  wire signed [`W-1:0] n1187_i0;
  wire signed [`W-1:0] n1187_i1;
  wire signed [`W-1:0] n1187_i2;
  wire signed [`W-1:0] n1187_v;
  wire signed [`W-1:0] n1184_i0;
  wire signed [`W-1:0] n1184_i1;
  wire signed [`W-1:0] n1184_i2;
  wire signed [`W-1:0] n1184_i3;
  wire signed [`W-1:0] n1184_i4;
  wire signed [`W-1:0] n1184_v;
  wire signed [`W-1:0] short_circuit_idx_add_i0;
  wire signed [`W-1:0] short_circuit_idx_add_i1;
  wire signed [`W-1:0] short_circuit_idx_add_i2;
  wire signed [`W-1:0] short_circuit_idx_add_v;
  wire signed [`W-1:0] notir2_i0;
  wire signed [`W-1:0] notir2_i1;
  wire signed [`W-1:0] notir2_i2;
  wire signed [`W-1:0] notir2_i3;
  wire signed [`W-1:0] notir2_i4;
  wire signed [`W-1:0] notir2_i5;
  wire signed [`W-1:0] notir2_i6;
  wire signed [`W-1:0] notir2_i7;
  wire signed [`W-1:0] notir2_i8;
  wire signed [`W-1:0] notir2_i9;
  wire signed [`W-1:0] notir2_i10;
  wire signed [`W-1:0] notir2_i11;
  wire signed [`W-1:0] notir2_i12;
  wire signed [`W-1:0] notir2_i13;
  wire signed [`W-1:0] notir2_i14;
  wire signed [`W-1:0] notir2_i15;
  wire signed [`W-1:0] notir2_i16;
  wire signed [`W-1:0] notir2_i17;
  wire signed [`W-1:0] notir2_i18;
  wire signed [`W-1:0] notir2_i19;
  wire signed [`W-1:0] notir2_i20;
  wire signed [`W-1:0] notir2_v;
  wire signed [`W-1:0] n1180_i0;
  wire signed [`W-1:0] n1180_i1;
  wire signed [`W-1:0] n1180_i2;
  wire signed [`W-1:0] n1180_v;
  wire signed [`W-1:0] n1181_i0;
  wire signed [`W-1:0] n1181_i1;
  wire signed [`W-1:0] n1181_i2;
  wire signed [`W-1:0] n1181_v;
  wire signed [`W-1:0] n726_i0;
  wire signed [`W-1:0] n726_i1;
  wire signed [`W-1:0] n726_i2;
  wire signed [`W-1:0] n726_v;
  wire signed [`W-1:0] a4_i0;
  wire signed [`W-1:0] a4_i1;
  wire signed [`W-1:0] a4_i2;
  wire signed [`W-1:0] a4_v;
  wire signed [`W-1:0] dpc22__DSA_i0;
  wire signed [`W-1:0] dpc22__DSA_i1;
  wire signed [`W-1:0] dpc22__DSA_i2;
  wire signed [`W-1:0] dpc22__DSA_i3;
  wire signed [`W-1:0] dpc22__DSA_v;
  wire signed [`W-1:0] n722_i0;
  wire signed [`W-1:0] n722_i1;
  wire signed [`W-1:0] n722_i2;
  wire signed [`W-1:0] n722_i3;
  wire signed [`W-1:0] n722_i4;
  wire signed [`W-1:0] n722_i5;
  wire signed [`W-1:0] n722_v;
  wire signed [`W-1:0] n723_i0;
  wire signed [`W-1:0] n723_i1;
  wire signed [`W-1:0] n723_i2;
  wire signed [`W-1:0] n723_i3;
  wire signed [`W-1:0] n723_i4;
  wire signed [`W-1:0] n723_v;
  wire signed [`W-1:0] n720_i0;
  wire signed [`W-1:0] n720_i1;
  wire signed [`W-1:0] n720_i2;
  wire signed [`W-1:0] n720_v;
  wire signed [`W-1:0] n721_i0;
  wire signed [`W-1:0] n721_i1;
  wire signed [`W-1:0] n721_i2;
  wire signed [`W-1:0] n721_i3;
  wire signed [`W-1:0] n721_i4;
  wire signed [`W-1:0] n721_v;
  wire signed [`W-1:0] n728_i0;
  wire signed [`W-1:0] n728_i1;
  wire signed [`W-1:0] n728_i2;
  wire signed [`W-1:0] n728_v;
  wire signed [`W-1:0] pipeUNK36_i0;
  wire signed [`W-1:0] pipeUNK36_i1;
  wire signed [`W-1:0] pipeUNK36_v;
  wire signed [`W-1:0] op_clv_i0;
  wire signed [`W-1:0] op_clv_i1;
  wire signed [`W-1:0] op_clv_i2;
  wire signed [`W-1:0] op_clv_v;
  wire signed [`W-1:0] notalucin_i0;
  wire signed [`W-1:0] notalucin_i1;
  wire signed [`W-1:0] notalucin_i2;
  wire signed [`W-1:0] notalucin_i3;
  wire signed [`W-1:0] notalucin_i4;
  wire signed [`W-1:0] notalucin_v;
  wire signed [`W-1:0] n1166_i0;
  wire signed [`W-1:0] n1166_i1;
  wire signed [`W-1:0] n1166_i2;
  wire signed [`W-1:0] n1166_i3;
  wire signed [`W-1:0] n1166_v;
  wire signed [`W-1:0] alua0_i0;
  wire signed [`W-1:0] alua0_i1;
  wire signed [`W-1:0] alua0_i2;
  wire signed [`W-1:0] alua0_i3;
  wire signed [`W-1:0] alua0_v;
  wire signed [`W-1:0] adh4_i0;
  wire signed [`W-1:0] adh4_i1;
  wire signed [`W-1:0] adh4_i2;
  wire signed [`W-1:0] adh4_i3;
  wire signed [`W-1:0] adh4_i4;
  wire signed [`W-1:0] adh4_i5;
  wire signed [`W-1:0] adh4_i6;
  wire signed [`W-1:0] adh4_v;
  wire signed [`W-1:0] n1161_i0;
  wire signed [`W-1:0] n1161_i1;
  wire signed [`W-1:0] n1161_v;
  wire signed [`W-1:0] n1162_i0;
  wire signed [`W-1:0] n1162_i1;
  wire signed [`W-1:0] n1162_v;
  wire signed [`W-1:0] clk1out_i0;
  wire signed [`W-1:0] clk1out_i1;
  wire signed [`W-1:0] clk1out_i2;
  wire signed [`W-1:0] clk1out_v;
  wire signed [`W-1:0] op_T5_ind_y_i0;
  wire signed [`W-1:0] op_T5_ind_y_i1;
  wire signed [`W-1:0] op_T5_ind_y_i2;
  wire signed [`W-1:0] op_T5_ind_y_v;
  wire signed [`W-1:0] n1169_i0;
  wire signed [`W-1:0] n1169_i1;
  wire signed [`W-1:0] n1169_i2;
  wire signed [`W-1:0] n1169_i3;
  wire signed [`W-1:0] n1169_v;
  wire signed [`W-1:0] dpc30_ADHPCH_i0;
  wire signed [`W-1:0] dpc30_ADHPCH_i1;
  wire signed [`W-1:0] dpc30_ADHPCH_i2;
  wire signed [`W-1:0] dpc30_ADHPCH_i3;
  wire signed [`W-1:0] dpc30_ADHPCH_i4;
  wire signed [`W-1:0] dpc30_ADHPCH_i5;
  wire signed [`W-1:0] dpc30_ADHPCH_i6;
  wire signed [`W-1:0] dpc30_ADHPCH_i7;
  wire signed [`W-1:0] dpc30_ADHPCH_i8;
  wire signed [`W-1:0] dpc30_ADHPCH_i9;
  wire signed [`W-1:0] dpc30_ADHPCH_v;
  wire signed [`W-1:0] pch5_i0;
  wire signed [`W-1:0] pch5_i1;
  wire signed [`W-1:0] pch5_i2;
  wire signed [`W-1:0] pch5_v;
  wire signed [`W-1:0] n46_i0;
  wire signed [`W-1:0] n46_i1;
  wire signed [`W-1:0] n46_i2;
  wire signed [`W-1:0] n46_v;
  wire signed [`W-1:0] n47_i0;
  wire signed [`W-1:0] n47_i1;
  wire signed [`W-1:0] n47_v;
  wire signed [`W-1:0] pipeUNK05_i0;
  wire signed [`W-1:0] pipeUNK05_i1;
  wire signed [`W-1:0] pipeUNK05_v;
  wire signed [`W-1:0] pipeVectorA2_i0;
  wire signed [`W-1:0] pipeVectorA2_i1;
  wire signed [`W-1:0] pipeVectorA2_v;
  wire signed [`W-1:0] n42_i0;
  wire signed [`W-1:0] n42_i1;
  wire signed [`W-1:0] n42_i2;
  wire signed [`W-1:0] n42_v;
  wire signed [`W-1:0] n43_i0;
  wire signed [`W-1:0] n43_i1;
  wire signed [`W-1:0] n43_i2;
  wire signed [`W-1:0] n43_i3;
  wire signed [`W-1:0] n43_i4;
  wire signed [`W-1:0] n43_i5;
  wire signed [`W-1:0] n43_i6;
  wire signed [`W-1:0] n43_i7;
  wire signed [`W-1:0] n43_i8;
  wire signed [`W-1:0] n43_i9;
  wire signed [`W-1:0] n43_i10;
  wire signed [`W-1:0] n43_i11;
  wire signed [`W-1:0] n43_i12;
  wire signed [`W-1:0] n43_i13;
  wire signed [`W-1:0] n43_i14;
  wire signed [`W-1:0] n43_i15;
  wire signed [`W-1:0] n43_v;
  wire signed [`W-1:0] pipeT2out_i0;
  wire signed [`W-1:0] pipeT2out_i1;
  wire signed [`W-1:0] pipeT2out_i2;
  wire signed [`W-1:0] pipeT2out_v;
  wire signed [`W-1:0] dpc42_DL_ADH_i0;
  wire signed [`W-1:0] dpc42_DL_ADH_i1;
  wire signed [`W-1:0] dpc42_DL_ADH_i2;
  wire signed [`W-1:0] dpc42_DL_ADH_i3;
  wire signed [`W-1:0] dpc42_DL_ADH_i4;
  wire signed [`W-1:0] dpc42_DL_ADH_i5;
  wire signed [`W-1:0] dpc42_DL_ADH_i6;
  wire signed [`W-1:0] dpc42_DL_ADH_i7;
  wire signed [`W-1:0] dpc42_DL_ADH_i8;
  wire signed [`W-1:0] dpc42_DL_ADH_i9;
  wire signed [`W-1:0] dpc42_DL_ADH_v;
  wire signed [`W-1:0] x_op_T4_rti_i0;
  wire signed [`W-1:0] x_op_T4_rti_i1;
  wire signed [`W-1:0] x_op_T4_rti_i2;
  wire signed [`W-1:0] x_op_T4_rti_v;
  wire signed [`W-1:0] adl7_i0;
  wire signed [`W-1:0] adl7_i1;
  wire signed [`W-1:0] adl7_i2;
  wire signed [`W-1:0] adl7_i3;
  wire signed [`W-1:0] adl7_i4;
  wire signed [`W-1:0] adl7_i5;
  wire signed [`W-1:0] adl7_i6;
  wire signed [`W-1:0] adl7_i7;
  wire signed [`W-1:0] adl7_v;
  wire signed [`W-1:0] op_T0_cli_sei_i0;
  wire signed [`W-1:0] op_T0_cli_sei_i1;
  wire signed [`W-1:0] op_T0_cli_sei_i2;
  wire signed [`W-1:0] op_T0_cli_sei_v;
  wire signed [`W-1:0] n1561_i0;
  wire signed [`W-1:0] n1561_i1;
  wire signed [`W-1:0] n1561_i2;
  wire signed [`W-1:0] n1561_v;
  wire signed [`W-1:0] n1290_i0;
  wire signed [`W-1:0] n1290_i1;
  wire signed [`W-1:0] n1290_i2;
  wire signed [`W-1:0] n1290_v;
  wire signed [`W-1:0] dpc41_DL_ADL_i0;
  wire signed [`W-1:0] dpc41_DL_ADL_i1;
  wire signed [`W-1:0] dpc41_DL_ADL_i2;
  wire signed [`W-1:0] dpc41_DL_ADL_i3;
  wire signed [`W-1:0] dpc41_DL_ADL_i4;
  wire signed [`W-1:0] dpc41_DL_ADL_i5;
  wire signed [`W-1:0] dpc41_DL_ADL_i6;
  wire signed [`W-1:0] dpc41_DL_ADL_i7;
  wire signed [`W-1:0] dpc41_DL_ADL_i8;
  wire signed [`W-1:0] dpc41_DL_ADL_i9;
  wire signed [`W-1:0] dpc41_DL_ADL_v;
  wire signed [`W-1:0] nmi_i0;
  wire signed [`W-1:0] nmi_i1;
  wire signed [`W-1:0] nmi_v;
  wire signed [`W-1:0] n1566_i0;
  wire signed [`W-1:0] n1566_i1;
  wire signed [`W-1:0] n1566_i2;
  wire signed [`W-1:0] n1566_i3;
  wire signed [`W-1:0] n1566_v;
  wire signed [`W-1:0] t3_i0;
  wire signed [`W-1:0] t3_i1;
  wire signed [`W-1:0] t3_i2;
  wire signed [`W-1:0] t3_i3;
  wire signed [`W-1:0] t3_i4;
  wire signed [`W-1:0] t3_i5;
  wire signed [`W-1:0] t3_i6;
  wire signed [`W-1:0] t3_i7;
  wire signed [`W-1:0] t3_i8;
  wire signed [`W-1:0] t3_i9;
  wire signed [`W-1:0] t3_i10;
  wire signed [`W-1:0] t3_i11;
  wire signed [`W-1:0] t3_i12;
  wire signed [`W-1:0] t3_i13;
  wire signed [`W-1:0] t3_i14;
  wire signed [`W-1:0] t3_i15;
  wire signed [`W-1:0] t3_i16;
  wire signed [`W-1:0] t3_v;
  wire signed [`W-1:0] pipeUNK35_i0;
  wire signed [`W-1:0] pipeUNK35_i1;
  wire signed [`W-1:0] pipeUNK35_v;
  wire signed [`W-1:0] n474_i0;
  wire signed [`W-1:0] n474_i1;
  wire signed [`W-1:0] n474_i2;
  wire signed [`W-1:0] n474_v;
  wire signed [`W-1:0] n1712_i0;
  wire signed [`W-1:0] n1712_i1;
  wire signed [`W-1:0] n1712_i2;
  wire signed [`W-1:0] n1712_v;
  wire signed [`W-1:0] n1711_i0;
  wire signed [`W-1:0] n1711_i1;
  wire signed [`W-1:0] n1711_i2;
  wire signed [`W-1:0] n1711_v;
  wire signed [`W-1:0] op_T__cpx_cpy_imm_zp_i0;
  wire signed [`W-1:0] op_T__cpx_cpy_imm_zp_i1;
  wire signed [`W-1:0] op_T__cpx_cpy_imm_zp_i2;
  wire signed [`W-1:0] op_T__cpx_cpy_imm_zp_v;
  wire signed [`W-1:0] _TWOCYCLE_phi1_i0;
  wire signed [`W-1:0] _TWOCYCLE_phi1_i1;
  wire signed [`W-1:0] _TWOCYCLE_phi1_v;
  wire signed [`W-1:0] n1715_i0;
  wire signed [`W-1:0] n1715_i1;
  wire signed [`W-1:0] n1715_i2;
  wire signed [`W-1:0] n1715_i3;
  wire signed [`W-1:0] n1715_v;
  wire signed [`W-1:0] dpc18__DAA_i0;
  wire signed [`W-1:0] dpc18__DAA_i1;
  wire signed [`W-1:0] dpc18__DAA_i2;
  wire signed [`W-1:0] dpc18__DAA_i3;
  wire signed [`W-1:0] dpc18__DAA_i4;
  wire signed [`W-1:0] dpc18__DAA_v;
  wire signed [`W-1:0] n1714_i0;
  wire signed [`W-1:0] n1714_i1;
  wire signed [`W-1:0] n1714_i2;
  wire signed [`W-1:0] n1714_v;
  wire signed [`W-1:0] n472_i0;
  wire signed [`W-1:0] n472_i1;
  wire signed [`W-1:0] n472_i2;
  wire signed [`W-1:0] n472_v;
  wire signed [`W-1:0] n470_i0;
  wire signed [`W-1:0] n470_i1;
  wire signed [`W-1:0] n470_i2;
  wire signed [`W-1:0] n470_i3;
  wire signed [`W-1:0] n470_v;
  wire signed [`W-1:0] n471_i0;
  wire signed [`W-1:0] n471_i1;
  wire signed [`W-1:0] n471_i2;
  wire signed [`W-1:0] n471_v;
  wire signed [`W-1:0] n476_i0;
  wire signed [`W-1:0] n476_i1;
  wire signed [`W-1:0] n476_i2;
  wire signed [`W-1:0] n476_i3;
  wire signed [`W-1:0] n476_v;
  wire signed [`W-1:0] n477_i0;
  wire signed [`W-1:0] n477_i1;
  wire signed [`W-1:0] n477_i2;
  wire signed [`W-1:0] n477_i3;
  wire signed [`W-1:0] n477_i4;
  wire signed [`W-1:0] n477_v;
  wire signed [`W-1:0] n1360_i0;
  wire signed [`W-1:0] n1360_i1;
  wire signed [`W-1:0] n1360_v;
  wire signed [`W-1:0] n475_i0;
  wire signed [`W-1:0] n475_i1;
  wire signed [`W-1:0] n475_i2;
  wire signed [`W-1:0] n475_v;
  wire signed [`W-1:0] n478_i0;
  wire signed [`W-1:0] n478_i1;
  wire signed [`W-1:0] n478_i2;
  wire signed [`W-1:0] n478_v;
  wire signed [`W-1:0] n479_i0;
  wire signed [`W-1:0] n479_i1;
  wire signed [`W-1:0] n479_i2;
  wire signed [`W-1:0] n479_v;
  wire signed [`W-1:0] n1368_i0;
  wire signed [`W-1:0] n1368_i1;
  wire signed [`W-1:0] n1368_i2;
  wire signed [`W-1:0] n1368_v;
  wire signed [`W-1:0] n1369_i0;
  wire signed [`W-1:0] n1369_i1;
  wire signed [`W-1:0] n1369_i2;
  wire signed [`W-1:0] n1369_i3;
  wire signed [`W-1:0] n1369_v;

  spice_pin_input pin_irq(irq, irq_v, irq_i1);
  spice_pin_input pin_clk0(clk0, clk0_v, clk0_i2);
  spice_pin_input pin_rdy(rdy, rdy_v, rdy_i2);
  spice_pin_input pin_res(res, res_v, res_i1);
  spice_pin_input pin_so(so, so_v, so_i2);
  spice_pin_input pin_nmi(nmi, nmi_v, nmi_i1);

  spice_pin_output pin_clk1out(clk1out, clk1out_v, clk1out_i2);
  spice_pin_output pin_ab4(ab4, ab4_v, ab4_i2);
  spice_pin_output pin_ab5(ab5, ab5_v, ab5_i2);
  spice_pin_output pin_ab6(ab6, ab6_v, ab6_i2);
  spice_pin_output pin_ab7(ab7, ab7_v, ab7_i2);
  spice_pin_output pin_ab0(ab0, ab0_v, ab0_i2);
  spice_pin_output pin_ab1(ab1, ab1_v, ab1_i2);
  spice_pin_output pin_ab2(ab2, ab2_v, ab2_i2);
  spice_pin_output pin_ab3(ab3, ab3_v, ab3_i2);
  spice_pin_output pin_ab8(ab8, ab8_v, ab8_i2);
  spice_pin_output pin_ab9(ab9, ab9_v, ab9_i2);
  spice_pin_output pin_ab15(ab15, ab15_v, ab15_i2);
  spice_pin_output pin_ab14(ab14, ab14_v, ab14_i2);
  spice_pin_output pin_ab12(ab12, ab12_v, ab12_i2);
  spice_pin_output pin_ab13(ab13, ab13_v, ab13_i2);
  spice_pin_output pin_ab10(ab10, ab10_v, ab10_i2);
  spice_pin_output pin_rw(rw, rw_v, rw_i2);
  spice_pin_output pin_sync(sync, sync_v, sync_i2);
  spice_pin_output pin_ab11(ab11, ab11_v, ab11_i2);
  spice_pin_output pin_clk2out(clk2out, clk2out_v, clk2out_i2);

  spice_pin_bidirectional pin_db5(db5_i, db5_o, db5_t, db5_v, db5_i4);
  spice_pin_bidirectional pin_db7(db7_i, db7_o, db7_t, db7_v, db7_i4);
  spice_pin_bidirectional pin_db1(db1_i, db1_o, db1_t, db1_v, db1_i4);
  spice_pin_bidirectional pin_db0(db0_i, db0_o, db0_t, db0_v, db0_i4);
  spice_pin_bidirectional pin_db4(db4_i, db4_o, db4_t, db4_v, db4_i4);
  spice_pin_bidirectional pin_db6(db6_i, db6_o, db6_t, db6_v, db6_i4);
  spice_pin_bidirectional pin_db3(db3_i, db3_o, db3_t, db3_v, db3_i4);
  spice_pin_bidirectional pin_db2(db2_i, db2_o, db2_t, db2_v, db2_i4);

  spice_transistor_nmos t3489(~dpc13_ORS_v[`W-1], aluanorb1_v, notaluoutmux1_v, aluanorb1_i1, notaluoutmux1_i5);
  spice_transistor_nmos t3485(~cclk_v[`W-1], n1594_v, n688_v, n1594_i0, n688_i0);
  spice_transistor_nmos_gnd t3486(~n1395_v[`W-1], Reset0_v, Reset0_i2);
  spice_transistor_nmos_vdd t176(~n714_v[`W-1], dpc19_ADDSB7_v, dpc19_ADDSB7_i0);
  spice_transistor_nmos t170(~cclk_v[`W-1], _ABL5_v, n210_v, _ABL5_i0, n210_i0);
  spice_transistor_nmos_vdd t2572(~n1639_v[`W-1], ab15_v, ab15_i1);
  spice_transistor_nmos_vdd t2570(~n1541_v[`W-1], dpc10_ADLADD_v, dpc10_ADLADD_i2);
  spice_transistor_nmos_gnd g_1303((~n600_v[`W-1]|~n8_v[`W-1]), n36_v, n36_i1);
  spice_transistor_nmos t2683(~dpc9_DBADD_v[`W-1], alub7_v, idb7_v, alub7_i0, idb7_i7);
  spice_transistor_nmos_gnd t2682(~idb1_v[`W-1], n243_v, n243_i0);
  spice_transistor_nmos g_1429((~ADH_ABH_v[`W-1]&~cp1_v[`W-1]), _ABH4_v, n212_v, _ABH4_i2, n212_i2);
  spice_transistor_nmos t2684(~dpc9_DBADD_v[`W-1], alub6_v, idb6_v, alub6_i0, idb6_i9);
  spice_transistor_nmos_gnd g_1399((~n1720_v[`W-1]|~RnWstretched_v[`W-1]), n373_v, n373_i2);
  spice_transistor_nmos_gnd g_1398((~n689_v[`W-1]|~notRdy0_v[`W-1]), VEC0_v, VEC0_i4);
  spice_transistor_nmos_gnd g_1397((~clearIR_v[`W-1]|~pd3_v[`W-1]), pd3_clearIR_v, pd3_clearIR_i3);
  spice_transistor_nmos_gnd g_1396((~notalucout_v[`W-1]|~n1218_v[`W-1]), n1257_v, n1257_i2);
  spice_transistor_nmos_gnd t613(~clock1_v[`W-1], op_T0_v, op_T0_i1);
  spice_transistor_nmos_gnd g_1082((~alucout_v[`W-1]|~n838_v[`W-1]), n811_v, n811_i1);
  spice_transistor_nmos_gnd g_1393((~n1002_v[`W-1]|~op_T2_abs_access_v[`W-1]|~nnT2BR_v[`W-1]|~n1286_v[`W-1]|~n862_v[`W-1]), n1211_v, n1211_i4);
  spice_transistor_nmos_gnd g_1392((~n783_v[`W-1]|~n1542_v[`W-1]), n1253_v, n1253_i1);
  spice_transistor_nmos_gnd g_1391((~op_T__iny_dey_v[`W-1]|~op_T0_tay_ldy_not_idx_v[`W-1]|~op_T0_ldy_mem_v[`W-1]), n616_v, n616_i2);
  spice_transistor_nmos_gnd g_1390((~n105_v[`W-1]|~__AxB_0_v[`W-1]), _AxB_0__C0in_v, _AxB_0__C0in_i1);
  spice_transistor_nmos t2371(~dpc5_SADL_v[`W-1], adl1_v, n694_v, adl1_i4, n694_i3);
  spice_transistor_nmos t2370(~dpc24_ACSB_v[`W-1], n1592_v, sb7_v, n1592_i3, sb7_i9);
  spice_transistor_nmos_gnd t2373(~pchp0_v[`W-1], n1722_v, n1722_i0);
  spice_transistor_nmos t2372(~cclk_v[`W-1], _ABL2_v, n642_v, _ABL2_i1, n642_i1);
  spice_transistor_nmos t2878(~cclk_v[`W-1], n1693_v, n264_v, n1693_i0, n264_i1);
  spice_transistor_nmos t3178(~dpc39_PCLPCL_v[`W-1], pcl0_v, n488_v, pcl0_i1, n488_i3);
  spice_transistor_nmos t3179(~dpc39_PCLPCL_v[`W-1], pcl3_v, n723_v, pcl3_i1, n723_i3);
  spice_transistor_nmos t3174(~dpc39_PCLPCL_v[`W-1], pcl4_v, n208_v, pcl4_i1, n208_i3);
  spice_transistor_nmos t2476(~dpc31_PCHPCH_v[`W-1], pch7_v, n1206_v, pch7_i2, n1206_i1);
  spice_transistor_nmos t3176(~dpc39_PCLPCL_v[`W-1], pcl6_v, n1458_v, pcl6_i1, n1458_i3);
  spice_transistor_nmos t3177(~dpc39_PCLPCL_v[`W-1], pcl1_v, n976_v, pcl1_i1, n976_i2);
  spice_transistor_nmos_gnd t3172(~n366_v[`W-1], op_SRS_v, op_SRS_i2);
  spice_transistor_nmos t3173(~dpc39_PCLPCL_v[`W-1], pcl5_v, n72_v, pcl5_i1, n72_i3);
  spice_transistor_nmos_gnd t505(~pipeUNK21_v[`W-1], n572_v, n572_i0);
  spice_transistor_nmos_gnd g_1648(((~_DA_ADD1_v[`W-1]&~n600_v[`W-1])|(~n1682_v[`W-1]&~n8_v[`W-1])), n613_v, n613_i3);
  spice_transistor_nmos_gnd t507(~n1100_v[`W-1], ab0_v, ab0_i0);
  spice_transistor_nmos_gnd t506(~sb6_v[`W-1], n61_v, n61_i0);
  spice_transistor_nmos_gnd t501(~n1676_v[`W-1], n634_v, n634_i0);
  spice_transistor_nmos t503(~cclk_v[`W-1], notir0_v, n310_v, notir0_i1, n310_i0);
  spice_transistor_nmos_vdd t502(~n1676_v[`W-1], n86_v, n86_i0);
  spice_transistor_nmos_gnd g_1641(((~n1269_v[`W-1]&~DBNeg_v[`W-1])|(~pipeUNK01_v[`W-1]&~n1401_v[`W-1])), n626_v, n626_i2);
  spice_transistor_nmos_gnd g_1640(((~n79_v[`W-1]&(~n1343_v[`W-1]|~n877_v[`W-1]))|~n_0_ADL0_v[`W-1]), n696_v, n696_i2);
  spice_transistor_nmos_gnd g_1643((~n975_v[`W-1]|(~cclk_v[`W-1]&~n312_v[`W-1])), n854_v, n854_i3);
  spice_transistor_nmos_gnd g_1642(((~DBNeg_v[`W-1]&~n754_v[`W-1])|(~n1595_v[`W-1]&~pipeUNK13_v[`W-1])), n1181_v, n1181_i2);
  spice_transistor_nmos_gnd g_1645(((~n440_v[`W-1]&~op_inc_nop_v[`W-1])|(~op_T3_ind_x_v[`W-1]|~op_T4_ind_y_v[`W-1]|~op_plp_pla_v[`W-1]|~op_T2_ind_y_v[`W-1]|~op_T3_abs_idx_v[`W-1])), n1107_v, n1107_i2);
  spice_transistor_nmos t2478(~dpc31_PCHPCH_v[`W-1], pch5_v, n1301_v, pch5_i2, n1301_i1);
  spice_transistor_nmos_gnd g_1647((~n637_v[`W-1]|(~n1398_v[`W-1]&~C67_v[`W-1])), notaluvout_v, notaluvout_i2);
  spice_transistor_nmos_gnd g_1646(((~AxB7_v[`W-1]&~_C67_v[`W-1])|~__AxB7__C67_v[`W-1]), __AxBxC_7_v, __AxBxC_7_i2);
  spice_transistor_nmos_gnd t2645(~notidl3_v[`W-1], idl3_v, idl3_i0);
  spice_transistor_nmos t2199(~dpc27_SBADH_v[`W-1], adh2_v, sb2_v, adh2_i4, sb2_i8);
  spice_transistor_nmos t2198(~dpc27_SBADH_v[`W-1], adh3_v, sb3_v, adh3_i3, sb3_i9);
  spice_transistor_nmos_gnd t2195(~cp1_v[`W-1], n1247_v, n1247_i1);
  spice_transistor_nmos_gnd t2194(~cp1_v[`W-1], n38_v, n38_i1);
  spice_transistor_nmos t2197(~dpc27_SBADH_v[`W-1], adh4_v, dasb4_v, adh4_i4, dasb4_i9);
  spice_transistor_nmos t2191(~dpc27_SBADH_v[`W-1], sb6_v, adh6_v, sb6_i9, adh6_i3);
  spice_transistor_nmos t2190(~dpc27_SBADH_v[`W-1], adh7_v, sb7_v, adh7_i3, sb7_i7);
  spice_transistor_nmos t2193(~dpc27_SBADH_v[`W-1], adh0_v, dasb0_v, adh0_i2, dasb0_i9);
  spice_transistor_nmos t2192(~dpc1_SBY_v[`W-1], y0_v, dasb0_v, y0_i0, dasb0_i8);
  spice_transistor_nmos t2753(~cclk_v[`W-1], pipeUNK01_v, n1110_v, pipeUNK01_i0, n1110_i2);
  spice_transistor_nmos_vdd t2752(~n21_v[`W-1], dpc30_ADHPCH_v, dpc30_ADHPCH_i8);
  spice_transistor_nmos_gnd t2751(~n21_v[`W-1], n228_v, n228_i0);
  spice_transistor_nmos_gnd t2209(~n75_v[`W-1], dpc20_ADDSB06_v, dpc20_ADDSB06_i5);
  spice_transistor_nmos_vdd t2208(~n834_v[`W-1], n102_v, n102_i2);
  spice_transistor_nmos_gnd t2754(~notalu7_v[`W-1], alu7_v, alu7_i2);
  spice_transistor_nmos t1882(~cp1_v[`W-1], n1181_v, n69_v, n1181_i0, n69_i0);
  spice_transistor_nmos t1883(~cclk_v[`W-1], _ABL7_v, n171_v, _ABL7_i1, n171_i1);
  spice_transistor_nmos_vdd t1880(~n1295_v[`W-1], dpc25_SBDB_v, dpc25_SBDB_i9);
  spice_transistor_nmos t1881(~cclk_v[`W-1], n1209_v, n663_v, n1209_i0, n663_i0);
  spice_transistor_nmos_gnd t1886(~n799_v[`W-1], n1339_v, n1339_i1);
  spice_transistor_nmos_gnd t1887(~n643_v[`W-1], db3_v, db3_i2);
  spice_transistor_nmos_gnd g_1359((~notir1_v[`W-1]|~notir7_v[`W-1]|~ir5_v[`W-1]|~ir6_v[`W-1]), op_from_x_v, op_from_x_i1);
  spice_transistor_nmos_vdd t2643(~n625_v[`W-1], dpc3_SBX_v, dpc3_SBX_i8);
  spice_transistor_nmos_gnd t1408(~nots1_v[`W-1], n694_v, n694_i2);
  spice_transistor_nmos_gnd t1409(~n321_v[`W-1], n849_v, n849_i0);
  spice_transistor_nmos t1407(~cp1_v[`W-1], n533_v, n599_v, n533_i0, n599_i1);
  spice_transistor_nmos_gnd t1404(~nots3_v[`W-1], n998_v, n998_i2);
  spice_transistor_nmos_gnd t1402(~ir7_v[`W-1], notir7_v, notir7_i0);
  spice_transistor_nmos_gnd t1403(~n1304_v[`W-1], n1688_v, n1688_i0);
  spice_transistor_nmos_gnd t1400(~db0_v[`W-1], n93_v, n93_i0);
  spice_transistor_nmos_gnd t1401(~a2_v[`W-1], n419_v, n419_i0);
  spice_transistor_nmos_gnd t967(~n368_v[`W-1], n218_v, n218_i0);
  spice_transistor_nmos t1331(~cclk_v[`W-1], n831_v, a5_v, n831_i0, a5_i0);
  spice_transistor_nmos_gnd t1996(~n334_v[`W-1], n118_v, n118_i0);
  spice_transistor_nmos_gnd t1082(~dpc12_0ADD_v[`W-1], alua6_v, alua6_i1);
  spice_transistor_nmos_gnd t1083(~dpc12_0ADD_v[`W-1], alua5_v, alua5_i1);
  spice_transistor_nmos_gnd t1080(~dpc12_0ADD_v[`W-1], alua1_v, alua1_i1);
  spice_transistor_nmos_gnd t1081(~dpc12_0ADD_v[`W-1], alua4_v, alua4_i1);
  spice_transistor_nmos_gnd t1086(~notalucin_v[`W-1], n105_v, n105_i0);
  spice_transistor_nmos t963(~dpc6_SBS_v[`W-1], dasb0_v, s0_v, dasb0_i3, s0_i1);
  spice_transistor_nmos_gnd t1089(~n37_v[`W-1], db2_v, db2_i1);
  spice_transistor_nmos t962(~cclk_v[`W-1], n1694_v, x2_v, n1694_i0, x2_i0);
  spice_transistor_nmos_gnd t1310(~idb1_v[`W-1], n1474_v, n1474_i0);
  spice_transistor_nmos_gnd t985(~n790_v[`W-1], op_rmw_v, op_rmw_i0);
  spice_transistor_nmos t1315(~cclk_v[`W-1], _ABL3_v, n138_v, _ABL3_i0, n138_i2);
  spice_transistor_nmos t989(~dpc37_PCLDB_v[`W-1], idb0_v, n488_v, idb0_i6, n488_i1);
  spice_transistor_nmos_gnd t988(~sb1_v[`W-1], n320_v, n320_i0);
  spice_transistor_nmos_gnd t1319(~n653_v[`W-1], n390_v, n390_i0);
  spice_transistor_nmos_gnd t2577(~pipeUNK29_v[`W-1], n1511_v, n1511_i0);
  spice_transistor_nmos_gnd t1538(~pipeUNK42_v[`W-1], n253_v, n253_i0);
  spice_transistor_nmos_gnd t1531(~_ABL2_v[`W-1], abl2_v, abl2_i3);
  spice_transistor_nmos_vdd t1536(~n520_v[`W-1], db2_v, db2_i2);
  spice_transistor_nmos_gnd t1534(~a5_v[`W-1], n1719_v, n1719_i0);
  spice_transistor_nmos_vdd t1515(~n288_v[`W-1], n794_v, n794_i0);
  spice_transistor_nmos_vdd t1516(~abh0_v[`W-1], n826_v, n826_i1);
  spice_transistor_nmos_gnd t1474(~n595_v[`W-1], n992_v, n992_i0);
  spice_transistor_nmos_gnd t1693(~n1124_v[`W-1], n1662_v, n1662_i0);
  spice_transistor_nmos t3418(~cclk_v[`W-1], n696_v, n610_v, n696_i0, n610_i1);
  spice_transistor_nmos_gnd g_1238((~ir4_v[`W-1]|~t3_v[`W-1]|~notir3_v[`W-1]|~notir2_v[`W-1]), op_T3_mem_abs_v, op_T3_mem_abs_i2);
  spice_transistor_nmos_gnd g_1239((~ir6_v[`W-1]|~ir2_v[`W-1]|~notir1_v[`W-1]|~notir3_v[`W-1]|~clock2_v[`W-1]|~ir4_v[`W-1]|~ir7_v[`W-1]), op_T__asl_rol_a_v, op_T__asl_rol_a_i1);
  spice_transistor_nmos t1690(~cp1_v[`W-1], n1093_v, n226_v, n1093_i0, n226_i0);
  spice_transistor_nmos_gnd g_1307((~notir1_v[`W-1]|~notir7_v[`W-1]|~notir5_v[`W-1]|~notir6_v[`W-1]), op_inc_nop_v, op_inc_nop_i1);
  spice_transistor_nmos_gnd t1697(~n226_v[`W-1], n1593_v, n1593_i2);
  spice_transistor_nmos_gnd t1626(~db5_v[`W-1], n1588_v, n1588_i1);
  spice_transistor_nmos_gnd t1627(~n747_v[`W-1], n1417_v, n1417_i2);
  spice_transistor_nmos t1624(~cclk_v[`W-1], notaluoutmux1_v, notalu1_v, notaluoutmux1_i3, notalu1_i1);
  spice_transistor_nmos t1620(~cclk_v[`W-1], pipeUNK26_v, n132_v, pipeUNK26_i1, n132_i0);
  spice_transistor_nmos t1621(~cclk_v[`W-1], n1254_v, _ABL6_v, n1254_i1, _ABL6_i1);
  spice_transistor_nmos_gnd t1694(~n1269_v[`W-1], n1401_v, n1401_i0);
  spice_transistor_nmos_gnd g_1236((~n1002_v[`W-1]|~n952_v[`W-1]|~n630_v[`W-1]|~op_T2_v[`W-1]), n152_v, n152_i1);
  spice_transistor_nmos_gnd t1628(~pd6_clearIR_v[`W-1], n1309_v, n1309_i0);
  spice_transistor_nmos_gnd t1629(~_op_branch_bit7_v[`W-1], n201_v, n201_i0);
  spice_transistor_nmos_gnd t3410(~n794_v[`W-1], db1_v, db1_i3);
  spice_transistor_nmos_gnd g_1230((~ir4_v[`W-1]|~ir2_v[`W-1]|~t2_v[`W-1]|~irline3_v[`W-1]|~ir7_v[`W-1]), op_T2_stack_access_v, op_T2_stack_access_i2);
  spice_transistor_nmos_gnd g_1353((~n1398_v[`W-1]|~n748_v[`W-1]), AxB7_v, AxB7_i3);
  spice_transistor_nmos_gnd g_1111((~ir3_v[`W-1]|~ir6_v[`W-1]|~ir7_v[`W-1]|~ir2_v[`W-1]|~ir4_v[`W-1]|~notir5_v[`W-1]|~irline3_v[`W-1]), op_jsr_v, op_jsr_i2);
  spice_transistor_nmos t2632(~cp1_v[`W-1], p1_v, n566_v, p1_i1, n566_i0);
  spice_transistor_nmos_gnd g_1351((~dor7_v[`W-1]|~RnWstretched_v[`W-1]), n1501_v, n1501_i2);
  spice_transistor_nmos_gnd t189(~n408_v[`W-1], aluvout_v, aluvout_i0);
  spice_transistor_nmos g_1436((~ADL_ABL_v[`W-1]&~cp1_v[`W-1]), _ABL5_v, n1094_v, _ABL5_i2, n1094_i2);
  spice_transistor_nmos t181(~cp1_v[`W-1], n1141_v, n101_v, n1141_i0, n101_i0);
  spice_transistor_nmos t180(~cclk_v[`W-1], n779_v, n805_v, n779_i0, n805_i0);
  spice_transistor_nmos t182(~cclk_v[`W-1], n408_v, notaluvout_v, n408_i0, notaluvout_i0);
  spice_transistor_nmos_gnd t185(~notidl6_v[`W-1], idl6_v, idl6_i0);
  spice_transistor_nmos_gnd t349(~ir0_v[`W-1], notir0_v, notir0_i0);
  spice_transistor_nmos_gnd t347(~op_T3_jmp_v[`W-1], n980_v, n980_i0);
  spice_transistor_nmos_vdd t345(~n525_v[`W-1], dpc26_ACDB_v, dpc26_ACDB_i0);
  spice_transistor_nmos_gnd t344(~n525_v[`W-1], n800_v, n800_i0);
  spice_transistor_nmos_gnd t343(~n1305_v[`W-1], dpc17_SUMS_v, dpc17_SUMS_i0);
  spice_transistor_nmos_gnd t340(~n1452_v[`W-1], n861_v, n861_i0);
  spice_transistor_nmos t1958(~dpc13_ORS_v[`W-1], aluanorb0_v, notaluoutmux0_v, aluanorb0_i0, notaluoutmux0_i3);
  spice_transistor_nmos_gnd g_1437((~n523_v[`W-1]&(~dpc35_PCHC_v[`W-1]|~n83_v[`W-1])), n1657_v, n1657_i2);
  spice_transistor_nmos_gnd t1959(~n947_v[`W-1], n1654_v, n1654_i1);
  spice_transistor_nmos_gnd t3365(~adl5_v[`W-1], n1094_v, n1094_i0);
  spice_transistor_nmos_gnd g_1394((~n1113_v[`W-1]|~cclk_v[`W-1]), n161_v, n161_i3);
  spice_transistor_nmos_gnd g_1421((~n813_v[`W-1]&~n46_v[`W-1]), n1101_v, n1101_i2);
  spice_transistor_nmos_gnd t1955(~n1230_v[`W-1], n708_v, n708_i0);
  spice_transistor_nmos t72(~dpc1_SBY_v[`W-1], y6_v, sb6_v, y6_i1, sb6_i1);
  spice_transistor_nmos t73(~cp1_v[`W-1], n920_v, n785_v, n920_i0, n785_i0);
  spice_transistor_nmos_vdd t76(~n127_v[`W-1], clk2out_v, clk2out_i0);
  spice_transistor_nmos t77(~dpc1_SBY_v[`W-1], y4_v, dasb4_v, y4_i0, dasb4_i2);
  spice_transistor_nmos_gnd t74(~n1318_v[`W-1], n748_v, n748_i0);
  spice_transistor_nmos_vdd t75(~dpc14_SRS_v[`W-1], n304_v, n304_i0);
  spice_transistor_nmos_gnd g_1258((~notir0_v[`W-1]|~notir6_v[`W-1]|~clock2_v[`W-1]|~notir5_v[`W-1]), x_op_T__adc_sbc_v, x_op_T__adc_sbc_i2);
  spice_transistor_nmos_gnd g_1259((~notir0_v[`W-1]|~ir5_v[`W-1]|~clock2_v[`W-1]|~notir6_v[`W-1]|~notir7_v[`W-1]), op_T__cmp_v, op_T__cmp_i1);
  spice_transistor_nmos_gnd g_1256((~notir0_v[`W-1]|~clock2_v[`W-1]|~notir6_v[`W-1]|~notir5_v[`W-1]), op_T__adc_sbc_v, op_T__adc_sbc_i2);
  spice_transistor_nmos_gnd g_1257((~ir4_v[`W-1]|~ir2_v[`W-1]|~notir3_v[`W-1]|~irline3_v[`W-1]|~ir5_v[`W-1]|~notir7_v[`W-1]|~clock2_v[`W-1]), op_T__iny_dey_v, op_T__iny_dey_i1);
  spice_transistor_nmos_gnd g_1252((~n964_v[`W-1]|~n732_v[`W-1]), clock1_v, clock1_i33);
  spice_transistor_nmos_gnd g_1253((~n604_v[`W-1]|~n1377_v[`W-1]), n385_v, n385_i2);
  spice_transistor_nmos_gnd g_1250((~t3_v[`W-1]|~notir3_v[`W-1]|~notir4_v[`W-1]), x_op_T3_abs_idx_v, x_op_T3_abs_idx_i2);
  spice_transistor_nmos_vdd t3501(~n951_v[`W-1], n642_v, n642_i3);
  spice_transistor_nmos_gnd t2569(~n1541_v[`W-1], n491_v, n491_i0);
  spice_transistor_nmos_vdd t167(~dor5_v[`W-1], n373_v, n373_i0);
  spice_transistor_nmos_vdd t166(~n1296_v[`W-1], ab11_v, ab11_i0);
  spice_transistor_nmos_gnd t162(~n272_v[`W-1], n952_v, n952_i0);
  spice_transistor_nmos_vdd t2270(~cclk_v[`W-1], idb5_v, idb5_i5);
  spice_transistor_nmos t2272(~cclk_v[`W-1], n440_v, pipeUNK39_v, n440_i0, pipeUNK39_i0);
  spice_transistor_nmos_gnd g_1277((~n1357_v[`W-1]|~n18_v[`W-1]), n378_v, n378_i3);
  spice_transistor_nmos_gnd t2274(~op_T3_branch_v[`W-1], n1708_v, n1708_i1);
  spice_transistor_nmos_gnd t2276(~pclp4_v[`W-1], n208_v, n208_i0);
  spice_transistor_nmos_gnd g_1410((~n1357_v[`W-1]|~n1360_v[`W-1]), n1575_v, n1575_i3);
  spice_transistor_nmos_gnd g_1412((~RnWstretched_v[`W-1]|~dor1_v[`W-1]), n794_v, n794_i2);
  spice_transistor_nmos_gnd g_1413((~n266_v[`W-1]|~cclk_v[`W-1]), n525_v, n525_i3);
  spice_transistor_nmos_gnd g_1414((~n923_v[`W-1]|~n293_v[`W-1]), n810_v, n810_i1);
  spice_transistor_nmos_gnd g_1416((~n1177_v[`W-1]|~pipeUNK03_v[`W-1]|~n1111_v[`W-1]), n1614_v, n1614_i1);
  spice_transistor_nmos t2363(~dpc24_ACSB_v[`W-1], dasb0_v, n146_v, dasb0_i10, n146_i2);
  spice_transistor_nmos t2366(~dpc24_ACSB_v[`W-1], sb3_v, n1654_v, sb3_i10, n1654_i3);
  spice_transistor_nmos t2367(~dpc24_ACSB_v[`W-1], dasb4_v, n1344_v, dasb4_i11, n1344_i1);
  spice_transistor_nmos t2364(~dpc24_ACSB_v[`W-1], sb1_v, n929_v, sb1_i9, n929_i3);
  spice_transistor_nmos t2365(~dpc24_ACSB_v[`W-1], n1618_v, sb2_v, n1618_i1, sb2_i9);
  spice_transistor_nmos t2368(~dpc24_ACSB_v[`W-1], sb5_v, n831_v, sb5_i8, n831_i2);
  spice_transistor_nmos t2369(~dpc24_ACSB_v[`W-1], n326_v, sb6_v, n326_i3, sb6_i11);
  spice_transistor_nmos_gnd g_1098((~clearIR_v[`W-1]|~pd0_v[`W-1]), pd0_clearIR_v, pd0_clearIR_i2);
  spice_transistor_nmos_gnd g_1099((~clearIR_v[`W-1]|~pd5_v[`W-1]), pd5_clearIR_v, pd5_clearIR_i2);
  spice_transistor_nmos_gnd g_1094((~x_op_T4_ind_y_v[`W-1]|~x_op_T3_abs_idx_v[`W-1]), n261_v, n261_i2);
  spice_transistor_nmos_gnd t3103(~n1254_v[`W-1], ab6_v, ab6_i1);
  spice_transistor_nmos_gnd t3102(~pipeUNK41_v[`W-1], n1497_v, n1497_i1);
  spice_transistor_nmos_gnd g_1090((~n1130_v[`W-1]|~n267_v[`W-1]), n80_v, n80_i2);
  spice_transistor_nmos_gnd g_1091((~n1708_v[`W-1]|~n771_v[`W-1]), n1055_v, n1055_i1);
  spice_transistor_nmos_gnd g_1674(((~_C56_v[`W-1]&~n336_v[`W-1])|~n1084_v[`W-1]), C67_v, C67_i5);
  spice_transistor_nmos_gnd g_1676((((~n646_v[`W-1]|(~nnT2BR_v[`W-1]&~BRtaken_v[`W-1]))&~n372_v[`W-1])|(~n862_v[`W-1]&~notRdy0_v[`W-1])), n1085_v, n1085_i2);
  spice_transistor_nmos_gnd g_1671(((~notRdy0_v[`W-1]&~pipeT3out_v[`W-1])|(~n16_v[`W-1]&~pipeT2out_v[`W-1])), n428_v, n428_i2);
  spice_transistor_nmos_gnd g_1672(((~op_T2_ADL_ADD_v[`W-1]&~n638_v[`W-1])|(~op_T2_stack_v[`W-1]|~notRdy0_v[`W-1]|~op_T4_brk_jsr_v[`W-1]|~op_T3_ind_x_v[`W-1]|~op_T4_rti_v[`W-1]|~op_T3_stack_bit_jmp_v[`W-1])), n604_v, n604_i4);
  spice_transistor_nmos_gnd g_1673((~op_T2_stack_v[`W-1]|(~n1289_v[`W-1]&~op_T0_jsr_v[`W-1])), n632_v, n632_i2);
  spice_transistor_nmos_gnd g_1095((~op_T3_abs_idx_ind_v[`W-1]|~x_op_T4_ind_y_v[`W-1]|~op_T5_rts_v[`W-1]|~op_T5_ind_x_v[`W-1]), n726_v, n726_i2);
  spice_transistor_nmos_vdd t570(~n772_v[`W-1], dpc17_SUMS_v, dpc17_SUMS_i1);
  spice_transistor_nmos_gnd t571(~s5_v[`W-1], n496_v, n496_i1);
  spice_transistor_nmos_gnd t572(~pclp2_v[`W-1], n481_v, n481_i0);
  spice_transistor_nmos_gnd g_1070((~n1247_v[`W-1]|~cclk_v[`W-1]|~n800_v[`W-1]), dpc26_ACDB_v, dpc26_ACDB_i9);
  spice_transistor_nmos_vdd t578(~dor2_v[`W-1], n520_v, n520_i0);
  spice_transistor_nmos_gnd g_1078((~alub3_v[`W-1]|~alua3_v[`W-1]), n649_v, n649_i3);
  spice_transistor_nmos_gnd g_1079((~n71_v[`W-1]|~cclk_v[`W-1]|~n1247_v[`W-1]), dpc7_SS_v, dpc7_SS_i9);
  spice_transistor_nmos_gnd t2189(~n890_v[`W-1], n1694_v, n1694_i1);
  spice_transistor_nmos_gnd t2184(~p3_v[`W-1], n1194_v, n1194_i2);
  spice_transistor_nmos_gnd t2185(~n350_v[`W-1], n988_v, n988_i0);
  spice_transistor_nmos_gnd t2180(~n398_v[`W-1], n321_v, n321_i2);
  spice_transistor_nmos_gnd t2748(~n698_v[`W-1], VEC1_v, VEC1_i1);
  spice_transistor_nmos t2218(~dpc15_ANDS_v[`W-1], n336_v, n722_v, n336_i1, n722_i5);
  spice_transistor_nmos t2219(~dpc15_ANDS_v[`W-1], n304_v, n1318_v, n304_i4, n1318_i2);
  spice_transistor_nmos t2216(~dpc15_ANDS_v[`W-1], n1063_v, n296_v, n1063_i1, n296_i4);
  spice_transistor_nmos t2217(~dpc15_ANDS_v[`W-1], n277_v, n477_v, n277_i4, n477_i2);
  spice_transistor_nmos t2214(~dpc15_ANDS_v[`W-1], n681_v, n740_v, n681_i1, n740_i4);
  spice_transistor_nmos t2212(~dpc15_ANDS_v[`W-1], aluanandb0_v, notaluoutmux0_v, aluanandb0_i0, notaluoutmux0_i5);
  spice_transistor_nmos t2213(~dpc15_ANDS_v[`W-1], aluanandb1_v, notaluoutmux1_v, aluanandb1_i1, notaluoutmux1_i4);
  spice_transistor_nmos_gnd t2210(~C45_v[`W-1], _C45_v, _C45_i1);
  spice_transistor_nmos_gnd g_1097((~n954_v[`W-1]|~op_T__bit_v[`W-1]|~n885_v[`W-1]), n513_v, n513_i2);
  spice_transistor_nmos_gnd t880(~idb2_v[`W-1], n458_v, n458_i0);
  spice_transistor_nmos_gnd t881(~pchp4_v[`W-1], n27_v, n27_i0);
  spice_transistor_nmos_gnd t883(~pcl5_v[`W-1], n386_v, n386_i0);
  spice_transistor_nmos_gnd t404(~db3_v[`W-1], n1281_v, n1281_i0);
  spice_transistor_nmos_gnd t405(~_C56_v[`W-1], C56_v, C56_i0);
  spice_transistor_nmos t407(~cclk_v[`W-1], n878_v, n462_v, n878_i0, n462_i0);
  spice_transistor_nmos t402(~cp1_v[`W-1], p2_v, n845_v, p2_i0, n845_i0);
  spice_transistor_nmos_gnd t1983(~n1033_v[`W-1], dpc21_ADDADL_v, dpc21_ADDADL_i9);
  spice_transistor_nmos_gnd t1982(~idb3_v[`W-1], n457_v, n457_i1);
  spice_transistor_nmos_gnd t1980(~adh4_v[`W-1], n212_v, n212_i0);
  spice_transistor_nmos_gnd t978(~n1585_v[`W-1], n962_v, n962_i0);
  spice_transistor_nmos_gnd t1329(~dpc22__DSA_v[`W-1], n306_v, n306_i0);
  spice_transistor_nmos_gnd t1327(~n1484_v[`W-1], n1491_v, n1491_i1);
  spice_transistor_nmos_vdd t1322(~n866_v[`W-1], n9_v, n9_i0);
  spice_transistor_nmos_gnd g_1192((~ir4_v[`W-1]|~ir2_v[`W-1]|~t5_v[`W-1]|~ir5_v[`W-1]|~irline3_v[`W-1]|~ir6_v[`W-1]|~ir3_v[`W-1]|~ir7_v[`W-1]), op_T5_brk_v, op_T5_brk_i2);
  spice_transistor_nmos t1508(~dpc0_YSB_v[`W-1], sb3_v, n1531_v, sb3_i5, n1531_i0);
  spice_transistor_nmos_gnd g_1331((~n1691_v[`W-1]|~DA_AB2_v[`W-1]), DA_AxB2_v, DA_AxB2_i2);
  spice_transistor_nmos_gnd g_1160((~notir2_v[`W-1]|~t2_v[`W-1]|~notir4_v[`W-1]), op_T2_idx_x_xy_v, op_T2_idx_x_xy_i1);
  spice_transistor_nmos_gnd t3153(~n130_v[`W-1], ADL_ABL_v, ADL_ABL_i1);
  spice_transistor_nmos_gnd g_1161((~ir4_v[`W-1]|~notir3_v[`W-1]|~notir2_v[`W-1]|~t2_v[`W-1]), op_T2_abs_v, op_T2_abs_i1);
  spice_transistor_nmos_gnd g_1162((~notir2_v[`W-1]|~ir7_v[`W-1]|~ir4_v[`W-1]|~notir6_v[`W-1]|~notir3_v[`W-1]|~irline3_v[`W-1]), op_jmp_v, op_jmp_i1);
  spice_transistor_nmos_gnd t1189(~n526_v[`W-1], pclp0_v, pclp0_i1);
  spice_transistor_nmos_gnd t1188(~n1392_v[`W-1], n284_v, n284_i0);
  spice_transistor_nmos t1183(~cclk_v[`W-1], x1_v, n1709_v, x1_i0, n1709_i0);
  spice_transistor_nmos_vdd t1182(~abl1_v[`W-1], n1479_v, n1479_i0);
  spice_transistor_nmos_gnd t1181(~abl1_v[`W-1], n842_v, n842_i0);
  spice_transistor_nmos_gnd t1180(~abl1_v[`W-1], n66_v, n66_i1);
  spice_transistor_nmos t1185(~cp1_v[`W-1], n562_v, n645_v, n562_i0, n645_i0);
  spice_transistor_nmos_gnd t1184(~n_0_ADL1_v[`W-1], adl1_v, adl1_i1);
  spice_transistor_nmos_gnd g_1166((~ir4_v[`W-1]|~notir2_v[`W-1]|~ir7_v[`W-1]|~clock1_v[`W-1]|~irline3_v[`W-1]|~ir6_v[`W-1]|~notir5_v[`W-1]), op_T0_bit_v, op_T0_bit_i1);
  spice_transistor_nmos_gnd g_1194((~cclk_v[`W-1]|~n1247_v[`W-1]|~n441_v[`W-1]), dpc1_SBY_v, dpc1_SBY_i9);
  spice_transistor_nmos_gnd g_1167((~ir7_v[`W-1]|~ir4_v[`W-1]|~notir2_v[`W-1]|~notir3_v[`W-1]|~notir6_v[`W-1]|~t3_v[`W-1]|~irline3_v[`W-1]), op_T3_jmp_v, op_T3_jmp_i2);
  spice_transistor_nmos t1616(~cclk_v[`W-1], n896_v, notidl3_v, n896_i0, notidl3_i0);
  spice_transistor_nmos t1615(~cclk_v[`W-1], n436_v, x4_v, n436_i1, x4_i1);
  spice_transistor_nmos_gnd t1619(~n1045_v[`W-1], Pout7_v, Pout7_i1);
  spice_transistor_nmos_gnd t1618(~db7_v[`W-1], n588_v, n588_i0);
  spice_transistor_nmos_gnd g_1197((~n781_v[`W-1]|~n1492_v[`W-1]), n1457_v, n1457_i1);
  spice_transistor_nmos_gnd g_1666(((~n1070_v[`W-1]&~n919_v[`W-1])|~n200_v[`W-1]), n1486_v, n1486_i2);
  spice_transistor_nmos_gnd g_1196((~n662_v[`W-1]|~cclk_v[`W-1]|~n1247_v[`W-1]), dpc3_SBX_v, dpc3_SBX_i9);
  spice_transistor_nmos_gnd t3009(~n312_v[`W-1], n995_v, n995_i0);
  spice_transistor_nmos_gnd t1929(~n1450_v[`W-1], n1499_v, n1499_i0);
  spice_transistor_nmos_gnd t1928(~n1609_v[`W-1], ir5_v, ir5_i0);
  spice_transistor_nmos_gnd g_1344((~n1258_v[`W-1]|~n440_v[`W-1]), n813_v, n813_i1);
  spice_transistor_nmos_gnd t916(~n726_v[`W-1], n630_v, n630_i0);
  spice_transistor_nmos_gnd t917(~n1195_v[`W-1], n1191_v, n1191_i0);
  spice_transistor_nmos_gnd t914(~nots7_v[`W-1], n721_v, n721_i2);
  spice_transistor_nmos_gnd g_1345((~notRdy0_v[`W-1]|~pipeUNK34_v[`W-1]), n720_v, n720_i2);
  spice_transistor_nmos t915(~cclk_v[`W-1], n1225_v, pipedpc28_v, n1225_i1, pipedpc28_i0);
  spice_transistor_nmos t372(~dpc10_ADLADD_v[`W-1], adl0_v, alub0_v, adl0_i1, alub0_i0);
  spice_transistor_nmos_gnd t373(~C1x5Reset_v[`W-1], n1054_v, n1054_i0);
  spice_transistor_nmos_gnd t370(~n198_v[`W-1], n424_v, n424_i1);
  spice_transistor_nmos t374(~dpc4_SSB_v[`W-1], n694_v, sb1_v, n694_i1, sb1_i2);
  spice_transistor_nmos_gnd t375(~n869_v[`W-1], ab13_v, ab13_i1);
  spice_transistor_nmos_gnd g_1047((~notir7_v[`W-1]|~ir4_v[`W-1]|~notir6_v[`W-1]|~clock1_v[`W-1]|~irline3_v[`W-1]), op_T0_cpx_cpy_inx_iny_v, op_T0_cpx_cpy_inx_iny_i1);
  spice_transistor_nmos t2757(~cclk_v[`W-1], n1121_v, n1225_v, n1121_i1, n1225_i2);
  spice_transistor_nmos_gnd t3448(~sb7_v[`W-1], n852_v, n852_i0);
  spice_transistor_nmos t2547(~dpc32_PCHADH_v[`W-1], adh7_v, n1206_v, adh7_i5, n1206_i2);
  spice_transistor_nmos_gnd t3372(~_ABH1_v[`W-1], abh1_v, abh1_i3);
  spice_transistor_nmos_gnd t3370(~pipeUNK35_v[`W-1], n238_v, n238_i0);
  spice_transistor_nmos t3376(~dpc40_ADLPCL_v[`W-1], adl2_v, pcl2_v, adl2_i8, pcl2_i2);
  spice_transistor_nmos t3377(~dpc40_ADLPCL_v[`W-1], pcl5_v, adl5_v, pcl5_i2, adl5_i7);
  spice_transistor_nmos_gnd t2204(~y6_v[`W-1], n1439_v, n1439_i1);
  spice_transistor_nmos_gnd g_1340((~RnWstretched_v[`W-1]|~dor3_v[`W-1]), n1613_v, n1613_i2);
  spice_transistor_nmos t3378(~dpc40_ADLPCL_v[`W-1], adl4_v, pcl4_v, adl4_i7, pcl4_i2);
  spice_transistor_nmos t3379(~dpc40_ADLPCL_v[`W-1], adl6_v, pcl6_v, adl6_i7, pcl6_i2);
  spice_transistor_nmos_vdd t2544(~n839_v[`W-1], n43_v, n43_i0);
  spice_transistor_nmos_gnd t3440(~n1338_v[`W-1], n462_v, n462_i1);
  spice_transistor_nmos t2545(~cclk_v[`W-1], n484_v, pclp7_v, n484_i0, pclp7_i1);
  spice_transistor_nmos_gnd g_1249((~t3_v[`W-1]|~notir3_v[`W-1]|~notir4_v[`W-1]), op_T3_abs_idx_v, op_T3_abs_idx_i1);
  spice_transistor_nmos_gnd g_1245((~RnWstretched_v[`W-1]|~n769_v[`W-1]), n1325_v, n1325_i2);
  spice_transistor_nmos_gnd g_1244((~n1257_v[`W-1]|~n811_v[`W-1]), n753_v, n753_i1);
  spice_transistor_nmos_gnd g_1247((~ir3_v[`W-1]|~ir2_v[`W-1]|~notir0_v[`W-1]|~t5_v[`W-1]), op_T5_mem_ind_idx_v, op_T5_mem_ind_idx_i2);
  spice_transistor_nmos_gnd g_1246((~n1708_v[`W-1]|~n770_v[`W-1]), n19_v, n19_i2);
  spice_transistor_nmos_gnd g_1241((~__AxB_6_v[`W-1]|~C56_v[`W-1]), _AxB_6__C56_v, _AxB_6__C56_i1);
  spice_transistor_nmos_gnd g_1240((~dor1_v[`W-1]|~RnWstretched_v[`W-1]), n288_v, n288_i3);
  spice_transistor_nmos_gnd g_1243((~RnWstretched_v[`W-1]|~n224_v[`W-1]), n520_v, n520_i2);
  spice_transistor_nmos_gnd t3445(~n680_v[`W-1], n1526_v, n1526_i1);
  spice_transistor_nmos_gnd t2511(~idb3_v[`W-1], n1621_v, n1621_i1);
  spice_transistor_nmos_gnd t2517(~_DA_ADD1_v[`W-1], n1682_v, n1682_i0);
  spice_transistor_nmos_vdd t2516(~n1613_v[`W-1], n643_v, n643_i1);
  spice_transistor_nmos t794(~cclk_v[`W-1], pipeUNK14_v, n318_v, pipeUNK14_i0, n318_i0);
  spice_transistor_nmos_gnd t791(~notalu2_v[`W-1], alu2_v, alu2_i1);
  spice_transistor_nmos_gnd t153(~pch0_v[`W-1], n1010_v, n1010_i0);
  spice_transistor_nmos_gnd t157(~_ABL7_v[`W-1], n567_v, n567_i0);
  spice_transistor_nmos_vdd t154(~n798_v[`W-1], db1_v, db1_i1);
  spice_transistor_nmos_gnd t158(~adl6_v[`W-1], n1548_v, n1548_i0);
  spice_transistor_nmos_gnd t2543(~adl3_v[`W-1], n1507_v, n1507_i0);
  spice_transistor_nmos_gnd g_1130((~n1083_v[`W-1]|~pd2_clearIR_v[`W-1]|~n409_v[`W-1]|~pd4_clearIR_v[`W-1]), PD_xxx010x1_v, PD_xxx010x1_i1);
  spice_transistor_nmos_gnd g_1407((~n1247_v[`W-1]|~cclk_v[`W-1]|~n1335_v[`W-1]), dpc24_ACSB_v, dpc24_ACSB_i9);
  spice_transistor_nmos_gnd g_1405((~n919_v[`W-1]|~n1070_v[`W-1]), n200_v, n200_i1);
  spice_transistor_nmos_gnd g_1403((~RnWstretched_v[`W-1]|~n1463_v[`W-1]), n1076_v, n1076_i2);
  spice_transistor_nmos_gnd g_1402((~RnWstretched_v[`W-1]|~n1613_v[`W-1]), n42_v, n42_i2);
  spice_transistor_nmos_gnd g_1401((~n23_v[`W-1]|~RnWstretched_v[`W-1]), n298_v, n298_i2);
  spice_transistor_nmos_gnd g_1400((~C34_v[`W-1]|~dpc22__DSA_v[`W-1]), n1179_v, n1179_i2);
  spice_transistor_nmos_gnd g_1409((~n1697_v[`W-1]|~n773_v[`W-1]), n275_v, n275_i2);
  spice_transistor_nmos_gnd t2894(~n541_v[`W-1], ir7_v, ir7_i2);
  spice_transistor_nmos_gnd t2093(~abh4_v[`W-1], n1677_v, n1677_i2);
  spice_transistor_nmos_gnd g_1029((~irline3_v[`W-1]|~notir2_v[`W-1]|~ir6_v[`W-1]|~notir5_v[`W-1]|~ir7_v[`W-1]|~ir4_v[`W-1]|~clock2_v[`W-1]), op_T__bit_v, op_T__bit_i2);
  spice_transistor_nmos_gnd t2357(~n659_v[`W-1], ab15_v, ab15_i0);
  spice_transistor_nmos_gnd t2424(~n1255_v[`W-1], dpc13_ORS_v, dpc13_ORS_i5);
  spice_transistor_nmos_gnd t2427(~n897_v[`W-1], n1369_v, n1369_i2);
  spice_transistor_nmos_vdd t2353(~n298_v[`W-1], db7_v, db7_i2);
  spice_transistor_nmos t2351(~cclk_v[`W-1], pclp3_v, n1631_v, pclp3_i1, n1631_i0);
  spice_transistor_nmos t3118(~dpc2_XSB_v[`W-1], n1694_v, sb2_v, n1694_i2, sb2_i10);
  spice_transistor_nmos_gnd g_1088((~notRdy0_v[`W-1]|~n347_v[`W-1]|~n790_v[`W-1]), n191_v, n191_i2);
  spice_transistor_nmos_gnd t2541(~n1400_v[`W-1], n83_v, n83_i0);
  spice_transistor_nmos t3116(~dpc2_XSB_v[`W-1], n1724_v, sb6_v, n1724_i2, sb6_i12);
  spice_transistor_nmos_gnd t3117(~n1256_v[`W-1], dpc15_ANDS_v, dpc15_ANDS_i9);
  spice_transistor_nmos t3115(~dpc2_XSB_v[`W-1], n578_v, sb5_v, n578_i1, sb5_i10);
  spice_transistor_nmos_gnd g_1663((~pipeUNK40_v[`W-1]|(~notRdy0_v[`W-1]&~pipeUNK39_v[`W-1])), n1039_v, n1039_i2);
  spice_transistor_nmos_gnd g_1662(((~pipeT5out_v[`W-1]&~notRdy0_v[`W-1])|(~pipeT4out_v[`W-1]&~n16_v[`W-1])), n468_v, n468_i2);
  spice_transistor_nmos_gnd g_1661(((~n986_v[`W-1]&~n600_v[`W-1])|(~n8_v[`W-1]&~n876_v[`W-1])), n345_v, n345_i3);
  spice_transistor_nmos_gnd g_1660((~_AxB_6__C56_v[`W-1]|(~C56_v[`W-1]&~__AxB_6_v[`W-1])), __AxBxC_6_v, __AxBxC_6_i2);
  spice_transistor_nmos_gnd g_1667(((~PD_1xx000x0_v[`W-1]|~PD_xxx010x1_v[`W-1])|(~PD_xxxx10x0_v[`W-1]&~PD_n_0xx0xx0x_v[`W-1])), _TWOCYCLE_v, _TWOCYCLE_i2);
  spice_transistor_nmos_gnd g_1665(((~op_from_x_v[`W-1]&~n335_v[`W-1])|(~op_sty_cpy_mem_v[`W-1]&~n335_v[`W-1])), n1303_v, n1303_i2);
  spice_transistor_nmos_gnd g_1664(((~pipeUNK09_v[`W-1]&~pipeUNK06_v[`W-1])|~n1673_v[`W-1]), n754_v, n754_i3);
  spice_transistor_nmos_gnd g_1669((~n260_v[`W-1]|(~n852_v[`W-1]&~n1205_v[`W-1])), dasb7_v, dasb7_i2);
  spice_transistor_nmos_gnd g_1668((~n735_v[`W-1]|(~n320_v[`W-1]&~n36_v[`W-1])), dasb1_v, dasb1_i2);
  spice_transistor_nmos_gnd t567(~__AxB_6_v[`W-1], n122_v, n122_i0);
  spice_transistor_nmos_gnd t565(~n664_v[`W-1], n1697_v, n1697_i0);
  spice_transistor_nmos_gnd t569(~n772_v[`W-1], n1305_v, n1305_i1);
  spice_transistor_nmos_gnd g_1069((~clearIR_v[`W-1]|~pd2_v[`W-1]), pd2_clearIR_v, pd2_clearIR_i2);
  spice_transistor_nmos_gnd g_1068((~op_jsr_v[`W-1]|~op_brk_rti_v[`W-1]|~x_op_jmp_v[`W-1]), n134_v, n134_i1);
  spice_transistor_nmos_gnd t2738(~n1441_v[`W-1], dpc42_DL_ADH_v, dpc42_DL_ADH_i8);
  spice_transistor_nmos_gnd t2228(~n1549_v[`W-1], n929_v, n929_i1);
  spice_transistor_nmos t2731(~cclk_v[`W-1], x5_v, n578_v, x5_i2, n578_i0);
  spice_transistor_nmos_vdd t2222(~n1191_v[`W-1], ab6_v, ab6_i0);
  spice_transistor_nmos_vdd t2221(~cclk_v[`W-1], adl1_v, adl1_i3);
  spice_transistor_nmos_vdd t2227(~n1499_v[`W-1], dpc18__DAA_v, dpc18__DAA_i0);
  spice_transistor_nmos_gnd t2226(~n1499_v[`W-1], n709_v, n709_i0);
  spice_transistor_nmos t2737(~cclk_v[`W-1], n1229_v, pchp0_v, n1229_i0, pchp0_i1);
  spice_transistor_nmos_vdd t2736(~cclk_v[`W-1], adl0_v, adl0_i6);
  spice_transistor_nmos t892(~cclk_v[`W-1], pipeT4out_v, n188_v, pipeT4out_i0, n188_i0);
  spice_transistor_nmos t890(~cp1_v[`W-1], n1132_v, n1087_v, n1132_i0, n1087_i0);
  spice_transistor_nmos_gnd t896(~abh6_v[`W-1], n635_v, n635_i1);
  spice_transistor_nmos_gnd t895(~abh6_v[`W-1], n1523_v, n1523_i2);
  spice_transistor_nmos_vdd t894(~abh6_v[`W-1], n963_v, n963_i2);
  spice_transistor_nmos_gnd t418(~idb5_v[`W-1], n1383_v, n1383_i0);
  spice_transistor_nmos t417(~cclk_v[`W-1], n1187_v, nots6_v, n1187_i1, nots6_i0);
  spice_transistor_nmos_vdd t416(~cclk_v[`W-1], sb6_v, sb6_i4);
  spice_transistor_nmos t415(~dpc30_ADHPCH_v[`W-1], pch6_v, adh6_v, pch6_i0, adh6_i1);
  spice_transistor_nmos t414(~dpc30_ADHPCH_v[`W-1], pch7_v, adh7_v, pch7_i1, adh7_i1);
  spice_transistor_nmos t413(~dpc30_ADHPCH_v[`W-1], pch4_v, adh4_v, pch4_i1, adh4_i1);
  spice_transistor_nmos t412(~dpc30_ADHPCH_v[`W-1], pch5_v, adh5_v, pch5_i0, adh5_i1);
  spice_transistor_nmos t411(~dpc30_ADHPCH_v[`W-1], pch2_v, adh2_v, pch2_i0, adh2_i1);
  spice_transistor_nmos t410(~dpc30_ADHPCH_v[`W-1], pch3_v, adh3_v, pch3_i1, adh3_i2);
  spice_transistor_nmos t1338(~dpc3_SBX_v[`W-1], x1_v, sb1_v, x1_i1, sb1_i4);
  spice_transistor_nmos_gnd g_1237((~ir3_v[`W-1]|~t2_v[`W-1]|~notir2_v[`W-1]|~ir4_v[`W-1]), op_T2_mem_zp_v, op_T2_mem_zp_i2);
  spice_transistor_nmos_gnd t1999(~n1129_v[`W-1], n1467_v, n1467_i1);
  spice_transistor_nmos_gnd t1334(~n172_v[`W-1], n1633_v, n1633_i0);
  spice_transistor_nmos_vdd t1335(~n172_v[`W-1], n210_v, n210_i1);
  spice_transistor_nmos_vdd t961(~cclk_v[`W-1], idb3_v, idb3_i1);
  spice_transistor_nmos_gnd t1046(~pchp2_v[`W-1], n1496_v, n1496_i0);
  spice_transistor_nmos t1047(~cclk_v[`W-1], n1251_v, y7_v, n1251_i0, y7_i0);
  spice_transistor_nmos_gnd t1040(~adh1_v[`W-1], n1267_v, n1267_i0);
  spice_transistor_nmos_gnd t1518(~s3_v[`W-1], n34_v, n34_i1);
  spice_transistor_nmos_gnd t1519(~pchp6_v[`W-1], n652_v, n652_i0);
  spice_transistor_nmos t2798(~dpc8_nDBADD_v[`W-1], alub5_v, n1383_v, alub5_i1, n1383_i1);
  spice_transistor_nmos_gnd t1048(~adl4_v[`W-1], n1519_v, n1519_i0);
  spice_transistor_nmos t1049(~cp1_v[`W-1], n262_v, n1447_v, n262_i0, n1447_i0);
  spice_transistor_nmos_gnd g_1281((~notir3_v[`W-1]|~ir7_v[`W-1]|~ir2_v[`W-1]|~notir1_v[`W-1]|~clock1_v[`W-1]|~ir4_v[`W-1]), op_T0_shift_a_v, op_T0_shift_a_i2);
  spice_transistor_nmos_gnd t1194(~_ABH3_v[`W-1], abh3_v, abh3_i3);
  spice_transistor_nmos t1197(~cclk_v[`W-1], pipeUNK37_v, n944_v, pipeUNK37_i0, n944_i0);
  spice_transistor_nmos_gnd t1191(~_C34_v[`W-1], C34_v, C34_i0);
  spice_transistor_nmos_gnd g_1360((~ir6_v[`W-1]|~notir1_v[`W-1]|~notir7_v[`W-1]), op_xy_v, op_xy_i2);
  spice_transistor_nmos t1199(~cp1_v[`W-1], n1684_v, notdor6_v, n1684_i0, notdor6_i0);
  spice_transistor_nmos_gnd g_1067((~x_op_jmp_v[`W-1]|~n347_v[`W-1]|~op_rmw_v[`W-1]), n510_v, n510_i2);
  spice_transistor_nmos_gnd g_1287((~op_T2_jmp_abs_v[`W-1]|~op_T2_php_pha_v[`W-1]|~x_op_T3_plp_pla_v[`W-1]|~op_T5_rti_rts_v[`W-1]|~xx_op_T5_jsr_v[`W-1]|~op_T4_jmp_v[`W-1]), n368_v, n368_i2);
  spice_transistor_nmos_gnd g_1286((~alua2_v[`W-1]|~alub2_v[`W-1]), n1691_v, n1691_i3);
  spice_transistor_nmos_gnd t1317(~so_v[`W-1], n1650_v, n1650_i0);
  spice_transistor_nmos_gnd g_1427((~alub3_v[`W-1]&~alua3_v[`W-1]), n350_v, n350_i4);
  spice_transistor_nmos_gnd t1608(~n334_v[`W-1], Pout2_v, Pout2_i1);
  spice_transistor_nmos t1604(~cclk_v[`W-1], C78_phi2_v, alurawcout_v, C78_phi2_i0, alurawcout_i0);
  spice_transistor_nmos_vdd t1602(~cclk_v[`W-1], idb7_v, idb7_i3);
  spice_transistor_nmos t1603(~cclk_v[`W-1], VEC1_v, n1452_v, VEC1_i0, n1452_i1);
  spice_transistor_nmos_gnd t1937(~_ABH6_v[`W-1], abh6_v, abh6_i3);
  spice_transistor_nmos t2108(~cp1_v[`W-1], n1387_v, idl5_v, n1387_i3, idl5_i0);
  spice_transistor_nmos_gnd t2109(~n815_v[`W-1], n_0_ADL2_v, n_0_ADL2_i0);
  spice_transistor_nmos_gnd t2556(~dpc18__DAA_v[`W-1], n700_v, n700_i0);
  spice_transistor_nmos_gnd t2495(~pipeUNK37_v[`W-1], n198_v, n198_i2);
  spice_transistor_nmos_vdd t1934(~n466_v[`W-1], n471_v, n471_i1);
  spice_transistor_nmos t2550(~dpc32_PCHADH_v[`W-1], adh4_v, n27_v, adh4_i6, n27_i2);
  spice_transistor_nmos t2553(~dpc32_PCHADH_v[`W-1], adh1_v, n209_v, adh1_i6, n209_i1);
  spice_transistor_nmos_vdd t2000(~n1633_v[`W-1], ab5_v, ab5_i1);
  spice_transistor_nmos_gnd g_1213((~n1533_v[`W-1]|~pipe_T0_v[`W-1]), n964_v, n964_i2);
  spice_transistor_nmos_gnd t3439(~n1017_v[`W-1], n578_v, n578_i2);
  spice_transistor_nmos_gnd t3438(~n906_v[`W-1], dpc19_ADDSB7_v, dpc19_ADDSB7_i2);
  spice_transistor_nmos_vdd t367(~n424_v[`W-1], notRdy0_v, notRdy0_i0);
  spice_transistor_nmos_gnd t363(~n1333_v[`W-1], n906_v, n906_i0);
  spice_transistor_nmos_vdd t362(~n1129_v[`W-1], cclk_v, cclk_i24);
  spice_transistor_nmos_gnd g_1171((~C78_phi2_v[`W-1]|~DC78_phi2_v[`W-1]), notalucout_v, notalucout_i2);
  spice_transistor_nmos_gnd g_1215((~DA_AxB2_v[`W-1]|~AxB1_v[`W-1]|~n936_v[`W-1]|~DA_C01_v[`W-1]), n388_v, n388_i1);
  spice_transistor_nmos_gnd t369(~n198_v[`W-1], notRdy0_v, notRdy0_i1);
  spice_transistor_nmos_gnd g_1352((~n785_v[`W-1]|~n1175_v[`W-1]|~n544_v[`W-1]), n267_v, n267_i2);
  spice_transistor_nmos_gnd t3437(~n906_v[`W-1], n714_v, n714_i1);
  spice_transistor_nmos_gnd g_1350((~n988_v[`W-1]|~n649_v[`W-1]), AxB3_v, AxB3_i4);
  spice_transistor_nmos_gnd g_1357((~dor6_v[`W-1]|~RnWstretched_v[`W-1]), n466_v, n466_i3);
  spice_transistor_nmos t3216(~cclk_v[`W-1], n1618_v, a2_v, n1618_i3, a2_i2);
  spice_transistor_nmos_gnd g_1356((~pipeUNK19_v[`W-1]|~notRdy0_v[`W-1]|~ONEBYTE_v[`W-1]), n1275_v, n1275_i2);
  spice_transistor_nmos_gnd t1539(~n1552_v[`W-1], dpc14_SRS_v, dpc14_SRS_i2);
  spice_transistor_nmos_gnd g_1355((~n358_v[`W-1]|~cp1_v[`W-1]), n1129_v, n1129_i3);
  spice_transistor_nmos_gnd t3432(~cclk_v[`W-1], n1585_v, n1585_i1);
  spice_transistor_nmos_gnd g_1316((~notRdy0_v[`W-1]|~pipe_WR_phi2_v[`W-1]|~C1x5Reset_v[`W-1]), notRnWprepad_v, notRnWprepad_i4);
  spice_transistor_nmos_gnd t2641(~idb2_v[`W-1], n1573_v, n1573_i0);
  spice_transistor_nmos_gnd t3349(~n598_v[`W-1], n1260_v, n1260_i2);
  spice_transistor_nmos t1533(~dpc3_SBX_v[`W-1], x7_v, sb7_v, x7_i1, sb7_i2);
  spice_transistor_nmos t3347(~dpc11_SBADD_v[`W-1], sb7_v, alua7_v, sb7_i10, alua7_i1);
  spice_transistor_nmos_gnd t3346(~pipeUNK08_v[`W-1], n954_v, n954_i0);
  spice_transistor_nmos_gnd t3345(~n1049_v[`W-1], n507_v, n507_i0);
  spice_transistor_nmos_gnd t3344(~cp1_v[`W-1], n839_v, n839_i1);
  spice_transistor_nmos t3342(~cp1_v[`W-1], n1095_v, idl4_v, n1095_i3, idl4_i1);
  spice_transistor_nmos t3341(~cclk_v[`W-1], n548_v, nots7_v, n548_i1, nots7_i1);
  spice_transistor_nmos_vdd t3340(~cclk_v[`W-1], sb5_v, sb5_i12);
  spice_transistor_nmos_gnd g_1134((~n1047_v[`W-1]|~cclk_v[`W-1]|~n1247_v[`W-1]), dpc23_SBAC_v, dpc23_SBAC_i9);
  spice_transistor_nmos_vdd t15(~n1140_v[`W-1], ab9_v, ab9_i0);
  spice_transistor_nmos t17(~cp1_v[`W-1], p0_v, n1082_v, p0_i0, n1082_i0);
  spice_transistor_nmos_gnd t10(~n190_v[`W-1], n220_v, n220_i0);
  spice_transistor_nmos_vdd t11(~n38_v[`W-1], n1247_v, n1247_i0);
  spice_transistor_nmos_gnd g_1139((~n1371_v[`W-1]|~n1433_v[`W-1]|~n1293_v[`W-1]|~n307_v[`W-1]), n620_v, n620_i1);
  spice_transistor_nmos_gnd g_1278((~t2_v[`W-1]|~op_push_pull_v[`W-1]|~notir3_v[`W-1]), op_T2_abs_access_v, op_T2_abs_access_i2);
  spice_transistor_nmos_gnd g_1279((~op_push_pull_v[`W-1]|~t3_v[`W-1]|~notir3_v[`W-1]), op_T3_abs_idx_ind_v, op_T3_abs_idx_ind_i2);
  spice_transistor_nmos_gnd g_1270((~brk_done_v[`W-1]|~n238_v[`W-1]|~short_circuit_idx_add_v[`W-1]), n1215_v, n1215_i3);
  spice_transistor_nmos_gnd g_1272((~n221_v[`W-1]|~_DBE_v[`W-1]), n251_v, n251_i3);
  spice_transistor_nmos_gnd g_1273((~_op_branch_bit7_v[`W-1]|~n31_v[`W-1]|~n846_v[`W-1]), n307_v, n307_i2);
  spice_transistor_nmos_gnd g_1274((~n134_v[`W-1]|~n1276_v[`W-1]), n930_v, n930_i1);
  spice_transistor_nmos_gnd g_1275((~n1404_v[`W-1]|~cclk_v[`W-1]), n133_v, n133_i3);
  spice_transistor_nmos_gnd g_1064((~t4_v[`W-1]|~irline3_v[`W-1]|~ir2_v[`W-1]|~ir5_v[`W-1]|~ir7_v[`W-1]|~ir3_v[`W-1]|~ir4_v[`W-1]|~notir6_v[`W-1]), x_op_T4_rti_v, x_op_T4_rti_i1);
  spice_transistor_nmos t2557(~cclk_v[`W-1], _ABH0_v, n381_v, _ABH0_i1, n381_i2);
  spice_transistor_nmos t2503(~dpc8_nDBADD_v[`W-1], alub1_v, n583_v, alub1_i0, n583_i0);
  spice_transistor_nmos_gnd t2501(~adh0_v[`W-1], n1668_v, n1668_i0);
  spice_transistor_nmos t2506(~cclk_v[`W-1], n126_v, n1486_v, n126_i1, n1486_i0);
  spice_transistor_nmos_gnd t789(~n1300_v[`W-1], ir2_v, ir2_i0);
  spice_transistor_nmos_vdd t149(~n154_v[`W-1], dpc20_ADDSB06_v, dpc20_ADDSB06_i0);
  spice_transistor_nmos_gnd t148(~n154_v[`W-1], n75_v, n75_i0);
  spice_transistor_nmos_gnd t145(~idb7_v[`W-1], n789_v, n789_i0);
  spice_transistor_nmos_gnd t144(~op_T0_lda_v[`W-1], n397_v, n397_i0);
  spice_transistor_nmos_gnd t147(~idb0_v[`W-1], n624_v, n624_i0);
  spice_transistor_nmos_gnd t146(~AxB3_v[`W-1], n884_v, n884_i0);
  spice_transistor_nmos_gnd t141(~x5_v[`W-1], n1017_v, n1017_i0);
  spice_transistor_nmos t142(~cp1_v[`W-1], n1424_v, idl2_v, n1424_i0, idl2_i1);
  spice_transistor_nmos_gnd g_1472((~DA_C01_v[`W-1]&~n936_v[`W-1]), n319_v, n319_i1);
  spice_transistor_nmos g_1471((~ADH_ABH_v[`W-1]&~cp1_v[`W-1]), _ABH3_v, n883_v, _ABH3_i2, n883_i2);
  spice_transistor_nmos g_1476((~cp1_v[`W-1]&~ADH_ABH_v[`W-1]), n494_v, _ABH7_v, n494_i2, _ABH7_i2);
  spice_transistor_nmos_gnd g_1474((~n1120_v[`W-1]&~n440_v[`W-1]), n504_v, n504_i2);
  spice_transistor_nmos_gnd t1975(~n119_v[`W-1], ir1_v, ir1_i1);
  spice_transistor_nmos_gnd g_1520((~n595_v[`W-1]&~_op_branch_done_v[`W-1]), n192_v, n192_i4);
  spice_transistor_nmos_gnd t1978(~n188_v[`W-1], t4_v, t4_i0);
  spice_transistor_nmos t2348(~cclk_v[`W-1], n795_v, n360_v, n795_i1, n360_i0);
  spice_transistor_nmos_gnd t3125(~ir5_v[`W-1], notir5_v, notir5_i2);
  spice_transistor_nmos g_1523((~cp1_v[`W-1]&~fetch_v[`W-1]), n1309_v, n1675_v, n1309_i2, n1675_i2);
  spice_transistor_nmos_gnd t3123(~n1719_v[`W-1], n831_v, n831_i3);
  spice_transistor_nmos_vdd t3122(~n224_v[`W-1], n37_v, n37_i1);
  spice_transistor_nmos t3120(~dpc2_XSB_v[`W-1], n436_v, dasb4_v, n436_i2, dasb4_i12);
  spice_transistor_nmos t2340(~cclk_v[`W-1], n740_v, notalu2_v, n740_i5, notalu2_i1);
  spice_transistor_nmos_gnd t2345(~n24_v[`W-1], n440_v, n440_i1);
  spice_transistor_nmos_gnd t2346(~y0_v[`W-1], n1025_v, n1025_i1);
  spice_transistor_nmos_gnd g_1525(((~dpc34_PCLC_v[`W-1]|~n311_v[`W-1])&~n919_v[`W-1]), n1229_v, n1229_i2);
  spice_transistor_nmos_gnd g_1526(((~n200_v[`W-1]|~n1202_v[`W-1])&~n293_v[`W-1]), n1402_v, n1402_i2);
  spice_transistor_nmos_vdd t2179(~n1399_v[`W-1], cp1_v, cp1_i57);
  spice_transistor_nmos_vdd t2250(~abh2_v[`W-1], n1545_v, n1545_i1);
  spice_transistor_nmos_gnd g_1050((~notir0_v[`W-1]|~notir4_v[`W-1]|~ir2_v[`W-1]|~notir3_v[`W-1]|~t2_v[`W-1]), op_T2_abs_y_v, op_T2_abs_y_i1);
  spice_transistor_nmos_gnd g_1051((~n329_v[`W-1]|~dpc36_IPC_v[`W-1]|~n641_v[`W-1]|~n783_v[`W-1]|~n1643_v[`W-1]|~n937_v[`W-1]|~n249_v[`W-1]|~n232_v[`W-1]|~n386_v[`W-1]), dpc34_PCLC_v, dpc34_PCLC_i2);
  spice_transistor_nmos_gnd g_1052((~notir4_v[`W-1]|~notir3_v[`W-1]|~ir6_v[`W-1]|~notir7_v[`W-1]|~ir2_v[`W-1]|~ir5_v[`W-1]|~irline3_v[`W-1]|~clock1_v[`W-1]), x_op_T0_tya_v, x_op_T0_tya_i1);
  spice_transistor_nmos_gnd t2251(~abh2_v[`W-1], n1034_v, n1034_i0);
  spice_transistor_nmos_gnd g_1054((~notir7_v[`W-1]|~notir6_v[`W-1]|~ir4_v[`W-1]|~ir2_v[`W-1]|~notir3_v[`W-1]|~notir1_v[`W-1]|~clock1_v[`W-1]|~ir5_v[`W-1]), op_T0_dex_v, op_T0_dex_i1);
  spice_transistor_nmos_gnd g_1055((~notir7_v[`W-1]|~ir4_v[`W-1]|~ir2_v[`W-1]|~ir6_v[`W-1]|~notir1_v[`W-1]|~notir3_v[`W-1]|~clock1_v[`W-1]|~ir5_v[`W-1]), x_op_T0_txa_v, x_op_T0_txa_i1);
  spice_transistor_nmos_gnd g_1509((~n1345_v[`W-1]&~n1166_v[`W-1]), n1542_v, n1542_i3);
  spice_transistor_nmos t556(~cclk_v[`W-1], n718_v, notidl0_v, n718_i0, notidl0_i0);
  spice_transistor_nmos g_1504((~ADH_ABH_v[`W-1]&~cp1_v[`W-1]), _ABH1_v, n1267_v, _ABH1_i2, n1267_i2);
  spice_transistor_nmos g_1505((~cp1_v[`W-1]&~fetch_v[`W-1]), n1641_v, n119_v, n1641_i2, n119_i2);
  spice_transistor_nmos g_1502((~fetch_v[`W-1]&~cp1_v[`W-1]), n541_v, n1605_v, n541_i2, n1605_i3);
  spice_transistor_nmos g_1500((~ADH_ABH_v[`W-1]&~cp1_v[`W-1]), _ABH5_v, n254_v, _ABH5_i2, n254_i2);
  spice_transistor_nmos_gnd t551(~n1417_v[`W-1], clk1out_v, clk1out_i0);
  spice_transistor_nmos_gnd t2234(~n756_v[`W-1], n1110_v, n1110_i1);
  spice_transistor_nmos t2235(~dpc26_ACDB_v[`W-1], n146_v, idb0_v, n146_i1, idb0_i8);
  spice_transistor_nmos t2236(~dpc26_ACDB_v[`W-1], n929_v, idb1_v, n929_i2, idb1_i4);
  spice_transistor_nmos t2237(~dpc26_ACDB_v[`W-1], n1618_v, idb2_v, n1618_i0, idb2_i6);
  spice_transistor_nmos t1859(~dpc25_SBDB_v[`W-1], idb4_v, dasb4_v, idb4_i3, dasb4_i8);
  spice_transistor_nmos t1858(~dpc25_SBDB_v[`W-1], sb3_v, idb3_v, sb3_i7, idb3_i3);
  spice_transistor_nmos t1855(~dpc25_SBDB_v[`W-1], dasb0_v, idb0_v, dasb0_i6, idb0_i7);
  spice_transistor_nmos t1857(~dpc25_SBDB_v[`W-1], idb2_v, sb2_v, idb2_i5, sb2_i7);
  spice_transistor_nmos t1856(~dpc25_SBDB_v[`W-1], sb1_v, idb1_v, sb1_i7, idb1_i3);
  spice_transistor_nmos t2238(~dpc26_ACDB_v[`W-1], n1654_v, idb3_v, n1654_i2, idb3_i6);
  spice_transistor_nmos_gnd t1850(~n251_v[`W-1], RnWstretched_v, RnWstretched_i0);
  spice_transistor_nmos_gnd g_1182((~n755_v[`W-1]|~n781_v[`W-1]), n1170_v, n1170_i1);
  spice_transistor_nmos_gnd g_1183((~RnWstretched_v[`W-1]|~dor0_v[`W-1]), n769_v, n769_i2);
  spice_transistor_nmos t2728(~dpc9_DBADD_v[`W-1], alub5_v, idb5_v, alub5_i0, idb5_i7);
  spice_transistor_nmos t2729(~dpc9_DBADD_v[`W-1], alub4_v, idb4_v, alub4_i1, idb4_i7);
  spice_transistor_nmos_gnd g_1186((~n318_v[`W-1]|~_op_branch_bit7_v[`W-1]|~_op_branch_bit6_v[`W-1]), n1293_v, n1293_i2);
  spice_transistor_nmos_gnd g_1187((~brk_done_v[`W-1]|~n760_v[`W-1]), INTG_v, INTG_i2);
  spice_transistor_nmos_gnd g_1184((~n902_v[`W-1]|~n1464_v[`W-1]), n1109_v, n1109_i3);
  spice_transistor_nmos_gnd g_1185((~n761_v[`W-1]|~n149_v[`W-1]), n762_v, n762_i2);
  spice_transistor_nmos_gnd g_1188((~n1258_v[`W-1]|~op_ANDS_v[`W-1]|~n946_v[`W-1]|~n1412_v[`W-1]), n384_v, n384_i2);
  spice_transistor_nmos t2726(~dpc9_DBADD_v[`W-1], alub3_v, idb3_v, alub3_i1, idb3_i8);
  spice_transistor_nmos_gnd t2258(~pcl0_v[`W-1], n937_v, n937_i0);
  spice_transistor_nmos t2725(~dpc9_DBADD_v[`W-1], alub1_v, idb1_v, alub1_i1, idb1_i6);
  spice_transistor_nmos g_1451((~ADL_ABL_v[`W-1]&~cp1_v[`W-1]), _ABL0_v, n123_v, _ABL0_i2, n123_i2);
  spice_transistor_nmos_gnd t2621(~n1153_v[`W-1], n1639_v, n1639_i2);
  spice_transistor_nmos_gnd t429(~_ABH4_v[`W-1], abh4_v, abh4_i0);
  spice_transistor_nmos_gnd t422(~n135_v[`W-1], clk2out_v, clk2out_i1);
  spice_transistor_nmos t420(~cclk_v[`W-1], n1090_v, n1683_v, n1090_i0, n1683_i0);
  spice_transistor_nmos_gnd t421(~n762_v[`W-1], n1018_v, n1018_i0);
  spice_transistor_nmos_vdd t426(~cclk_v[`W-1], adh4_v, adh4_i2);
  spice_transistor_nmos_vdd t427(~cclk_v[`W-1], adl5_v, adl5_i0);
  spice_transistor_nmos t2656(~cclk_v[`W-1], pipe_T0_v, n17_v, pipe_T0_i0, n17_i2);
  spice_transistor_nmos_gnd t2653(~n1145_v[`W-1], op_ORS_v, op_ORS_i1);
  spice_transistor_nmos_vdd t2651(~dor0_v[`W-1], n1325_v, n1325_i1);
  spice_transistor_nmos t1079(~cp1_v[`W-1], _TWOCYCLE_v, _TWOCYCLE_phi1_v, _TWOCYCLE_i0, _TWOCYCLE_phi1_i0);
  spice_transistor_nmos_gnd t1078(~dpc12_0ADD_v[`W-1], alua0_v, alua0_i1);
  spice_transistor_nmos t1932(~cclk_v[`W-1], pclp5_v, n1073_v, pclp5_i1, n1073_i0);
  spice_transistor_nmos_gnd t2099(~_C78_v[`W-1], alurawcout_v, alurawcout_i1);
  spice_transistor_nmos t1453(~cclk_v[`W-1], n586_v, pipeUNK19_v, n586_i0, pipeUNK19_i0);
  spice_transistor_nmos t1452(~cclk_v[`W-1], n14_v, pipeUNK20_v, n14_i0, pipeUNK20_i0);
  spice_transistor_nmos_vdd t1679(~n42_v[`W-1], db3_v, db3_i1);
  spice_transistor_nmos t1678(~cclk_v[`W-1], n1037_v, n266_v, n1037_i0, n266_i0);
  spice_transistor_nmos t1677(~dpc41_DL_ADL_v[`W-1], adl5_v, n1387_v, adl5_i2, n1387_i2);
  spice_transistor_nmos t1676(~dpc41_DL_ADL_v[`W-1], adl6_v, n1014_v, adl6_i2, n1014_i2);
  spice_transistor_nmos_gnd g_1313((~RnWstretched_v[`W-1]|~dor5_v[`W-1]), n1720_v, n1720_i2);
  spice_transistor_nmos t1704(~cp1_v[`W-1], n1275_v, n1581_v, n1275_i0, n1581_i0);
  spice_transistor_nmos_gnd t1706(~ir1_v[`W-1], notir1_v, notir1_i0);
  spice_transistor_nmos_vdd t1701(~n475_v[`W-1], ab12_v, ab12_i1);
  spice_transistor_nmos_gnd t1700(~n1708_v[`W-1], n236_v, n236_i1);
  spice_transistor_nmos t1703(~cp1_v[`W-1], D1x1_v, n1472_v, D1x1_i0, n1472_i0);
  spice_transistor_nmos_gnd t1709(~n1399_v[`W-1], n1105_v, n1105_i2);
  spice_transistor_nmos_gnd g_1144((~op_T5_mem_ind_idx_v[`W-1]|~op_T3_mem_abs_v[`W-1]|~op_T4_mem_abs_idx_v[`W-1]|~op_T3_mem_zp_idx_v[`W-1]|~op_T2_mem_zp_v[`W-1]), n347_v, n347_i3);
  spice_transistor_nmos_gnd g_1145((~ir3_v[`W-1]|~ir2_v[`W-1]|~notir0_v[`W-1]|~t2_v[`W-1]), op_T2_ind_v, op_T2_ind_i1);
  spice_transistor_nmos_gnd t1927(~n1560_v[`W-1], n1081_v, n1081_i1);
  spice_transistor_nmos_gnd g_1142((~ir3_v[`W-1]|~ir7_v[`W-1]|~t2_v[`W-1]|~ir4_v[`W-1]|~ir6_v[`W-1]|~irline3_v[`W-1]|~ir2_v[`W-1]|~notir5_v[`W-1]), op_T2_jsr_v, op_T2_jsr_i3);
  spice_transistor_nmos_gnd g_1143((~n201_v[`W-1]|~n846_v[`W-1]|~n1045_v[`W-1]), n1371_v, n1371_i2);
  spice_transistor_nmos_gnd g_1364((~n644_v[`W-1]|~n1357_v[`W-1]), n678_v, n678_i3);
  spice_transistor_nmos_gnd t312(~n445_v[`W-1], sync_v, sync_i0);
  spice_transistor_nmos_gnd g_1140((~n460_v[`W-1]|~n43_v[`W-1]), n692_v, n692_i3);
  spice_transistor_nmos_gnd t317(~_ABH2_v[`W-1], abh2_v, abh2_i0);
  spice_transistor_nmos_gnd g_1141((~ir7_v[`W-1]|~notir6_v[`W-1]|~ir4_v[`W-1]|~irline3_v[`W-1]|~ir2_v[`W-1]|~ir3_v[`W-1]), op_rti_rts_v, op_rti_rts_i3);
  spice_transistor_nmos t2940(~cp1_v[`W-1], n666_v, n1380_v, n666_i1, n1380_i1);
  spice_transistor_nmos_gnd g_1361((~alub4_v[`W-1]|~alua4_v[`W-1]), n404_v, n404_i3);
  spice_transistor_nmos_gnd g_1365((~op_T__inx_v[`W-1]|~op_T__dex_v[`W-1]|~op_T0_ldx_tax_tsx_v[`W-1]), n844_v, n844_i2);
  spice_transistor_nmos t3119(~dpc2_XSB_v[`W-1], n242_v, sb3_v, n242_i2, sb3_i11);
  spice_transistor_nmos_gnd t3158(~notRdy0_v[`W-1], n1120_v, n1120_i0);
  spice_transistor_nmos_gnd g_1271((~notRdy0_v[`W-1]|~n959_v[`W-1]), n1154_v, n1154_i2);
  spice_transistor_nmos t684(~cclk_v[`W-1], pipeUNK32_v, n1081_v, pipeUNK32_i0, n1081_i0);
  spice_transistor_nmos t3358(~cclk_v[`W-1], n1199_v, notidl2_v, n1199_i1, notidl2_i1);
  spice_transistor_nmos_gnd t1920(~alu1_v[`W-1], _DA_ADD1_v, _DA_ADD1_i0);
  spice_transistor_nmos_gnd t228(~n621_v[`W-1], n355_v, n355_i0);
  spice_transistor_nmos_gnd g_1276((~alub5_v[`W-1]|~alua5_v[`W-1]), n1632_v, n1632_i4);
  spice_transistor_nmos_gnd t225(~n1061_v[`W-1], pchp3_v, pchp3_i0);
  spice_transistor_nmos t226(~dpc7_SS_v[`W-1], n332_v, s0_v, n332_i0, s0_i0);
  spice_transistor_nmos_vdd t227(~cclk_v[`W-1], idb0_v, idb0_i1);
  spice_transistor_nmos_gnd g_1312((~op_T2_php_v[`W-1]|~op_T4_brk_v[`W-1]), n1391_v, n1391_i2);
  spice_transistor_nmos t937(~dpc16_EORS_v[`W-1], notaluoutmux1_v, n953_v, notaluoutmux1_i0, n953_i0);
  spice_transistor_nmos t526(~dpc21_ADDADL_v[`W-1], alu7_v, adl7_v, alu7_i0, adl7_i0);
  spice_transistor_nmos t21(~cclk_v[`W-1], n983_v, nots0_v, n983_i0, nots0_i0);
  spice_transistor_nmos t20(~cclk_v[`W-1], n1162_v, n272_v, n1162_i0, n272_i0);
  spice_transistor_nmos_gnd t25(~abl0_v[`W-1], n1100_v, n1100_i0);
  spice_transistor_nmos t24(~cp1_v[`W-1], n1495_v, p3_v, n1495_i0, p3_i0);
  spice_transistor_nmos_vdd t27(~abl0_v[`W-1], n855_v, n855_i0);
  spice_transistor_nmos_gnd t26(~abl0_v[`W-1], n1660_v, n1660_i0);
  spice_transistor_nmos_gnd t524(~db5_v[`W-1], n568_v, n568_i1);
  spice_transistor_nmos t2504(~dpc8_nDBADD_v[`W-1], alub3_v, n1621_v, alub3_i0, n1621_i0);
  spice_transistor_nmos t523(~cclk_v[`W-1], n844_v, n459_v, n844_i0, n459_i0);
  spice_transistor_nmos_vdd t1922(~n1152_v[`W-1], ab2_v, ab2_i0);
  spice_transistor_nmos t522(~dpc21_ADDADL_v[`W-1], adl4_v, alu4_v, adl4_i1, alu4_i1);
  spice_transistor_nmos t521(~dpc21_ADDADL_v[`W-1], adl3_v, alu3_v, adl3_i0, alu3_i0);
  spice_transistor_nmos_gnd t2538(~idb6_v[`W-1], n1416_v, n1416_i0);
  spice_transistor_nmos_gnd t2537(~n_0_ADL2_v[`W-1], adl2_v, adl2_i6);
  spice_transistor_nmos t2535(~cclk_v[`W-1], n635_v, _ABH6_v, n635_i3, _ABH6_i1);
  spice_transistor_nmos t520(~cp1_v[`W-1], n87_v, idl1_v, n87_i1, idl1_i0);
  spice_transistor_nmos_gnd t2508(~pipeUNK02_v[`W-1], n1492_v, n1492_i0);
  spice_transistor_nmos t2531(~dpc38_PCLADL_v[`W-1], adl2_v, n481_v, adl2_i5, n481_i2);
  spice_transistor_nmos t2530(~dpc38_PCLADL_v[`W-1], n976_v, adl1_v, n976_i0, adl1_i5);
  spice_transistor_nmos_gnd g_1060((~n491_v[`W-1]|~cclk_v[`W-1]|~n1247_v[`W-1]), dpc10_ADLADD_v, dpc10_ADLADD_i9);
  spice_transistor_nmos_vdd t130(~n1369_v[`W-1], dpc38_PCLADL_v, dpc38_PCLADL_i0);
  spice_transistor_nmos t132(~dpc4_SSB_v[`W-1], n721_v, sb7_v, n721_i0, sb7_i0);
  spice_transistor_nmos t133(~dpc4_SSB_v[`W-1], n618_v, sb6_v, n618_i0, sb6_i2);
  spice_transistor_nmos_gnd t134(~n818_v[`W-1], n1043_v, n1043_i0);
  spice_transistor_nmos_vdd t135(~n818_v[`W-1], dpc40_ADLPCL_v, dpc40_ADLPCL_i0);
  spice_transistor_nmos t136(~dpc4_SSB_v[`W-1], n3_v, dasb4_v, n3_i0, dasb4_i3);
  spice_transistor_nmos g_1463((~cp1_v[`W-1]&~ADL_ABL_v[`W-1]), n1016_v, _ABL1_v, n1016_i2, _ABL1_i2);
  spice_transistor_nmos_gnd g_1464((~alua5_v[`W-1]&~alub5_v[`W-1]), n477_v, n477_i4);
  spice_transistor_nmos_gnd g_1468((~alub7_v[`W-1]&~alua7_v[`W-1]), n1318_v, n1318_i5);
  spice_transistor_nmos_gnd t2890(~pchp1_v[`W-1], n209_v, n209_i2);
  spice_transistor_nmos t2891(~cp1_v[`W-1], notRnWprepad_v, n759_v, notRnWprepad_i2, n759_i0);
  spice_transistor_nmos_gnd g_1317((~x_op_push_pull_v[`W-1]|~notir3_v[`W-1]|~ir2_v[`W-1]|~ir0_v[`W-1]), op_implied_v, op_implied_i2);
  spice_transistor_nmos_gnd t2892(~idb0_v[`W-1], n1687_v, n1687_i1);
  spice_transistor_nmos t3130(~cclk_v[`W-1], n1391_v, pipeUNK15_v, n1391_i0, pipeUNK15_i1);
  spice_transistor_nmos_gnd t3131(~n531_v[`W-1], n1255_v, n1255_i1);
  spice_transistor_nmos t3134(~cclk_v[`W-1], _ABH4_v, n999_v, _ABH4_i1, n999_i3);
  spice_transistor_nmos t3136(~cclk_v[`W-1], n1106_v, n1404_v, n1106_i0, n1404_i0);
  spice_transistor_nmos_gnd t3137(~notidl5_v[`W-1], idl5_v, idl5_i1);
  spice_transistor_nmos_gnd g_1267((~cclk_v[`W-1]|~n255_v[`W-1]|~n1247_v[`W-1]), dpc31_PCHPCH_v, dpc31_PCHPCH_i9);
  spice_transistor_nmos_gnd g_1266((~ir4_v[`W-1]|~irline3_v[`W-1]|~t3_v[`W-1]|~ir7_v[`W-1]), op_T3_stack_bit_jmp_v, op_T3_stack_bit_jmp_i1);
  spice_transistor_nmos_gnd g_1265((~ir7_v[`W-1]|~ir4_v[`W-1]|~ir2_v[`W-1]|~notir3_v[`W-1]|~notir5_v[`W-1]|~t3_v[`W-1]|~irline3_v[`W-1]), op_T3_plp_pla_v, op_T3_plp_pla_i2);
  spice_transistor_nmos_gnd g_1264((~RnWstretched_v[`W-1]|~dor5_v[`W-1]), n612_v, n612_i2);
  spice_transistor_nmos_gnd g_1263((~cclk_v[`W-1]|~n1247_v[`W-1]|~n282_v[`W-1]), dpc6_SBS_v, dpc6_SBS_i9);
  spice_transistor_nmos_gnd t2896(~pipeUNK12_v[`W-1], n587_v, n587_i0);
  spice_transistor_nmos_gnd g_1261((~cclk_v[`W-1]|~n708_v[`W-1]|~n1247_v[`W-1]), dpc11_SBADD_v, dpc11_SBADD_i9);
  spice_transistor_nmos_gnd g_1260((~notir3_v[`W-1]|~ir7_v[`W-1]|~ir4_v[`W-1]|~ir2_v[`W-1]|~notir1_v[`W-1]|~clock2_v[`W-1]), op_T__shift_a_v, op_T__shift_a_i2);
  spice_transistor_nmos t2897(~dpc20_ADDSB06_v[`W-1], alu0_v, dasb0_v, alu0_i2, dasb0_i11);
  spice_transistor_nmos_gnd g_1269((~cp1_v[`W-1]|~n519_v[`W-1]), n127_v, n127_i3);
  spice_transistor_nmos_gnd g_1268((~C1x5Reset_v[`W-1]|~INTG_v[`W-1]), D1x1_v, D1x1_i3);
  spice_transistor_nmos t2895(~dpc20_ADDSB06_v[`W-1], alu1_v, sb1_v, alu1_i3, sb1_i10);
  spice_transistor_nmos t549(~cclk_v[`W-1], n1071_v, notalu3_v, n1071_i1, notalu3_i0);
  spice_transistor_nmos g_1518((~cp1_v[`W-1]&~ADL_ABL_v[`W-1]), n935_v, _ABL2_v, n935_i2, _ABL2_i2);
  spice_transistor_nmos_gnd g_1049((~notir7_v[`W-1]|~notir6_v[`W-1]|~notir0_v[`W-1]|~notir5_v[`W-1]|~clock1_v[`W-1]), op_T0_sbc_v, op_T0_sbc_i1);
  spice_transistor_nmos_gnd g_1048((~notir0_v[`W-1]|~notir6_v[`W-1]|~clock1_v[`W-1]|~notir5_v[`W-1]), op_T0_adc_sbc_v, op_T0_adc_sbc_i1);
  spice_transistor_nmos g_1515((~ADH_ABH_v[`W-1]&~cp1_v[`W-1]), _ABH2_v, n168_v, _ABH2_i2, n168_i2);
  spice_transistor_nmos_gnd t540(~n1635_v[`W-1], dpc29_0ADH17_v, dpc29_0ADH17_i1);
  spice_transistor_nmos_gnd g_1517((~Pout3_v[`W-1]&~op_T0_sbc_v[`W-1]), n29_v, n29_i2);
  spice_transistor_nmos g_1516((~fetch_v[`W-1]&~cp1_v[`W-1]), n1300_v, n571_v, n1300_i2, n571_i2);
  spice_transistor_nmos t546(~dpc13_ORS_v[`W-1], n649_v, n1071_v, n649_i0, n1071_i0);
  spice_transistor_nmos t2241(~dpc26_ACDB_v[`W-1], n326_v, idb6_v, n326_i2, idb6_i6);
  spice_transistor_nmos t2240(~dpc26_ACDB_v[`W-1], n831_v, idb5_v, n831_i1, idb5_i4);
  spice_transistor_nmos t2242(~dpc26_ACDB_v[`W-1], n1592_v, idb7_v, n1592_i2, idb7_i6);
  spice_transistor_nmos t1848(~dpc23_SBAC_v[`W-1], dasb7_v, a7_v, dasb7_i0, a7_i2);
  spice_transistor_nmos_gnd t1849(~n251_v[`W-1], n1028_v, n1028_i0);
  spice_transistor_nmos t1846(~dpc23_SBAC_v[`W-1], dasb5_v, a5_v, dasb5_i0, a5_i2);
  spice_transistor_nmos t1847(~dpc23_SBAC_v[`W-1], dasb6_v, a6_v, dasb6_i0, a6_i2);
  spice_transistor_nmos t1844(~dpc23_SBAC_v[`W-1], dasb3_v, a3_v, dasb3_i0, a3_i1);
  spice_transistor_nmos t1845(~dpc23_SBAC_v[`W-1], dasb4_v, a4_v, dasb4_i7, a4_i0);
  spice_transistor_nmos t1842(~dpc23_SBAC_v[`W-1], dasb1_v, a1_v, dasb1_i0, a1_i1);
  spice_transistor_nmos t1843(~dpc23_SBAC_v[`W-1], a2_v, dasb2_v, a2_i1, dasb2_i0);
  spice_transistor_nmos t1841(~dpc23_SBAC_v[`W-1], dasb0_v, a0_v, dasb0_i5, a0_i1);
  spice_transistor_nmos_gnd t2086(~a4_v[`W-1], n556_v, n556_i0);
  spice_transistor_nmos t2085(~cclk_v[`W-1], n1194_v, pipeUNK04_v, n1194_i1, pipeUNK04_i0);
  spice_transistor_nmos_gnd t2084(~n646_v[`W-1], n470_v, n470_i0);
  spice_transistor_nmos_gnd g_1195((~op_T2_zp_zp_idx_v[`W-1]|~op_T2_ind_v[`W-1]), n1225_v, n1225_i4);
  spice_transistor_nmos t2082(~cclk_v[`W-1], pipeUNK30_v, n385_v, pipeUNK30_i0, n385_i0);
  spice_transistor_nmos_gnd g_1199((~n61_v[`W-1]|~n739_v[`W-1]), n479_v, n479_i1);
  spice_transistor_nmos_gnd g_1198((~n862_v[`W-1]|~op_T5_rts_v[`W-1]|~nnT2BR_v[`W-1]|~n646_v[`W-1]|~n236_v[`W-1]|~op_T2_abs_access_v[`W-1]), n272_v, n272_i3);
  spice_transistor_nmos_gnd t2089(~n1121_v[`W-1], n291_v, n291_i2);
  spice_transistor_nmos_gnd t1280(~pd5_clearIR_v[`W-1], n928_v, n928_i0);
  spice_transistor_nmos_gnd t1282(~pch1_v[`W-1], n1070_v, n1070_i0);
  spice_transistor_nmos_vdd t435(~n1523_v[`W-1], n635_v, n635_i0);
  spice_transistor_nmos_gnd t434(~n1523_v[`W-1], n963_v, n963_i1);
  spice_transistor_nmos_vdd t437(~n1260_v[`W-1], dpc32_PCHADH_v, dpc32_PCHADH_i1);
  spice_transistor_nmos_gnd t436(~n1260_v[`W-1], n1413_v, n1413_i1);
  spice_transistor_nmos t431(~cclk_v[`W-1], n474_v, n15_v, n474_i0, n15_i0);
  spice_transistor_nmos t432(~dpc2_XSB_v[`W-1], n1169_v, dasb0_v, n1169_i0, dasb0_i2);
  spice_transistor_nmos_vdd t439(~n220_v[`W-1], ADL_ABL_v, ADL_ABL_i0);
  spice_transistor_nmos_gnd t438(~n220_v[`W-1], n130_v, n130_i0);
  spice_transistor_nmos t941(~dpc16_EORS_v[`W-1], n1469_v, n277_v, n1469_i0, n277_i1);
  spice_transistor_nmos t940(~dpc16_EORS_v[`W-1], __AxB_4_v, n296_v, __AxB_4_i0, n296_i0);
  spice_transistor_nmos t943(~dpc16_EORS_v[`W-1], n304_v, n177_v, n304_i1, n177_i1);
  spice_transistor_nmos t942(~dpc16_EORS_v[`W-1], __AxB_6_v, n722_v, __AxB_6_i1, n722_i1);
  spice_transistor_nmos_gnd g_1649((~n1691_v[`W-1]|(~n681_v[`W-1]&~_C12_v[`W-1])), C23_v, C23_i2);
  spice_transistor_nmos_gnd t2667(~db6_v[`W-1], n1638_v, n1638_i1);
  spice_transistor_nmos_gnd t2669(~n206_v[`W-1], n465_v, n465_i0);
  spice_transistor_nmos t2883(~n771_v[`W-1], n430_v, n465_v, n430_i3, n465_i1);
  spice_transistor_nmos_gnd t2881(~n745_v[`W-1], n241_v, n241_i2);
  spice_transistor_nmos t2864(~cclk_v[`W-1], n1575_v, pipeT2out_v, n1575_i1, pipeT2out_i0);
  spice_transistor_nmos_gnd t2867(~x4_v[`W-1], n485_v, n485_i1);
  spice_transistor_nmos t2259(~cclk_v[`W-1], n1500_v, n526_v, n1500_i0, n526_i1);
  spice_transistor_nmos_gnd t2869(~notdor4_v[`W-1], dor4_v, dor4_i1);
  spice_transistor_nmos_gnd t1448(~op_implied_v[`W-1], n664_v, n664_i1);
  spice_transistor_nmos t1449(~cp1_v[`W-1], n675_v, n330_v, n675_i1, n330_i0);
  spice_transistor_nmos_gnd g_1219((~op_T0_jsr_v[`W-1]|~op_T0_php_pha_v[`W-1]|~op_T5_rti_v[`W-1]|~op_T5_brk_v[`W-1]|~op_T4_rts_v[`W-1]|~op_T3_plp_pla_v[`W-1]), n1464_v, n1464_i2);
  spice_transistor_nmos t1716(~cp1_v[`W-1], n50_v, INTG_v, n50_i0, INTG_i0);
  spice_transistor_nmos_vdd t1712(~n1325_v[`W-1], db0_v, db0_i1);
  spice_transistor_nmos_gnd t1718(~op_branch_done_v[`W-1], _op_branch_done_v, _op_branch_done_i0);
  spice_transistor_nmos_gnd t2437(~n1696_v[`W-1], rw_v, rw_i1);
  spice_transistor_nmos_gnd g_1118((~op_T5_rti_v[`W-1]|~op_T3_v[`W-1]|~op_T4_v[`W-1]|~op_T0_jmp_v[`W-1]|~op_T0_brk_rti_v[`W-1]|~op_T5_ind_x_v[`W-1]|~op_T5_rts_v[`W-1]), n256_v, n256_i1);
  spice_transistor_nmos_gnd t3127(~n1599_v[`W-1], n538_v, n538_i0);
  spice_transistor_nmos_gnd t301(~n612_v[`W-1], db5_v, db5_i0);
  spice_transistor_nmos_gnd t300(~n730_v[`W-1], n1724_v, n1724_i0);
  spice_transistor_nmos_gnd t1479(~op_T0_clc_sec_v[`W-1], n889_v, n889_i1);
  spice_transistor_nmos_gnd t309(~n445_v[`W-1], n417_v, n417_i0);
  spice_transistor_nmos_gnd t308(~n445_v[`W-1], n317_v, n317_i0);
  spice_transistor_nmos_vdd t1477(~n17_v[`W-1], clock1_v, clock1_i1);
  spice_transistor_nmos t1476(~cclk_v[`W-1], n676_v, _ABH1_v, n676_i0, _ABH1_i0);
  spice_transistor_nmos_gnd t1472(~n339_v[`W-1], n543_v, n543_i0);
  spice_transistor_nmos g_1506((~cp1_v[`W-1]&~fetch_v[`W-1]), n409_v, n310_v, n409_i3, n310_i2);
  spice_transistor_nmos_vdd t1471(~n91_v[`W-1], dpc15_ANDS_v, dpc15_ANDS_i0);
  spice_transistor_nmos_gnd t1470(~n91_v[`W-1], n1256_v, n1256_i0);
  spice_transistor_nmos_gnd t2143(~n108_v[`W-1], dpc16_EORS_v, dpc16_EORS_i8);
  spice_transistor_nmos_gnd t1656(~n126_v[`W-1], pchp1_v, pchp1_i0);
  spice_transistor_nmos_gnd t239(~op_T5_brk_v[`W-1], n689_v, n689_i0);
  spice_transistor_nmos t238(~dpc42_DL_ADH_v[`W-1], adh7_v, n1147_v, adh7_i0, n1147_i0);
  spice_transistor_nmos t237(~dpc42_DL_ADH_v[`W-1], adh6_v, n1014_v, adh6_i0, n1014_i0);
  spice_transistor_nmos t236(~dpc42_DL_ADH_v[`W-1], adh5_v, n1387_v, adh5_i0, n1387_i0);
  spice_transistor_nmos t235(~dpc42_DL_ADH_v[`W-1], adh4_v, n1095_v, adh4_i0, n1095_i0);
  spice_transistor_nmos t234(~dpc42_DL_ADH_v[`W-1], adh3_v, n1661_v, adh3_i0, n1661_i0);
  spice_transistor_nmos t233(~dpc42_DL_ADH_v[`W-1], adh2_v, n1424_v, adh2_i0, n1424_i1);
  spice_transistor_nmos t232(~dpc42_DL_ADH_v[`W-1], adh1_v, n87_v, adh1_i0, n87_i0);
  spice_transistor_nmos t231(~dpc42_DL_ADH_v[`W-1], adh0_v, n719_v, adh0_i0, n719_i0);
  spice_transistor_nmos_gnd g_1119((~ir2_v[`W-1]|~ir7_v[`W-1]|~t4_v[`W-1]|~ir4_v[`W-1]|~ir3_v[`W-1]|~ir6_v[`W-1]|~irline3_v[`W-1]), op_T4_brk_jsr_v, op_T4_brk_jsr_i1);
  spice_transistor_nmos_gnd t1651(~n95_v[`W-1], n531_v, n531_i0);
  spice_transistor_nmos_gnd g_1370((~n344_v[`W-1]|~n232_v[`W-1]), n1316_v, n1316_i1);
  spice_transistor_nmos_gnd t1650(~n987_v[`W-1], n1169_v, n1169_i1);
  spice_transistor_nmos_gnd g_1373((~ir5_v[`W-1]|~notir7_v[`W-1]|~ir6_v[`W-1]), op_store_v, op_store_i2);
  spice_transistor_nmos_vdd t36(~cclk_v[`W-1], dasb4_v, dasb4_i0);
  spice_transistor_nmos t37(~cclk_v[`W-1], n973_v, nots4_v, n973_i0, nots4_i0);
  spice_transistor_nmos t34(~cclk_v[`W-1], n518_v, y6_v, n518_i0, y6_i0);
  spice_transistor_nmos_gnd t35(~p0_v[`W-1], n31_v, n31_i0);
  spice_transistor_nmos_gnd g_1374((~n345_v[`W-1]|~n432_v[`W-1]), n1097_v, n1097_i1);
  spice_transistor_nmos_gnd g_1376((~alua7_v[`W-1]|~alub7_v[`W-1]), n1398_v, n1398_i4);
  spice_transistor_nmos t2528(~dpc38_PCLADL_v[`W-1], n1647_v, adl7_v, n1647_i1, adl7_i5);
  spice_transistor_nmos t2529(~dpc38_PCLADL_v[`W-1], adl0_v, n488_v, adl0_i5, n488_i2);
  spice_transistor_nmos_gnd g_1378((~RnWstretched_v[`W-1]|~dor4_v[`W-1]), n147_v, n147_i2);
  spice_transistor_nmos_gnd t2521(~notRdy0_v[`W-1], n1718_v, n1718_i1);
  spice_transistor_nmos_gnd t2522(~op_T0_eor_v[`W-1], n837_v, n837_i0);
  spice_transistor_nmos_vdd t2523(~n747_v[`W-1], clk1out_v, clk1out_i1);
  spice_transistor_nmos_gnd t2524(~n358_v[`W-1], n1715_v, n1715_i2);
  spice_transistor_nmos t2525(~dpc38_PCLADL_v[`W-1], adl4_v, n208_v, adl4_i5, n208_i2);
  spice_transistor_nmos t2526(~dpc38_PCLADL_v[`W-1], n72_v, adl5_v, n72_i2, adl5_i4);
  spice_transistor_nmos t2527(~dpc38_PCLADL_v[`W-1], adl6_v, n1458_v, adl6_i4, n1458_i1);
  spice_transistor_nmos_gnd t129(~n1369_v[`W-1], n1462_v, n1462_i0);
  spice_transistor_nmos t128(~dpc4_SSB_v[`W-1], n1389_v, sb2_v, n1389_i0, sb2_i1);
  spice_transistor_nmos t2629(~cclk_v[`W-1], pipeUNK09_v, n327_v, pipeUNK09_i0, n327_i0);
  spice_transistor_nmos_gnd t121(~pclp7_v[`W-1], n1647_v, n1647_i0);
  spice_transistor_nmos t127(~dpc4_SSB_v[`W-1], n998_v, sb3_v, n998_i0, sb3_i1);
  spice_transistor_nmos t126(~cclk_v[`W-1], n1179_v, n393_v, n1179_i0, n393_i0);
  spice_transistor_nmos t125(~cp1_v[`W-1], n430_v, n1570_v, n430_i0, n1570_i0);
  spice_transistor_nmos_gnd t124(~DBZ_v[`W-1], _DBZ_v, _DBZ_i0);
  spice_transistor_nmos_gnd g_1644(((~op_T0_acc_v[`W-1]&~n397_v[`W-1])|(~op_T0_tay_v[`W-1]|~op_ANDS_v[`W-1]|~op_T0_tax_v[`W-1]|~op_T0_shift_a_v[`W-1])), n11_v, n11_i2);
  spice_transistor_nmos g_1459((~cp1_v[`W-1]&~fetch_v[`W-1]), n227_v, n927_v, n227_i2, n927_i2);
  spice_transistor_nmos_gnd g_1328((~dor6_v[`W-1]|~RnWstretched_v[`W-1]), n471_v, n471_i2);
  spice_transistor_nmos_gnd g_1329((~_op_branch_bit6_v[`W-1]|~n90_v[`W-1]|~n201_v[`W-1]), n1433_v, n1433_i2);
  spice_transistor_nmos_gnd g_1326((~alub0_v[`W-1]|~alua0_v[`W-1]), aluanorb0_v, aluanorb0_i3);
  spice_transistor_nmos_gnd g_1327((~n43_v[`W-1]|~n688_v[`W-1]), n1223_v, n1223_i3);
  spice_transistor_nmos_gnd g_1322((~n1010_v[`W-1]|~n1007_v[`W-1]|~n923_v[`W-1]|~n1070_v[`W-1]|~n1265_v[`W-1]), dpc35_PCHC_v, dpc35_PCHC_i1);
  spice_transistor_nmos_gnd g_1323((~n796_v[`W-1]|~n43_v[`W-1]), n35_v, n35_i3);
  spice_transistor_nmos_gnd g_1320((~op_T2_abs_access_v[`W-1]|~n646_v[`W-1]), n773_v, n773_i1);
  spice_transistor_nmos_gnd g_1321((~n620_v[`W-1]|~n270_v[`W-1]), n1115_v, n1115_i1);
  spice_transistor_nmos_gnd t3383(~res_v[`W-1], n312_v, n312_i1);
  spice_transistor_nmos_gnd t3382(~n1271_v[`W-1], dpc27_SBADH_v, dpc27_SBADH_i9);
  spice_transistor_nmos_gnd g_1210((~AxB3_v[`W-1]|~_C23_v[`W-1]), __AxB3__C23_v, __AxB3__C23_i1);
  spice_transistor_nmos_gnd g_1211((~pipe_T0_v[`W-1]|~notRdy0_v[`W-1]), n1180_v, n1180_i2);
  spice_transistor_nmos_gnd g_1216((~n1448_v[`W-1]|~n182_v[`W-1]), n1619_v, n1619_i1);
  spice_transistor_nmos_gnd g_1217((~irline3_v[`W-1]|~notir7_v[`W-1]|~ir4_v[`W-1]|~ir3_v[`W-1]|~notir6_v[`W-1]|~clock2_v[`W-1]), op_T__cpx_cpy_imm_zp_v, op_T__cpx_cpy_imm_zp_i1);
  spice_transistor_nmos t3384(~dpc20_ADDSB06_v[`W-1], alu2_v, sb2_v, alu2_i3, sb2_i11);
  spice_transistor_nmos_gnd t3435(~sb3_v[`W-1], n432_v, n432_i0);
  spice_transistor_nmos_vdd t3434(~n1270_v[`W-1], dpc39_PCLPCL_v, dpc39_PCLPCL_i8);
  spice_transistor_nmos t3389(~cclk_v[`W-1], n1341_v, n695_v, n1341_i1, n695_i0);
  spice_transistor_nmos_gnd t3388(~nots6_v[`W-1], n618_v, n618_i3);
  spice_transistor_nmos_gnd t3433(~n1270_v[`W-1], n1518_v, n1518_i0);
  spice_transistor_nmos_gnd g_1528((~n616_v[`W-1]&~n844_v[`W-1]), n946_v, n946_i2);
  spice_transistor_nmos_gnd g_1038((~notir3_v[`W-1]|~ir2_v[`W-1]|~ir4_v[`W-1]|~clock1_v[`W-1]|~notir1_v[`W-1]|~ir5_v[`W-1]|~ir6_v[`W-1]|~notir7_v[`W-1]), op_T0_txa_v, op_T0_txa_i1);
  spice_transistor_nmos_gnd g_1039((~notir3_v[`W-1]|~notir4_v[`W-1]|~ir2_v[`W-1]|~clock1_v[`W-1]|~ir5_v[`W-1]|~irline3_v[`W-1]|~ir6_v[`W-1]|~notir7_v[`W-1]), op_T0_tya_v, op_T0_tya_i1);
  spice_transistor_nmos t2935(~cp1_v[`W-1], n47_v, n420_v, n47_i1, n420_i0);
  spice_transistor_nmos_gnd g_1032((~n265_v[`W-1]|~n43_v[`W-1]), n818_v, n818_i3);
  spice_transistor_nmos_gnd g_1033((~n937_v[`W-1]|~dpc36_IPC_v[`W-1]), n1345_v, n1345_i1);
  spice_transistor_nmos_gnd g_1031((~n819_v[`W-1]|~n1154_v[`W-1]), n1380_v, n1380_i3);
  spice_transistor_nmos_gnd g_1036((~n862_v[`W-1]|~n1258_v[`W-1]|~n192_v[`W-1]|~n1002_v[`W-1]|~n1109_v[`W-1]), n1130_v, n1130_i2);
  spice_transistor_nmos_gnd g_1037((~dor0_v[`W-1]|~RnWstretched_v[`W-1]), n1072_v, n1072_i2);
  spice_transistor_nmos_gnd g_1034((~ir6_v[`W-1]|~irline3_v[`W-1]|~ir2_v[`W-1]|~notir3_v[`W-1]|~notir4_v[`W-1]|~notir5_v[`W-1]|~notir7_v[`W-1]), op_clv_v, op_clv_i2);
  spice_transistor_nmos_gnd t2252(~abh2_v[`W-1], n994_v, n994_i1);
  spice_transistor_nmos_gnd t1879(~n1295_v[`W-1], n1238_v, n1238_i1);
  spice_transistor_nmos_gnd t2256(~n610_v[`W-1], n582_v, n582_i2);
  spice_transistor_nmos t2257(~dpc0_YSB_v[`W-1], n1251_v, sb7_v, n1251_i1, sb7_i8);
  spice_transistor_nmos t2254(~dpc27_SBADH_v[`W-1], sb1_v, adh1_v, sb1_i8, adh1_i4);
  spice_transistor_nmos_gnd t1873(~op_T0_cld_sed_v[`W-1], n774_v, n774_i0);
  spice_transistor_nmos_gnd t1870(~_ABL3_v[`W-1], abl3_v, abl3_i3);
  spice_transistor_nmos t1876(~dpc41_DL_ADL_v[`W-1], n1147_v, adl7_v, n1147_i2, adl7_i3);
  spice_transistor_nmos_gnd t1875(~notdor6_v[`W-1], dor6_v, dor6_i0);
  spice_transistor_nmos_gnd t1874(~n390_v[`W-1], n1258_v, n1258_i0);
  spice_transistor_nmos_gnd t2090(~n981_v[`W-1], n733_v, n733_i0);
  spice_transistor_nmos t2091(~cclk_v[`W-1], _ABL1_v, n66_v, _ABL1_i1, n66_i2);
  spice_transistor_nmos_vdd t2092(~abh4_v[`W-1], n475_v, n475_i2);
  spice_transistor_nmos_gnd t1917(~n663_v[`W-1], pchp7_v, pchp7_i0);
  spice_transistor_nmos_gnd t2094(~abh4_v[`W-1], n999_v, n999_i2);
  spice_transistor_nmos t2095(~cclk_v[`W-1], notaluoutmux0_v, notalu0_v, notaluoutmux0_i4, notalu0_i1);
  spice_transistor_nmos_gnd t2096(~C01_v[`W-1], _C01_v, _C01_i0);
  spice_transistor_nmos_gnd t2098(~n1447_v[`W-1], n1175_v, n1175_i0);
  spice_transistor_nmos_vdd t1911(~cclk_v[`W-1], adh2_v, adh2_i3);
  spice_transistor_nmos t1279(~cclk_v[`W-1], n296_v, notalu4_v, n296_i2, notalu4_i1);
  spice_transistor_nmos_gnd t1274(~n1010_v[`W-1], n311_v, n311_i0);
  spice_transistor_nmos t1271(~cclk_v[`W-1], n340_v, pipeUNK12_v, n340_i1, pipeUNK12_i0);
  spice_transistor_nmos t1273(~n1446_v[`W-1], n430_v, n206_v, n430_i1, n206_i1);
  spice_transistor_nmos_gnd t440(~n400_v[`W-1], n102_v, n102_i0);
  spice_transistor_nmos_vdd t441(~n400_v[`W-1], n1696_v, n1696_i0);
  spice_transistor_nmos_gnd t442(~n834_v[`W-1], n1696_v, n1696_i1);
  spice_transistor_nmos_gnd t443(~n834_v[`W-1], n400_v, n400_i2);
  spice_transistor_nmos_gnd t444(~x7_v[`W-1], n1561_v, n1561_i0);
  spice_transistor_nmos_vdd t446(~n1545_v[`W-1], ab10_v, ab10_i0);
  spice_transistor_nmos_gnd g_1148((~ir2_v[`W-1]|~notir4_v[`W-1]|~notir0_v[`W-1]|~ir3_v[`W-1]|~t5_v[`W-1]), op_T5_ind_y_v, op_T5_ind_y_i1);
  spice_transistor_nmos_gnd g_1149((~clock1_v[`W-1]|~notir0_v[`W-1]), op_T0_acc_v, op_T0_acc_i1);
  spice_transistor_nmos_gnd t932(~alu2_v[`W-1], _DA_ADD2_v, _DA_ADD2_i0);
  spice_transistor_nmos_gnd t934(~n1593_v[`W-1], n1552_v, n1552_i0);
  spice_transistor_nmos_vdd t935(~n1593_v[`W-1], dpc14_SRS_v, dpc14_SRS_i1);
  spice_transistor_nmos t936(~dpc16_EORS_v[`W-1], __AxB_0_v, notaluoutmux0_v, __AxB_0_i0, notaluoutmux0_i0);
  spice_transistor_nmos t681(~cclk_v[`W-1], n473_v, pipeUNK33_v, n473_i0, pipeUNK33_i0);
  spice_transistor_nmos t938(~dpc16_EORS_v[`W-1], __AxB_2_v, n740_v, __AxB_2_i0, n740_i1);
  spice_transistor_nmos t939(~dpc16_EORS_v[`W-1], n884_v, n1071_v, n884_i1, n1071_i2);
  spice_transistor_nmos_gnd t2678(~cp1_v[`W-1], n43_v, n43_i1);
  spice_transistor_nmos_gnd t2674(~abl5_v[`W-1], n210_v, n210_i3);
  spice_transistor_nmos_gnd t2675(~abl5_v[`W-1], n172_v, n172_i2);
  spice_transistor_nmos_vdd t2676(~abl5_v[`W-1], n1633_v, n1633_i2);
  spice_transistor_nmos_gnd t2677(~n419_v[`W-1], n1618_v, n1618_i2);
  spice_transistor_nmos_gnd t1011(~n25_v[`W-1], n674_v, n674_i0);
  spice_transistor_nmos t1010(~cclk_v[`W-1], n1675_v, notir6_v, n1675_i0, notir6_i1);
  spice_transistor_nmos t1013(~cclk_v[`W-1], pd3_v, n1281_v, pd3_i0, n1281_i1);
  spice_transistor_nmos t1012(~cclk_v[`W-1], n1588_v, pd5_v, n1588_i0, pd5_i0);
  spice_transistor_nmos t1015(~cclk_v[`W-1], n929_v, a1_v, n929_i0, a1_i0);
  spice_transistor_nmos t1014(~cclk_v[`W-1], pd4_v, n1075_v, pd4_i0, n1075_i0);
  spice_transistor_nmos t1017(~cclk_v[`W-1], n1638_v, notidl6_v, n1638_i0, notidl6_i1);
  spice_transistor_nmos_gnd t1388(~notalu0_v[`W-1], alu0_v, alu0_i1);
  spice_transistor_nmos_vdd t2873(~n1315_v[`W-1], n381_v, n381_i3);
  spice_transistor_nmos_gnd t2871(~notdor3_v[`W-1], dor3_v, dor3_i1);
  spice_transistor_nmos_gnd t1385(~n1356_v[`W-1], n326_v, n326_i1);
  spice_transistor_nmos t1384(~dpc37_PCLDB_v[`W-1], n1458_v, idb6_v, n1458_i0, idb6_i2);
  spice_transistor_nmos t592(~dpc43_DL_DB_v[`W-1], idb7_v, n1147_v, idb7_i2, n1147_i1);
  spice_transistor_nmos t590(~dpc43_DL_DB_v[`W-1], idb5_v, n1387_v, idb5_i1, n1387_i1);
  spice_transistor_nmos t591(~dpc43_DL_DB_v[`W-1], idb6_v, n1014_v, idb6_i0, n1014_i1);
  spice_transistor_nmos_vdd t594(~n322_v[`W-1], ab7_v, ab7_i0);
  spice_transistor_nmos_gnd t1478(~n17_v[`W-1], n646_v, n646_i0);
  spice_transistor_nmos t1125(~cclk_v[`W-1], n442_v, n509_v, n442_i1, n509_i0);
  spice_transistor_nmos_gnd t1126(~n1025_v[`W-1], n564_v, n564_i1);
  spice_transistor_nmos t1121(~cp1_v[`W-1], n1339_v, n597_v, n1339_i0, n597_i0);
  spice_transistor_nmos_gnd t1120(~pclp5_v[`W-1], n72_v, n72_i0);
  spice_transistor_nmos_gnd t1123(~n485_v[`W-1], n436_v, n436_i0);
  spice_transistor_nmos_gnd t1122(~n402_v[`W-1], n834_v, n834_i2);
  spice_transistor_nmos_gnd t1496(~n1105_v[`W-1], cp1_v, cp1_i35);
  spice_transistor_nmos_gnd g_1658(((~A_B3_v[`W-1]&~C23_v[`W-1])|(~DC34_v[`W-1]|~n988_v[`W-1])), _C34_v, _C34_i3);
  spice_transistor_nmos t1493(~cclk_v[`W-1], pipe_VEC_v, _VEC_v, pipe_VEC_i0, _VEC_i0);
  spice_transistor_nmos_gnd g_1180((~notir4_v[`W-1]|~ir3_v[`W-1]|~n603_v[`W-1]|~ir2_v[`W-1]|~irline3_v[`W-1]|~clock1_v[`W-1]), op_branch_done_v, op_branch_done_i2);
  spice_transistor_nmos_gnd g_1659(((~op_from_x_v[`W-1]&~n335_v[`W-1])|(~op_T2_idx_x_xy_v[`W-1]&~n1244_v[`W-1])|(~op_T2_ind_x_v[`W-1]|~op_T0_dex_v[`W-1]|~op_T0_cpx_inx_v[`W-1]|~x_op_T0_txa_v[`W-1]|~op_T0_txs_v[`W-1])), n1106_v, n1106_i2);
  spice_transistor_nmos_gnd g_1181((~notir3_v[`W-1]|~ir2_v[`W-1]|~ir6_v[`W-1]|~ir4_v[`W-1]|~notir5_v[`W-1]|~notir7_v[`W-1]|~clock1_v[`W-1]|~irline3_v[`W-1]), op_T0_tay_v, op_T0_tay_i1);
  spice_transistor_nmos_gnd t2487(~dpc29_0ADH17_v[`W-1], adh5_v, adh5_i3);
  spice_transistor_nmos_gnd t2486(~dpc29_0ADH17_v[`W-1], adh2_v, adh2_i5);
  spice_transistor_nmos t3446(~cclk_v[`W-1], n629_v, n760_v, n629_i0, n760_i0);
  spice_transistor_nmos t1723(~dpc5_SADL_v[`W-1], adl3_v, n998_v, adl3_i3, n998_i3);
  spice_transistor_nmos t1722(~dpc5_SADL_v[`W-1], adl4_v, n3_v, adl4_i4, n3_i3);
  spice_transistor_nmos t1721(~dpc5_SADL_v[`W-1], adl5_v, n280_v, adl5_i3, n280_i3);
  spice_transistor_nmos_gnd t1720(~notir5_v[`W-1], n503_v, n503_i0);
  spice_transistor_nmos t1727(~dpc5_SADL_v[`W-1], n721_v, adl7_v, n721_i3, adl7_i2);
  spice_transistor_nmos t1724(~dpc5_SADL_v[`W-1], adl2_v, n1389_v, adl2_i3, n1389_i2);
  spice_transistor_nmos_gnd t1729(~_ABL1_v[`W-1], abl1_v, abl1_i3);
  spice_transistor_nmos_gnd t2488(~dpc29_0ADH17_v[`W-1], adh4_v, adh4_i5);
  spice_transistor_nmos t3142(~dpc0_YSB_v[`W-1], n767_v, sb1_v, n767_i2, sb1_i11);
  spice_transistor_nmos t2727(~dpc9_DBADD_v[`W-1], idb2_v, alub2_v, idb2_i8, alub2_i2);
  spice_transistor_nmos t2724(~cp1_v[`W-1], n1147_v, idl7_v, n1147_i3, idl7_i1);
  spice_transistor_nmos_gnd t3030(~n90_v[`W-1], Pout6_v, Pout6_i1);
  spice_transistor_nmos_gnd t338(~pclp0_v[`W-1], n488_v, n488_i0);
  spice_transistor_nmos t334(~cclk_v[`W-1], n261_v, pipeUNK36_v, n261_i0, pipeUNK36_i0);
  spice_transistor_nmos t335(~cp1_v[`W-1], n959_v, n323_v, n959_i0, n323_i0);
  spice_transistor_nmos_gnd t332(~n182_v[`W-1], n442_v, n442_i0);
  spice_transistor_nmos_vdd t333(~dor1_v[`W-1], n798_v, n798_i1);
  spice_transistor_nmos_gnd t331(~n1602_v[`W-1], n1596_v, n1596_i0);
  spice_transistor_nmos t2804(~cclk_v[`W-1], n871_v, x7_v, n871_i1, x7_i2);
  spice_transistor_nmos t2800(~dpc8_nDBADD_v[`W-1], alub7_v, n423_v, alub7_i1, n423_i0);
  spice_transistor_nmos_gnd t1462(~t3_v[`W-1], op_T3_v, op_T3_i0);
  spice_transistor_nmos_gnd t205(~n999_v[`W-1], ab12_v, ab12_i0);
  spice_transistor_nmos_gnd g_1020((~ir6_v[`W-1]|~ir3_v[`W-1]|~ir4_v[`W-1]|~irline3_v[`W-1]|~t5_v[`W-1]|~notir5_v[`W-1]|~ir7_v[`W-1]|~ir2_v[`W-1]), xx_op_T5_jsr_v, xx_op_T5_jsr_i1);
  spice_transistor_nmos t117(~cp1_v[`W-1], n653_v, n1497_v, n653_i0, n1497_i0);
  spice_transistor_nmos_gnd t115(~notdor1_v[`W-1], dor1_v, dor1_i0);
  spice_transistor_nmos_gnd t112(~dpc12_0ADD_v[`W-1], alua3_v, alua3_i1);
  spice_transistor_nmos_gnd t110(~abh3_v[`W-1], n1346_v, n1346_i0);
  spice_transistor_nmos_gnd t111(~abh3_v[`W-1], n359_v, n359_i0);
  spice_transistor_nmos_gnd t118(~_ABH7_v[`W-1], abh7_v, abh7_i0);
  spice_transistor_nmos_gnd t2152(~n1534_v[`W-1], n763_v, n763_i0);
  spice_transistor_nmos t2554(~dpc32_PCHADH_v[`W-1], adh0_v, n1722_v, adh0_i6, n1722_i2);
  spice_transistor_nmos_gnd g_1254((~n453_v[`W-1]|~n609_v[`W-1]), n1213_v, n1213_i1);
  spice_transistor_nmos_gnd g_1255((~clock2_v[`W-1]|~notir0_v[`W-1]|~ir7_v[`W-1]), op_T__ora_and_eor_adc_v, op_T__ora_and_eor_adc_i2);
  spice_transistor_nmos_gnd g_1339((~op_T5_ind_y_v[`W-1]|~op_T4_abs_idx_v[`W-1]), n595_v, n595_i2);
  spice_transistor_nmos_gnd g_1338((~DA_AB2_v[`W-1]|~AxB3_v[`W-1]), n1610_v, n1610_i1);
  spice_transistor_nmos_gnd g_1335((~ir6_v[`W-1]|~notir1_v[`W-1]|~ir7_v[`W-1]), op_asl_rol_v, op_asl_rol_i2);
  spice_transistor_nmos_gnd g_1334((~notir7_v[`W-1]|~notir6_v[`W-1]|~ir4_v[`W-1]|~irline3_v[`W-1]|~ir5_v[`W-1]|~clock1_v[`W-1]), op_T0_cpy_iny_v, op_T0_cpy_iny_i1);
  spice_transistor_nmos_gnd g_1337((~_VEC_v[`W-1]|~C1x5Reset_v[`W-1]|~n264_v[`W-1]), n1712_v, n1712_i2);
  spice_transistor_nmos_gnd g_1336((~pd1_v[`W-1]|~clearIR_v[`W-1]), pd1_clearIR_v, pd1_clearIR_i3);
  spice_transistor_nmos_gnd g_1330((~_C01_v[`W-1]|~AxB1_v[`W-1]), __AxB1__C01_v, __AxB1__C01_i1);
  spice_transistor_nmos_gnd g_1333((~n1374_v[`W-1]|~n1578_v[`W-1]|~n645_v[`W-1]), n1368_v, n1368_i2);
  spice_transistor_nmos_gnd g_1332((~C67_v[`W-1]|~n1318_v[`W-1]), n637_v, n637_i1);
  spice_transistor_nmos_gnd t2461(~AxB5_v[`W-1], n1469_v, n1469_i1);
  spice_transistor_nmos_gnd t2462(~n231_v[`W-1], ONEBYTE_v, ONEBYTE_i0);
  spice_transistor_nmos_gnd t2467(~n133_v[`W-1], n602_v, n602_i0);
  spice_transistor_nmos_gnd t2466(~n300_v[`W-1], n847_v, n847_i0);
  spice_transistor_nmos_gnd t2469(~n709_v[`W-1], dpc18__DAA_v, dpc18__DAA_i1);
  spice_transistor_nmos_vdd t2468(~n133_v[`W-1], dpc2_XSB_v, dpc2_XSB_i2);
  spice_transistor_nmos_gnd g_1251((~t4_v[`W-1]|~notir0_v[`W-1]|~ir2_v[`W-1]|~ir3_v[`W-1]|~notir4_v[`W-1]), x_op_T4_ind_y_v, x_op_T4_ind_y_i3);
  spice_transistor_nmos_gnd g_1024((~notir3_v[`W-1]|~ir6_v[`W-1]|~ir7_v[`W-1]|~ir4_v[`W-1]|~irline3_v[`W-1]|~t2_v[`W-1]|~ir5_v[`W-1]|~ir2_v[`W-1]), op_T2_php_v, op_T2_php_i1);
  spice_transistor_nmos_gnd t2565(~abl7_v[`W-1], n1254_v, n1254_i2);
  spice_transistor_nmos_gnd g_1109((~t5_v[`W-1]|~notir0_v[`W-1]|~ir2_v[`W-1]|~ir3_v[`W-1]|~ir4_v[`W-1]), op_T5_ind_x_v, op_T5_ind_x_i2);
  spice_transistor_nmos_gnd t2566(~abl7_v[`W-1], n1195_v, n1195_i2);
  spice_transistor_nmos_gnd g_1201((~n236_v[`W-1]|~n192_v[`W-1]), n506_v, n506_i3);
  spice_transistor_nmos_gnd g_1200((~n1580_v[`W-1]|~n613_v[`W-1]), n1159_v, n1159_i1);
  spice_transistor_nmos_gnd g_1203((~n55_v[`W-1]|~cclk_v[`W-1]), n628_v, n628_i3);
  spice_transistor_nmos_vdd t2567(~abl7_v[`W-1], n1191_v, n1191_i2);
  spice_transistor_nmos t3398(~cclk_v[`W-1], pipeUNK17_v, n334_v, pipeUNK17_i0, n334_i2);
  spice_transistor_nmos_vdd t3399(~n1479_v[`W-1], ab1_v, ab1_i1);
  spice_transistor_nmos_vdd t2560(~n1041_v[`W-1], ab3_v, ab3_i0);
  spice_transistor_nmos t3391(~dpc6_SBS_v[`W-1], s7_v, sb7_v, s7_i2, sb7_i11);
  spice_transistor_nmos_gnd t3392(~n642_v[`W-1], ab2_v, ab2_i1);
  spice_transistor_nmos_gnd t3421(~aluanandb1_v[`W-1], n936_v, n936_i0);
  spice_transistor_nmos_gnd g_1537((~n1202_v[`W-1]&~n200_v[`W-1]), n293_v, n293_i3);
  spice_transistor_nmos_gnd g_1535((~n604_v[`W-1]&~n779_v[`W-1]), n1594_v, n1594_i2);
  spice_transistor_nmos_gnd g_1533((~n1262_v[`W-1]&~n572_v[`W-1]), n933_v, n933_i2);
  spice_transistor_nmos_gnd g_1532((~n1184_v[`W-1]&(~n1253_v[`W-1]|~n163_v[`W-1])), n1631_v, n1631_i2);
  spice_transistor_nmos_gnd g_1599(((~aluanandb0_v[`W-1]&~notalucin_v[`W-1])|~aluanorb0_v[`W-1]), DA_C01_v, DA_C01_i3);
  spice_transistor_nmos_gnd g_1539((~alua0_v[`W-1]&~alub0_v[`W-1]), aluanandb0_v, aluanandb0_i3);
  spice_transistor_nmos_gnd t1864(~_C45_v[`W-1], DA_C45_v, DA_C45_i0);
  spice_transistor_nmos_gnd t1865(~n1194_v[`W-1], Pout3_v, Pout3_i0);
  spice_transistor_nmos t1867(~cclk_v[`W-1], n824_v, n398_v, n824_i0, n398_i0);
  spice_transistor_nmos t1860(~dpc25_SBDB_v[`W-1], idb5_v, sb5_v, idb5_i3, sb5_i6);
  spice_transistor_nmos t1861(~dpc25_SBDB_v[`W-1], idb6_v, sb6_v, idb6_i4, sb6_i8);
  spice_transistor_nmos t1862(~dpc25_SBDB_v[`W-1], sb7_v, idb7_v, sb7_i5, idb7_i4);
  spice_transistor_nmos t1863(~cclk_v[`W-1], n1065_v, n1124_v, n1065_i0, n1124_i1);
  spice_transistor_nmos_gnd g_1021((~notir2_v[`W-1]|~ir4_v[`W-1]|~irline3_v[`W-1]|~ir5_v[`W-1]|~notir3_v[`W-1]|~t2_v[`W-1]|~notir6_v[`W-1]|~ir7_v[`W-1]), op_T2_jmp_abs_v, op_T2_jmp_abs_i1);
  spice_transistor_nmos_vdd t2942(~n617_v[`W-1], n676_v, n676_i3);
  spice_transistor_nmos_gnd g_1023((~ir7_v[`W-1]|~ir3_v[`W-1]|~notir6_v[`W-1]|~irline3_v[`W-1]|~ir4_v[`W-1]|~t5_v[`W-1]|~ir2_v[`W-1]), op_T5_rti_rts_v, op_T5_rti_rts_i1);
  spice_transistor_nmos_gnd g_1022((~ir7_v[`W-1]|~t4_v[`W-1]|~notir6_v[`W-1]|~notir2_v[`W-1]|~irline3_v[`W-1]|~ir4_v[`W-1]|~notir3_v[`W-1]), op_T4_jmp_v, op_T4_jmp_i1);
  spice_transistor_nmos_gnd t1868(~VEC0_v[`W-1], n728_v, n728_i0);
  spice_transistor_nmos_gnd g_1027((~ir3_v[`W-1]|~t4_v[`W-1]|~ir7_v[`W-1]|~ir6_v[`W-1]|~irline3_v[`W-1]|~ir4_v[`W-1]|~ir5_v[`W-1]|~ir2_v[`W-1]), op_T4_brk_v, op_T4_brk_i1);
  spice_transistor_nmos_gnd g_1026((~ir2_v[`W-1]|~notir3_v[`W-1]|~ir7_v[`W-1]|~ir4_v[`W-1]|~irline3_v[`W-1]), op_push_pull_v, op_push_pull_i1);
  spice_transistor_nmos_gnd t2444(~op_store_v[`W-1], _op_store_v, _op_store_i0);
  spice_transistor_nmos_gnd g_1319((~n1184_v[`W-1]|~n1643_v[`W-1]), n410_v, n410_i1);
  spice_transistor_nmos_gnd t2266(~n862_v[`W-1], n445_v, n445_i3);
  spice_transistor_nmos_gnd t2264(~pch5_v[`W-1], n499_v, n499_i0);
  spice_transistor_nmos t2263(~dpc0_YSB_v[`W-1], n733_v, sb5_v, n733_i1, sb5_i7);
  spice_transistor_nmos t2262(~dpc0_YSB_v[`W-1], n518_v, sb6_v, n518_i2, sb6_i10);
  spice_transistor_nmos_gnd t2261(~n47_v[`W-1], n603_v, n603_i0);
  spice_transistor_nmos t2260(~dpc0_YSB_v[`W-1], n658_v, dasb4_v, n658_i1, dasb4_i10);
  spice_transistor_nmos_gnd t2068(~pipe_VEC_v[`W-1], n1578_v, n1578_i0);
  spice_transistor_nmos t3175(~dpc39_PCLPCL_v[`W-1], pcl7_v, n1647_v, pcl7_i2, n1647_i3);
  spice_transistor_nmos_vdd t2066(~n1028_v[`W-1], RnWstretched_v, RnWstretched_i1);
  spice_transistor_nmos t2281(~cclk_v[`W-1], n616_v, n460_v, n616_i0, n460_i0);
  spice_transistor_nmos_vdd t2280(~n628_v[`W-1], dpc24_ACSB_v, dpc24_ACSB_i0);
  spice_transistor_nmos t1266(~cclk_v[`W-1], pipeUNK29_v, n169_v, pipeUNK29_i0, n169_i0);
  spice_transistor_nmos_gnd t1267(~pipeUNK26_v[`W-1], n1714_v, n1714_i0);
  spice_transistor_nmos t1264(~cp1_v[`W-1], n1687_v, notdor0_v, n1687_i0, notdor0_i0);
  spice_transistor_nmos t1265(~cp1_v[`W-1], n299_v, n1625_v, n299_i0, n1625_i0);
  spice_transistor_nmos_gnd t1262(~n1620_v[`W-1], ir3_v, ir3_i1);
  spice_transistor_nmos t1263(~cclk_v[`W-1], pipeUNK11_v, n862_v, pipeUNK11_i1, n862_i0);
  spice_transistor_nmos_gnd g_1155((~n562_v[`W-1]|~n882_v[`W-1]), n1374_v, n1374_i2);
  spice_transistor_nmos t451(~cp1_v[`W-1], n402_v, notRnWprepad_v, n402_i0, notRnWprepad_i0);
  spice_transistor_nmos t450(~dpc9_DBADD_v[`W-1], alub0_v, idb0_v, alub0_i1, idb0_i4);
  spice_transistor_nmos t457(~cclk_v[`W-1], n568_v, notidl5_v, n568_i0, notidl5_i0);
  spice_transistor_nmos_vdd t456(~cclk_v[`W-1], adh1_v, adh1_i2);
  spice_transistor_nmos t455(~dpc2_XSB_v[`W-1], n871_v, sb7_v, n871_i0, sb7_i1);
  spice_transistor_nmos t454(~cclk_v[`W-1], n1717_v, n1113_v, n1717_i0, n1113_i0);
  spice_transistor_nmos_gnd t459(~abl3_v[`W-1], n990_v, n990_i0);
  spice_transistor_nmos_gnd t458(~abl3_v[`W-1], n138_v, n138_i0);
  spice_transistor_nmos_gnd g_1159((~op_T__ora_and_eor_adc_v[`W-1]|~op_T__shift_a_v[`W-1]|~op_T0_lda_v[`W-1]|~op_T0_tya_v[`W-1]|~op_T__adc_sbc_v[`W-1]|~op_T0_pla_v[`W-1]|~op_T0_txa_v[`W-1]), n1455_v, n1455_i3);
  spice_transistor_nmos_vdd t2153(~n1534_v[`W-1], dpc8_nDBADD_v, dpc8_nDBADD_i3);
  spice_transistor_nmos_gnd t691(~pch6_v[`W-1], n278_v, n278_i0);
  spice_transistor_nmos_gnd t922(~notRdy0_v[`W-1], n372_v, n372_i0);
  spice_transistor_nmos_gnd t693(~n567_v[`W-1], n1026_v, n1026_i0);
  spice_transistor_nmos_gnd t692(~n567_v[`W-1], n171_v, n171_i0);
  spice_transistor_nmos t926(~cp1_v[`W-1], n457_v, notdor3_v, n457_i0, notdor3_i0);
  spice_transistor_nmos t924(~cclk_v[`W-1], n359_v, _ABH3_v, n359_i1, _ABH3_i0);
  spice_transistor_nmos_gnd t929(~notdor2_v[`W-1], dor2_v, dor2_i1);
  spice_transistor_nmos_gnd t2658(~n359_v[`W-1], ab11_v, ab11_i1);
  spice_transistor_nmos t2601(~cclk_v[`W-1], n862_v, pipeT_SYNC_v, n862_i3, pipeT_SYNC_i0);
  spice_transistor_nmos t2600(~cclk_v[`W-1], n213_v, notidl1_v, n213_i1, notidl1_i0);
  spice_transistor_nmos t2602(~cp1_v[`W-1], n789_v, notdor7_v, n789_i1, notdor7_i0);
  spice_transistor_nmos_gnd t2605(~n1660_v[`W-1], n855_v, n855_i2);
  spice_transistor_nmos_vdd t2606(~n1660_v[`W-1], n1100_v, n1100_i3);
  spice_transistor_nmos t1008(~cp1_v[`W-1], notRdy0_v, n902_v, notRdy0_i5, n902_i0);
  spice_transistor_nmos_gnd t1009(~ir2_v[`W-1], notir2_v, notir2_i0);
  spice_transistor_nmos_gnd t1000(~n1110_v[`W-1], n771_v, n771_i0);
  spice_transistor_nmos_gnd t1006(~pipeUNK27_v[`W-1], n920_v, n920_i1);
  spice_transistor_nmos_gnd t1398(~op_T2_branch_v[`W-1], n636_v, n636_i0);
  spice_transistor_nmos t1392(~cclk_v[`W-1], n111_v, pd2_v, n111_i0, pd2_i0);
  spice_transistor_nmos t1393(~cclk_v[`W-1], n62_v, pd7_v, n62_i0, pd7_i0);
  spice_transistor_nmos t1391(~cp1_v[`W-1], n1290_v, n698_v, n1290_i0, n698_i0);
  spice_transistor_nmos_gnd t1397(~notalu1_v[`W-1], alu1_v, alu1_i1);
  spice_transistor_nmos t1394(~cclk_v[`W-1], n374_v, pd6_v, n374_i0, pd6_i0);
  spice_transistor_nmos_gnd t1395(~n675_v[`W-1], n888_v, n888_i0);
  spice_transistor_nmos t589(~dpc43_DL_DB_v[`W-1], idb4_v, n1095_v, idb4_i0, n1095_i1);
  spice_transistor_nmos t588(~dpc43_DL_DB_v[`W-1], idb3_v, n1661_v, idb3_i0, n1661_i1);
  spice_transistor_nmos_gnd t855(~_op_branch_bit6_v[`W-1], n846_v, n846_i0);
  spice_transistor_nmos_gnd g_1318((~notir4_v[`W-1]|~notir3_v[`W-1]|~t4_v[`W-1]), op_T4_mem_abs_idx_v, op_T4_mem_abs_idx_i2);
  spice_transistor_nmos t3359(~cclk_v[`W-1], n824_v, pipeUNK34_v, n824_i1, pipeUNK34_i0);
  spice_transistor_nmos t1484(~dpc41_DL_ADL_v[`W-1], adl2_v, n1424_v, adl2_i2, n1424_i3);
  spice_transistor_nmos t1485(~dpc41_DL_ADL_v[`W-1], adl0_v, n719_v, adl0_i3, n719_i3);
  spice_transistor_nmos t1482(~dpc41_DL_ADL_v[`W-1], adl4_v, n1095_v, adl4_i3, n1095_i2);
  spice_transistor_nmos t1483(~dpc41_DL_ADL_v[`W-1], adl1_v, n87_v, adl1_i2, n87_i3);
  spice_transistor_nmos t1481(~dpc41_DL_ADL_v[`W-1], adl3_v, n1661_v, adl3_i2, n1661_i2);
  spice_transistor_nmos_gnd g_1288((~op_SRS_v[`W-1]|~n781_v[`W-1]), n160_v, n160_i2);
  spice_transistor_nmos_gnd t1337(~idb3_v[`W-1], n1600_v, n1600_i0);
  spice_transistor_nmos_vdd t1739(~cclk_v[`W-1], sb1_v, sb1_i6);
  spice_transistor_nmos_gnd t1735(~notidl7_v[`W-1], idl7_v, idl7_i0);
  spice_transistor_nmos_gnd t1731(~pchp3_v[`W-1], n141_v, n141_i0);
  spice_transistor_nmos t1732(~cp1_v[`W-1], n1528_v, n1215_v, n1528_i0, n1215_i1);
  spice_transistor_nmos t1733(~cp1_v[`W-1], n1161_v, n109_v, n1161_i0, n109_i1);
  spice_transistor_nmos_gnd g_1315((~__AxB_4_v[`W-1]|~C34_v[`W-1]), _AxB_4__C34_v, _AxB_4__C34_i1);
  spice_transistor_nmos t329(~dpc0_YSB_v[`W-1], n564_v, dasb0_v, n564_i0, dasb0_i1);
  spice_transistor_nmos t321(~dpc21_ADDADL_v[`W-1], alu2_v, adl2_v, alu2_i0, adl2_i0);
  spice_transistor_nmos t323(~dpc21_ADDADL_v[`W-1], adl0_v, alu0_v, adl0_i0, alu0_i0);
  spice_transistor_nmos t322(~dpc21_ADDADL_v[`W-1], adl1_v, alu1_v, adl1_i0, alu1_i0);
  spice_transistor_nmos_gnd t326(~n1699_v[`W-1], n913_v, n913_i0);
  spice_transistor_nmos_gnd g_1105((~ir3_v[`W-1]|~ir7_v[`W-1]|~ir6_v[`W-1]|~ir4_v[`W-1]|~irline3_v[`W-1]|~t3_v[`W-1]|~ir2_v[`W-1]|~notir5_v[`W-1]), op_T3_jsr_v, op_T3_jsr_i1);
  spice_transistor_nmos_gnd t3450(~n138_v[`W-1], ab3_v, ab3_i1);
  spice_transistor_nmos t2129(~H1x1_v[`W-1], Pout3_v, idb3_v, Pout3_i1, idb3_i5);
  spice_transistor_nmos t2551(~dpc32_PCHADH_v[`W-1], adh3_v, n141_v, adh3_i6, n141_i2);
  spice_transistor_nmos_gnd t215(~alucout_v[`W-1], n206_v, n206_i0);
  spice_transistor_nmos_gnd t217(~n241_v[`W-1], n1033_v, n1033_i0);
  spice_transistor_nmos_gnd t213(~n867_v[`W-1], n876_v, n876_i0);
  spice_transistor_nmos t212(~cclk_v[`W-1], pipeUNK22_v, n29_v, pipeUNK22_i0, n29_i0);
  spice_transistor_nmos_vdd t218(~n241_v[`W-1], dpc21_ADDADL_v, dpc21_ADDADL_i0);
  spice_transistor_nmos_gnd g_1411((~n852_v[`W-1]|~n1205_v[`W-1]), n260_v, n260_i1);
  spice_transistor_nmos_gnd g_1415((~op_T0_bit_v[`W-1]|~op_T0_and_v[`W-1]), n669_v, n669_i2);
  spice_transistor_nmos_gnd g_1081((~n459_v[`W-1]|~n43_v[`W-1]), n625_v, n625_i3);
  spice_transistor_nmos_gnd g_1417((~pipeUNK10_v[`W-1]&~pipeUNK09_v[`W-1]), n1111_v, n1111_i2);
  spice_transistor_nmos_gnd t103(~y1_v[`W-1], n1138_v, n1138_i0);
  spice_transistor_nmos_vdd t104(~n963_v[`W-1], ab14_v, ab14_i0);
  spice_transistor_nmos_vdd t109(~abh3_v[`W-1], n1296_v, n1296_i0);
  spice_transistor_nmos_gnd t57(~pch4_v[`W-1], n1400_v, n1400_i0);
  spice_transistor_nmos_gnd g_1283((~notir5_v[`W-1]|~notir3_v[`W-1]|~ir2_v[`W-1]|~ir6_v[`W-1]|~ir4_v[`W-1]|~notir1_v[`W-1]|~notir7_v[`W-1]|~clock1_v[`W-1]), op_T0_tax_v, op_T0_tax_i1);
  spice_transistor_nmos_vdd t3353(~cclk_v[`W-1], adl7_v, adl7_i7);
  spice_transistor_nmos_gnd t1640(~n1521_v[`W-1], n242_v, n242_i1);
  spice_transistor_nmos_gnd g_1308((~notRdy0_v[`W-1]|~n1214_v[`W-1]), fetch_v, fetch_i1);
  spice_transistor_nmos_gnd g_1309((~AxB5_v[`W-1]|~DA_C45_v[`W-1]|~n647_v[`W-1]|~n122_v[`W-1]), n570_v, n570_i1);
  spice_transistor_nmos_gnd g_1300((~n43_v[`W-1]|~n1477_v[`W-1]), n1541_v, n1541_i3);
  spice_transistor_nmos_gnd g_1301((~brk_done_v[`W-1]|~p2_v[`W-1]), n334_v, n334_i4);
  spice_transistor_nmos_gnd g_1302((~ir4_v[`W-1]|~t2_v[`W-1]|~ir2_v[`W-1]|~ir7_v[`W-1]|~irline3_v[`W-1]), op_T2_stack_v, op_T2_stack_i1);
  spice_transistor_nmos_gnd g_1304((~n43_v[`W-1]|~n1509_v[`W-1]), n611_v, n611_i3);
  spice_transistor_nmos_gnd g_1306((~aluanorb1_v[`W-1]|~n936_v[`W-1]), AxB1_v, AxB1_i3);
  spice_transistor_nmos_gnd t2472(~db4_v[`W-1], n1075_v, n1075_i1);
  spice_transistor_nmos_gnd t2473(~dpc34_PCLC_v[`W-1], n1007_v, n1007_i0);
  spice_transistor_nmos_gnd t2470(~x0_v[`W-1], n987_v, n987_i1);
  spice_transistor_nmos_gnd t2246(~n1649_v[`W-1], n795_v, n795_i0);
  spice_transistor_nmos t2477(~dpc31_PCHPCH_v[`W-1], pch4_v, n27_v, pch4_i2, n27_i1);
  spice_transistor_nmos t2475(~dpc31_PCHPCH_v[`W-1], pch6_v, n652_v, pch6_i2, n652_i1);
  spice_transistor_nmos t1641(~dpc1_SBY_v[`W-1], y1_v, sb1_v, y1_i2, sb1_i5);
  spice_transistor_nmos t2479(~dpc31_PCHPCH_v[`W-1], pch2_v, n1496_v, pch2_i1, n1496_i1);
  spice_transistor_nmos_gnd t3066(~n1462_v[`W-1], dpc38_PCLADL_v, dpc38_PCLADL_i9);
  spice_transistor_nmos_gnd t3234(~pch2_v[`W-1], n1265_v, n1265_i1);
  spice_transistor_nmos t2010(~cp1_v[`W-1], n1409_v, n916_v, n1409_i0, n916_i0);
  spice_transistor_nmos_gnd t3064(~adl2_v[`W-1], n935_v, n935_i0);
  spice_transistor_nmos_gnd t3355(~pclp1_v[`W-1], n976_v, n976_i3);
  spice_transistor_nmos_gnd t3065(~n5_v[`W-1], n146_v, n146_i3);
  spice_transistor_nmos_gnd g_1235((~op_T2_brk_v[`W-1]|~op_T3_jsr_v[`W-1]), n824_v, n824_i3);
  spice_transistor_nmos t3417(~cclk_v[`W-1], x_op_T__adc_sbc_v, pipeUNK03_v, x_op_T__adc_sbc_i0, pipeUNK03_i0);
  spice_transistor_nmos_gnd g_1231((~RnWstretched_v[`W-1]|~n466_v[`W-1]), n7_v, n7_i2);
  spice_transistor_nmos_gnd g_1232((~ir3_v[`W-1]|~notir2_v[`W-1]|~t2_v[`W-1]), op_T2_zp_zp_idx_v, op_T2_zp_zp_idx_i2);
  spice_transistor_nmos_gnd g_1233((~alub1_v[`W-1]|~alua1_v[`W-1]), aluanorb1_v, aluanorb1_i3);
  spice_transistor_nmos_gnd g_1543((~n1408_v[`W-1]&~n980_v[`W-1]), n473_v, n473_i2);
  spice_transistor_nmos_gnd g_1540((~n110_v[`W-1]&~n681_v[`W-1]), __AxB_2_v, __AxB_2_i3);
  spice_transistor_nmos_gnd t2011(~n666_v[`W-1], n862_v, n862_i1);
  spice_transistor_nmos_gnd g_1546(((~n118_v[`W-1]|~n888_v[`W-1])&~n264_v[`W-1]), n480_v, n480_i1);
  spice_transistor_nmos_gnd g_1548((~alua2_v[`W-1]&~alub2_v[`W-1]), n681_v, n681_i5);
  spice_transistor_nmos_gnd g_1018((~n510_v[`W-1]|~n218_v[`W-1]|~op_T3_branch_v[`W-1]|~n1258_v[`W-1]), n1716_v, n1716_i1);
  spice_transistor_nmos_gnd g_1019((~AxB5_v[`W-1]|~_C45_v[`W-1]), __AxB5__C45_v, __AxB5__C45_i1);
  spice_transistor_nmos_gnd g_1075((~RnWstretched_v[`W-1]|~dor2_v[`W-1]), n37_v, n37_i2);
  spice_transistor_nmos t2278(~cclk_v[`W-1], n927_v, notir4_v, n927_i0, notir4_i0);
  spice_transistor_nmos_gnd t2279(~n628_v[`W-1], n1335_v, n1335_i0);
  spice_transistor_nmos t2592(~dpc13_ORS_v[`W-1], n404_v, n296_v, n404_i0, n296_i5);
  spice_transistor_nmos_gnd t8(~db2_v[`W-1], n1199_v, n1199_i0);
  spice_transistor_nmos_vdd t4(~n826_v[`W-1], ab8_v, ab8_i0);
  spice_transistor_nmos_gnd t5(~db1_v[`W-1], n1319_v, n1319_i0);
  spice_transistor_nmos_gnd t2(~notalucout_v[`W-1], alucout_v, alucout_i0);
  spice_transistor_nmos_gnd t0(~pipeVectorA0_v[`W-1], n_0_ADL0_v, n_0_ADL0_i0);
  spice_transistor_nmos_vdd t1(~n1608_v[`W-1], ab13_v, ab13_i0);
  spice_transistor_nmos t2079(~cclk_v[`W-1], n728_v, pipeVectorA0_v, n728_i1, pipeVectorA0_i1);
  spice_transistor_nmos_gnd t2076(~abh0_v[`W-1], n381_v, n381_i1);
  spice_transistor_nmos t2077(~cclk_v[`W-1], pipeUNK13_v, n1045_v, pipeUNK13_i0, n1045_i1);
  spice_transistor_nmos t2074(~cclk_v[`W-1], n1177_v, n1069_v, n1177_i0, n1069_i0);
  spice_transistor_nmos_gnd t2075(~abh0_v[`W-1], n1315_v, n1315_i0);
  spice_transistor_nmos_gnd t2013(~pchp7_v[`W-1], n1206_v, n1206_i0);
  spice_transistor_nmos_gnd t1258(~n1632_v[`W-1], A_B5_v, A_B5_i0);
  spice_transistor_nmos_gnd t1253(~n31_v[`W-1], Pout0_v, Pout0_i1);
  spice_transistor_nmos t1257(~cclk_v[`W-1], Reset0_v, pipephi2Reset0x_v, Reset0_i0, pipephi2Reset0x_i0);
  spice_transistor_nmos_vdd t1254(~dor3_v[`W-1], n42_v, n42_i0);
  spice_transistor_nmos_gnd g_1112((~brk_done_v[`W-1]|~op_rti_rts_v[`W-1]|~op_T4_ind_x_v[`W-1]|~x_op_T3_ind_y_v[`W-1]|~op_T2_jsr_v[`W-1]|~n389_v[`W-1]), n300_v, n300_i2);
  spice_transistor_nmos_gnd g_1163((~op_EORS_v[`W-1]|~op_SRS_v[`W-1]|~op_ORS_v[`W-1]|~op_ANDS_v[`W-1]), op_SUMS_v, op_SUMS_i2);
  spice_transistor_nmos_gnd g_1164((~notir7_v[`W-1]|~ir6_v[`W-1]|~ir5_v[`W-1]|~notir2_v[`W-1]|~irline3_v[`W-1]), op_sty_cpy_mem_v, op_sty_cpy_mem_i1);
  spice_transistor_nmos_gnd g_1165((~C12_v[`W-1]|~__AxB_2_v[`W-1]), _AxB_2__C12_v, _AxB_2__C12_i1);
  spice_transistor_nmos_vdd t466(~n35_v[`W-1], dpc7_SS_v, dpc7_SS_i7);
  spice_transistor_nmos_gnd g_1670(((~notRdy0_v[`W-1]&~pipeT2out_v[`W-1])|(~pipeT_SYNC_v[`W-1]&~n16_v[`W-1])), n1091_v, n1091_i2);
  spice_transistor_nmos_gnd t464(~n378_v[`W-1], t5_v, t5_i0);
  spice_transistor_nmos_gnd t465(~n35_v[`W-1], n71_v, n71_i0);
  spice_transistor_nmos_gnd t463(~a6_v[`W-1], n1356_v, n1356_i0);
  spice_transistor_nmos_vdd t460(~abl3_v[`W-1], n1041_v, n1041_i0);
  spice_transistor_nmos_gnd t461(~pipeUNK11_v[`W-1], n1214_v, n1214_i0);
  spice_transistor_nmos_gnd g_1492((~n1303_v[`W-1]&~n383_v[`W-1]), n782_v, n782_i2);
  spice_transistor_nmos_gnd g_1495((~n918_v[`W-1]&~n1063_v[`W-1]), __AxB_4_v, __AxB_4_i3);
  spice_transistor_nmos_vdd t918(~n1195_v[`W-1], n1254_v, n1254_i0);
  spice_transistor_nmos_gnd g_1179((~ir4_v[`W-1]|~ir2_v[`W-1]|~notir6_v[`W-1]|~notir3_v[`W-1]|~ir7_v[`W-1]|~t2_v[`W-1]|~irline3_v[`W-1]|~ir5_v[`W-1]), op_T2_pha_v, op_T2_pha_i1);
  spice_transistor_nmos_gnd t2618(~notdor7_v[`W-1], dor7_v, dor7_i0);
  spice_transistor_nmos_gnd t2613(~n1315_v[`W-1], n826_v, n826_i2);
  spice_transistor_nmos_gnd t2611(~n556_v[`W-1], n1344_v, n1344_i2);
  spice_transistor_nmos t2616(~cclk_v[`W-1], n733_v, y5_v, n733_i2, y5_i1);
  spice_transistor_nmos_gnd t2614(~n1265_v[`W-1], n1202_v, n1202_i0);
  spice_transistor_nmos t2916(~dpc33_PCHDB_v[`W-1], n1301_v, idb5_v, n1301_i3, idb5_i8);
  spice_transistor_nmos_gnd g_1074((~n43_v[`W-1]|~n509_v[`W-1]), n1270_v, n1270_i3);
  spice_transistor_nmos_gnd t2107(~n1138_v[`W-1], n767_v, n767_i1);
  spice_transistor_nmos_gnd t869(~n291_v[`W-1], n1157_v, n1157_i0);
  spice_transistor_nmos_gnd t860(~adl7_v[`W-1], n1046_v, n1046_i0);
  spice_transistor_nmos_gnd t861(~n1107_v[`W-1], n389_v, n389_i1);
  spice_transistor_nmos_gnd t866(~y2_v[`W-1], n1484_v, n1484_i0);
  spice_transistor_nmos t1103(~cclk_v[`W-1], n1724_v, x6_v, n1724_i1, x6_i0);
  spice_transistor_nmos_vdd t1101(~cclk_v[`W-1], adl3_v, adl3_i1);
  spice_transistor_nmos t1107(~dpc17_SUMS_v[`W-1], __AxBxC_1_v, notaluoutmux1_v, __AxBxC_1_i0, notaluoutmux1_i1);
  spice_transistor_nmos t1106(~dpc17_SUMS_v[`W-1], __AxBxC_0_v, notaluoutmux0_v, __AxBxC_0_i0, notaluoutmux0_i1);
  spice_transistor_nmos_gnd t1105(~n1238_v[`W-1], dpc25_SBDB_v, dpc25_SBDB_i0);
  spice_transistor_nmos t1109(~dpc17_SUMS_v[`W-1], __AxBxC_3_v, n1071_v, __AxBxC_3_i0, n1071_i3);
  spice_transistor_nmos t1108(~dpc17_SUMS_v[`W-1], __AxBxC_2_v, n740_v, __AxBxC_2_i0, n740_i2);
  spice_transistor_nmos t2118(~cclk_v[`W-1], n1231_v, pipeUNK21_v, n1231_i0, pipeUNK21_i1);
  spice_transistor_nmos_gnd g_1174((~irline3_v[`W-1]|~notir3_v[`W-1]|~notir6_v[`W-1]|~clock1_v[`W-1]|~notir7_v[`W-1]|~ir2_v[`W-1]|~notir4_v[`W-1]), op_T0_cld_sed_v, op_T0_cld_sed_i2);
  spice_transistor_nmos_gnd g_1175((~clock1_v[`W-1]|~notir7_v[`W-1]|~notir1_v[`W-1]|~ir6_v[`W-1]|~notir5_v[`W-1]), op_T0_ldx_tax_tsx_v, op_T0_ldx_tax_tsx_i1);
  spice_transistor_nmos_gnd g_1173((~notRdy0_v[`W-1]|~n1716_v[`W-1]), n180_v, n180_i1);
  spice_transistor_nmos_vdd t1035(~n358_v[`W-1], n1467_v, n1467_i0);
  spice_transistor_nmos_vdd t481(~n670_v[`W-1], n1417_v, n1417_i0);
  spice_transistor_nmos_gnd t482(~n994_v[`W-1], ab10_v, ab10_i1);
  spice_transistor_nmos_gnd t489(~n1439_v[`W-1], n518_v, n518_i1);
  spice_transistor_nmos t2552(~dpc32_PCHADH_v[`W-1], adh2_v, n1496_v, adh2_i6, n1496_i2);
  spice_transistor_nmos t2625(~cclk_v[`W-1], nnT2BR_v, n1269_v, nnT2BR_i1, n1269_i1);
  spice_transistor_nmos_vdd t1749(~n1596_v[`W-1], dpc27_SBADH_v, dpc27_SBADH_i0);
  spice_transistor_nmos_gnd t1748(~n1596_v[`W-1], n1271_v, n1271_i0);
  spice_transistor_nmos t1741(~cclk_v[`W-1], n897_v, n1211_v, n897_i0, n1211_i0);
  spice_transistor_nmos t1740(~cclk_v[`W-1], n182_v, n265_v, n182_i1, n265_i0);
  spice_transistor_nmos_gnd t1745(~n966_v[`W-1], n1635_v, n1635_i1);
  spice_transistor_nmos_gnd t1747(~n559_v[`W-1], n770_v, n770_i0);
  spice_transistor_nmos_vdd t1746(~n966_v[`W-1], dpc29_0ADH17_v, dpc29_0ADH17_i2);
  spice_transistor_nmos t1938(~cclk_v[`W-1], n1358_v, n521_v, n1358_i0, n521_i0);
  spice_transistor_nmos_gnd t1939(~n318_v[`W-1], Pout1_v, Pout1_i1);
  spice_transistor_nmos_gnd g_1086((~idb1_v[`W-1]|~idb4_v[`W-1]|~idb2_v[`W-1]|~idb7_v[`W-1]|~idb5_v[`W-1]|~idb0_v[`W-1]|~idb6_v[`W-1]|~idb3_v[`W-1]), DBZ_v, DBZ_i2);
  spice_transistor_nmos_gnd g_1172((~pipeUNK36_v[`W-1]|~n1137_v[`W-1]|~n916_v[`W-1]|~notRdy0_v[`W-1]), short_circuit_idx_add_v, short_circuit_idx_add_i1);
  spice_transistor_nmos t2130(~H1x1_v[`W-1], Pout6_v, idb6_v, Pout6_i0, idb6_i5);
  spice_transistor_nmos_gnd t2459(~abh7_v[`W-1], n659_v, n659_i1);
  spice_transistor_nmos t260(~cp1_v[`W-1], n931_v, n1674_v, n931_i0, n1674_i0);
  spice_transistor_nmos t261(~cp1_v[`W-1], n1526_v, n1450_v, n1526_i0, n1450_i0);
  spice_transistor_nmos_gnd t262(~op_T0_v[`W-1], n638_v, n638_i0);
  spice_transistor_nmos_gnd t263(~n512_v[`W-1], n154_v, n154_i2);
  spice_transistor_nmos_gnd t265(~n1427_v[`W-1], n1448_v, n1448_i0);
  spice_transistor_nmos_gnd t266(~n223_v[`W-1], n1357_v, n1357_i0);
  spice_transistor_nmos_gnd t267(~n1219_v[`W-1], n1002_v, n1002_i0);
  spice_transistor_nmos t268(~H1x1_v[`W-1], idb0_v, Pout0_v, idb0_i2, Pout0_i0);
  spice_transistor_nmos t269(~cclk_v[`W-1], n604_v, n1477_v, n604_i0, n1477_i0);
  spice_transistor_nmos t3308(~cclk_v[`W-1], n1712_v, pipeVectorA2_v, n1712_i0, pipeVectorA2_i1);
  spice_transistor_nmos t2745(~dpc37_PCLDB_v[`W-1], n723_v, idb3_v, n723_i2, idb3_i9);
  spice_transistor_nmos t2746(~dpc37_PCLDB_v[`W-1], n976_v, idb1_v, n976_i1, idb1_i7);
  spice_transistor_nmos t2215(~dpc15_ANDS_v[`W-1], n350_v, n1071_v, n350_i2, n1071_i5);
  spice_transistor_nmos_gnd t3348(~y5_v[`W-1], n981_v, n981_i1);
  spice_transistor_nmos t3195(~dpc4_SSB_v[`W-1], n332_v, dasb0_v, n332_i3, dasb0_i12);
  spice_transistor_nmos_gnd t2743(~n519_v[`W-1], n670_v, n670_i2);
  spice_transistor_nmos_gnd g_1085((~n1624_v[`W-1]|~n139_v[`W-1]), n169_v, n169_i2);
  spice_transistor_nmos t86(~cclk_v[`W-1], n490_v, notidl4_v, n490_i0, notidl4_i0);
  spice_transistor_nmos t85(~cclk_v[`W-1], n1673_v, op_T__bit_v, n1673_i0, op_T__bit_i0);
  spice_transistor_nmos t84(~cclk_v[`W-1], n513_v, pipeUNK06_v, n513_i0, pipeUNK06_i0);
  spice_transistor_nmos t83(~H1x1_v[`W-1], idb2_v, Pout2_v, idb2_i0, Pout2_i0);
  spice_transistor_nmos t82(~H1x1_v[`W-1], Pout7_v, idb7_v, Pout7_i0, idb7_i0);
  spice_transistor_nmos t2591(~cp1_v[`W-1], n468_v, n18_v, n468_i0, n18_i0);
  spice_transistor_nmos_gnd g_1046((~notir6_v[`W-1]|~notir7_v[`W-1]|~clock1_v[`W-1]|~notir0_v[`W-1]|~ir5_v[`W-1]), op_T0_cmp_v, op_T0_cmp_i1);
  spice_transistor_nmos_gnd t886(~pipeUNK18_v[`W-1], n850_v, n850_i0);
  spice_transistor_nmos_gnd t2449(~n754_v[`W-1], n1595_v, n1595_i0);
  spice_transistor_nmos t2446(~cclk_v[`W-1], nots1_v, n1711_v, nots1_i1, n1711_i0);
  spice_transistor_nmos_gnd t2445(~op_SRS_v[`W-1], n139_v, n139_i0);
  spice_transistor_nmos_gnd t2442(~dpc28_0ADH0_v[`W-1], adh0_v, adh0_i3);
  spice_transistor_nmos_gnd t3404(~x3_v[`W-1], n1521_v, n1521_i1);
  spice_transistor_nmos_gnd t2829(~x2_v[`W-1], n890_v, n890_i1);
  spice_transistor_nmos_gnd t3406(~n355_v[`W-1], n593_v, n593_i1);
  spice_transistor_nmos_vdd t3407(~n355_v[`W-1], dpc4_SSB_v, dpc4_SSB_i9);
  spice_transistor_nmos_gnd g_1229((~_DA_ADD1_v[`W-1]|~_DA_ADD2_v[`W-1]), n867_v, n867_i2);
  spice_transistor_nmos_gnd g_1228((~n647_v[`W-1]|~n1632_v[`W-1]), AxB5_v, AxB5_i3);
  spice_transistor_nmos_gnd t2255(~dpc12_0ADD_v[`W-1], alua2_v, alua2_i1);
  spice_transistor_nmos_gnd g_1223((~n1132_v[`W-1]|~pipephi2Reset0x_v[`W-1]), n717_v, n717_i2);
  spice_transistor_nmos_gnd g_1222((~notir0_v[`W-1]|~ir2_v[`W-1]|~t4_v[`W-1]|~ir4_v[`W-1]|~ir3_v[`W-1]), op_T4_ind_x_v, op_T4_ind_x_i2);
  spice_transistor_nmos_gnd g_1220((~n507_v[`W-1]|~n954_v[`W-1]|~n253_v[`W-1]), n279_v, n279_i1);
  spice_transistor_nmos_gnd g_1227((~n853_v[`W-1]|~n572_v[`W-1]), n1517_v, n1517_i1);
  spice_transistor_nmos_gnd g_1226((~dor3_v[`W-1]|~RnWstretched_v[`W-1]), n643_v, n643_i2);
  spice_transistor_nmos_gnd g_1225((~ir3_v[`W-1]|~ir7_v[`W-1]|~ir4_v[`W-1]|~notir5_v[`W-1]|~ir6_v[`W-1]|~ir2_v[`W-1]|~t5_v[`W-1]|~irline3_v[`W-1]), op_T5_jsr_v, op_T5_jsr_i2);
  spice_transistor_nmos_gnd g_1224((~pipeUNK09_v[`W-1]|~notRdy0_v[`W-1]), n781_v, n781_i3);
  spice_transistor_nmos_gnd g_1550((~n163_v[`W-1]&~n1253_v[`W-1]), n1184_v, n1184_i3);
  spice_transistor_nmos_gnd t2808(~n1211_v[`W-1], n1655_v, n1655_i0);
  spice_transistor_nmos_gnd g_1557((~n336_v[`W-1]&~n803_v[`W-1]), __AxB_6_v, __AxB_6_i4);
  spice_transistor_nmos t2747(~dpc37_PCLDB_v[`W-1], idb7_v, n1647_v, idb7_i8, n1647_i2);
  spice_transistor_nmos g_1559((~ADH_ABH_v[`W-1]&~cp1_v[`W-1]), _ABH6_v, n880_v, _ABH6_i2, n880_i2);
  spice_transistor_nmos t1802(~cclk_v[`W-1], pipeUNK35_v, n501_v, pipeUNK35_i0, n501_i0);
  spice_transistor_nmos t1801(~cp1_v[`W-1], notRdy0_v, n1276_v, notRdy0_i7, n1276_i0);
  spice_transistor_nmos_gnd t1806(~t2_v[`W-1], op_T2_v, op_T2_i0);
  spice_transistor_nmos_gnd t711(~n1529_v[`W-1], n91_v, n91_i0);
  spice_transistor_nmos t713(~cp1_v[`W-1], n854_v, n1395_v, n854_i0, n1395_i0);
  spice_transistor_nmos_vdd t2598(~cclk_v[`W-1], idb6_v, idb6_i8);
  spice_transistor_nmos_gnd t2049(~n1455_v[`W-1], n1412_v, n1412_i0);
  spice_transistor_nmos_gnd g_1314((~n1357_v[`W-1]|~n1606_v[`W-1]), n188_v, n188_i3);
  spice_transistor_nmos_gnd g_1311((~n152_v[`W-1]|~notRdy0_v[`W-1]), n1343_v, n1343_i1);
  spice_transistor_nmos t2042(~cp1_v[`W-1], n1039_v, n24_v, n1039_i0, n24_i0);
  spice_transistor_nmos_gnd t2040(~n196_v[`W-1], dpc5_SADL_v, dpc5_SADL_i7);
  spice_transistor_nmos t2047(~cclk_v[`W-1], n993_v, n20_v, n993_i0, n20_i0);
  spice_transistor_nmos_gnd g_1441((~n715_v[`W-1]&~n1316_v[`W-1]), n1386_v, n1386_i1);
  spice_transistor_nmos t2045(~cclk_v[`W-1], n1101_v, n190_v, n1101_i0, n190_i1);
  spice_transistor_nmos_gnd t2044(~op_rti_rts_v[`W-1], n1377_v, n1377_i0);
  spice_transistor_nmos t2919(~cclk_v[`W-1], _ABH5_v, n869_v, _ABH5_i1, n869_i3);
  spice_transistor_nmos t2918(~dpc33_PCHDB_v[`W-1], idb7_v, n1206_v, idb7_i9, n1206_i3);
  spice_transistor_nmos t2915(~dpc33_PCHDB_v[`W-1], n27_v, idb4_v, n27_i3, idb4_i8);
  spice_transistor_nmos t2914(~dpc33_PCHDB_v[`W-1], n141_v, idb3_v, n141_i3, idb3_i10);
  spice_transistor_nmos t2917(~dpc33_PCHDB_v[`W-1], idb6_v, n652_v, idb6_i10, n652_i3);
  spice_transistor_nmos_gnd t2128(~db6_v[`W-1], n374_v, n374_i1);
  spice_transistor_nmos t2911(~dpc33_PCHDB_v[`W-1], n1722_v, idb0_v, n1722_i3, idb0_i10);
  spice_transistor_nmos t2913(~dpc33_PCHDB_v[`W-1], idb2_v, n1496_v, idb2_i9, n1496_i3);
  spice_transistor_nmos t2912(~dpc33_PCHDB_v[`W-1], idb1_v, n209_v, idb1_i8, n209_i3);
  spice_transistor_nmos t478(~cclk_v[`W-1], DC78_phi2_v, DC78_v, DC78_phi2_i0, DC78_i0);
  spice_transistor_nmos_gnd g_1294((~clearIR_v[`W-1]|~pd6_v[`W-1]), pd6_clearIR_v, pd6_clearIR_i2);
  spice_transistor_nmos_gnd g_1445((~n743_v[`W-1]&~n1488_v[`W-1]), n609_v, n609_i2);
  spice_transistor_nmos_gnd g_1041((~ir4_v[`W-1]|~clock1_v[`W-1]|~ir2_v[`W-1]|~notir5_v[`W-1]|~ir6_v[`W-1]|~ir3_v[`W-1]|~irline3_v[`W-1]|~ir7_v[`W-1]), op_T0_jsr_v, op_T0_jsr_i1);
  spice_transistor_nmos_gnd g_1178((~pipeUNK33_v[`W-1]|~pipeUNK32_v[`W-1]|~pipeUNK31_v[`W-1]|~pipeUNK30_v[`W-1]), n1178_v, n1178_i2);
  spice_transistor_nmos_gnd g_1177((~n43_v[`W-1]|~n521_v[`W-1]), n6_v, n6_i3);
  spice_transistor_nmos_gnd g_1176((~n43_v[`W-1]|~n805_v[`W-1]), n1534_v, n1534_i3);
  spice_transistor_nmos t473(~cclk_v[`W-1], n207_v, n1061_v, n207_i0, n1061_i1);
  spice_transistor_nmos_gnd t475(~rdy_v[`W-1], n958_v, n958_i0);
  spice_transistor_nmos_gnd t477(~n1240_v[`W-1], dpc43_DL_DB_v, dpc43_DL_DB_i0);
  spice_transistor_nmos_gnd g_1170((~n467_v[`W-1]|~n630_v[`W-1]), n1705_v, n1705_i2);
  spice_transistor_nmos t1653(~cp1_v[`W-1], n1368_v, n1149_v, n1368_i0, n1149_i0);
  spice_transistor_nmos_gnd t2623(~alu5_v[`W-1], n761_v, n761_i1);
  spice_transistor_nmos_vdd t2622(~n1153_v[`W-1], n659_v, n659_i2);
  spice_transistor_nmos_gnd t679(~ir6_v[`W-1], _op_branch_bit6_v, _op_branch_bit6_i0);
  spice_transistor_nmos_gnd g_1488((~op_shift_v[`W-1]&~n440_v[`W-1]), n905_v, n905_i2);
  spice_transistor_nmos_gnd g_1487((~alua1_v[`W-1]&~alub1_v[`W-1]), aluanandb1_v, aluanandb1_i4);
  spice_transistor_nmos_gnd t900(~aluanorb1_v[`W-1], aluaorb1_v, aluaorb1_i0);
  spice_transistor_nmos_gnd g_1485((~n1440_v[`W-1]&(~n1081_v[`W-1]|~op_T0_sbc_v[`W-1]|~n1002_v[`W-1])), n779_v, n779_i2);
  spice_transistor_nmos_gnd t905(~n635_v[`W-1], ab14_v, ab14_i1);
  spice_transistor_nmos_gnd g_1482((~_DA_ADD1_v[`W-1]&~_DA_ADD2_v[`W-1]), n986_v, n986_i1);
  spice_transistor_nmos_gnd g_1481((~aluaorb0_v[`W-1]&~aluanandb0_v[`W-1]), __AxB_0_v, __AxB_0_i3);
  spice_transistor_nmos_gnd g_1480((~n647_v[`W-1]&~DA_C45_v[`W-1]), n757_v, n757_i1);
  spice_transistor_nmos_gnd g_1040((~ir3_v[`W-1]|~notir4_v[`W-1]|~notir0_v[`W-1]|~t3_v[`W-1]|~ir2_v[`W-1]), op_T3_ind_y_v, op_T3_ind_y_i1);
  spice_transistor_nmos t1652(~cclk_v[`W-1], n31_v, pipeUNK16_v, n31_i2, pipeUNK16_i0);
  spice_transistor_nmos_gnd g_1136((~n732_v[`W-1]|~n964_v[`W-1]), n17_v, n17_i4);
  spice_transistor_nmos_gnd t3188(~notidl1_v[`W-1], idl1_v, idl1_i1);
  spice_transistor_nmos_gnd t2455(~abh1_v[`W-1], n676_v, n676_i2);
  spice_transistor_nmos_gnd t2822(~a1_v[`W-1], n1549_v, n1549_i1);
  spice_transistor_nmos t2825(~cclk_v[`W-1], n1602_v, n506_v, n1602_i1, n506_i0);
  spice_transistor_nmos t2824(~cp1_v[`W-1], n1650_v, n94_v, n1650_i1, n94_i1);
  spice_transistor_nmos_gnd t2827(~n249_v[`W-1], n163_v, n163_i0);
  spice_transistor_nmos_gnd t2826(~n770_v[`W-1], n853_v, n853_i0);
  spice_transistor_nmos_gnd t875(~n599_v[`W-1], dpc22__DSA_v, dpc22__DSA_i0);
  spice_transistor_nmos_vdd t877(~n692_v[`W-1], dpc1_SBY_v, dpc1_SBY_i2);
  spice_transistor_nmos_gnd t876(~n692_v[`W-1], n441_v, n441_i0);
  spice_transistor_nmos_vdd t870(~n291_v[`W-1], dpc41_DL_ADL_v, dpc41_DL_ADL_i0);
  spice_transistor_nmos_gnd t873(~n278_v[`W-1], n1488_v, n1488_i0);
  spice_transistor_nmos t2139(~cclk_v[`W-1], n952_v, n1509_v, n952_i1, n1509_i0);
  spice_transistor_nmos t1986(~cclk_v[`W-1], n11_v, n55_v, n11_i0, n55_i0);
  spice_transistor_nmos_vdd t1118(~cclk_v[`W-1], sb3_v, sb3_i3);
  spice_transistor_nmos_vdd t3016(~n1034_v[`W-1], n994_v, n994_i3);
  spice_transistor_nmos t1114(~cp1_v[`W-1], n1376_v, notdor2_v, n1376_i0, notdor2_i1);
  spice_transistor_nmos t1117(~cclk_v[`W-1], n34_v, nots3_v, n34_i0, nots3_i0);
  spice_transistor_nmos t1110(~dpc17_SUMS_v[`W-1], __AxBxC_4_v, n296_v, __AxBxC_4_i0, n296_i1);
  spice_transistor_nmos t1111(~dpc17_SUMS_v[`W-1], __AxBxC_5_v, n277_v, __AxBxC_5_i0, n277_i2);
  spice_transistor_nmos t1112(~dpc17_SUMS_v[`W-1], n722_v, __AxBxC_6_v, n722_i2, __AxBxC_6_i0);
  spice_transistor_nmos t1113(~dpc17_SUMS_v[`W-1], n304_v, __AxBxC_7_v, n304_i2, __AxBxC_7_i0);
  spice_transistor_nmos_gnd t974(~_ABL0_v[`W-1], abl0_v, abl0_i3);
  spice_transistor_nmos t1333(~H1x1_v[`W-1], Pout1_v, idb1_v, Pout1_i0, idb1_i2);
  spice_transistor_nmos_gnd t3236(~n865_v[`W-1], n420_v, n420_i1);
  spice_transistor_nmos_gnd t495(~pd3_clearIR_v[`W-1], n1083_v, n1083_i0);
  spice_transistor_nmos_gnd t492(~n670_v[`W-1], n747_v, n747_i0);
  spice_transistor_nmos_gnd t491(~adh6_v[`W-1], n880_v, n880_i0);
  spice_transistor_nmos t490(~dpc7_SS_v[`W-1], s7_v, n721_v, s7_i0, n721_i1);
  spice_transistor_nmos_gnd g_1169((~notir6_v[`W-1]|~notir7_v[`W-1]|~ir4_v[`W-1]|~irline3_v[`W-1]|~clock1_v[`W-1]|~notir5_v[`W-1]), op_T0_cpx_inx_v, op_T0_cpx_inx_i1);
  spice_transistor_nmos_gnd t2012(~n1323_v[`W-1], dpc37_PCLDB_v, dpc37_PCLDB_i4);
  spice_transistor_nmos t499(~dpc13_ORS_v[`W-1], n722_v, n1084_v, n722_i0, n1084_i0);
  spice_transistor_nmos t1507(~cclk_v[`W-1], n146_v, a0_v, n146_i0, a0_i0);
  spice_transistor_nmos t3181(~dpc27_SBADH_v[`W-1], adh5_v, sb5_v, adh5_i5, sb5_i11);
  spice_transistor_nmos t1505(~dpc0_YSB_v[`W-1], n1491_v, sb2_v, n1491_i2, sb2_i3);
  spice_transistor_nmos_gnd g_1395((~n861_v[`W-1]|~notRdy0_v[`W-1]), brk_done_v, brk_done_i8);
  spice_transistor_nmos_gnd t2016(~idb7_v[`W-1], DBNeg_v, DBNeg_i0);
  spice_transistor_nmos t1752(~cp1_v[`W-1], n1014_v, idl6_v, n1014_i3, idl6_i1);
  spice_transistor_nmos_gnd t1503(~pipeVectorA2_v[`W-1], n815_v, n815_i0);
  spice_transistor_nmos_vdd t1750(~cclk_v[`W-1], adl2_v, adl2_i4);
  spice_transistor_nmos t1751(~cclk_v[`W-1], n1402_v, pchp2_v, n1402_i0, pchp2_i1);
  spice_transistor_nmos_gnd t1756(~n1533_v[`W-1], clock2_v, clock2_i0);
  spice_transistor_nmos_vdd t1757(~n373_v[`W-1], db5_v, db5_i3);
  spice_transistor_nmos t3373(~dpc40_ADLPCL_v[`W-1], pcl1_v, adl1_v, pcl1_i2, adl1_i8);
  spice_transistor_nmos t3180(~dpc39_PCLPCL_v[`W-1], pcl2_v, n481_v, pcl2_i1, n481_i3);
  spice_transistor_nmos_gnd g_1202((~pipeUNK20_v[`W-1]|~n430_v[`W-1]), n959_v, n959_i2);
  spice_transistor_nmos_gnd g_1205((~dor2_v[`W-1]|~RnWstretched_v[`W-1]), n224_v, n224_i2);
  spice_transistor_nmos_gnd g_1204((~n10_v[`W-1]|~n236_v[`W-1]), n176_v, n176_i2);
  spice_transistor_nmos_gnd t1687(~op_xy_v[`W-1], n1244_v, n1244_i0);
  spice_transistor_nmos_gnd g_1207((~n347_v[`W-1]|~_op_store_v[`W-1]), n335_v, n335_i1);
  spice_transistor_nmos_gnd g_1206((~VEC0_v[`W-1]|~VEC1_v[`W-1]), _VEC_v, _VEC_i3);
  spice_transistor_nmos_gnd g_1209((~n1247_v[`W-1]|~cclk_v[`W-1]|~n1043_v[`W-1]), dpc40_ADLPCL_v, dpc40_ADLPCL_i9);
  spice_transistor_nmos_gnd t3427(~n649_v[`W-1], A_B3_v, A_B3_i0);
  spice_transistor_nmos_gnd t3420(~notRdy0_v[`W-1], n1440_v, n1440_i0);
  spice_transistor_nmos_gnd g_1053((~notir3_v[`W-1]|~ir4_v[`W-1]|~notir7_v[`W-1]|~ir2_v[`W-1]|~irline3_v[`W-1]|~ir5_v[`W-1]|~clock1_v[`W-1]), op_T0_iny_dey_v, op_T0_iny_dey_i1);
  spice_transistor_nmos_gnd t272(~n1575_v[`W-1], t2_v, t2_i0);
  spice_transistor_nmos_vdd t276(~n631_v[`W-1], dpc37_PCLDB_v, dpc37_PCLDB_i0);
  spice_transistor_nmos_gnd t275(~n631_v[`W-1], n1323_v, n1323_i0);
  spice_transistor_nmos_gnd g_1536((~dpc35_PCHC_v[`W-1]&~n83_v[`W-1]), n523_v, n523_i3);
  spice_transistor_nmos_vdd t279(~cclk_v[`W-1], adl4_v, adl4_i0);
  spice_transistor_nmos_gnd t2759(~pcl2_v[`W-1], n783_v, n783_i0);
  spice_transistor_nmos_gnd g_1056((~n979_v[`W-1]|~n550_v[`W-1]|~op_T0_shift_a_v[`W-1]|~nnT2BR_v[`W-1]|~n862_v[`W-1]|~n782_v[`W-1]), n1347_v, n1347_i2);
  spice_transistor_nmos_gnd t92(~n381_v[`W-1], ab8_v, ab8_i1);
  spice_transistor_nmos_gnd g_1057((~notRdy0_v[`W-1]|~n992_v[`W-1]), n46_v, n46_i1);
  spice_transistor_nmos_gnd t2101(~n171_v[`W-1], ab7_v, ab7_i1);
  spice_transistor_nmos_gnd t1949(~n94_v[`W-1], n1024_v, n1024_i0);
  spice_transistor_nmos_gnd t2458(~abh7_v[`W-1], n1153_v, n1153_i0);
  spice_transistor_nmos_gnd t1947(~n849_v[`W-1], dpc33_PCHDB_v, dpc33_PCHDB_i1);
  spice_transistor_nmos_gnd t3183(~adh5_v[`W-1], n254_v, n254_i0);
  spice_transistor_nmos t3182(~dpc5_SADL_v[`W-1], n618_v, adl6_v, n618_i2, adl6_i5);
  spice_transistor_nmos_gnd t3184(~n336_v[`W-1], n1038_v, n1038_i0);
  spice_transistor_nmos_gnd t1946(~n1411_v[`W-1], pclp2_v, pclp2_i1);
  spice_transistor_nmos t2450(~dpc30_ADHPCH_v[`W-1], pch1_v, adh1_v, pch1_i1, adh1_i5);
  spice_transistor_nmos t2451(~cp1_v[`W-1], n590_v, n1178_v, n590_i0, n1178_i0);
  spice_transistor_nmos_gnd t2452(~_ABH5_v[`W-1], abh5_v, abh5_i3);
  spice_transistor_nmos t2453(~dpc30_ADHPCH_v[`W-1], pch0_v, adh0_v, pch0_i1, adh0_i4);
  spice_transistor_nmos_gnd t2454(~abh1_v[`W-1], n617_v, n617_i0);
  spice_transistor_nmos_gnd t1945(~y3_v[`W-1], n184_v, n184_i0);
  spice_transistor_nmos t2456(~cclk_v[`W-1], pchp6_v, n1192_v, pchp6_i1, n1192_i0);
  spice_transistor_nmos_vdd t2457(~abh7_v[`W-1], n1639_v, n1639_i0);
  spice_transistor_nmos_gnd t3473(~n1072_v[`W-1], db0_v, db0_i3);
  spice_transistor_nmos_gnd t1944(~op_T5_jsr_v[`W-1], n1219_v, n1219_i1);
  spice_transistor_nmos_gnd t1943(~n1574_v[`W-1], n1089_v, n1089_i1);
  spice_transistor_nmos_gnd g_1059((~n1252_v[`W-1]|~n597_v[`W-1]), n882_v, n882_i1);
  spice_transistor_nmos_gnd t1942(~clk0_v[`W-1], n519_v, n519_i1);
  spice_transistor_nmos t1941(~cp1_v[`W-1], n644_v, n428_v, n644_i0, n428_i0);
  spice_transistor_nmos_gnd t1024(~n471_v[`W-1], db6_v, db6_i0);
  spice_transistor_nmos t2247(~cp1_v[`W-1], n1180_v, n1533_v, n1180_i0, n1533_i1);
  spice_transistor_nmos_gnd g_1567((~n311_v[`W-1]&~dpc34_PCLC_v[`W-1]), n919_v, n919_i3);
  spice_transistor_nmos_gnd g_1560(((~op_rol_ror_v[`W-1]|~op_T0_adc_sbc_v[`W-1])&~n1044_v[`W-1]), n1408_v, n1408_i2);
  spice_transistor_nmos_gnd g_1562(((~n410_v[`W-1]|~n392_v[`W-1])&~n344_v[`W-1]), n1073_v, n1073_i2);
  spice_transistor_nmos_gnd g_1563(((~n1581_v[`W-1]|~n1570_v[`W-1])&~n1472_v[`W-1]), dpc36_IPC_v, dpc36_IPC_i3);
  spice_transistor_nmos_gnd t1835(~idb6_v[`W-1], n1684_v, n1684_i1);
  spice_transistor_nmos_gnd t1834(~n503_v[`W-1], n270_v, n270_i0);
  spice_transistor_nmos t1833(~cp1_v[`W-1], notRdy0_v, n1272_v, notRdy0_i8, n1272_i1);
  spice_transistor_nmos t705(~cclk_v[`W-1], n277_v, notalu5_v, n277_i0, notalu5_i0);
  spice_transistor_nmos_vdd t702(~abl2_v[`W-1], n1152_v, n1152_i0);
  spice_transistor_nmos_gnd t701(~abl2_v[`W-1], n951_v, n951_i0);
  spice_transistor_nmos_gnd t700(~abl2_v[`W-1], n642_v, n642_i0);
  spice_transistor_nmos_gnd t709(~idb6_v[`W-1], n351_v, n351_i0);
  spice_transistor_nmos_gnd t708(~AxB7_v[`W-1], n177_v, n177_i0);
  spice_transistor_nmos t3053(~cclk_v[`W-1], n632_v, n339_v, n632_i0, n339_i1);
  spice_transistor_nmos_gnd g_1363((~x_op_T4_rti_v[`W-1]|~op_T0_plp_v[`W-1]), n327_v, n327_i2);
  spice_transistor_nmos_gnd t2588(~nmi_v[`W-1], n1392_v, n1392_i1);
  spice_transistor_nmos t2589(~cclk_v[`W-1], n1699_v, n1024_v, n1699_i1, n1024_i1);
  spice_transistor_nmos_gnd t3057(~n1467_v[`W-1], cclk_v, cclk_i207);
  spice_transistor_nmos_gnd g_1367((~alub6_v[`W-1]|~alua6_v[`W-1]), n1084_v, n1084_i3);
  spice_transistor_nmos_vdd t3055(~n1364_v[`W-1], dpc16_EORS_v, dpc16_EORS_i9);
  spice_transistor_nmos_gnd t3054(~n1364_v[`W-1], n108_v, n108_i1);
  spice_transistor_nmos t2582(~cclk_v[`W-1], pipeT3out_v, n678_v, pipeT3out_i0, n678_i0);
  spice_transistor_nmos_gnd t2583(~pipeUNK22_v[`W-1], n533_v, n533_i1);
  spice_transistor_nmos_gnd g_1369((~notir1_v[`W-1]|~ir7_v[`W-1]|~notir6_v[`W-1]|~notir5_v[`W-1]), op_ror_v, op_ror_i2);
  spice_transistor_nmos_vdd t2586(~n1423_v[`W-1], n869_v, n869_i2);
  spice_transistor_nmos_gnd t2585(~n1423_v[`W-1], n1608_v, n1608_i2);
  spice_transistor_nmos t2909(~cclk_v[`W-1], n1379_v, pipeUNK10_v, n1379_i0, pipeUNK10_i0);
  spice_transistor_nmos_vdd t2902(~n830_v[`W-1], dpc23_SBAC_v, dpc23_SBAC_i8);
  spice_transistor_nmos_gnd t2900(~n902_v[`W-1], n1289_v, n1289_i0);
  spice_transistor_nmos_gnd t2901(~n830_v[`W-1], n1047_v, n1047_i0);
  spice_transistor_nmos_gnd t3350(~n310_v[`W-1], ir0_v, ir0_i1);
  spice_transistor_nmos_gnd g_1108((~ir3_v[`W-1]|~ir7_v[`W-1]|~irline3_v[`W-1]|~ir2_v[`W-1]|~ir4_v[`W-1]|~ir5_v[`W-1]), op_brk_rti_v, op_brk_rti_i2);
  spice_transistor_nmos_gnd t3351(~adh7_v[`W-1], n494_v, n494_i0);
  spice_transistor_nmos_gnd g_1102((~ir3_v[`W-1]|~ir7_v[`W-1]|~ir6_v[`W-1]|~ir4_v[`W-1]|~t2_v[`W-1]|~irline3_v[`W-1]|~ir2_v[`W-1]|~ir5_v[`W-1]), op_T2_brk_v, op_T2_brk_i1);
  spice_transistor_nmos_gnd g_1101((~n1247_v[`W-1]|~n763_v[`W-1]|~cclk_v[`W-1]), dpc8_nDBADD_v, dpc8_nDBADD_i9);
  spice_transistor_nmos_gnd g_1106((~notir6_v[`W-1]|~notir3_v[`W-1]|~ir7_v[`W-1]|~notir2_v[`W-1]|~clock1_v[`W-1]|~irline3_v[`W-1]|~ir4_v[`W-1]), op_T0_jmp_v, op_T0_jmp_i1);
  spice_transistor_nmos_vdd t3352(~cclk_v[`W-1], adh6_v, adh6_i6);
  spice_transistor_nmos_gnd g_1104((~notir6_v[`W-1]|~ir7_v[`W-1]|~ir3_v[`W-1]|~ir4_v[`W-1]|~irline3_v[`W-1]|~t5_v[`W-1]|~notir5_v[`W-1]|~ir2_v[`W-1]), op_T5_rts_v, op_T5_rts_i2);
  spice_transistor_nmos_gnd t2654(~a0_v[`W-1], n5_v, n5_i0);
  spice_transistor_nmos t2630(~cclk_v[`W-1], _op_set_C_v, pipeUNK08_v, _op_set_C_i0, pipeUNK08_i0);
  spice_transistor_nmos_gnd t2248(~s0_v[`W-1], n983_v, n983_i1);
  spice_transistor_nmos t2634(~cclk_v[`W-1], n306_v, n581_v, n306_i1, n581_i1);
  spice_transistor_nmos_gnd t2635(~n1157_v[`W-1], dpc41_DL_ADL_v, dpc41_DL_ADL_i9);
  spice_transistor_nmos_gnd t2637(~notdor5_v[`W-1], dor5_v, dor5_i1);
  spice_transistor_nmos_gnd t3357(~n184_v[`W-1], n1531_v, n1531_i2);
  spice_transistor_nmos t1349(~cclk_v[`W-1], n396_v, n796_v, n396_i0, n796_i0);
  spice_transistor_nmos_vdd t1344(~n1715_v[`W-1], n1105_v, n1105_i0);
  spice_transistor_nmos_gnd t1347(~pcl1_v[`W-1], n329_v, n329_i0);
  spice_transistor_nmos_gnd t1346(~y4_v[`W-1], n565_v, n565_i0);
  spice_transistor_nmos_gnd t1341(~dpc12_0ADD_v[`W-1], alua7_v, alua7_i0);
  spice_transistor_nmos_gnd t1340(~alu6_v[`W-1], n149_v, n149_i0);
  spice_transistor_nmos_gnd t1342(~n1715_v[`W-1], n1399_v, n1399_i0);
  spice_transistor_nmos_gnd g_1151((~irline3_v[`W-1]|~notir4_v[`W-1]|~ir2_v[`W-1]|~ir3_v[`W-1]|~t3_v[`W-1]), op_T3_branch_v, op_T3_branch_i3);
  spice_transistor_nmos_gnd g_1617(((~x_op_T0_tya_v[`W-1]|~op_T2_abs_y_v[`W-1]|~op_T0_iny_dey_v[`W-1]|~op_T0_cpy_iny_v[`W-1]|~op_T3_ind_y_v[`W-1])|(~n335_v[`W-1]&~op_sty_cpy_mem_v[`W-1])|(~op_T2_idx_x_xy_v[`W-1]&~op_xy_v[`W-1])), n1717_v, n1717_i2);
  spice_transistor_nmos_gnd g_1614(((~n440_v[`W-1]&~op_shift_right_v[`W-1])|~op_T0_shift_right_a_v[`W-1]), n366_v, n366_i2);
  spice_transistor_nmos_gnd g_1615((((~n1610_v[`W-1]|~n388_v[`W-1])&(~n319_v[`W-1]|~n1691_v[`W-1]))|~dpc18__DAA_v[`W-1]), DC34_v, DC34_i1);
  spice_transistor_nmos_gnd g_1612(((~AxB3_v[`W-1]&~_C23_v[`W-1])|~__AxB3__C23_v[`W-1]), __AxBxC_3_v, __AxBxC_3_i2);
  spice_transistor_nmos_gnd g_1613(((~pipeUNK17_v[`W-1]&~n553_v[`W-1])|(~n1573_v[`W-1]&~n781_v[`W-1])|(~n270_v[`W-1]&~n1662_v[`W-1])), n845_v, n845_i2);
  spice_transistor_nmos_gnd g_1610((~n743_v[`W-1]|(~n523_v[`W-1]&~n499_v[`W-1])), n875_v, n875_i2);
  spice_transistor_nmos_gnd g_1611((~n936_v[`W-1]|(~C01_v[`W-1]&~aluaorb1_v[`W-1])), _C12_v, _C12_i2);
  spice_transistor_nmos_gnd g_1618((~NMIP_v[`W-1]|(~n1392_v[`W-1]&~cclk_v[`W-1])), n297_v, n297_i1);
  spice_transistor_nmos_gnd g_1619((~_AxB_2__C12_v[`W-1]|(~C12_v[`W-1]&~__AxB_2_v[`W-1])), __AxBxC_2_v, __AxBxC_2_i2);
  spice_transistor_nmos_gnd g_1585((~alub4_v[`W-1]&~alua4_v[`W-1]), n1063_v, n1063_i4);
  spice_transistor_nmos_gnd g_1582(((~n715_v[`W-1]|~n1316_v[`W-1])&~n1386_v[`W-1]), n484_v, n484_i2);
  spice_transistor_nmos g_1580((~ADH_ABH_v[`W-1]&~cp1_v[`W-1]), _ABH0_v, n1668_v, _ABH0_i2, n1668_i2);
  spice_transistor_nmos_gnd t2126(~n1579_v[`W-1], n221_v, n221_i0);
  spice_transistor_nmos t2127(~H1x1_v[`W-1], Pout4_v, idb4_v, Pout4_i1, idb4_i4);
  spice_transistor_nmos_gnd t2120(~clk0_v[`W-1], n358_v, n358_i1);
  spice_transistor_nmos t2123(~dpc3_SBX_v[`W-1], x0_v, dasb0_v, x0_i0, dasb0_i7);
  spice_transistor_nmos_vdd t1169(~n519_v[`W-1], n135_v, n135_i1);
  spice_transistor_nmos_vdd t1699(~n543_v[`W-1], dpc5_SADL_v, dpc5_SADL_i0);
  spice_transistor_nmos_gnd t1698(~n543_v[`W-1], n196_v, n196_i0);
  spice_transistor_nmos_gnd t1161(~n236_v[`W-1], n79_v, n79_i0);
  spice_transistor_nmos t1160(~dpc8_nDBADD_v[`W-1], alub0_v, n624_v, alub0_i2, n624_i1);
  spice_transistor_nmos_gnd t1162(~C23_v[`W-1], _C23_v, _C23_i0);
  spice_transistor_nmos t1165(~dpc8_nDBADD_v[`W-1], alub2_v, n458_v, alub2_i0, n458_i1);
  spice_transistor_nmos t1164(~dpc8_nDBADD_v[`W-1], alub4_v, n478_v, alub4_i0, n478_i0);
  spice_transistor_nmos_gnd t3129(~irq_v[`W-1], n1599_v, n1599_i1);
  spice_transistor_nmos t1588(~cclk_v[`W-1], n722_v, notalu6_v, n722_i3, notalu6_i1);
  spice_transistor_nmos_vdd t1587(~cclk_v[`W-1], dasb0_v, dasb0_i4);
  spice_transistor_nmos t1583(~cclk_v[`W-1], n559_v, n608_v, n559_i0, n608_i1);
  spice_transistor_nmos_gnd g_1343((~n180_v[`W-1]|~n819_v[`W-1]|~Reset0_v[`W-1]), n501_v, n501_i2);
  spice_transistor_nmos_gnd t1580(~pipedpc28_v[`W-1], dpc28_0ADH0_v, dpc28_0ADH0_i0);
  spice_transistor_nmos t1767(~cclk_v[`W-1], pclp1_v, n1099_v, pclp1_i0, n1099_i0);
  spice_transistor_nmos t1766(~cclk_v[`W-1], n1130_v, n512_v, n1130_i0, n512_i1);
  spice_transistor_nmos t1765(~cclk_v[`W-1], n674_v, n745_v, n674_i1, n745_i0);
  spice_transistor_nmos_gnd t1762(~n761_v[`W-1], n1056_v, n1056_i0);
  spice_transistor_nmos_vdd t1760(~cclk_v[`W-1], idb2_v, idb2_i4);
  spice_transistor_nmos_gnd t1566(~n128_v[`W-1], n1592_v, n1592_i1);
  spice_transistor_nmos_gnd t1561(~n210_v[`W-1], ab5_v, ab5_i0);
  spice_transistor_nmos_vdd t3149(~abl4_v[`W-1], n634_v, n634_i1);
  spice_transistor_nmos_gnd g_1154((~pipeUNK23_v[`W-1]|~pipephi2Reset0_v[`W-1]), n819_v, n819_i2);
  spice_transistor_nmos_gnd g_1157((~n1038_v[`W-1]|~AxB7_v[`W-1]), n269_v, n269_i1);
  spice_transistor_nmos_gnd g_1156((~nnT2BR_v[`W-1]|~n847_v[`W-1]|~n440_v[`W-1]|~n275_v[`W-1]|~op_T4_jmp_v[`W-1]), n104_v, n104_i2);
  spice_transistor_nmos_gnd t3148(~abl4_v[`W-1], n1676_v, n1676_i2);
  spice_transistor_nmos_gnd g_1150((~notir7_v[`W-1]|~clock1_v[`W-1]|~notir5_v[`W-1]|~ir6_v[`W-1]|~notir0_v[`W-1]), op_T0_lda_v, op_T0_lda_i2);
  spice_transistor_nmos_gnd g_1153((~RnWstretched_v[`W-1]|~dor4_v[`W-1]), n1463_v, n1463_i2);
  spice_transistor_nmos_gnd g_1152((~notir4_v[`W-1]|~irline3_v[`W-1]|~t2_v[`W-1]|~ir3_v[`W-1]|~ir2_v[`W-1]), op_T2_branch_v, op_T2_branch_i2);
  spice_transistor_nmos_vdd t1956(~n1230_v[`W-1], dpc11_SBADD_v, dpc11_SBADD_i7);
  spice_transistor_nmos t2115(~cp1_v[`W-1], n1718_v, n671_v, n1718_i0, n671_i0);
  spice_transistor_nmos t1957(~dpc13_ORS_v[`W-1], n304_v, n1398_v, n304_i3, n1398_i0);
  spice_transistor_nmos_gnd t3015(~n1034_v[`W-1], n1545_v, n1545_i2);
  spice_transistor_nmos t248(~dpc6_SBS_v[`W-1], s5_v, sb5_v, s5_i0, sb5_i1);
  spice_transistor_nmos t249(~dpc6_SBS_v[`W-1], s6_v, sb6_v, s6_i0, sb6_i3);
  spice_transistor_nmos t242(~cclk_v[`W-1], n1117_v, pipeVectorA1_v, n1117_i0, pipeVectorA1_i0);
  spice_transistor_nmos t243(~cp1_v[`W-1], n797_v, notdor4_v, n797_i0, notdor4_i0);
  spice_transistor_nmos t241(~cclk_v[`W-1], n326_v, a6_v, n326_i0, a6_i0);
  spice_transistor_nmos_gnd t695(~n551_v[`W-1], n8_v, n8_i0);
  spice_transistor_nmos_gnd g_1158((~n1055_v[`W-1]|~op_T0_cpx_cpy_inx_iny_v[`W-1]|~op_T0_cmp_v[`W-1]), n1560_v, n1560_i2);
  spice_transistor_nmos_vdd t694(~n567_v[`W-1], n322_v, n322_i1);
  spice_transistor_nmos t925(~cp1_v[`W-1], n626_v, n756_v, n626_i0, n756_i0);
  spice_transistor_nmos_gnd t2681(~a3_v[`W-1], n947_v, n947_i1);
  spice_transistor_nmos t696(~cclk_v[`W-1], n1620_v, notir3_v, n1620_i0, notir3_i1);
  spice_transistor_nmos_gnd g_1479(((~n1345_v[`W-1]|~n1166_v[`W-1])&~n1542_v[`W-1]), n1099_v, n1099_i2);
  spice_transistor_nmos t527(~dpc21_ADDADL_v[`W-1], adl5_v, alu5_v, adl5_i1, alu5_i0);
  spice_transistor_nmos_gnd t398(~dpc29_0ADH17_v[`W-1], adh1_v, adh1_i1);
  spice_transistor_nmos t2943(~cp1_v[`W-1], n1474_v, notdor1_v, n1474_i1, notdor1_i1);
  spice_transistor_nmos_gnd t390(~notRdy0_v[`W-1], n16_v, n16_i0);
  spice_transistor_nmos_gnd t391(~db1_v[`W-1], n213_v, n213_i0);
  spice_transistor_nmos_gnd t392(~pipeVectorA1_v[`W-1], n_0_ADL1_v, n_0_ADL1_i0);
  spice_transistor_nmos_gnd t393(~nots5_v[`W-1], n280_v, n280_i2);
  spice_transistor_nmos t394(~cclk_v[`W-1], n1654_v, a3_v, n1654_i0, a3_i0);
  spice_transistor_nmos_vdd t397(~n317_v[`W-1], n417_v, n417_i1);
  spice_transistor_nmos_gnd t2110(~op_T0_cli_sei_v[`W-1], n1065_v, n1065_i1);
  spice_transistor_nmos t2532(~dpc38_PCLADL_v[`W-1], n723_v, adl3_v, n723_i1, adl3_i4);
  spice_transistor_nmos_gnd g_1063((~op_T0_ora_v[`W-1]|~notRdy0_v[`W-1]), n1145_v, n1145_i2);
  spice_transistor_nmos_gnd t3193(~n837_v[`W-1], op_EORS_v, op_EORS_i1);
  spice_transistor_nmos_gnd t3196(~idb7_v[`W-1], n423_v, n423_i1);
  spice_transistor_nmos t3197(~cclk_v[`W-1], pipeUNK02_v, n774_v, pipeUNK02_i1, n774_i1);
  spice_transistor_nmos_gnd t3194(~n590_v[`W-1], alucin_v, alucin_i1);
  spice_transistor_nmos_vdd t1991(~n23_v[`W-1], n1501_v, n1501_i1);
  spice_transistor_nmos t3198(~cclk_v[`W-1], op_SRS_v, n968_v, op_SRS_i3, n968_i1);
  spice_transistor_nmos t3199(~cclk_v[`W-1], op_SUMS_v, n415_v, op_SUMS_i0, n415_i1);
  spice_transistor_nmos_gnd t3466(~D1x1_v[`W-1], n1471_v, n1471_i1);
  spice_transistor_nmos_gnd t3467(~n386_v[`W-1], n392_v, n392_i0);
  spice_transistor_nmos t3469(~cclk_v[`W-1], n700_v, n1565_v, n700_i1, n1565_i1);
  spice_transistor_nmos_gnd t2112(~x1_v[`W-1], n1434_v, n1434_i0);
  spice_transistor_nmos_gnd t1992(~n968_v[`W-1], n1093_v, n1093_i1);
  spice_transistor_nmos_gnd g_1579((~C34_v[`W-1]&~n700_v[`W-1]), n695_v, n695_i2);
  spice_transistor_nmos t3454(~cclk_v[`W-1], n1649_v, n1027_v, n1649_i1, n1027_i0);
  spice_transistor_nmos_gnd g_1574((~n462_v[`W-1]&~n824_v[`W-1]), n1642_v, n1642_i2);
  spice_transistor_nmos_gnd t1828(~y7_v[`W-1], n1640_v, n1640_i0);
  spice_transistor_nmos t1829(~cclk_v[`W-1], n119_v, notir1_v, n119_i0, notir1_i1);
  spice_transistor_nmos t1993(~cclk_v[`W-1], n1705_v, n1020_v, n1705_i0, n1020_i1);
  spice_transistor_nmos_gnd t2231(~n31_v[`W-1], n132_v, n132_i1);
  spice_transistor_nmos t1823(~cp1_v[`W-1], n1360_v, n1091_v, n1360_i0, n1091_i0);
  spice_transistor_nmos_gnd t1825(~n1679_v[`W-1], n1262_v, n1262_i0);
  spice_transistor_nmos t1826(~cclk_v[`W-1], pipeUNK41_v, n504_v, pipeUNK41_i0, n504_i0);
  spice_transistor_nmos t1827(~cclk_v[`W-1], op_ANDS_v, n1574_v, op_ANDS_i0, n1574_i0);
  spice_transistor_nmos_gnd t2029(~n878_v[`W-1], n631_v, n631_i2);
  spice_transistor_nmos_vdd t2028(~cclk_v[`W-1], adh7_v, adh7_i2);
  spice_transistor_nmos_gnd g_1371((~n1247_v[`W-1]|~n969_v[`W-1]|~cclk_v[`W-1]), dpc0_YSB_v, dpc0_YSB_i9);
  spice_transistor_nmos_gnd g_1372((~n673_v[`W-1]|~op_T0_sbc_v[`W-1]), n1304_v, n1304_i2);
  spice_transistor_nmos_gnd t3049(~n993_v[`W-1], pclp6_v, pclp6_i0);
  spice_transistor_nmos_gnd g_1379((~notir6_v[`W-1]|~notir1_v[`W-1]|~ir7_v[`W-1]), op_shift_right_v, op_shift_right_i1);
  spice_transistor_nmos_gnd t3046(~idb2_v[`W-1], n1376_v, n1376_i1);
  spice_transistor_nmos_gnd t3047(~PD_0xx0xx0x_v[`W-1], PD_n_0xx0xx0x_v, PD_n_0xx0xx0x_i0);
  spice_transistor_nmos_gnd t1755(~n905_v[`W-1], n979_v, n979_i0);
  spice_transistor_nmos_gnd g_1146((~notir0_v[`W-1]|~ir6_v[`W-1]|~notir7_v[`W-1]|~ir5_v[`W-1]), op_sta_cmp_v, op_sta_cmp_i1);
  spice_transistor_nmos t2930(~cclk_v[`W-1], n104_v, n1221_v, n104_i0, n1221_i1);
  spice_transistor_nmos_gnd g_1110((~notir6_v[`W-1]|~ir7_v[`W-1]|~notir3_v[`W-1]|~notir2_v[`W-1]|~ir4_v[`W-1]|~irline3_v[`W-1]), x_op_jmp_v, x_op_jmp_i3);
  spice_transistor_nmos_gnd g_1115((~cclk_v[`W-1]|~n962_v[`W-1]), _DBE_v, _DBE_i1);
  spice_transistor_nmos_gnd g_1114((~n1054_v[`W-1]|~_VEC_v[`W-1]), n70_v, n70_i2);
  spice_transistor_nmos_gnd g_1117((~n1149_v[`W-1]|~n1312_v[`W-1]), n264_v, n264_i3);
  spice_transistor_nmos_gnd g_1116((~n440_v[`W-1]|~n646_v[`W-1]), n812_v, n812_i1);
  spice_transistor_nmos_gnd g_1147((~n383_v[`W-1]|~notRdy0_v[`W-1]), n917_v, n917_i2);
  spice_transistor_nmos t2483(~cclk_v[`W-1], n515_v, n1411_v, n515_i0, n1411_i1);
  spice_transistor_nmos t2482(~dpc31_PCHPCH_v[`W-1], pch1_v, n209_v, pch1_i2, n209_i0);
  spice_transistor_nmos t2481(~dpc31_PCHPCH_v[`W-1], pch0_v, n1722_v, pch0_i2, n1722_i1);
  spice_transistor_nmos t2480(~dpc31_PCHPCH_v[`W-1], pch3_v, n141_v, pch3_i2, n141_i1);
  spice_transistor_nmos_gnd t2339(~nots0_v[`W-1], n332_v, n332_i2);
  spice_transistor_nmos_gnd t2485(~dpc29_0ADH17_v[`W-1], adh3_v, adh3_i5);
  spice_transistor_nmos t2334(~dpc37_PCLDB_v[`W-1], idb4_v, n208_v, idb4_i6, n208_i1);
  spice_transistor_nmos_vdd t2336(~cclk_v[`W-1], adh3_v, adh3_i4);
  spice_transistor_nmos_gnd t2331(~n581_v[`W-1], n838_v, n838_i0);
  spice_transistor_nmos_gnd t2119(~_ABH0_v[`W-1], abh0_v, abh0_i3);
  spice_transistor_nmos_gnd t2803(~n958_v[`W-1], n1449_v, n1449_i0);
  spice_transistor_nmos_gnd t2802(~n927_v[`W-1], ir4_v, ir4_i0);
  spice_transistor_nmos_gnd g_1460((~n761_v[`W-1]&~n149_v[`W-1]), n233_v, n233_i1);
  spice_transistor_nmos_gnd t1352(~n1380_v[`W-1], n109_v, n109_i0);
  spice_transistor_nmos t1350(~cclk_v[`W-1], _ABL0_v, n1100_v, _ABL0_i1, n1100_i2);
  spice_transistor_nmos_gnd g_1605(((~n1511_v[`W-1]&~pipeUNK28_v[`W-1])|(~pipeUNK29_v[`W-1]&~n1714_v[`W-1])), n262_v, n262_i2);
  spice_transistor_nmos_gnd g_1604((~n1619_v[`W-1]|(~nnT2BR_v[`W-1]&~BRtaken_v[`W-1])), n586_v, n586_i2);
  spice_transistor_nmos_gnd g_1607((~n330_v[`W-1]|(~cclk_v[`W-1]&~n1599_v[`W-1])), n807_v, n807_i1);
  spice_transistor_nmos_gnd g_1606(((~notalucin_v[`W-1]&~aluanandb0_v[`W-1])|~aluanorb0_v[`W-1]), C01_v, C01_i2);
  spice_transistor_nmos_gnd g_1601((((~n757_v[`W-1]|~__AxB_6_v[`W-1])&(~n570_v[`W-1]|~n269_v[`W-1]))|~dpc18__DAA_v[`W-1]), DC78_v, DC78_i2);
  spice_transistor_nmos_gnd g_1603(((~AxB1_v[`W-1]&~_C01_v[`W-1])|~__AxB1__C01_v[`W-1]), __AxBxC_1_v, __AxBxC_1_i2);
  spice_transistor_nmos_gnd g_1602((~n1629_v[`W-1]|(~n1135_v[`W-1]&~n753_v[`W-1])), dasb5_v, dasb5_i2);
  spice_transistor_nmos g_1489((~cp1_v[`W-1]&~fetch_v[`W-1]), n1083_v, n1620_v, n1083_i4, n1620_i2);
  spice_transistor_nmos_gnd g_1609((~__AxB5__C45_v[`W-1]|(~_C45_v[`W-1]&~AxB5_v[`W-1])), __AxBxC_5_v, __AxBxC_5_i2);
  spice_transistor_nmos_gnd g_1608((~n50_v[`W-1]|((~n646_v[`W-1]|~nnT2BR_v[`W-1])&~n480_v[`W-1])), n629_v, n629_i2);
  spice_transistor_nmos_gnd g_1375((~AxB7_v[`W-1]|~_C67_v[`W-1]), __AxB7__C67_v, __AxB7__C67_i1);
  spice_transistor_nmos_gnd g_1597(((~n755_v[`W-1]&~_DBZ_v[`W-1])|(~n243_v[`W-1]&~n781_v[`W-1])|(~pipeUNK14_v[`W-1]&~n1170_v[`W-1])), n566_v, n566_i2);
  spice_transistor_nmos_gnd g_1590((~alub6_v[`W-1]&~alua6_v[`W-1]), n336_v, n336_i5);
  spice_transistor_nmos_gnd g_1593((~n609_v[`W-1]&(~n1488_v[`W-1]|~n743_v[`W-1])), n1192_v, n1192_i2);
  spice_transistor_nmos_gnd g_1598((~n1345_v[`W-1]|(~dpc36_IPC_v[`W-1]&~n937_v[`W-1])), n1500_v, n1500_i2);
  spice_transistor_nmos_gnd t1222(~n1675_v[`W-1], ir6_v, ir6_i2);
  spice_transistor_nmos t1227(~cclk_v[`W-1], n176_v, n598_v, n176_i0, n598_i0);
  spice_transistor_nmos_gnd t1225(~n384_v[`W-1], n885_v, n885_i0);
  spice_transistor_nmos t1228(~cclk_v[`W-1], n1592_v, a7_v, n1592_i0, a7_i1);
  spice_transistor_nmos_gnd t2154(~n69_v[`W-1], n1045_v, n1045_i2);
  spice_transistor_nmos_vdd t2157(~n417_v[`W-1], sync_v, sync_i1);
  spice_transistor_nmos_gnd t1178(~a7_v[`W-1], n128_v, n128_i0);
  spice_transistor_nmos_gnd t1176(~_ABL5_v[`W-1], abl5_v, abl5_i0);
  spice_transistor_nmos_gnd t2640(~notalu5_v[`W-1], alu5_v, alu5_i3);
  spice_transistor_nmos t1599(~dpc1_SBY_v[`W-1], y2_v, sb2_v, y2_i2, sb2_i6);
  spice_transistor_nmos t1590(~dpc14_SRS_v[`W-1], aluanandb1_v, notaluoutmux0_v, aluanandb1_i0, notaluoutmux0_i2);
  spice_transistor_nmos t1591(~dpc14_SRS_v[`W-1], notaluoutmux1_v, n681_v, notaluoutmux1_i2, n681_i0);
  spice_transistor_nmos t1592(~dpc14_SRS_v[`W-1], n350_v, n740_v, n350_i0, n740_i3);
  spice_transistor_nmos t1593(~dpc14_SRS_v[`W-1], n1071_v, n1063_v, n1071_i4, n1063_i0);
  spice_transistor_nmos t1594(~dpc14_SRS_v[`W-1], n296_v, n477_v, n296_i3, n477_i0);
  spice_transistor_nmos t1595(~dpc14_SRS_v[`W-1], n277_v, n336_v, n277_i3, n336_i0);
  spice_transistor_nmos t1596(~dpc14_SRS_v[`W-1], n722_v, n1318_v, n722_i4, n1318_i1);
  spice_transistor_nmos t1597(~cclk_v[`W-1], n469_v, n875_v, n469_i0, n875_i0);
  spice_transistor_nmos_gnd t1773(~n161_v[`W-1], n969_v, n969_i0);
  spice_transistor_nmos_vdd t1774(~n161_v[`W-1], dpc0_YSB_v, dpc0_YSB_i3);
  spice_transistor_nmos_gnd t1775(~n641_v[`W-1], n715_v, n715_i0);
  spice_transistor_nmos_gnd g_1404((~cclk_v[`W-1]|~n1247_v[`W-1]|~n602_v[`W-1]), dpc2_XSB_v, dpc2_XSB_i9);
  spice_transistor_nmos t1779(~dpc1_SBY_v[`W-1], y5_v, sb5_v, y5_i0, sb5_i5);
  spice_transistor_nmos t1576(~cclk_v[`W-1], y3_v, n1531_v, y3_i0, n1531_i1);
  spice_transistor_nmos_gnd t1573(~n15_v[`W-1], pclp4_v, pclp4_i0);
  spice_transistor_nmos_gnd t1570(~alucin_v[`W-1], notalucin_v, notalucin_i1);
  spice_transistor_nmos t1571(~cclk_v[`W-1], n658_v, y4_v, n658_i0, y4_i2);
  spice_transistor_nmos t1578(~cp1_v[`W-1], n472_v, n1606_v, n472_i0, n1606_i0);
  spice_transistor_nmos t1579(~cclk_v[`W-1], pipeUNK05_v, n90_v, pipeUNK05_i0, n90_i0);
  spice_transistor_nmos_gnd t2642(~n625_v[`W-1], n662_v, n662_i0);
  spice_transistor_nmos_gnd t1685(~n476_v[`W-1], n956_v, n956_i0);
  spice_transistor_nmos_vdd t1686(~n476_v[`W-1], dpc12_0ADD_v, dpc12_0ADD_i7);
  spice_transistor_nmos_gnd t1681(~s4_v[`W-1], n973_v, n973_i1);
  spice_transistor_nmos_gnd t1682(~n1471_v[`W-1], Pout4_v, Pout4_i0);
  spice_transistor_nmos t1683(~cclk_v[`W-1], n1586_v, n621_v, n1586_i0, n621_i1);
  spice_transistor_nmos_gnd t1689(~idb5_v[`W-1], n961_v, n961_i0);
  spice_transistor_nmos t993(~dpc37_PCLDB_v[`W-1], idb2_v, n481_v, idb2_i3, n481_i1);
  spice_transistor_nmos_gnd t1307(~adh2_v[`W-1], n168_v, n168_i0);
  spice_transistor_nmos_gnd t2033(~pd2_clearIR_v[`W-1], n571_v, n571_i0);
  spice_transistor_nmos_gnd t991(~abh5_v[`W-1], n1423_v, n1423_i0);
  spice_transistor_nmos_vdd t3132(~n531_v[`W-1], dpc13_ORS_v, dpc13_ORS_i8);
  spice_transistor_nmos t585(~dpc43_DL_DB_v[`W-1], idb0_v, n719_v, idb0_i5, n719_i2);
  spice_transistor_nmos_vdd t3133(~dor7_v[`W-1], n298_v, n298_i1);
  spice_transistor_nmos t587(~dpc43_DL_DB_v[`W-1], idb2_v, n1424_v, idb2_i1, n1424_i2);
  spice_transistor_nmos_gnd t2037(~notidl4_v[`W-1], idl4_v, idl4_i0);
  spice_transistor_nmos_gnd g_1212((~n1247_v[`W-1]|~n225_v[`W-1]|~cclk_v[`W-1]), dpc9_DBADD_v, dpc9_DBADD_i9);
  spice_transistor_nmos t586(~dpc43_DL_DB_v[`W-1], idb1_v, n87_v, idb1_i0, n87_i2);
  spice_transistor_nmos t581(~cp1_v[`W-1], notRdy0_v, n1679_v, notRdy0_i3, n1679_i0);
  spice_transistor_nmos_gnd t852(~ir7_v[`W-1], _op_branch_bit7_v, _op_branch_bit7_i0);
  spice_transistor_nmos_gnd t2590(~_ABL4_v[`W-1], abl4_v, abl4_i0);
  spice_transistor_nmos t1985(~dpc1_SBY_v[`W-1], y3_v, sb3_v, y3_i2, sb3_i8);
  spice_transistor_nmos t582(~cp1_v[`W-1], n223_v, n1215_v, n223_i1, n1215_i0);
  spice_transistor_nmos t259(~cclk_v[`W-1], n242_v, x3_v, n242_i0, x3_i0);
  spice_transistor_nmos t251(~dpc6_SBS_v[`W-1], dasb4_v, s4_v, dasb4_i4, s4_i0);
  spice_transistor_nmos t250(~dpc6_SBS_v[`W-1], s3_v, sb3_v, s3_i0, sb3_i2);
  spice_transistor_nmos t253(~dpc6_SBS_v[`W-1], s2_v, sb2_v, s2_i0, sb2_i2);
  spice_transistor_nmos t252(~dpc6_SBS_v[`W-1], s1_v, sb1_v, s1_i0, sb1_i1);
  spice_transistor_nmos t1984(~dpc40_ADLPCL_v[`W-1], pcl7_v, adl7_v, pcl7_i1, adl7_i4);
  spice_transistor_nmos_gnd g_1077((~irline3_v[`W-1]|~ir6_v[`W-1]|~notir2_v[`W-1]|~notir5_v[`W-1]|~clock1_v[`W-1]|~ir7_v[`W-1]|~ir4_v[`W-1]), x_op_T0_bit_v, x_op_T0_bit_i2);
  spice_transistor_nmos_gnd g_1262((~cclk_v[`W-1]|~n956_v[`W-1]|~n1247_v[`W-1]), dpc12_0ADD_v, dpc12_0ADD_i9);
  spice_transistor_nmos t2133(~cp1_v[`W-1], n961_v, notdor5_v, n961_i1, notdor5_i0);
  spice_transistor_nmos t3211(~cclk_v[`W-1], n19_v, pipeUNK18_v, n19_i0, pipeUNK18_i1);
  spice_transistor_nmos t3210(~dpc10_ADLADD_v[`W-1], adl3_v, alub3_v, adl3_i6, alub3_i2);
  spice_transistor_nmos_gnd t3214(~db0_v[`W-1], n718_v, n718_i1);
  spice_transistor_nmos_gnd t3217(~db2_v[`W-1], n111_v, n111_i1);
  spice_transistor_nmos_gnd t2648(~_C12_v[`W-1], C12_v, C12_i0);
  spice_transistor_nmos_gnd t3219(~db3_v[`W-1], n896_v, n896_i1);
  spice_transistor_nmos t3218(~cclk_v[`W-1], n304_v, notalu7_v, n304_i5, notalu7_i1);
  spice_transistor_nmos_gnd g_1346((~n753_v[`W-1]|~n1135_v[`W-1]), n1629_v, n1629_i1);
  spice_transistor_nmos_vdd t382(~n1076_v[`W-1], db4_v, db4_i0);
  spice_transistor_nmos_gnd t386(~op_ror_v[`W-1], n544_v, n544_i0);
  spice_transistor_nmos t385(~dpc4_SSB_v[`W-1], n280_v, sb5_v, n280_i1, sb5_i2);
  spice_transistor_nmos_gnd t384(~pcl7_v[`W-1], n641_v, n641_i0);
  spice_transistor_nmos_gnd t3036(~pcl4_v[`W-1], n1643_v, n1643_i0);
  spice_transistor_nmos_gnd g_1124((~ir4_v[`W-1]|~notir0_v[`W-1]|~ir2_v[`W-1]|~ir3_v[`W-1]|~t3_v[`W-1]), op_T3_ind_x_v, op_T3_ind_x_i1);
  spice_transistor_nmos t1988(~cp1_v[`W-1], n913_v, n1274_v, n913_i1, n1274_i0);
  spice_transistor_nmos_gnd g_1121((~ir7_v[`W-1]|~ir4_v[`W-1]|~ir2_v[`W-1]|~notir6_v[`W-1]|~ir5_v[`W-1]|~ir3_v[`W-1]|~t5_v[`W-1]|~irline3_v[`W-1]), op_T5_rti_v, op_T5_rti_i2);
  spice_transistor_nmos t3328(~cclk_v[`W-1], pipephi2Reset0_v, Reset0_v, pipephi2Reset0_i0, Reset0_i1);
  spice_transistor_nmos_vdd t3458(~n634_v[`W-1], ab4_v, ab4_i1);
  spice_transistor_nmos_gnd t3457(~n1358_v[`W-1], n396_v, n396_i1);
  spice_transistor_nmos_gnd t2056(~n676_v[`W-1], ab9_v, ab9_i1);
  spice_transistor_nmos_gnd t3321(~notalu3_v[`W-1], alu3_v, alu3_i2);
  spice_transistor_nmos_vdd t3323(~n1277_v[`W-1], dpc42_DL_ADH_v, dpc42_DL_ADH_i9);
  spice_transistor_nmos_gnd t3322(~n1277_v[`W-1], n1441_v, n1441_i1);
  spice_transistor_nmos_gnd g_1066((~notir2_v[`W-1]|~irline3_v[`W-1]|~ir4_v[`W-1]|~clock2_v[`W-1]|~notir7_v[`W-1]|~notir3_v[`W-1]|~notir6_v[`W-1]), op_T__cpx_cpy_abs_v, op_T__cpx_cpy_abs_i1);
  spice_transistor_nmos_gnd g_1071((~cclk_v[`W-1]|~n1247_v[`W-1]|~n228_v[`W-1]), dpc30_ADHPCH_v, dpc30_ADHPCH_i9);
  spice_transistor_nmos_gnd g_1298((~n1449_v[`W-1]|~n759_v[`W-1]), n944_v, n944_i2);
  spice_transistor_nmos_gnd g_1299((~n43_v[`W-1]|~n1027_v[`W-1]), n476_v, n476_i3);
  spice_transistor_nmos_gnd g_1292((~n43_v[`W-1]|~n1162_v[`W-1]), n21_v, n21_i3);
  spice_transistor_nmos_gnd g_1293((~notir6_v[`W-1]|~ir2_v[`W-1]|~ir4_v[`W-1]|~clock2_v[`W-1]|~notir3_v[`W-1]|~notir7_v[`W-1]|~ir5_v[`W-1]|~notir1_v[`W-1]), op_T__dex_v, op_T__dex_i1);
  spice_transistor_nmos_gnd g_1290((~notir7_v[`W-1]|~notir4_v[`W-1]|~ir6_v[`W-1]|~ir2_v[`W-1]|~notir3_v[`W-1]|~notir1_v[`W-1]|~clock1_v[`W-1]|~ir5_v[`W-1]), op_T0_txs_v, op_T0_txs_i2);
  spice_transistor_nmos_gnd g_1291((~ir6_v[`W-1]|~ir2_v[`W-1]|~notir4_v[`W-1]|~notir3_v[`W-1]|~notir5_v[`W-1]|~notir1_v[`W-1]|~notir7_v[`W-1]|~clock1_v[`W-1]), op_T0_tsx_v, op_T0_tsx_i2);
  spice_transistor_nmos_gnd g_1296((~notir2_v[`W-1]|~notir4_v[`W-1]|~ir3_v[`W-1]|~t3_v[`W-1]), op_T3_mem_zp_idx_v, op_T3_mem_zp_idx_i2);
  spice_transistor_nmos_gnd g_1297((~n192_v[`W-1]|~n256_v[`W-1]), n25_v, n25_i2);
  spice_transistor_nmos_gnd g_1295((~n771_v[`W-1]|~n850_v[`W-1]), n1446_v, n1446_i2);
  spice_transistor_nmos t2032(~cclk_v[`W-1], n80_v, n1333_v, n80_i0, n1333_i1);
  spice_transistor_nmos t1961(~dpc5_SADL_v[`W-1], adl0_v, n332_v, adl0_i4, n332_i1);
  spice_transistor_nmos_gnd t1960(~pcl6_v[`W-1], n232_v, n232_i0);
  spice_transistor_nmos_gnd t3038(~n147_v[`W-1], db4_v, db4_i3);
  spice_transistor_nmos_gnd g_1348((~op_branch_done_v[`W-1]|~n1211_v[`W-1]|~n467_v[`W-1]), n10_v, n10_i2);
  spice_transistor_nmos_gnd g_1349((~n930_v[`W-1]|~n470_v[`W-1]), n1286_v, n1286_i1);
  spice_transistor_nmos_vdd t3035(~n769_v[`W-1], n1072_v, n1072_i0);
  spice_transistor_nmos_gnd g_1341((~n1662_v[`W-1]|~n781_v[`W-1]), n553_v, n553_i1);
  spice_transistor_nmos_gnd g_1342((~op_ANDS_v[`W-1]|~n384_v[`W-1]), n550_v, n550_i2);
  spice_transistor_nmos t1964(~cclk_v[`W-1], n1300_v, notir2_v, n1300_i1, notir2_i1);
  spice_transistor_nmos_gnd g_1125((~notir4_v[`W-1]|~ir2_v[`W-1]|~t4_v[`W-1]|~ir3_v[`W-1]|~notir0_v[`W-1]), op_T4_ind_y_v, op_T4_ind_y_i1);
  spice_transistor_nmos_gnd g_1126((~t3_v[`W-1]|~ir2_v[`W-1]|~ir3_v[`W-1]|~notir0_v[`W-1]|~notir4_v[`W-1]), x_op_T3_ind_y_v, x_op_T3_ind_y_i2);
  spice_transistor_nmos_gnd g_1127((~pd4_clearIR_v[`W-1]|~pd0_clearIR_v[`W-1]|~pd3_clearIR_v[`W-1]|~pd2_clearIR_v[`W-1]|~n1605_v[`W-1]), PD_1xx000x0_v, PD_1xx000x0_i1);
  spice_transistor_nmos_gnd g_1120((~notir6_v[`W-1]|~ir2_v[`W-1]|~ir4_v[`W-1]|~ir3_v[`W-1]|~ir5_v[`W-1]|~t4_v[`W-1]|~irline3_v[`W-1]|~ir7_v[`W-1]), op_T4_rti_v, op_T4_rti_i1);
  spice_transistor_nmos_gnd t1967(~n1691_v[`W-1], n110_v, n110_i0);
  spice_transistor_nmos_gnd g_1122((~t2_v[`W-1]|~ir3_v[`W-1]), op_T2_ADL_ADD_v, op_T2_ADL_ADD_i1);
  spice_transistor_nmos_gnd g_1123((~t2_v[`W-1]|~notir0_v[`W-1]|~ir3_v[`W-1]|~ir2_v[`W-1]|~notir4_v[`W-1]), op_T2_ind_y_v, op_T2_ind_y_i1);
  spice_transistor_nmos_gnd g_1128((~pd4_clearIR_v[`W-1]|~pd1_clearIR_v[`W-1]|~pd7_clearIR_v[`W-1]), PD_0xx0xx0x_v, PD_0xx0xx0x_i2);
  spice_transistor_nmos_gnd g_1129((~irline3_v[`W-1]|~ir6_v[`W-1]|~ir2_v[`W-1]|~notir3_v[`W-1]|~ir7_v[`W-1]|~clock1_v[`W-1]|~notir5_v[`W-1]|~ir4_v[`W-1]), op_T0_plp_v, op_T0_plp_i1);
  spice_transistor_nmos_gnd g_1089((~ir1_v[`W-1]|~ir0_v[`W-1]), n1133_v, n1133_i2);
  spice_transistor_nmos_gnd g_1514((~Pout3_v[`W-1]&~op_T0_adc_sbc_v[`W-1]), n673_v, n673_i2);
  spice_transistor_nmos_gnd g_1045((~clock1_v[`W-1]|~ir5_v[`W-1]|~ir7_v[`W-1]|~ir6_v[`W-1]|~notir0_v[`W-1]), op_T0_ora_v, op_T0_ora_i1);
  spice_transistor_nmos_gnd g_1044((~ir4_v[`W-1]|~notir3_v[`W-1]|~ir2_v[`W-1]|~ir5_v[`W-1]|~ir7_v[`W-1]|~irline3_v[`W-1]|~clock1_v[`W-1]), op_T0_php_pha_v, op_T0_php_pha_i1);
  spice_transistor_nmos_gnd g_1043((~clock1_v[`W-1]|~ir5_v[`W-1]|~ir7_v[`W-1]|~notir6_v[`W-1]|~notir0_v[`W-1]), op_T0_eor_v, op_T0_eor_i2);
  spice_transistor_nmos_gnd g_1042((~ir3_v[`W-1]|~ir2_v[`W-1]|~notir0_v[`W-1]|~ir4_v[`W-1]|~t2_v[`W-1]), op_T2_ind_x_v, op_T2_ind_x_i1);
  spice_transistor_nmos_gnd t3147(~abl4_v[`W-1], n86_v, n86_i3);
  spice_transistor_nmos_gnd t3146(~n469_v[`W-1], pchp5_v, pchp5_i1);
  spice_transistor_nmos_gnd t2328(~n1133_v[`W-1], irline3_v, irline3_i0);
  spice_transistor_nmos_vdd t2326(~n1566_v[`W-1], dpc43_DL_DB_v, dpc43_DL_DB_i9);
  spice_transistor_nmos t2324(~cclk_v[`W-1], n1455_v, n1505_v, n1455_i1, n1505_i0);
  spice_transistor_nmos_gnd t2325(~n1566_v[`W-1], n1240_v, n1240_i1);
  spice_transistor_nmos t2320(~dpc37_PCLDB_v[`W-1], n72_v, idb5_v, n72_i1, idb5_i6);
  spice_transistor_nmos_gnd t2321(~aluanorb0_v[`W-1], aluaorb0_v, aluaorb0_i0);
  spice_transistor_nmos_gnd t1369(~notidl0_v[`W-1], idl0_v, idl0_i1);
  spice_transistor_nmos_gnd t1365(~idb4_v[`W-1], n478_v, n478_i1);
  spice_transistor_nmos_gnd g_1630(((~pipeUNK04_v[`W-1]&~n1457_v[`W-1])|(~n1600_v[`W-1]&~n781_v[`W-1])|(~n270_v[`W-1]&~n1492_v[`W-1])), n1495_v, n1495_i2);
  spice_transistor_nmos_gnd g_1631(((~n609_v[`W-1]&~n453_v[`W-1])|~n1213_v[`W-1]), n1209_v, n1209_i2);
  spice_transistor_nmos_gnd g_1632(((~n1416_v[`W-1]&~n1111_v[`W-1])|~n587_v[`W-1]|(~n1614_v[`W-1]&~pipeUNK05_v[`W-1])|(~n1245_v[`W-1]&~pipeUNK03_v[`W-1])), n299_v, n299_i2);
  spice_transistor_nmos_gnd g_1633((~n1159_v[`W-1]|(~n1580_v[`W-1]&~n613_v[`W-1])), dasb2_v, dasb2_i2);
  spice_transistor_nmos_gnd g_1634(((~n233_v[`W-1]&~n1257_v[`W-1])|(~n1018_v[`W-1]&~n811_v[`W-1])), n1205_v, n1205_i2);
  spice_transistor_nmos_gnd g_1635(((~n761_v[`W-1]&~n1257_v[`W-1])|(~n1056_v[`W-1]&~n811_v[`W-1])), n739_v, n739_i2);
  spice_transistor_nmos_gnd g_1636((~n297_v[`W-1]|(~n284_v[`W-1]&~cclk_v[`W-1])), NMIP_v, NMIP_i3);
  spice_transistor_nmos_gnd g_1637((~n1126_v[`W-1]|(~VEC1_v[`W-1]&~notRdy0_v[`W-1])), n1290_v, n1290_i2);
  spice_transistor_nmos_gnd g_1638(((~x_op_T__adc_sbc_v[`W-1]|~op_T__cpx_cpy_abs_v[`W-1]|~op_T__asl_rol_a_v[`W-1]|~op_T__cmp_v[`W-1]|~op_T__cpx_cpy_imm_zp_v[`W-1])|(~op_asl_rol_v[`W-1]&~n1258_v[`W-1])), _op_set_C_v, _op_set_C_i2);
  spice_transistor_nmos_gnd g_1639(((~n739_v[`W-1]&~n61_v[`W-1])|~n479_v[`W-1]), dasb6_v, dasb6_i2);
  spice_transistor_nmos t538(~dpc13_ORS_v[`W-1], n740_v, n1691_v, n740_i0, n1691_i0);
  spice_transistor_nmos_gnd t534(~n990_v[`W-1], n1041_v, n1041_i1);
  spice_transistor_nmos_vdd t535(~n990_v[`W-1], n138_v, n138_i1);
  spice_transistor_nmos_vdd t2148(~cclk_v[`W-1], adh5_v, adh5_i2);
  spice_transistor_nmos_vdd t2149(~cclk_v[`W-1], adl6_v, adl6_i3);
  spice_transistor_nmos_gnd t2920(~n1674_v[`W-1], n772_v, n772_i2);
  spice_transistor_nmos_gnd t1217(~adl0_v[`W-1], n123_v, n123_i0);
  spice_transistor_nmos_gnd t1216(~n1272_v[`W-1], n608_v, n608_i0);
  spice_transistor_nmos t1214(~cclk_v[`W-1], pchp4_v, n1657_v, pchp4_i1, n1657_i0);
  spice_transistor_nmos t1211(~dpc20_ADDSB06_v[`W-1], alu3_v, sb3_v, alu3_i1, sb3_i4);
  spice_transistor_nmos t1210(~dpc20_ADDSB06_v[`W-1], dasb4_v, alu4_v, dasb4_i5, alu4_i2);
  spice_transistor_nmos t3374(~dpc40_ADLPCL_v[`W-1], adl0_v, pcl0_v, adl0_i8, pcl0_i2);
  spice_transistor_nmos t3375(~dpc40_ADLPCL_v[`W-1], pcl3_v, adl3_v, pcl3_i2, adl3_i7);
  spice_transistor_nmos_vdd t2778(~n842_v[`W-1], n66_v, n66_i3);
  spice_transistor_nmos_gnd g_1191((~ir7_v[`W-1]|~ir6_v[`W-1]|~notir5_v[`W-1]|~notir1_v[`W-1]), op_rol_ror_v, op_rol_ror_i1);
  spice_transistor_nmos_gnd g_1190((~notir6_v[`W-1]|~ir4_v[`W-1]|~t4_v[`W-1]|~ir2_v[`W-1]|~notir5_v[`W-1]|~irline3_v[`W-1]|~ir7_v[`W-1]|~ir3_v[`W-1]), op_T4_rts_v, op_T4_rts_i1);
  spice_transistor_nmos t2595(~dpc13_ORS_v[`W-1], n1632_v, n277_v, n1632_i1, n277_i5);
  spice_transistor_nmos_gnd t1785(~db4_v[`W-1], n490_v, n490_i1);
  spice_transistor_nmos_gnd t1780(~pipeUNK15_v[`W-1], H1x1_v, H1x1_i4);
  spice_transistor_nmos t1782(~dpc1_SBY_v[`W-1], y7_v, sb7_v, y7_i1, sb7_i4);
  spice_transistor_nmos_gnd t1543(~n1084_v[`W-1], n803_v, n803_i0);
  spice_transistor_nmos_gnd t1540(~idb4_v[`W-1], n797_v, n797_i1);
  spice_transistor_nmos t1547(~cclk_v[`W-1], op_EORS_v, n982_v, op_EORS_i0, n982_i1);
  spice_transistor_nmos t1549(~cclk_v[`W-1], op_ORS_v, n88_v, op_ORS_i0, n88_i1);
  spice_transistor_nmos_vdd t1548(~cclk_v[`W-1], sb7_v, sb7_i3);
  spice_transistor_nmos_gnd t2490(~dpc29_0ADH17_v[`W-1], adh7_v, adh7_i4);
  spice_transistor_nmos_gnd t2491(~dpc29_0ADH17_v[`W-1], adh6_v, adh6_i4);
  spice_transistor_nmos_gnd g_1096((~n523_v[`W-1]|~n499_v[`W-1]), n743_v, n743_i1);
  spice_transistor_nmos_vdd t2818(~dor6_v[`W-1], n7_v, n7_i0);
  spice_transistor_nmos_gnd g_1620((~n404_v[`W-1]|(~_C34_v[`W-1]&~n1063_v[`W-1])), C45_v, C45_i2);
  spice_transistor_nmos_gnd t2819(~n_0_ADL0_v[`W-1], adl0_v, adl0_i7);
  spice_transistor_nmos_gnd g_1438((~fetch_v[`W-1]&~D1x1_v[`W-1]), clearIR_v, clearIR_i9);
  spice_transistor_nmos_gnd g_1093((~n506_v[`W-1]|~n933_v[`W-1]), n877_v, n877_i1);
  spice_transistor_nmos t49(~dpc11_SBADD_v[`W-1], alua4_v, dasb4_v, alua4_i0, dasb4_i1);
  spice_transistor_nmos t48(~dpc11_SBADD_v[`W-1], alua3_v, sb3_v, alua3_i0, sb3_i0);
  spice_transistor_nmos_gnd t42(~pd0_clearIR_v[`W-1], n409_v, n409_i0);
  spice_transistor_nmos t47(~dpc11_SBADD_v[`W-1], sb2_v, alua2_v, sb2_i0, alua2_i0);
  spice_transistor_nmos t46(~dpc11_SBADD_v[`W-1], sb1_v, alua1_v, sb1_i0, alua1_i0);
  spice_transistor_nmos t45(~cclk_v[`W-1], y1_v, n767_v, y1_i0, n767_i0);
  spice_transistor_nmos_gnd t44(~notalu4_v[`W-1], alu4_v, alu4_i0);
  spice_transistor_nmos t3203(~dpc10_ADLADD_v[`W-1], adl6_v, alub6_v, adl6_i6, alub6_i2);
  spice_transistor_nmos t3200(~cclk_v[`W-1], n680_v, n1688_v, n680_i0, n1688_i1);
  spice_transistor_nmos t3206(~dpc10_ADLADD_v[`W-1], adl1_v, alub1_v, adl1_i7, alub1_i2);
  spice_transistor_nmos t3207(~dpc10_ADLADD_v[`W-1], adl4_v, alub4_v, adl4_i6, alub4_i2);
  spice_transistor_nmos t3204(~dpc10_ADLADD_v[`W-1], adl7_v, alub7_v, adl7_i6, alub7_i2);
  spice_transistor_nmos t3208(~dpc10_ADLADD_v[`W-1], alub5_v, adl5_v, alub5_i2, adl5_i5);
  spice_transistor_nmos t3209(~cclk_v[`W-1], n1126_v, VEC0_v, n1126_i0, VEC0_i1);
  spice_transistor_nmos_gnd g_1248((~notir3_v[`W-1]|~notir4_v[`W-1]|~t4_v[`W-1]), op_T4_abs_idx_v, op_T4_abs_idx_i1);
  spice_transistor_nmos_gnd g_1242((~cclk_v[`W-1]|~n1247_v[`W-1]|~n1518_v[`W-1]), dpc39_PCLPCL_v, dpc39_PCLPCL_i9);
  spice_transistor_nmos t283(~dpc7_SS_v[`W-1], n618_v, s6_v, n618_i1, s6_i1);
  spice_transistor_nmos_gnd t280(~n101_v[`W-1], n1364_v, n1364_i0);
  spice_transistor_nmos t286(~dpc7_SS_v[`W-1], n998_v, s3_v, n998_i1, s3_i1);
  spice_transistor_nmos t287(~dpc7_SS_v[`W-1], n1389_v, s2_v, n1389_i1, s2_i1);
  spice_transistor_nmos t284(~dpc7_SS_v[`W-1], n280_v, s5_v, n280_i0, s5_i1);
  spice_transistor_nmos t285(~dpc7_SS_v[`W-1], n3_v, s4_v, n3_i1, s4_i1);
  spice_transistor_nmos_gnd t3336(~db7_v[`W-1], n62_v, n62_i1);
  spice_transistor_nmos t3337(~cp1_v[`W-1], n1338_v, n720_v, n1338_i0, n720_i0);
  spice_transistor_nmos t288(~dpc7_SS_v[`W-1], n694_v, s1_v, n694_i0, s1_i1);
  spice_transistor_nmos_gnd t289(~adh3_v[`W-1], n883_v, n883_i0);
  spice_transistor_nmos_gnd t3332(~pd1_clearIR_v[`W-1], n1641_v, n1641_i0);
  spice_transistor_nmos_vdd t3331(~cclk_v[`W-1], idb1_v, idb1_i9);
  spice_transistor_nmos g_1522((~cp1_v[`W-1]&~fetch_v[`W-1]), n928_v, n1609_v, n928_i2, n1609_i2);
  spice_transistor_nmos_gnd g_1289((~n1642_v[`W-1]|~n335_v[`W-1]|~n1258_v[`W-1]|~n440_v[`W-1]|~op_T4_brk_v[`W-1]|~op_T2_php_pha_v[`W-1]), _WR_v, _WR_i2);
  spice_transistor_nmos t2519(~cclk_v[`W-1], pipeT5out_v, n378_v, pipeT5out_i0, n378_i1);
  spice_transistor_nmos t2799(~dpc8_nDBADD_v[`W-1], alub6_v, n351_v, alub6_i1, n351_i1);
  spice_transistor_nmos_gnd t2797(~n565_v[`W-1], n658_v, n658_i2);
  spice_transistor_nmos_gnd g_1280((~ir7_v[`W-1]|~ir4_v[`W-1]|~notir3_v[`W-1]|~ir2_v[`W-1]|~notir5_v[`W-1]|~irline3_v[`W-1]), op_plp_pla_v, op_plp_pla_i1);
  spice_transistor_nmos_gnd g_1282((~notir6_v[`W-1]|~notir3_v[`W-1]|~ir2_v[`W-1]|~ir7_v[`W-1]|~ir4_v[`W-1]|~clock1_v[`W-1]|~irline3_v[`W-1]|~notir5_v[`W-1]), op_T0_pla_v, op_T0_pla_i2);
  spice_transistor_nmos_gnd g_1284((~clearIR_v[`W-1]|~pd4_v[`W-1]), pd4_clearIR_v, pd4_clearIR_i5);
  spice_transistor_nmos t2009(~cclk_v[`W-1], n541_v, notir7_v, n541_i0, notir7_i1);
  spice_transistor_nmos_gnd t2008(~n1067_v[`W-1], ADH_ABH_v, ADH_ABH_i1);
  spice_transistor_nmos_gnd g_1358((~n1024_v[`W-1]|~n1274_v[`W-1]), n1069_v, n1069_i2);
  spice_transistor_nmos_gnd t3022(~n393_v[`W-1], n551_v, n551_i1);
  spice_transistor_nmos t3023(~cclk_v[`W-1], pipeUNK23_v, n1085_v, pipeUNK23_i0, n1085_i0);
  spice_transistor_nmos_gnd t3021(~adl1_v[`W-1], n1016_v, n1016_i0);
  spice_transistor_nmos t3024(~cclk_v[`W-1], n1175_v, pipeUNK28_v, n1175_i1, pipeUNK28_i0);
  spice_transistor_nmos_gnd g_1133((~notir2_v[`W-1]|~ir6_v[`W-1]|~notir7_v[`W-1]|~clock1_v[`W-1]|~notir5_v[`W-1]|~irline3_v[`W-1]), op_T0_ldy_mem_v, op_T0_ldy_mem_i1);
  spice_transistor_nmos_gnd g_1132((~ir4_v[`W-1]|~irline3_v[`W-1]|~ir6_v[`W-1]|~notir5_v[`W-1]|~notir7_v[`W-1]|~clock1_v[`W-1]), op_T0_tay_ldy_not_idx_v, op_T0_tay_ldy_not_idx_i1);
  spice_transistor_nmos_gnd g_1131((~notir6_v[`W-1]|~ir4_v[`W-1]|~ir2_v[`W-1]|~notir3_v[`W-1]|~notir7_v[`W-1]|~irline3_v[`W-1]|~notir5_v[`W-1]|~clock2_v[`W-1]), op_T__inx_v, op_T__inx_i1);
  spice_transistor_nmos_gnd g_1137((~notir3_v[`W-1]|~irline3_v[`W-1]|~ir6_v[`W-1]|~clock1_v[`W-1]|~notir4_v[`W-1]|~ir7_v[`W-1]|~ir2_v[`W-1]), op_T0_clc_sec_v, op_T0_clc_sec_i2);
  spice_transistor_nmos_gnd t2889(~ir4_v[`W-1], notir4_v, notir4_i1);
  spice_transistor_nmos_gnd g_1135((~n43_v[`W-1]|~n1505_v[`W-1]), n830_v, n830_i3);
  spice_transistor_nmos_gnd t3470(~n329_v[`W-1], n1166_v, n1166_i0);
  spice_transistor_nmos t637(~cclk_v[`W-1], y2_v, n1491_v, y2_i0, n1491_i0);
  spice_transistor_nmos_gnd t2140(~notdor0_v[`W-1], dor0_v, dor0_i0);
  spice_transistor_nmos_gnd t2141(~aluvout_v[`W-1], n1245_v, n1245_i0);
  spice_transistor_nmos_gnd g_1214((~op_T2_stack_access_v[`W-1]|~n1222_v[`W-1]), n1090_v, n1090_i2);
  spice_transistor_nmos t2146(~cclk_v[`W-1], n1169_v, x0_v, n1169_i2, x0_i1);
  spice_transistor_nmos t2239(~dpc26_ACDB_v[`W-1], idb4_v, n1344_v, idb4_i5, n1344_i0);
  spice_transistor_nmos_gnd t1963(~s2_v[`W-1], n1190_v, n1190_i0);
  spice_transistor_nmos t2147(~cclk_v[`W-1], n588_v, notidl7_v, n588_i1, notidl7_i1);
  spice_transistor_nmos_gnd t3156(~PD_xxxx10x0_v[`W-1], n231_v, n231_i1);
  spice_transistor_nmos_gnd t3157(~pclp6_v[`W-1], n1458_v, n1458_i2);
  spice_transistor_nmos_gnd t3152(~n681_v[`W-1], DA_AB2_v, DA_AB2_i0);
  spice_transistor_nmos_gnd t3150(~n1434_v[`W-1], n1709_v, n1709_i1);
  spice_transistor_nmos_gnd t3151(~nots2_v[`W-1], n1389_v, n1389_i3);
  spice_transistor_nmos_gnd t2145(~n850_v[`W-1], n430_v, n430_i2);
  spice_transistor_nmos_gnd g_1629((~n854_v[`W-1]|(~n995_v[`W-1]&~cclk_v[`W-1])), n975_v, n975_i1);
  spice_transistor_nmos_gnd g_1628(((~n783_v[`W-1]&~n1542_v[`W-1])|~n1253_v[`W-1]), n515_v, n515_i2);
  spice_transistor_nmos_gnd g_1627(((~n335_v[`W-1]&~op_sta_cmp_v[`W-1])|~op_T2_pha_v[`W-1]), n1037_v, n1037_i2);
  spice_transistor_nmos_gnd g_1626(((~n206_v[`W-1]&~n853_v[`W-1])|~n1517_v[`W-1]), n916_v, n916_i3);
  spice_transistor_nmos_gnd g_1625((~n410_v[`W-1]|(~n1184_v[`W-1]&~n1643_v[`W-1])), n474_v, n474_i2);
  spice_transistor_nmos_gnd g_1624(((~C34_v[`W-1]&~__AxB_4_v[`W-1])|~_AxB_4__C34_v[`W-1]), __AxBxC_4_v, __AxBxC_4_i2);
  spice_transistor_nmos_gnd g_1623(((~cclk_v[`W-1]&~n538_v[`W-1])|~n807_v[`W-1]), n330_v, n330_i3);
  spice_transistor_nmos_gnd g_1622(((~A_B7_v[`W-1]&~C67_v[`W-1])|~n748_v[`W-1]), _C78_v, _C78_i2);
  spice_transistor_nmos_gnd g_1621(((~n253_v[`W-1]&~n270_v[`W-1])|(~n279_v[`W-1]&~pipeUNK16_v[`W-1])|(~n1224_v[`W-1]&~n507_v[`W-1])|(~n954_v[`W-1]&~n206_v[`W-1])), n1082_v, n1082_i2);
  spice_transistor_nmos_gnd t2173(~t4_v[`W-1], op_T4_v, op_T4_i0);
  spice_transistor_nmos t528(~dpc21_ADDADL_v[`W-1], adl6_v, alu6_v, adl6_i1, alu6_i1);
  spice_transistor_nmos t1208(~dpc20_ADDSB06_v[`W-1], alu6_v, sb6_v, alu6_i2, sb6_i6);
  spice_transistor_nmos t1209(~dpc20_ADDSB06_v[`W-1], alu5_v, sb5_v, alu5_i1, sb5_i3);
  spice_transistor_nmos_gnd t2777(~n842_v[`W-1], n1479_v, n1479_i1);
  spice_transistor_nmos t2771(~cclk_v[`W-1], pipeUNK40_v, n191_v, pipeUNK40_i0, n191_i0);
  spice_transistor_nmos_gnd t2773(~n404_v[`W-1], n918_v, n918_i0);
  spice_transistor_nmos_gnd t1201(~n1221_v[`W-1], n1566_v, n1566_i0);
  spice_transistor_nmos t1203(~cclk_v[`W-1], _WR_v, pipe_WR_phi2_v, _WR_i0, pipe_WR_phi2_i0);
  spice_transistor_nmos t1205(~cp1_v[`W-1], n1375_v, n95_v, n1375_i1, n95_i0);
  spice_transistor_nmos t1206(~cp1_v[`W-1], n1089_v, n1529_v, n1089_i0, n1529_i1);
  spice_transistor_nmos_gnd t1375(~p1_v[`W-1], n318_v, n318_i1);
  spice_transistor_nmos_gnd t1372(~n1683_v[`W-1], n966_v, n966_i0);
  spice_transistor_nmos_gnd t1379(~pchp5_v[`W-1], n1301_v, n1301_i0);
  spice_transistor_nmos t2863(~cclk_v[`W-1], n633_v, n1059_v, n633_i0, n1059_i0);
  spice_transistor_nmos_gnd t1799(~n1565_v[`W-1], n1218_v, n1218_i0);
  spice_transistor_nmos t1796(~cclk_v[`W-1], n1049_v, n160_v, n1049_i0, n160_i0);
  spice_transistor_nmos_gnd t1797(~n477_v[`W-1], n647_v, n647_i0);
  spice_transistor_nmos_gnd t1792(~n1501_v[`W-1], db7_v, db7_i1);
  spice_transistor_nmos t1790(~cclk_v[`W-1], pipeUNK27_v, op_SRS_v, pipeUNK27_i1, op_SRS_i0);
  spice_transistor_nmos t1558(~cp1_v[`W-1], n1624_v, notRdy0_v, n1624_i0, notRdy0_i6);
  spice_transistor_nmos_gnd t1554(~n86_v[`W-1], ab4_v, ab4_i0);
  spice_transistor_nmos_gnd t1552(~sb2_v[`W-1], n1580_v, n1580_i0);
  spice_transistor_nmos_gnd t1969(~pclp3_v[`W-1], n723_v, n723_i0);
  spice_transistor_nmos_vdd t3442(~n7_v[`W-1], db6_v, db6_i3);
  spice_transistor_nmos_gnd g_1025((~notir3_v[`W-1]|~ir7_v[`W-1]|~ir4_v[`W-1]|~irline3_v[`W-1]|~t2_v[`W-1]|~ir5_v[`W-1]|~ir2_v[`W-1]), op_T2_php_pha_v, op_T2_php_pha_i1);
  spice_transistor_nmos_gnd g_1408((~n1693_v[`W-1]|~n1291_v[`W-1]), n1312_v, n1312_i2);
  spice_transistor_nmos_gnd g_1028((~ir2_v[`W-1]|~ir4_v[`W-1]|~notir3_v[`W-1]|~notir5_v[`W-1]|~irline3_v[`W-1]|~ir7_v[`W-1]|~t3_v[`W-1]), x_op_T3_plp_pla_v, x_op_T3_plp_pla_i1);
  spice_transistor_nmos_gnd g_1368((~op_T4_ind_x_v[`W-1]|~op_T2_abs_v[`W-1]|~op_jmp_v[`W-1]|~notRdy0_v[`W-1]|~n1109_v[`W-1]|~brk_done_v[`W-1]|~op_T2_jsr_v[`W-1]|~op_rti_rts_v[`W-1]|~n389_v[`W-1]), n1649_v, n1649_i3);
  spice_transistor_nmos_vdd t196(~n1720_v[`W-1], n612_v, n612_i0);
  spice_transistor_nmos_vdd t2779(~abh1_v[`W-1], n1140_v, n1140_i1);
  spice_transistor_nmos_vdd t197(~dor4_v[`W-1], n1076_v, n1076_i0);
  spice_transistor_nmos_gnd t192(~pch7_v[`W-1], n453_v, n453_i0);
  spice_transistor_nmos_gnd t52(~n593_v[`W-1], dpc4_SSB_v, dpc4_SSB_i0);
  spice_transistor_nmos t53(~dpc11_SBADD_v[`W-1], alua0_v, dasb0_v, alua0_i0, dasb0_i0);
  spice_transistor_nmos t55(~dpc11_SBADD_v[`W-1], alua5_v, sb5_v, alua5_i0, sb5_i0);
  spice_transistor_nmos t56(~dpc11_SBADD_v[`W-1], alua6_v, sb6_v, alua6_i0, sb6_i0);
  spice_transistor_nmos_gnd t60(~pch3_v[`W-1], n923_v, n923_i0);
  spice_transistor_nmos_gnd t190(~ir3_v[`W-1], notir3_v, notir3_i0);
  spice_transistor_nmos_gnd t3237(~NMIP_v[`W-1], n645_v, n645_i1);
  spice_transistor_nmos_gnd t2050(~n1346_v[`W-1], n1296_v, n1296_i2);
  spice_transistor_nmos_gnd t3235(~n1640_v[`W-1], n1251_v, n1251_i2);
  spice_transistor_nmos t191(~cclk_v[`W-1], n1609_v, notir5_v, n1609_i0, notir5_i0);
  spice_transistor_nmos t3233(~cclk_v[`W-1], a4_v, n1344_v, a4_i2, n1344_i3);
  spice_transistor_nmos_vdd t2051(~n1346_v[`W-1], n359_v, n359_i2);
  spice_transistor_nmos t2053(~dpc19_ADDSB7_v[`W-1], alu7_v, sb7_v, alu7_i1, sb7_i6);
  spice_transistor_nmos_gnd g_1362((~n320_v[`W-1]|~n36_v[`W-1]), n735_v, n735_i1);
  spice_transistor_nmos_gnd t3309(~n1561_v[`W-1], n871_v, n871_i2);
  spice_transistor_nmos_vdd t299(~cclk_v[`W-1], adh0_v, adh0_i1);
  spice_transistor_nmos_gnd t295(~s6_v[`W-1], n1187_v, n1187_i0);
  spice_transistor_nmos_gnd t297(~pd7_clearIR_v[`W-1], n1605_v, n1605_i0);
  spice_transistor_nmos t296(~cp1_v[`W-1], n719_v, idl0_v, n719_i1, idl0_i0);
  spice_transistor_nmos_gnd t290(~_ABL6_v[`W-1], abl7_v, abl7_i0);
  spice_transistor_nmos_gnd t293(~n1413_v[`W-1], dpc32_PCHADH_v, dpc32_PCHADH_i0);
  spice_transistor_nmos_gnd t3056(~AxB1_v[`W-1], n953_v, n953_i1);
  spice_transistor_nmos_vdd t3492(~n6_v[`W-1], dpc6_SBS_v, dpc6_SBS_i8);
  spice_transistor_nmos_gnd t3491(~n6_v[`W-1], n282_v, n282_i0);
  spice_transistor_nmos_gnd t3497(~n678_v[`W-1], t3_v, t3_i1);
  spice_transistor_nmos_gnd t3496(~x6_v[`W-1], n730_v, n730_i1);
  spice_transistor_nmos_gnd t3495(~idb1_v[`W-1], n583_v, n583_i1);
  spice_transistor_nmos t3499(~cclk_v[`W-1], pd0_v, n93_v, pd0_i0, n93_i1);
  spice_transistor_nmos t3498(~cclk_v[`W-1], pd1_v, n1319_v, pd1_i0, n1319_i1);
  spice_transistor_nmos_gnd g_1083((~n323_v[`W-1]|~n671_v[`W-1]|~Reset0_v[`W-1]), n14_v, n14_i2);
  spice_transistor_nmos_vdd t3504(~cclk_v[`W-1], idb4_v, idb4_i9);
  spice_transistor_nmos_gnd t2780(~n1409_v[`W-1], n1231_v, n1231_i1);
  spice_transistor_nmos_gnd t2782(~sb5_v[`W-1], n1135_v, n1135_i0);
  spice_transistor_nmos t2785(~cclk_v[`W-1], _ABL4_v, n86_v, _ABL4_i1, n86_i2);
  spice_transistor_nmos_gnd t2786(~n70_v[`W-1], n1117_v, n1117_i1);
  spice_transistor_nmos_gnd t2018(~n636_v[`W-1], nnT2BR_v, nnT2BR_i0);
  spice_transistor_nmos_vdd t2019(~n855_v[`W-1], ab0_v, ab0_i1);
  spice_transistor_nmos_gnd g_1080((~n288_v[`W-1]|~RnWstretched_v[`W-1]), n798_v, n798_i2);
  spice_transistor_nmos_gnd t3013(~n717_v[`W-1], C1x5Reset_v, C1x5Reset_i1);
  spice_transistor_nmos t3012(~cp1_v[`W-1], n1291_v, brk_done_v, n1291_i0, brk_done_i0);
  spice_transistor_nmos t2548(~dpc32_PCHADH_v[`W-1], adh6_v, n652_v, adh6_i5, n652_i2);
  spice_transistor_nmos t2549(~dpc32_PCHADH_v[`W-1], adh5_v, n1301_v, adh5_i4, n1301_i2);
  spice_transistor_nmos t3503(~cclk_v[`W-1], n1190_v, nots2_v, n1190_i1, nots2_i1);
  spice_transistor_nmos_vdd t3502(~cclk_v[`W-1], sb2_v, sb2_i12);
  spice_transistor_nmos_gnd g_1380((~ir6_v[`W-1]|~notir1_v[`W-1]|~ir7_v[`W-1]), op_shift_v, op_shift_i1);
  spice_transistor_nmos_gnd g_1381((~notir6_v[`W-1]|~notir1_v[`W-1]), op_lsr_ror_dec_inc_v, op_lsr_ror_dec_inc_i2);
  spice_transistor_nmos_gnd g_1382((~clearIR_v[`W-1]|~pd7_v[`W-1]), pd7_clearIR_v, pd7_clearIR_i3);
  spice_transistor_nmos_gnd g_1383((~brk_done_v[`W-1]|~n717_v[`W-1]), n1087_v, n1087_i2);
  spice_transistor_nmos_gnd g_1384((~pd0_clearIR_v[`W-1]|~pd2_clearIR_v[`W-1]|~n1083_v[`W-1]), PD_xxxx10x0_v, PD_xxxx10x0_i2);
  spice_transistor_nmos_gnd g_1386((~n470_v[`W-1]|~n134_v[`W-1]), n467_v, n467_i3);
  spice_transistor_nmos_gnd g_1387((~n812_v[`W-1]|~n31_v[`W-1]), n1044_v, n1044_i1);
  spice_transistor_nmos_gnd g_1388((~n43_v[`W-1]|~n360_v[`W-1]), n1230_v, n1230_i3);
  spice_transistor_nmos_gnd g_1389((~RnWstretched_v[`W-1]|~dor7_v[`W-1]), n23_v, n23_i2);
  spice_transistor_nmos g_1434((~ADL_ABL_v[`W-1]&~cp1_v[`W-1]), _ABL4_v, n1519_v, _ABL4_i2, n1519_i2);
  spice_transistor_nmos g_1435((~ADL_ABL_v[`W-1]&~cp1_v[`W-1]), _ABL7_v, n1046_v, _ABL7_i2, n1046_i2);
  spice_transistor_nmos g_1433((~ADL_ABL_v[`W-1]&~cp1_v[`W-1]), _ABL6_v, n1548_v, _ABL6_i2, n1548_i2);
  spice_transistor_nmos g_1430((~ADL_ABL_v[`W-1]&~cp1_v[`W-1]), _ABL3_v, n1507_v, _ABL3_i2, n1507_i2);
  spice_transistor_nmos_gnd g_1431((~n790_v[`W-1]&~_op_store_v[`W-1]), n1137_v, n1137_i2);
  spice_transistor_nmos_gnd t3163(~n617_v[`W-1], n1140_v, n1140_i2);
  spice_transistor_nmos_gnd t3161(~n1398_v[`W-1], A_B7_v, A_B7_i0);
  spice_transistor_nmos_gnd t3167(~x_op_T0_bit_v[`W-1], n1379_v, n1379_i1);
  spice_transistor_nmos_gnd t3166(~n1625_v[`W-1], n90_v, n90_i2);
  spice_transistor_nmos_gnd t3164(~n1527_v[`W-1], n1295_v, n1295_i2);
  spice_transistor_nmos_gnd g_1218((~n236_v[`W-1]|~nnT2BR_v[`W-1]), n1427_v, n1427_i2);
  spice_transistor_nmos_gnd g_1168((~ir2_v[`W-1]|~ir4_v[`W-1]|~irline3_v[`W-1]|~notir3_v[`W-1]|~ir7_v[`W-1]), x_op_push_pull_v, x_op_push_pull_i1);
  spice_transistor_nmos_gnd t3500(~n951_v[`W-1], n1152_v, n1152_i2);
  spice_transistor_nmos_gnd g_1652(((~C45_v[`W-1]&~A_B5_v[`W-1])|~n647_v[`W-1]), _C56_v, _C56_i2);
  spice_transistor_nmos_gnd g_1653((~n1316_v[`W-1]|(~n232_v[`W-1]&~n344_v[`W-1])), n20_v, n20_i2);
  spice_transistor_nmos_gnd g_1650((~n1115_v[`W-1]|(~n620_v[`W-1]&~n270_v[`W-1])), BRtaken_v, BRtaken_i2);
  spice_transistor_nmos_gnd g_1651(((~pipeT3out_v[`W-1]&~n16_v[`W-1])|(~pipeT4out_v[`W-1]&~notRdy0_v[`W-1])), n472_v, n472_i2);
  spice_transistor_nmos_gnd g_1656((~n810_v[`W-1]|(~n293_v[`W-1]&~n923_v[`W-1])), n207_v, n207_i2);
  spice_transistor_nmos_gnd g_1657((~_AxB_0__C0in_v[`W-1]|(~n105_v[`W-1]&~__AxB_0_v[`W-1])), __AxBxC_0_v, __AxBxC_0_i2);
  spice_transistor_nmos_gnd g_1654((~n1097_v[`W-1]|(~n345_v[`W-1]&~n432_v[`W-1])), dasb3_v, dasb3_i2);
  spice_transistor_nmos_gnd g_1655(((~n646_v[`W-1]|~n1655_v[`W-1]|~op_T5_rts_v[`W-1])|(~n236_v[`W-1]&~n1262_v[`W-1])), n182_v, n182_i4);
  spice_transistor_nmos_gnd g_1065((~ir2_v[`W-1]|~notir4_v[`W-1]|~clock1_v[`W-1]|~notir3_v[`W-1]|~ir7_v[`W-1]|~notir6_v[`W-1]|~irline3_v[`W-1]), op_T0_cli_sei_v, op_T0_cli_sei_i2);
  spice_transistor_nmos_gnd t518(~ir6_v[`W-1], notir6_v, notir6_i0);
  spice_transistor_nmos_gnd t519(~n1225_v[`W-1], n1222_v, n1222_i0);
  spice_transistor_nmos_gnd t512(~nots4_v[`W-1], n3_v, n3_i2);
  spice_transistor_nmos_gnd t510(~op_T2_jsr_v[`W-1], n383_v, n383_i0);
  spice_transistor_nmos_gnd t516(~n1223_v[`W-1], n225_v, n225_i0);
  spice_transistor_nmos_vdd t517(~n1223_v[`W-1], dpc9_DBADD_v, dpc9_DBADD_i1);
  spice_transistor_nmos_gnd t514(~pipeUNK06_v[`W-1], n755_v, n755_i0);
  spice_transistor_nmos t515(~cclk_v[`W-1], n496_v, nots5_v, n496_i0, nots5_i1);
  spice_transistor_nmos_gnd t2767(~n1026_v[`W-1], n322_v, n322_i2);
  spice_transistor_nmos_vdd t2764(~n611_v[`W-1], dpc31_PCHPCH_v, dpc31_PCHPCH_i8);
  spice_transistor_nmos t2762(~cp1_v[`W-1], n1661_v, idl3_v, n1661_i3, idl3_i1);
  spice_transistor_nmos_gnd t2763(~n611_v[`W-1], n255_v, n255_i0);
  spice_transistor_nmos_gnd t2760(~pd4_clearIR_v[`W-1], n227_v, n227_i0);
  spice_transistor_nmos_vdd t1894(~n102_v[`W-1], rw_v, rw_i0);
  spice_transistor_nmos_vdd t2768(~n1026_v[`W-1], n171_v, n171_i3);
  spice_transistor_nmos_vdd t1410(~n321_v[`W-1], dpc33_PCHDB_v, dpc33_PCHDB_i0);
  spice_transistor_nmos_gnd g_1103((~ir2_v[`W-1]|~notir6_v[`W-1]|~ir7_v[`W-1]|~ir4_v[`W-1]|~notir1_v[`W-1]|~clock1_v[`W-1]|~notir3_v[`W-1]), op_T0_shift_right_a_v, op_T0_shift_right_a_i1);
  spice_transistor_nmos_gnd g_1100((~op_lsr_ror_dec_inc_v[`W-1]|~op_asl_rol_v[`W-1]), n790_v, n790_i3);
  spice_transistor_nmos t682(~cclk_v[`W-1], pipeUNK31_v, n389_v, pipeUNK31_i0, n389_i0);
  spice_transistor_nmos_gnd g_1107((~ir3_v[`W-1]|~ir7_v[`W-1]|~irline3_v[`W-1]|~clock1_v[`W-1]|~ir4_v[`W-1]|~ir5_v[`W-1]|~ir2_v[`W-1]), op_T0_brk_rti_v, op_T0_brk_rti_i1);
  spice_transistor_nmos_gnd t994(~op_clv_v[`W-1], n340_v, n340_i0);
  spice_transistor_nmos_gnd t992(~abh5_v[`W-1], n869_v, n869_i1);
  spice_transistor_nmos_vdd t990(~abh5_v[`W-1], n1608_v, n1608_i1);
  spice_transistor_nmos t1309(~cclk_v[`W-1], n889_v, pipeUNK42_v, n889_i0, pipeUNK42_i0);
  spice_transistor_nmos t1308(~dpc10_ADLADD_v[`W-1], adl2_v, alub2_v, adl2_i1, alub2_i1);
  spice_transistor_nmos_gnd t683(~pcl3_v[`W-1], n249_v, n249_i0);
  spice_transistor_nmos_gnd t998(~n415_v[`W-1], n931_v, n931_i1);
  spice_transistor_nmos_gnd t999(~n88_v[`W-1], n1375_v, n1375_i0);
  spice_transistor_nmos t2631(~cp1_v[`W-1], notRnWprepad_v, n1579_v, notRnWprepad_i1, n1579_i1);
  spice_transistor_nmos t1529(~dpc3_SBX_v[`W-1], x5_v, sb5_v, x5_i1, sb5_i4);
  spice_transistor_nmos t1528(~dpc3_SBX_v[`W-1], sb6_v, x6_v, sb6_i7, x6_i1);
  spice_transistor_nmos_vdd t1521(~n1677_v[`W-1], n999_v, n999_i1);
  spice_transistor_nmos_gnd t1520(~n1677_v[`W-1], n475_v, n475_i0);
  spice_transistor_nmos t1523(~dpc3_SBX_v[`W-1], dasb4_v, x4_v, dasb4_i6, x4_i0);
  spice_transistor_nmos t1522(~cclk_v[`W-1], n865_v, n958_v, n865_i0, n958_i1);
  spice_transistor_nmos t1525(~dpc3_SBX_v[`W-1], x2_v, sb2_v, x2_i1, sb2_i4);
  spice_transistor_nmos t1524(~dpc3_SBX_v[`W-1], x3_v, sb3_v, x3_i1, sb3_i6);
  spice_transistor_nmos_vdd t1527(~n582_v[`W-1], ADH_ABH_v, ADH_ABH_i0);
  spice_transistor_nmos_gnd t1526(~n582_v[`W-1], n1067_v, n1067_i0);
  spice_transistor_nmos t2877(~cclk_v[`W-1], n799_v, n264_v, n799_i1, n264_i0);
  spice_transistor_nmos_gnd t1901(~C67_v[`W-1], _C67_v, _C67_i0);
  spice_transistor_nmos_gnd t1907(~n1020_v[`W-1], n1277_v, n1277_i0);
  spice_transistor_nmos_gnd t1906(~s7_v[`W-1], n548_v, n548_i0);
  spice_transistor_nmos t2733(~cclk_v[`W-1], _ABH2_v, n994_v, _ABH2_i1, n994_i2);
  spice_transistor_nmos_gnd t2732(~op_T0_tsx_v[`W-1], n1586_v, n1586_i1);
  spice_transistor_nmos_gnd g_1424((~n410_v[`W-1]&~n392_v[`W-1]), n344_v, n344_i2);
  spice_transistor_nmos_gnd t199(~n982_v[`W-1], n1141_v, n1141_i1);
  spice_transistor_nmos_gnd t64(~notalu6_v[`W-1], alu6_v, alu6_i0);
  spice_transistor_nmos_gnd t67(~notidl2_v[`W-1], idl2_v, idl2_i0);
  spice_transistor_nmos t63(~cclk_v[`W-1], n1347_v, n1527_v, n1347_i0, n1527_i0);
  spice_transistor_nmos t3228(~cclk_v[`W-1], n1374_v, n1252_v, n1374_i0, n1252_i0);
  spice_transistor_nmos_gnd t358(~idb0_v[`W-1], n1224_v, n1224_i0);
  spice_transistor_nmos_gnd t356(~n1341_v[`W-1], n600_v, n600_i0);
  spice_transistor_nmos_gnd t350(~n66_v[`W-1], ab1_v, ab1_i0);
  spice_transistor_nmos t3225(~dpc2_XSB_v[`W-1], n1709_v, sb1_v, n1709_i2, sb1_i12);
  spice_transistor_nmos_gnd t3226(~n669_v[`W-1], op_ANDS_v, op_ANDS_i1);
  spice_transistor_nmos_gnd g_1084((~n917_v[`W-1]|~op_T0_txs_v[`W-1]|~n1109_v[`W-1]), n1358_v, n1358_i3);
  spice_transistor_nmos_gnd t1919(~n127_v[`W-1], n135_v, n135_i2);
  spice_transistor_nmos_gnd t3314(~s1_v[`W-1], n1711_v, n1711_i1);
  spice_transistor_nmos t3316(~cclk_v[`W-1], y0_v, n564_v, y0_i2, n564_i2);
  spice_transistor_nmos t3317(~cclk_v[`W-1], n659_v, _ABH7_v, n659_i3, _ABH7_i1);
  spice_transistor_nmos_vdd t3313(~n1463_v[`W-1], n147_v, n147_i1);
  spice_transistor_nmos_gnd g_1616(((~_TWOCYCLE_phi1_v[`W-1]&~n1528_v[`W-1])|~n1161_v[`W-1]), n732_v, n732_i3);
  spice_transistor_nmos_gnd g_1366((~ir6_v[`W-1]|~ir7_v[`W-1]|~notir0_v[`W-1]|~notir5_v[`W-1]|~clock1_v[`W-1]), op_T0_and_v, op_T0_and_i1);

  spice_pullup p_888(n1640_v, n1640_i2);
  spice_pullup p_283(aluanorb0_v, aluanorb0_i2);
  spice_pullup p_715(pd7_clearIR_v, pd7_clearIR_i1);
  spice_pullup p_825(n133_v, n133_i2);
  spice_pullup p_192(n1159_v, n1159_i0);
  spice_pullup p_828(n130_v, n130_i2);
  spice_pullup p_1000(n1293_v, n1293_i0);
  spice_pullup p_1001(n1290_v, n1290_i1);
  spice_pullup p_1004(n474_v, n474_i1);
  spice_pullup p_309(n1718_v, n1718_i2);
  spice_pullup p_308(n1719_v, n1719_i2);
  spice_pullup p_6(n299_v, n299_i1);
  spice_pullup p_4(op_T4_v, op_T4_i1);
  spice_pullup p_5(x_op_T3_ind_y_v, x_op_T3_ind_y_i0);
  spice_pullup p_0(n344_v, n344_i0);
  spice_pullup p_233(op_T5_rts_v, op_T5_rts_i0);
  spice_pullup p_232(n818_v, n818_i2);
  spice_pullup p_231(n1526_v, n1526_i2);
  spice_pullup p_230(__AxB_0_v, __AxB_0_i1);
  spice_pullup p_541(n1491_v, n1491_i3);
  spice_pullup p_543(x_op_T0_bit_v, x_op_T0_bit_i1);
  spice_pullup p_545(dasb3_v, dasb3_i1);
  spice_pullup p_544(n1474_v, n1474_i2);
  spice_pullup p_547(n1304_v, n1304_i1);
  spice_pullup p_405(n637_v, n637_i0);
  spice_pullup p_787(n441_v, n441_i1);
  spice_pullup p_786(n442_v, n442_i2);
  spice_pullup p_783(n1401_v, n1401_i1);
  spice_pullup p_782(n1402_v, n1402_i1);
  spice_pullup p_781(n1408_v, n1408_i0);
  spice_pullup p_780(dor4_v, dor4_i2);
  spice_pullup p_905(op_T3_ind_x_v, op_T3_ind_x_i0);
  spice_pullup p_9(n293_v, n293_i0);
  spice_pullup p_904(abh0_v, abh0_i4);
  spice_pullup p_169(n256_v, n256_i0);
  spice_pullup p_493(abh7_v, abh7_i4);
  spice_pullup p_492(op_T0_cmp_v, op_T0_cmp_i0);
  spice_pullup p_491(n1357_v, n1357_i1);
  spice_pullup p_497(n485_v, n485_i2);
  spice_pullup p_496(__AxBxC_5_v, __AxBxC_5_i1);
  spice_pullup p_494(n488_v, n488_i4);
  spice_pullup p_499(n480_v, n480_i0);
  spice_pullup p_498(n481_v, n481_i4);
  spice_pullup p_525(n747_v, n747_i3);
  spice_pullup p_420(n213_v, n213_i2);
  spice_pullup p_7(n297_v, n297_i0);
  spice_pullup p_89(op_T5_brk_v, op_T5_brk_i1);
  spice_pullup p_88(__AxBxC_0_v, __AxBxC_0_i1);
  spice_pullup p_83(n1343_v, n1343_i0);
  spice_pullup p_82(n409_v, n409_i1);
  spice_pullup p_81(op_T0_acc_v, op_T0_acc_i0);
  spice_pullup p_80(n1219_v, n1219_i2);
  spice_pullup p_87(n378_v, n378_i2);
  spice_pullup p_86(dpc36_IPC_v, dpc36_IPC_i0);
  spice_pullup p_85(n1347_v, n1347_i1);
  spice_pullup p_84(n1346_v, n1346_i3);
  spice_pullup p_909(n732_v, n732_i0);
  spice_pullup p_767(n1065_v, n1065_i2);
  spice_pullup p_763(op_T2_jsr_v, op_T2_jsr_i1);
  spice_pullup p_908(n733_v, n733_i3);
  spice_pullup p_822(n946_v, n946_i0);
  spice_pullup p_823(n947_v, n947_i2);
  spice_pullup p_820(n8_v, n8_i1);
  spice_pullup p_821(n1462_v, n1462_i2);
  spice_pullup p_826(n132_v, n132_i2);
  spice_pullup p_827(op_T0_pla_v, op_T0_pla_i0);
  spice_pullup p_44(n1192_v, n1192_i1);
  spice_pullup p_42(n1190_v, n1190_i2);
  spice_pullup p_3(n340_v, n340_i2);
  spice_pullup p_1008(n1717_v, n1717_i1);
  spice_pullup p_40(n1439_v, n1439_i2);
  spice_pullup p_421(n218_v, n218_i1);
  spice_pullup p_412(n1101_v, n1101_i1);
  spice_pullup p_361(C1x5Reset_v, C1x5Reset_i2);
  spice_pullup p_958(n986_v, n986_i0);
  spice_pullup p_360(_op_store_v, _op_store_i1);
  spice_pullup p_956(n980_v, n980_i1);
  spice_pullup p_954(n988_v, n988_i1);
  spice_pullup p_955(n983_v, n983_i2);
  spice_pullup p_952(n1566_v, n1566_i3);
  spice_pullup p_363(n831_v, n831_i4);
  spice_pullup p_1(n345_v, n345_i0);
  spice_pullup p_365(n834_v, n834_i4);
  spice_pullup p_364(n837_v, n837_i2);
  spice_pullup p_408(n1376_v, n1376_i2);
  spice_pullup p_367(n839_v, n839_i2);
  spice_pullup p_960(op_T0_ldx_tax_tsx_v, op_T0_ldx_tax_tsx_i0);
  spice_pullup p_366(n838_v, n838_i1);
  spice_pullup p_911(n739_v, n739_i0);
  spice_pullup p_917(n1356_v, n1356_i2);
  spice_pullup p_660(op_T0_cpx_cpy_inx_iny_v, op_T0_cpx_cpy_inx_iny_i0);
  spice_pullup p_914(_WR_v, _WR_i1);
  spice_pullup p_661(n630_v, n630_i1);
  spice_pullup p_915(INTG_v, INTG_i1);
  spice_pullup p_662(n631_v, n631_i3);
  spice_pullup p_664(n964_v, n964_i0);
  spice_pullup p_918(n462_v, n462_i2);
  spice_pullup p_665(__AxBxC_1_v, __AxBxC_1_i1);
  spice_pullup p_919(op_T0_v, op_T0_i2);
  spice_pullup p_669(n962_v, n962_i1);
  spice_pullup p_1010(n1715_v, n1715_i3);
  spice_pullup p_1013(n477_v, n477_i3);
  spice_pullup p_1012(n1364_v, n1364_i3);
  spice_pullup p_1015(n479_v, n479_i0);
  spice_pullup p_634(n1267_v, n1267_i1);
  spice_pullup p_103(n243_v, n243_i1);
  spice_pullup p_102(idl5_v, idl5_i2);
  spice_pullup p_558(n490_v, n490_i2);
  spice_pullup p_559(n491_v, n491_i1);
  spice_pullup p_790(op_T5_rti_rts_v, op_T5_rti_rts_i0);
  spice_pullup p_791(n445_v, n445_i4);
  spice_pullup p_792(dor3_v, dor3_i2);
  spice_pullup p_793(op_plp_pla_v, op_plp_pla_i0);
  spice_pullup p_794(n1542_v, n1542_i0);
  spice_pullup p_796(pclp4_v, pclp4_i2);
  spice_pullup p_797(n38_v, n38_i2);
  spice_pullup p_798(op_from_x_v, op_from_x_i0);
  spice_pullup p_710(n674_v, n674_i2);
  spice_pullup p_741(PD_xxx010x1_v, PD_xxx010x1_i0);
  spice_pullup p_514(t5_v, t5_i1);
  spice_pullup p_315(n1137_v, n1137_i0);
  spice_pullup p_310(n1270_v, n1270_i2);
  spice_pullup p_311(n1271_v, n1271_i2);
  spice_pullup p_312(n1138_v, n1138_i2);
  spice_pullup p_313(n1133_v, n1133_i1);
  spice_pullup p_515(n854_v, n854_i1);
  spice_pullup p_629(n669_v, n669_i1);
  spice_pullup p_174(n169_v, n169_i1);
  spice_pullup p_170(op_T0_tya_v, op_T0_tya_i0);
  spice_pullup p_171(n254_v, n254_i1);
  spice_pullup p_172(n255_v, n255_i1);
  spice_pullup p_173(n168_v, n168_i1);
  spice_pullup p_488(n1449_v, n1449_i1);
  spice_pullup p_489(n1448_v, n1448_i1);
  spice_pullup p_484(n1117_v, n1117_i2);
  spice_pullup p_485(idl3_v, idl3_i2);
  spice_pullup p_486(Pout4_v, Pout4_i2);
  spice_pullup p_487(n467_v, n467_i0);
  spice_pullup p_480(n1110_v, n1110_i3);
  spice_pullup p_481(ir4_v, ir4_i2);
  spice_pullup p_482(n1115_v, n1115_i0);
  spice_pullup p_483(op_T0_clc_sec_v, op_T0_clc_sec_i1);
  spice_pullup p_746(n470_v, n470_i1);
  spice_pullup p_1003(n1295_v, n1295_i3);
  spice_pullup p_972(alu2_v, alu2_i4);
  spice_pullup p_745(n473_v, n473_i1);
  spice_pullup p_726(ir5_v, ir5_i2);
  spice_pullup p_1005(n1712_v, n1712_i1);
  spice_pullup p_130(aluaorb0_v, aluaorb0_i1);
  spice_pullup p_865(n326_v, n326_i4);
  spice_pullup p_220(n224_v, n224_i1);
  spice_pullup p_819(n1026_v, n1026_i3);
  spice_pullup p_818(n332_v, n332_i4);
  spice_pullup p_813(ir6_v, ir6_i3);
  spice_pullup p_812(n334_v, n334_i3);
  spice_pullup p_838(n80_v, n80_i1);
  spice_pullup p_969(n484_v, n484_i1);
  spice_pullup p_963(n110_v, n110_i1);
  spice_pullup p_961(A_B7_v, A_B7_i1);
  spice_pullup p_967(n1631_v, n1631_i1);
  spice_pullup p_966(_DBE_v, _DBE_i0);
  spice_pullup p_965(n118_v, n118_i1);
  spice_pullup p_616(n1043_v, n1043_i1);
  spice_pullup p_784(n1400_v, n1400_i2);
  spice_pullup p_427(n916_v, n916_i1);
  spice_pullup p_613(n70_v, n70_i1);
  spice_pullup p_619(n1046_v, n1046_i1);
  spice_pullup p_618(n1047_v, n1047_i1);
  spice_pullup p_303(n1488_v, n1488_i1);
  spice_pullup p_789(x_op_T3_abs_idx_v, x_op_T3_abs_idx_i0);
  spice_pullup p_900(op_T0_lda_v, op_T0_lda_i1);
  spice_pullup p_302(n1484_v, n1484_i2);
  spice_pullup p_301(n1486_v, n1486_i1);
  spice_pullup p_300(op_T3_plp_pla_v, op_T3_plp_pla_i0);
  spice_pullup p_306(op_push_pull_v, op_push_pull_i0);
  spice_pullup p_882(PD_n_0xx0xx0x_v, PD_n_0xx0xx0x_i1);
  spice_pullup p_305(n795_v, n795_i2);
  spice_pullup p_239(__AxB5__C45_v, __AxB5__C45_i0);
  spice_pullup p_304(n797_v, n797_i2);
  spice_pullup p_8(__AxB1__C01_v, __AxB1__C01_i0);
  spice_pullup p_509(_DA_ADD1_v, _DA_ADD1_i2);
  spice_pullup p_132(op_asl_rol_v, op_asl_rol_i0);
  spice_pullup p_2(n347_v, n347_i0);
  spice_pullup p_160(n385_v, n385_i1);
  spice_pullup p_565(n21_v, n21_i2);
  spice_pullup p_563(n27_v, n27_i4);
  spice_pullup p_562(notir4_v, notir4_i2);
  spice_pullup p_769(idl2_v, idl2_i2);
  spice_pullup p_768(n1067_v, n1067_i2);
  spice_pullup p_765(n1069_v, n1069_i1);
  spice_pullup p_764(op_T3_branch_v, op_T3_branch_i1);
  spice_pullup p_201(pchp7_v, pchp7_i2);
  spice_pullup p_766(n1063_v, n1063_i2);
  spice_pullup p_761(n714_v, n714_i2);
  spice_pullup p_760(n715_v, n715_i1);
  spice_pullup p_762(abh1_v, abh1_i4);
  spice_pullup p_707(n1090_v, n1090_i1);
  spice_pullup p_369(op_T5_rti_v, op_T5_rti_i0);
  spice_pullup p_109(n176_v, n176_i1);
  spice_pullup p_108(n177_v, n177_i2);
  spice_pullup p_236(n812_v, n812_i0);
  spice_pullup p_234(n810_v, n810_i0);
  spice_pullup p_307(n790_v, n790_i1);
  spice_pullup p_279(n233_v, n233_i0);
  spice_pullup p_540(n617_v, n617_i3);
  spice_pullup p_615(C34_v, C34_i1);
  spice_pullup p_614(n79_v, n79_i1);
  spice_pullup p_617(H1x1_v, H1x1_i8);
  spice_pullup p_542(n1471_v, n1471_i2);
  spice_pullup p_611(n72_v, n72_i4);
  spice_pullup p_446(n1595_v, n1595_i1);
  spice_pullup p_612(n71_v, n71_i1);
  spice_pullup p_278(n232_v, n232_i1);
  spice_pullup p_585(n184_v, n184_i2);
  spice_pullup p_584(notRnWprepad_v, notRnWprepad_i3);
  spice_pullup p_587(n1464_v, n1464_i0);
  spice_pullup p_586(n188_v, n188_i2);
  spice_pullup p_581(n979_v, n979_i1);
  spice_pullup p_580(t2_v, t2_i2);
  spice_pullup p_583(n180_v, n180_i0);
  spice_pullup p_804(n34_v, n34_i2);
  spice_pullup p_546(op_T0_brk_rti_v, op_T0_brk_rti_i0);
  spice_pullup p_589(__AxB3__C23_v, __AxB3__C23_i0);
  spice_pullup p_588(n861_v, n861_i1);
  spice_pullup p_805(n641_v, n641_i2);
  spice_pullup p_549(idl4_v, idl4_i2);
  spice_pullup p_357(n929_v, n929_i4);
  spice_pullup p_806(AxB3_v, AxB3_i1);
  spice_pullup p_548(n1305_v, n1305_i2);
  spice_pullup p_503(n191_v, n191_i1);
  spice_pullup p_808(n647_v, n647_i1);
  spice_pullup p_809(op_shift_right_v, op_shift_right_i0);
  spice_pullup p_439(n662_v, n662_i1);
  spice_pullup p_800(n31_v, n31_i4);
  spice_pullup p_802(n36_v, n36_i0);
  spice_pullup p_698(n1070_v, n1070_i1);
  spice_pullup p_807(n645_v, n645_i2);
  spice_pullup p_502(n196_v, n196_i2);
  spice_pullup p_438(pd3_clearIR_v, pd3_clearIR_i1);
  spice_pullup p_314(n1130_v, n1130_i1);
  spice_pullup p_839(op_T2_ind_x_v, op_T2_ind_x_i0);
  spice_pullup p_974(n568_v, n568_i2);
  spice_pullup p_426(n917_v, n917_i0);
  spice_pullup p_976(n565_v, n565_i2);
  spice_pullup p_970(dor2_v, dor2_i2);
  spice_pullup p_971(n1635_v, n1635_i2);
  spice_pullup p_978(n567_v, n567_i4);
  spice_pullup p_425(n918_v, n918_i1);
  spice_pullup p_422(op_T2_mem_zp_v, op_T2_mem_zp_i0);
  spice_pullup p_973(n1638_v, n1638_i2);
  spice_pullup p_423(op_T0_tay_v, op_T0_tay_i0);
  spice_pullup p_228(op_T2_ind_v, op_T2_ind_i0);
  spice_pullup p_352(n1573_v, n1573_i1);
  spice_pullup p_678(op_T__ora_and_eor_adc_v, op_T__ora_and_eor_adc_i0);
  spice_pullup p_355(n1575_v, n1575_i2);
  spice_pullup p_276(n236_v, n236_i2);
  spice_pullup p_1006(n1711_v, n1711_i2);
  spice_pullup p_570(n1087_v, n1087_i1);
  spice_pullup p_571(op_T2_pha_v, op_T2_pha_i0);
  spice_pullup p_574(n1083_v, n1083_i1);
  spice_pullup p_221(n221_v, n221_i1);
  spice_pullup p_577(n975_v, n975_i0);
  spice_pullup p_778(op_T0_jmp_v, op_T0_jmp_i0);
  spice_pullup p_776(_C67_v, _C67_i1);
  spice_pullup p_777(n595_v, n595_i1);
  spice_pullup p_774(n1660_v, n1660_i3);
  spice_pullup p_775(n593_v, n593_i2);
  spice_pullup p_772(op_T__inx_v, op_T__inx_i0);
  spice_pullup p_773(n1662_v, n1662_i1);
  spice_pullup p_770(n1668_v, n1668_i1);
  spice_pullup p_771(op_T__asl_rol_a_v, op_T__asl_rol_a_i0);
  spice_pullup p_163(n389_v, n389_i2);
  spice_pullup p_162(n388_v, n388_i0);
  spice_pullup p_222(n220_v, n220_i3);
  spice_pullup p_161(n386_v, n386_i2);
  spice_pullup p_372(n781_v, n781_i0);
  spice_pullup p_378(n1720_v, n1720_i1);
  spice_pullup p_877(n998_v, n998_i4);
  spice_pullup p_166(_op_set_C_v, _op_set_C_i1);
  spice_pullup p_703(so_v, so_i1);
  spice_pullup p_165(op_jsr_v, op_jsr_i0);
  spice_pullup p_223(n152_v, n152_i0);
  spice_pullup p_436(_op_branch_bit6_v, _op_branch_bit6_i2);
  spice_pullup p_164(op_T2_idx_x_xy_v, op_T2_idx_x_xy_i0);
  spice_pullup p_870(n1594_v, n1594_i1);
  spice_pullup p_118(n1618_v, n1618_i4);
  spice_pullup p_119(n1619_v, n1619_i0);
  spice_pullup p_873(abh6_v, abh6_i4);
  spice_pullup p_643(n1316_v, n1316_i0);
  spice_pullup p_168(n251_v, n251_i2);
  spice_pullup p_224(aluanorb1_v, aluanorb1_i2);
  spice_pullup p_646(A_B3_v, A_B3_i1);
  spice_pullup p_647(n1312_v, n1312_i0);
  spice_pullup p_644(n1315_v, n1315_i3);
  spice_pullup p_645(C67_v, C67_i1);
  spice_pullup p_335(n1229_v, n1229_i1);
  spice_pullup p_225(n154_v, n154_i3);
  spice_pullup p_608(Pout6_v, Pout6_i2);
  spice_pullup p_609(op_T0_dex_v, op_T0_dex_i0);
  spice_pullup p_596(n884_v, n884_i2);
  spice_pullup p_597(n889_v, n889_i2);
  spice_pullup p_285(n149_v, n149_i1);
  spice_pullup p_226(op_T2_stack_access_v, op_T2_stack_access_i0);
  spice_pullup p_592(n883_v, n883_i1);
  spice_pullup p_495(op_T2_brk_v, op_T2_brk_i0);
  spice_pullup p_590(n862_v, n862_i4);
  spice_pullup p_591(n867_v, n867_i1);
  spice_pullup p_1002(PD_1xx000x0_v, PD_1xx000x0_i0);
  spice_pullup p_598(n888_v, n888_i1);
  spice_pullup p_599(abh5_v, abh5_i4);
  spice_pullup p_196(n1153_v, n1153_i3);
  spice_pullup p_333(n629_v, n629_i1);
  spice_pullup p_533(n1697_v, n1697_i1);
  spice_pullup p_197(n1552_v, n1552_i2);
  spice_pullup p_330(n626_v, n626_i1);
  spice_pullup p_901(n1423_v, n1423_i3);
  spice_pullup p_58(n1281_v, n1281_i2);
  spice_pullup p_59(_C23_v, _C23_i1);
  spice_pullup p_54(n1178_v, n1178_i1);
  spice_pullup p_55(n510_v, n510_i0);
  spice_pullup p_56(n513_v, n513_i1);
  spice_pullup p_57(C01_v, C01_i1);
  spice_pullup p_50(_op_branch_bit7_v, _op_branch_bit7_i2);
  spice_pullup p_51(x_op_T0_tya_v, x_op_T0_tya_i0);
  spice_pullup p_52(n1170_v, n1170_i0);
  spice_pullup p_53(n1179_v, n1179_i1);
  spice_pullup p_348(n207_v, n207_i1);
  spice_pullup p_903(n1427_v, n1427_i1);
  spice_pullup p_907(n730_v, n730_i2);
  spice_pullup p_906(pclp6_v, pclp6_i2);
  spice_pullup p_863(n320_v, n320_i1);
  spice_pullup p_666(n966_v, n966_i3);
  spice_pullup p_667(nnT2BR_v, nnT2BR_i2);
  spice_pullup p_344(n1534_v, n1534_i2);
  spice_pullup p_722(notir7_v, notir7_i2);
  spice_pullup p_713(n673_v, n673_i0);
  spice_pullup p_131(t4_v, t4_i2);
  spice_pullup p_452(n1599_v, n1599_i2);
  spice_pullup p_450(n1593_v, n1593_i3);
  spice_pullup p_984(n1181_v, n1181_i1);
  spice_pullup p_18(n279_v, n279_i0);
  spice_pullup p_289(n931_v, n931_i2);
  spice_pullup p_135(n695_v, n695_i1);
  spice_pullup p_291(n937_v, n937_i1);
  spice_pullup p_290(n930_v, n930_i0);
  spice_pullup p_293(n935_v, n935_i1);
  spice_pullup p_292(n936_v, n936_i1);
  spice_pullup p_136(_DA_ADD2_v, _DA_ADD2_i1);
  spice_pullup p_296(D1x1_v, D1x1_i2);
  spice_pullup p_281(op_sta_cmp_v, op_sta_cmp_i0);
  spice_pullup p_286(aluvout_v, aluvout_i2);
  spice_pullup p_287(n933_v, n933_i0);
  spice_pullup p_347(op_T2_ADL_ADD_v, op_T2_ADL_ADD_i0);
  spice_pullup p_346(n200_v, n200_i0);
  spice_pullup p_137(n1548_v, n1548_i1);
  spice_pullup p_342(n16_v, n16_i1);
  spice_pullup p_341(n17_v, n17_i3);
  spice_pullup p_340(n14_v, n14_i1);
  spice_pullup p_127(DA_C45_v, DA_C45_i1);
  spice_pullup p_126(alucout_v, alucout_i2);
  spice_pullup p_125(n1141_v, n1141_i2);
  spice_pullup p_124(abh4_v, abh4_i4);
  spice_pullup p_123(n1610_v, n1610_i0);
  spice_pullup p_122(n1613_v, n1613_i1);
  spice_pullup p_121(op_T4_rts_v, op_T4_rts_i0);
  spice_pullup p_120(n1614_v, n1614_i0);
  spice_pullup p_129(n692_v, n692_i2);
  spice_pullup p_128(n1145_v, n1145_i1);
  spice_pullup p_182(op_sty_cpy_mem_v, op_sty_cpy_mem_i0);
  spice_pullup p_351(n208_v, n208_i4);
  spice_pullup p_700(n1676_v, n1676_i3);
  spice_pullup p_444(n755_v, n755_i1);
  spice_pullup p_799(pchp5_v, pchp5_i2);
  spice_pullup p_636(n1469_v, n1469_i2);
  spice_pullup p_638(n1018_v, n1018_i1);
  spice_pullup p_211(abh3_v, abh3_i4);
  spice_pullup p_210(n423_v, n423_i2);
  spice_pullup p_959(n987_v, n987_i2);
  spice_pullup p_213(n424_v, n424_i2);
  spice_pullup p_212(AxB1_v, AxB1_i1);
  spice_pullup p_575(n1082_v, n1082_i1);
  spice_pullup p_676(n875_v, n875_i1);
  spice_pullup p_49(n1175_v, n1175_i2);
  spice_pullup p_47(__AxBxC_6_v, __AxBxC_6_i1);
  spice_pullup p_46(n1194_v, n1194_i3);
  spice_pullup p_45(n1195_v, n1195_i3);
  spice_pullup p_43(n_0_ADL2_v, n_0_ADL2_i2);
  spice_pullup p_41(n1199_v, n1199_i2);
  spice_pullup p_824(n944_v, n944_i1);
  spice_pullup p_912(n1358_v, n1358_i2);
  spice_pullup p_913(n468_v, n468_i1);
  spice_pullup p_910(n735_v, n735_i0);
  spice_pullup p_916(x_op_T4_ind_y_v, x_op_T4_ind_y_i0);
  spice_pullup p_829(n134_v, n134_i0);
  spice_pullup p_801(n1541_v, n1541_i2);
  spice_pullup p_1007(op_T__cpx_cpy_imm_zp_v, op_T__cpx_cpy_imm_zp_i0);
  spice_pullup p_670(n969_v, n969_i1);
  spice_pullup p_950(n269_v, n269_i0);
  spice_pullup p_184(n1605_v, n1605_i1);
  spice_pullup p_951(op_xy_v, op_xy_i1);
  spice_pullup p_202(n533_v, n533_i2);
  spice_pullup p_353(_C45_v, _C45_i2);
  spice_pullup p_527(x_op_push_pull_v, x_op_push_pull_i0);
  spice_pullup p_254(n1120_v, n1120_i1);
  spice_pullup p_526(n748_v, n748_i1);
  spice_pullup p_200(op_lsr_ror_dec_inc_v, op_lsr_ror_dec_inc_i0);
  spice_pullup p_866(n327_v, n327_i1);
  spice_pullup p_867(op_inc_nop_v, op_inc_nop_i0);
  spice_pullup p_785(n1339_v, n1339_i2);
  spice_pullup p_207(n1399_v, n1399_i3);
  spice_pullup p_756(n1440_v, n1440_i1);
  spice_pullup p_757(n1260_v, n1260_i3);
  spice_pullup p_750(n951_v, n951_i3);
  spice_pullup p_751(op_T__cpx_cpy_abs_v, op_T__cpx_cpy_abs_i0);
  spice_pullup p_752(n953_v, n953_i2);
  spice_pullup p_753(n952_v, n952_i2);
  spice_pullup p_238(n815_v, n815_i2);
  spice_pullup p_205(n538_v, n538_i1);
  spice_pullup p_138(n1549_v, n1549_i2);
  spice_pullup p_139(n543_v, n543_i3);
  spice_pullup p_273(n432_v, n432_i1);
  spice_pullup p_229(BRtaken_v, BRtaken_i0);
  spice_pullup p_624(n1684_v, n1684_i2);
  spice_pullup p_625(n1687_v, n1687_i2);
  spice_pullup p_424(n919_v, n919_i0);
  spice_pullup p_622(_op_branch_done_v, _op_branch_done_i1);
  spice_pullup p_623(n1682_v, n1682_i1);
  spice_pullup p_891(n1649_v, n1649_i2);
  spice_pullup p_890(n1642_v, n1642_i0);
  spice_pullup p_957(n981_v, n981_i2);
  spice_pullup p_927(op_T4_brk_v, op_T4_brk_i0);
  spice_pullup p_280(n146_v, n146_i4);
  spice_pullup p_237(n813_v, n813_i0);
  spice_pullup p_899(Pout2_v, Pout2_i2);
  spice_pullup p_898(n1209_v, n1209_i1);
  spice_pullup p_626(op_EORS_v, op_EORS_i2);
  spice_pullup p_627(n1688_v, n1688_i2);
  spice_pullup p_620(n1045_v, n1045_i3);
  spice_pullup p_362(n830_v, n830_i2);
  spice_pullup p_621(n1044_v, n1044_i0);
  spice_pullup p_78(n400_v, n400_i3);
  spice_pullup p_79(n1379_v, n1379_i2);
  spice_pullup p_272(op_rmw_v, op_rmw_i1);
  spice_pullup p_72(n1222_v, n1222_i1);
  spice_pullup p_73(AxB5_v, AxB5_i1);
  spice_pullup p_70(n1224_v, n1224_i1);
  spice_pullup p_71(n1223_v, n1223_i2);
  spice_pullup p_76(n1374_v, n1374_i1);
  spice_pullup p_77(n1377_v, n1377_i1);
  spice_pullup p_74(DC34_v, DC34_i0);
  spice_pullup p_75(n1375_v, n1375_i2);
  spice_pullup p_453(n504_v, n504_i1);
  spice_pullup p_270(Pout3_v, Pout3_i2);
  spice_pullup p_277(n231_v, n231_i2);
  spice_pullup p_929(n350_v, n350_i3);
  spice_pullup p_928(n351_v, n351_i2);
  spice_pullup p_923(op_T2_abs_y_v, op_T2_abs_y_i0);
  spice_pullup p_922(n1517_v, n1517_i0);
  spice_pullup p_356(n928_v, n928_i1);
  spice_pullup p_748(n959_v, n959_i1);
  spice_pullup p_593(n882_v, n882_i0);
  spice_pullup p_788(n440_v, n440_i2);
  spice_pullup p_271(n436_v, n436_i3);
  spice_pullup p_368(n3_v, n3_i4);
  spice_pullup p_681(n1245_v, n1245_i1);
  spice_pullup p_953(t3_v, t3_i2);
  spice_pullup p_628(_DBZ_v, _DBZ_i1);
  spice_pullup p_977(n566_v, n566_i1);
  spice_pullup p_875(n990_v, n990_i3);
  spice_pullup p_721(n1323_v, n1323_i2);
  spice_pullup p_578(n973_v, n973_i2);
  spice_pullup p_724(op_T__shift_a_v, op_T__shift_a_i0);
  spice_pullup p_727(n5_v, n5_i2);
  spice_pullup p_579(n1081_v, n1081_i2);
  spice_pullup p_435(aluanandb1_v, aluanandb1_i3);
  spice_pullup p_434(n842_v, n842_i3);
  spice_pullup p_389(Pout7_v, Pout7_i2);
  spice_pullup p_216(dpc28_0ADH0_v, dpc28_0ADH0_i2);
  spice_pullup p_431(n846_v, n846_i1);
  spice_pullup p_430(n847_v, n847_i1);
  spice_pullup p_432(n845_v, n845_i1);
  spice_pullup p_871(n1592_v, n1592_i4);
  spice_pullup p_153(n1383_v, n1383_i2);
  spice_pullup p_569(n1709_v, n1709_i3);
  spice_pullup p_779(n1089_v, n1089_i2);
  spice_pullup p_659(dpc35_PCHC_v, dpc35_PCHC_i0);
  spice_pullup p_658(n1335_v, n1335_i1);
  spice_pullup p_218(n227_v, n227_i1);
  spice_pullup p_653(n318_v, n318_i3);
  spice_pullup p_652(n319_v, n319_i0);
  spice_pullup p_648(op_T4_rti_v, op_T4_rti_i0);
  spice_pullup p_872(n995_v, n995_i1);
  spice_pullup p_65(n_0_ADL1_v, n_0_ADL1_i2);
  spice_pullup p_64(Pout0_v, Pout0_i2);
  spice_pullup p_67(op_T0_tsx_v, op_T0_tsx_i1);
  spice_pullup p_66(n681_v, n681_i3);
  spice_pullup p_61(n1289_v, n1289_i1);
  spice_pullup p_60(fetch_v, fetch_i0);
  spice_pullup p_63(n689_v, n689_i1);
  spice_pullup p_69(op_T0_plp_v, op_T0_plp_i0);
  spice_pullup p_68(n458_v, n458_i2);
  spice_pullup p_316(n1135_v, n1135_i1);
  spice_pullup p_938(op_T2_zp_zp_idx_v, op_T2_zp_zp_idx_i0);
  spice_pullup p_939(n284_v, n284_i1);
  spice_pullup p_930(n358_v, n358_i3);
  spice_pullup p_931(n1033_v, n1033_i2);
  spice_pullup p_932(n1446_v, n1446_i1);
  spice_pullup p_933(n288_v, n288_i1);
  spice_pullup p_934(Pout1_v, Pout1_i2);
  spice_pullup p_935(op_T4_mem_abs_idx_v, op_T4_mem_abs_idx_i0);
  spice_pullup p_936(n280_v, n280_i4);
  spice_pullup p_937(n282_v, n282_i1);
  spice_pullup p_373(n782_v, n782_i0);
  spice_pullup p_370(op_T__dex_v, op_T__dex_i0);
  spice_pullup p_371(op_T0_sbc_v, op_T0_sbc_i0);
  spice_pullup p_376(op_T2_v, op_T2_i1);
  spice_pullup p_377(n789_v, n789_i2);
  spice_pullup p_374(n783_v, n783_i1);
  spice_pullup p_375(n1724_v, n1724_i3);
  spice_pullup p_642(PD_xxxx10x0_v, PD_xxxx10x0_i1);
  spice_pullup p_379(op_branch_done_v, op_branch_done_i1);
  spice_pullup p_113(n1500_v, n1500_i1);
  spice_pullup p_840(op_T0_cpx_inx_v, op_T0_cpx_inx_i0);
  spice_pullup p_841(n1650_v, n1650_i2);
  spice_pullup p_842(n1657_v, n1657_i1);
  spice_pullup p_843(n1654_v, n1654_i4);
  spice_pullup p_876(n992_v, n992_i1);
  spice_pullup p_699(n1561_v, n1561_i2);
  spice_pullup p_640(pd6_clearIR_v, pd6_clearIR_i1);
  spice_pullup p_925(n355_v, n355_i3);
  spice_pullup p_275(abl5_v, abl5_i4);
  spice_pullup p_848(n583_v, n583_i2);
  spice_pullup p_849(n588_v, n588_i2);
  spice_pullup p_610(n75_v, n75_i2);
  spice_pullup p_695(op_T0_shift_right_a_v, op_T0_shift_right_a_i0);
  spice_pullup p_554(n1309_v, n1309_i1);
  spice_pullup p_921(n1518_v, n1518_i1);
  spice_pullup p_694(clearIR_v, clearIR_i0);
  spice_pullup p_641(n1463_v, n1463_i1);
  spice_pullup p_705(abl0_v, abl0_i4);
  spice_pullup p_112(abl2_v, abl2_i4);
  spice_pullup p_235(n811_v, n811_i0);
  spice_pullup p_111(n172_v, n172_i3);
  spice_pullup p_114(_C01_v, _C01_i1);
  spice_pullup p_732(n1253_v, n1253_i0);
  spice_pullup p_733(abl3_v, abl3_i4);
  spice_pullup p_730(n1257_v, n1257_i0);
  spice_pullup p_736(op_T4_ind_x_v, op_T4_ind_x_i0);
  spice_pullup p_737(__AxB_4_v, __AxB_4_i1);
  spice_pullup p_734(n1251_v, n1251_i3);
  spice_pullup p_319(n519_v, n519_i3);
  spice_pullup p_738(op_T2_jmp_abs_v, op_T2_jmp_abs_i0);
  spice_pullup p_739(n300_v, n300_i1);
  spice_pullup p_398(C12_v, C12_i1);
  spice_pullup p_399(n503_v, n503_i2);
  spice_pullup p_428(alucin_v, alucin_i2);
  spice_pullup p_429(n913_v, n913_i2);
  spice_pullup p_394(n1038_v, n1038_i1);
  spice_pullup p_395(n404_v, n404_i2);
  spice_pullup p_396(NMIP_v, NMIP_i1);
  spice_pullup p_397(op_T0_ora_v, op_T0_ora_i0);
  spice_pullup p_390(op_T2_stack_v, op_T2_stack_i0);
  spice_pullup p_391(n1580_v, n1580_i1);
  spice_pullup p_392(n1586_v, n1586_i2);
  spice_pullup p_393(n1585_v, n1585_i2);
  spice_pullup p_181(n670_v, n670_i3);
  spice_pullup p_180(dasb6_v, dasb6_i1);
  spice_pullup p_183(n1600_v, n1600_i1);
  spice_pullup p_1011(n1714_v, n1714_i1);
  spice_pullup p_187(n803_v, n803_i1);
  spice_pullup p_186(alurawcout_v, alurawcout_i2);
  spice_pullup p_110(_AxB_6__C56_v, _AxB_6__C56_i0);
  spice_pullup p_649(n1319_v, n1319_i2);
  spice_pullup p_188(n800_v, n800_i1);
  spice_pullup p_902(_C34_v, _C34_i1);
  spice_pullup p_116(op_T0_and_v, op_T0_and_i0);
  spice_pullup p_10(n291_v, n291_i3);
  spice_pullup p_11(n270_v, n270_i1);
  spice_pullup p_12(op_T0_jsr_v, op_T0_jsr_i0);
  spice_pullup p_13(n272_v, n272_i2);
  spice_pullup p_14(op_T2_abs_access_v, op_T2_abs_access_i0);
  spice_pullup p_15(__AxBxC_3_v, __AxBxC_3_i1);
  spice_pullup p_16(n275_v, n275_i0);
  spice_pullup p_17(n278_v, n278_i2);
  spice_pullup p_19(n108_v, n108_i2);
  spice_pullup p_117(pclp0_v, pclp0_i2);
  spice_pullup p_350(n209_v, n209_i4);
  spice_pullup p_606(n779_v, n779_i1);
  spice_pullup p_564(n20_v, n20_i1);
  spice_pullup p_607(ONEBYTE_v, ONEBYTE_i1);
  spice_pullup p_115(n1507_v, n1507_i1);
  spice_pullup p_604(n773_v, n773_i0);
  spice_pullup p_602(n771_v, n771_i2);
  spice_pullup p_603(n770_v, n770_i2);
  spice_pullup p_600(n774_v, n774_i2);
  spice_pullup p_601(op_T5_jsr_v, op_T5_jsr_i1);
  spice_pullup p_874(irline3_v, irline3_i1);
  spice_pullup p_897(op_T0_adc_sbc_v, op_T0_adc_sbc_i0);
  spice_pullup p_896(n570_v, n570_i0);
  spice_pullup p_895(n571_v, n571_i1);
  spice_pullup p_894(n572_v, n572_i1);
  spice_pullup p_893(n578_v, n578_i3);
  spice_pullup p_892(op_T3_jsr_v, op_T3_jsr_i0);
  spice_pullup p_594(n880_v, n880_i1);
  spice_pullup p_595(n885_v, n885_i1);
  spice_pullup p_133(n696_v, n696_i1);
  spice_pullup p_22(n105_v, n105_i1);
  spice_pullup p_731(n1255_v, n1255_i2);
  spice_pullup p_572(n1085_v, n1085_i1);
  spice_pullup p_206(n428_v, n428_i1);
  spice_pullup p_134(n694_v, n694_i4);
  spice_pullup p_259(n523_v, n523_i0);
  spice_pullup p_258(op_ORS_v, op_ORS_i2);
  spice_pullup p_709(n1093_v, n1093_i2);
  spice_pullup p_708(n1091_v, n1091_i1);
  spice_pullup p_255(_C12_v, _C12_i1);
  spice_pullup p_257(n525_v, n525_i2);
  spice_pullup p_256(notir3_v, notir3_i2);
  spice_pullup p_251(n1392_v, n1392_i2);
  spice_pullup p_250(n1708_v, n1708_i2);
  spice_pullup p_253(n1129_v, n1129_i2);
  spice_pullup p_252(n1391_v, n1391_i1);
  spice_pullup p_419(n212_v, n212_i1);
  spice_pullup p_413(n1458_v, n1458_i4);
  spice_pullup p_411(n1107_v, n1107_i1);
  spice_pullup p_410(n1106_v, n1106_i1);
  spice_pullup p_417(DA_AB2_v, DA_AB2_i1);
  spice_pullup p_414(__AxB_6_v, __AxB_6_i2);
  spice_pullup p_345(n201_v, n201_i1);
  spice_pullup p_576(n976_v, n976_i4);
  spice_pullup p_677(alu1_v, alu1_i4);
  spice_pullup p_675(n877_v, n877_i0);
  spice_pullup p_101(n241_v, n241_i3);
  spice_pullup p_672(AxB7_v, AxB7_i1);
  spice_pullup p_671(n1560_v, n1560_i1);
  spice_pullup p_679(idl1_v, idl1_i2);
  spice_pullup p_100(op_ror_v, op_ror_i1);
  spice_pullup p_555(n499_v, n499_i1);
  spice_pullup p_883(n127_v, n127_i2);
  spice_pullup p_552(n1497_v, n1497_i2);
  spice_pullup p_440(n1039_v, n1039_i1);
  spice_pullup p_418(n_0_ADL0_v, n_0_ADL0_i2);
  spice_pullup p_105(n249_v, n249_i2);
  spice_pullup p_725(ir7_v, ir7_i3);
  spice_pullup p_795(x_op_T0_txa_v, x_op_T0_txa_i0);
  spice_pullup p_441(n753_v, n753_i0);
  spice_pullup p_979(n1187_v, n1187_i2);
  spice_pullup p_104(n242_v, n242_i3);
  spice_pullup p_204(n531_v, n531_i3);
  spice_pullup p_416(n1722_v, n1722_i4);
  spice_pullup p_415(n1109_v, n1109_i0);
  spice_pullup p_107(abl7_v, abl7_i4);
  spice_pullup p_443(n757_v, n757_i0);
  spice_pullup p_742(op_T0_bit_v, op_T0_bit_i0);
  spice_pullup p_106(op_T0_txa_v, op_T0_txa_i0);
  spice_pullup p_880(n123_v, n123_i1);
  spice_pullup p_881(pchp3_v, pchp3_i2);
  spice_pullup p_884(n128_v, n128_i2);
  spice_pullup p_885(n1647_v, n1647_i4);
  spice_pullup p_886(op_T__bit_v, op_T__bit_i1);
  spice_pullup p_887(n1641_v, n1641_i1);
  spice_pullup p_445(n754_v, n754_i1);
  spice_pullup p_317(_VEC_v, _VEC_i1);
  spice_pullup p_288(op_T2_php_pha_v, op_T2_php_pha_i0);
  spice_pullup p_282(C45_v, C45_i1);
  spice_pullup p_318(n1277_v, n1277_i3);
  spice_pullup p_568(n29_v, n29_i1);
  spice_pullup p_674(n876_v, n876_i1);
  spice_pullup p_673(n1240_v, n1240_i2);
  spice_pullup p_975(n564_v, n564_i3);
  spice_pullup p_711(op_T3_abs_idx_ind_v, op_T3_abs_idx_ind_i0);
  spice_pullup p_566(__AxBxC_2_v, __AxBxC_2_i1);
  spice_pullup p_719(dor6_v, dor6_i2);
  spice_pullup p_248(dpc34_PCLC_v, dpc34_PCLC_i1);
  spice_pullup p_249(n1705_v, n1705_i1);
  spice_pullup p_240(n1523_v, n1523_i3);
  spice_pullup p_869(n329_v, n329_i2);
  spice_pullup p_284(n141_v, n141_i4);
  spice_pullup p_400(C56_v, C56_i1);
  spice_pullup p_401(n1213_v, n1213_i0);
  spice_pullup p_402(n632_v, n632_i1);
  spice_pullup p_403(alu0_v, alu0_i3);
  spice_pullup p_860(__AxBxC_4_v, __AxBxC_4_i1);
  spice_pullup p_179(n678_v, n678_i2);
  spice_pullup p_861(n658_v, n658_i3);
  spice_pullup p_176(n160_v, n160_i1);
  spice_pullup p_177(n161_v, n161_i2);
  spice_pullup p_227(clock2_v, clock2_i1);
  spice_pullup p_668(n961_v, n961_i2);
  spice_pullup p_561(n25_v, n25_i1);
  spice_pullup p_717(n1413_v, n1413_i2);
  spice_pullup p_560(op_T4_ind_y_v, op_T4_ind_y_i0);
  spice_pullup p_175(op_T0_tax_v, op_T0_tax_i0);
  spice_pullup p_556(n494_v, n494_i1);
  spice_pullup p_38(n553_v, n553_i0);
  spice_pullup p_39(op_T0_php_pha_v, op_T0_php_pha_i0);
  spice_pullup p_36(n551_v, n551_i2);
  spice_pullup p_37(n550_v, n550_i0);
  spice_pullup p_35(n556_v, n556_i2);
  spice_pullup p_32(n1629_v, n1629_i0);
  spice_pullup p_33(aluanandb0_v, aluanandb0_i1);
  spice_pullup p_30(n1621_v, n1621_i2);
  spice_pullup p_31(ir1_v, ir1_i2);
  spice_pullup p_1017(n1369_v, n1369_i3);
  spice_pullup p_457(aluaorb1_v, aluaorb1_i1);
  spice_pullup p_456(op_T3_stack_bit_jmp_v, op_T3_stack_bit_jmp_i0);
  spice_pullup p_879(n122_v, n122_i1);
  spice_pullup p_878(op_T3_v, op_T3_i1);
  spice_pullup p_454(n1025_v, n1025_i2);
  spice_pullup p_178(n163_v, n163_i1);
  spice_pullup p_553(notaluvout_v, notaluvout_i1);
  spice_pullup p_550(n1301_v, n1301_i4);
  spice_pullup p_728(n1531_v, n1531_i3);
  spice_pullup p_989(n721_v, n721_i4);
  spice_pullup p_988(n720_v, n720_i1);
  spice_pullup p_981(short_circuit_idx_add_v, short_circuit_idx_add_i0);
  spice_pullup p_551(n1303_v, n1303_i0);
  spice_pullup p_982(notir2_v, notir2_i2);
  spice_pullup p_985(n726_v, n726_i1);
  spice_pullup p_987(n723_v, n723_i4);
  spice_pullup p_986(dpc22__DSA_v, dpc22__DSA_i2);
  spice_pullup p_720(n1416_v, n1416_i1);
  spice_pullup p_451(n507_v, n507_i1);
  spice_pullup p_723(_C78_v, _C78_i1);
  spice_pullup p_48(op_SUMS_v, op_SUMS_i1);
  spice_pullup p_336(op_ANDS_v, op_ANDS_i2);
  spice_pullup p_191(n608_v, n608_i2);
  spice_pullup p_557(n496_v, n496_i2);
  spice_pullup p_337(n1286_v, n1286_i0);
  spice_pullup p_889(n1643_v, n1643_i1);
  spice_pullup p_442(op_T2_php_v, op_T2_php_i0);
  spice_pullup p_447(n506_v, n506_i1);
  spice_pullup p_639(op_rol_ror_v, op_rol_ror_i0);
  spice_pullup p_996(n472_v, n472_i1);
  spice_pullup p_706(n1097_v, n1097_i0);
  spice_pullup p_471(n1206_v, n1206_i4);
  spice_pullup p_470(op_T2_ind_y_v, op_T2_ind_y_i0);
  spice_pullup p_475(n1211_v, n1211_i2);
  spice_pullup p_474(n1202_v, n1202_i1);
  spice_pullup p_477(n1214_v, n1214_i1);
  spice_pullup p_476(__AxB7__C67_v, __AxB7__C67_i0);
  spice_pullup p_297(op_T__adc_sbc_v, op_T__adc_sbc_i0);
  spice_pullup p_167(n253_v, n253_i1);
  spice_pullup p_697(n1073_v, n1073_i1);
  spice_pullup p_696(n1075_v, n1075_i2);
  spice_pullup p_691(op_jmp_v, op_jmp_i0);
  spice_pullup p_690(n767_v, n767_i3);
  spice_pullup p_693(pclp2_v, pclp2_i2);
  spice_pullup p_692(alu7_v, alu7_i3);
  spice_pullup p_505(n192_v, n192_i0);
  spice_pullup p_504(_AxB_2__C12_v, _AxB_2__C12_i0);
  spice_pullup p_507(n1457_v, n1457_i0);
  spice_pullup p_506(n1455_v, n1455_i2);
  spice_pullup p_501(notir0_v, notir0_i2);
  spice_pullup p_500(n198_v, n198_i3);
  spice_pullup p_702(pd2_clearIR_v, pd2_clearIR_i1);
  spice_pullup p_185(pd1_clearIR_v, pd1_clearIR_i1);
  spice_pullup p_189(n807_v, n807_i0);
  spice_pullup p_701(n1677_v, n1677_i3);
  spice_pullup p_508(dor5_v, dor5_i2);
  spice_pullup p_29(pd0_clearIR_v, pd0_clearIR_i1);
  spice_pullup p_28(op_T0_eor_v, op_T0_eor_i1);
  spice_pullup p_21(n104_v, n104_i1);
  spice_pullup p_23(op_T5_ind_x_v, op_T5_ind_x_i0);
  spice_pullup p_25(n90_v, n90_i3);
  spice_pullup p_24(n91_v, n91_i3);
  spice_pullup p_27(dor0_v, dor0_i2);
  spice_pullup p_816(n330_v, n330_i1);
  spice_pullup p_663(n1521_v, n1521_i2);
  spice_pullup p_815(alu6_v, alu6_i4);
  spice_pullup p_747(n476_v, n476_i2);
  spice_pullup p_811(n335_v, n335_i0);
  spice_pullup p_810(n649_v, n649_i2);
  spice_pullup p_539(n616_v, n616_i1);
  spice_pullup p_383(dor7_v, dor7_i2);
  spice_pullup p_868(ir0_v, ir0_i2);
  spice_pullup p_382(n62_v, n62_i2);
  spice_pullup p_567(n23_v, n23_i1);
  spice_pullup p_864(n321_v, n321_i3);
  spice_pullup p_380(op_T3_ind_y_v, op_T3_ind_y_i0);
  spice_pullup p_387(n1588_v, n1588_i2);
  spice_pullup p_386(n1371_v, n1371_i0);
  spice_pullup p_605(n772_v, n772_i3);
  spice_pullup p_385(Reset0_v, Reset0_i3);
  spice_pullup p_384(_AxB_4__C34_v, _AxB_4__C34_i0);
  spice_pullup p_437(n849_v, n849_i2);
  spice_pullup p_388(op_T4_jmp_v, op_T4_jmp_i0);
  spice_pullup p_998(x_op_T4_rti_v, x_op_T4_rti_i0);
  spice_pullup p_999(op_T0_cli_sei_v, op_T0_cli_sei_i1);
  spice_pullup p_433(n844_v, n844_i1);
  spice_pullup p_34(_AxB_0__C0in_v, _AxB_0__C0in_i0);
  spice_pullup p_992(notalucin_v, notalucin_i2);
  spice_pullup p_993(n1166_v, n1166_i1);
  spice_pullup p_990(n728_v, n728_i2);
  spice_pullup p_991(op_clv_v, op_clv_i1);
  spice_pullup p_997(n46_v, n46_i0);
  spice_pullup p_994(op_T5_ind_y_v, op_T5_ind_y_i0);
  spice_pullup p_995(n1169_v, n1169_i3);
  spice_pullup p_735(n1258_v, n1258_i1);
  spice_pullup p_462(n501_v, n501_i1);
  spice_pullup p_463(n604_v, n604_i1);
  spice_pullup p_460(n1037_v, n1037_i1);
  spice_pullup p_461(n1034_v, n1034_i3);
  spice_pullup p_466(n600_v, n600_i1);
  spice_pullup p_464(op_T3_mem_abs_v, op_T3_mem_abs_i0);
  spice_pullup p_465(alu4_v, alu4_i3);
  spice_pullup p_468(n602_v, n602_i1);
  spice_pullup p_381(n61_v, n61_i1);
  spice_pullup p_264(n1230_v, n1230_i2);
  spice_pullup p_265(n1231_v, n1231_i2);
  spice_pullup p_266(abl4_v, abl4_i4);
  spice_pullup p_267(op_T0_cpy_iny_v, op_T0_cpy_iny_i0);
  spice_pullup p_261(n1017_v, n1017_i2);
  spice_pullup p_262(xx_op_T5_jsr_v, xx_op_T5_jsr_i0);
  spice_pullup p_263(A_B5_v, A_B5_i1);
  spice_pullup p_155(n366_v, n366_i1);
  spice_pullup p_268(n1238_v, n1238_i2);
  spice_pullup p_269(op_T2_branch_v, op_T2_branch_i1);
  spice_pullup p_358(n920_v, n920_i2);
  spice_pullup p_688(n763_v, n763_i1);
  spice_pullup p_689(n761_v, n761_i2);
  spice_pullup p_684(n896_v, n896_i2);
  spice_pullup p_516(op_rti_rts_v, op_rti_rts_i1);
  spice_pullup p_517(n850_v, n850_i2);
  spice_pullup p_512(n905_v, n905_i1);
  spice_pullup p_513(n1511_v, n1511_i1);
  spice_pullup p_510(n906_v, n906_i3);
  spice_pullup p_511(op_T3_mem_zp_idx_v, op_T3_mem_zp_idx_i0);
  spice_pullup p_156(PD_0xx0xx0x_v, PD_0xx0xx0x_i1);
  spice_pullup p_157(op_T0_iny_dey_v, op_T0_iny_dey_i0);
  spice_pullup p_154(n368_v, n368_i1);
  spice_pullup p_198(op_T3_abs_idx_v, op_T3_abs_idx_i0);
  spice_pullup p_473(DBNeg_v, DBNeg_i1);
  spice_pullup p_150(n1380_v, n1380_i2);
  spice_pullup p_151(op_T3_jmp_v, op_T3_jmp_i1);
  spice_pullup p_651(n1010_v, n1010_i2);
  spice_pullup p_650(n1318_v, n1318_i3);
  spice_pullup p_964(pchp1_v, pchp1_i2);
  spice_pullup p_472(n609_v, n609_i0);
  spice_pullup p_655(n311_v, n311_i1);
  spice_pullup p_657(alu5_v, alu5_i4);
  spice_pullup p_656(n317_v, n317_i2);
  spice_pullup p_582(n182_v, n182_i2);
  spice_pullup p_523(DBZ_v, DBZ_i1);
  spice_pullup p_859(n652_v, n652_i4);
  spice_pullup p_858(n457_v, n457_i2);
  spice_pullup p_853(n419_v, n419_i2);
  spice_pullup p_852(x_op_T3_plp_pla_v, x_op_T3_plp_pla_i0);
  spice_pullup p_851(n1433_v, n1433_i0);
  spice_pullup p_850(n1434_v, n1434_i2);
  spice_pullup p_857(n1345_v, n1345_i0);
  spice_pullup p_856(n1344_v, n1344_i4);
  spice_pullup p_855(n453_v, n453_i1);
  spice_pullup p_854(dasb2_v, dasb2_i1);
  spice_pullup p_479(n1111_v, n1111_i0);
  spice_pullup p_716(n1412_v, n1412_i1);
  spice_pullup p_862(DA_AxB2_v, DA_AxB2_i0);
  spice_pullup p_478(n1215_v, n1215_i2);
  spice_pullup p_962(n111_v, n111_i2);
  spice_pullup p_534(n1694_v, n1694_i3);
  spice_pullup p_455(n1024_v, n1024_i2);
  spice_pullup p_803(n35_v, n35_i2);
  spice_pullup p_531(n1056_v, n1056_i1);
  spice_pullup p_467(n603_v, n603_i1);
  spice_pullup p_469(n1205_v, n1205_i0);
  spice_pullup p_329(n620_v, n620_i0);
  spice_pullup p_328(n1225_v, n1225_i3);
  spice_pullup p_459(n1028_v, n1028_i2);
  spice_pullup p_458(C23_v, C23_i1);
  spice_pullup p_325(n1002_v, n1002_i1);
  spice_pullup p_324(n515_v, n515_i1);
  spice_pullup p_327(DA_C01_v, DA_C01_i0);
  spice_pullup p_326(op_store_v, op_store_i1);
  spice_pullup p_321(dasb1_v, dasb1_i1);
  spice_pullup p_320(n518_v, n518_i3);
  spice_pullup p_323(op_implied_v, op_implied_i1);
  spice_pullup p_322(n1007_v, n1007_i1);
  spice_pullup p_299(VEC1_v, VEC1_i2);
  spice_pullup p_298(op_T__iny_dey_v, op_T__iny_dey_i0);
  spice_pullup p_729(n1256_v, n1256_i2);
  spice_pullup p_62(n1578_v, n1578_i1);
  spice_pullup p_749(n958_v, n958_i3);
  spice_pullup p_215(n853_v, n853_i1);
  spice_pullup p_214(_C56_v, _C56_i1);
  spice_pullup p_219(n225_v, n225_i1);
  spice_pullup p_217(n228_v, n228_i1);
  spice_pullup p_332(n624_v, n624_i2);
  spice_pullup p_743(n306_v, n306_i2);
  spice_pullup p_529(n1054_v, n1054_i1);
  spice_pullup p_528(x_op_jmp_v, x_op_jmp_i0);
  spice_pullup p_522(n743_v, n743_i0);
  spice_pullup p_521(n6_v, n6_i2);
  spice_pullup p_520(n819_v, n819_i0);
  spice_pullup p_524(dor1_v, dor1_i2);
  spice_pullup p_740(op_T__cmp_v, op_T__cmp_i0);
  spice_pullup p_295(n824_v, n824_i2);
  spice_pullup p_294(op_SRS_v, op_SRS_i4);
  spice_pullup p_744(n307_v, n307_i0);
  spice_pullup p_145(n1389_v, n1389_i4);
  spice_pullup p_144(n410_v, n410_i0);
  spice_pullup p_147(ir2_v, ir2_i2);
  spice_pullup p_146(notalucout_v, notalucout_i1);
  spice_pullup p_141(op_shift_v, op_shift_i0);
  spice_pullup p_140(pd4_clearIR_v, pd4_clearIR_i1);
  spice_pullup p_143(n548_v, n548_i2);
  spice_pullup p_142(n544_v, n544_i1);
  spice_pullup p_149(n1386_v, n1386_i0);
  spice_pullup p_148(op_T5_mem_ind_idx_v, op_T5_mem_ind_idx_i0);
  spice_pullup p_926(op_T4_abs_idx_v, op_T4_abs_idx_i0);
  spice_pullup p_20(n109_v, n109_i2);
  spice_pullup p_406(n638_v, n638_i1);
  spice_pullup p_685(n646_v, n646_i2);
  spice_pullup p_274(n238_v, n238_i1);
  spice_pullup p_407(n1218_v, n1218_i1);
  spice_pullup p_754(n954_v, n954_i1);
  spice_pullup p_924(n1275_v, n1275_i1);
  spice_pullup p_1009(n1716_v, n1716_i0);
  spice_pullup p_359(n923_v, n923_i1);
  spice_pullup p_260(n1016_v, n1016_i1);
  spice_pullup p_349(n206_v, n206_i3);
  spice_pullup p_844(n1655_v, n1655_i1);
  spice_pullup p_845(n586_v, n586_i1);
  spice_pullup p_846(n587_v, n587_i1);
  spice_pullup p_847(n582_v, n582_i3);
  spice_pullup p_573(n1084_v, n1084_i2);
  spice_pullup p_831(n708_v, n708_i1);
  spice_pullup p_830(n139_v, n139_i1);
  spice_pullup p_343(n19_v, n19_i1);
  spice_pullup p_354(ir3_v, ir3_i2);
  spice_pullup p_835(notir1_v, notir1_i2);
  spice_pullup p_834(__AxB_2_v, __AxB_2_i1);
  spice_pullup p_920(n1519_v, n1519_i1);
  spice_pullup p_686(n769_v, n769_i1);
  spice_pullup p_687(n762_v, n762_i1);
  spice_pullup p_682(n1244_v, n1244_i1);
  spice_pullup p_683(n890_v, n890_i2);
  spice_pullup p_680(n871_v, n871_i3);
  spice_pullup p_817(DC78_v, DC78_i1);
  spice_pullup p_518(_TWOCYCLE_v, _TWOCYCLE_i1);
  spice_pullup p_755(n956_v, n956_i1);
  spice_pullup p_519(n852_v, n852_i1);
  spice_pullup p_409(n465_v, n465_i2);
  spice_pullup p_814(n336_v, n336_i3);
  spice_pullup p_26(n93_v, n93_i2);
  spice_pullup p_448(idl0_v, idl0_i2);
  spice_pullup p_449(n1596_v, n1596_i3);
  spice_pullup p_712(n1099_v, n1099_i1);
  spice_pullup p_338(n11_v, n11_i1);
  spice_pullup p_339(n10_v, n10_i0);
  spice_pullup p_334(n628_v, n628_i2);
  spice_pullup p_331(n625_v, n625_i2);
  spice_pullup p_193(x_op_T__adc_sbc_v, x_op_T__adc_sbc_i1);
  spice_pullup p_190(op_T4_brk_jsr_v, op_T4_brk_jsr_i0);
  spice_pullup p_208(n1398_v, n1398_i2);
  spice_pullup p_209(n420_v, n420_i2);
  spice_pullup p_490(n466_v, n466_i1);
  spice_pullup p_535(n1691_v, n1691_i2);
  spice_pullup p_536(n618_v, n618_i4);
  spice_pullup p_537(n613_v, n613_i0);
  spice_pullup p_530(n1055_v, n1055_i0);
  spice_pullup p_194(n1154_v, n1154_i0);
  spice_pullup p_532(op_T2_abs_v, op_T2_abs_i0);
  spice_pullup p_195(n1157_v, n1157_i2);
  spice_pullup p_538(n611_v, n611_i2);
  spice_pullup p_980(n1184_v, n1184_i0);
  spice_pullup p_199(op_brk_rti_v, op_brk_rti_i0);
  spice_pullup p_1014(n478_v, n478_i2);
  spice_pullup p_704(n1094_v, n1094_i1);
  spice_pullup p_152(brk_done_v, brk_done_i1);
  spice_pullup p_158(n383_v, n383_i1);
  spice_pullup p_159(n384_v, n384_i1);
  spice_pullup p_1016(n1368_v, n1368_i1);
  spice_pullup p_404(n636_v, n636_i2);
  spice_pullup p_98(notir6_v, notir6_i2);
  spice_pullup p_99(op_T0_txs_v, op_T0_txs_i0);
  spice_pullup p_90(n372_v, n372_i1);
  spice_pullup p_91(n374_v, n374_i2);
  spice_pullup p_92(abl1_v, abl1_i4);
  spice_pullup p_93(n392_v, n392_i1);
  spice_pullup p_94(idl7_v, idl7_i2);
  spice_pullup p_95(n390_v, n390_i2);
  spice_pullup p_96(n397_v, n397_i1);
  spice_pullup p_97(n396_v, n396_i2);
  spice_pullup p_758(n718_v, n718_i2);
  spice_pullup p_633(n664_v, n664_i2);
  spice_pullup p_632(op_T0_ldy_mem_v, op_T0_ldy_mem_i0);
  spice_pullup p_983(n1180_v, n1180_i1);
  spice_pullup p_631(n1262_v, n1262_i1);
  spice_pullup p_759(n717_v, n717_i1);
  spice_pullup p_630(pd5_clearIR_v, pd5_clearIR_i1);
  spice_pullup p_637(VEC0_v, VEC0_i2);
  spice_pullup p_718(alu3_v, alu3_i3);
  spice_pullup p_635(n1265_v, n1265_i2);
  spice_pullup p_833(n700_v, n700_i2);
  spice_pullup p_832(n709_v, n709_i2);
  spice_pullup p_837(n83_v, n83_i1);
  spice_pullup p_836(rdy_v, rdy_i1);
  spice_pullup p_714(op_T0_cld_sed_v, op_T0_cld_sed_i1);
  spice_pullup p_246(n1499_v, n1499_i3);
  spice_pullup p_247(notir5_v, notir5_i3);
  spice_pullup p_244(n1496_v, n1496_i4);
  spice_pullup p_203(__AxBxC_7_v, __AxBxC_7_i1);
  spice_pullup p_245(op_T0_shift_a_v, op_T0_shift_a_i0);
  spice_pullup p_242(dasb7_v, dasb7_i1);
  spice_pullup p_243(n1495_v, n1495_i1);
  spice_pullup p_241(n1492_v, n1492_i1);
  spice_pullup p_654(n312_v, n312_i2);
  spice_pullup p_949(n264_v, n264_i2);
  spice_pullup p_948(n267_v, n267_i0);
  spice_pullup p_945(n262_v, n262_i1);
  spice_pullup p_944(dasb5_v, dasb5_i1);
  spice_pullup p_947(n260_v, n260_i0);
  spice_pullup p_946(n261_v, n261_i1);
  spice_pullup p_941(op_T0_tay_ldy_not_idx_v, op_T0_tay_ldy_not_idx_i0);
  spice_pullup p_940(abh2_v, abh2_i4);
  spice_pullup p_943(idl6_v, idl6_i2);
  spice_pullup p_942(n1441_v, n1441_i2);
  spice_pullup p_968(n1632_v, n1632_i2);

  spice_node_2 n_DBNeg(eclk, ereset, DBNeg_i0,DBNeg_i1, DBNeg_v);
  spice_node_2 n_n344(eclk, ereset, n344_i0,n344_i2, n344_v);
  spice_node_2 n_n345(eclk, ereset, n345_i0,n345_i3, n345_v);
  spice_node_2 n_n347(eclk, ereset, n347_i0,n347_i3, n347_v);
  spice_node_3 n_n340(eclk, ereset, n340_i0,n340_i1,n340_i2, n340_v);
  spice_node_2 n_op_T4(eclk, ereset, op_T4_i0,op_T4_i1, op_T4_v);
  spice_node_2 n_x_op_T3_ind_y(eclk, ereset, x_op_T3_ind_y_i0,x_op_T3_ind_y_i2, x_op_T3_ind_y_v);
  spice_node_1 n_p3(eclk, ereset, p3_i0, p3_v);
  spice_node_3 n_ab13(eclk, ereset, ab13_i0,ab13_i1,ab13_i2, ab13_v);
  spice_node_2 n_n298(eclk, ereset, n298_i1,n298_i2, n298_v);
  spice_node_3 n_n299(eclk, ereset, n299_i0,n299_i1,n299_i2, n299_v);
  spice_node_6 n_n296(eclk, ereset, n296_i0,n296_i1,n296_i2,n296_i3,n296_i4,n296_i5, n296_v);
  spice_node_2 n_n297(eclk, ereset, n297_i0,n297_i1, n297_v);
  spice_node_1 n_pipeUNK20(eclk, ereset, pipeUNK20_i0, pipeUNK20_v);
  spice_node_2 n___AxB1__C01(eclk, ereset, __AxB1__C01_i0,__AxB1__C01_i1, __AxB1__C01_v);
  spice_node_2 n_pch1(eclk, ereset, pch1_i1,pch1_i2, pch1_v);
  spice_node_2 n_n293(eclk, ereset, n293_i0,n293_i3, n293_v);
  spice_node_1 n_n597(eclk, ereset, n597_i0, n597_v);
  spice_node_2 n_n291(eclk, ereset, n291_i2,n291_i3, n291_v);
  spice_node_2 n_n270(eclk, ereset, n270_i0,n270_i1, n270_v);
  spice_node_2 n_op_T0_jsr(eclk, ereset, op_T0_jsr_i0,op_T0_jsr_i1, op_T0_jsr_v);
  spice_node_3 n_n272(eclk, ereset, n272_i0,n272_i2,n272_i3, n272_v);
  spice_node_2 n_op_T2_abs_access(eclk, ereset, op_T2_abs_access_i0,op_T2_abs_access_i2, op_T2_abs_access_v);
  spice_node_3 n___AxBxC_3(eclk, ereset, __AxBxC_3_i0,__AxBxC_3_i1,__AxBxC_3_i2, __AxBxC_3_v);
  spice_node_2 n_n275(eclk, ereset, n275_i0,n275_i2, n275_v);
  spice_node_1 n_notalu2(eclk, ereset, notalu2_i1, notalu2_v);
  spice_node_6 n_n277(eclk, ereset, n277_i0,n277_i1,n277_i2,n277_i3,n277_i4,n277_i5, n277_v);
  spice_node_2 n_n278(eclk, ereset, n278_i0,n278_i2, n278_v);
  spice_node_2 n_n279(eclk, ereset, n279_i0,n279_i1, n279_v);
  spice_node_2 n_n108(eclk, ereset, n108_i1,n108_i2, n108_v);
  spice_node_3 n_n109(eclk, ereset, n109_i0,n109_i1,n109_i2, n109_v);
  spice_node_2 n_n102(eclk, ereset, n102_i0,n102_i2, n102_v);
  spice_node_1 n_irq(eclk, ereset, irq_i1, irq_v);
  spice_node_1 n_n101(eclk, ereset, n101_i0, n101_v);
  spice_node_2 n__ABL1(eclk, ereset, _ABL1_i1,_ABL1_i2, _ABL1_v);
  spice_node_3 n_n104(eclk, ereset, n104_i0,n104_i1,n104_i2, n104_v);
  spice_node_2 n_n105(eclk, ereset, n105_i0,n105_i1, n105_v);
  spice_node_1 n_pipeUNK04(eclk, ereset, pipeUNK04_i0, pipeUNK04_v);
  spice_node_2 n_x1(eclk, ereset, x1_i0,x1_i1, x1_v);
  spice_node_2 n_n91(eclk, ereset, n91_i0,n91_i3, n91_v);
  spice_node_3 n_n90(eclk, ereset, n90_i0,n90_i2,n90_i3, n90_v);
  spice_node_3 n_n93(eclk, ereset, n93_i0,n93_i1,n93_i2, n93_v);
  spice_node_2 n__ABH3(eclk, ereset, _ABH3_i0,_ABH3_i2, _ABH3_v);
  spice_node_1 n_n95(eclk, ereset, n95_i0, n95_v);
  spice_node_1 n_n94(eclk, ereset, n94_i1, n94_v);
  spice_node_2 n_dor0(eclk, ereset, dor0_i0,dor0_i2, dor0_v);
  spice_node_3 n_alub3(eclk, ereset, alub3_i0,alub3_i1,alub3_i2, alub3_v);
  spice_node_2 n_op_T0_eor(eclk, ereset, op_T0_eor_i1,op_T0_eor_i2, op_T0_eor_v);
  spice_node_2 n_pd0_clearIR(eclk, ereset, pd0_clearIR_i1,pd0_clearIR_i2, pd0_clearIR_v);
  spice_node_3 n_n1621(eclk, ereset, n1621_i0,n1621_i1,n1621_i2, n1621_v);
  spice_node_2 n_n1620(eclk, ereset, n1620_i0,n1620_i2, n1620_v);
  spice_node_2 n_alua6(eclk, ereset, alua6_i0,alua6_i1, alua6_v);
  spice_node_2 n_ir1(eclk, ereset, ir1_i1,ir1_i2, ir1_v);
  spice_node_1 n_n1625(eclk, ereset, n1625_i0, n1625_v);
  spice_node_1 n_n1624(eclk, ereset, n1624_i0, n1624_v);
  spice_node_2 n_n1629(eclk, ereset, n1629_i0,n1629_i1, n1629_v);
  spice_node_3 n_aluanandb0(eclk, ereset, aluanandb0_i0,aluanandb0_i1,aluanandb0_i3, aluanandb0_v);
  spice_node_1 n_n559(eclk, ereset, n559_i0, n559_v);
  spice_node_2 n__AxB_0__C0in(eclk, ereset, _AxB_0__C0in_i0,_AxB_0__C0in_i1, _AxB_0__C0in_v);
  spice_node_1 n_pipe_T0(eclk, ereset, pipe_T0_i0, pipe_T0_v);
  spice_node_2 n_n556(eclk, ereset, n556_i0,n556_i2, n556_v);
  spice_node_2 n_n551(eclk, ereset, n551_i1,n551_i2, n551_v);
  spice_node_2 n_n550(eclk, ereset, n550_i0,n550_i2, n550_v);
  spice_node_2 n_n553(eclk, ereset, n553_i0,n553_i1, n553_v);
  spice_node_2 n_op_T0_php_pha(eclk, ereset, op_T0_php_pha_i0,op_T0_php_pha_i1, op_T0_php_pha_v);
  spice_node_3 n_n1199(eclk, ereset, n1199_i0,n1199_i1,n1199_i2, n1199_v);
  spice_node_2 n_n1191(eclk, ereset, n1191_i0,n1191_i2, n1191_v);
  spice_node_3 n_n1190(eclk, ereset, n1190_i0,n1190_i1,n1190_i2, n1190_v);
  spice_node_2 n_n_0_ADL2(eclk, ereset, n_0_ADL2_i0,n_0_ADL2_i2, n_0_ADL2_v);
  spice_node_3 n_n1192(eclk, ereset, n1192_i0,n1192_i1,n1192_i2, n1192_v);
  spice_node_2 n_n1195(eclk, ereset, n1195_i2,n1195_i3, n1195_v);
  spice_node_3 n_n1194(eclk, ereset, n1194_i1,n1194_i2,n1194_i3, n1194_v);
  spice_node_3 n___AxBxC_6(eclk, ereset, __AxBxC_6_i0,__AxBxC_6_i1,__AxBxC_6_i2, __AxBxC_6_v);
  spice_node_3 n_op_SUMS(eclk, ereset, op_SUMS_i0,op_SUMS_i1,op_SUMS_i2, op_SUMS_v);
  spice_node_1 n_n1177(eclk, ereset, n1177_i0, n1177_v);
  spice_node_1 n_pipeUNK21(eclk, ereset, pipeUNK21_i1, pipeUNK21_v);
  spice_node_3 n_n1175(eclk, ereset, n1175_i0,n1175_i1,n1175_i2, n1175_v);
  spice_node_2 n__op_branch_bit7(eclk, ereset, _op_branch_bit7_i0,_op_branch_bit7_i2, _op_branch_bit7_v);
  spice_node_2 n_x_op_T0_tya(eclk, ereset, x_op_T0_tya_i0,x_op_T0_tya_i1, x_op_T0_tya_v);
  spice_node_1 n_clk0(eclk, ereset, clk0_i2, clk0_v);
  spice_node_2 n_n1170(eclk, ereset, n1170_i0,n1170_i1, n1170_v);
  spice_node_3 n_n1179(eclk, ereset, n1179_i0,n1179_i1,n1179_i2, n1179_v);
  spice_node_3 n_n1178(eclk, ereset, n1178_i0,n1178_i1,n1178_i2, n1178_v);
  spice_node_2 n_n510(eclk, ereset, n510_i0,n510_i2, n510_v);
  spice_node_3 n_n513(eclk, ereset, n513_i0,n513_i1,n513_i2, n513_v);
  spice_node_2 n_C01(eclk, ereset, C01_i1,C01_i2, C01_v);
  spice_node_1 n_notidl3(eclk, ereset, notidl3_i0, notidl3_v);
  spice_node_12 n_sb2(eclk, ereset, sb2_i0,sb2_i1,sb2_i2,sb2_i3,sb2_i4,sb2_i6,sb2_i7,sb2_i8,sb2_i9,sb2_i10,sb2_i11,sb2_i12, sb2_v);
  spice_node_1 n_n512(eclk, ereset, n512_i1, n512_v);
  spice_node_3 n_n1281(eclk, ereset, n1281_i0,n1281_i1,n1281_i2, n1281_v);
  spice_node_1 n_pipeUNK12(eclk, ereset, pipeUNK12_i0, pipeUNK12_v);
  spice_node_8 n_adl1(eclk, ereset, adl1_i0,adl1_i1,adl1_i2,adl1_i3,adl1_i4,adl1_i5,adl1_i7,adl1_i8, adl1_v);
  spice_node_3 n_n515(eclk, ereset, n515_i0,n515_i1,n515_i2, n515_v);
  spice_node_2 n_fetch(eclk, ereset, fetch_i0,fetch_i1, fetch_v);
  spice_node_2 n_n1289(eclk, ereset, n1289_i0,n1289_i1, n1289_v);
  spice_node_1 n_notdor2(eclk, ereset, notdor2_i1, notdor2_v);
  spice_node_1 n_n1579(eclk, ereset, n1579_i1, n1579_v);
  spice_node_2 n_n1578(eclk, ereset, n1578_i0,n1578_i1, n1578_v);
  spice_node_2 n_n689(eclk, ereset, n689_i0,n689_i1, n689_v);
  spice_node_12 n_sb7(eclk, ereset, sb7_i0,sb7_i1,sb7_i2,sb7_i3,sb7_i4,sb7_i5,sb7_i6,sb7_i7,sb7_i8,sb7_i9,sb7_i10,sb7_i11, sb7_v);
  spice_node_1 n_pipeUNK28(eclk, ereset, pipeUNK28_i0, pipeUNK28_v);
  spice_node_3 n_Pout0(eclk, ereset, Pout0_i0,Pout0_i1,Pout0_i2, Pout0_v);
  spice_node_1 n_n1570(eclk, ereset, n1570_i0, n1570_v);
  spice_node_4 n_n681(eclk, ereset, n681_i0,n681_i1,n681_i3,n681_i5, n681_v);
  spice_node_2 n_ir3(eclk, ereset, ir3_i1,ir3_i2, ir3_v);
  spice_node_3 n_n1575(eclk, ereset, n1575_i1,n1575_i2,n1575_i3, n1575_v);
  spice_node_2 n_op_T0_tsx(eclk, ereset, op_T0_tsx_i1,op_T0_tsx_i2, op_T0_tsx_v);
  spice_node_3 n_n458(eclk, ereset, n458_i0,n458_i1,n458_i2, n458_v);
  spice_node_2 n_pcl5(eclk, ereset, pcl5_i1,pcl5_i2, pcl5_v);
  spice_node_1 n_n621(eclk, ereset, n621_i1, n621_v);
  spice_node_1 n_notdor4(eclk, ereset, notdor4_i0, notdor4_v);
  spice_node_2 n_n1224(eclk, ereset, n1224_i0,n1224_i1, n1224_v);
  spice_node_1 n_p1(eclk, ereset, p1_i1, p1_v);
  spice_node_2 n_n1222(eclk, ereset, n1222_i0,n1222_i1, n1222_v);
  spice_node_1 n_n1221(eclk, ereset, n1221_i1, n1221_v);
  spice_node_3 n_n624(eclk, ereset, n624_i0,n624_i1,n624_i2, n624_v);
  spice_node_2 n_n1371(eclk, ereset, n1371_i0,n1371_i2, n1371_v);
  spice_node_3 n_Pout7(eclk, ereset, Pout7_i0,Pout7_i1,Pout7_i2, Pout7_v);
  spice_node_3 n_n404(eclk, ereset, n404_i0,n404_i2,n404_i3, n404_v);
  spice_node_3 n_n1375(eclk, ereset, n1375_i0,n1375_i1,n1375_i2, n1375_v);
  spice_node_3 n_n1374(eclk, ereset, n1374_i0,n1374_i1,n1374_i2, n1374_v);
  spice_node_4 n_alu0(eclk, ereset, alu0_i0,alu0_i1,alu0_i2,alu0_i3, alu0_v);
  spice_node_3 n_ab1(eclk, ereset, ab1_i0,ab1_i1,ab1_i2, ab1_v);
  spice_node_3 n_n1379(eclk, ereset, n1379_i0,n1379_i1,n1379_i2, n1379_v);
  spice_node_3 n_n409(eclk, ereset, n409_i0,n409_i1,n409_i3, n409_v);
  spice_node_1 n_n408(eclk, ereset, n408_i0, n408_v);
  spice_node_2 n_n453(eclk, ereset, n453_i0,n453_i1, n453_v);
  spice_node_5 n_n1344(eclk, ereset, n1344_i0,n1344_i1,n1344_i2,n1344_i3,n1344_i4, n1344_v);
  spice_node_2 n_n1345(eclk, ereset, n1345_i0,n1345_i1, n1345_v);
  spice_node_2 n_n1346(eclk, ereset, n1346_i0,n1346_i3, n1346_v);
  spice_node_3 n_n1347(eclk, ereset, n1347_i0,n1347_i1,n1347_i2, n1347_v);
  spice_node_2 n_n1245(eclk, ereset, n1245_i0,n1245_i1, n1245_v);
  spice_node_2 n_dpc36_IPC(eclk, ereset, dpc36_IPC_i0,dpc36_IPC_i3, dpc36_IPC_v);
  spice_node_3 n_n378(eclk, ereset, n378_i1,n378_i2,n378_i3, n378_v);
  spice_node_3 n___AxBxC_0(eclk, ereset, __AxBxC_0_i0,__AxBxC_0_i1,__AxBxC_0_i2, __AxBxC_0_v);
  spice_node_2 n_op_T5_brk(eclk, ereset, op_T5_brk_i1,op_T5_brk_i2, op_T5_brk_v);
  spice_node_2 n_n373(eclk, ereset, n373_i0,n373_i2, n373_v);
  spice_node_2 n_n372(eclk, ereset, n372_i0,n372_i1, n372_v);
  spice_node_3 n_n374(eclk, ereset, n374_i0,n374_i1,n374_i2, n374_v);
  spice_node_2 n_pcl6(eclk, ereset, pcl6_i1,pcl6_i2, pcl6_v);
  spice_node_2 n_abl1(eclk, ereset, abl1_i3,abl1_i4, abl1_v);
  spice_node_1 n_n393(eclk, ereset, n393_i0, n393_v);
  spice_node_2 n_n392(eclk, ereset, n392_i0,n392_i1, n392_v);
  spice_node_3 n_idl7(eclk, ereset, idl7_i0,idl7_i1,idl7_i2, idl7_v);
  spice_node_2 n_n390(eclk, ereset, n390_i0,n390_i2, n390_v);
  spice_node_2 n_n397(eclk, ereset, n397_i0,n397_i1, n397_v);
  spice_node_3 n_n396(eclk, ereset, n396_i0,n396_i1,n396_i2, n396_v);
  spice_node_1 n_notalu0(eclk, ereset, notalu0_i1, notalu0_v);
  spice_node_3 n_ab11(eclk, ereset, ab11_i0,ab11_i1,ab11_i2, ab11_v);
  spice_node_1 n_n398(eclk, ereset, n398_i0, n398_v);
  spice_node_3 n_notir6(eclk, ereset, notir6_i0,notir6_i1,notir6_i2, notir6_v);
  spice_node_2 n_op_shift_right(eclk, ereset, op_shift_right_i0,op_shift_right_i1, op_shift_right_v);
  spice_node_2 n_op_T0_txs(eclk, ereset, op_T0_txs_i0,op_T0_txs_i2, op_T0_txs_v);
  spice_node_2 n_op_ror(eclk, ereset, op_ror_i1,op_ror_i2, op_ror_v);
  spice_node_2 n_dpc33_PCHDB(eclk, ereset, dpc33_PCHDB_i0,dpc33_PCHDB_i1, dpc33_PCHDB_v);
  spice_node_2 n_n241(eclk, ereset, n241_i2,n241_i3, n241_v);
  spice_node_3 n_idl5(eclk, ereset, idl5_i0,idl5_i1,idl5_i2, idl5_v);
  spice_node_2 n_n243(eclk, ereset, n243_i0,n243_i1, n243_v);
  spice_node_4 n_n242(eclk, ereset, n242_i0,n242_i1,n242_i2,n242_i3, n242_v);
  spice_node_2 n_n249(eclk, ereset, n249_i0,n249_i2, n249_v);
  spice_node_7 n_notRdy0(eclk, ereset, notRdy0_i0,notRdy0_i1,notRdy0_i3,notRdy0_i5,notRdy0_i6,notRdy0_i7,notRdy0_i8, notRdy0_v);
  spice_node_2 n_op_T0_txa(eclk, ereset, op_T0_txa_i0,op_T0_txa_i1, op_T0_txa_v);
  spice_node_2 n_abl7(eclk, ereset, abl7_i0,abl7_i4, abl7_v);
  spice_node_3 n_n177(eclk, ereset, n177_i0,n177_i1,n177_i2, n177_v);
  spice_node_3 n_n176(eclk, ereset, n176_i0,n176_i1,n176_i2, n176_v);
  spice_node_3 n_db5(eclk, ereset, db5_i0,db5_i3,db5_i4, db5_v);
  spice_node_2 n__AxB_6__C56(eclk, ereset, _AxB_6__C56_i0,_AxB_6__C56_i1, _AxB_6__C56_v);
  spice_node_2 n_n172(eclk, ereset, n172_i2,n172_i3, n172_v);
  spice_node_3 n_n171(eclk, ereset, n171_i0,n171_i1,n171_i3, n171_v);
  spice_node_1 n_pipeVectorA1(eclk, ereset, pipeVectorA1_i0, pipeVectorA1_v);
  spice_node_2 n_abl2(eclk, ereset, abl2_i3,abl2_i4, abl2_v);
  spice_node_3 n_n1500(eclk, ereset, n1500_i0,n1500_i1,n1500_i2, n1500_v);
  spice_node_2 n_pcl2(eclk, ereset, pcl2_i1,pcl2_i2, pcl2_v);
  spice_node_5 n_n652(eclk, ereset, n652_i0,n652_i1,n652_i2,n652_i3,n652_i4, n652_v);
  spice_node_3 n_n1507(eclk, ereset, n1507_i0,n1507_i1,n1507_i2, n1507_v);
  spice_node_2 n_op_T0_and(eclk, ereset, op_T0_and_i0,op_T0_and_i1, op_T0_and_v);
  spice_node_1 n_n1505(eclk, ereset, n1505_i0, n1505_v);
  spice_node_2 n_n1364(eclk, ereset, n1364_i0,n1364_i3, n1364_v);
  spice_node_3 n_n659(eclk, ereset, n659_i1,n659_i2,n659_i3, n659_v);
  spice_node_2 n_n1115(eclk, ereset, n1115_i0,n1115_i1, n1115_v);
  spice_node_5 n_n1618(eclk, ereset, n1618_i0,n1618_i1,n1618_i2,n1618_i3,n1618_i4, n1618_v);
  spice_node_2 n_n1619(eclk, ereset, n1619_i0,n1619_i1, n1619_v);
  spice_node_2 n_n1614(eclk, ereset, n1614_i0,n1614_i1, n1614_v);
  spice_node_2 n_op_T4_rts(eclk, ereset, op_T4_rts_i0,op_T4_rts_i1, op_T4_rts_v);
  spice_node_2 n_n1613(eclk, ereset, n1613_i1,n1613_i2, n1613_v);
  spice_node_2 n_n1610(eclk, ereset, n1610_i0,n1610_i1, n1610_v);
  spice_node_2 n_pcl7(eclk, ereset, pcl7_i1,pcl7_i2, pcl7_v);
  spice_node_2 n_op_T0_clc_sec(eclk, ereset, op_T0_clc_sec_i1,op_T0_clc_sec_i2, op_T0_clc_sec_v);
  spice_node_2 n_alua4(eclk, ereset, alua4_i0,alua4_i1, alua4_v);
  spice_node_2 n_abh4(eclk, ereset, abh4_i0,abh4_i4, abh4_v);
  spice_node_2 n_n1140(eclk, ereset, n1140_i1,n1140_i2, n1140_v);
  spice_node_3 n_n1141(eclk, ereset, n1141_i0,n1141_i1,n1141_i2, n1141_v);
  spice_node_2 n_alucout(eclk, ereset, alucout_i0,alucout_i2, alucout_v);
  spice_node_4 n_n1147(eclk, ereset, n1147_i0,n1147_i1,n1147_i2,n1147_i3, n1147_v);
  spice_node_2 n_DA_C45(eclk, ereset, DA_C45_i0,DA_C45_i1, DA_C45_v);
  spice_node_2 n_n1145(eclk, ereset, n1145_i1,n1145_i2, n1145_v);
  spice_node_2 n_y1(eclk, ereset, y1_i0,y1_i2, y1_v);
  spice_node_1 n_n1149(eclk, ereset, n1149_i0, n1149_v);
  spice_node_2 n_n692(eclk, ereset, n692_i2,n692_i3, n692_v);
  spice_node_2 n_BRtaken(eclk, ereset, BRtaken_i0,BRtaken_i2, BRtaken_v);
  spice_node_2 n_op_asl_rol(eclk, ereset, op_asl_rol_i0,op_asl_rol_i2, op_asl_rol_v);
  spice_node_3 n_n696(eclk, ereset, n696_i0,n696_i1,n696_i2, n696_v);
  spice_node_1 n_notalu1(eclk, ereset, notalu1_i1, notalu1_v);
  spice_node_5 n_n694(eclk, ereset, n694_i0,n694_i1,n694_i2,n694_i3,n694_i4, n694_v);
  spice_node_2 n_n1541(eclk, ereset, n1541_i2,n1541_i3, n1541_v);
  spice_node_1 n_n698(eclk, ereset, n698_i0, n698_v);
  spice_node_2 n__DA_ADD2(eclk, ereset, _DA_ADD2_i0,_DA_ADD2_i1, _DA_ADD2_v);
  spice_node_3 n_n1548(eclk, ereset, n1548_i0,n1548_i1,n1548_i2, n1548_v);
  spice_node_2 n_n1549(eclk, ereset, n1549_i1,n1549_i2, n1549_v);
  spice_node_2 n_n543(eclk, ereset, n543_i0,n543_i3, n543_v);
  spice_node_2 n_pd4_clearIR(eclk, ereset, pd4_clearIR_i1,pd4_clearIR_i5, pd4_clearIR_v);
  spice_node_2 n_n541(eclk, ereset, n541_i0,n541_i2, n541_v);
  spice_node_2 n_op_shift(eclk, ereset, op_shift_i0,op_shift_i1, op_shift_v);
  spice_node_2 n_n544(eclk, ereset, n544_i0,n544_i1, n544_v);
  spice_node_3 n_n548(eclk, ereset, n548_i0,n548_i1,n548_i2, n548_v);
  spice_node_2 n_dpc11_SBADD(eclk, ereset, dpc11_SBADD_i7,dpc11_SBADD_i9, dpc11_SBADD_v);
  spice_node_2 n_n761(eclk, ereset, n761_i1,n761_i2, n761_v);
  spice_node_2 n_dpc40_ADLPCL(eclk, ereset, dpc40_ADLPCL_i0,dpc40_ADLPCL_i9, dpc40_ADLPCL_v);
  spice_node_1 n_n415(eclk, ereset, n415_i1, n415_v);
  spice_node_2 n_n417(eclk, ereset, n417_i0,n417_i1, n417_v);
  spice_node_5 n_n1389(eclk, ereset, n1389_i0,n1389_i1,n1389_i2,n1389_i3,n1389_i4, n1389_v);
  spice_node_2 n_notalucout(eclk, ereset, notalucout_i1,notalucout_i2, notalucout_v);
  spice_node_8 n_adl0(eclk, ereset, adl0_i0,adl0_i1,adl0_i3,adl0_i4,adl0_i5,adl0_i6,adl0_i7,adl0_i8, adl0_v);
  spice_node_2 n_ir2(eclk, ereset, ir2_i0,ir2_i2, ir2_v);
  spice_node_2 n_op_T5_mem_ind_idx(eclk, ereset, op_T5_mem_ind_idx_i0,op_T5_mem_ind_idx_i2, op_T5_mem_ind_idx_v);
  spice_node_2 n_n1386(eclk, ereset, n1386_i0,n1386_i1, n1386_v);
  spice_node_4 n_n1387(eclk, ereset, n1387_i0,n1387_i1,n1387_i2,n1387_i3, n1387_v);
  spice_node_3 n_n1380(eclk, ereset, n1380_i1,n1380_i2,n1380_i3, n1380_v);
  spice_node_2 n_op_T3_jmp(eclk, ereset, op_T3_jmp_i1,op_T3_jmp_i2, op_T3_jmp_v);
  spice_node_3 n_brk_done(eclk, ereset, brk_done_i0,brk_done_i1,brk_done_i8, brk_done_v);
  spice_node_3 n_n1383(eclk, ereset, n1383_i0,n1383_i1,n1383_i2, n1383_v);
  spice_node_2 n_n368(eclk, ereset, n368_i1,n368_i2, n368_v);
  spice_node_1 n_pd4(eclk, ereset, pd4_i0, pd4_v);
  spice_node_2 n_n366(eclk, ereset, n366_i1,n366_i2, n366_v);
  spice_node_2 n__ABL4(eclk, ereset, _ABL4_i1,_ABL4_i2, _ABL4_v);
  spice_node_2 n_PD_0xx0xx0x(eclk, ereset, PD_0xx0xx0x_i1,PD_0xx0xx0x_i2, PD_0xx0xx0x_v);
  spice_node_2 n_dpc14_SRS(eclk, ereset, dpc14_SRS_i1,dpc14_SRS_i2, dpc14_SRS_v);
  spice_node_1 n_n360(eclk, ereset, n360_i0, n360_v);
  spice_node_1 n_pd1(eclk, ereset, pd1_i0, pd1_v);
  spice_node_3 n_n381(eclk, ereset, n381_i1,n381_i2,n381_i3, n381_v);
  spice_node_2 n_op_T0_iny_dey(eclk, ereset, op_T0_iny_dey_i0,op_T0_iny_dey_i1, op_T0_iny_dey_v);
  spice_node_2 n_n383(eclk, ereset, n383_i0,n383_i1, n383_v);
  spice_node_2 n_n384(eclk, ereset, n384_i1,n384_i2, n384_v);
  spice_node_3 n_n385(eclk, ereset, n385_i0,n385_i1,n385_i2, n385_v);
  spice_node_2 n_n386(eclk, ereset, n386_i0,n386_i2, n386_v);
  spice_node_2 n_n388(eclk, ereset, n388_i0,n388_i1, n388_v);
  spice_node_3 n_n389(eclk, ereset, n389_i0,n389_i1,n389_i2, n389_v);
  spice_node_2 n_op_T2_idx_x_xy(eclk, ereset, op_T2_idx_x_xy_i0,op_T2_idx_x_xy_i1, op_T2_idx_x_xy_v);
  spice_node_2 n_op_jsr(eclk, ereset, op_jsr_i0,op_jsr_i2, op_jsr_v);
  spice_node_3 n__op_set_C(eclk, ereset, _op_set_C_i0,_op_set_C_i1,_op_set_C_i2, _op_set_C_v);
  spice_node_2 n_n253(eclk, ereset, n253_i0,n253_i1, n253_v);
  spice_node_6 n_notaluoutmux1(eclk, ereset, notaluoutmux1_i0,notaluoutmux1_i1,notaluoutmux1_i2,notaluoutmux1_i3,notaluoutmux1_i4,notaluoutmux1_i5, notaluoutmux1_v);
  spice_node_2 n_n251(eclk, ereset, n251_i2,n251_i3, n251_v);
  spice_node_2 n_n256(eclk, ereset, n256_i0,n256_i1, n256_v);
  spice_node_2 n_op_T0_tya(eclk, ereset, op_T0_tya_i0,op_T0_tya_i1, op_T0_tya_v);
  spice_node_3 n_n254(eclk, ereset, n254_i0,n254_i1,n254_i2, n254_v);
  spice_node_2 n_n255(eclk, ereset, n255_i0,n255_i1, n255_v);
  spice_node_3 n_n168(eclk, ereset, n168_i0,n168_i1,n168_i2, n168_v);
  spice_node_3 n_n169(eclk, ereset, n169_i0,n169_i1,n169_i2, n169_v);
  spice_node_1 n_DC78_phi2(eclk, ereset, DC78_phi2_i0, DC78_phi2_v);
  spice_node_12 n_sb5(eclk, ereset, sb5_i0,sb5_i1,sb5_i2,sb5_i3,sb5_i4,sb5_i5,sb5_i6,sb5_i7,sb5_i8,sb5_i10,sb5_i11,sb5_i12, sb5_v);
  spice_node_2 n_op_T0_tax(eclk, ereset, op_T0_tax_i0,op_T0_tax_i1, op_T0_tax_v);
  spice_node_3 n_n160(eclk, ereset, n160_i0,n160_i1,n160_i2, n160_v);
  spice_node_2 n_n161(eclk, ereset, n161_i2,n161_i3, n161_v);
  spice_node_2 n_a3(eclk, ereset, a3_i0,a3_i1, a3_v);
  spice_node_2 n_n163(eclk, ereset, n163_i0,n163_i1, n163_v);
  spice_node_3 n_n1090(eclk, ereset, n1090_i0,n1090_i1,n1090_i2, n1090_v);
  spice_node_3 n_dasb6(eclk, ereset, dasb6_i0,dasb6_i1,dasb6_i2, dasb6_v);
  spice_node_3 n_n1093(eclk, ereset, n1093_i0,n1093_i1,n1093_i2, n1093_v);
  spice_node_2 n_s5(eclk, ereset, s5_i0,s5_i1, s5_v);
  spice_node_3 n_n1099(eclk, ereset, n1099_i0,n1099_i1,n1099_i2, n1099_v);
  spice_node_2 n_n1609(eclk, ereset, n1609_i0,n1609_i2, n1609_v);
  spice_node_2 n_n1608(eclk, ereset, n1608_i1,n1608_i2, n1608_v);
  spice_node_2 n_op_sty_cpy_mem(eclk, ereset, op_sty_cpy_mem_i0,op_sty_cpy_mem_i1, op_sty_cpy_mem_v);
  spice_node_2 n_n1600(eclk, ereset, n1600_i0,n1600_i1, n1600_v);
  spice_node_1 n_nots4(eclk, ereset, nots4_i0, nots4_v);
  spice_node_1 n_n1602(eclk, ereset, n1602_i1, n1602_v);
  spice_node_3 n_n1605(eclk, ereset, n1605_i0,n1605_i1,n1605_i3, n1605_v);
  spice_node_1 n_pipeUNK14(eclk, ereset, pipeUNK14_i0, pipeUNK14_v);
  spice_node_1 n_n1606(eclk, ereset, n1606_i0, n1606_v);
  spice_node_2 n_pd1_clearIR(eclk, ereset, pd1_clearIR_i1,pd1_clearIR_i3, pd1_clearIR_v);
  spice_node_3 n_alurawcout(eclk, ereset, alurawcout_i0,alurawcout_i1,alurawcout_i2, alurawcout_v);
  spice_node_2 n_n803(eclk, ereset, n803_i0,n803_i1, n803_v);
  spice_node_2 n_dpc0_YSB(eclk, ereset, dpc0_YSB_i3,dpc0_YSB_i9, dpc0_YSB_v);
  spice_node_2 n_n800(eclk, ereset, n800_i0,n800_i1, n800_v);
  spice_node_2 n_n807(eclk, ereset, n807_i0,n807_i1, n807_v);
  spice_node_0 n_n806(eclk, ereset,  n806_v);
  spice_node_1 n_n805(eclk, ereset, n805_i0, n805_v);
  spice_node_2 n_op_T4_brk_jsr(eclk, ereset, op_T4_brk_jsr_i0,op_T4_brk_jsr_i1, op_T4_brk_jsr_v);
  spice_node_2 n_n1159(eclk, ereset, n1159_i0,n1159_i1, n1159_v);
  spice_node_3 n_x_op_T__adc_sbc(eclk, ereset, x_op_T__adc_sbc_i0,x_op_T__adc_sbc_i1,x_op_T__adc_sbc_i2, x_op_T__adc_sbc_v);
  spice_node_2 n_n1154(eclk, ereset, n1154_i0,n1154_i2, n1154_v);
  spice_node_2 n_n1157(eclk, ereset, n1157_i0,n1157_i2, n1157_v);
  spice_node_3 n_rw(eclk, ereset, rw_i0,rw_i1,rw_i2, rw_v);
  spice_node_12 n_sb1(eclk, ereset, sb1_i0,sb1_i1,sb1_i2,sb1_i4,sb1_i5,sb1_i6,sb1_i7,sb1_i8,sb1_i9,sb1_i10,sb1_i11,sb1_i12, sb1_v);
  spice_node_2 n_n1153(eclk, ereset, n1153_i0,n1153_i3, n1153_v);
  spice_node_2 n_n1152(eclk, ereset, n1152_i0,n1152_i2, n1152_v);
  spice_node_2 n_dpc13_ORS(eclk, ereset, dpc13_ORS_i5,dpc13_ORS_i8, dpc13_ORS_v);
  spice_node_2 n_pch6(eclk, ereset, pch6_i0,pch6_i2, pch6_v);
  spice_node_1 n_p2(eclk, ereset, p2_i0, p2_v);
  spice_node_2 n_n1552(eclk, ereset, n1552_i0,n1552_i2, n1552_v);
  spice_node_2 n_op_T3_abs_idx(eclk, ereset, op_T3_abs_idx_i0,op_T3_abs_idx_i1, op_T3_abs_idx_v);
  spice_node_2 n_op_brk_rti(eclk, ereset, op_brk_rti_i0,op_brk_rti_i2, op_brk_rti_v);
  spice_node_1 n_pipeUNK34(eclk, ereset, pipeUNK34_i0, pipeUNK34_v);
  spice_node_1 n_n50(eclk, ereset, n50_i0, n50_v);
  spice_node_2 n_op_lsr_ror_dec_inc(eclk, ereset, op_lsr_ror_dec_inc_i0,op_lsr_ror_dec_inc_i2, op_lsr_ror_dec_inc_v);
  spice_node_6 n_adh1(eclk, ereset, adh1_i0,adh1_i1,adh1_i2,adh1_i4,adh1_i5,adh1_i6, adh1_v);
  spice_node_1 n_pipeT_SYNC(eclk, ereset, pipeT_SYNC_i0, pipeT_SYNC_v);
  spice_node_1 n_pclp7(eclk, ereset, pclp7_i1, pclp7_v);
  spice_node_2 n_pchp7(eclk, ereset, pchp7_i0,pchp7_i2, pchp7_v);
  spice_node_2 n_dpc23_SBAC(eclk, ereset, dpc23_SBAC_i8,dpc23_SBAC_i9, dpc23_SBAC_v);
  spice_node_3 n_n533(eclk, ereset, n533_i0,n533_i1,n533_i2, n533_v);
  spice_node_3 n___AxBxC_7(eclk, ereset, __AxBxC_7_i0,__AxBxC_7_i1,__AxBxC_7_i2, __AxBxC_7_v);
  spice_node_2 n_n531(eclk, ereset, n531_i0,n531_i3, n531_v);
  spice_node_13 n_dasb0(eclk, ereset, dasb0_i0,dasb0_i1,dasb0_i2,dasb0_i3,dasb0_i4,dasb0_i5,dasb0_i6,dasb0_i7,dasb0_i8,dasb0_i9,dasb0_i10,dasb0_i11,dasb0_i12, dasb0_v);
  spice_node_3 n_sync(eclk, ereset, sync_i0,sync_i1,sync_i2, sync_v);
  spice_node_2 n_n538(eclk, ereset, n538_i0,n538_i1, n538_v);
  spice_node_2 n__ABH7(eclk, ereset, _ABH7_i1,_ABH7_i2, _ABH7_v);
  spice_node_3 n_n428(eclk, ereset, n428_i0,n428_i1,n428_i2, n428_v);
  spice_node_2 n_n1399(eclk, ereset, n1399_i0,n1399_i3, n1399_v);
  spice_node_3 n_n1398(eclk, ereset, n1398_i0,n1398_i2,n1398_i4, n1398_v);
  spice_node_2 n_op_T0_shift_a(eclk, ereset, op_T0_shift_a_i0,op_T0_shift_a_i2, op_T0_shift_a_v);
  spice_node_1 n_n1395(eclk, ereset, n1395_i0, n1395_v);
  spice_node_3 n_notir5(eclk, ereset, notir5_i0,notir5_i2,notir5_i3, notir5_v);
  spice_node_3 n_db4(eclk, ereset, db4_i0,db4_i3,db4_i4, db4_v);
  spice_node_2 n_n1392(eclk, ereset, n1392_i1,n1392_i2, n1392_v);
  spice_node_2 n__C56(eclk, ereset, _C56_i1,_C56_i2, _C56_v);
  spice_node_2 n_alua5(eclk, ereset, alua5_i0,alua5_i1, alua5_v);
  spice_node_3 n__TWOCYCLE(eclk, ereset, _TWOCYCLE_i0,_TWOCYCLE_i1,_TWOCYCLE_i2, _TWOCYCLE_v);
  spice_node_2 n_n853(eclk, ereset, n853_i0,n853_i1, n853_v);
  spice_node_1 n_pipeUNK26(eclk, ereset, pipeUNK26_i1, pipeUNK26_v);
  spice_node_2 n_dpc28_0ADH0(eclk, ereset, dpc28_0ADH0_i0,dpc28_0ADH0_i2, dpc28_0ADH0_v);
  spice_node_2 n_n228(eclk, ereset, n228_i0,n228_i1, n228_v);
  spice_node_3 n_n227(eclk, ereset, n227_i0,n227_i1,n227_i2, n227_v);
  spice_node_1 n_n226(eclk, ereset, n226_i0, n226_v);
  spice_node_2 n_n225(eclk, ereset, n225_i0,n225_i1, n225_v);
  spice_node_2 n_n224(eclk, ereset, n224_i1,n224_i2, n224_v);
  spice_node_1 n_n223(eclk, ereset, n223_i1, n223_v);
  spice_node_1 n_notdor0(eclk, ereset, notdor0_i0, notdor0_v);
  spice_node_2 n_n221(eclk, ereset, n221_i0,n221_i1, n221_v);
  spice_node_2 n_n220(eclk, ereset, n220_i0,n220_i3, n220_v);
  spice_node_1 n_pipeUNK39(eclk, ereset, pipeUNK39_i0, pipeUNK39_v);
  spice_node_2 n__ABL0(eclk, ereset, _ABL0_i1,_ABL0_i2, _ABL0_v);
  spice_node_2 n_n152(eclk, ereset, n152_i0,n152_i1, n152_v);
  spice_node_3 n_aluanorb1(eclk, ereset, aluanorb1_i1,aluanorb1_i2,aluanorb1_i3, aluanorb1_v);
  spice_node_2 n_n154(eclk, ereset, n154_i2,n154_i3, n154_v);
  spice_node_2 n_op_T2_stack_access(eclk, ereset, op_T2_stack_access_i0,op_T2_stack_access_i2, op_T2_stack_access_v);
  spice_node_2 n_clock2(eclk, ereset, clock2_i0,clock2_i1, clock2_v);
  spice_node_1 n_res(eclk, ereset, res_i1, res_v);
  spice_node_1 n_notdor7(eclk, ereset, notdor7_i0, notdor7_v);
  spice_node_2 n_n1293(eclk, ereset, n1293_i0,n1293_i2, n1293_v);
  spice_node_2 n_n1256(eclk, ereset, n1256_i0,n1256_i2, n1256_v);
  spice_node_2 n_t4(eclk, ereset, t4_i0,t4_i2, t4_v);
  spice_node_3 n___AxB_0(eclk, ereset, __AxB_0_i0,__AxB_0_i1,__AxB_0_i3, __AxB_0_v);
  spice_node_3 n_n1526(eclk, ereset, n1526_i0,n1526_i1,n1526_i2, n1526_v);
  spice_node_2 n_n818(eclk, ereset, n818_i2,n818_i3, n818_v);
  spice_node_2 n_n819(eclk, ereset, n819_i0,n819_i2, n819_v);
  spice_node_2 n_n1255(eclk, ereset, n1255_i1,n1255_i2, n1255_v);
  spice_node_2 n_n810(eclk, ereset, n810_i0,n810_i1, n810_v);
  spice_node_2 n_n811(eclk, ereset, n811_i0,n811_i1, n811_v);
  spice_node_2 n_n812(eclk, ereset, n812_i0,n812_i1, n812_v);
  spice_node_2 n_n813(eclk, ereset, n813_i0,n813_i1, n813_v);
  spice_node_2 n_n815(eclk, ereset, n815_i0,n815_i2, n815_v);
  spice_node_2 n___AxB5__C45(eclk, ereset, __AxB5__C45_i0,__AxB5__C45_i1, __AxB5__C45_v);
  spice_node_2 n_abl3(eclk, ereset, abl3_i3,abl3_i4, abl3_v);
  spice_node_4 n_n1251(eclk, ereset, n1251_i0,n1251_i1,n1251_i2,n1251_i3, n1251_v);
  spice_node_1 n_notalu4(eclk, ereset, notalu4_i1, notalu4_v);
  spice_node_4 n_n1491(eclk, ereset, n1491_i0,n1491_i1,n1491_i2,n1491_i3, n1491_v);
  spice_node_2 n_n1492(eclk, ereset, n1492_i0,n1492_i1, n1492_v);
  spice_node_3 n_ab7(eclk, ereset, ab7_i0,ab7_i1,ab7_i2, ab7_v);
  spice_node_3 n_dasb7(eclk, ereset, dasb7_i0,dasb7_i1,dasb7_i2, dasb7_v);
  spice_node_3 n_n1495(eclk, ereset, n1495_i0,n1495_i1,n1495_i2, n1495_v);
  spice_node_5 n_n1496(eclk, ereset, n1496_i0,n1496_i1,n1496_i2,n1496_i3,n1496_i4, n1496_v);
  spice_node_3 n_n1497(eclk, ereset, n1497_i0,n1497_i1,n1497_i2, n1497_v);
  spice_node_2 n_n1499(eclk, ereset, n1499_i0,n1499_i3, n1499_v);
  spice_node_3 n_n423(eclk, ereset, n423_i0,n423_i1,n423_i2, n423_v);
  spice_node_2 n_dpc4_SSB(eclk, ereset, dpc4_SSB_i0,dpc4_SSB_i9, dpc4_SSB_v);
  spice_node_2 n_s4(eclk, ereset, s4_i0,s4_i1, s4_v);
  spice_node_2 n_dpc34_PCLC(eclk, ereset, dpc34_PCLC_i1,dpc34_PCLC_i2, dpc34_PCLC_v);
  spice_node_3 n_n1705(eclk, ereset, n1705_i0,n1705_i1,n1705_i2, n1705_v);
  spice_node_2 n_n1708(eclk, ereset, n1708_i1,n1708_i2, n1708_v);
  spice_node_4 n_n1709(eclk, ereset, n1709_i0,n1709_i1,n1709_i2,n1709_i3, n1709_v);
  spice_node_2 n_n424(eclk, ereset, n424_i1,n424_i2, n424_v);
  spice_node_3 n_n1391(eclk, ereset, n1391_i0,n1391_i1,n1391_i2, n1391_v);
  spice_node_2 n__ABH5(eclk, ereset, _ABH5_i1,_ABH5_i2, _ABH5_v);
  spice_node_2 n_n1129(eclk, ereset, n1129_i2,n1129_i3, n1129_v);
  spice_node_2 n_n1120(eclk, ereset, n1120_i0,n1120_i1, n1120_v);
  spice_node_1 n_n1121(eclk, ereset, n1121_i1, n1121_v);
  spice_node_2 n__C12(eclk, ereset, _C12_i1,_C12_i2, _C12_v);
  spice_node_1 n_notalu7(eclk, ereset, notalu7_i1, notalu7_v);
  spice_node_1 n_n1124(eclk, ereset, n1124_i1, n1124_v);
  spice_node_3 n_notir3(eclk, ereset, notir3_i0,notir3_i1,notir3_i2, notir3_v);
  spice_node_1 n_n1126(eclk, ereset, n1126_i0, n1126_v);
  spice_node_2 n_n525(eclk, ereset, n525_i2,n525_i3, n525_v);
  spice_node_1 n_n526(eclk, ereset, n526_i1, n526_v);
  spice_node_1 n_notdor1(eclk, ereset, notdor1_i1, notdor1_v);
  spice_node_2 n_n520(eclk, ereset, n520_i0,n520_i2, n520_v);
  spice_node_1 n_n521(eclk, ereset, n521_i0, n521_v);
  spice_node_3 n_op_ORS(eclk, ereset, op_ORS_i0,op_ORS_i1,op_ORS_i2, op_ORS_v);
  spice_node_2 n_n523(eclk, ereset, n523_i0,n523_i3, n523_v);
  spice_node_4 n_n1014(eclk, ereset, n1014_i0,n1014_i1,n1014_i2,n1014_i3, n1014_v);
  spice_node_2 n_dpc21_ADDADL(eclk, ereset, dpc21_ADDADL_i0,dpc21_ADDADL_i9, dpc21_ADDADL_v);
  spice_node_3 n_n1016(eclk, ereset, n1016_i0,n1016_i1,n1016_i2, n1016_v);
  spice_node_2 n_n1017(eclk, ereset, n1017_i0,n1017_i2, n1017_v);
  spice_node_2 n_n1010(eclk, ereset, n1010_i0,n1010_i2, n1010_v);
  spice_node_1 n_pipeUNK11(eclk, ereset, pipeUNK11_i1, pipeUNK11_v);
  spice_node_2 n_a1(eclk, ereset, a1_i0,a1_i1, a1_v);
  spice_node_2 n_dpc32_PCHADH(eclk, ereset, dpc32_PCHADH_i0,dpc32_PCHADH_i1, dpc32_PCHADH_v);
  spice_node_2 n_A_B5(eclk, ereset, A_B5_i0,A_B5_i1, A_B5_v);
  spice_node_3 n_ab12(eclk, ereset, ab12_i0,ab12_i1,ab12_i2, ab12_v);
  spice_node_2 n_n1230(eclk, ereset, n1230_i2,n1230_i3, n1230_v);
  spice_node_3 n_n1231(eclk, ereset, n1231_i0,n1231_i1,n1231_i2, n1231_v);
  spice_node_2 n_abl4(eclk, ereset, abl4_i0,abl4_i4, abl4_v);
  spice_node_2 n_op_T0_cpy_iny(eclk, ereset, op_T0_cpy_iny_i0,op_T0_cpy_iny_i1, op_T0_cpy_iny_v);
  spice_node_2 n_n1238(eclk, ereset, n1238_i1,n1238_i2, n1238_v);
  spice_node_2 n_op_T2_branch(eclk, ereset, op_T2_branch_i1,op_T2_branch_i2, op_T2_branch_v);
  spice_node_2 n_dpc38_PCLADL(eclk, ereset, dpc38_PCLADL_i0,dpc38_PCLADL_i9, dpc38_PCLADL_v);
  spice_node_3 n_Pout3(eclk, ereset, Pout3_i0,Pout3_i1,Pout3_i2, Pout3_v);
  spice_node_4 n_n436(eclk, ereset, n436_i0,n436_i1,n436_i2,n436_i3, n436_v);
  spice_node_2 n_dpc10_ADLADD(eclk, ereset, dpc10_ADLADD_i2,dpc10_ADLADD_i9, dpc10_ADLADD_v);
  spice_node_2 n_op_rmw(eclk, ereset, op_rmw_i0,op_rmw_i1, op_rmw_v);
  spice_node_3 n_ab4(eclk, ereset, ab4_i0,ab4_i1,ab4_i2, ab4_v);
  spice_node_2 n_n432(eclk, ereset, n432_i0,n432_i1, n432_v);
  spice_node_4 n_n430(eclk, ereset, n430_i0,n430_i1,n430_i2,n430_i3, n430_v);
  spice_node_2 n_n238(eclk, ereset, n238_i0,n238_i1, n238_v);
  spice_node_2 n_abl5(eclk, ereset, abl5_i0,abl5_i4, abl5_v);
  spice_node_3 n_alub6(eclk, ereset, alub6_i0,alub6_i1,alub6_i2, alub6_v);
  spice_node_2 n_n236(eclk, ereset, n236_i1,n236_i2, n236_v);
  spice_node_3 n_ab8(eclk, ereset, ab8_i0,ab8_i1,ab8_i2, ab8_v);
  spice_node_2 n_n231(eclk, ereset, n231_i1,n231_i2, n231_v);
  spice_node_2 n_n232(eclk, ereset, n232_i0,n232_i1, n232_v);
  spice_node_2 n_n233(eclk, ereset, n233_i0,n233_i1, n233_v);
  spice_node_2 n_x2(eclk, ereset, x2_i0,x2_i1, x2_v);
  spice_node_5 n_n146(eclk, ereset, n146_i0,n146_i1,n146_i2,n146_i3,n146_i4, n146_v);
  spice_node_2 n_n147(eclk, ereset, n147_i1,n147_i2, n147_v);
  spice_node_2 n_op_sta_cmp(eclk, ereset, op_sta_cmp_i0,op_sta_cmp_i1, op_sta_cmp_v);
  spice_node_2 n_C45(eclk, ereset, C45_i1,C45_i2, C45_v);
  spice_node_3 n_aluanorb0(eclk, ereset, aluanorb0_i0,aluanorb0_i2,aluanorb0_i3, aluanorb0_v);
  spice_node_2 n_dpc27_SBADH(eclk, ereset, dpc27_SBADH_i0,dpc27_SBADH_i9, dpc27_SBADH_v);
  spice_node_5 n_n141(eclk, ereset, n141_i0,n141_i1,n141_i2,n141_i3,n141_i4, n141_v);
  spice_node_3 n_ab9(eclk, ereset, ab9_i0,ab9_i1,ab9_i2, ab9_v);
  spice_node_2 n_n149(eclk, ereset, n149_i0,n149_i1, n149_v);
  spice_node_2 n_aluvout(eclk, ereset, aluvout_i0,aluvout_i2, aluvout_v);
  spice_node_2 n_n933(eclk, ereset, n933_i0,n933_i2, n933_v);
  spice_node_2 n_op_T2_php_pha(eclk, ereset, op_T2_php_pha_i0,op_T2_php_pha_i1, op_T2_php_pha_v);
  spice_node_3 n_n931(eclk, ereset, n931_i0,n931_i1,n931_i2, n931_v);
  spice_node_2 n_n930(eclk, ereset, n930_i0,n930_i1, n930_v);
  spice_node_2 n_n937(eclk, ereset, n937_i0,n937_i1, n937_v);
  spice_node_2 n_n936(eclk, ereset, n936_i0,n936_i1, n936_v);
  spice_node_3 n_n935(eclk, ereset, n935_i0,n935_i1,n935_i2, n935_v);
  spice_node_4 n_op_SRS(eclk, ereset, op_SRS_i0,op_SRS_i2,op_SRS_i3,op_SRS_i4, op_SRS_v);
  spice_node_1 n_pd5(eclk, ereset, pd5_i0, pd5_v);
  spice_node_1 n_nots3(eclk, ereset, nots3_i0, nots3_v);
  spice_node_2 n__ABL3(eclk, ereset, _ABL3_i0,_ABL3_i2, _ABL3_v);
  spice_node_4 n_n824(eclk, ereset, n824_i0,n824_i1,n824_i2,n824_i3, n824_v);
  spice_node_3 n_D1x1(eclk, ereset, D1x1_i0,D1x1_i2,D1x1_i3, D1x1_v);
  spice_node_2 n_n826(eclk, ereset, n826_i1,n826_i2, n826_v);
  spice_node_2 n_ADH_ABH(eclk, ereset, ADH_ABH_i0,ADH_ABH_i1, ADH_ABH_v);
  spice_node_1 n_pchp4(eclk, ereset, pchp4_i1, pchp4_v);
  spice_node_1 n_notdor3(eclk, ereset, notdor3_i0, notdor3_v);
  spice_node_2 n_op_T__adc_sbc(eclk, ereset, op_T__adc_sbc_i0,op_T__adc_sbc_i2, op_T__adc_sbc_v);
  spice_node_2 n_op_T__iny_dey(eclk, ereset, op_T__iny_dey_i0,op_T__iny_dey_i1, op_T__iny_dey_v);
  spice_node_3 n_VEC1(eclk, ereset, VEC1_i0,VEC1_i1,VEC1_i2, VEC1_v);
  spice_node_2 n_op_T3_plp_pla(eclk, ereset, op_T3_plp_pla_i0,op_T3_plp_pla_i2, op_T3_plp_pla_v);
  spice_node_3 n_n1486(eclk, ereset, n1486_i0,n1486_i1,n1486_i2, n1486_v);
  spice_node_1 n_notidl2(eclk, ereset, notidl2_i1, notidl2_v);
  spice_node_2 n_n1484(eclk, ereset, n1484_i0,n1484_i2, n1484_v);
  spice_node_2 n_n1488(eclk, ereset, n1488_i0,n1488_i1, n1488_v);
  spice_node_3 n_n797(eclk, ereset, n797_i0,n797_i1,n797_i2, n797_v);
  spice_node_1 n_n796(eclk, ereset, n796_i0, n796_v);
  spice_node_3 n_n795(eclk, ereset, n795_i0,n795_i1,n795_i2, n795_v);
  spice_node_2 n_n794(eclk, ereset, n794_i0,n794_i2, n794_v);
  spice_node_3 n_n1717(eclk, ereset, n1717_i0,n1717_i1,n1717_i2, n1717_v);
  spice_node_2 n_n1716(eclk, ereset, n1716_i0,n1716_i1, n1716_v);
  spice_node_2 n_op_push_pull(eclk, ereset, op_push_pull_i0,op_push_pull_i1, op_push_pull_v);
  spice_node_2 n_n790(eclk, ereset, n790_i1,n790_i3, n790_v);
  spice_node_2 n_n1719(eclk, ereset, n1719_i0,n1719_i2, n1719_v);
  spice_node_3 n_n1718(eclk, ereset, n1718_i0,n1718_i1,n1718_i2, n1718_v);
  spice_node_1 n_n799(eclk, ereset, n799_i1, n799_v);
  spice_node_2 n_n798(eclk, ereset, n798_i1,n798_i2, n798_v);
  spice_node_2 n_n1270(eclk, ereset, n1270_i2,n1270_i3, n1270_v);
  spice_node_2 n_n1271(eclk, ereset, n1271_i0,n1271_i2, n1271_v);
  spice_node_1 n_n610(eclk, ereset, n610_i1, n610_v);
  spice_node_2 n_pcl0(eclk, ereset, pcl0_i1,pcl0_i2, pcl0_v);
  spice_node_2 n_n1138(eclk, ereset, n1138_i0,n1138_i2, n1138_v);
  spice_node_2 n_n1133(eclk, ereset, n1133_i1,n1133_i2, n1133_v);
  spice_node_1 n_n1132(eclk, ereset, n1132_i0, n1132_v);
  spice_node_1 n_pipe_WR_phi2(eclk, ereset, pipe_WR_phi2_i0, pipe_WR_phi2_v);
  spice_node_3 n_n1130(eclk, ereset, n1130_i0,n1130_i1,n1130_i2, n1130_v);
  spice_node_2 n_n1137(eclk, ereset, n1137_i0,n1137_i2, n1137_v);
  spice_node_2 n_a6(eclk, ereset, a6_i0,a6_i2, a6_v);
  spice_node_2 n_n1135(eclk, ereset, n1135_i0,n1135_i1, n1135_v);
  spice_node_3 n__VEC(eclk, ereset, _VEC_i0,_VEC_i1,_VEC_i3, _VEC_v);
  spice_node_1 n_n1276(eclk, ereset, n1276_i0, n1276_v);
  spice_node_2 n_n1277(eclk, ereset, n1277_i0,n1277_i3, n1277_v);
  spice_node_2 n_n519(eclk, ereset, n519_i1,n519_i3, n519_v);
  spice_node_4 n_n518(eclk, ereset, n518_i0,n518_i1,n518_i2,n518_i3, n518_v);
  spice_node_3 n_dasb1(eclk, ereset, dasb1_i0,dasb1_i1,dasb1_i2, dasb1_v);
  spice_node_1 n_pipeUNK29(eclk, ereset, pipeUNK29_i0, pipeUNK29_v);
  spice_node_2 n_n1007(eclk, ereset, n1007_i0,n1007_i1, n1007_v);
  spice_node_2 n_op_implied(eclk, ereset, op_implied_i1,op_implied_i2, op_implied_v);
  spice_node_3 n_db0(eclk, ereset, db0_i1,db0_i3,db0_i4, db0_v);
  spice_node_2 n__C23(eclk, ereset, _C23_i0,_C23_i1, _C23_v);
  spice_node_2 n_n1002(eclk, ereset, n1002_i0,n1002_i1, n1002_v);
  spice_node_2 n_op_store(eclk, ereset, op_store_i1,op_store_i2, op_store_v);
  spice_node_2 n_pclp0(eclk, ereset, pclp0_i1,pclp0_i2, pclp0_v);
  spice_node_2 n_op_T0_plp(eclk, ereset, op_T0_plp_i0,op_T0_plp_i1, op_T0_plp_v);
  spice_node_4 n_n1225(eclk, ereset, n1225_i1,n1225_i2,n1225_i3,n1225_i4, n1225_v);
  spice_node_2 n_n620(eclk, ereset, n620_i0,n620_i1, n620_v);
  spice_node_2 n_n1223(eclk, ereset, n1223_i2,n1223_i3, n1223_v);
  spice_node_3 n_n626(eclk, ereset, n626_i0,n626_i1,n626_i2, n626_v);
  spice_node_2 n_n625(eclk, ereset, n625_i2,n625_i3, n625_v);
  spice_node_2 n_AxB5(eclk, ereset, AxB5_i1,AxB5_i3, AxB5_v);
  spice_node_3 n_n629(eclk, ereset, n629_i0,n629_i1,n629_i2, n629_v);
  spice_node_2 n_n628(eclk, ereset, n628_i2,n628_i3, n628_v);
  spice_node_3 n_n1229(eclk, ereset, n1229_i0,n1229_i1,n1229_i2, n1229_v);
  spice_node_3 n_op_ANDS(eclk, ereset, op_ANDS_i0,op_ANDS_i1,op_ANDS_i2, op_ANDS_v);
  spice_node_3 n_alub7(eclk, ereset, alub7_i0,alub7_i1,alub7_i2, alub7_v);
  spice_node_2 n_n1286(eclk, ereset, n1286_i0,n1286_i1, n1286_v);
  spice_node_3 n_n11(eclk, ereset, n11_i0,n11_i1,n11_i2, n11_v);
  spice_node_2 n_n10(eclk, ereset, n10_i0,n10_i2, n10_v);
  spice_node_6 n_adh6(eclk, ereset, adh6_i0,adh6_i1,adh6_i3,adh6_i4,adh6_i5,adh6_i6, adh6_v);
  spice_node_1 n_n15(eclk, ereset, n15_i0, n15_v);
  spice_node_3 n_n14(eclk, ereset, n14_i0,n14_i1,n14_i2, n14_v);
  spice_node_3 n_n17(eclk, ereset, n17_i2,n17_i3,n17_i4, n17_v);
  spice_node_2 n_n16(eclk, ereset, n16_i0,n16_i1, n16_v);
  spice_node_3 n_n19(eclk, ereset, n19_i0,n19_i1,n19_i2, n19_v);
  spice_node_1 n_n18(eclk, ereset, n18_i0, n18_v);
  spice_node_1 n_n688(eclk, ereset, n688_i0, n688_v);
  spice_node_2 n_n201(eclk, ereset, n201_i0,n201_i1, n201_v);
  spice_node_2 n_n200(eclk, ereset, n200_i0,n200_i1, n200_v);
  spice_node_2 n_dpc29_0ADH17(eclk, ereset, dpc29_0ADH17_i1,dpc29_0ADH17_i2, dpc29_0ADH17_v);
  spice_node_2 n_pch7(eclk, ereset, pch7_i1,pch7_i2, pch7_v);
  spice_node_2 n_op_T2_ADL_ADD(eclk, ereset, op_T2_ADL_ADD_i0,op_T2_ADL_ADD_i1, op_T2_ADL_ADD_v);
  spice_node_3 n_n207(eclk, ereset, n207_i0,n207_i1,n207_i2, n207_v);
  spice_node_3 n_n206(eclk, ereset, n206_i0,n206_i1,n206_i3, n206_v);
  spice_node_5 n_n209(eclk, ereset, n209_i0,n209_i1,n209_i2,n209_i3,n209_i4, n209_v);
  spice_node_5 n_n208(eclk, ereset, n208_i0,n208_i1,n208_i2,n208_i3,n208_i4, n208_v);
  spice_node_2 n_n1573(eclk, ereset, n1573_i0,n1573_i1, n1573_v);
  spice_node_7 n_adl3(eclk, ereset, adl3_i0,adl3_i1,adl3_i2,adl3_i3,adl3_i4,adl3_i6,adl3_i7, adl3_v);
  spice_node_2 n__C45(eclk, ereset, _C45_i1,_C45_i2, _C45_v);
  spice_node_2 n_n_0_ADL1(eclk, ereset, n_0_ADL1_i0,n_0_ADL1_i2, n_0_ADL1_v);
  spice_node_1 n_pipeUNK15(eclk, ereset, pipeUNK15_i1, pipeUNK15_v);
  spice_node_1 n_n680(eclk, ereset, n680_i0, n680_v);
  spice_node_1 n_pipedpc28(eclk, ereset, pipedpc28_i0, pipedpc28_v);
  spice_node_1 n_n1574(eclk, ereset, n1574_i0, n1574_v);
  spice_node_3 n_n928(eclk, ereset, n928_i0,n928_i1,n928_i2, n928_v);
  spice_node_5 n_n929(eclk, ereset, n929_i0,n929_i1,n929_i2,n929_i3,n929_i4, n929_v);
  spice_node_3 n_n920(eclk, ereset, n920_i0,n920_i1,n920_i2, n920_v);
  spice_node_2 n_dpc17_SUMS(eclk, ereset, dpc17_SUMS_i0,dpc17_SUMS_i1, dpc17_SUMS_v);
  spice_node_2 n_n923(eclk, ereset, n923_i0,n923_i1, n923_v);
  spice_node_2 n__op_store(eclk, ereset, _op_store_i0,_op_store_i1, _op_store_v);
  spice_node_2 n_C1x5Reset(eclk, ereset, C1x5Reset_i1,C1x5Reset_i2, C1x5Reset_v);
  spice_node_2 n_n927(eclk, ereset, n927_i0,n927_i2, n927_v);
  spice_node_1 n_pipeUNK19(eclk, ereset, pipeUNK19_i0, pipeUNK19_v);
  spice_node_8 n_idb6(eclk, ereset, idb6_i0,idb6_i2,idb6_i4,idb6_i5,idb6_i6,idb6_i8,idb6_i9,idb6_i10, idb6_v);
  spice_node_2 n_n830(eclk, ereset, n830_i2,n830_i3, n830_v);
  spice_node_5 n_n831(eclk, ereset, n831_i0,n831_i1,n831_i2,n831_i3,n831_i4, n831_v);
  spice_node_2 n_n837(eclk, ereset, n837_i0,n837_i2, n837_v);
  spice_node_2 n_n834(eclk, ereset, n834_i2,n834_i4, n834_v);
  spice_node_2 n_n838(eclk, ereset, n838_i0,n838_i1, n838_v);
  spice_node_2 n_n839(eclk, ereset, n839_i1,n839_i2, n839_v);
  spice_node_5 n_n3(eclk, ereset, n3_i0,n3_i1,n3_i2,n3_i3,n3_i4, n3_v);
  spice_node_2 n_op_T5_rti(eclk, ereset, op_T5_rti_i0,op_T5_rti_i2, op_T5_rti_v);
  spice_node_1 n_n785(eclk, ereset, n785_i0, n785_v);
  spice_node_2 n_op_T__dex(eclk, ereset, op_T__dex_i0,op_T__dex_i1, op_T__dex_v);
  spice_node_2 n_op_T0_sbc(eclk, ereset, op_T0_sbc_i0,op_T0_sbc_i1, op_T0_sbc_v);
  spice_node_1 n_pchp0(eclk, ereset, pchp0_i1, pchp0_v);
  spice_node_2 n_n781(eclk, ereset, n781_i0,n781_i3, n781_v);
  spice_node_2 n_n782(eclk, ereset, n782_i0,n782_i2, n782_v);
  spice_node_2 n_n783(eclk, ereset, n783_i0,n783_i1, n783_v);
  spice_node_4 n_n1724(eclk, ereset, n1724_i0,n1724_i1,n1724_i2,n1724_i3, n1724_v);
  spice_node_2 n_op_T2(eclk, ereset, op_T2_i0,op_T2_i1, op_T2_v);
  spice_node_3 n_n789(eclk, ereset, n789_i0,n789_i1,n789_i2, n789_v);
  spice_node_2 n_n1720(eclk, ereset, n1720_i1,n1720_i2, n1720_v);
  spice_node_2 n_op_branch_done(eclk, ereset, op_branch_done_i1,op_branch_done_i2, op_branch_done_v);
  spice_node_2 n_op_T3_ind_y(eclk, ereset, op_T3_ind_y_i0,op_T3_ind_y_i1, op_T3_ind_y_v);
  spice_node_2 n_n61(eclk, ereset, n61_i0,n61_i1, n61_v);
  spice_node_3 n_n62(eclk, ereset, n62_i0,n62_i1,n62_i2, n62_v);
  spice_node_2 n_dor7(eclk, ereset, dor7_i0,dor7_i2, dor7_v);
  spice_node_2 n_y0(eclk, ereset, y0_i0,y0_i2, y0_v);
  spice_node_2 n__AxB_4__C34(eclk, ereset, _AxB_4__C34_i0,_AxB_4__C34_i1, _AxB_4__C34_v);
  spice_node_3 n_n66(eclk, ereset, n66_i1,n66_i2,n66_i3, n66_v);
  spice_node_4 n_Reset0(eclk, ereset, Reset0_i0,Reset0_i1,Reset0_i2,Reset0_i3, Reset0_v);
  spice_node_1 n_notalu6(eclk, ereset, notalu6_i1, notalu6_v);
  spice_node_1 n_n69(eclk, ereset, n69_i0, n69_v);
  spice_node_6 n_adh0(eclk, ereset, adh0_i0,adh0_i1,adh0_i2,adh0_i3,adh0_i4,adh0_i6, adh0_v);
  spice_node_3 n_n1588(eclk, ereset, n1588_i0,n1588_i1,n1588_i2, n1588_v);
  spice_node_2 n_op_T4_jmp(eclk, ereset, op_T4_jmp_i0,op_T4_jmp_i1, op_T4_jmp_v);
  spice_node_2 n_op_T2_stack(eclk, ereset, op_T2_stack_i0,op_T2_stack_i1, op_T2_stack_v);
  spice_node_2 n_n1580(eclk, ereset, n1580_i0,n1580_i1, n1580_v);
  spice_node_1 n_n1581(eclk, ereset, n1581_i0, n1581_v);
  spice_node_3 n_n1586(eclk, ereset, n1586_i0,n1586_i1,n1586_i2, n1586_v);
  spice_node_1 n_pipeT4out(eclk, ereset, pipeT4out_i0, pipeT4out_v);
  spice_node_2 n_n1585(eclk, ereset, n1585_i1,n1585_i2, n1585_v);
  spice_node_2 n_n1038(eclk, ereset, n1038_i0,n1038_i1, n1038_v);
  spice_node_2 n_DC34(eclk, ereset, DC34_i0,DC34_i1, DC34_v);
  spice_node_1 n_n509(eclk, ereset, n509_i0, n509_v);
  spice_node_2 n_NMIP(eclk, ereset, NMIP_i1,NMIP_i3, NMIP_v);
  spice_node_2 n_op_T0_ora(eclk, ereset, op_T0_ora_i0,op_T0_ora_i1, op_T0_ora_v);
  spice_node_2 n_op_T3_stack_bit_jmp(eclk, ereset, op_T3_stack_bit_jmp_i0,op_T3_stack_bit_jmp_i1, op_T3_stack_bit_jmp_v);
  spice_node_2 n_pch2(eclk, ereset, pch2_i0,pch2_i1, pch2_v);
  spice_node_3 n_n1037(eclk, ereset, n1037_i0,n1037_i1,n1037_i2, n1037_v);
  spice_node_2 n_C56(eclk, ereset, C56_i0,C56_i1, C56_v);
  spice_node_1 n_n402(eclk, ereset, n402_i0, n402_v);
  spice_node_2 n_n630(eclk, ereset, n630_i0,n630_i1, n630_v);
  spice_node_2 n_n631(eclk, ereset, n631_i2,n631_i3, n631_v);
  spice_node_2 n_op_T5_ind_x(eclk, ereset, op_T5_ind_x_i0,op_T5_ind_x_i2, op_T5_ind_x_v);
  spice_node_3 n_n1211(eclk, ereset, n1211_i0,n1211_i2,n1211_i4, n1211_v);
  spice_node_2 n_n634(eclk, ereset, n634_i0,n634_i1, n634_v);
  spice_node_2 n___AxB7__C67(eclk, ereset, __AxB7__C67_i0,__AxB7__C67_i1, __AxB7__C67_v);
  spice_node_2 n_n1214(eclk, ereset, n1214_i0,n1214_i1, n1214_v);
  spice_node_2 n_n637(eclk, ereset, n637_i0,n637_i1, n637_v);
  spice_node_2 n_n638(eclk, ereset, n638_i0,n638_i1, n638_v);
  spice_node_2 n_ADL_ABL(eclk, ereset, ADL_ABL_i0,ADL_ABL_i1, ADL_ABL_v);
  spice_node_2 n_n1218(eclk, ereset, n1218_i0,n1218_i1, n1218_v);
  spice_node_3 n_n1376(eclk, ereset, n1376_i0,n1376_i1,n1376_i2, n1376_v);
  spice_node_3 n_n465(eclk, ereset, n465_i0,n465_i1,n465_i2, n465_v);
  spice_node_2 n_n1107(eclk, ereset, n1107_i1,n1107_i2, n1107_v);
  spice_node_1 n_pipeUNK42(eclk, ereset, pipeUNK42_i0, pipeUNK42_v);
  spice_node_2 n_n1105(eclk, ereset, n1105_i0,n1105_i2, n1105_v);
  spice_node_1 n_n1450(eclk, ereset, n1450_i0, n1450_v);
  spice_node_1 n_n1452(eclk, ereset, n1452_i1, n1452_v);
  spice_node_2 n_dor5(eclk, ereset, dor5_i1,dor5_i2, dor5_v);
  spice_node_5 n_n1458(eclk, ereset, n1458_i0,n1458_i1,n1458_i2,n1458_i3,n1458_i4, n1458_v);
  spice_node_3 n___AxB_6(eclk, ereset, __AxB_6_i1,__AxB_6_i2,__AxB_6_i4, __AxB_6_v);
  spice_node_8 n_idb0(eclk, ereset, idb0_i1,idb0_i2,idb0_i4,idb0_i5,idb0_i6,idb0_i7,idb0_i8,idb0_i10, idb0_v);
  spice_node_2 n_n1109(eclk, ereset, n1109_i0,n1109_i3, n1109_v);
  spice_node_5 n_n1722(eclk, ereset, n1722_i0,n1722_i1,n1722_i2,n1722_i3,n1722_i4, n1722_v);
  spice_node_2 n_DA_AB2(eclk, ereset, DA_AB2_i0,DA_AB2_i1, DA_AB2_v);
  spice_node_2 n_n_0_ADL0(eclk, ereset, n_0_ADL0_i0,n_0_ADL0_i2, n_0_ADL0_v);
  spice_node_2 n_dpc19_ADDSB7(eclk, ereset, dpc19_ADDSB7_i0,dpc19_ADDSB7_i2, dpc19_ADDSB7_v);
  spice_node_1 n_pipeUNK10(eclk, ereset, pipeUNK10_i0, pipeUNK10_v);
  spice_node_3 n_n212(eclk, ereset, n212_i0,n212_i1,n212_i2, n212_v);
  spice_node_3 n_n213(eclk, ereset, n213_i0,n213_i1,n213_i2, n213_v);
  spice_node_3 n_n210(eclk, ereset, n210_i0,n210_i1,n210_i3, n210_v);
  spice_node_3 n_ab3(eclk, ereset, ab3_i0,ab3_i1,ab3_i2, ab3_v);
  spice_node_2 n_n218(eclk, ereset, n218_i0,n218_i1, n218_v);
  spice_node_2 n_op_T2_mem_zp(eclk, ereset, op_T2_mem_zp_i0,op_T2_mem_zp_i2, op_T2_mem_zp_v);
  spice_node_2 n_op_T0_tay(eclk, ereset, op_T0_tay_i0,op_T0_tay_i1, op_T0_tay_v);
  spice_node_2 n_n919(eclk, ereset, n919_i0,n919_i3, n919_v);
  spice_node_2 n_n918(eclk, ereset, n918_i0,n918_i1, n918_v);
  spice_node_2 n_n917(eclk, ereset, n917_i0,n917_i2, n917_v);
  spice_node_3 n_n916(eclk, ereset, n916_i0,n916_i1,n916_i3, n916_v);
  spice_node_2 n_alucin(eclk, ereset, alucin_i1,alucin_i2, alucin_v);
  spice_node_3 n_n913(eclk, ereset, n913_i0,n913_i1,n913_i2, n913_v);
  spice_node_2 n_n847(eclk, ereset, n847_i0,n847_i1, n847_v);
  spice_node_2 n_n846(eclk, ereset, n846_i0,n846_i1, n846_v);
  spice_node_3 n_n845(eclk, ereset, n845_i0,n845_i1,n845_i2, n845_v);
  spice_node_3 n_n844(eclk, ereset, n844_i0,n844_i1,n844_i2, n844_v);
  spice_node_2 n_y7(eclk, ereset, y7_i0,y7_i1, y7_v);
  spice_node_2 n_n842(eclk, ereset, n842_i0,n842_i3, n842_v);
  spice_node_4 n_aluanandb1(eclk, ereset, aluanandb1_i0,aluanandb1_i1,aluanandb1_i3,aluanandb1_i4, aluanandb1_v);
  spice_node_2 n__op_branch_bit6(eclk, ereset, _op_branch_bit6_i0,_op_branch_bit6_i2, _op_branch_bit6_v);
  spice_node_2 n_n849(eclk, ereset, n849_i0,n849_i2, n849_v);
  spice_node_1 n_pipeUNK33(eclk, ereset, pipeUNK33_i0, pipeUNK33_v);
  spice_node_1 n_n663(eclk, ereset, n663_i0, n663_v);
  spice_node_2 n_pd3_clearIR(eclk, ereset, pd3_clearIR_i1,pd3_clearIR_i3, pd3_clearIR_v);
  spice_node_2 n_n662(eclk, ereset, n662_i0,n662_i1, n662_v);
  spice_node_3 n_n1039(eclk, ereset, n1039_i0,n1039_i1,n1039_i2, n1039_v);
  spice_node_2 n_n753(eclk, ereset, n753_i0,n753_i1, n753_v);
  spice_node_1 n_nots2(eclk, ereset, nots2_i1, nots2_v);
  spice_node_1 n_pchp6(eclk, ereset, pchp6_i1, pchp6_v);
  spice_node_2 n_op_T2_php(eclk, ereset, op_T2_php_i0,op_T2_php_i1, op_T2_php_v);
  spice_node_2 n_n757(eclk, ereset, n757_i0,n757_i1, n757_v);
  spice_node_1 n_n756(eclk, ereset, n756_i0, n756_v);
  spice_node_2 n_n755(eclk, ereset, n755_i0,n755_i1, n755_v);
  spice_node_2 n_n754(eclk, ereset, n754_i1,n754_i3, n754_v);
  spice_node_1 n_n759(eclk, ereset, n759_i0, n759_v);
  spice_node_1 n_pd0(eclk, ereset, pd0_i0, pd0_v);
  spice_node_2 n_n1595(eclk, ereset, n1595_i0,n1595_i1, n1595_v);
  spice_node_3 n_n506(eclk, ereset, n506_i0,n506_i1,n506_i3, n506_v);
  spice_node_3 n_idl0(eclk, ereset, idl0_i0,idl0_i1,idl0_i2, idl0_v);
  spice_node_2 n_n1596(eclk, ereset, n1596_i0,n1596_i3, n1596_v);
  spice_node_3 n_db6(eclk, ereset, db6_i0,db6_i3,db6_i4, db6_v);
  spice_node_2 n_n1593(eclk, ereset, n1593_i2,n1593_i3, n1593_v);
  spice_node_2 n_n1033(eclk, ereset, n1033_i0,n1033_i2, n1033_v);
  spice_node_2 n_n1599(eclk, ereset, n1599_i1,n1599_i2, n1599_v);
  spice_node_2 n_n1025(eclk, ereset, n1025_i1,n1025_i2, n1025_v);
  spice_node_3 n_n1024(eclk, ereset, n1024_i0,n1024_i1,n1024_i2, n1024_v);
  spice_node_1 n_n1027(eclk, ereset, n1027_i0, n1027_v);
  spice_node_2 n_C12(eclk, ereset, C12_i0,C12_i1, C12_v);
  spice_node_2 n_aluaorb1(eclk, ereset, aluaorb1_i0,aluaorb1_i1, aluaorb1_v);
  spice_node_1 n_n1020(eclk, ereset, n1020_i1, n1020_v);
  spice_node_2 n_C23(eclk, ereset, C23_i1,C23_i2, C23_v);
  spice_node_2 n_pcl1(eclk, ereset, pcl1_i1,pcl1_i2, pcl1_v);
  spice_node_1 n_pipephi2Reset0x(eclk, ereset, pipephi2Reset0x_i0, pipephi2Reset0x_v);
  spice_node_1 n_nots6(eclk, ereset, nots6_i0, nots6_v);
  spice_node_2 n_n1028(eclk, ereset, n1028_i0,n1028_i2, n1028_v);
  spice_node_2 n_n503(eclk, ereset, n503_i0,n503_i2, n503_v);
  spice_node_2 n_n1034(eclk, ereset, n1034_i0,n1034_i3, n1034_v);
  spice_node_3 n_n501(eclk, ereset, n501_i0,n501_i1,n501_i2, n501_v);
  spice_node_2 n_s6(eclk, ereset, s6_i0,s6_i1, s6_v);
  spice_node_2 n_op_T3_mem_abs(eclk, ereset, op_T3_mem_abs_i0,op_T3_mem_abs_i2, op_T3_mem_abs_v);
  spice_node_4 n_alu4(eclk, ereset, alu4_i0,alu4_i1,alu4_i2,alu4_i3, alu4_v);
  spice_node_1 n_nots5(eclk, ereset, nots5_i1, nots5_v);
  spice_node_2 n_n600(eclk, ereset, n600_i0,n600_i1, n600_v);
  spice_node_2 n_n603(eclk, ereset, n603_i0,n603_i1, n603_v);
  spice_node_2 n_n1213(eclk, ereset, n1213_i0,n1213_i1, n1213_v);
  spice_node_2 n_n1205(eclk, ereset, n1205_i0,n1205_i2, n1205_v);
  spice_node_2 n_op_T2_ind_y(eclk, ereset, op_T2_ind_y_i0,op_T2_ind_y_i1, op_T2_ind_y_v);
  spice_node_5 n_n1206(eclk, ereset, n1206_i0,n1206_i1,n1206_i2,n1206_i3,n1206_i4, n1206_v);
  spice_node_2 n_n609(eclk, ereset, n609_i0,n609_i2, n609_v);
  spice_node_3 n_n608(eclk, ereset, n608_i0,n608_i1,n608_i2, n608_v);
  spice_node_2 n_n1202(eclk, ereset, n1202_i0,n1202_i1, n1202_v);
  spice_node_2 n_n1560(eclk, ereset, n1560_i1,n1560_i2, n1560_v);
  spice_node_2 n_x0(eclk, ereset, x0_i0,x0_i1, x0_v);
  spice_node_3 n_n635(eclk, ereset, n635_i0,n635_i1,n635_i3, n635_v);
  spice_node_2 n_n636(eclk, ereset, n636_i0,n636_i2, n636_v);
  spice_node_4 n_n1215(eclk, ereset, n1215_i0,n1215_i1,n1215_i2,n1215_i3, n1215_v);
  spice_node_1 n_n1447(eclk, ereset, n1447_i0, n1447_v);
  spice_node_2 n_n1446(eclk, ereset, n1446_i1,n1446_i2, n1446_v);
  spice_node_2 n_ir4(eclk, ereset, ir4_i0,ir4_i2, ir4_v);
  spice_node_3 n_ab10(eclk, ereset, ab10_i0,ab10_i1,ab10_i2, ab10_v);
  spice_node_1 n_pipeUNK13(eclk, ereset, pipeUNK13_i0, pipeUNK13_v);
  spice_node_3 n_n1117(eclk, ereset, n1117_i0,n1117_i1,n1117_i2, n1117_v);
  spice_node_3 n_idl6(eclk, ereset, idl6_i0,idl6_i1,idl6_i2, idl6_v);
  spice_node_3 n_Pout4(eclk, ereset, Pout4_i0,Pout4_i1,Pout4_i2, Pout4_v);
  spice_node_2 n_n1449(eclk, ereset, n1449_i0,n1449_i1, n1449_v);
  spice_node_2 n_n1448(eclk, ereset, n1448_i0,n1448_i1, n1448_v);
  spice_node_2 n_n1219(eclk, ereset, n1219_i1,n1219_i2, n1219_v);
  spice_node_2 n_x_op_T4_ind_y(eclk, ereset, x_op_T4_ind_y_i0,x_op_T4_ind_y_i3, x_op_T4_ind_y_v);
  spice_node_1 n_n460(eclk, ereset, n460_i0, n460_v);
  spice_node_2 n_abh7(eclk, ereset, abh7_i0,abh7_i4, abh7_v);
  spice_node_5 n_n488(eclk, ereset, n488_i0,n488_i1,n488_i2,n488_i3,n488_i4, n488_v);
  spice_node_2 n_op_T2_brk(eclk, ereset, op_T2_brk_i0,op_T2_brk_i1, op_T2_brk_v);
  spice_node_3 n___AxBxC_5(eclk, ereset, __AxBxC_5_i0,__AxBxC_5_i1,__AxBxC_5_i2, __AxBxC_5_v);
  spice_node_2 n_n485(eclk, ereset, n485_i1,n485_i2, n485_v);
  spice_node_3 n_n484(eclk, ereset, n484_i0,n484_i1,n484_i2, n484_v);
  spice_node_6 n_adh5(eclk, ereset, adh5_i0,adh5_i1,adh5_i2,adh5_i3,adh5_i4,adh5_i5, adh5_v);
  spice_node_5 n_n481(eclk, ereset, n481_i0,n481_i1,n481_i2,n481_i3,n481_i4, n481_v);
  spice_node_2 n_n480(eclk, ereset, n480_i0,n480_i1, n480_v);
  spice_node_1 n_pipeUNK09(eclk, ereset, pipeUNK09_i0, pipeUNK09_v);
  spice_node_2 n_n198(eclk, ereset, n198_i2,n198_i3, n198_v);
  spice_node_3 n_ab15(eclk, ereset, ab15_i0,ab15_i1,ab15_i2, ab15_v);
  spice_node_3 n_notir0(eclk, ereset, notir0_i0,notir0_i1,notir0_i2, notir0_v);
  spice_node_1 n_pipeUNK37(eclk, ereset, pipeUNK37_i0, pipeUNK37_v);
  spice_node_2 n_n196(eclk, ereset, n196_i0,n196_i2, n196_v);
  spice_node_3 n_n191(eclk, ereset, n191_i0,n191_i1,n191_i2, n191_v);
  spice_node_1 n_n190(eclk, ereset, n190_i1, n190_v);
  spice_node_2 n__AxB_2__C12(eclk, ereset, _AxB_2__C12_i0,_AxB_2__C12_i1, _AxB_2__C12_v);
  spice_node_2 n_n192(eclk, ereset, n192_i0,n192_i4, n192_v);
  spice_node_3 n_n1106(eclk, ereset, n1106_i0,n1106_i1,n1106_i2, n1106_v);
  spice_node_3 n_n1455(eclk, ereset, n1455_i1,n1455_i2,n1455_i3, n1455_v);
  spice_node_1 n_n1274(eclk, ereset, n1274_i0, n1274_v);
  spice_node_2 n_n1457(eclk, ereset, n1457_i0,n1457_i1, n1457_v);
  spice_node_1 n_pclp1(eclk, ereset, pclp1_i0, pclp1_v);
  spice_node_3 n_n1100(eclk, ereset, n1100_i0,n1100_i2,n1100_i3, n1100_v);
  spice_node_3 n_n1101(eclk, ereset, n1101_i0,n1101_i1,n1101_i2, n1101_v);
  spice_node_1 n_n902(eclk, ereset, n902_i0, n902_v);
  spice_node_2 n_pcl4(eclk, ereset, pcl4_i1,pcl4_i2, pcl4_v);
  spice_node_2 n__DA_ADD1(eclk, ereset, _DA_ADD1_i0,_DA_ADD1_i2, _DA_ADD1_v);
  spice_node_2 n_n906(eclk, ereset, n906_i0,n906_i3, n906_v);
  spice_node_2 n__ABH1(eclk, ereset, _ABH1_i0,_ABH1_i2, _ABH1_v);
  spice_node_2 n_op_T3_mem_zp_idx(eclk, ereset, op_T3_mem_zp_idx_i0,op_T3_mem_zp_idx_i2, op_T3_mem_zp_idx_v);
  spice_node_2 n_n905(eclk, ereset, n905_i1,n905_i2, n905_v);
  spice_node_3 n_n420(eclk, ereset, n420_i0,n420_i1,n420_i2, n420_v);
  spice_node_2 n_t5(eclk, ereset, t5_i0,t5_i1, t5_v);
  spice_node_3 n_n854(eclk, ereset, n854_i0,n854_i1,n854_i3, n854_v);
  spice_node_2 n_n855(eclk, ereset, n855_i0,n855_i2, n855_v);
  spice_node_2 n_op_rti_rts(eclk, ereset, op_rti_rts_i1,op_rti_rts_i3, op_rti_rts_v);
  spice_node_2 n_n850(eclk, ereset, n850_i0,n850_i2, n850_v);
  spice_node_2 n_abh3(eclk, ereset, abh3_i3,abh3_i4, abh3_v);
  spice_node_2 n_n852(eclk, ereset, n852_i0,n852_i1, n852_v);
  spice_node_2 n_op_T5_rts(eclk, ereset, op_T5_rts_i0,op_T5_rts_i2, op_T5_rts_v);
  spice_node_2 n_a5(eclk, ereset, a5_i0,a5_i2, a5_v);
  spice_node_2 n_dpc9_DBADD(eclk, ereset, dpc9_DBADD_i1,dpc9_DBADD_i9, dpc9_DBADD_v);
  spice_node_2 n_n6(eclk, ereset, n6_i2,n6_i3, n6_v);
  spice_node_2 n_AxB1(eclk, ereset, AxB1_i1,AxB1_i3, AxB1_v);
  spice_node_2 n_n611(eclk, ereset, n611_i2,n611_i3, n611_v);
  spice_node_6 n_n740(eclk, ereset, n740_i0,n740_i1,n740_i2,n740_i3,n740_i4,n740_i5, n740_v);
  spice_node_2 n_dpc31_PCHPCH(eclk, ereset, dpc31_PCHPCH_i8,dpc31_PCHPCH_i9, dpc31_PCHPCH_v);
  spice_node_2 n_n743(eclk, ereset, n743_i0,n743_i1, n743_v);
  spice_node_2 n_DBZ(eclk, ereset, DBZ_i1,DBZ_i2, DBZ_v);
  spice_node_1 n_n745(eclk, ereset, n745_i0, n745_v);
  spice_node_2 n_dor1(eclk, ereset, dor1_i0,dor1_i2, dor1_v);
  spice_node_2 n_n747(eclk, ereset, n747_i0,n747_i3, n747_v);
  spice_node_2 n_n748(eclk, ereset, n748_i0,n748_i1, n748_v);
  spice_node_2 n_n617(eclk, ereset, n617_i0,n617_i3, n617_v);
  spice_node_2 n_x_op_push_pull(eclk, ereset, x_op_push_pull_i0,x_op_push_pull_i1, x_op_push_pull_v);
  spice_node_1 n_pipeUNK16(eclk, ereset, pipeUNK16_i0, pipeUNK16_v);
  spice_node_2 n_x_op_jmp(eclk, ereset, x_op_jmp_i0,x_op_jmp_i3, x_op_jmp_v);
  spice_node_2 n_n1054(eclk, ereset, n1054_i0,n1054_i1, n1054_v);
  spice_node_2 n_n1055(eclk, ereset, n1055_i0,n1055_i1, n1055_v);
  spice_node_2 n_n1056(eclk, ereset, n1056_i0,n1056_i1, n1056_v);
  spice_node_2 n_op_T2_abs(eclk, ereset, op_T2_abs_i0,op_T2_abs_i1, op_T2_abs_v);
  spice_node_1 n_n1059(eclk, ereset, n1059_i0, n1059_v);
  spice_node_2 n_n1696(eclk, ereset, n1696_i0,n1696_i1, n1696_v);
  spice_node_2 n_n1697(eclk, ereset, n1697_i0,n1697_i1, n1697_v);
  spice_node_4 n_n1694(eclk, ereset, n1694_i0,n1694_i1,n1694_i2,n1694_i3, n1694_v);
  spice_node_1 n_n1693(eclk, ereset, n1693_i0, n1693_v);
  spice_node_1 n_pd7(eclk, ereset, pd7_i0, pd7_v);
  spice_node_3 n_n1691(eclk, ereset, n1691_i0,n1691_i2,n1691_i3, n1691_v);
  spice_node_2 n_dpc24_ACSB(eclk, ereset, dpc24_ACSB_i0,dpc24_ACSB_i9, dpc24_ACSB_v);
  spice_node_1 n_n1699(eclk, ereset, n1699_i1, n1699_v);
  spice_node_5 n_n618(eclk, ereset, n618_i0,n618_i1,n618_i2,n618_i3,n618_i4, n618_v);
  spice_node_2 n_n612(eclk, ereset, n612_i0,n612_i2, n612_v);
  spice_node_2 n_n613(eclk, ereset, n613_i0,n613_i3, n613_v);
  spice_node_1 n_n1272(eclk, ereset, n1272_i1, n1272_v);
  spice_node_2 n_op_T0(eclk, ereset, op_T0_i1,op_T0_i2, op_T0_v);
  spice_node_3 n_n616(eclk, ereset, n616_i0,n616_i1,n616_i2, n616_v);
  spice_node_3 n_n1275(eclk, ereset, n1275_i0,n1275_i1,n1275_i2, n1275_v);
  spice_node_1 n_pipeUNK31(eclk, ereset, pipeUNK31_i0, pipeUNK31_v);
  spice_node_2 n_y5(eclk, ereset, y5_i0,y5_i1, y5_v);
  spice_node_1 n_n1472(eclk, ereset, n1472_i0, n1472_v);
  spice_node_8 n_idb2(eclk, ereset, idb2_i0,idb2_i1,idb2_i3,idb2_i4,idb2_i5,idb2_i6,idb2_i8,idb2_i9, idb2_v);
  spice_node_2 n_n1471(eclk, ereset, n1471_i1,n1471_i2, n1471_v);
  spice_node_2 n_x_op_T0_bit(eclk, ereset, x_op_T0_bit_i1,x_op_T0_bit_i2, x_op_T0_bit_v);
  spice_node_1 n_n1477(eclk, ereset, n1477_i0, n1477_v);
  spice_node_3 n_n1474(eclk, ereset, n1474_i0,n1474_i1,n1474_i2, n1474_v);
  spice_node_3 n_dasb3(eclk, ereset, dasb3_i0,dasb3_i1,dasb3_i2, dasb3_v);
  spice_node_2 n_op_T0_brk_rti(eclk, ereset, op_T0_brk_rti_i0,op_T0_brk_rti_i1, op_T0_brk_rti_v);
  spice_node_2 n_n1479(eclk, ereset, n1479_i0,n1479_i1, n1479_v);
  spice_node_2 n_n1304(eclk, ereset, n1304_i1,n1304_i2, n1304_v);
  spice_node_2 n_n1305(eclk, ereset, n1305_i1,n1305_i2, n1305_v);
  spice_node_3 n_idl4(eclk, ereset, idl4_i0,idl4_i1,idl4_i2, idl4_v);
  spice_node_2 n__ABL6(eclk, ereset, _ABL6_i1,_ABL6_i2, _ABL6_v);
  spice_node_2 n_n1300(eclk, ereset, n1300_i1,n1300_i2, n1300_v);
  spice_node_5 n_n1301(eclk, ereset, n1301_i0,n1301_i1,n1301_i2,n1301_i3,n1301_i4, n1301_v);
  spice_node_8 n_idb3(eclk, ereset, idb3_i0,idb3_i1,idb3_i3,idb3_i5,idb3_i6,idb3_i8,idb3_i9,idb3_i10, idb3_v);
  spice_node_2 n_n1303(eclk, ereset, n1303_i0,n1303_i2, n1303_v);
  spice_node_3 n_notaluvout(eclk, ereset, notaluvout_i0,notaluvout_i1,notaluvout_i2, notaluvout_v);
  spice_node_3 n_n1309(eclk, ereset, n1309_i0,n1309_i1,n1309_i2, n1309_v);
  spice_node_1 n_notidl5(eclk, ereset, notidl5_i0, notidl5_v);
  spice_node_2 n_n499(eclk, ereset, n499_i0,n499_i1, n499_v);
  spice_node_3 n_n494(eclk, ereset, n494_i0,n494_i1,n494_i2, n494_v);
  spice_node_1 n_notalu3(eclk, ereset, notalu3_i0, notalu3_v);
  spice_node_3 n_n496(eclk, ereset, n496_i0,n496_i1,n496_i2, n496_v);
  spice_node_3 n_n490(eclk, ereset, n490_i0,n490_i1,n490_i2, n490_v);
  spice_node_2 n_n491(eclk, ereset, n491_i0,n491_i1, n491_v);
  spice_node_2 n_op_T4_ind_y(eclk, ereset, op_T4_ind_y_i0,op_T4_ind_y_i1, op_T4_ind_y_v);
  spice_node_8 n_idb7(eclk, ereset, idb7_i0,idb7_i2,idb7_i3,idb7_i4,idb7_i6,idb7_i7,idb7_i8,idb7_i9, idb7_v);
  spice_node_1 n_n24(eclk, ereset, n24_i0, n24_v);
  spice_node_2 n_n25(eclk, ereset, n25_i1,n25_i2, n25_v);
  spice_node_3 n_notir4(eclk, ereset, notir4_i0,notir4_i1,notir4_i2, notir4_v);
  spice_node_5 n_n27(eclk, ereset, n27_i0,n27_i1,n27_i2,n27_i3,n27_i4, n27_v);
  spice_node_3 n_n20(eclk, ereset, n20_i0,n20_i1,n20_i2, n20_v);
  spice_node_2 n_n21(eclk, ereset, n21_i2,n21_i3, n21_v);
  spice_node_3 n___AxBxC_2(eclk, ereset, __AxBxC_2_i0,__AxBxC_2_i1,__AxBxC_2_i2, __AxBxC_2_v);
  spice_node_2 n_n23(eclk, ereset, n23_i1,n23_i2, n23_v);
  spice_node_2 n__ABL7(eclk, ereset, _ABL7_i1,_ABL7_i2, _ABL7_v);
  spice_node_3 n_n29(eclk, ereset, n29_i0,n29_i1,n29_i2, n29_v);
  spice_node_2 n_n7(eclk, ereset, n7_i0,n7_i2, n7_v);
  spice_node_2 n_n410(eclk, ereset, n410_i0,n410_i1, n410_v);
  spice_node_1 n_n590(eclk, ereset, n590_i0, n590_v);
  spice_node_3 n_n1085(eclk, ereset, n1085_i0,n1085_i1,n1085_i2, n1085_v);
  spice_node_2 n__C67(eclk, ereset, _C67_i0,_C67_i1, _C67_v);
  spice_node_3 n_n1083(eclk, ereset, n1083_i0,n1083_i1,n1083_i4, n1083_v);
  spice_node_2 n_op_T0_jmp(eclk, ereset, op_T0_jmp_i0,op_T0_jmp_i1, op_T0_jmp_v);
  spice_node_3 n_alub0(eclk, ereset, alub0_i0,alub0_i1,alub0_i2, alub0_v);
  spice_node_5 n_n976(eclk, ereset, n976_i0,n976_i1,n976_i2,n976_i3,n976_i4, n976_v);
  spice_node_2 n_n975(eclk, ereset, n975_i0,n975_i1, n975_v);
  spice_node_1 n_pipeUNK02(eclk, ereset, pipeUNK02_i1, pipeUNK02_v);
  spice_node_3 n_n973(eclk, ereset, n973_i0,n973_i1,n973_i2, n973_v);
  spice_node_2 n_t2(eclk, ereset, t2_i0,t2_i2, t2_v);
  spice_node_1 n_pipeUNK23(eclk, ereset, pipeUNK23_i0, pipeUNK23_v);
  spice_node_2 n_n979(eclk, ereset, n979_i0,n979_i1, n979_v);
  spice_node_2 n_a2(eclk, ereset, a2_i1,a2_i2, a2_v);
  spice_node_3 n_n182(eclk, ereset, n182_i1,n182_i2,n182_i4, n182_v);
  spice_node_2 n_s1(eclk, ereset, s1_i0,s1_i1, s1_v);
  spice_node_2 n_n180(eclk, ereset, n180_i0,n180_i1, n180_v);
  spice_node_1 n_nots7(eclk, ereset, nots7_i1, nots7_v);
  spice_node_5 n_notRnWprepad(eclk, ereset, notRnWprepad_i0,notRnWprepad_i1,notRnWprepad_i2,notRnWprepad_i3,notRnWprepad_i4, notRnWprepad_v);
  spice_node_2 n_n184(eclk, ereset, n184_i0,n184_i2, n184_v);
  spice_node_3 n_n188(eclk, ereset, n188_i0,n188_i2,n188_i3, n188_v);
  spice_node_2 n_n1464(eclk, ereset, n1464_i0,n1464_i2, n1464_v);
  spice_node_3 n_n869(eclk, ereset, n869_i1,n869_i2,n869_i3, n869_v);
  spice_node_1 n_pclp3(eclk, ereset, pclp3_i1, pclp3_v);
  spice_node_2 n_n861(eclk, ereset, n861_i0,n861_i1, n861_v);
  spice_node_2 n___AxB3__C23(eclk, ereset, __AxB3__C23_i0,__AxB3__C23_i1, __AxB3__C23_v);
  spice_node_2 n_dpc43_DL_DB(eclk, ereset, dpc43_DL_DB_i0,dpc43_DL_DB_i9, dpc43_DL_DB_v);
  spice_node_4 n_n862(eclk, ereset, n862_i0,n862_i1,n862_i3,n862_i4, n862_v);
  spice_node_1 n_n865(eclk, ereset, n865_i0, n865_v);
  spice_node_2 n_n867(eclk, ereset, n867_i1,n867_i2, n867_v);
  spice_node_0 n_n866(eclk, ereset,  n866_v);
  spice_node_3 n_n883(eclk, ereset, n883_i0,n883_i1,n883_i2, n883_v);
  spice_node_2 n_n882(eclk, ereset, n882_i0,n882_i1, n882_v);
  spice_node_3 n_n880(eclk, ereset, n880_i0,n880_i1,n880_i2, n880_v);
  spice_node_3 n_ab6(eclk, ereset, ab6_i0,ab6_i1,ab6_i2, ab6_v);
  spice_node_2 n_n885(eclk, ereset, n885_i0,n885_i1, n885_v);
  spice_node_3 n_n884(eclk, ereset, n884_i0,n884_i1,n884_i2, n884_v);
  spice_node_3 n_n889(eclk, ereset, n889_i0,n889_i1,n889_i2, n889_v);
  spice_node_2 n_n888(eclk, ereset, n888_i0,n888_i1, n888_v);
  spice_node_2 n_abh5(eclk, ereset, abh5_i3,abh5_i4, abh5_v);
  spice_node_3 n_n774(eclk, ereset, n774_i0,n774_i1,n774_i2, n774_v);
  spice_node_2 n_x7(eclk, ereset, x7_i1,x7_i2, x7_v);
  spice_node_2 n_op_T5_jsr(eclk, ereset, op_T5_jsr_i1,op_T5_jsr_i2, op_T5_jsr_v);
  spice_node_2 n_n771(eclk, ereset, n771_i0,n771_i2, n771_v);
  spice_node_2 n_n770(eclk, ereset, n770_i0,n770_i2, n770_v);
  spice_node_2 n_n773(eclk, ereset, n773_i0,n773_i1, n773_v);
  spice_node_2 n_n772(eclk, ereset, n772_i2,n772_i3, n772_v);
  spice_node_3 n_n779(eclk, ereset, n779_i0,n779_i1,n779_i2, n779_v);
  spice_node_2 n_ONEBYTE(eclk, ereset, ONEBYTE_i0,ONEBYTE_i1, ONEBYTE_v);
  spice_node_2 n_n419(eclk, ereset, n419_i0,n419_i2, n419_v);
  spice_node_3 n_Pout6(eclk, ereset, Pout6_i0,Pout6_i1,Pout6_i2, Pout6_v);
  spice_node_2 n_op_T0_dex(eclk, ereset, op_T0_dex_i0,op_T0_dex_i1, op_T0_dex_v);
  spice_node_2 n_n75(eclk, ereset, n75_i0,n75_i2, n75_v);
  spice_node_1 n_pipeUNK27(eclk, ereset, pipeUNK27_i1, pipeUNK27_v);
  spice_node_5 n_n72(eclk, ereset, n72_i0,n72_i1,n72_i2,n72_i3,n72_i4, n72_v);
  spice_node_2 n_n71(eclk, ereset, n71_i0,n71_i1, n71_v);
  spice_node_2 n_n70(eclk, ereset, n70_i1,n70_i2, n70_v);
  spice_node_2 n_n79(eclk, ereset, n79_i0,n79_i1, n79_v);
  spice_node_2 n_C34(eclk, ereset, C34_i0,C34_i1, C34_v);
  spice_node_2 n_n1043(eclk, ereset, n1043_i0,n1043_i1, n1043_v);
  spice_node_2 n_H1x1(eclk, ereset, H1x1_i4,H1x1_i8, H1x1_v);
  spice_node_2 n_n1041(eclk, ereset, n1041_i0,n1041_i1, n1041_v);
  spice_node_2 n_n1047(eclk, ereset, n1047_i0,n1047_i1, n1047_v);
  spice_node_3 n_n1046(eclk, ereset, n1046_i0,n1046_i1,n1046_i2, n1046_v);
  spice_node_3 n_n1045(eclk, ereset, n1045_i1,n1045_i2,n1045_i3, n1045_v);
  spice_node_2 n_n1044(eclk, ereset, n1044_i0,n1044_i1, n1044_v);
  spice_node_1 n_n1049(eclk, ereset, n1049_i0, n1049_v);
  spice_node_2 n__op_branch_done(eclk, ereset, _op_branch_done_i0,_op_branch_done_i1, _op_branch_done_v);
  spice_node_2 n_alua3(eclk, ereset, alua3_i0,alua3_i1, alua3_v);
  spice_node_1 n_n1683(eclk, ereset, n1683_i0, n1683_v);
  spice_node_2 n_n1682(eclk, ereset, n1682_i0,n1682_i1, n1682_v);
  spice_node_3 n_n1684(eclk, ereset, n1684_i0,n1684_i1,n1684_i2, n1684_v);
  spice_node_3 n_n1687(eclk, ereset, n1687_i0,n1687_i1,n1687_i2, n1687_v);
  spice_node_3 n_op_EORS(eclk, ereset, op_EORS_i0,op_EORS_i1,op_EORS_i2, op_EORS_v);
  spice_node_3 n_n1688(eclk, ereset, n1688_i0,n1688_i1,n1688_i2, n1688_v);
  spice_node_1 n_n1269(eclk, ereset, n1269_i1, n1269_v);
  spice_node_2 n__DBZ(eclk, ereset, _DBZ_i0,_DBZ_i1, _DBZ_v);
  spice_node_2 n_n669(eclk, ereset, n669_i1,n669_i2, n669_v);
  spice_node_2 n__ABH4(eclk, ereset, _ABH4_i1,_ABH4_i2, _ABH4_v);
  spice_node_2 n_pd5_clearIR(eclk, ereset, pd5_clearIR_i1,pd5_clearIR_i2, pd5_clearIR_v);
  spice_node_2 n_n1262(eclk, ereset, n1262_i0,n1262_i1, n1262_v);
  spice_node_2 n_op_T0_ldy_mem(eclk, ereset, op_T0_ldy_mem_i0,op_T0_ldy_mem_i1, op_T0_ldy_mem_v);
  spice_node_2 n_n664(eclk, ereset, n664_i1,n664_i2, n664_v);
  spice_node_3 n_n1267(eclk, ereset, n1267_i0,n1267_i1,n1267_i2, n1267_v);
  spice_node_1 n_notdor5(eclk, ereset, notdor5_i0, notdor5_v);
  spice_node_2 n_op_T3_branch(eclk, ereset, op_T3_branch_i1,op_T3_branch_i3, op_T3_branch_v);
  spice_node_3 n_clk2out(eclk, ereset, clk2out_i0,clk2out_i1,clk2out_i2, clk2out_v);
  spice_node_3 n_n1469(eclk, ereset, n1469_i0,n1469_i1,n1469_i2, n1469_v);
  spice_node_2 n_dpc5_SADL(eclk, ereset, dpc5_SADL_i0,dpc5_SADL_i7, dpc5_SADL_v);
  spice_node_3 n_VEC0(eclk, ereset, VEC0_i1,VEC0_i2,VEC0_i4, VEC0_v);
  spice_node_2 n_n1018(eclk, ereset, n1018_i0,n1018_i1, n1018_v);
  spice_node_2 n_n1467(eclk, ereset, n1467_i0,n1467_i1, n1467_v);
  spice_node_2 n_op_rol_ror(eclk, ereset, op_rol_ror_i0,op_rol_ror_i1, op_rol_ror_v);
  spice_node_2 n_pd6_clearIR(eclk, ereset, pd6_clearIR_i1,pd6_clearIR_i2, pd6_clearIR_v);
  spice_node_2 n_n1463(eclk, ereset, n1463_i1,n1463_i2, n1463_v);
  spice_node_2 n_PD_xxxx10x0(eclk, ereset, PD_xxxx10x0_i1,PD_xxxx10x0_i2, PD_xxxx10x0_v);
  spice_node_2 n_n1316(eclk, ereset, n1316_i0,n1316_i1, n1316_v);
  spice_node_2 n_n1315(eclk, ereset, n1315_i0,n1315_i3, n1315_v);
  spice_node_2 n_C67(eclk, ereset, C67_i1,C67_i5, C67_v);
  spice_node_2 n_A_B3(eclk, ereset, A_B3_i0,A_B3_i1, A_B3_v);
  spice_node_2 n_n1312(eclk, ereset, n1312_i0,n1312_i2, n1312_v);
  spice_node_2 n_op_T4_rti(eclk, ereset, op_T4_rti_i0,op_T4_rti_i1, op_T4_rti_v);
  spice_node_3 n_n1319(eclk, ereset, n1319_i0,n1319_i1,n1319_i2, n1319_v);
  spice_node_4 n_n1318(eclk, ereset, n1318_i1,n1318_i2,n1318_i3,n1318_i5, n1318_v);
  spice_node_2 n_xx_op_T5_jsr(eclk, ereset, xx_op_T5_jsr_i0,xx_op_T5_jsr_i1, xx_op_T5_jsr_v);
  spice_node_3 n_idl3(eclk, ereset, idl3_i0,idl3_i1,idl3_i2, idl3_v);
  spice_node_1 n_notidl7(eclk, ereset, notidl7_i1, notidl7_v);
  spice_node_2 n_n319(eclk, ereset, n319_i0,n319_i1, n319_v);
  spice_node_3 n_n318(eclk, ereset, n318_i0,n318_i1,n318_i3, n318_v);
  spice_node_2 n_n312(eclk, ereset, n312_i1,n312_i2, n312_v);
  spice_node_2 n_n311(eclk, ereset, n311_i0,n311_i1, n311_v);
  spice_node_2 n_n310(eclk, ereset, n310_i0,n310_i2, n310_v);
  spice_node_2 n_n317(eclk, ereset, n317_i0,n317_i2, n317_v);
  spice_node_6 n_adh3(eclk, ereset, adh3_i0,adh3_i2,adh3_i3,adh3_i4,adh3_i5,adh3_i6, adh3_v);
  spice_node_4 n_alu5(eclk, ereset, alu5_i0,alu5_i1,alu5_i3,alu5_i4, alu5_v);
  spice_node_2 n_n1335(eclk, ereset, n1335_i0,n1335_i1, n1335_v);
  spice_node_2 n_dpc35_PCHC(eclk, ereset, dpc35_PCHC_i0,dpc35_PCHC_i1, dpc35_PCHC_v);
  spice_node_2 n_n441(eclk, ereset, n441_i0,n441_i1, n441_v);
  spice_node_3 n_n440(eclk, ereset, n440_i0,n440_i1,n440_i2, n440_v);
  spice_node_2 n_dpc26_ACDB(eclk, ereset, dpc26_ACDB_i0,dpc26_ACDB_i9, dpc26_ACDB_v);
  spice_node_1 n_n1333(eclk, ereset, n1333_i1, n1333_v);
  spice_node_2 n_dor3(eclk, ereset, dor3_i1,dor3_i2, dor3_v);
  spice_node_3 n_n632(eclk, ereset, n632_i0,n632_i1,n632_i2, n632_v);
  spice_node_2 n_n1521(eclk, ereset, n1521_i1,n1521_i2, n1521_v);
  spice_node_1 n_n633(eclk, ereset, n633_i0, n633_v);
  spice_node_2 n_n964(eclk, ereset, n964_i0,n964_i2, n964_v);
  spice_node_3 n___AxBxC_1(eclk, ereset, __AxBxC_1_i0,__AxBxC_1_i1,__AxBxC_1_i2, __AxBxC_1_v);
  spice_node_2 n_n966(eclk, ereset, n966_i0,n966_i3, n966_v);
  spice_node_3 n_nnT2BR(eclk, ereset, nnT2BR_i0,nnT2BR_i1,nnT2BR_i2, nnT2BR_v);
  spice_node_1 n_pipeUNK32(eclk, ereset, pipeUNK32_i0, pipeUNK32_v);
  spice_node_3 n_n961(eclk, ereset, n961_i0,n961_i1,n961_i2, n961_v);
  spice_node_2 n_n962(eclk, ereset, n962_i0,n962_i1, n962_v);
  spice_node_2 n_n963(eclk, ereset, n963_i1,n963_i2, n963_v);
  spice_node_1 n_n968(eclk, ereset, n968_i1, n968_v);
  spice_node_2 n_n969(eclk, ereset, n969_i0,n969_i1, n969_v);
  spice_node_2 n_n400(eclk, ereset, n400_i2,n400_i3, n400_v);
  spice_node_2 n_AxB7(eclk, ereset, AxB7_i1,AxB7_i3, AxB7_v);
  spice_node_1 n_n878(eclk, ereset, n878_i0, n878_v);
  spice_node_2 n_n1240(eclk, ereset, n1240_i1,n1240_i2, n1240_v);
  spice_node_2 n_n876(eclk, ereset, n876_i0,n876_i1, n876_v);
  spice_node_2 n_n877(eclk, ereset, n877_i0,n877_i1, n877_v);
  spice_node_2 n_dpc6_SBS(eclk, ereset, dpc6_SBS_i8,dpc6_SBS_i9, dpc6_SBS_v);
  spice_node_3 n_n875(eclk, ereset, n875_i0,n875_i1,n875_i2, n875_v);
  spice_node_4 n_alu1(eclk, ereset, alu1_i0,alu1_i1,alu1_i3,alu1_i4, alu1_v);
  spice_node_2 n_op_T__ora_and_eor_adc(eclk, ereset, op_T__ora_and_eor_adc_i0,op_T__ora_and_eor_adc_i2, op_T__ora_and_eor_adc_v);
  spice_node_3 n_idl1(eclk, ereset, idl1_i0,idl1_i1,idl1_i2, idl1_v);
  spice_node_4 n_n871(eclk, ereset, n871_i0,n871_i1,n871_i2,n871_i3, n871_v);
  spice_node_8 n_adl2(eclk, ereset, adl2_i0,adl2_i1,adl2_i2,adl2_i3,adl2_i4,adl2_i5,adl2_i6,adl2_i8, adl2_v);
  spice_node_1 n_n9(eclk, ereset, n9_i0, n9_v);
  spice_node_1 n_n1533(eclk, ereset, n1533_i1, n1533_v);
  spice_node_1 n_n644(eclk, ereset, n644_i0, n644_v);
  spice_node_2 n_n890(eclk, ereset, n890_i1,n890_i2, n890_v);
  spice_node_8 n_idb4(eclk, ereset, idb4_i0,idb4_i3,idb4_i4,idb4_i5,idb4_i6,idb4_i7,idb4_i8,idb4_i9, idb4_v);
  spice_node_1 n_notalu5(eclk, ereset, notalu5_i0, notalu5_v);
  spice_node_1 n_pd3(eclk, ereset, pd3_i0, pd3_v);
  spice_node_2 n_n1247(eclk, ereset, n1247_i0,n1247_i1, n1247_v);
  spice_node_3 n_n896(eclk, ereset, n896_i0,n896_i1,n896_i2, n896_v);
  spice_node_1 n_n897(eclk, ereset, n897_i0, n897_v);
  spice_node_2 n_dpc39_PCLPCL(eclk, ereset, dpc39_PCLPCL_i8,dpc39_PCLPCL_i9, dpc39_PCLPCL_v);
  spice_node_1 n_pipeUNK18(eclk, ereset, pipeUNK18_i1, pipeUNK18_v);
  spice_node_1 n_pipeUNK01(eclk, ereset, pipeUNK01_i0, pipeUNK01_v);
  spice_node_2 n_n641(eclk, ereset, n641_i0,n641_i2, n641_v);
  spice_node_2 n__ABH2(eclk, ereset, _ABH2_i1,_ABH2_i2, _ABH2_v);
  spice_node_2 n_n769(eclk, ereset, n769_i1,n769_i2, n769_v);
  spice_node_2 n_n762(eclk, ereset, n762_i1,n762_i2, n762_v);
  spice_node_2 n_n763(eclk, ereset, n763_i0,n763_i1, n763_v);
  spice_node_1 n_n760(eclk, ereset, n760_i0, n760_v);
  spice_node_2 n_clock1(eclk, ereset, clock1_i1,clock1_i33, clock1_v);
  spice_node_4 n_n767(eclk, ereset, n767_i0,n767_i1,n767_i2,n767_i3, n767_v);
  spice_node_2 n_op_jmp(eclk, ereset, op_jmp_i0,op_jmp_i1, op_jmp_v);
  spice_node_4 n_alu7(eclk, ereset, alu7_i0,alu7_i1,alu7_i2,alu7_i3, alu7_v);
  spice_node_1 n_pipeUNK17(eclk, ereset, pipeUNK17_i0, pipeUNK17_v);
  spice_node_2 n_pclp2(eclk, ereset, pclp2_i1,pclp2_i2, pclp2_v);
  spice_node_2 n_n1076(eclk, ereset, n1076_i0,n1076_i2, n1076_v);
  spice_node_2 n_clearIR(eclk, ereset, clearIR_i0,clearIR_i9, clearIR_v);
  spice_node_2 n_op_T0_shift_right_a(eclk, ereset, op_T0_shift_right_a_i0,op_T0_shift_right_a_i1, op_T0_shift_right_a_v);
  spice_node_3 n_n1075(eclk, ereset, n1075_i0,n1075_i1,n1075_i2, n1075_v);
  spice_node_2 n_n1072(eclk, ereset, n1072_i0,n1072_i2, n1072_v);
  spice_node_3 n_n1073(eclk, ereset, n1073_i0,n1073_i1,n1073_i2, n1073_v);
  spice_node_2 n_n1070(eclk, ereset, n1070_i0,n1070_i1, n1070_v);
  spice_node_6 n_n1071(eclk, ereset, n1071_i0,n1071_i1,n1071_i2,n1071_i3,n1071_i4,n1071_i5, n1071_v);
  spice_node_3 n_alub5(eclk, ereset, alub5_i0,alub5_i1,alub5_i2, alub5_v);
  spice_node_1 n_n1679(eclk, ereset, n1679_i0, n1679_v);
  spice_node_1 n_n1674(eclk, ereset, n1674_i0, n1674_v);
  spice_node_2 n_n1675(eclk, ereset, n1675_i0,n1675_i2, n1675_v);
  spice_node_2 n_n1676(eclk, ereset, n1676_i2,n1676_i3, n1676_v);
  spice_node_2 n_n1677(eclk, ereset, n1677_i2,n1677_i3, n1677_v);
  spice_node_2 n_pch0(eclk, ereset, pch0_i1,pch0_i2, pch0_v);
  spice_node_2 n_pd2_clearIR(eclk, ereset, pd2_clearIR_i1,pd2_clearIR_i2, pd2_clearIR_v);
  spice_node_2 n_so(eclk, ereset, so_i1,so_i2, so_v);
  spice_node_1 n_n1673(eclk, ereset, n1673_i0, n1673_v);
  spice_node_3 n_n1094(eclk, ereset, n1094_i0,n1094_i1,n1094_i2, n1094_v);
  spice_node_4 n_n1095(eclk, ereset, n1095_i0,n1095_i1,n1095_i2,n1095_i3, n1095_v);
  spice_node_2 n_abl0(eclk, ereset, abl0_i3,abl0_i4, abl0_v);
  spice_node_2 n_n1097(eclk, ereset, n1097_i0,n1097_i1, n1097_v);
  spice_node_3 n_n678(eclk, ereset, n678_i0,n678_i2,n678_i3, n678_v);
  spice_node_3 n_n1091(eclk, ereset, n1091_i0,n1091_i1,n1091_i2, n1091_v);
  spice_node_3 n_n642(eclk, ereset, n642_i0,n642_i1,n642_i3, n642_v);
  spice_node_3 n_n674(eclk, ereset, n674_i0,n674_i1,n674_i2, n674_v);
  spice_node_1 n_n675(eclk, ereset, n675_i1, n675_v);
  spice_node_3 n_n676(eclk, ereset, n676_i0,n676_i2,n676_i3, n676_v);
  spice_node_2 n_op_T3_abs_idx_ind(eclk, ereset, op_T3_abs_idx_ind_i0,op_T3_abs_idx_ind_i2, op_T3_abs_idx_ind_v);
  spice_node_2 n_n670(eclk, ereset, n670_i2,n670_i3, n670_v);
  spice_node_1 n_n671(eclk, ereset, n671_i0, n671_v);
  spice_node_3 n_ab14(eclk, ereset, ab14_i0,ab14_i1,ab14_i2, ab14_v);
  spice_node_2 n_n673(eclk, ereset, n673_i0,n673_i2, n673_v);
  spice_node_1 n_notdor6(eclk, ereset, notdor6_i0, notdor6_v);
  spice_node_2 n_op_T0_cld_sed(eclk, ereset, op_T0_cld_sed_i1,op_T0_cld_sed_i2, op_T0_cld_sed_v);
  spice_node_2 n_pd7_clearIR(eclk, ereset, pd7_clearIR_i1,pd7_clearIR_i3, pd7_clearIR_v);
  spice_node_1 n_n1411(eclk, ereset, n1411_i1, n1411_v);
  spice_node_2 n_n1412(eclk, ereset, n1412_i0,n1412_i1, n1412_v);
  spice_node_2 n_n1413(eclk, ereset, n1413_i1,n1413_i2, n1413_v);
  spice_node_4 n_alu3(eclk, ereset, alu3_i0,alu3_i1,alu3_i2,alu3_i3, alu3_v);
  spice_node_2 n_dor6(eclk, ereset, dor6_i0,dor6_i2, dor6_v);
  spice_node_2 n_n1416(eclk, ereset, n1416_i0,n1416_i1, n1416_v);
  spice_node_2 n_n1417(eclk, ereset, n1417_i0,n1417_i2, n1417_v);
  spice_node_2 n_n1323(eclk, ereset, n1323_i0,n1323_i2, n1323_v);
  spice_node_3 n_notir7(eclk, ereset, notir7_i0,notir7_i1,notir7_i2, notir7_v);
  spice_node_2 n_s3(eclk, ereset, s3_i0,s3_i1, s3_v);
  spice_node_1 n_pclp5(eclk, ereset, pclp5_i1, pclp5_v);
  spice_node_2 n__C78(eclk, ereset, _C78_i1,_C78_i2, _C78_v);
  spice_node_2 n_op_T__shift_a(eclk, ereset, op_T__shift_a_i0,op_T__shift_a_i2, op_T__shift_a_v);
  spice_node_2 n_n1325(eclk, ereset, n1325_i1,n1325_i2, n1325_v);
  spice_node_2 n_ir7(eclk, ereset, ir7_i2,ir7_i3, ir7_v);
  spice_node_2 n_ir5(eclk, ereset, ir5_i0,ir5_i2, ir5_v);
  spice_node_2 n_n5(eclk, ereset, n5_i0,n5_i2, n5_v);
  spice_node_2 n_n647(eclk, ereset, n647_i0,n647_i1, n647_v);
  spice_node_2 n_op_T2_ind(eclk, ereset, op_T2_ind_i0,op_T2_ind_i1, op_T2_ind_v);
  spice_node_2 n_n1257(eclk, ereset, n1257_i0,n1257_i2, n1257_v);
  spice_node_3 n_n1254(eclk, ereset, n1254_i0,n1254_i1,n1254_i2, n1254_v);
  spice_node_1 n_n1527(eclk, ereset, n1527_i0, n1527_v);
  spice_node_2 n_op_plp_pla(eclk, ereset, op_plp_pla_i0,op_plp_pla_i1, op_plp_pla_v);
  spice_node_2 n_n1253(eclk, ereset, n1253_i0,n1253_i1, n1253_v);
  spice_node_2 n_alua7(eclk, ereset, alua7_i0,alua7_i1, alua7_v);
  spice_node_2 n_n1523(eclk, ereset, n1523_i2,n1523_i3, n1523_v);
  spice_node_1 n_n1528(eclk, ereset, n1528_i0, n1528_v);
  spice_node_1 n_n1529(eclk, ereset, n1529_i1, n1529_v);
  spice_node_2 n_n1258(eclk, ereset, n1258_i0,n1258_i1, n1258_v);
  spice_node_2 n_op_T4_ind_x(eclk, ereset, op_T4_ind_x_i0,op_T4_ind_x_i2, op_T4_ind_x_v);
  spice_node_3 n___AxB_4(eclk, ereset, __AxB_4_i0,__AxB_4_i1,__AxB_4_i3, __AxB_4_v);
  spice_node_2 n_op_T2_jmp_abs(eclk, ereset, op_T2_jmp_abs_i0,op_T2_jmp_abs_i1, op_T2_jmp_abs_v);
  spice_node_2 n_n300(eclk, ereset, n300_i1,n300_i2, n300_v);
  spice_node_2 n_op_T__cmp(eclk, ereset, op_T__cmp_i0,op_T__cmp_i1, op_T__cmp_v);
  spice_node_2 n_PD_xxx010x1(eclk, ereset, PD_xxx010x1_i0,PD_xxx010x1_i1, PD_xxx010x1_v);
  spice_node_2 n_op_T0_bit(eclk, ereset, op_T0_bit_i0,op_T0_bit_i1, op_T0_bit_v);
  spice_node_6 n_n304(eclk, ereset, n304_i0,n304_i1,n304_i2,n304_i3,n304_i4,n304_i5, n304_v);
  spice_node_2 n_y3(eclk, ereset, y3_i0,y3_i2, y3_v);
  spice_node_3 n_n306(eclk, ereset, n306_i0,n306_i1,n306_i2, n306_v);
  spice_node_2 n_n307(eclk, ereset, n307_i0,n307_i2, n307_v);
  spice_node_3 n_n473(eclk, ereset, n473_i0,n473_i1,n473_i2, n473_v);
  spice_node_2 n_DA_C01(eclk, ereset, DA_C01_i0,DA_C01_i3, DA_C01_v);
  spice_node_3 n_n959(eclk, ereset, n959_i0,n959_i1,n959_i2, n959_v);
  spice_node_3 n_n958(eclk, ereset, n958_i0,n958_i1,n958_i3, n958_v);
  spice_node_2 n_n951(eclk, ereset, n951_i0,n951_i3, n951_v);
  spice_node_2 n_op_T__cpx_cpy_abs(eclk, ereset, op_T__cpx_cpy_abs_i0,op_T__cpx_cpy_abs_i1, op_T__cpx_cpy_abs_v);
  spice_node_3 n_n953(eclk, ereset, n953_i0,n953_i1,n953_i2, n953_v);
  spice_node_3 n_n952(eclk, ereset, n952_i0,n952_i1,n952_i2, n952_v);
  spice_node_1 n_pd2(eclk, ereset, pd2_i0, pd2_v);
  spice_node_2 n_n954(eclk, ereset, n954_i0,n954_i1, n954_v);
  spice_node_6 n_notaluoutmux0(eclk, ereset, notaluoutmux0_i0,notaluoutmux0_i1,notaluoutmux0_i2,notaluoutmux0_i3,notaluoutmux0_i4,notaluoutmux0_i5, notaluoutmux0_v);
  spice_node_2 n_n956(eclk, ereset, n956_i0,n956_i1, n956_v);
  spice_node_2 n_n507(eclk, ereset, n507_i0,n507_i1, n507_v);
  spice_node_2 n_dpc2_XSB(eclk, ereset, dpc2_XSB_i2,dpc2_XSB_i9, dpc2_XSB_v);
  spice_node_1 n_n666(eclk, ereset, n666_i1, n666_v);
  spice_node_3 n_n504(eclk, ereset, n504_i0,n504_i1,n504_i2, n504_v);
  spice_node_2 n_n1260(eclk, ereset, n1260_i2,n1260_i3, n1260_v);
  spice_node_4 n_n719(eclk, ereset, n719_i0,n719_i1,n719_i2,n719_i3, n719_v);
  spice_node_3 n_n718(eclk, ereset, n718_i0,n718_i1,n718_i2, n718_v);
  spice_node_2 n_n717(eclk, ereset, n717_i1,n717_i2, n717_v);
  spice_node_2 n_n715(eclk, ereset, n715_i0,n715_i1, n715_v);
  spice_node_2 n_n714(eclk, ereset, n714_i1,n714_i2, n714_v);
  spice_node_2 n_abh1(eclk, ereset, abh1_i3,abh1_i4, abh1_v);
  spice_node_2 n_op_T2_jsr(eclk, ereset, op_T2_jsr_i1,op_T2_jsr_i3, op_T2_jsr_v);
  spice_node_2 n_cp1(eclk, ereset, cp1_i35,cp1_i57, cp1_v);
  spice_node_2 n_n1265(eclk, ereset, n1265_i1,n1265_i2, n1265_v);
  spice_node_3 n_n1069(eclk, ereset, n1069_i0,n1069_i1,n1069_i2, n1069_v);
  spice_node_2 n_dpc8_nDBADD(eclk, ereset, dpc8_nDBADD_i3,dpc8_nDBADD_i9, dpc8_nDBADD_v);
  spice_node_1 n_n1061(eclk, ereset, n1061_i1, n1061_v);
  spice_node_2 n_dpc25_SBDB(eclk, ereset, dpc25_SBDB_i0,dpc25_SBDB_i9, dpc25_SBDB_v);
  spice_node_4 n_n1063(eclk, ereset, n1063_i0,n1063_i1,n1063_i2,n1063_i4, n1063_v);
  spice_node_2 n__ABH0(eclk, ereset, _ABH0_i1,_ABH0_i2, _ABH0_v);
  spice_node_3 n_n1065(eclk, ereset, n1065_i0,n1065_i1,n1065_i2, n1065_v);
  spice_node_1 n_nots1(eclk, ereset, nots1_i1, nots1_v);
  spice_node_2 n_n1067(eclk, ereset, n1067_i0,n1067_i2, n1067_v);
  spice_node_3 n_idl2(eclk, ereset, idl2_i0,idl2_i1,idl2_i2, idl2_v);
  spice_node_1 n_pd6(eclk, ereset, pd6_i0, pd6_v);
  spice_node_3 n_n1668(eclk, ereset, n1668_i0,n1668_i1,n1668_i2, n1668_v);
  spice_node_2 n_dpc16_EORS(eclk, ereset, dpc16_EORS_i8,dpc16_EORS_i9, dpc16_EORS_v);
  spice_node_2 n_op_T__asl_rol_a(eclk, ereset, op_T__asl_rol_a_i0,op_T__asl_rol_a_i1, op_T__asl_rol_a_v);
  spice_node_2 n_op_T__inx(eclk, ereset, op_T__inx_i0,op_T__inx_i1, op_T__inx_v);
  spice_node_2 n_n1662(eclk, ereset, n1662_i0,n1662_i1, n1662_v);
  spice_node_4 n_n1661(eclk, ereset, n1661_i0,n1661_i1,n1661_i2,n1661_i3, n1661_v);
  spice_node_2 n_n1660(eclk, ereset, n1660_i0,n1660_i3, n1660_v);
  spice_node_3 n_n1087(eclk, ereset, n1087_i0,n1087_i1,n1087_i2, n1087_v);
  spice_node_2 n_op_T2_pha(eclk, ereset, op_T2_pha_i0,op_T2_pha_i1, op_T2_pha_v);
  spice_node_2 n_n593(eclk, ereset, n593_i1,n593_i2, n593_v);
  spice_node_3 n_n1084(eclk, ereset, n1084_i0,n1084_i2,n1084_i3, n1084_v);
  spice_node_2 n_n595(eclk, ereset, n595_i1,n595_i2, n595_v);
  spice_node_3 n_n1082(eclk, ereset, n1082_i0,n1082_i1,n1082_i2, n1082_v);
  spice_node_3 n_n1081(eclk, ereset, n1081_i0,n1081_i1,n1081_i2, n1081_v);
  spice_node_1 n_n599(eclk, ereset, n599_i1, n599_v);
  spice_node_1 n_n598(eclk, ereset, n598_i0, n598_v);
  spice_node_3 n_n1089(eclk, ereset, n1089_i0,n1089_i1,n1089_i2, n1089_v);
  spice_node_2 n_dor4(eclk, ereset, dor4_i1,dor4_i2, dor4_v);
  spice_node_1 n_n1409(eclk, ereset, n1409_i0, n1409_v);
  spice_node_2 n_n1408(eclk, ereset, n1408_i0,n1408_i2, n1408_v);
  spice_node_2 n_s0(eclk, ereset, s0_i0,s0_i1, s0_v);
  spice_node_3 n_n1402(eclk, ereset, n1402_i0,n1402_i1,n1402_i2, n1402_v);
  spice_node_2 n_n1401(eclk, ereset, n1401_i0,n1401_i1, n1401_v);
  spice_node_2 n_n1400(eclk, ereset, n1400_i0,n1400_i2, n1400_v);
  spice_node_13 n_dasb4(eclk, ereset, dasb4_i0,dasb4_i1,dasb4_i2,dasb4_i3,dasb4_i4,dasb4_i5,dasb4_i6,dasb4_i7,dasb4_i8,dasb4_i9,dasb4_i10,dasb4_i11,dasb4_i12, dasb4_v);
  spice_node_1 n_n1404(eclk, ereset, n1404_i0, n1404_v);
  spice_node_1 n_pipephi2Reset0(eclk, ereset, pipephi2Reset0_i0, pipephi2Reset0_v);
  spice_node_2 n_x6(eclk, ereset, x6_i0,x6_i1, x6_v);
  spice_node_3 n_n1339(eclk, ereset, n1339_i0,n1339_i1,n1339_i2, n1339_v);
  spice_node_1 n_n1338(eclk, ereset, n1338_i0, n1338_v);
  spice_node_2 n_aluaorb0(eclk, ereset, aluaorb0_i0,aluaorb0_i1, aluaorb0_v);
  spice_node_1 n_pipeUNK06(eclk, ereset, pipeUNK06_i0, pipeUNK06_v);
  spice_node_3 n_n442(eclk, ereset, n442_i0,n442_i1,n442_i2, n442_v);
  spice_node_2 n_op_T0_cpx_cpy_inx_iny(eclk, ereset, op_T0_cpx_cpy_inx_iny_i0,op_T0_cpx_cpy_inx_iny_i1, op_T0_cpx_cpy_inx_iny_v);
  spice_node_12 n_sb6(eclk, ereset, sb6_i0,sb6_i1,sb6_i2,sb6_i3,sb6_i4,sb6_i6,sb6_i7,sb6_i8,sb6_i9,sb6_i10,sb6_i11,sb6_i12, sb6_v);
  spice_node_2 n_x_op_T3_abs_idx(eclk, ereset, x_op_T3_abs_idx_i0,x_op_T3_abs_idx_i2, x_op_T3_abs_idx_v);
  spice_node_2 n_op_T5_rti_rts(eclk, ereset, op_T5_rti_rts_i0,op_T5_rti_rts_i1, op_T5_rti_rts_v);
  spice_node_2 n_n445(eclk, ereset, n445_i3,n445_i4, n445_v);
  spice_node_2 n_alua2(eclk, ereset, alua2_i0,alua2_i1, alua2_v);
  spice_node_2 n_n1545(eclk, ereset, n1545_i1,n1545_i2, n1545_v);
  spice_node_2 n_n1542(eclk, ereset, n1542_i0,n1542_i3, n1542_v);
  spice_node_2 n_x_op_T0_txa(eclk, ereset, x_op_T0_txa_i0,x_op_T0_txa_i1, x_op_T0_txa_v);
  spice_node_2 n_pclp4(eclk, ereset, pclp4_i0,pclp4_i2, pclp4_v);
  spice_node_2 n_n38(eclk, ereset, n38_i1,n38_i2, n38_v);
  spice_node_2 n_op_from_x(eclk, ereset, op_from_x_i0,op_from_x_i1, op_from_x_v);
  spice_node_2 n_pchp5(eclk, ereset, pchp5_i1,pchp5_i2, pchp5_v);
  spice_node_1 n_p0(eclk, ereset, p0_i0, p0_v);
  spice_node_3 n_n31(eclk, ereset, n31_i0,n31_i2,n31_i4, n31_v);
  spice_node_3 n_n695(eclk, ereset, n695_i0,n695_i1,n695_i2, n695_v);
  spice_node_2 n_n37(eclk, ereset, n37_i1,n37_i2, n37_v);
  spice_node_2 n_n36(eclk, ereset, n36_i0,n36_i1, n36_v);
  spice_node_2 n_n35(eclk, ereset, n35_i2,n35_i3, n35_v);
  spice_node_3 n_n34(eclk, ereset, n34_i0,n34_i1,n34_i2, n34_v);
  spice_node_1 n_notidl6(eclk, ereset, notidl6_i1, notidl6_v);
  spice_node_2 n_AxB3(eclk, ereset, AxB3_i1,AxB3_i4, AxB3_v);
  spice_node_2 n_n643(eclk, ereset, n643_i1,n643_i2, n643_v);
  spice_node_2 n_n1534(eclk, ereset, n1534_i2,n1534_i3, n1534_v);
  spice_node_3 n_n645(eclk, ereset, n645_i0,n645_i1,n645_i2, n645_v);
  spice_node_2 n_n1244(eclk, ereset, n1244_i0,n1244_i1, n1244_v);
  spice_node_4 n_n1531(eclk, ereset, n1531_i0,n1531_i1,n1531_i2,n1531_i3, n1531_v);
  spice_node_2 n_n646(eclk, ereset, n646_i0,n646_i2, n646_v);
  spice_node_3 n_n649(eclk, ereset, n649_i0,n649_i2,n649_i3, n649_v);
  spice_node_2 n_alua1(eclk, ereset, alua1_i0,alua1_i1, alua1_v);
  spice_node_6 n_adh7(eclk, ereset, adh7_i0,adh7_i1,adh7_i2,adh7_i3,adh7_i4,adh7_i5, adh7_v);
  spice_node_1 n_n339(eclk, ereset, n339_i1, n339_v);
  spice_node_1 n_pipeUNK08(eclk, ereset, pipeUNK08_i0, pipeUNK08_v);
  spice_node_2 n_n335(eclk, ereset, n335_i0,n335_i1, n335_v);
  spice_node_3 n_n334(eclk, ereset, n334_i2,n334_i3,n334_i4, n334_v);
  spice_node_2 n_ir6(eclk, ereset, ir6_i2,ir6_i3, ir6_v);
  spice_node_4 n_n336(eclk, ereset, n336_i0,n336_i1,n336_i3,n336_i5, n336_v);
  spice_node_4 n_alu6(eclk, ereset, alu6_i0,alu6_i1,alu6_i2,alu6_i4, alu6_v);
  spice_node_3 n_n330(eclk, ereset, n330_i0,n330_i1,n330_i3, n330_v);
  spice_node_3 n_DC78(eclk, ereset, DC78_i0,DC78_i1,DC78_i2, DC78_v);
  spice_node_5 n_n332(eclk, ereset, n332_i0,n332_i1,n332_i2,n332_i3,n332_i4, n332_v);
  spice_node_2 n_n1026(eclk, ereset, n1026_i0,n1026_i3, n1026_v);
  spice_node_2 n_n8(eclk, ereset, n8_i0,n8_i1, n8_v);
  spice_node_2 n_n1462(eclk, ereset, n1462_i0,n1462_i2, n1462_v);
  spice_node_3 n_INTG(eclk, ereset, INTG_i0,INTG_i1,INTG_i2, INTG_v);
  spice_node_2 n_pch4(eclk, ereset, pch4_i1,pch4_i2, pch4_v);
  spice_node_2 n_n946(eclk, ereset, n946_i0,n946_i2, n946_v);
  spice_node_2 n_n947(eclk, ereset, n947_i1,n947_i2, n947_v);
  spice_node_3 n_n944(eclk, ereset, n944_i0,n944_i1,n944_i2, n944_v);
  spice_node_3 n_db2(eclk, ereset, db2_i1,db2_i2,db2_i4, db2_v);
  spice_node_2 n_cclk(eclk, ereset, cclk_i24,cclk_i207, cclk_v);
  spice_node_1 n_pipeT5out(eclk, ereset, pipeT5out_i0, pipeT5out_v);
  spice_node_2 n_n133(eclk, ereset, n133_i2,n133_i3, n133_v);
  spice_node_3 n_n132(eclk, ereset, n132_i0,n132_i1,n132_i2, n132_v);
  spice_node_2 n_op_T0_pla(eclk, ereset, op_T0_pla_i0,op_T0_pla_i2, op_T0_pla_v);
  spice_node_2 n_n130(eclk, ereset, n130_i0,n130_i2, n130_v);
  spice_node_2 n_n135(eclk, ereset, n135_i1,n135_i2, n135_v);
  spice_node_2 n_n134(eclk, ereset, n134_i0,n134_i1, n134_v);
  spice_node_2 n_n139(eclk, ereset, n139_i0,n139_i1, n139_v);
  spice_node_3 n_n138(eclk, ereset, n138_i0,n138_i1,n138_i2, n138_v);
  spice_node_2 n_n708(eclk, ereset, n708_i0,n708_i1, n708_v);
  spice_node_2 n_n709(eclk, ereset, n709_i0,n709_i2, n709_v);
  spice_node_3 n_alub2(eclk, ereset, alub2_i0,alub2_i1,alub2_i2, alub2_v);
  spice_node_1 n_pipeT3out(eclk, ereset, pipeT3out_i0, pipeT3out_v);
  spice_node_2 n__ABL2(eclk, ereset, _ABL2_i1,_ABL2_i2, _ABL2_v);
  spice_node_3 n_n700(eclk, ereset, n700_i0,n700_i1,n700_i2, n700_v);
  spice_node_3 n___AxB_2(eclk, ereset, __AxB_2_i0,__AxB_2_i1,__AxB_2_i3, __AxB_2_v);
  spice_node_3 n_notir1(eclk, ereset, notir1_i0,notir1_i1,notir1_i2, notir1_v);
  spice_node_1 n_n88(eclk, ereset, n88_i1, n88_v);
  spice_node_2 n_rdy(eclk, ereset, rdy_i1,rdy_i2, rdy_v);
  spice_node_3 n_db1(eclk, ereset, db1_i1,db1_i3,db1_i4, db1_v);
  spice_node_2 n_n83(eclk, ereset, n83_i0,n83_i1, n83_v);
  spice_node_3 n_n80(eclk, ereset, n80_i0,n80_i1,n80_i2, n80_v);
  spice_node_2 n_s2(eclk, ereset, s2_i0,s2_i1, s2_v);
  spice_node_3 n_n86(eclk, ereset, n86_i0,n86_i2,n86_i3, n86_v);
  spice_node_4 n_n87(eclk, ereset, n87_i0,n87_i1,n87_i2,n87_i3, n87_v);
  spice_node_2 n_op_T2_ind_x(eclk, ereset, op_T2_ind_x_i0,op_T2_ind_x_i1, op_T2_ind_x_v);
  spice_node_2 n_x4(eclk, ereset, x4_i0,x4_i1, x4_v);
  spice_node_2 n_op_T0_cpx_inx(eclk, ereset, op_T0_cpx_inx_i0,op_T0_cpx_inx_i1, op_T0_cpx_inx_v);
  spice_node_1 n_pipeUNK30(eclk, ereset, pipeUNK30_i0, pipeUNK30_v);
  spice_node_2 n_a7(eclk, ereset, a7_i1,a7_i2, a7_v);
  spice_node_3 n_n1650(eclk, ereset, n1650_i0,n1650_i1,n1650_i2, n1650_v);
  spice_node_6 n_adh2(eclk, ereset, adh2_i0,adh2_i1,adh2_i3,adh2_i4,adh2_i5,adh2_i6, adh2_v);
  spice_node_3 n_n1657(eclk, ereset, n1657_i0,n1657_i1,n1657_i2, n1657_v);
  spice_node_5 n_n1654(eclk, ereset, n1654_i0,n1654_i1,n1654_i2,n1654_i3,n1654_i4, n1654_v);
  spice_node_2 n_n1655(eclk, ereset, n1655_i0,n1655_i1, n1655_v);
  spice_node_3 n_n586(eclk, ereset, n586_i0,n586_i1,n586_i2, n586_v);
  spice_node_2 n_n587(eclk, ereset, n587_i0,n587_i1, n587_v);
  spice_node_2 n_pch3(eclk, ereset, pch3_i1,pch3_i2, pch3_v);
  spice_node_2 n_n582(eclk, ereset, n582_i2,n582_i3, n582_v);
  spice_node_3 n_n583(eclk, ereset, n583_i0,n583_i1,n583_i2, n583_v);
  spice_node_1 n_n581(eclk, ereset, n581_i1, n581_v);
  spice_node_3 n_n588(eclk, ereset, n588_i0,n588_i1,n588_i2, n588_v);
  spice_node_2 n_x5(eclk, ereset, x5_i1,x5_i2, x5_v);
  spice_node_1 n_pipeUNK03(eclk, ereset, pipeUNK03_i0, pipeUNK03_v);
  spice_node_7 n_adl4(eclk, ereset, adl4_i0,adl4_i1,adl4_i3,adl4_i4,adl4_i5,adl4_i6,adl4_i7, adl4_v);
  spice_node_2 n_n1434(eclk, ereset, n1434_i0,n1434_i2, n1434_v);
  spice_node_2 n_s7(eclk, ereset, s7_i0,s7_i2, s7_v);
  spice_node_3 n_alub1(eclk, ereset, alub1_i0,alub1_i1,alub1_i2, alub1_v);
  spice_node_2 n_n1433(eclk, ereset, n1433_i0,n1433_i2, n1433_v);
  spice_node_2 n_x_op_T3_plp_pla(eclk, ereset, x_op_T3_plp_pla_i0,x_op_T3_plp_pla_i1, x_op_T3_plp_pla_v);
  spice_node_1 n_pipe_VEC(eclk, ereset, pipe_VEC_i0, pipe_VEC_v);
  spice_node_1 n_nots0(eclk, ereset, nots0_i0, nots0_v);
  spice_node_1 n_pipeUNK41(eclk, ereset, pipeUNK41_i0, pipeUNK41_v);
  spice_node_2 n_n1439(eclk, ereset, n1439_i1,n1439_i2, n1439_v);
  spice_node_3 n_db7(eclk, ereset, db7_i1,db7_i2,db7_i4, db7_v);
  spice_node_1 n_n459(eclk, ereset, n459_i0, n459_v);
  spice_node_3 n_dasb2(eclk, ereset, dasb2_i0,dasb2_i1,dasb2_i2, dasb2_v);
  spice_node_1 n_n1341(eclk, ereset, n1341_i1, n1341_v);
  spice_node_2 n_op_T0_acc(eclk, ereset, op_T0_acc_i0,op_T0_acc_i1, op_T0_acc_v);
  spice_node_2 n_n1343(eclk, ereset, n1343_i0,n1343_i1, n1343_v);
  spice_node_1 n_pipeUNK40(eclk, ereset, pipeUNK40_i0, pipeUNK40_v);
  spice_node_3 n_n457(eclk, ereset, n457_i0,n457_i1,n457_i2, n457_v);
  spice_node_2 n_n1377(eclk, ereset, n1377_i0,n1377_i1, n1377_v);
  spice_node_7 n_idb5(eclk, ereset, idb5_i1,idb5_i3,idb5_i4,idb5_i5,idb5_i6,idb5_i7,idb5_i8, idb5_v);
  spice_node_2 n_dpc7_SS(eclk, ereset, dpc7_SS_i7,dpc7_SS_i9, dpc7_SS_v);
  spice_node_2 n_n1501(eclk, ereset, n1501_i1,n1501_i2, n1501_v);
  spice_node_2 n__C01(eclk, ereset, _C01_i0,_C01_i1, _C01_v);
  spice_node_1 n_n653(eclk, ereset, n653_i0, n653_v);
  spice_node_3 n_db3(eclk, ereset, db3_i1,db3_i2,db3_i4, db3_v);
  spice_node_3 n___AxBxC_4(eclk, ereset, __AxBxC_4_i0,__AxBxC_4_i1,__AxBxC_4_i2, __AxBxC_4_v);
  spice_node_1 n_n1509(eclk, ereset, n1509_i0, n1509_v);
  spice_node_4 n_n658(eclk, ereset, n658_i0,n658_i1,n658_i2,n658_i3, n658_v);
  spice_node_2 n_DA_AxB2(eclk, ereset, DA_AxB2_i0,DA_AxB2_i2, DA_AxB2_v);
  spice_node_1 n_n55(eclk, ereset, n55_i0, n55_v);
  spice_node_2 n_n322(eclk, ereset, n322_i1,n322_i2, n322_v);
  spice_node_1 n_n323(eclk, ereset, n323_i0, n323_v);
  spice_node_2 n_n320(eclk, ereset, n320_i0,n320_i1, n320_v);
  spice_node_2 n_n321(eclk, ereset, n321_i2,n321_i3, n321_v);
  spice_node_5 n_n326(eclk, ereset, n326_i0,n326_i1,n326_i2,n326_i3,n326_i4, n326_v);
  spice_node_3 n_n327(eclk, ereset, n327_i0,n327_i1,n327_i2, n327_v);
  spice_node_2 n_op_inc_nop(eclk, ereset, op_inc_nop_i0,op_inc_nop_i1, op_inc_nop_v);
  spice_node_2 n_dpc1_SBY(eclk, ereset, dpc1_SBY_i2,dpc1_SBY_i9, dpc1_SBY_v);
  spice_node_2 n_ir0(eclk, ereset, ir0_i1,ir0_i2, ir0_v);
  spice_node_2 n_n329(eclk, ereset, n329_i0,n329_i2, n329_v);
  spice_node_3 n_ab2(eclk, ereset, ab2_i0,ab2_i1,ab2_i2, ab2_v);
  spice_node_3 n_n1594(eclk, ereset, n1594_i0,n1594_i1,n1594_i2, n1594_v);
  spice_node_5 n_n1592(eclk, ereset, n1592_i0,n1592_i1,n1592_i2,n1592_i3,n1592_i4, n1592_v);
  spice_node_2 n_n995(eclk, ereset, n995_i0,n995_i1, n995_v);
  spice_node_3 n_n994(eclk, ereset, n994_i1,n994_i2,n994_i3, n994_v);
  spice_node_2 n_abh6(eclk, ereset, abh6_i3,abh6_i4, abh6_v);
  spice_node_2 n_irline3(eclk, ereset, irline3_i0,irline3_i1, irline3_v);
  spice_node_8 n_idb1(eclk, ereset, idb1_i0,idb1_i2,idb1_i3,idb1_i4,idb1_i6,idb1_i7,idb1_i8,idb1_i9, idb1_v);
  spice_node_2 n_n990(eclk, ereset, n990_i0,n990_i3, n990_v);
  spice_node_1 n_n993(eclk, ereset, n993_i0, n993_v);
  spice_node_2 n_n992(eclk, ereset, n992_i0,n992_i1, n992_v);
  spice_node_3 n_n999(eclk, ereset, n999_i1,n999_i2,n999_i3, n999_v);
  spice_node_5 n_n998(eclk, ereset, n998_i0,n998_i1,n998_i2,n998_i3,n998_i4, n998_v);
  spice_node_2 n_op_T3(eclk, ereset, op_T3_i0,op_T3_i1, op_T3_v);
  spice_node_7 n_adl6(eclk, ereset, adl6_i1,adl6_i2,adl6_i3,adl6_i4,adl6_i5,adl6_i6,adl6_i7, adl6_v);
  spice_node_2 n_n122(eclk, ereset, n122_i0,n122_i1, n122_v);
  spice_node_3 n_n123(eclk, ereset, n123_i0,n123_i1,n123_i2, n123_v);
  spice_node_2 n_pchp3(eclk, ereset, pchp3_i0,pchp3_i2, pchp3_v);
  spice_node_2 n_PD_n_0xx0xx0x(eclk, ereset, PD_n_0xx0xx0x_i0,PD_n_0xx0xx0x_i1, PD_n_0xx0xx0x_v);
  spice_node_1 n_n126(eclk, ereset, n126_i1, n126_v);
  spice_node_2 n_n127(eclk, ereset, n127_i2,n127_i3, n127_v);
  spice_node_2 n_n128(eclk, ereset, n128_i0,n128_i2, n128_v);
  spice_node_2 n_dpc20_ADDSB06(eclk, ereset, dpc20_ADDSB06_i0,dpc20_ADDSB06_i5, dpc20_ADDSB06_v);
  spice_node_3 n_alub4(eclk, ereset, alub4_i0,alub4_i1,alub4_i2, alub4_v);
  spice_node_5 n_n1647(eclk, ereset, n1647_i0,n1647_i1,n1647_i2,n1647_i3,n1647_i4, n1647_v);
  spice_node_3 n_op_T__bit(eclk, ereset, op_T__bit_i0,op_T__bit_i1,op_T__bit_i2, op_T__bit_v);
  spice_node_3 n_n1641(eclk, ereset, n1641_i0,n1641_i1,n1641_i2, n1641_v);
  spice_node_2 n_n1640(eclk, ereset, n1640_i0,n1640_i2, n1640_v);
  spice_node_2 n_n1643(eclk, ereset, n1643_i0,n1643_i1, n1643_v);
  spice_node_2 n_n1642(eclk, ereset, n1642_i0,n1642_i2, n1642_v);
  spice_node_3 n_n1649(eclk, ereset, n1649_i1,n1649_i2,n1649_i3, n1649_v);
  spice_node_2 n_x3(eclk, ereset, x3_i0,x3_i1, x3_v);
  spice_node_1 n_n1252(eclk, ereset, n1252_i0, n1252_v);
  spice_node_2 n_op_T3_jsr(eclk, ereset, op_T3_jsr_i0,op_T3_jsr_i1, op_T3_jsr_v);
  spice_node_4 n_n578(eclk, ereset, n578_i0,n578_i1,n578_i2,n578_i3, n578_v);
  spice_node_3 n_n604(eclk, ereset, n604_i0,n604_i1,n604_i4, n604_v);
  spice_node_2 n_y2(eclk, ereset, y2_i0,y2_i2, y2_v);
  spice_node_2 n_n572(eclk, ereset, n572_i0,n572_i1, n572_v);
  spice_node_3 n_n571(eclk, ereset, n571_i0,n571_i1,n571_i2, n571_v);
  spice_node_2 n_n570(eclk, ereset, n570_i0,n570_i1, n570_v);
  spice_node_1 n_notidl1(eclk, ereset, notidl1_i0, notidl1_v);
  spice_node_2 n_op_T0_adc_sbc(eclk, ereset, op_T0_adc_sbc_i0,op_T0_adc_sbc_i1, op_T0_adc_sbc_v);
  spice_node_2 n_dpc15_ANDS(eclk, ereset, dpc15_ANDS_i0,dpc15_ANDS_i9, dpc15_ANDS_v);
  spice_node_3 n_n1209(eclk, ereset, n1209_i0,n1209_i1,n1209_i2, n1209_v);
  spice_node_3 n_Pout2(eclk, ereset, Pout2_i0,Pout2_i1,Pout2_i2, Pout2_v);
  spice_node_2 n_op_T0_lda(eclk, ereset, op_T0_lda_i1,op_T0_lda_i2, op_T0_lda_v);
  spice_node_2 n_n1423(eclk, ereset, n1423_i0,n1423_i3, n1423_v);
  spice_node_2 n__C34(eclk, ereset, _C34_i1,_C34_i3, _C34_v);
  spice_node_4 n_n1424(eclk, ereset, n1424_i0,n1424_i1,n1424_i2,n1424_i3, n1424_v);
  spice_node_2 n_n1427(eclk, ereset, n1427_i1,n1427_i2, n1427_v);
  spice_node_2 n_abh0(eclk, ereset, abh0_i3,abh0_i4, abh0_v);
  spice_node_2 n_op_T3_ind_x(eclk, ereset, op_T3_ind_x_i0,op_T3_ind_x_i1, op_T3_ind_x_v);
  spice_node_2 n_n602(eclk, ereset, n602_i0,n602_i1, n602_v);
  spice_node_2 n_pclp6(eclk, ereset, pclp6_i0,pclp6_i2, pclp6_v);
  spice_node_2 n_n730(eclk, ereset, n730_i1,n730_i2, n730_v);
  spice_node_4 n_n733(eclk, ereset, n733_i0,n733_i1,n733_i2,n733_i3, n733_v);
  spice_node_2 n_n732(eclk, ereset, n732_i0,n732_i3, n732_v);
  spice_node_2 n_n735(eclk, ereset, n735_i0,n735_i1, n735_v);
  spice_node_2 n_a0(eclk, ereset, a0_i0,a0_i1, a0_v);
  spice_node_3 n_ab5(eclk, ereset, ab5_i0,ab5_i1,ab5_i2, ab5_v);
  spice_node_2 n_n739(eclk, ereset, n739_i0,n739_i2, n739_v);
  spice_node_2 n_pcl3(eclk, ereset, pcl3_i1,pcl3_i2, pcl3_v);
  spice_node_3 n_n1358(eclk, ereset, n1358_i0,n1358_i2,n1358_i3, n1358_v);
  spice_node_1 n_n469(eclk, ereset, n469_i0, n469_v);
  spice_node_3 n_n468(eclk, ereset, n468_i0,n468_i1,n468_i2, n468_v);
  spice_node_3 n__WR(eclk, ereset, _WR_i0,_WR_i1,_WR_i2, _WR_v);
  spice_node_2 n_n467(eclk, ereset, n467_i0,n467_i3, n467_v);
  spice_node_2 n_n466(eclk, ereset, n466_i1,n466_i3, n466_v);
  spice_node_2 n_n1357(eclk, ereset, n1357_i0,n1357_i1, n1357_v);
  spice_node_2 n_n1356(eclk, ereset, n1356_i0,n1356_i2, n1356_v);
  spice_node_2 n_op_T0_cmp(eclk, ereset, op_T0_cmp_i0,op_T0_cmp_i1, op_T0_cmp_v);
  spice_node_3 n_n462(eclk, ereset, n462_i0,n462_i1,n462_i2, n462_v);
  spice_node_3 n_n1519(eclk, ereset, n1519_i0,n1519_i1,n1519_i2, n1519_v);
  spice_node_2 n_n1518(eclk, ereset, n1518_i0,n1518_i1, n1518_v);
  spice_node_2 n_n1517(eclk, ereset, n1517_i0,n1517_i1, n1517_v);
  spice_node_1 n_notidl4(eclk, ereset, notidl4_i0, notidl4_v);
  spice_node_2 n_n1511(eclk, ereset, n1511_i0,n1511_i1, n1511_v);
  spice_node_2 n__ABL5(eclk, ereset, _ABL5_i0,_ABL5_i2, _ABL5_v);
  spice_node_2 n_op_T2_abs_y(eclk, ereset, op_T2_abs_y_i0,op_T2_abs_y_i1, op_T2_abs_y_v);
  spice_node_1 n_pipeVectorA0(eclk, ereset, pipeVectorA0_i1, pipeVectorA0_v);
  spice_node_2 n_n355(eclk, ereset, n355_i0,n355_i3, n355_v);
  spice_node_2 n_op_T4_abs_idx(eclk, ereset, op_T4_abs_idx_i0,op_T4_abs_idx_i1, op_T4_abs_idx_v);
  spice_node_2 n_RnWstretched(eclk, ereset, RnWstretched_i0,RnWstretched_i1, RnWstretched_v);
  spice_node_2 n_op_T4_brk(eclk, ereset, op_T4_brk_i0,op_T4_brk_i1, op_T4_brk_v);
  spice_node_3 n_n351(eclk, ereset, n351_i0,n351_i1,n351_i2, n351_v);
  spice_node_4 n_n350(eclk, ereset, n350_i0,n350_i2,n350_i3,n350_i4, n350_v);
  spice_node_3 n_n359(eclk, ereset, n359_i0,n359_i1,n359_i2, n359_v);
  spice_node_2 n_n358(eclk, ereset, n358_i1,n358_i3, n358_v);
  spice_node_2 n_n1111(eclk, ereset, n1111_i0,n1111_i2, n1111_v);
  spice_node_3 n_n1110(eclk, ereset, n1110_i1,n1110_i2,n1110_i3, n1110_v);
  spice_node_1 n_n1113(eclk, ereset, n1113_i0, n1113_v);
  spice_node_2 n__ABH6(eclk, ereset, _ABH6_i1,_ABH6_i2, _ABH6_v);
  spice_node_2 n_n288(eclk, ereset, n288_i1,n288_i3, n288_v);
  spice_node_3 n_Pout1(eclk, ereset, Pout1_i0,Pout1_i1,Pout1_i2, Pout1_v);
  spice_node_2 n_op_T4_mem_abs_idx(eclk, ereset, op_T4_mem_abs_idx_i0,op_T4_mem_abs_idx_i2, op_T4_mem_abs_idx_v);
  spice_node_5 n_n280(eclk, ereset, n280_i0,n280_i1,n280_i2,n280_i3,n280_i4, n280_v);
  spice_node_2 n_dpc37_PCLDB(eclk, ereset, dpc37_PCLDB_i0,dpc37_PCLDB_i4, dpc37_PCLDB_v);
  spice_node_2 n_n282(eclk, ereset, n282_i0,n282_i1, n282_v);
  spice_node_2 n_op_T2_zp_zp_idx(eclk, ereset, op_T2_zp_zp_idx_i0,op_T2_zp_zp_idx_i2, op_T2_zp_zp_idx_v);
  spice_node_2 n_n284(eclk, ereset, n284_i0,n284_i1, n284_v);
  spice_node_2 n_abh2(eclk, ereset, abh2_i0,abh2_i4, abh2_v);
  spice_node_2 n_op_T0_tay_ldy_not_idx(eclk, ereset, op_T0_tay_ldy_not_idx_i0,op_T0_tay_ldy_not_idx_i1, op_T0_tay_ldy_not_idx_v);
  spice_node_2 n_n1441(eclk, ereset, n1441_i1,n1441_i2, n1441_v);
  spice_node_2 n_n1440(eclk, ereset, n1440_i0,n1440_i1, n1440_v);
  spice_node_3 n_dasb5(eclk, ereset, dasb5_i0,dasb5_i1,dasb5_i2, dasb5_v);
  spice_node_3 n_n262(eclk, ereset, n262_i0,n262_i1,n262_i2, n262_v);
  spice_node_3 n_n261(eclk, ereset, n261_i0,n261_i1,n261_i2, n261_v);
  spice_node_2 n_n260(eclk, ereset, n260_i0,n260_i1, n260_v);
  spice_node_2 n_n267(eclk, ereset, n267_i0,n267_i2, n267_v);
  spice_node_1 n_n266(eclk, ereset, n266_i0, n266_v);
  spice_node_1 n_n265(eclk, ereset, n265_i0, n265_v);
  spice_node_4 n_n264(eclk, ereset, n264_i0,n264_i1,n264_i2,n264_i3, n264_v);
  spice_node_2 n_n269(eclk, ereset, n269_i0,n269_i1, n269_v);
  spice_node_3 n_ab0(eclk, ereset, ab0_i0,ab0_i1,ab0_i2, ab0_v);
  spice_node_2 n_op_xy(eclk, ereset, op_xy_i1,op_xy_i2, op_xy_v);
  spice_node_1 n_n1291(eclk, ereset, n1291_i0, n1291_v);
  spice_node_2 n_n1296(eclk, ereset, n1296_i0,n1296_i2, n1296_v);
  spice_node_1 n_n1565(eclk, ereset, n1565_i1, n1565_v);
  spice_node_2 n_PD_1xx000x0(eclk, ereset, PD_1xx000x0_i0,PD_1xx000x0_i1, PD_1xx000x0_v);
  spice_node_2 n_n1295(eclk, ereset, n1295_i2,n1295_i3, n1295_v);
  spice_node_2 n_n988(eclk, ereset, n988_i0,n988_i1, n988_v);
  spice_node_2 n_y4(eclk, ereset, y4_i0,y4_i2, y4_v);
  spice_node_1 n_n982(eclk, ereset, n982_i1, n982_v);
  spice_node_3 n_n983(eclk, ereset, n983_i0,n983_i1,n983_i2, n983_v);
  spice_node_2 n_n980(eclk, ereset, n980_i0,n980_i1, n980_v);
  spice_node_2 n_n981(eclk, ereset, n981_i1,n981_i2, n981_v);
  spice_node_2 n_n986(eclk, ereset, n986_i0,n986_i1, n986_v);
  spice_node_2 n_n987(eclk, ereset, n987_i1,n987_i2, n987_v);
  spice_node_2 n_dpc12_0ADD(eclk, ereset, dpc12_0ADD_i7,dpc12_0ADD_i9, dpc12_0ADD_v);
  spice_node_2 n_op_T0_ldx_tax_tsx(eclk, ereset, op_T0_ldx_tax_tsx_i0,op_T0_ldx_tax_tsx_i1, op_T0_ldx_tax_tsx_v);
  spice_node_2 n_y6(eclk, ereset, y6_i0,y6_i1, y6_v);
  spice_node_1 n_pchp2(eclk, ereset, pchp2_i1, pchp2_v);
  spice_node_2 n_A_B7(eclk, ereset, A_B7_i0,A_B7_i1, A_B7_v);
  spice_node_1 n_notidl0(eclk, ereset, notidl0_i0, notidl0_v);
  spice_node_3 n_n111(eclk, ereset, n111_i0,n111_i1,n111_i2, n111_v);
  spice_node_2 n_n110(eclk, ereset, n110_i0,n110_i1, n110_v);
  spice_node_2 n_pchp1(eclk, ereset, pchp1_i0,pchp1_i2, pchp1_v);
  spice_node_2 n_n119(eclk, ereset, n119_i0,n119_i2, n119_v);
  spice_node_2 n_n118(eclk, ereset, n118_i0,n118_i1, n118_v);
  spice_node_2 n__DBE(eclk, ereset, _DBE_i0,_DBE_i1, _DBE_v);
  spice_node_7 n_adl5(eclk, ereset, adl5_i0,adl5_i1,adl5_i2,adl5_i3,adl5_i4,adl5_i5,adl5_i7, adl5_v);
  spice_node_3 n_n1631(eclk, ereset, n1631_i0,n1631_i1,n1631_i2, n1631_v);
  spice_node_3 n_n1632(eclk, ereset, n1632_i1,n1632_i2,n1632_i4, n1632_v);
  spice_node_2 n_n1633(eclk, ereset, n1633_i0,n1633_i2, n1633_v);
  spice_node_2 n_dor2(eclk, ereset, dor2_i1,dor2_i2, dor2_v);
  spice_node_2 n_n1635(eclk, ereset, n1635_i1,n1635_i2, n1635_v);
  spice_node_4 n_alu2(eclk, ereset, alu2_i0,alu2_i1,alu2_i3,alu2_i4, alu2_v);
  spice_node_3 n_n1638(eclk, ereset, n1638_i0,n1638_i1,n1638_i2, n1638_v);
  spice_node_2 n_n1639(eclk, ereset, n1639_i0,n1639_i2, n1639_v);
  spice_node_3 n_n568(eclk, ereset, n568_i0,n568_i1,n568_i2, n568_v);
  spice_node_1 n_C78_phi2(eclk, ereset, C78_phi2_i0, C78_phi2_v);
  spice_node_1 n_pipeUNK22(eclk, ereset, pipeUNK22_i0, pipeUNK22_v);
  spice_node_1 n_n562(eclk, ereset, n562_i0, n562_v);
  spice_node_4 n_n564(eclk, ereset, n564_i0,n564_i1,n564_i2,n564_i3, n564_v);
  spice_node_2 n_n565(eclk, ereset, n565_i0,n565_i2, n565_v);
  spice_node_3 n_n566(eclk, ereset, n566_i0,n566_i1,n566_i2, n566_v);
  spice_node_2 n_n567(eclk, ereset, n567_i0,n567_i4, n567_v);
  spice_node_12 n_sb3(eclk, ereset, sb3_i0,sb3_i1,sb3_i2,sb3_i3,sb3_i4,sb3_i5,sb3_i6,sb3_i7,sb3_i8,sb3_i9,sb3_i10,sb3_i11, sb3_v);
  spice_node_2 n_dpc3_SBX(eclk, ereset, dpc3_SBX_i8,dpc3_SBX_i9, dpc3_SBX_v);
  spice_node_3 n_n1187(eclk, ereset, n1187_i0,n1187_i1,n1187_i2, n1187_v);
  spice_node_2 n_n1184(eclk, ereset, n1184_i0,n1184_i3, n1184_v);
  spice_node_2 n_short_circuit_idx_add(eclk, ereset, short_circuit_idx_add_i0,short_circuit_idx_add_i1, short_circuit_idx_add_v);
  spice_node_3 n_notir2(eclk, ereset, notir2_i0,notir2_i1,notir2_i2, notir2_v);
  spice_node_3 n_n1180(eclk, ereset, n1180_i0,n1180_i1,n1180_i2, n1180_v);
  spice_node_3 n_n1181(eclk, ereset, n1181_i0,n1181_i1,n1181_i2, n1181_v);
  spice_node_2 n_n726(eclk, ereset, n726_i1,n726_i2, n726_v);
  spice_node_2 n_a4(eclk, ereset, a4_i0,a4_i2, a4_v);
  spice_node_2 n_dpc22__DSA(eclk, ereset, dpc22__DSA_i0,dpc22__DSA_i2, dpc22__DSA_v);
  spice_node_6 n_n722(eclk, ereset, n722_i0,n722_i1,n722_i2,n722_i3,n722_i4,n722_i5, n722_v);
  spice_node_5 n_n723(eclk, ereset, n723_i0,n723_i1,n723_i2,n723_i3,n723_i4, n723_v);
  spice_node_3 n_n720(eclk, ereset, n720_i0,n720_i1,n720_i2, n720_v);
  spice_node_5 n_n721(eclk, ereset, n721_i0,n721_i1,n721_i2,n721_i3,n721_i4, n721_v);
  spice_node_3 n_n728(eclk, ereset, n728_i0,n728_i1,n728_i2, n728_v);
  spice_node_1 n_pipeUNK36(eclk, ereset, pipeUNK36_i0, pipeUNK36_v);
  spice_node_2 n_op_clv(eclk, ereset, op_clv_i1,op_clv_i2, op_clv_v);
  spice_node_2 n_notalucin(eclk, ereset, notalucin_i1,notalucin_i2, notalucin_v);
  spice_node_2 n_n1166(eclk, ereset, n1166_i0,n1166_i1, n1166_v);
  spice_node_2 n_alua0(eclk, ereset, alua0_i0,alua0_i1, alua0_v);
  spice_node_6 n_adh4(eclk, ereset, adh4_i0,adh4_i1,adh4_i2,adh4_i4,adh4_i5,adh4_i6, adh4_v);
  spice_node_1 n_n1161(eclk, ereset, n1161_i0, n1161_v);
  spice_node_1 n_n1162(eclk, ereset, n1162_i0, n1162_v);
  spice_node_3 n_clk1out(eclk, ereset, clk1out_i0,clk1out_i1,clk1out_i2, clk1out_v);
  spice_node_2 n_op_T5_ind_y(eclk, ereset, op_T5_ind_y_i0,op_T5_ind_y_i1, op_T5_ind_y_v);
  spice_node_4 n_n1169(eclk, ereset, n1169_i0,n1169_i1,n1169_i2,n1169_i3, n1169_v);
  spice_node_2 n_dpc30_ADHPCH(eclk, ereset, dpc30_ADHPCH_i8,dpc30_ADHPCH_i9, dpc30_ADHPCH_v);
  spice_node_2 n_pch5(eclk, ereset, pch5_i0,pch5_i2, pch5_v);
  spice_node_2 n_n46(eclk, ereset, n46_i0,n46_i1, n46_v);
  spice_node_1 n_n47(eclk, ereset, n47_i1, n47_v);
  spice_node_1 n_pipeUNK05(eclk, ereset, pipeUNK05_i0, pipeUNK05_v);
  spice_node_1 n_pipeVectorA2(eclk, ereset, pipeVectorA2_i1, pipeVectorA2_v);
  spice_node_2 n_n42(eclk, ereset, n42_i0,n42_i2, n42_v);
  spice_node_2 n_n43(eclk, ereset, n43_i0,n43_i1, n43_v);
  spice_node_1 n_pipeT2out(eclk, ereset, pipeT2out_i0, pipeT2out_v);
  spice_node_2 n_dpc42_DL_ADH(eclk, ereset, dpc42_DL_ADH_i8,dpc42_DL_ADH_i9, dpc42_DL_ADH_v);
  spice_node_2 n_x_op_T4_rti(eclk, ereset, x_op_T4_rti_i0,x_op_T4_rti_i1, x_op_T4_rti_v);
  spice_node_7 n_adl7(eclk, ereset, adl7_i0,adl7_i2,adl7_i3,adl7_i4,adl7_i5,adl7_i6,adl7_i7, adl7_v);
  spice_node_2 n_op_T0_cli_sei(eclk, ereset, op_T0_cli_sei_i1,op_T0_cli_sei_i2, op_T0_cli_sei_v);
  spice_node_2 n_n1561(eclk, ereset, n1561_i0,n1561_i2, n1561_v);
  spice_node_3 n_n1290(eclk, ereset, n1290_i0,n1290_i1,n1290_i2, n1290_v);
  spice_node_2 n_dpc41_DL_ADL(eclk, ereset, dpc41_DL_ADL_i0,dpc41_DL_ADL_i9, dpc41_DL_ADL_v);
  spice_node_1 n_nmi(eclk, ereset, nmi_i1, nmi_v);
  spice_node_2 n_n1566(eclk, ereset, n1566_i0,n1566_i3, n1566_v);
  spice_node_2 n_t3(eclk, ereset, t3_i1,t3_i2, t3_v);
  spice_node_1 n_pipeUNK35(eclk, ereset, pipeUNK35_i0, pipeUNK35_v);
  spice_node_3 n_n474(eclk, ereset, n474_i0,n474_i1,n474_i2, n474_v);
  spice_node_3 n_n1712(eclk, ereset, n1712_i0,n1712_i1,n1712_i2, n1712_v);
  spice_node_3 n_n1711(eclk, ereset, n1711_i0,n1711_i1,n1711_i2, n1711_v);
  spice_node_2 n_op_T__cpx_cpy_imm_zp(eclk, ereset, op_T__cpx_cpy_imm_zp_i0,op_T__cpx_cpy_imm_zp_i1, op_T__cpx_cpy_imm_zp_v);
  spice_node_1 n__TWOCYCLE_phi1(eclk, ereset, _TWOCYCLE_phi1_i0, _TWOCYCLE_phi1_v);
  spice_node_2 n_n1715(eclk, ereset, n1715_i2,n1715_i3, n1715_v);
  spice_node_2 n_dpc18__DAA(eclk, ereset, dpc18__DAA_i0,dpc18__DAA_i1, dpc18__DAA_v);
  spice_node_2 n_n1714(eclk, ereset, n1714_i0,n1714_i1, n1714_v);
  spice_node_3 n_n472(eclk, ereset, n472_i0,n472_i1,n472_i2, n472_v);
  spice_node_2 n_n470(eclk, ereset, n470_i0,n470_i1, n470_v);
  spice_node_2 n_n471(eclk, ereset, n471_i1,n471_i2, n471_v);
  spice_node_2 n_n476(eclk, ereset, n476_i2,n476_i3, n476_v);
  spice_node_4 n_n477(eclk, ereset, n477_i0,n477_i2,n477_i3,n477_i4, n477_v);
  spice_node_1 n_n1360(eclk, ereset, n1360_i0, n1360_v);
  spice_node_2 n_n475(eclk, ereset, n475_i0,n475_i2, n475_v);
  spice_node_3 n_n478(eclk, ereset, n478_i0,n478_i1,n478_i2, n478_v);
  spice_node_2 n_n479(eclk, ereset, n479_i0,n479_i1, n479_v);
  spice_node_3 n_n1368(eclk, ereset, n1368_i0,n1368_i1,n1368_i2, n1368_v);
  spice_node_2 n_n1369(eclk, ereset, n1369_i2,n1369_i3, n1369_v);

endmodule
