* SPICE3 file created from 4001.ext - technology: nmos

.option scale=1u

M1000 clk2 GND GND GND efet w=241 l=16
+ ad=39724 pd=3842 as=1.32121e+06 ps=97808 
M1001 clk1 GND GND GND efet w=241 l=16
+ ad=26307 pd=2800 as=0 ps=0 
M1002 d2 GND d2 GND efet w=443 l=275
+ ad=94881 pd=7472 as=0 ps=0 
M1003 d3 GND d3 GND efet w=448 l=283
+ ad=120243 pd=10236 as=0 ps=0 
M1004 sync GND GND GND efet w=226 l=16
+ ad=59770 pd=6506 as=0 ps=0 
M1005 GND diff_847_4156# d3 GND efet w=2335 l=8
+ ad=0 pd=0 as=0 ps=0 
M1006 GND diff_1237_4156# d2 GND efet w=2332 l=8
+ ad=0 pd=0 as=0 ps=0 
M1007 Vdd diff_889_3418# d3 GND efet w=1075 l=23
+ ad=423648 pd=37992 as=0 ps=0 
M1008 GND diff_1624_4156# d1 GND efet w=2332 l=8
+ ad=0 pd=0 as=94236 ps=7574 
M1009 GND diff_2011_4156# d0 GND efet w=2332 l=8
+ ad=0 pd=0 as=93441 ps=7526 
M1010 GND diff_6085_4357# diff_6094_4246# GND efet w=889 l=13
+ ad=0 pd=0 as=59323 ps=3682 
M1011 GND clk1 diff_6535_4298# GND efet w=61 l=16
+ ad=0 pd=0 as=2729 ps=228 
M1012 GND sync diff_6085_4357# GND efet w=190 l=16
+ ad=0 pd=0 as=17550 ps=1502 
M1013 diff_7004_4333# diff_6880_4216# GND GND efet w=67 l=13
+ ad=3020 pd=456 as=0 ps=0 
M1014 diff_6625_3571# diff_7004_4333# GND GND efet w=100 l=13
+ ad=4496 pd=510 as=0 ps=0 
M1015 diff_6535_4298# Vdd Vdd GND efet w=16 l=22
+ ad=0 pd=0 as=0 ps=0 
M1016 GND diff_2509_4258# diff_2521_4214# GND efet w=1546 l=16
+ ad=0 pd=0 as=123880 ps=7204 
M1017 Vdd diff_4144_4258# diff_2521_4214# GND efet w=1606 l=16
+ ad=0 pd=0 as=0 ps=0 
M1018 diff_2521_4214# diff_2512_4201# diff_2521_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1019 diff_2521_4214# diff_2512_4201# diff_2572_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1020 diff_2521_4214# diff_2512_4201# diff_2623_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1021 diff_2521_4214# diff_2512_4201# diff_2674_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1022 diff_2521_4214# diff_2512_4201# diff_2725_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1023 diff_2521_4214# diff_2512_4201# diff_2776_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1024 diff_2521_4214# diff_2512_4201# diff_2827_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1025 diff_2521_4214# diff_2512_4201# diff_2878_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1026 diff_2521_4214# diff_2512_4201# diff_2929_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1027 diff_2521_4214# diff_2512_4201# diff_2980_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1028 diff_2521_4214# diff_2512_4201# diff_3031_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1029 diff_2521_4214# diff_2512_4201# diff_3082_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1030 diff_2521_4214# diff_2512_4201# diff_3133_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1031 diff_2521_4214# diff_2512_4201# diff_3184_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1032 diff_2521_4214# diff_2512_4201# diff_3235_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1033 diff_2521_4214# diff_2512_4201# diff_3286_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1034 diff_2521_4214# diff_2512_4201# diff_3337_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1035 diff_2521_4214# diff_2512_4201# diff_3388_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1036 diff_2521_4214# diff_2512_4201# diff_3439_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1037 diff_2521_4214# diff_2512_4201# diff_3490_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1038 diff_2521_4214# diff_2512_4201# diff_3541_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1039 diff_2521_4214# diff_2512_4201# diff_3592_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1040 diff_2521_4214# diff_2512_4201# diff_3643_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1041 diff_2521_4214# diff_2512_4201# diff_3694_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1042 diff_2521_4214# diff_2512_4201# diff_3745_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1043 diff_2521_4214# diff_2512_4201# diff_3796_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1044 diff_2521_4214# diff_2512_4201# diff_3847_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1045 diff_2521_4214# diff_2512_4201# diff_3898_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1046 diff_2521_4214# diff_2512_4201# diff_3949_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1047 diff_2521_4214# diff_2512_4201# diff_4000_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1048 diff_2521_4214# diff_2512_4201# diff_4051_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1049 diff_2521_4214# diff_2512_4201# diff_4102_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1050 diff_2521_4214# diff_2512_4201# diff_4153_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1051 diff_2521_4214# diff_2512_4201# diff_4204_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1052 diff_2521_4214# diff_2512_4201# diff_4255_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1053 diff_2521_4214# diff_2512_4201# diff_4306_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1054 diff_2521_4214# diff_2512_4201# diff_4357_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1055 diff_2521_4214# diff_2512_4201# diff_4408_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1056 diff_2521_4214# diff_2512_4201# diff_4459_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1057 diff_2521_4214# diff_2512_4201# diff_4510_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1058 diff_2521_4214# diff_2512_4201# diff_4561_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1059 diff_2521_4214# diff_2512_4201# diff_4612_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1060 diff_2521_4214# diff_2512_4201# diff_4663_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1061 diff_2521_4214# diff_2512_4201# diff_4714_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1062 diff_2521_4214# diff_2512_4201# diff_4765_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1063 diff_2521_4214# diff_2512_4201# diff_4816_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1064 diff_2521_4214# diff_2512_4201# diff_4867_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1065 diff_2521_4214# diff_2512_4201# diff_4918_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1066 diff_2521_4214# diff_2512_4201# diff_4969_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1067 diff_2521_4214# diff_2512_4201# diff_5020_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1068 diff_2521_4214# diff_2512_4201# diff_5071_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1069 diff_2521_4214# diff_2512_4201# diff_5122_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1070 diff_2521_4214# diff_2512_4201# diff_5173_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1071 diff_2521_4214# diff_2512_4201# diff_5224_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1072 diff_2521_4214# diff_2512_4201# diff_5275_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1073 diff_2521_4214# diff_2512_4201# diff_5326_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1074 diff_2521_4214# diff_2512_4201# diff_5377_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1075 diff_2521_4214# diff_2512_4201# diff_5428_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1076 diff_2521_4214# diff_2512_4201# diff_5479_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1077 diff_2521_4214# diff_2512_4201# diff_5530_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1078 diff_2521_4214# diff_2512_4201# diff_5581_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1079 diff_2521_4214# diff_2512_4201# diff_5632_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1080 diff_2521_4214# diff_2512_4201# diff_5683_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1081 diff_2521_4214# diff_2512_4201# diff_5734_4157# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1082 diff_5918_4184# diff_5905_1069# diff_2512_4201# GND efet w=221 l=16
+ ad=23284 pd=1722 as=5882 ps=576 
M1083 Vdd Vdd diff_916_3763# GND efet w=22 l=22
+ ad=0 pd=0 as=1471 ps=176 
M1084 Vdd Vdd diff_1072_3769# GND efet w=19 l=25
+ ad=0 pd=0 as=1166 ps=164 
M1085 Vdd diff_1276_3418# d2 GND efet w=1071 l=25
+ ad=0 pd=0 as=0 ps=0 
M1086 diff_916_3763# diff_916_3763# diff_916_3763# GND efet w=3 l=7
+ ad=0 pd=0 as=0 ps=0 
M1087 Vdd diff_916_3763# diff_889_3418# GND efet w=19 l=16
+ ad=0 pd=0 as=19135 ps=1622 
M1088 Vdd diff_1072_3769# diff_847_4156# GND efet w=19 l=16
+ ad=0 pd=0 as=23632 ps=1916 
M1089 diff_1072_3769# diff_1072_3769# diff_1072_3769# GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M1090 diff_916_3763# diff_916_3763# diff_916_3763# GND efet w=2 l=6
+ ad=0 pd=0 as=0 ps=0 
M1091 diff_889_3418# diff_916_3763# diff_889_3418# GND efet w=103 l=33
+ ad=0 pd=0 as=0 ps=0 
M1092 diff_1072_3769# diff_1072_3769# diff_1072_3769# GND efet w=3 l=13
+ ad=0 pd=0 as=0 ps=0 
M1093 Vdd Vdd diff_1303_3760# GND efet w=16 l=22
+ ad=0 pd=0 as=1232 ps=178 
M1094 Vdd Vdd diff_1459_3766# GND efet w=22 l=25
+ ad=0 pd=0 as=1327 ps=190 
M1095 diff_1303_3760# diff_1303_3760# diff_1303_3760# GND efet w=4 l=5
+ ad=0 pd=0 as=0 ps=0 
M1096 Vdd diff_1303_3760# diff_1276_3418# GND efet w=19 l=16
+ ad=0 pd=0 as=19156 ps=1622 
M1097 Vdd diff_1459_3766# diff_1237_4156# GND efet w=19 l=16
+ ad=0 pd=0 as=24019 ps=1922 
M1098 diff_1459_3766# diff_1459_3766# diff_1459_3766# GND efet w=7 l=8
+ ad=0 pd=0 as=0 ps=0 
M1099 diff_1303_3760# diff_1303_3760# diff_1303_3760# GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M1100 diff_847_4156# diff_1072_3769# diff_847_4156# GND efet w=139 l=15
+ ad=0 pd=0 as=0 ps=0 
M1101 diff_1276_3418# diff_1303_3760# diff_1276_3418# GND efet w=106 l=33
+ ad=0 pd=0 as=0 ps=0 
M1102 diff_1459_3766# diff_1459_3766# diff_1459_3766# GND efet w=2 l=15
+ ad=0 pd=0 as=0 ps=0 
M1103 Vdd diff_1663_3415# d1 GND efet w=1075 l=16
+ ad=0 pd=0 as=0 ps=0 
M1104 Vdd Vdd diff_1684_3766# GND efet w=19 l=25
+ ad=0 pd=0 as=1051 ps=154 
M1105 Vdd Vdd diff_1846_3766# GND efet w=19 l=25
+ ad=0 pd=0 as=1105 ps=152 
M1106 Vdd diff_2053_3415# d0 GND efet w=1068 l=23
+ ad=0 pd=0 as=0 ps=0 
M1107 Vdd diff_1684_3766# diff_1663_3415# GND efet w=16 l=16
+ ad=0 pd=0 as=19396 ps=1736 
M1108 diff_1684_3766# diff_1684_3766# diff_1684_3766# GND efet w=4 l=10
+ ad=0 pd=0 as=0 ps=0 
M1109 diff_1237_4156# diff_1459_3766# diff_1237_4156# GND efet w=139 l=15
+ ad=0 pd=0 as=0 ps=0 
M1110 Vdd diff_1846_3766# diff_1624_4156# GND efet w=17 l=17
+ ad=0 pd=0 as=23389 ps=1910 
M1111 diff_1846_3766# diff_1846_3766# diff_1846_3766# GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M1112 diff_1684_3766# diff_1684_3766# diff_1684_3766# GND efet w=2 l=9
+ ad=0 pd=0 as=0 ps=0 
M1113 diff_1846_3766# diff_1846_3766# diff_1846_3766# GND efet w=0 l=1
+ ad=0 pd=0 as=0 ps=0 
M1114 Vdd Vdd diff_2080_3763# GND efet w=19 l=22
+ ad=0 pd=0 as=1249 ps=164 
M1115 Vdd Vdd diff_2218_3868# GND efet w=19 l=22
+ ad=0 pd=0 as=1030 ps=146 
M1116 diff_2521_4157# diff_2512_4144# diff_2521_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1117 diff_2572_4157# diff_2512_4144# diff_2572_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1118 diff_2623_4157# diff_2512_4144# diff_2623_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1119 diff_2674_4157# diff_2512_4144# diff_2674_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1120 diff_2725_4157# diff_2512_4144# diff_2725_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1121 diff_2776_4157# diff_2512_4144# diff_2776_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1122 diff_2827_4157# diff_2512_4144# diff_2827_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1123 diff_2878_4157# diff_2512_4144# diff_2878_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1124 diff_2929_4157# diff_2512_4144# diff_2929_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1125 diff_2980_4157# diff_2512_4144# diff_2980_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1126 diff_3031_4157# diff_2512_4144# diff_3031_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1127 diff_3082_4157# diff_2512_4144# diff_3082_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1128 diff_3133_4157# diff_2512_4144# diff_3133_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1129 diff_3184_4157# diff_2512_4144# diff_3184_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1130 diff_3235_4157# diff_2512_4144# diff_3235_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1131 diff_3286_4157# diff_2512_4144# diff_3286_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1132 diff_3337_4157# diff_2512_4144# diff_3337_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1133 diff_3388_4157# diff_2512_4144# diff_3388_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1134 diff_3439_4157# diff_2512_4144# diff_3439_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1135 diff_3490_4157# diff_2512_4144# diff_3490_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1136 diff_3541_4157# diff_2512_4144# diff_3541_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1137 diff_3592_4157# diff_2512_4144# diff_3592_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1138 diff_3643_4157# diff_2512_4144# diff_3643_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1139 diff_3694_4157# diff_2512_4144# diff_3694_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1140 diff_3745_4157# diff_2512_4144# diff_3745_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1141 diff_3796_4157# diff_2512_4144# diff_3796_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1142 diff_3847_4157# diff_2512_4144# diff_3847_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1143 diff_3898_4157# diff_2512_4144# diff_3898_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1144 diff_3949_4157# diff_2512_4144# diff_3949_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1145 diff_4000_4157# diff_2512_4144# diff_4000_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1146 diff_4051_4157# diff_2512_4144# diff_4051_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1147 diff_4102_4157# diff_2512_4144# diff_4102_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1148 diff_4153_4157# diff_2512_4144# diff_4153_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1149 diff_4204_4157# diff_2512_4144# diff_4204_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1150 diff_4255_4157# diff_2512_4144# diff_4255_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1151 diff_4306_4157# diff_2512_4144# diff_4306_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1152 diff_4357_4157# diff_2512_4144# diff_4357_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1153 diff_4408_4157# diff_2512_4144# diff_4408_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1154 diff_4459_4157# diff_2512_4144# diff_4459_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1155 diff_4510_4157# diff_2512_4144# diff_4510_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1156 diff_4561_4157# diff_2512_4144# diff_4561_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1157 diff_4612_4157# diff_2512_4144# diff_4612_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1158 diff_4663_4157# diff_2512_4144# diff_4663_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1159 diff_4714_4157# diff_2512_4144# diff_4714_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1160 diff_4765_4157# diff_2512_4144# diff_4765_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1161 diff_4816_4157# diff_2512_4144# diff_4816_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1162 diff_4867_4157# diff_2512_4144# diff_4867_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1163 diff_4918_4157# diff_2512_4144# diff_4918_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1164 diff_4969_4157# diff_2512_4144# diff_4969_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1165 diff_5020_4157# diff_2512_4144# diff_5020_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1166 diff_5071_4157# diff_2512_4144# diff_5071_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1167 diff_5122_4157# diff_2512_4144# diff_5122_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1168 diff_5173_4157# diff_2512_4144# diff_5173_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1169 diff_5224_4157# diff_2512_4144# diff_5224_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1170 diff_5275_4157# diff_2512_4144# diff_5275_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1171 diff_5326_4157# diff_2512_4144# diff_5326_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1172 diff_5377_4157# diff_2512_4144# diff_5377_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1173 diff_5428_4157# diff_2512_4144# diff_5428_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1174 diff_5479_4157# diff_2512_4144# diff_5479_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1175 diff_5530_4157# diff_2512_4144# diff_5530_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1176 diff_5581_4157# diff_2512_4144# diff_5581_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1177 diff_5632_4157# diff_2512_4144# diff_5632_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1178 diff_5683_4157# diff_2512_4144# diff_5683_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1179 diff_5734_4157# diff_2512_4144# diff_5734_4103# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1180 diff_2512_4201# Vdd Vdd GND efet w=13 l=28
+ ad=0 pd=0 as=0 ps=0 
M1181 diff_2521_4103# diff_2512_4090# diff_2521_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1182 diff_2572_4103# diff_2512_4090# diff_2572_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1183 diff_2623_4103# diff_2512_4090# diff_2623_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1184 diff_2674_4103# diff_2512_4090# diff_2674_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1185 diff_2725_4103# diff_2512_4090# diff_2725_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1186 diff_2776_4103# diff_2512_4090# diff_2776_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1187 diff_2827_4103# diff_2512_4090# diff_2827_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1188 diff_2878_4103# diff_2512_4090# diff_2878_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1189 diff_2929_4103# diff_2512_4090# diff_2929_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1190 diff_2980_4103# diff_2512_4090# diff_2980_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1191 diff_3031_4103# diff_2512_4090# diff_3031_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1192 diff_3082_4103# diff_2512_4090# diff_3082_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1193 diff_3133_4103# diff_2512_4090# diff_3133_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1194 diff_3184_4103# diff_2512_4090# diff_3184_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1195 diff_3235_4103# diff_2512_4090# diff_3235_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1196 diff_3286_4103# diff_2512_4090# diff_3286_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1197 diff_3337_4103# diff_2512_4090# diff_3337_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1198 diff_3388_4103# diff_2512_4090# diff_3388_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1199 diff_3439_4103# diff_2512_4090# diff_3439_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1200 diff_3490_4103# diff_2512_4090# diff_3490_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1201 diff_3541_4103# diff_2512_4090# diff_3541_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1202 diff_3592_4103# diff_2512_4090# diff_3592_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1203 diff_3643_4103# diff_2512_4090# diff_3643_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1204 diff_3694_4103# diff_2512_4090# diff_3694_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1205 diff_3745_4103# diff_2512_4090# diff_3745_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1206 diff_3796_4103# diff_2512_4090# diff_3796_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1207 diff_3847_4103# diff_2512_4090# diff_3847_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1208 diff_3898_4103# diff_2512_4090# diff_3898_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1209 diff_3949_4103# diff_2512_4090# diff_3949_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1210 diff_4000_4103# diff_2512_4090# diff_4000_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1211 diff_4051_4103# diff_2512_4090# diff_4051_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1212 diff_4102_4103# diff_2512_4090# diff_4102_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1213 diff_4153_4103# diff_2512_4090# diff_4153_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1214 diff_4204_4103# diff_2512_4090# diff_4204_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1215 diff_4255_4103# diff_2512_4090# diff_4255_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1216 diff_4306_4103# diff_2512_4090# diff_4306_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1217 diff_4357_4103# diff_2512_4090# diff_4357_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1218 diff_4408_4103# diff_2512_4090# diff_4408_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1219 diff_4459_4103# diff_2512_4090# diff_4459_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1220 diff_4510_4103# diff_2512_4090# diff_4510_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1221 diff_4561_4103# diff_2512_4090# diff_4561_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1222 diff_4612_4103# diff_2512_4090# diff_4612_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1223 diff_4663_4103# diff_2512_4090# diff_4663_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1224 diff_4714_4103# diff_2512_4090# diff_4714_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1225 diff_4765_4103# diff_2512_4090# diff_4765_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1226 diff_4816_4103# diff_2512_4090# diff_4816_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1227 diff_4867_4103# diff_2512_4090# diff_4867_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1228 diff_4918_4103# diff_2512_4090# diff_4918_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1229 diff_4969_4103# diff_2512_4090# diff_4969_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1230 diff_5020_4103# diff_2512_4090# diff_5020_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1231 diff_5071_4103# diff_2512_4090# diff_5071_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1232 diff_5122_4103# diff_2512_4090# diff_5122_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1233 diff_5173_4103# diff_2512_4090# diff_5173_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1234 diff_5224_4103# diff_2512_4090# diff_5224_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1235 diff_5275_4103# diff_2512_4090# diff_5275_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1236 diff_5326_4103# diff_2512_4090# diff_5326_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1237 diff_5377_4103# diff_2512_4090# diff_5377_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1238 diff_5428_4103# diff_2512_4090# diff_5428_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1239 diff_5479_4103# diff_2512_4090# diff_5479_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1240 diff_5530_4103# diff_2512_4090# diff_5530_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1241 diff_5581_4103# diff_2512_4090# diff_5581_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1242 diff_5632_4103# diff_2512_4090# diff_5632_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1243 diff_5683_4103# diff_2512_4090# diff_5683_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1244 diff_5734_4103# diff_2512_4090# diff_5734_4046# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1245 Vdd Vdd diff_2512_4033# GND efet w=13 l=28
+ ad=0 pd=0 as=5073 ps=640 
M1246 diff_2521_4046# diff_2512_4033# diff_2521_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1247 diff_2572_4046# diff_2512_4033# diff_2572_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1248 diff_2623_4046# diff_2512_4033# diff_2623_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1249 diff_2674_4046# diff_2512_4033# diff_2674_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1250 diff_2725_4046# diff_2512_4033# diff_2725_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1251 diff_2776_4046# diff_2512_4033# diff_2776_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1252 diff_2827_4046# diff_2512_4033# diff_2827_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1253 diff_2878_4046# diff_2512_4033# diff_2878_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1254 diff_2929_4046# diff_2512_4033# diff_2929_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1255 diff_2980_4046# diff_2512_4033# diff_2980_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1256 diff_3031_4046# diff_2512_4033# diff_3031_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1257 diff_3082_4046# diff_2512_4033# diff_3082_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1258 diff_3133_4046# diff_2512_4033# diff_3133_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1259 diff_3184_4046# diff_2512_4033# diff_3184_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1260 diff_3235_4046# diff_2512_4033# diff_3235_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1261 diff_3286_4046# diff_2512_4033# diff_3286_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1262 diff_3337_4046# diff_2512_4033# diff_3337_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1263 diff_3388_4046# diff_2512_4033# diff_3388_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1264 diff_3439_4046# diff_2512_4033# diff_3439_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1265 diff_3490_4046# diff_2512_4033# diff_3490_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1266 diff_3541_4046# diff_2512_4033# diff_3541_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1267 diff_3592_4046# diff_2512_4033# diff_3592_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1268 diff_3643_4046# diff_2512_4033# diff_3643_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1269 diff_3694_4046# diff_2512_4033# diff_3694_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1270 diff_3745_4046# diff_2512_4033# diff_3745_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1271 diff_3796_4046# diff_2512_4033# diff_3796_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1272 diff_3847_4046# diff_2512_4033# diff_3847_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1273 diff_3898_4046# diff_2512_4033# diff_3898_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1274 diff_3949_4046# diff_2512_4033# diff_3949_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1275 diff_4000_4046# diff_2512_4033# diff_4000_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1276 diff_4051_4046# diff_2512_4033# diff_4051_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1277 diff_4102_4046# diff_2512_4033# diff_4102_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1278 diff_4153_4046# diff_2512_4033# diff_4153_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1279 diff_4204_4046# diff_2512_4033# diff_4204_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1280 diff_4255_4046# diff_2512_4033# diff_4255_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1281 diff_4306_4046# diff_2512_4033# diff_4306_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1282 diff_4357_4046# diff_2512_4033# diff_4357_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1283 diff_4408_4046# diff_2512_4033# diff_4408_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1284 diff_4459_4046# diff_2512_4033# diff_4459_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1285 diff_4510_4046# diff_2512_4033# diff_4510_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1286 diff_4561_4046# diff_2512_4033# diff_4561_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1287 diff_4612_4046# diff_2512_4033# diff_4612_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1288 diff_4663_4046# diff_2512_4033# diff_4663_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1289 diff_4714_4046# diff_2512_4033# diff_4714_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1290 diff_4765_4046# diff_2512_4033# diff_4765_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1291 diff_4816_4046# diff_2512_4033# diff_4816_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1292 diff_4867_4046# diff_2512_4033# diff_4867_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1293 diff_4918_4046# diff_2512_4033# diff_4918_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1294 diff_4969_4046# diff_2512_4033# diff_4969_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1295 diff_5020_4046# diff_2512_4033# diff_5020_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1296 diff_5071_4046# diff_2512_4033# diff_5071_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1297 diff_5122_4046# diff_2512_4033# diff_5122_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1298 diff_5173_4046# diff_2512_4033# diff_5173_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1299 diff_5224_4046# diff_2512_4033# diff_5224_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1300 diff_5275_4046# diff_2512_4033# diff_5275_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1301 diff_5326_4046# diff_2512_4033# diff_5326_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1302 diff_5377_4046# diff_2512_4033# diff_5377_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1303 diff_5428_4046# diff_2512_4033# diff_5428_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1304 diff_5479_4046# diff_2512_4033# diff_5479_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1305 diff_5530_4046# diff_2512_4033# diff_5530_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1306 diff_5581_4046# diff_2512_4033# diff_5581_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1307 diff_5632_4046# diff_2512_4033# diff_5632_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1308 diff_5683_4046# diff_2512_4033# diff_5683_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1309 diff_5734_4046# diff_2512_4033# diff_5734_3992# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1310 diff_2512_4033# diff_5962_1069# diff_5918_4184# GND efet w=184 l=13
+ ad=0 pd=0 as=0 ps=0 
M1311 diff_5918_4184# diff_6034_2491# diff_2512_4144# GND efet w=205 l=16
+ ad=0 pd=0 as=6638 ps=558 
M1312 diff_2512_4144# Vdd Vdd GND efet w=16 l=28
+ ad=0 pd=0 as=0 ps=0 
M1313 Vdd Vdd diff_2512_4090# GND efet w=16 l=28
+ ad=0 pd=0 as=5700 ps=610 
M1314 diff_2521_3992# diff_2512_3979# diff_2521_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1315 diff_2572_3992# diff_2512_3979# diff_2572_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1316 diff_2623_3992# diff_2512_3979# diff_2623_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1317 diff_2674_3992# diff_2512_3979# diff_2674_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1318 diff_2725_3992# diff_2512_3979# diff_2725_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1319 diff_2776_3992# diff_2512_3979# diff_2776_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1320 diff_2827_3992# diff_2512_3979# diff_2827_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1321 diff_2878_3992# diff_2512_3979# diff_2878_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1322 diff_2929_3992# diff_2512_3979# diff_2929_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1323 diff_2980_3992# diff_2512_3979# diff_2980_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1324 diff_3031_3992# diff_2512_3979# diff_3031_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1325 diff_3082_3992# diff_2512_3979# diff_3082_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1326 diff_3133_3992# diff_2512_3979# diff_3133_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1327 diff_3184_3992# diff_2512_3979# diff_3184_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1328 diff_3235_3992# diff_2512_3979# diff_3235_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1329 diff_3286_3992# diff_2512_3979# diff_3286_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1330 diff_3337_3992# diff_2512_3979# diff_3337_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1331 diff_3388_3992# diff_2512_3979# diff_3388_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1332 diff_3439_3992# diff_2512_3979# diff_3439_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1333 diff_3490_3992# diff_2512_3979# diff_3490_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1334 diff_3541_3992# diff_2512_3979# diff_3541_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1335 diff_3592_3992# diff_2512_3979# diff_3592_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1336 diff_3643_3992# diff_2512_3979# diff_3643_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1337 diff_3694_3992# diff_2512_3979# diff_3694_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1338 diff_3745_3992# diff_2512_3979# diff_3745_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1339 diff_3796_3992# diff_2512_3979# diff_3796_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1340 diff_3847_3992# diff_2512_3979# diff_3847_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1341 diff_3898_3992# diff_2512_3979# diff_3898_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1342 diff_3949_3992# diff_2512_3979# diff_3949_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1343 diff_4000_3992# diff_2512_3979# diff_4000_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1344 diff_4051_3992# diff_2512_3979# diff_4051_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1345 diff_4102_3992# diff_2512_3979# diff_4102_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1346 diff_4153_3992# diff_2512_3979# diff_4153_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1347 diff_4204_3992# diff_2512_3979# diff_4204_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1348 diff_4255_3992# diff_2512_3979# diff_4255_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1349 diff_4306_3992# diff_2512_3979# diff_4306_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1350 diff_4357_3992# diff_2512_3979# diff_4357_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1351 diff_4408_3992# diff_2512_3979# diff_4408_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1352 diff_4459_3992# diff_2512_3979# diff_4459_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1353 diff_4510_3992# diff_2512_3979# diff_4510_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1354 diff_4561_3992# diff_2512_3979# diff_4561_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1355 diff_4612_3992# diff_2512_3979# diff_4612_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1356 diff_4663_3992# diff_2512_3979# diff_4663_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1357 diff_4714_3992# diff_2512_3979# diff_4714_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1358 diff_4765_3992# diff_2512_3979# diff_4765_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1359 diff_4816_3992# diff_2512_3979# diff_4816_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1360 diff_4867_3992# diff_2512_3979# diff_4867_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1361 diff_4918_3992# diff_2512_3979# diff_4918_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1362 diff_4969_3992# diff_2512_3979# diff_4969_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1363 diff_5020_3992# diff_2512_3979# diff_5020_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1364 diff_5071_3992# diff_2512_3979# diff_5071_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1365 diff_5122_3992# diff_2512_3979# diff_5122_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1366 diff_5173_3992# diff_2512_3979# diff_5173_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1367 diff_5224_3992# diff_2512_3979# diff_5224_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1368 diff_5275_3992# diff_2512_3979# diff_5275_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1369 diff_5326_3992# diff_2512_3979# diff_5326_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1370 diff_5377_3992# diff_2512_3979# diff_5377_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1371 diff_5428_3992# diff_2512_3979# diff_5428_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1372 diff_5479_3992# diff_2512_3979# diff_5479_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1373 diff_5530_3992# diff_2512_3979# diff_5530_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1374 diff_5581_3992# diff_2512_3979# diff_5581_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1375 diff_5632_3992# diff_2512_3979# diff_5632_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1376 diff_5683_3992# diff_2512_3979# diff_5683_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1377 diff_5734_3992# diff_2512_3979# diff_5734_3935# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1378 diff_5918_3962# diff_5905_1069# diff_2512_3979# GND efet w=217 l=14
+ ad=24457 pd=1826 as=5462 ps=564 
M1379 diff_2512_4090# diff_6079_2449# diff_5918_4184# GND efet w=196 l=13
+ ad=0 pd=0 as=0 ps=0 
M1380 diff_2521_3935# diff_2512_3922# diff_2521_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1381 diff_2572_3935# diff_2512_3922# diff_2572_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1382 diff_2623_3935# diff_2512_3922# diff_2623_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1383 diff_2674_3935# diff_2512_3922# diff_2674_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1384 diff_2725_3935# diff_2512_3922# diff_2725_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1385 diff_2776_3935# diff_2512_3922# diff_2776_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1386 diff_2827_3935# diff_2512_3922# diff_2827_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1387 diff_2878_3935# diff_2512_3922# diff_2878_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1388 diff_2929_3935# diff_2512_3922# diff_2929_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1389 diff_2980_3935# diff_2512_3922# diff_2980_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1390 diff_3031_3935# diff_2512_3922# diff_3031_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1391 diff_3082_3935# diff_2512_3922# diff_3082_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1392 diff_3133_3935# diff_2512_3922# diff_3133_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1393 diff_3184_3935# diff_2512_3922# diff_3184_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1394 diff_3235_3935# diff_2512_3922# diff_3235_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1395 diff_3286_3935# diff_2512_3922# diff_3286_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1396 diff_3337_3935# diff_2512_3922# diff_3337_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1397 diff_3388_3935# diff_2512_3922# diff_3388_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1398 diff_3439_3935# diff_2512_3922# diff_3439_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1399 diff_3490_3935# diff_2512_3922# diff_3490_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1400 diff_3541_3935# diff_2512_3922# diff_3541_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1401 diff_3592_3935# diff_2512_3922# diff_3592_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1402 diff_3643_3935# diff_2512_3922# diff_3643_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1403 diff_3694_3935# diff_2512_3922# diff_3694_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1404 diff_3745_3935# diff_2512_3922# diff_3745_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1405 diff_3796_3935# diff_2512_3922# diff_3796_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1406 diff_3847_3935# diff_2512_3922# diff_3847_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1407 diff_3898_3935# diff_2512_3922# diff_3898_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1408 diff_3949_3935# diff_2512_3922# diff_3949_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1409 diff_4000_3935# diff_2512_3922# diff_4000_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1410 diff_4051_3935# diff_2512_3922# diff_4051_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1411 diff_4102_3935# diff_2512_3922# diff_4102_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1412 diff_4153_3935# diff_2512_3922# diff_4153_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1413 diff_4204_3935# diff_2512_3922# diff_4204_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1414 diff_4255_3935# diff_2512_3922# diff_4255_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1415 diff_4306_3935# diff_2512_3922# diff_4306_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1416 diff_4357_3935# diff_2512_3922# diff_4357_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1417 diff_4408_3935# diff_2512_3922# diff_4408_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1418 diff_4459_3935# diff_2512_3922# diff_4459_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1419 diff_4510_3935# diff_2512_3922# diff_4510_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1420 diff_4561_3935# diff_2512_3922# diff_4561_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1421 diff_4612_3935# diff_2512_3922# diff_4612_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1422 diff_4663_3935# diff_2512_3922# diff_4663_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1423 diff_4714_3935# diff_2512_3922# diff_4714_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1424 diff_4765_3935# diff_2512_3922# diff_4765_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1425 diff_4816_3935# diff_2512_3922# diff_4816_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1426 diff_4867_3935# diff_2512_3922# diff_4867_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1427 diff_4918_3935# diff_2512_3922# diff_4918_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1428 diff_4969_3935# diff_2512_3922# diff_4969_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1429 diff_5020_3935# diff_2512_3922# diff_5020_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1430 diff_5071_3935# diff_2512_3922# diff_5071_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1431 diff_5122_3935# diff_2512_3922# diff_5122_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1432 diff_5173_3935# diff_2512_3922# diff_5173_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1433 diff_5224_3935# diff_2512_3922# diff_5224_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1434 diff_5275_3935# diff_2512_3922# diff_5275_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1435 diff_5326_3935# diff_2512_3922# diff_5326_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1436 diff_5377_3935# diff_2512_3922# diff_5377_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1437 diff_5428_3935# diff_2512_3922# diff_5428_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1438 diff_5479_3935# diff_2512_3922# diff_5479_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1439 diff_5530_3935# diff_2512_3922# diff_5530_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1440 diff_5581_3935# diff_2512_3922# diff_5581_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1441 diff_5632_3935# diff_2512_3922# diff_5632_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1442 diff_5683_3935# diff_2512_3922# diff_5683_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1443 diff_5734_3935# diff_2512_3922# diff_5734_3881# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1444 diff_2080_3763# diff_2080_3763# diff_2080_3763# GND efet w=0 l=1
+ ad=0 pd=0 as=0 ps=0 
M1445 Vdd diff_2080_3763# diff_2053_3415# GND efet w=16 l=16
+ ad=0 pd=0 as=19261 ps=1616 
M1446 Vdd diff_2218_3868# diff_2011_4156# GND efet w=16 l=16
+ ad=0 pd=0 as=23767 ps=1868 
M1447 diff_2218_3868# diff_2218_3868# diff_2218_3868# GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M1448 diff_2080_3763# diff_2080_3763# diff_2080_3763# GND efet w=0 l=1
+ ad=0 pd=0 as=0 ps=0 
M1449 diff_889_3418# diff_847_4156# GND GND efet w=241 l=16
+ ad=0 pd=0 as=0 ps=0 
M1450 diff_847_4156# diff_1021_3622# GND GND efet w=466 l=16
+ ad=0 pd=0 as=0 ps=0 
M1451 diff_1663_3415# diff_1684_3766# diff_1663_3415# GND efet w=150 l=8
+ ad=0 pd=0 as=0 ps=0 
M1452 diff_1624_4156# diff_1846_3766# diff_1624_4156# GND efet w=139 l=18
+ ad=0 pd=0 as=0 ps=0 
M1453 GND diff_475_2011# diff_889_3418# GND efet w=472 l=16
+ ad=0 pd=0 as=0 ps=0 
M1454 diff_1276_3418# diff_1237_4156# GND GND efet w=241 l=16
+ ad=0 pd=0 as=0 ps=0 
M1455 diff_1237_4156# diff_1408_3622# GND GND efet w=469 l=16
+ ad=0 pd=0 as=0 ps=0 
M1456 diff_2053_3415# diff_2080_3763# diff_2053_3415# GND efet w=103 l=33
+ ad=0 pd=0 as=0 ps=0 
M1457 diff_2218_3868# diff_2218_3868# diff_2218_3868# GND efet w=0 l=1
+ ad=0 pd=0 as=0 ps=0 
M1458 diff_2512_3979# Vdd Vdd GND efet w=13 l=31
+ ad=0 pd=0 as=0 ps=0 
M1459 diff_2521_3881# diff_2512_3868# diff_2521_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1460 diff_2572_3881# diff_2512_3868# diff_2572_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1461 diff_2623_3881# diff_2512_3868# diff_2623_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1462 diff_2674_3881# diff_2512_3868# diff_2674_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1463 diff_2725_3881# diff_2512_3868# diff_2725_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1464 diff_2776_3881# diff_2512_3868# diff_2776_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1465 diff_2827_3881# diff_2512_3868# diff_2827_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1466 diff_2878_3881# diff_2512_3868# diff_2878_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1467 diff_2929_3881# diff_2512_3868# diff_2929_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1468 diff_2980_3881# diff_2512_3868# diff_2980_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1469 diff_3031_3881# diff_2512_3868# diff_3031_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1470 diff_3082_3881# diff_2512_3868# diff_3082_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1471 diff_3133_3881# diff_2512_3868# diff_3133_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1472 diff_3184_3881# diff_2512_3868# diff_3184_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1473 diff_3235_3881# diff_2512_3868# diff_3235_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1474 diff_3286_3881# diff_2512_3868# diff_3286_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1475 diff_3337_3881# diff_2512_3868# diff_3337_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1476 diff_3388_3881# diff_2512_3868# diff_3388_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1477 diff_3439_3881# diff_2512_3868# diff_3439_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1478 diff_3490_3881# diff_2512_3868# diff_3490_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1479 diff_3541_3881# diff_2512_3868# diff_3541_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1480 diff_3592_3881# diff_2512_3868# diff_3592_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1481 diff_3643_3881# diff_2512_3868# diff_3643_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1482 diff_3694_3881# diff_2512_3868# diff_3694_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1483 diff_3745_3881# diff_2512_3868# diff_3745_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1484 diff_3796_3881# diff_2512_3868# diff_3796_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1485 diff_3847_3881# diff_2512_3868# diff_3847_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1486 diff_3898_3881# diff_2512_3868# diff_3898_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1487 diff_3949_3881# diff_2512_3868# diff_3949_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1488 diff_4000_3881# diff_2512_3868# diff_4000_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1489 diff_4051_3881# diff_2512_3868# diff_4051_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1490 diff_4102_3881# diff_2512_3868# diff_4102_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1491 diff_4153_3881# diff_2512_3868# diff_4153_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1492 diff_4204_3881# diff_2512_3868# diff_4204_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1493 diff_4255_3881# diff_2512_3868# diff_4255_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1494 diff_4306_3881# diff_2512_3868# diff_4306_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1495 diff_4357_3881# diff_2512_3868# diff_4357_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1496 diff_4408_3881# diff_2512_3868# diff_4408_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1497 diff_4459_3881# diff_2512_3868# diff_4459_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1498 diff_4510_3881# diff_2512_3868# diff_4510_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1499 diff_4561_3881# diff_2512_3868# diff_4561_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1500 diff_4612_3881# diff_2512_3868# diff_4612_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1501 diff_4663_3881# diff_2512_3868# diff_4663_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1502 diff_4714_3881# diff_2512_3868# diff_4714_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1503 diff_4765_3881# diff_2512_3868# diff_4765_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1504 diff_4816_3881# diff_2512_3868# diff_4816_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1505 diff_4867_3881# diff_2512_3868# diff_4867_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1506 diff_4918_3881# diff_2512_3868# diff_4918_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1507 diff_4969_3881# diff_2512_3868# diff_4969_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1508 diff_5020_3881# diff_2512_3868# diff_5020_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1509 diff_5071_3881# diff_2512_3868# diff_5071_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1510 diff_5122_3881# diff_2512_3868# diff_5122_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1511 diff_5173_3881# diff_2512_3868# diff_5173_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1512 diff_5224_3881# diff_2512_3868# diff_5224_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1513 diff_5275_3881# diff_2512_3868# diff_5275_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1514 diff_5326_3881# diff_2512_3868# diff_5326_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1515 diff_5377_3881# diff_2512_3868# diff_5377_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1516 diff_5428_3881# diff_2512_3868# diff_5428_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1517 diff_5479_3881# diff_2512_3868# diff_5479_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1518 diff_5530_3881# diff_2512_3868# diff_5530_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1519 diff_5581_3881# diff_2512_3868# diff_5581_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1520 diff_5632_3881# diff_2512_3868# diff_5632_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1521 diff_5683_3881# diff_2512_3868# diff_5683_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1522 diff_5734_3881# diff_2512_3868# diff_5734_3824# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1523 diff_2011_4156# diff_2218_3868# diff_2011_4156# GND efet w=123 l=24
+ ad=0 pd=0 as=0 ps=0 
M1524 Vdd Vdd diff_2512_3811# GND efet w=13 l=31
+ ad=0 pd=0 as=5073 ps=640 
M1525 diff_2521_3824# diff_2512_3811# diff_2521_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1526 diff_2572_3824# diff_2512_3811# diff_2572_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1527 diff_2623_3824# diff_2512_3811# diff_2623_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1528 diff_2674_3824# diff_2512_3811# diff_2674_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1529 diff_2725_3824# diff_2512_3811# diff_2725_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1530 diff_2776_3824# diff_2512_3811# diff_2776_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1531 diff_2827_3824# diff_2512_3811# diff_2827_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1532 diff_2878_3824# diff_2512_3811# diff_2878_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1533 diff_2929_3824# diff_2512_3811# diff_2929_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1534 diff_2980_3824# diff_2512_3811# diff_2980_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1535 diff_3031_3824# diff_2512_3811# diff_3031_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1536 diff_3082_3824# diff_2512_3811# diff_3082_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1537 diff_3133_3824# diff_2512_3811# diff_3133_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1538 diff_3184_3824# diff_2512_3811# diff_3184_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1539 diff_3235_3824# diff_2512_3811# diff_3235_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1540 diff_3286_3824# diff_2512_3811# diff_3286_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1541 diff_3337_3824# diff_2512_3811# diff_3337_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1542 diff_3388_3824# diff_2512_3811# diff_3388_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1543 diff_3439_3824# diff_2512_3811# diff_3439_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1544 diff_3490_3824# diff_2512_3811# diff_3490_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1545 diff_3541_3824# diff_2512_3811# diff_3541_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1546 diff_3592_3824# diff_2512_3811# diff_3592_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1547 diff_3643_3824# diff_2512_3811# diff_3643_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1548 diff_3694_3824# diff_2512_3811# diff_3694_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1549 diff_3745_3824# diff_2512_3811# diff_3745_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1550 diff_3796_3824# diff_2512_3811# diff_3796_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1551 diff_3847_3824# diff_2512_3811# diff_3847_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1552 diff_3898_3824# diff_2512_3811# diff_3898_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1553 diff_3949_3824# diff_2512_3811# diff_3949_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1554 diff_4000_3824# diff_2512_3811# diff_4000_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1555 diff_4051_3824# diff_2512_3811# diff_4051_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1556 diff_4102_3824# diff_2512_3811# diff_4102_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1557 diff_4153_3824# diff_2512_3811# diff_4153_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1558 diff_4204_3824# diff_2512_3811# diff_4204_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1559 diff_4255_3824# diff_2512_3811# diff_4255_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1560 diff_4306_3824# diff_2512_3811# diff_4306_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1561 diff_4357_3824# diff_2512_3811# diff_4357_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1562 diff_4408_3824# diff_2512_3811# diff_4408_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1563 diff_4459_3824# diff_2512_3811# diff_4459_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1564 diff_4510_3824# diff_2512_3811# diff_4510_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1565 diff_4561_3824# diff_2512_3811# diff_4561_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1566 diff_4612_3824# diff_2512_3811# diff_4612_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1567 diff_4663_3824# diff_2512_3811# diff_4663_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1568 diff_4714_3824# diff_2512_3811# diff_4714_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1569 diff_4765_3824# diff_2512_3811# diff_4765_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1570 diff_4816_3824# diff_2512_3811# diff_4816_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1571 diff_4867_3824# diff_2512_3811# diff_4867_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1572 diff_4918_3824# diff_2512_3811# diff_4918_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1573 diff_4969_3824# diff_2512_3811# diff_4969_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1574 diff_5020_3824# diff_2512_3811# diff_5020_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1575 diff_5071_3824# diff_2512_3811# diff_5071_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1576 diff_5122_3824# diff_2512_3811# diff_5122_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1577 diff_5173_3824# diff_2512_3811# diff_5173_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1578 diff_5224_3824# diff_2512_3811# diff_5224_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1579 diff_5275_3824# diff_2512_3811# diff_5275_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1580 diff_5326_3824# diff_2512_3811# diff_5326_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1581 diff_5377_3824# diff_2512_3811# diff_5377_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1582 diff_5428_3824# diff_2512_3811# diff_5428_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1583 diff_5479_3824# diff_2512_3811# diff_5479_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1584 diff_5530_3824# diff_2512_3811# diff_5530_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1585 diff_5581_3824# diff_2512_3811# diff_5581_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1586 diff_5632_3824# diff_2512_3811# diff_5632_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1587 diff_5683_3824# diff_2512_3811# diff_5683_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1588 diff_5734_3824# diff_2512_3811# diff_5734_3770# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1589 diff_2512_3811# diff_5962_1069# diff_5918_3962# GND efet w=184 l=13
+ ad=0 pd=0 as=0 ps=0 
M1590 diff_5918_3962# diff_6034_2491# diff_2512_3922# GND efet w=209 l=14
+ ad=0 pd=0 as=6920 ps=558 
M1591 diff_2512_3922# Vdd Vdd GND efet w=16 l=34
+ ad=0 pd=0 as=0 ps=0 
M1592 Vdd Vdd diff_2512_3868# GND efet w=16 l=31
+ ad=0 pd=0 as=5700 ps=610 
M1593 diff_2521_3770# diff_2512_3757# diff_2521_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1594 diff_2572_3770# diff_2512_3757# diff_2572_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1595 diff_2623_3770# diff_2512_3757# diff_2623_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1596 diff_2674_3770# diff_2512_3757# diff_2674_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1597 diff_2725_3770# diff_2512_3757# diff_2725_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1598 diff_2776_3770# diff_2512_3757# diff_2776_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1599 diff_2827_3770# diff_2512_3757# diff_2827_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1600 diff_2878_3770# diff_2512_3757# diff_2878_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1601 diff_2929_3770# diff_2512_3757# diff_2929_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1602 diff_2980_3770# diff_2512_3757# diff_2980_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1603 diff_3031_3770# diff_2512_3757# diff_3031_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1604 diff_3082_3770# diff_2512_3757# diff_3082_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1605 diff_3133_3770# diff_2512_3757# diff_3133_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1606 diff_3184_3770# diff_2512_3757# diff_3184_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1607 diff_3235_3770# diff_2512_3757# diff_3235_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1608 diff_3286_3770# diff_2512_3757# diff_3286_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1609 diff_3337_3770# diff_2512_3757# diff_3337_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1610 diff_3388_3770# diff_2512_3757# diff_3388_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1611 diff_3439_3770# diff_2512_3757# diff_3439_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1612 diff_3490_3770# diff_2512_3757# diff_3490_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1613 diff_3541_3770# diff_2512_3757# diff_3541_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1614 diff_3592_3770# diff_2512_3757# diff_3592_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1615 diff_3643_3770# diff_2512_3757# diff_3643_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1616 diff_3694_3770# diff_2512_3757# diff_3694_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1617 diff_3745_3770# diff_2512_3757# diff_3745_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1618 diff_3796_3770# diff_2512_3757# diff_3796_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1619 diff_3847_3770# diff_2512_3757# diff_3847_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1620 diff_3898_3770# diff_2512_3757# diff_3898_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1621 diff_3949_3770# diff_2512_3757# diff_3949_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1622 diff_4000_3770# diff_2512_3757# diff_4000_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1623 diff_4051_3770# diff_2512_3757# diff_4051_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1624 diff_4102_3770# diff_2512_3757# diff_4102_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1625 diff_4153_3770# diff_2512_3757# diff_4153_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1626 diff_4204_3770# diff_2512_3757# diff_4204_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1627 diff_4255_3770# diff_2512_3757# diff_4255_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1628 diff_4306_3770# diff_2512_3757# diff_4306_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1629 diff_4357_3770# diff_2512_3757# diff_4357_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1630 diff_4408_3770# diff_2512_3757# diff_4408_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1631 diff_4459_3770# diff_2512_3757# diff_4459_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1632 diff_4510_3770# diff_2512_3757# diff_4510_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1633 diff_4561_3770# diff_2512_3757# diff_4561_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1634 diff_4612_3770# diff_2512_3757# diff_4612_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1635 diff_4663_3770# diff_2512_3757# diff_4663_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1636 diff_4714_3770# diff_2512_3757# diff_4714_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1637 diff_4765_3770# diff_2512_3757# diff_4765_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1638 diff_4816_3770# diff_2512_3757# diff_4816_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1639 diff_4867_3770# diff_2512_3757# diff_4867_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1640 diff_4918_3770# diff_2512_3757# diff_4918_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1641 diff_4969_3770# diff_2512_3757# diff_4969_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1642 diff_5020_3770# diff_2512_3757# diff_5020_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1643 diff_5071_3770# diff_2512_3757# diff_5071_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1644 diff_5122_3770# diff_2512_3757# diff_5122_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1645 diff_5173_3770# diff_2512_3757# diff_5173_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1646 diff_5224_3770# diff_2512_3757# diff_5224_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1647 diff_5275_3770# diff_2512_3757# diff_5275_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1648 diff_5326_3770# diff_2512_3757# diff_5326_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1649 diff_5377_3770# diff_2512_3757# diff_5377_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1650 diff_5428_3770# diff_2512_3757# diff_5428_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1651 diff_5479_3770# diff_2512_3757# diff_5479_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1652 diff_5530_3770# diff_2512_3757# diff_5530_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1653 diff_5581_3770# diff_2512_3757# diff_5581_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1654 diff_5632_3770# diff_2512_3757# diff_5632_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1655 diff_5683_3770# diff_2512_3757# diff_5683_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1656 diff_5734_3770# diff_2512_3757# diff_5734_3713# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1657 diff_847_4156# diff_475_2011# GND GND efet w=475 l=16
+ ad=0 pd=0 as=0 ps=0 
M1658 GND diff_475_2011# diff_1276_3418# GND efet w=472 l=16
+ ad=0 pd=0 as=0 ps=0 
M1659 diff_1663_3415# diff_1624_4156# GND GND efet w=241 l=16
+ ad=0 pd=0 as=0 ps=0 
M1660 diff_1624_4156# diff_1798_3622# GND GND efet w=469 l=16
+ ad=0 pd=0 as=0 ps=0 
M1661 diff_1237_4156# diff_475_2011# GND GND efet w=475 l=16
+ ad=0 pd=0 as=0 ps=0 
M1662 GND diff_475_2011# diff_1663_3415# GND efet w=475 l=16
+ ad=0 pd=0 as=0 ps=0 
M1663 diff_2053_3415# diff_2011_4156# GND GND efet w=241 l=16
+ ad=0 pd=0 as=0 ps=0 
M1664 diff_2011_4156# diff_2185_3622# GND GND efet w=469 l=16
+ ad=0 pd=0 as=0 ps=0 
M1665 diff_5918_3734# diff_5905_1069# diff_2512_3757# GND efet w=218 l=16
+ ad=24730 pd=1790 as=5786 ps=576 
M1666 diff_2512_3868# diff_6079_2449# diff_5918_3962# GND efet w=196 l=13
+ ad=0 pd=0 as=0 ps=0 
M1667 diff_6094_4246# diff_6223_2134# diff_5918_3962# GND efet w=385 l=16
+ ad=0 pd=0 as=0 ps=0 
M1668 diff_5918_4184# diff_6265_2299# diff_6094_4246# GND efet w=400 l=16
+ ad=0 pd=0 as=0 ps=0 
M1669 GND diff_6085_4357# diff_6859_4286# GND efet w=100 l=13
+ ad=0 pd=0 as=2600 ps=252 
M1670 diff_6085_4357# diff_6661_4216# GND GND efet w=115 l=16
+ ad=0 pd=0 as=0 ps=0 
M1671 diff_6085_4357# Vdd Vdd GND efet w=16 l=34
+ ad=0 pd=0 as=0 ps=0 
M1672 diff_6880_4216# diff_6880_4216# diff_6880_4216# GND efet w=2 l=2
+ ad=5055 pd=582 as=0 ps=0 
M1673 diff_6859_4286# diff_6661_3556# diff_6859_4258# GND efet w=100 l=13
+ ad=0 pd=0 as=2846 ps=300 
M1674 diff_6880_4216# diff_6880_4216# diff_6880_4216# GND efet w=0 l=1
+ ad=0 pd=0 as=0 ps=0 
M1675 GND diff_6706_4228# diff_6661_4216# GND efet w=55 l=13
+ ad=0 pd=0 as=4342 ps=532 
M1676 diff_6859_4258# diff_6625_3799# diff_6880_4216# GND efet w=103 l=13
+ ad=0 pd=0 as=0 ps=0 
M1677 diff_6661_4216# diff_6661_4216# diff_6661_4216# GND efet w=1 l=1
+ ad=0 pd=0 as=0 ps=0 
M1678 GND d3 diff_7072_2716# GND efet w=403 l=13
+ ad=0 pd=0 as=11408 ps=884 
M1679 diff_6661_4216# Vdd Vdd GND efet w=14 l=94
+ ad=0 pd=0 as=0 ps=0 
M1680 diff_6706_4228# diff_6706_4228# diff_6706_4228# GND efet w=3 l=7
+ ad=880 pd=122 as=0 ps=0 
M1681 Vdd Vdd Vdd GND efet w=0 l=1
+ ad=0 pd=0 as=0 ps=0 
M1682 Vdd Vdd Vdd GND efet w=1 l=3
+ ad=0 pd=0 as=0 ps=0 
M1683 diff_6706_4228# diff_6706_4228# diff_6706_4228# GND efet w=2 l=5
+ ad=0 pd=0 as=0 ps=0 
M1684 Vdd Vdd diff_6880_4216# GND efet w=16 l=79
+ ad=0 pd=0 as=0 ps=0 
M1685 diff_7004_4333# Vdd Vdd GND efet w=13 l=52
+ ad=0 pd=0 as=0 ps=0 
M1686 diff_6625_3571# Vdd Vdd GND efet w=16 l=28
+ ad=0 pd=0 as=0 ps=0 
M1687 diff_7072_2716# Vdd Vdd GND efet w=22 l=37
+ ad=0 pd=0 as=0 ps=0 
M1688 diff_6706_4228# diff_6535_4298# diff_6778_3391# GND efet w=28 l=16
+ ad=0 pd=0 as=9433 ps=902 
M1689 diff_7072_3184# Vdd Vdd GND efet w=22 l=37
+ ad=7286 pd=492 as=0 ps=0 
M1690 GND diff_7072_2716# diff_7072_3184# GND efet w=112 l=13
+ ad=0 pd=0 as=0 ps=0 
M1691 diff_6661_4216# diff_6625_3799# GND GND efet w=37 l=13
+ ad=0 pd=0 as=0 ps=0 
M1692 sync clk2 diff_6919_3958# GND efet w=28 l=13
+ ad=0 pd=0 as=904 ps=124 
M1693 diff_6919_3958# diff_6919_3958# diff_6919_3958# GND efet w=1 l=1
+ ad=0 pd=0 as=0 ps=0 
M1694 diff_6919_3958# diff_6919_3958# diff_6919_3958# GND efet w=0 l=1
+ ad=0 pd=0 as=0 ps=0 
M1695 GND diff_6625_3799# diff_4144_4258# GND efet w=733 l=13
+ ad=0 pd=0 as=32121 ps=2638 
M1696 diff_4144_4258# diff_6479_3832# diff_4144_4258# GND efet w=135 l=41
+ ad=0 pd=0 as=0 ps=0 
M1697 diff_4144_4258# diff_6479_3832# Vdd GND efet w=37 l=13
+ ad=0 pd=0 as=0 ps=0 
M1698 diff_1624_4156# diff_475_2011# GND GND efet w=472 l=16
+ ad=0 pd=0 as=0 ps=0 
M1699 GND diff_475_2011# diff_2053_3415# GND efet w=472 l=16
+ ad=0 pd=0 as=0 ps=0 
M1700 diff_2521_3713# diff_2512_3700# diff_2521_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1701 diff_2572_3713# diff_2512_3700# diff_2572_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1702 diff_2623_3713# diff_2512_3700# diff_2623_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1703 diff_2674_3713# diff_2512_3700# diff_2674_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1704 diff_2725_3713# diff_2512_3700# diff_2725_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1705 diff_2776_3713# diff_2512_3700# diff_2776_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1706 diff_2827_3713# diff_2512_3700# diff_2827_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1707 diff_2878_3713# diff_2512_3700# diff_2878_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1708 diff_2929_3713# diff_2512_3700# diff_2929_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1709 diff_2980_3713# diff_2512_3700# diff_2980_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1710 diff_3031_3713# diff_2512_3700# diff_3031_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1711 diff_3082_3713# diff_2512_3700# diff_3082_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1712 diff_3133_3713# diff_2512_3700# diff_3133_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1713 diff_3184_3713# diff_2512_3700# diff_3184_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1714 diff_3235_3713# diff_2512_3700# diff_3235_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1715 diff_3286_3713# diff_2512_3700# diff_3286_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1716 diff_3337_3713# diff_2512_3700# diff_3337_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1717 diff_3388_3713# diff_2512_3700# diff_3388_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1718 diff_3439_3713# diff_2512_3700# diff_3439_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1719 diff_3490_3713# diff_2512_3700# diff_3490_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1720 diff_3541_3713# diff_2512_3700# diff_3541_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1721 diff_3592_3713# diff_2512_3700# diff_3592_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1722 diff_3643_3713# diff_2512_3700# diff_3643_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1723 diff_3694_3713# diff_2512_3700# diff_3694_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1724 diff_3745_3713# diff_2512_3700# diff_3745_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1725 diff_3796_3713# diff_2512_3700# diff_3796_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1726 diff_3847_3713# diff_2512_3700# diff_3847_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1727 diff_3898_3713# diff_2512_3700# diff_3898_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1728 diff_3949_3713# diff_2512_3700# diff_3949_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1729 diff_4000_3713# diff_2512_3700# diff_4000_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1730 diff_4051_3713# diff_2512_3700# diff_4051_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1731 diff_4102_3713# diff_2512_3700# diff_4102_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1732 diff_4153_3713# diff_2512_3700# diff_4153_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1733 diff_4204_3713# diff_2512_3700# diff_4204_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1734 diff_4255_3713# diff_2512_3700# diff_4255_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1735 diff_4306_3713# diff_2512_3700# diff_4306_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1736 diff_4357_3713# diff_2512_3700# diff_4357_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1737 diff_4408_3713# diff_2512_3700# diff_4408_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1738 diff_4459_3713# diff_2512_3700# diff_4459_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1739 diff_4510_3713# diff_2512_3700# diff_4510_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1740 diff_4561_3713# diff_2512_3700# diff_4561_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1741 diff_4612_3713# diff_2512_3700# diff_4612_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1742 diff_4663_3713# diff_2512_3700# diff_4663_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1743 diff_4714_3713# diff_2512_3700# diff_4714_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1744 diff_4765_3713# diff_2512_3700# diff_4765_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1745 diff_4816_3713# diff_2512_3700# diff_4816_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1746 diff_4867_3713# diff_2512_3700# diff_4867_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1747 diff_4918_3713# diff_2512_3700# diff_4918_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1748 diff_4969_3713# diff_2512_3700# diff_4969_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1749 diff_5020_3713# diff_2512_3700# diff_5020_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1750 diff_5071_3713# diff_2512_3700# diff_5071_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1751 diff_5122_3713# diff_2512_3700# diff_5122_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1752 diff_5173_3713# diff_2512_3700# diff_5173_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1753 diff_5224_3713# diff_2512_3700# diff_5224_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1754 diff_5275_3713# diff_2512_3700# diff_5275_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1755 diff_5326_3713# diff_2512_3700# diff_5326_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1756 diff_5377_3713# diff_2512_3700# diff_5377_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1757 diff_5428_3713# diff_2512_3700# diff_5428_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1758 diff_5479_3713# diff_2512_3700# diff_5479_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1759 diff_5530_3713# diff_2512_3700# diff_5530_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1760 diff_5581_3713# diff_2512_3700# diff_5581_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1761 diff_5632_3713# diff_2512_3700# diff_5632_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1762 diff_5683_3713# diff_2512_3700# diff_5683_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1763 diff_5734_3713# diff_2512_3700# diff_5734_3659# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1764 diff_2512_3757# Vdd Vdd GND efet w=13 l=28
+ ad=0 pd=0 as=0 ps=0 
M1765 diff_2521_3659# diff_2512_3646# diff_2521_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1766 diff_2572_3659# diff_2512_3646# diff_2572_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1767 diff_2623_3659# diff_2512_3646# diff_2623_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1768 diff_2674_3659# diff_2512_3646# diff_2674_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1769 diff_2725_3659# diff_2512_3646# diff_2725_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1770 diff_2776_3659# diff_2512_3646# diff_2776_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1771 diff_2827_3659# diff_2512_3646# diff_2827_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1772 diff_2878_3659# diff_2512_3646# diff_2878_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1773 diff_2929_3659# diff_2512_3646# diff_2929_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1774 diff_2980_3659# diff_2512_3646# diff_2980_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1775 diff_3031_3659# diff_2512_3646# diff_3031_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1776 diff_3082_3659# diff_2512_3646# diff_3082_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1777 diff_3133_3659# diff_2512_3646# diff_3133_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1778 diff_3184_3659# diff_2512_3646# diff_3184_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1779 diff_3235_3659# diff_2512_3646# diff_3235_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1780 diff_3286_3659# diff_2512_3646# diff_3286_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1781 diff_3337_3659# diff_2512_3646# diff_3337_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1782 diff_3388_3659# diff_2512_3646# diff_3388_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1783 diff_3439_3659# diff_2512_3646# diff_3439_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1784 diff_3490_3659# diff_2512_3646# diff_3490_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1785 diff_3541_3659# diff_2512_3646# diff_3541_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1786 diff_3592_3659# diff_2512_3646# diff_3592_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1787 diff_3643_3659# diff_2512_3646# diff_3643_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1788 diff_3694_3659# diff_2512_3646# diff_3694_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1789 diff_3745_3659# diff_2512_3646# diff_3745_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1790 diff_3796_3659# diff_2512_3646# diff_3796_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1791 diff_3847_3659# diff_2512_3646# diff_3847_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1792 diff_3898_3659# diff_2512_3646# diff_3898_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1793 diff_3949_3659# diff_2512_3646# diff_3949_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1794 diff_4000_3659# diff_2512_3646# diff_4000_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1795 diff_4051_3659# diff_2512_3646# diff_4051_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1796 diff_4102_3659# diff_2512_3646# diff_4102_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1797 diff_4153_3659# diff_2512_3646# diff_4153_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1798 diff_4204_3659# diff_2512_3646# diff_4204_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1799 diff_4255_3659# diff_2512_3646# diff_4255_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1800 diff_4306_3659# diff_2512_3646# diff_4306_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1801 diff_4357_3659# diff_2512_3646# diff_4357_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1802 diff_4408_3659# diff_2512_3646# diff_4408_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1803 diff_4459_3659# diff_2512_3646# diff_4459_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1804 diff_4510_3659# diff_2512_3646# diff_4510_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1805 diff_4561_3659# diff_2512_3646# diff_4561_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1806 diff_4612_3659# diff_2512_3646# diff_4612_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1807 diff_4663_3659# diff_2512_3646# diff_4663_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1808 diff_4714_3659# diff_2512_3646# diff_4714_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1809 diff_4765_3659# diff_2512_3646# diff_4765_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1810 diff_4816_3659# diff_2512_3646# diff_4816_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1811 diff_4867_3659# diff_2512_3646# diff_4867_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1812 diff_4918_3659# diff_2512_3646# diff_4918_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1813 diff_4969_3659# diff_2512_3646# diff_4969_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1814 diff_5020_3659# diff_2512_3646# diff_5020_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1815 diff_5071_3659# diff_2512_3646# diff_5071_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1816 diff_5122_3659# diff_2512_3646# diff_5122_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1817 diff_5173_3659# diff_2512_3646# diff_5173_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1818 diff_5224_3659# diff_2512_3646# diff_5224_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1819 diff_5275_3659# diff_2512_3646# diff_5275_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1820 diff_5326_3659# diff_2512_3646# diff_5326_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1821 diff_5377_3659# diff_2512_3646# diff_5377_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1822 diff_5428_3659# diff_2512_3646# diff_5428_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1823 diff_5479_3659# diff_2512_3646# diff_5479_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1824 diff_5530_3659# diff_2512_3646# diff_5530_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1825 diff_5581_3659# diff_2512_3646# diff_5581_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1826 diff_5632_3659# diff_2512_3646# diff_5632_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1827 diff_5683_3659# diff_2512_3646# diff_5683_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1828 diff_5734_3659# diff_2512_3646# diff_5734_3602# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1829 Vdd Vdd diff_2512_3589# GND efet w=13 l=31
+ ad=0 pd=0 as=5073 ps=640 
M1830 diff_2521_3602# diff_2512_3589# diff_2521_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1831 diff_2572_3602# diff_2512_3589# diff_2572_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1832 diff_2623_3602# diff_2512_3589# diff_2623_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1833 diff_2674_3602# diff_2512_3589# diff_2674_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1834 diff_2725_3602# diff_2512_3589# diff_2725_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1835 diff_2776_3602# diff_2512_3589# diff_2776_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1836 diff_2827_3602# diff_2512_3589# diff_2827_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1837 diff_2878_3602# diff_2512_3589# diff_2878_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1838 diff_2929_3602# diff_2512_3589# diff_2929_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1839 diff_2980_3602# diff_2512_3589# diff_2980_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1840 diff_3031_3602# diff_2512_3589# diff_3031_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1841 diff_3082_3602# diff_2512_3589# diff_3082_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1842 diff_3133_3602# diff_2512_3589# diff_3133_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1843 diff_3184_3602# diff_2512_3589# diff_3184_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1844 diff_3235_3602# diff_2512_3589# diff_3235_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1845 diff_3286_3602# diff_2512_3589# diff_3286_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1846 diff_3337_3602# diff_2512_3589# diff_3337_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1847 diff_3388_3602# diff_2512_3589# diff_3388_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1848 diff_3439_3602# diff_2512_3589# diff_3439_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1849 diff_3490_3602# diff_2512_3589# diff_3490_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1850 diff_3541_3602# diff_2512_3589# diff_3541_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1851 diff_3592_3602# diff_2512_3589# diff_3592_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1852 diff_3643_3602# diff_2512_3589# diff_3643_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1853 diff_3694_3602# diff_2512_3589# diff_3694_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1854 diff_3745_3602# diff_2512_3589# diff_3745_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1855 diff_3796_3602# diff_2512_3589# diff_3796_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1856 diff_3847_3602# diff_2512_3589# diff_3847_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1857 diff_3898_3602# diff_2512_3589# diff_3898_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1858 diff_3949_3602# diff_2512_3589# diff_3949_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1859 diff_4000_3602# diff_2512_3589# diff_4000_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1860 diff_4051_3602# diff_2512_3589# diff_4051_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1861 diff_4102_3602# diff_2512_3589# diff_4102_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1862 diff_4153_3602# diff_2512_3589# diff_4153_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1863 diff_4204_3602# diff_2512_3589# diff_4204_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1864 diff_4255_3602# diff_2512_3589# diff_4255_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1865 diff_4306_3602# diff_2512_3589# diff_4306_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1866 diff_4357_3602# diff_2512_3589# diff_4357_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1867 diff_4408_3602# diff_2512_3589# diff_4408_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1868 diff_4459_3602# diff_2512_3589# diff_4459_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1869 diff_4510_3602# diff_2512_3589# diff_4510_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1870 diff_4561_3602# diff_2512_3589# diff_4561_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1871 diff_4612_3602# diff_2512_3589# diff_4612_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1872 diff_4663_3602# diff_2512_3589# diff_4663_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1873 diff_4714_3602# diff_2512_3589# diff_4714_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1874 diff_4765_3602# diff_2512_3589# diff_4765_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1875 diff_4816_3602# diff_2512_3589# diff_4816_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1876 diff_4867_3602# diff_2512_3589# diff_4867_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1877 diff_4918_3602# diff_2512_3589# diff_4918_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1878 diff_4969_3602# diff_2512_3589# diff_4969_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1879 diff_5020_3602# diff_2512_3589# diff_5020_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1880 diff_5071_3602# diff_2512_3589# diff_5071_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1881 diff_5122_3602# diff_2512_3589# diff_5122_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1882 diff_5173_3602# diff_2512_3589# diff_5173_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1883 diff_5224_3602# diff_2512_3589# diff_5224_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1884 diff_5275_3602# diff_2512_3589# diff_5275_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1885 diff_5326_3602# diff_2512_3589# diff_5326_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1886 diff_5377_3602# diff_2512_3589# diff_5377_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1887 diff_5428_3602# diff_2512_3589# diff_5428_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1888 diff_5479_3602# diff_2512_3589# diff_5479_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1889 diff_5530_3602# diff_2512_3589# diff_5530_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1890 diff_5581_3602# diff_2512_3589# diff_5581_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1891 diff_5632_3602# diff_2512_3589# diff_5632_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1892 diff_5683_3602# diff_2512_3589# diff_5683_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1893 diff_5734_3602# diff_2512_3589# diff_5734_3548# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1894 diff_2011_4156# diff_475_2011# GND GND efet w=475 l=16
+ ad=0 pd=0 as=0 ps=0 
M1895 diff_2512_3589# diff_5962_1069# diff_5918_3734# GND efet w=184 l=13
+ ad=0 pd=0 as=0 ps=0 
M1896 diff_5918_3734# diff_6034_2491# diff_2512_3700# GND efet w=208 l=13
+ ad=0 pd=0 as=7100 ps=570 
M1897 diff_2512_3700# Vdd Vdd GND efet w=16 l=25
+ ad=0 pd=0 as=0 ps=0 
M1898 Vdd Vdd diff_2512_3646# GND efet w=16 l=28
+ ad=0 pd=0 as=5700 ps=610 
M1899 diff_2521_3548# diff_2512_3535# diff_2521_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1900 diff_2572_3548# diff_2512_3535# diff_2572_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1901 diff_2623_3548# diff_2512_3535# diff_2623_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1902 diff_2674_3548# diff_2512_3535# diff_2674_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1903 diff_2725_3548# diff_2512_3535# diff_2725_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1904 diff_2776_3548# diff_2512_3535# diff_2776_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1905 diff_2827_3548# diff_2512_3535# diff_2827_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1906 diff_2878_3548# diff_2512_3535# diff_2878_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1907 diff_2929_3548# diff_2512_3535# diff_2929_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1908 diff_2980_3548# diff_2512_3535# diff_2980_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1909 diff_3031_3548# diff_2512_3535# diff_3031_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1910 diff_3082_3548# diff_2512_3535# diff_3082_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1911 diff_3133_3548# diff_2512_3535# diff_3133_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1912 diff_3184_3548# diff_2512_3535# diff_3184_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1913 diff_3235_3548# diff_2512_3535# diff_3235_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1914 diff_3286_3548# diff_2512_3535# diff_3286_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1915 diff_3337_3548# diff_2512_3535# diff_3337_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1916 diff_3388_3548# diff_2512_3535# diff_3388_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1917 diff_3439_3548# diff_2512_3535# diff_3439_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1918 diff_3490_3548# diff_2512_3535# diff_3490_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1919 diff_3541_3548# diff_2512_3535# diff_3541_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1920 diff_3592_3548# diff_2512_3535# diff_3592_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1921 diff_3643_3548# diff_2512_3535# diff_3643_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1922 diff_3694_3548# diff_2512_3535# diff_3694_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1923 diff_3745_3548# diff_2512_3535# diff_3745_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1924 diff_3796_3548# diff_2512_3535# diff_3796_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1925 diff_3847_3548# diff_2512_3535# diff_3847_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1926 diff_3898_3548# diff_2512_3535# diff_3898_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1927 diff_3949_3548# diff_2512_3535# diff_3949_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1928 diff_4000_3548# diff_2512_3535# diff_4000_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1929 diff_4051_3548# diff_2512_3535# diff_4051_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1930 diff_4102_3548# diff_2512_3535# diff_4102_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1931 diff_4153_3548# diff_2512_3535# diff_4153_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1932 diff_4204_3548# diff_2512_3535# diff_4204_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1933 diff_4255_3548# diff_2512_3535# diff_4255_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1934 diff_4306_3548# diff_2512_3535# diff_4306_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1935 diff_4357_3548# diff_2512_3535# diff_4357_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1936 diff_4408_3548# diff_2512_3535# diff_4408_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1937 diff_4459_3548# diff_2512_3535# diff_4459_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1938 diff_4510_3548# diff_2512_3535# diff_4510_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1939 diff_4561_3548# diff_2512_3535# diff_4561_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1940 diff_4612_3548# diff_2512_3535# diff_4612_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1941 diff_4663_3548# diff_2512_3535# diff_4663_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1942 diff_4714_3548# diff_2512_3535# diff_4714_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1943 diff_4765_3548# diff_2512_3535# diff_4765_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1944 diff_4816_3548# diff_2512_3535# diff_4816_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1945 diff_4867_3548# diff_2512_3535# diff_4867_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1946 diff_4918_3548# diff_2512_3535# diff_4918_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1947 diff_4969_3548# diff_2512_3535# diff_4969_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1948 diff_5020_3548# diff_2512_3535# diff_5020_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1949 diff_5071_3548# diff_2512_3535# diff_5071_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1950 diff_5122_3548# diff_2512_3535# diff_5122_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1951 diff_5173_3548# diff_2512_3535# diff_5173_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1952 diff_5224_3548# diff_2512_3535# diff_5224_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1953 diff_5275_3548# diff_2512_3535# diff_5275_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1954 diff_5326_3548# diff_2512_3535# diff_5326_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1955 diff_5377_3548# diff_2512_3535# diff_5377_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1956 diff_5428_3548# diff_2512_3535# diff_5428_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1957 diff_5479_3548# diff_2512_3535# diff_5479_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1958 diff_5530_3548# diff_2512_3535# diff_5530_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1959 diff_5581_3548# diff_2512_3535# diff_5581_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1960 diff_5632_3548# diff_2512_3535# diff_5632_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1961 diff_5683_3548# diff_2512_3535# diff_5683_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1962 diff_5734_3548# diff_2512_3535# diff_5734_3491# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M1963 diff_5918_3518# diff_5905_1069# diff_2512_3535# GND efet w=214 l=13
+ ad=24475 pd=1820 as=5930 ps=576 
M1964 diff_2512_3646# diff_6079_2449# diff_5918_3734# GND efet w=196 l=13
+ ad=0 pd=0 as=0 ps=0 
M1965 diff_2521_3491# diff_2512_3478# diff_2521_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1966 diff_2572_3491# diff_2512_3478# diff_2572_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1967 diff_2623_3491# diff_2512_3478# diff_2623_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1968 diff_2674_3491# diff_2512_3478# diff_2674_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1969 diff_2725_3491# diff_2512_3478# diff_2725_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1970 diff_2776_3491# diff_2512_3478# diff_2776_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1971 diff_2827_3491# diff_2512_3478# diff_2827_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1972 diff_2878_3491# diff_2512_3478# diff_2878_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1973 diff_2929_3491# diff_2512_3478# diff_2929_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1974 diff_2980_3491# diff_2512_3478# diff_2980_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1975 diff_3031_3491# diff_2512_3478# diff_3031_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1976 diff_3082_3491# diff_2512_3478# diff_3082_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1977 diff_3133_3491# diff_2512_3478# diff_3133_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1978 diff_3184_3491# diff_2512_3478# diff_3184_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1979 diff_3235_3491# diff_2512_3478# diff_3235_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1980 diff_3286_3491# diff_2512_3478# diff_3286_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1981 diff_3337_3491# diff_2512_3478# diff_3337_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1982 diff_3388_3491# diff_2512_3478# diff_3388_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1983 diff_3439_3491# diff_2512_3478# diff_3439_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1984 diff_3490_3491# diff_2512_3478# diff_3490_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1985 diff_3541_3491# diff_2512_3478# diff_3541_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1986 diff_3592_3491# diff_2512_3478# diff_3592_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1987 diff_3643_3491# diff_2512_3478# diff_3643_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1988 diff_3694_3491# diff_2512_3478# diff_3694_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1989 diff_3745_3491# diff_2512_3478# diff_3745_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1990 diff_3796_3491# diff_2512_3478# diff_3796_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1991 diff_3847_3491# diff_2512_3478# diff_3847_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1992 diff_3898_3491# diff_2512_3478# diff_3898_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1993 diff_3949_3491# diff_2512_3478# diff_3949_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1994 diff_4000_3491# diff_2512_3478# diff_4000_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1995 diff_4051_3491# diff_2512_3478# diff_4051_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1996 diff_4102_3491# diff_2512_3478# diff_4102_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1997 diff_4153_3491# diff_2512_3478# diff_4153_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1998 diff_4204_3491# diff_2512_3478# diff_4204_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M1999 diff_4255_3491# diff_2512_3478# diff_4255_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2000 diff_4306_3491# diff_2512_3478# diff_4306_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2001 diff_4357_3491# diff_2512_3478# diff_4357_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2002 diff_4408_3491# diff_2512_3478# diff_4408_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2003 diff_4459_3491# diff_2512_3478# diff_4459_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2004 diff_4510_3491# diff_2512_3478# diff_4510_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2005 diff_4561_3491# diff_2512_3478# diff_4561_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2006 diff_4612_3491# diff_2512_3478# diff_4612_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2007 diff_4663_3491# diff_2512_3478# diff_4663_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2008 diff_4714_3491# diff_2512_3478# diff_4714_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2009 diff_4765_3491# diff_2512_3478# diff_4765_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2010 diff_4816_3491# diff_2512_3478# diff_4816_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2011 diff_4867_3491# diff_2512_3478# diff_4867_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2012 diff_4918_3491# diff_2512_3478# diff_4918_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2013 diff_4969_3491# diff_2512_3478# diff_4969_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2014 diff_5020_3491# diff_2512_3478# diff_5020_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2015 diff_5071_3491# diff_2512_3478# diff_5071_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2016 diff_5122_3491# diff_2512_3478# diff_5122_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2017 diff_5173_3491# diff_2512_3478# diff_5173_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2018 diff_5224_3491# diff_2512_3478# diff_5224_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2019 diff_5275_3491# diff_2512_3478# diff_5275_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2020 diff_5326_3491# diff_2512_3478# diff_5326_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2021 diff_5377_3491# diff_2512_3478# diff_5377_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2022 diff_5428_3491# diff_2512_3478# diff_5428_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2023 diff_5479_3491# diff_2512_3478# diff_5479_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2024 diff_5530_3491# diff_2512_3478# diff_5530_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2025 diff_5581_3491# diff_2512_3478# diff_5581_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2026 diff_5632_3491# diff_2512_3478# diff_5632_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2027 diff_5683_3491# diff_2512_3478# diff_5683_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2028 diff_5734_3491# diff_2512_3478# diff_5734_3437# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2029 diff_2512_3535# Vdd Vdd GND efet w=13 l=28
+ ad=0 pd=0 as=0 ps=0 
M2030 diff_2521_3437# diff_2512_3424# diff_2521_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2031 diff_2572_3437# diff_2512_3424# diff_2572_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2032 diff_2623_3437# diff_2512_3424# diff_2623_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2033 diff_2674_3437# diff_2512_3424# diff_2674_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2034 diff_2725_3437# diff_2512_3424# diff_2725_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2035 diff_2776_3437# diff_2512_3424# diff_2776_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2036 diff_2827_3437# diff_2512_3424# diff_2827_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2037 diff_2878_3437# diff_2512_3424# diff_2878_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2038 diff_2929_3437# diff_2512_3424# diff_2929_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2039 diff_2980_3437# diff_2512_3424# diff_2980_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2040 diff_3031_3437# diff_2512_3424# diff_3031_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2041 diff_3082_3437# diff_2512_3424# diff_3082_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2042 diff_3133_3437# diff_2512_3424# diff_3133_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2043 diff_3184_3437# diff_2512_3424# diff_3184_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2044 diff_3235_3437# diff_2512_3424# diff_3235_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2045 diff_3286_3437# diff_2512_3424# diff_3286_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2046 diff_3337_3437# diff_2512_3424# diff_3337_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2047 diff_3388_3437# diff_2512_3424# diff_3388_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2048 diff_3439_3437# diff_2512_3424# diff_3439_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2049 diff_3490_3437# diff_2512_3424# diff_3490_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2050 diff_3541_3437# diff_2512_3424# diff_3541_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2051 diff_3592_3437# diff_2512_3424# diff_3592_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2052 diff_3643_3437# diff_2512_3424# diff_3643_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2053 diff_3694_3437# diff_2512_3424# diff_3694_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2054 diff_3745_3437# diff_2512_3424# diff_3745_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2055 diff_3796_3437# diff_2512_3424# diff_3796_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2056 diff_3847_3437# diff_2512_3424# diff_3847_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2057 diff_3898_3437# diff_2512_3424# diff_3898_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2058 diff_3949_3437# diff_2512_3424# diff_3949_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2059 diff_4000_3437# diff_2512_3424# diff_4000_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2060 diff_4051_3437# diff_2512_3424# diff_4051_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2061 diff_4102_3437# diff_2512_3424# diff_4102_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2062 diff_4153_3437# diff_2512_3424# diff_4153_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2063 diff_4204_3437# diff_2512_3424# diff_4204_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2064 diff_4255_3437# diff_2512_3424# diff_4255_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2065 diff_4306_3437# diff_2512_3424# diff_4306_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2066 diff_4357_3437# diff_2512_3424# diff_4357_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2067 diff_4408_3437# diff_2512_3424# diff_4408_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2068 diff_4459_3437# diff_2512_3424# diff_4459_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2069 diff_4510_3437# diff_2512_3424# diff_4510_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2070 diff_4561_3437# diff_2512_3424# diff_4561_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2071 diff_4612_3437# diff_2512_3424# diff_4612_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2072 diff_4663_3437# diff_2512_3424# diff_4663_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2073 diff_4714_3437# diff_2512_3424# diff_4714_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2074 diff_4765_3437# diff_2512_3424# diff_4765_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2075 diff_4816_3437# diff_2512_3424# diff_4816_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2076 diff_4867_3437# diff_2512_3424# diff_4867_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2077 diff_4918_3437# diff_2512_3424# diff_4918_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2078 diff_4969_3437# diff_2512_3424# diff_4969_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2079 diff_5020_3437# diff_2512_3424# diff_5020_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2080 diff_5071_3437# diff_2512_3424# diff_5071_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2081 diff_5122_3437# diff_2512_3424# diff_5122_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2082 diff_5173_3437# diff_2512_3424# diff_5173_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2083 diff_5224_3437# diff_2512_3424# diff_5224_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2084 diff_5275_3437# diff_2512_3424# diff_5275_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2085 diff_5326_3437# diff_2512_3424# diff_5326_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2086 diff_5377_3437# diff_2512_3424# diff_5377_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2087 diff_5428_3437# diff_2512_3424# diff_5428_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2088 diff_5479_3437# diff_2512_3424# diff_5479_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2089 diff_5530_3437# diff_2512_3424# diff_5530_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2090 diff_5581_3437# diff_2512_3424# diff_5581_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2091 diff_5632_3437# diff_2512_3424# diff_5632_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2092 diff_5683_3437# diff_2512_3424# diff_5683_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2093 diff_5734_3437# diff_2512_3424# diff_5734_3380# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2094 d3 clk2 diff_835_3365# GND efet w=28 l=16
+ ad=0 pd=0 as=644 ps=102 
M2095 d2 clk2 diff_1222_3365# GND efet w=28 l=16
+ ad=0 pd=0 as=644 ps=102 
M2096 d1 clk2 diff_1612_3365# GND efet w=28 l=16
+ ad=0 pd=0 as=644 ps=102 
M2097 d0 clk2 diff_1999_3365# GND efet w=28 l=16
+ ad=0 pd=0 as=644 ps=102 
M2098 Vdd Vdd diff_2512_3367# GND efet w=13 l=31
+ ad=0 pd=0 as=5073 ps=640 
M2099 diff_835_3365# diff_388_2056# diff_835_3196# GND efet w=28 l=16
+ ad=0 pd=0 as=10160 ps=880 
M2100 diff_1222_3365# diff_388_2056# diff_1222_3193# GND efet w=28 l=16
+ ad=0 pd=0 as=9935 ps=874 
M2101 diff_1612_3365# diff_388_2056# diff_1612_3193# GND efet w=28 l=16
+ ad=0 pd=0 as=10271 ps=874 
M2102 diff_1999_3365# diff_388_2056# diff_1999_3193# GND efet w=28 l=16
+ ad=0 pd=0 as=10232 ps=886 
M2103 diff_2521_3380# diff_2512_3367# diff_2521_3301# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2104 diff_2572_3380# diff_2512_3367# diff_2563_3160# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2105 diff_2623_3380# diff_2512_3367# diff_2623_3307# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2106 diff_2674_3380# diff_2512_3367# diff_2674_3205# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2107 diff_2725_3380# diff_2512_3367# diff_2725_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2108 diff_2776_3380# diff_2512_3367# diff_2776_3157# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2109 diff_2827_3380# diff_2512_3367# diff_2827_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2110 diff_2878_3380# diff_2512_3367# diff_2878_3205# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2111 diff_2929_3380# diff_2512_3367# diff_2929_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2112 diff_2980_3380# diff_2512_3367# diff_2980_3157# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2113 diff_3031_3380# diff_2512_3367# diff_3031_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2114 diff_3082_3380# diff_2512_3367# diff_3082_3205# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2115 diff_3133_3380# diff_2512_3367# diff_3133_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2116 diff_3184_3380# diff_2512_3367# diff_3184_3157# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2117 diff_3235_3380# diff_2512_3367# diff_3235_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2118 diff_3286_3380# diff_2512_3367# diff_3286_3205# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2119 diff_3337_3380# diff_2512_3367# diff_3337_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2120 diff_3388_3380# diff_2512_3367# diff_3388_3157# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2121 diff_3439_3380# diff_2512_3367# diff_3439_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2122 diff_3490_3380# diff_2512_3367# diff_3490_3205# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2123 diff_3541_3380# diff_2512_3367# diff_3541_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2124 diff_3592_3380# diff_2512_3367# diff_3592_3157# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2125 diff_3643_3380# diff_2512_3367# diff_3643_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2126 diff_3694_3380# diff_2512_3367# diff_3694_3205# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2127 diff_3745_3380# diff_2512_3367# diff_3745_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2128 diff_3796_3380# diff_2512_3367# diff_3796_3157# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2129 diff_3847_3380# diff_2512_3367# diff_3847_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2130 diff_3898_3380# diff_2512_3367# diff_3898_3205# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2131 diff_3949_3380# diff_2512_3367# diff_3949_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2132 diff_4000_3380# diff_2512_3367# diff_4000_3157# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2133 diff_4051_3380# diff_2512_3367# diff_4051_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2134 diff_4102_3380# diff_2512_3367# diff_4102_3205# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2135 diff_4153_3380# diff_2512_3367# diff_4153_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2136 diff_4204_3380# diff_2512_3367# diff_4204_3157# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2137 diff_4255_3380# diff_2512_3367# diff_4255_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2138 diff_4306_3380# diff_2512_3367# diff_4306_3205# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2139 diff_4357_3380# diff_2512_3367# diff_4357_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2140 diff_4408_3380# diff_2512_3367# diff_4408_3157# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2141 diff_4459_3380# diff_2512_3367# diff_4459_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2142 diff_4510_3380# diff_2512_3367# diff_4510_3205# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2143 diff_4561_3380# diff_2512_3367# diff_4561_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2144 diff_4612_3380# diff_2512_3367# diff_4612_3157# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2145 diff_4663_3380# diff_2512_3367# diff_4663_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2146 diff_4714_3380# diff_2512_3367# diff_4714_3205# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2147 diff_4765_3380# diff_2512_3367# diff_4765_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2148 diff_4816_3380# diff_2512_3367# diff_4816_3157# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2149 diff_4867_3380# diff_2512_3367# diff_4867_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2150 diff_4918_3380# diff_2512_3367# diff_4918_3205# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2151 diff_4969_3380# diff_2512_3367# diff_4969_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2152 diff_5020_3380# diff_2512_3367# diff_5020_3157# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2153 diff_5071_3380# diff_2512_3367# diff_5071_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2154 diff_5122_3380# diff_2512_3367# diff_5122_3205# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2155 diff_5173_3380# diff_2512_3367# diff_5173_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2156 diff_5224_3380# diff_2512_3367# diff_5224_3157# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2157 diff_5275_3380# diff_2512_3367# diff_5275_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2158 diff_5326_3380# diff_2512_3367# diff_5326_3205# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2159 diff_5377_3380# diff_2512_3367# diff_5377_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2160 diff_5428_3380# diff_2512_3367# diff_5428_3157# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2161 diff_5479_3380# diff_2512_3367# diff_5479_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2162 diff_5530_3380# diff_2512_3367# diff_5530_3205# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2163 diff_5581_3380# diff_2512_3367# diff_5581_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2164 diff_5632_3380# diff_2512_3367# diff_5632_3157# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2165 diff_5683_3380# diff_2512_3367# diff_5683_3304# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2166 diff_5734_3380# diff_2512_3367# diff_5734_3205# GND efet w=25 l=16
+ ad=0 pd=0 as=732 ps=110 
M2167 diff_701_3292# diff_388_2056# GND GND efet w=43 l=16
+ ad=1553 pd=180 as=0 ps=0 
M2168 diff_835_3196# diff_835_3196# diff_835_3196# GND efet w=7 l=7
+ ad=0 pd=0 as=0 ps=0 
M2169 Vdd Vdd diff_701_3292# GND efet w=8 l=101
+ ad=0 pd=0 as=0 ps=0 
M2170 GND GND sync GND efet w=287 l=17
+ ad=0 pd=0 as=0 ps=0 
M2171 diff_841_2926# diff_835_3196# GND GND efet w=190 l=16
+ ad=4560 pd=544 as=0 ps=0 
M2172 diff_1222_3193# diff_1222_3193# diff_1222_3193# GND efet w=7 l=7
+ ad=0 pd=0 as=0 ps=0 
M2173 diff_835_3196# diff_835_3196# diff_835_3196# GND efet w=4 l=4
+ ad=0 pd=0 as=0 ps=0 
M2174 GND diff_841_2926# diff_889_3250# GND efet w=124 l=13
+ ad=0 pd=0 as=8069 ps=860 
M2175 diff_889_3250# diff_701_3292# diff_835_3196# GND efet w=28 l=16
+ ad=0 pd=0 as=0 ps=0 
M2176 diff_1231_2926# diff_1222_3193# GND GND efet w=190 l=16
+ ad=4515 pd=544 as=0 ps=0 
M2177 diff_1612_3193# diff_1612_3193# diff_1612_3193# GND efet w=4 l=4
+ ad=0 pd=0 as=0 ps=0 
M2178 diff_1222_3193# diff_1222_3193# diff_1222_3193# GND efet w=4 l=4
+ ad=0 pd=0 as=0 ps=0 
M2179 GND diff_1231_2926# diff_1273_3250# GND efet w=124 l=13
+ ad=0 pd=0 as=8084 ps=854 
M2180 diff_1273_3250# diff_701_3292# diff_1222_3193# GND efet w=28 l=16
+ ad=0 pd=0 as=0 ps=0 
M2181 diff_1618_2926# diff_1612_3193# GND GND efet w=187 l=16
+ ad=4830 pd=538 as=0 ps=0 
M2182 diff_2512_3367# diff_5962_1069# diff_5918_3518# GND efet w=184 l=13
+ ad=0 pd=0 as=0 ps=0 
M2183 diff_5918_3518# diff_6034_2491# diff_2512_3478# GND efet w=211 l=13
+ ad=0 pd=0 as=7067 ps=570 
M2184 diff_2512_3478# Vdd Vdd GND efet w=16 l=25
+ ad=0 pd=0 as=0 ps=0 
M2185 Vdd Vdd diff_2512_3424# GND efet w=16 l=31
+ ad=0 pd=0 as=5700 ps=610 
M2186 diff_1999_3193# diff_1999_3193# diff_1999_3193# GND efet w=7 l=7
+ ad=0 pd=0 as=0 ps=0 
M2187 diff_1612_3193# diff_1612_3193# diff_1612_3193# GND efet w=1 l=1
+ ad=0 pd=0 as=0 ps=0 
M2188 GND diff_1618_2926# diff_1666_3250# GND efet w=124 l=16
+ ad=0 pd=0 as=7868 ps=848 
M2189 diff_1666_3250# diff_701_3292# diff_1612_3193# GND efet w=28 l=16
+ ad=0 pd=0 as=0 ps=0 
M2190 diff_2005_2926# diff_1999_3193# GND GND efet w=190 l=16
+ ad=4521 pd=538 as=0 ps=0 
M2191 diff_1999_3193# diff_1999_3193# diff_1999_3193# GND efet w=4 l=4
+ ad=0 pd=0 as=0 ps=0 
M2192 GND diff_2005_2926# diff_2053_3250# GND efet w=124 l=13
+ ad=0 pd=0 as=8030 ps=854 
M2193 diff_2053_3250# diff_701_3292# diff_1999_3193# GND efet w=28 l=16
+ ad=0 pd=0 as=0 ps=0 
M2194 diff_835_3196# cl GND GND efet w=88 l=16
+ ad=0 pd=0 as=0 ps=0 
M2195 GND cl diff_835_3196# GND efet w=88 l=19
+ ad=0 pd=0 as=0 ps=0 
M2196 diff_835_3196# diff_652_1966# GND GND efet w=116 l=17
+ ad=0 pd=0 as=0 ps=0 
M2197 diff_841_2926# Vdd Vdd GND efet w=13 l=37
+ ad=0 pd=0 as=0 ps=0 
M2198 diff_889_3250# Vdd Vdd GND efet w=13 l=34
+ ad=0 pd=0 as=0 ps=0 
M2199 Vdd Vdd Vdd GND efet w=4 l=4
+ ad=0 pd=0 as=0 ps=0 
M2200 Vdd Vdd Vdd GND efet w=3 l=4
+ ad=0 pd=0 as=0 ps=0 
M2201 diff_1222_3193# cl GND GND efet w=88 l=16
+ ad=0 pd=0 as=0 ps=0 
M2202 GND cl diff_1222_3193# GND efet w=88 l=19
+ ad=0 pd=0 as=0 ps=0 
M2203 GND diff_2521_3301# diff_2494_3091# GND efet w=70 l=13
+ ad=0 pd=0 as=4808 ps=486 
M2204 GND diff_2623_3307# diff_2593_3005# GND efet w=97 l=13
+ ad=0 pd=0 as=4578 ps=472 
M2205 diff_2687_3211# diff_2674_3205# GND GND efet w=97 l=13
+ ad=3891 pd=460 as=0 ps=0 
M2206 diff_2582_3167# diff_2563_3160# GND GND efet w=113 l=18
+ ad=2420 pd=264 as=0 ps=0 
M2207 GND diff_2725_3304# diff_2686_2951# GND efet w=87 l=16
+ ad=0 pd=0 as=4056 ps=434 
M2208 GND diff_2827_3304# diff_2791_3002# GND efet w=97 l=13
+ ad=0 pd=0 as=4611 ps=484 
M2209 diff_2891_3211# diff_2878_3205# GND GND efet w=97 l=13
+ ad=4023 pd=460 as=0 ps=0 
M2210 diff_2789_3164# diff_2776_3157# GND GND efet w=85 l=13
+ ad=2135 pd=234 as=0 ps=0 
M2211 GND diff_2929_3304# diff_2890_2951# GND efet w=87 l=16
+ ad=0 pd=0 as=4092 ps=434 
M2212 GND diff_3031_3304# diff_2995_3005# GND efet w=97 l=13
+ ad=0 pd=0 as=4713 ps=484 
M2213 diff_3095_3211# diff_3082_3205# GND GND efet w=97 l=13
+ ad=3987 pd=460 as=0 ps=0 
M2214 diff_2993_3164# diff_2980_3157# GND GND efet w=85 l=13
+ ad=2135 pd=234 as=0 ps=0 
M2215 GND diff_3133_3304# diff_3091_2951# GND efet w=87 l=16
+ ad=0 pd=0 as=4284 ps=440 
M2216 GND diff_3235_3304# diff_3196_3005# GND efet w=97 l=13
+ ad=0 pd=0 as=4830 ps=484 
M2217 diff_3299_3211# diff_3286_3205# GND GND efet w=97 l=13
+ ad=4191 pd=466 as=0 ps=0 
M2218 diff_3197_3164# diff_3184_3157# GND GND efet w=85 l=13
+ ad=2135 pd=234 as=0 ps=0 
M2219 GND diff_3337_3304# diff_3295_2951# GND efet w=87 l=16
+ ad=0 pd=0 as=4320 ps=440 
M2220 GND diff_3439_3304# diff_3400_3002# GND efet w=97 l=13
+ ad=0 pd=0 as=4950 ps=496 
M2221 diff_3503_3211# diff_3490_3205# GND GND efet w=97 l=13
+ ad=3624 pd=454 as=0 ps=0 
M2222 diff_3401_3164# diff_3388_3157# GND GND efet w=85 l=13
+ ad=2135 pd=234 as=0 ps=0 
M2223 GND diff_3541_3304# diff_3502_2951# GND efet w=87 l=16
+ ad=0 pd=0 as=3828 ps=428 
M2224 GND diff_3643_3304# diff_3607_3005# GND efet w=97 l=13
+ ad=0 pd=0 as=4374 ps=472 
M2225 diff_3707_3211# diff_3694_3205# GND GND efet w=97 l=13
+ ad=3783 pd=454 as=0 ps=0 
M2226 diff_3605_3164# diff_3592_3157# GND GND efet w=85 l=13
+ ad=2135 pd=234 as=0 ps=0 
M2227 GND diff_3745_3304# diff_3706_2951# GND efet w=87 l=16
+ ad=0 pd=0 as=3864 ps=428 
M2228 GND diff_3847_3304# diff_3811_3005# GND efet w=97 l=13
+ ad=0 pd=0 as=4485 ps=478 
M2229 diff_3911_3211# diff_3898_3205# GND GND efet w=97 l=13
+ ad=3624 pd=454 as=0 ps=0 
M2230 diff_3809_3164# diff_3796_3157# GND GND efet w=85 l=13
+ ad=2135 pd=234 as=0 ps=0 
M2231 GND diff_3949_3304# diff_3910_2951# GND efet w=87 l=16
+ ad=0 pd=0 as=3828 ps=428 
M2232 GND diff_4051_3304# diff_4015_3005# GND efet w=97 l=13
+ ad=0 pd=0 as=4374 ps=472 
M2233 diff_4115_3211# diff_4102_3205# GND GND efet w=97 l=13
+ ad=3804 pd=454 as=0 ps=0 
M2234 diff_4013_3164# diff_4000_3157# GND GND efet w=85 l=13
+ ad=2135 pd=234 as=0 ps=0 
M2235 GND diff_4153_3304# diff_4114_2951# GND efet w=87 l=16
+ ad=0 pd=0 as=3864 ps=428 
M2236 GND diff_4255_3304# diff_4219_3005# GND efet w=97 l=13
+ ad=0 pd=0 as=4485 ps=478 
M2237 diff_4319_3211# diff_4306_3205# GND GND efet w=97 l=13
+ ad=3858 pd=460 as=0 ps=0 
M2238 diff_4217_3164# diff_4204_3157# GND GND efet w=85 l=13
+ ad=2135 pd=234 as=0 ps=0 
M2239 GND diff_4357_3304# diff_4321_2951# GND efet w=87 l=16
+ ad=0 pd=0 as=4056 ps=434 
M2240 GND diff_4459_3304# diff_4426_3005# GND efet w=97 l=13
+ ad=0 pd=0 as=4602 ps=478 
M2241 diff_4523_3211# diff_4510_3205# GND GND efet w=97 l=13
+ ad=4035 pd=460 as=0 ps=0 
M2242 diff_4421_3164# diff_4408_3157# GND GND efet w=85 l=13
+ ad=2135 pd=234 as=0 ps=0 
M2243 GND diff_4561_3304# diff_4525_2951# GND efet w=87 l=16
+ ad=0 pd=0 as=4092 ps=434 
M2244 GND diff_4663_3304# diff_4630_3005# GND efet w=97 l=13
+ ad=0 pd=0 as=4713 ps=484 
M2245 diff_4727_3211# diff_4714_3205# GND GND efet w=97 l=13
+ ad=3855 pd=460 as=0 ps=0 
M2246 diff_4625_3164# diff_4612_3157# GND GND efet w=85 l=13
+ ad=2135 pd=234 as=0 ps=0 
M2247 GND diff_4765_3304# diff_4726_2951# GND efet w=87 l=16
+ ad=0 pd=0 as=4056 ps=434 
M2248 GND diff_4867_3304# diff_4831_3005# GND efet w=97 l=13
+ ad=0 pd=0 as=4602 ps=478 
M2249 diff_4931_3211# diff_4918_3205# GND GND efet w=97 l=13
+ ad=4023 pd=460 as=0 ps=0 
M2250 diff_4829_3164# diff_4816_3157# GND GND efet w=85 l=13
+ ad=2135 pd=234 as=0 ps=0 
M2251 GND diff_4969_3304# diff_4930_2951# GND efet w=87 l=16
+ ad=0 pd=0 as=4092 ps=434 
M2252 GND diff_5071_3304# diff_5035_3005# GND efet w=97 l=13
+ ad=0 pd=0 as=4713 ps=484 
M2253 diff_5135_3211# diff_5122_3205# GND GND efet w=97 l=13
+ ad=3855 pd=460 as=0 ps=0 
M2254 diff_5033_3164# diff_5020_3157# GND GND efet w=85 l=13
+ ad=2135 pd=234 as=0 ps=0 
M2255 GND diff_5173_3304# diff_5134_2951# GND efet w=87 l=16
+ ad=0 pd=0 as=4056 ps=434 
M2256 GND diff_5275_3304# diff_5239_3005# GND efet w=97 l=13
+ ad=0 pd=0 as=4602 ps=478 
M2257 diff_5339_3211# diff_5326_3205# GND GND efet w=97 l=13
+ ad=4023 pd=460 as=0 ps=0 
M2258 diff_5237_3164# diff_5224_3157# GND GND efet w=85 l=13
+ ad=2135 pd=234 as=0 ps=0 
M2259 GND diff_5377_3304# diff_5338_2951# GND efet w=87 l=16
+ ad=0 pd=0 as=4092 ps=434 
M2260 GND diff_5479_3304# diff_5443_3005# GND efet w=97 l=13
+ ad=0 pd=0 as=4713 ps=484 
M2261 diff_5543_3211# diff_5530_3205# GND GND efet w=97 l=13
+ ad=3747 pd=448 as=0 ps=0 
M2262 diff_5441_3164# diff_5428_3157# GND GND efet w=85 l=13
+ ad=2135 pd=234 as=0 ps=0 
M2263 GND diff_5581_3304# diff_5545_2951# GND efet w=87 l=16
+ ad=0 pd=0 as=4002 ps=428 
M2264 GND diff_5683_3304# diff_5650_3005# GND efet w=97 l=13
+ ad=0 pd=0 as=4467 ps=472 
M2265 diff_5747_3211# diff_5734_3205# GND GND efet w=97 l=13
+ ad=4860 pd=612 as=0 ps=0 
M2266 diff_5645_3164# diff_5632_3157# GND GND efet w=85 l=13
+ ad=2135 pd=234 as=0 ps=0 
M2267 diff_1222_3193# diff_652_1966# GND GND efet w=113 l=17
+ ad=0 pd=0 as=0 ps=0 
M2268 diff_1231_2926# Vdd Vdd GND efet w=13 l=37
+ ad=0 pd=0 as=0 ps=0 
M2269 diff_1273_3250# Vdd Vdd GND efet w=13 l=34
+ ad=0 pd=0 as=0 ps=0 
M2270 Vdd Vdd Vdd GND efet w=4 l=4
+ ad=0 pd=0 as=0 ps=0 
M2271 Vdd Vdd Vdd GND efet w=1 l=3
+ ad=0 pd=0 as=0 ps=0 
M2272 diff_1612_3193# cl GND GND efet w=88 l=16
+ ad=0 pd=0 as=0 ps=0 
M2273 GND cl diff_1612_3193# GND efet w=88 l=19
+ ad=0 pd=0 as=0 ps=0 
M2274 diff_1612_3193# diff_652_1966# GND GND efet w=119 l=17
+ ad=0 pd=0 as=0 ps=0 
M2275 diff_1618_2926# Vdd Vdd GND efet w=13 l=37
+ ad=0 pd=0 as=0 ps=0 
M2276 diff_1666_3250# Vdd Vdd GND efet w=13 l=34
+ ad=0 pd=0 as=0 ps=0 
M2277 Vdd Vdd Vdd GND efet w=1 l=1
+ ad=0 pd=0 as=0 ps=0 
M2278 Vdd Vdd Vdd GND efet w=1 l=1
+ ad=0 pd=0 as=0 ps=0 
M2279 diff_1999_3193# cl GND GND efet w=88 l=16
+ ad=0 pd=0 as=0 ps=0 
M2280 GND cl diff_1999_3193# GND efet w=88 l=19
+ ad=0 pd=0 as=0 ps=0 
M2281 diff_1999_3193# diff_652_1966# GND GND efet w=119 l=17
+ ad=0 pd=0 as=0 ps=0 
M2282 diff_2500_3043# diff_2623_2116# diff_2582_3167# GND efet w=76 l=16
+ ad=12363 pd=1180 as=0 ps=0 
M2283 diff_2695_3019# diff_2623_2116# diff_2789_3164# GND efet w=73 l=13
+ ad=10382 pd=1008 as=0 ps=0 
M2284 diff_2899_3019# diff_2623_2116# diff_2993_3164# GND efet w=73 l=13
+ ad=10668 pd=1126 as=0 ps=0 
M2285 diff_3100_3022# diff_2623_2116# diff_3197_3164# GND efet w=73 l=13
+ ad=9953 pd=996 as=0 ps=0 
M2286 diff_3304_3022# diff_2623_2116# diff_3401_3164# GND efet w=73 l=13
+ ad=10920 pd=1150 as=0 ps=0 
M2287 diff_3511_3016# diff_2623_2116# diff_3605_3164# GND efet w=73 l=13
+ ad=10703 pd=1020 as=0 ps=0 
M2288 diff_3715_3016# diff_2623_2116# diff_3809_3164# GND efet w=73 l=13
+ ad=11280 pd=1156 as=0 ps=0 
M2289 diff_3919_3016# diff_2623_2116# diff_4013_3164# GND efet w=73 l=13
+ ad=10703 pd=1020 as=0 ps=0 
M2290 diff_4123_3016# diff_2623_2116# diff_4217_3164# GND efet w=73 l=13
+ ad=11052 pd=1138 as=0 ps=0 
M2291 diff_4330_3019# diff_2623_2116# diff_4421_3164# GND efet w=73 l=13
+ ad=10394 pd=1008 as=0 ps=0 
M2292 diff_4534_3019# diff_2623_2116# diff_4625_3164# GND efet w=73 l=13
+ ad=10926 pd=1132 as=0 ps=0 
M2293 diff_4735_3019# diff_2623_2116# diff_4829_3164# GND efet w=73 l=13
+ ad=10364 pd=1008 as=0 ps=0 
M2294 diff_4939_3019# diff_2623_2116# diff_5033_3164# GND efet w=73 l=13
+ ad=10926 pd=1138 as=0 ps=0 
M2295 diff_5143_3019# diff_2623_2116# diff_5237_3164# GND efet w=73 l=13
+ ad=10364 pd=1008 as=0 ps=0 
M2296 diff_5347_3019# diff_2623_2116# diff_5441_3164# GND efet w=73 l=13
+ ad=11058 pd=1144 as=0 ps=0 
M2297 diff_5554_3016# diff_2623_2116# diff_5645_3164# GND efet w=73 l=13
+ ad=10892 pd=1054 as=0 ps=0 
M2298 diff_2512_3424# diff_6079_2449# diff_5918_3518# GND efet w=196 l=13
+ ad=0 pd=0 as=0 ps=0 
M2299 diff_6094_4246# diff_6130_2449# diff_5918_3518# GND efet w=385 l=16
+ ad=0 pd=0 as=0 ps=0 
M2300 diff_5918_3734# diff_6175_2281# diff_6094_4246# GND efet w=385 l=16
+ ad=0 pd=0 as=0 ps=0 
M2301 diff_2500_3043# diff_2488_3064# diff_2494_3091# GND efet w=100 l=13
+ ad=0 pd=0 as=0 ps=0 
M2302 diff_2005_2926# Vdd Vdd GND efet w=13 l=37
+ ad=0 pd=0 as=0 ps=0 
M2303 diff_2053_3250# Vdd Vdd GND efet w=13 l=34
+ ad=0 pd=0 as=0 ps=0 
M2304 diff_3299_3211# diff_2488_3064# diff_3304_3022# GND efet w=83 l=13
+ ad=0 pd=0 as=0 ps=0 
M2305 diff_3095_3211# diff_2488_3064# diff_3100_3022# GND efet w=76 l=14
+ ad=0 pd=0 as=0 ps=0 
M2306 diff_3503_3211# diff_2488_3064# diff_3511_3016# GND efet w=76 l=14
+ ad=0 pd=0 as=0 ps=0 
M2307 diff_3707_3211# diff_2488_3064# diff_3715_3016# GND efet w=79 l=13
+ ad=0 pd=0 as=0 ps=0 
M2308 diff_3911_3211# diff_2488_3064# diff_3919_3016# GND efet w=76 l=14
+ ad=0 pd=0 as=0 ps=0 
M2309 diff_2687_3211# diff_2488_3064# diff_2695_3019# GND efet w=74 l=14
+ ad=0 pd=0 as=0 ps=0 
M2310 Vdd Vdd Vdd GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M2311 Vdd Vdd Vdd GND efet w=1 l=1
+ ad=0 pd=0 as=0 ps=0 
M2312 diff_2891_3211# diff_2488_3064# diff_2899_3019# GND efet w=76 l=14
+ ad=0 pd=0 as=0 ps=0 
M2313 diff_2593_3005# diff_2584_2299# diff_2500_3043# GND efet w=70 l=13
+ ad=0 pd=0 as=0 ps=0 
M2314 diff_2791_3002# diff_2584_2299# diff_2695_3019# GND efet w=83 l=14
+ ad=0 pd=0 as=0 ps=0 
M2315 diff_2995_3005# diff_2584_2299# diff_2899_3019# GND efet w=82 l=19
+ ad=0 pd=0 as=0 ps=0 
M2316 diff_3196_3005# diff_2584_2299# diff_3100_3022# GND efet w=82 l=17
+ ad=0 pd=0 as=0 ps=0 
M2317 diff_3400_3002# diff_2584_2299# diff_3304_3022# GND efet w=85 l=13
+ ad=0 pd=0 as=0 ps=0 
M2318 diff_3607_3005# diff_2584_2299# diff_3511_3016# GND efet w=82 l=17
+ ad=0 pd=0 as=0 ps=0 
M2319 diff_4115_3211# diff_2488_3064# diff_4123_3016# GND efet w=76 l=14
+ ad=0 pd=0 as=0 ps=0 
M2320 diff_3811_3005# diff_2584_2299# diff_3715_3016# GND efet w=83 l=19
+ ad=0 pd=0 as=0 ps=0 
M2321 diff_4319_3211# diff_2488_3064# diff_4330_3019# GND efet w=73 l=13
+ ad=0 pd=0 as=0 ps=0 
M2322 diff_4523_3211# diff_2488_3064# diff_4534_3019# GND efet w=74 l=14
+ ad=0 pd=0 as=0 ps=0 
M2323 diff_4727_3211# diff_2488_3064# diff_4735_3019# GND efet w=74 l=14
+ ad=0 pd=0 as=0 ps=0 
M2324 diff_4931_3211# diff_2488_3064# diff_4939_3019# GND efet w=76 l=14
+ ad=0 pd=0 as=0 ps=0 
M2325 diff_5135_3211# diff_2488_3064# diff_5143_3019# GND efet w=74 l=14
+ ad=0 pd=0 as=0 ps=0 
M2326 diff_4015_3005# diff_2584_2299# diff_3919_3016# GND efet w=82 l=17
+ ad=0 pd=0 as=0 ps=0 
M2327 diff_4219_3005# diff_2584_2299# diff_4123_3016# GND efet w=82 l=19
+ ad=0 pd=0 as=0 ps=0 
M2328 diff_4426_3005# diff_2584_2299# diff_4330_3019# GND efet w=80 l=17
+ ad=0 pd=0 as=0 ps=0 
M2329 diff_4630_3005# diff_2584_2299# diff_4534_3019# GND efet w=80 l=17
+ ad=0 pd=0 as=0 ps=0 
M2330 diff_5339_3211# diff_2488_3064# diff_5347_3019# GND efet w=76 l=14
+ ad=0 pd=0 as=0 ps=0 
M2331 diff_4831_3005# diff_2584_2299# diff_4735_3019# GND efet w=82 l=19
+ ad=0 pd=0 as=0 ps=0 
M2332 diff_5035_3005# diff_2584_2299# diff_4939_3019# GND efet w=82 l=19
+ ad=0 pd=0 as=0 ps=0 
M2333 diff_5543_3211# diff_2488_3064# diff_5554_3016# GND efet w=70 l=13
+ ad=0 pd=0 as=0 ps=0 
M2334 diff_5239_3005# diff_2584_2299# diff_5143_3019# GND efet w=82 l=19
+ ad=0 pd=0 as=0 ps=0 
M2335 diff_5443_3005# diff_2584_2299# diff_5347_3019# GND efet w=82 l=19
+ ad=0 pd=0 as=0 ps=0 
M2336 diff_5650_3005# diff_2584_2299# diff_5554_3016# GND efet w=77 l=17
+ ad=0 pd=0 as=0 ps=0 
M2337 GND diff_841_2926# diff_844_2719# GND efet w=139 l=13
+ ad=0 pd=0 as=6708 ps=640 
M2338 GND diff_1231_2926# diff_1234_2719# GND efet w=139 l=13
+ ad=0 pd=0 as=6712 ps=632 
M2339 Vdd Vdd diff_844_2719# GND efet w=16 l=31
+ ad=0 pd=0 as=0 ps=0 
M2340 GND diff_1618_2926# diff_1621_2719# GND efet w=139 l=13
+ ad=0 pd=0 as=7051 ps=644 
M2341 diff_844_2719# diff_844_2719# diff_844_2719# GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M2342 diff_844_2719# diff_844_2719# diff_844_2719# GND efet w=7 l=7
+ ad=0 pd=0 as=0 ps=0 
M2343 Vdd Vdd diff_1234_2719# GND efet w=16 l=25
+ ad=0 pd=0 as=0 ps=0 
M2344 GND diff_2005_2926# diff_2008_2719# GND efet w=139 l=13
+ ad=0 pd=0 as=7074 ps=658 
M2345 diff_1234_2719# diff_1234_2719# diff_1234_2719# GND efet w=7 l=8
+ ad=0 pd=0 as=0 ps=0 
M2346 Vdd Vdd diff_1621_2719# GND efet w=16 l=25
+ ad=0 pd=0 as=0 ps=0 
M2347 diff_2686_2951# diff_2659_2353# diff_2500_3043# GND efet w=76 l=13
+ ad=0 pd=0 as=0 ps=0 
M2348 diff_2890_2951# diff_2659_2353# diff_2695_3019# GND efet w=76 l=13
+ ad=0 pd=0 as=0 ps=0 
M2349 diff_3091_2951# diff_2659_2353# diff_2899_3019# GND efet w=76 l=13
+ ad=0 pd=0 as=0 ps=0 
M2350 diff_3295_2951# diff_2659_2353# diff_3100_3022# GND efet w=76 l=13
+ ad=0 pd=0 as=0 ps=0 
M2351 diff_3502_2951# diff_2659_2353# diff_3304_3022# GND efet w=76 l=13
+ ad=0 pd=0 as=0 ps=0 
M2352 diff_3706_2951# diff_2659_2353# diff_3511_3016# GND efet w=76 l=13
+ ad=0 pd=0 as=0 ps=0 
M2353 diff_3910_2951# diff_2659_2353# diff_3715_3016# GND efet w=76 l=13
+ ad=0 pd=0 as=0 ps=0 
M2354 diff_4114_2951# diff_2659_2353# diff_3919_3016# GND efet w=76 l=13
+ ad=0 pd=0 as=0 ps=0 
M2355 diff_4321_2951# diff_2659_2353# diff_4123_3016# GND efet w=76 l=13
+ ad=0 pd=0 as=0 ps=0 
M2356 diff_4525_2951# diff_2659_2353# diff_4330_3019# GND efet w=76 l=13
+ ad=0 pd=0 as=0 ps=0 
M2357 diff_4726_2951# diff_2659_2353# diff_4534_3019# GND efet w=76 l=13
+ ad=0 pd=0 as=0 ps=0 
M2358 diff_4930_2951# diff_2659_2353# diff_4735_3019# GND efet w=76 l=13
+ ad=0 pd=0 as=0 ps=0 
M2359 diff_5134_2951# diff_2659_2353# diff_4939_3019# GND efet w=76 l=13
+ ad=0 pd=0 as=0 ps=0 
M2360 diff_5338_2951# diff_2659_2353# diff_5143_3019# GND efet w=76 l=13
+ ad=0 pd=0 as=0 ps=0 
M2361 diff_5545_2951# diff_2659_2353# diff_5347_3019# GND efet w=73 l=13
+ ad=0 pd=0 as=0 ps=0 
M2362 diff_5747_3211# diff_2659_2353# diff_5554_3016# GND efet w=113 l=14
+ ad=0 pd=0 as=0 ps=0 
M2363 diff_1621_2719# diff_1621_2719# diff_1621_2719# GND efet w=10 l=10
+ ad=0 pd=0 as=0 ps=0 
M2364 diff_2008_2719# diff_2008_2719# diff_2008_2719# GND efet w=4 l=4
+ ad=0 pd=0 as=0 ps=0 
M2365 Vdd Vdd diff_2008_2719# GND efet w=16 l=25
+ ad=0 pd=0 as=0 ps=0 
M2366 diff_2008_2719# diff_2008_2719# diff_2008_2719# GND efet w=8 l=8
+ ad=0 pd=0 as=0 ps=0 
M2367 diff_2500_3043# diff_2530_2884# diff_2542_2420# GND efet w=100 l=16
+ ad=0 pd=0 as=21374 ps=1712 
M2368 diff_2695_3019# diff_2812_2884# diff_2542_2420# GND efet w=100 l=13
+ ad=0 pd=0 as=0 ps=0 
M2369 diff_3100_3022# diff_2812_2884# diff_2953_2462# GND efet w=100 l=13
+ ad=0 pd=0 as=20093 ps=1622 
M2370 diff_3511_3016# diff_2812_2884# diff_3358_2806# GND efet w=100 l=13
+ ad=0 pd=0 as=22502 ps=1736 
M2371 diff_3919_3016# diff_2812_2884# diff_3769_2459# GND efet w=100 l=13
+ ad=0 pd=0 as=22766 ps=1718 
M2372 diff_4330_3019# diff_2812_2884# diff_4177_2459# GND efet w=100 l=13
+ ad=0 pd=0 as=20930 ps=1634 
M2373 diff_4735_3019# diff_2812_2884# diff_4588_2459# GND efet w=100 l=13
+ ad=0 pd=0 as=20513 ps=1574 
M2374 diff_5143_3019# diff_2812_2884# diff_4993_2459# GND efet w=100 l=13
+ ad=0 pd=0 as=22622 ps=1772 
M2375 diff_5554_3016# diff_2812_2884# diff_5401_2462# GND efet w=85 l=13
+ ad=0 pd=0 as=17987 ps=1424 
M2376 Vdd diff_844_2719# io3 GND efet w=439 l=16
+ ad=0 pd=0 as=61590 ps=4820 
M2377 d3 GND d3 GND efet w=443 l=275
+ ad=0 pd=0 as=0 ps=0 
M2378 GND diff_841_2926# io3 GND efet w=449 l=19
+ ad=0 pd=0 as=0 ps=0 
M2379 Vdd diff_1234_2719# io2 GND efet w=442 l=16
+ ad=0 pd=0 as=58522 ps=4794 
M2380 io2 GND io2 GND efet w=440 l=263
+ ad=0 pd=0 as=0 ps=0 
M2381 GND diff_1231_2926# io2 GND efet w=449 l=19
+ ad=0 pd=0 as=0 ps=0 
M2382 Vdd diff_1621_2719# io1 GND efet w=442 l=16
+ ad=0 pd=0 as=56491 ps=4608 
M2383 GND diff_1618_2926# io1 GND efet w=449 l=19
+ ad=0 pd=0 as=0 ps=0 
M2384 Vdd diff_2008_2719# io0 GND efet w=439 l=16
+ ad=0 pd=0 as=58402 ps=4818 
M2385 diff_1243_2417# diff_1018_1732# diff_1021_3622# GND efet w=55 l=16
+ ad=5341 pd=580 as=7119 ps=812 
M2386 diff_1358_2545# diff_1117_2257# diff_1243_2417# GND efet w=55 l=16
+ ad=6557 pd=608 as=0 ps=0 
M2387 diff_1621_2417# diff_1018_1732# diff_1408_3622# GND efet w=55 l=16
+ ad=5737 pd=604 as=5751 ps=650 
M2388 diff_1706_2587# diff_1117_2257# diff_1621_2417# GND efet w=55 l=16
+ ad=6284 pd=536 as=0 ps=0 
M2389 io1 GND io1 GND efet w=419 l=308
+ ad=0 pd=0 as=0 ps=0 
M2390 io3 GND io3 GND efet w=372 l=172
+ ad=0 pd=0 as=0 ps=0 
M2391 diff_1243_2417# diff_1030_2168# io3 GND efet w=52 l=13
+ ad=0 pd=0 as=0 ps=0 
M2392 GND diff_2005_2926# io0 GND efet w=449 l=19
+ ad=0 pd=0 as=0 ps=0 
M2393 diff_2899_3019# diff_2530_2884# diff_2953_2462# GND efet w=97 l=16
+ ad=0 pd=0 as=0 ps=0 
M2394 diff_3304_3022# diff_2530_2884# diff_3358_2806# GND efet w=100 l=16
+ ad=0 pd=0 as=0 ps=0 
M2395 diff_3715_3016# diff_2530_2884# diff_3769_2459# GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2396 diff_4123_3016# diff_2530_2884# diff_4177_2459# GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2397 diff_4534_3019# diff_2530_2884# diff_4588_2459# GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2398 diff_4939_3019# diff_2530_2884# diff_4993_2459# GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2399 diff_5347_3019# diff_2530_2884# diff_5401_2462# GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2400 diff_2254_2420# diff_1018_1732# diff_2185_3622# GND efet w=52 l=16
+ ad=8908 pd=1012 as=1698 ps=170 
M2401 diff_2417_2710# diff_1117_2257# diff_2254_2420# GND efet w=52 l=16
+ ad=4499 pd=402 as=0 ps=0 
M2402 diff_2008_2417# diff_1018_1732# diff_1798_3622# GND efet w=55 l=16
+ ad=6154 pd=664 as=5076 ps=578 
M2403 diff_2072_2599# diff_1117_2257# diff_2008_2417# GND efet w=55 l=16
+ ad=9719 pd=854 as=0 ps=0 
M2404 io0 GND io0 GND efet w=445 l=319
+ ad=0 pd=0 as=0 ps=0 
M2405 io3 GND io3 GND efet w=69 l=82
+ ad=0 pd=0 as=0 ps=0 
M2406 GND diff_1030_2168# diff_1117_2257# GND efet w=40 l=16
+ ad=0 pd=0 as=7424 ps=1060 
M2407 diff_1235_2224# io3 GND GND efet w=85 l=16
+ ad=5140 pd=460 as=0 ps=0 
M2408 GND io3 diff_1235_2224# GND efet w=85 l=16
+ ad=0 pd=0 as=0 ps=0 
M2409 diff_1621_2417# diff_1030_2168# io2 GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2410 io3 Vdd Vdd GND efet w=19 l=28
+ ad=0 pd=0 as=0 ps=0 
M2411 diff_1030_2168# diff_1030_2168# diff_1030_2168# GND efet w=0 l=1
+ ad=11099 pd=1352 as=0 ps=0 
M2412 diff_1420_2140# diff_1420_2140# diff_1420_2140# GND efet w=3 l=7
+ ad=1159 pd=188 as=0 ps=0 
M2413 diff_1030_2168# diff_1030_2168# diff_1030_2168# GND efet w=0 l=1
+ ad=0 pd=0 as=0 ps=0 
M2414 diff_1420_2140# diff_1420_2140# diff_1420_2140# GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M2415 diff_1030_2168# diff_1030_2168# diff_1030_2168# GND efet w=2 l=6
+ ad=0 pd=0 as=0 ps=0 
M2416 diff_1616_2221# io2 GND GND efet w=85 l=16
+ ad=5188 pd=466 as=0 ps=0 
M2417 GND io2 diff_1616_2221# GND efet w=85 l=16
+ ad=0 pd=0 as=0 ps=0 
M2418 diff_2953_2462# diff_1411_1187# diff_2500_2719# GND efet w=55 l=13
+ ad=0 pd=0 as=9307 ps=812 
M2419 diff_2417_2710# diff_2500_2719# GND GND efet w=124 l=13
+ ad=0 pd=0 as=0 ps=0 
M2420 diff_2500_2719# diff_2500_2719# diff_2500_2719# GND efet w=1 l=1
+ ad=0 pd=0 as=0 ps=0 
M2421 diff_2417_2710# Vdd Vdd GND efet w=22 l=61
+ ad=0 pd=0 as=0 ps=0 
M2422 diff_2500_2719# diff_2500_2719# diff_2500_2719# GND efet w=1 l=3
+ ad=0 pd=0 as=0 ps=0 
M2423 diff_3769_2459# diff_1411_1187# diff_3361_2519# GND efet w=58 l=13
+ ad=0 pd=0 as=8866 ps=776 
M2424 diff_4588_2459# diff_1411_1187# diff_4177_2519# GND efet w=52 l=13
+ ad=0 pd=0 as=10725 ps=826 
M2425 Vdd Vdd Vdd GND efet w=4 l=5
+ ad=0 pd=0 as=0 ps=0 
M2426 Vdd Vdd Vdd GND efet w=4 l=5
+ ad=0 pd=0 as=0 ps=0 
M2427 diff_1117_2257# diff_1117_2257# diff_1117_2257# GND efet w=6 l=13
+ ad=0 pd=0 as=0 ps=0 
M2428 Vdd Vdd Vdd GND efet w=2 l=15
+ ad=0 pd=0 as=0 ps=0 
M2429 Vdd Vdd diff_2953_2462# GND efet w=14 l=161
+ ad=0 pd=0 as=0 ps=0 
M2430 Vdd Vdd diff_2542_2420# GND efet w=13 l=163
+ ad=0 pd=0 as=0 ps=0 
M2431 Vdd Vdd Vdd GND efet w=2 l=10
+ ad=0 pd=0 as=0 ps=0 
M2432 diff_3361_2519# diff_3361_2519# diff_3361_2519# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M2433 diff_3361_2519# diff_3361_2519# diff_3361_2519# GND efet w=1 l=3
+ ad=0 pd=0 as=0 ps=0 
M2434 diff_3769_2459# Vdd Vdd GND efet w=14 l=157
+ ad=0 pd=0 as=0 ps=0 
M2435 Vdd Vdd diff_2072_2599# GND efet w=19 l=58
+ ad=0 pd=0 as=0 ps=0 
M2436 Vdd Vdd Vdd GND efet w=2 l=9
+ ad=0 pd=0 as=0 ps=0 
M2437 Vdd Vdd diff_3358_2806# GND efet w=13 l=161
+ ad=0 pd=0 as=0 ps=0 
M2438 Vdd Vdd Vdd GND efet w=5 l=10
+ ad=0 pd=0 as=0 ps=0 
M2439 diff_2072_2599# diff_3361_2519# GND GND efet w=103 l=16
+ ad=0 pd=0 as=0 ps=0 
M2440 diff_4177_2459# Vdd Vdd GND efet w=14 l=167
+ ad=0 pd=0 as=0 ps=0 
M2441 Vdd Vdd diff_1706_2587# GND efet w=19 l=97
+ ad=0 pd=0 as=0 ps=0 
M2442 diff_5401_2462# diff_1411_1187# diff_4993_2519# GND efet w=58 l=16
+ ad=0 pd=0 as=10317 ps=796 
M2443 diff_4588_2459# Vdd Vdd GND efet w=11 l=164
+ ad=0 pd=0 as=0 ps=0 
M2444 diff_1706_2587# diff_4177_2519# GND GND efet w=124 l=13
+ ad=0 pd=0 as=0 ps=0 
M2445 diff_3361_2519# diff_1561_1187# diff_3358_2806# GND efet w=55 l=13
+ ad=0 pd=0 as=0 ps=0 
M2446 Vdd Vdd Vdd GND efet w=2 l=7
+ ad=0 pd=0 as=0 ps=0 
M2447 diff_4177_2519# diff_1561_1187# diff_4177_2459# GND efet w=58 l=13
+ ad=0 pd=0 as=0 ps=0 
M2448 diff_4993_2459# Vdd Vdd GND efet w=16 l=167
+ ad=0 pd=0 as=0 ps=0 
M2449 diff_4993_2519# diff_1561_1187# diff_4993_2459# GND efet w=58 l=13
+ ad=0 pd=0 as=0 ps=0 
M2450 Vdd Vdd diff_1358_2545# GND efet w=19 l=61
+ ad=0 pd=0 as=0 ps=0 
M2451 diff_5401_2462# Vdd Vdd GND efet w=16 l=175
+ ad=0 pd=0 as=0 ps=0 
M2452 diff_1358_2545# diff_4993_2519# GND GND efet w=100 l=13
+ ad=0 pd=0 as=0 ps=0 
M2453 Vdd Vdd diff_1117_2257# GND efet w=16 l=109
+ ad=0 pd=0 as=0 ps=0 
M2454 diff_1117_2257# diff_1117_2257# diff_1117_2257# GND efet w=3 l=13
+ ad=0 pd=0 as=0 ps=0 
M2455 diff_2500_2719# diff_1561_1187# diff_2542_2420# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2456 diff_2008_2417# diff_1030_2168# io1 GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2457 diff_2254_2420# diff_1030_2168# io0 GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2458 io2 Vdd Vdd GND efet w=19 l=28
+ ad=0 pd=0 as=0 ps=0 
M2459 diff_1420_2140# Vdd Vdd GND efet w=16 l=16
+ ad=0 pd=0 as=0 ps=0 
M2460 diff_1030_2168# clk1 diff_1030_2134# GND efet w=25 l=16
+ ad=0 pd=0 as=1657 ps=268 
M2461 diff_1030_2134# diff_1030_2134# diff_1030_2134# GND efet w=3 l=8
+ ad=0 pd=0 as=0 ps=0 
M2462 GND diff_1030_2134# diff_1117_2257# GND efet w=89 l=14
+ ad=0 pd=0 as=0 ps=0 
M2463 Vdd Vdd diff_1235_2224# GND efet w=16 l=52
+ ad=0 pd=0 as=0 ps=0 
M2464 diff_1030_2134# diff_1030_2134# diff_1030_2134# GND efet w=2 l=4
+ ad=0 pd=0 as=0 ps=0 
M2465 Vdd Vdd Vdd GND efet w=2 l=6
+ ad=0 pd=0 as=0 ps=0 
M2466 Vdd diff_1420_2140# diff_1030_2168# GND efet w=20 l=52
+ ad=0 pd=0 as=0 ps=0 
M2467 Vdd Vdd diff_1202_2005# GND efet w=16 l=34
+ ad=0 pd=0 as=5053 ps=548 
M2468 diff_2003_2221# io1 GND GND efet w=85 l=16
+ ad=5140 pd=460 as=0 ps=0 
M2469 GND io1 diff_2003_2221# GND efet w=85 l=16
+ ad=0 pd=0 as=0 ps=0 
M2470 diff_2953_2462# diff_2536_2407# diff_2899_2270# GND efet w=97 l=16
+ ad=0 pd=0 as=10284 ps=1114 
M2471 diff_3358_2806# diff_2536_2407# diff_3304_2261# GND efet w=95 l=14
+ ad=0 pd=0 as=10419 ps=1132 
M2472 diff_3769_2459# diff_2536_2407# diff_3715_2267# GND efet w=97 l=13
+ ad=0 pd=0 as=10866 ps=1138 
M2473 diff_4177_2459# diff_2536_2407# diff_4123_2270# GND efet w=97 l=13
+ ad=0 pd=0 as=10668 ps=1126 
M2474 diff_2542_2420# diff_2536_2407# diff_2500_2240# GND efet w=100 l=16
+ ad=0 pd=0 as=11928 ps=1162 
M2475 diff_2542_2420# diff_2812_2410# diff_2695_2267# GND efet w=100 l=13
+ ad=0 pd=0 as=10007 ps=996 
M2476 diff_2953_2462# diff_2812_2410# diff_3100_2267# GND efet w=100 l=13
+ ad=0 pd=0 as=9578 ps=984 
M2477 diff_3358_2806# diff_2812_2410# diff_3511_2267# GND efet w=100 l=13
+ ad=0 pd=0 as=10328 ps=1008 
M2478 diff_3769_2459# diff_2812_2410# diff_3919_2267# GND efet w=100 l=13
+ ad=0 pd=0 as=10328 ps=1008 
M2479 diff_4588_2459# diff_2536_2407# diff_4534_2270# GND efet w=97 l=13
+ ad=0 pd=0 as=10542 ps=1120 
M2480 diff_4177_2459# diff_2812_2410# diff_4330_2267# GND efet w=100 l=13
+ ad=0 pd=0 as=10019 ps=996 
M2481 diff_4993_2459# diff_2536_2407# diff_4939_2270# GND efet w=97 l=13
+ ad=0 pd=0 as=10512 ps=1120 
M2482 diff_5401_2462# diff_2536_2407# diff_5347_2270# GND efet w=100 l=16
+ ad=0 pd=0 as=10392 ps=1126 
M2483 diff_4588_2459# diff_2812_2410# diff_4735_2267# GND efet w=100 l=13
+ ad=0 pd=0 as=9989 ps=996 
M2484 diff_4993_2459# diff_2812_2410# diff_5143_2267# GND efet w=100 l=13
+ ad=0 pd=0 as=9989 ps=996 
M2485 diff_5401_2462# diff_2812_2410# diff_5554_2267# GND efet w=85 l=10
+ ad=0 pd=0 as=10430 ps=1036 
M2486 diff_5747_2072# diff_2659_2353# diff_5554_2267# GND efet w=107 l=14
+ ad=5199 pd=612 as=0 ps=0 
M2487 diff_2500_2240# diff_2659_2353# diff_2686_2320# GND efet w=76 l=13
+ ad=0 pd=0 as=4293 ps=436 
M2488 diff_2695_2267# diff_2659_2353# diff_2890_2320# GND efet w=76 l=13
+ ad=0 pd=0 as=4329 ps=436 
M2489 diff_2899_2270# diff_2659_2353# diff_3091_2317# GND efet w=76 l=13
+ ad=0 pd=0 as=4521 ps=442 
M2490 diff_3100_2267# diff_2659_2353# diff_3295_2317# GND efet w=76 l=13
+ ad=0 pd=0 as=4557 ps=442 
M2491 diff_3304_2261# diff_2659_2353# diff_3502_2323# GND efet w=76 l=13
+ ad=0 pd=0 as=4065 ps=430 
M2492 diff_3511_2267# diff_2659_2353# diff_3706_2323# GND efet w=76 l=13
+ ad=0 pd=0 as=4101 ps=430 
M2493 diff_3715_2267# diff_2659_2353# diff_3910_2323# GND efet w=76 l=13
+ ad=0 pd=0 as=4065 ps=430 
M2494 diff_3919_2267# diff_2659_2353# diff_4114_2323# GND efet w=76 l=13
+ ad=0 pd=0 as=4101 ps=430 
M2495 diff_4123_2270# diff_2659_2353# diff_4321_2320# GND efet w=76 l=13
+ ad=0 pd=0 as=4293 ps=436 
M2496 diff_4330_2267# diff_2659_2353# diff_4525_2320# GND efet w=76 l=13
+ ad=0 pd=0 as=4329 ps=436 
M2497 diff_4534_2270# diff_2659_2353# diff_4726_2320# GND efet w=76 l=13
+ ad=0 pd=0 as=4293 ps=436 
M2498 diff_4735_2267# diff_2659_2353# diff_4930_2320# GND efet w=76 l=13
+ ad=0 pd=0 as=4329 ps=436 
M2499 diff_4939_2270# diff_2659_2353# diff_5134_2320# GND efet w=76 l=13
+ ad=0 pd=0 as=4293 ps=436 
M2500 diff_5143_2267# diff_2659_2353# diff_5338_2320# GND efet w=76 l=13
+ ad=0 pd=0 as=4329 ps=436 
M2501 diff_5347_2270# diff_2659_2353# diff_5545_2320# GND efet w=73 l=13
+ ad=0 pd=0 as=4230 ps=430 
M2502 io1 Vdd Vdd GND efet w=19 l=28
+ ad=0 pd=0 as=0 ps=0 
M2503 diff_2246_2221# io0 GND GND efet w=85 l=16
+ ad=5188 pd=466 as=0 ps=0 
M2504 GND io0 diff_2246_2221# GND efet w=85 l=16
+ ad=0 pd=0 as=0 ps=0 
M2505 io0 Vdd Vdd GND efet w=19 l=28
+ ad=0 pd=0 as=0 ps=0 
M2506 Vdd Vdd diff_1616_2221# GND efet w=16 l=55
+ ad=0 pd=0 as=0 ps=0 
M2507 Vdd Vdd diff_2003_2221# GND efet w=16 l=52
+ ad=0 pd=0 as=0 ps=0 
M2508 Vdd Vdd diff_2246_2221# GND efet w=16 l=49
+ ad=0 pd=0 as=0 ps=0 
M2509 diff_1030_2168# diff_1420_2140# diff_1030_2168# GND efet w=114 l=6
+ ad=0 pd=0 as=0 ps=0 
M2510 GND diff_1243_1996# diff_1202_2005# GND efet w=151 l=16
+ ad=0 pd=0 as=0 ps=0 
M2511 diff_1202_2005# diff_1018_1732# diff_1120_1930# GND efet w=28 l=16
+ ad=0 pd=0 as=972 ps=128 
M2512 diff_2695_2267# diff_2584_2299# diff_2791_2269# GND efet w=83 l=14
+ ad=0 pd=0 as=4803 ps=490 
M2513 diff_2899_2270# diff_2584_2299# diff_2995_2269# GND efet w=82 l=19
+ ad=0 pd=0 as=4905 ps=490 
M2514 diff_3304_2261# diff_2584_2299# diff_3400_2266# GND efet w=85 l=13
+ ad=0 pd=0 as=5142 ps=502 
M2515 diff_3100_2267# diff_2584_2299# diff_3196_2266# GND efet w=82 l=17
+ ad=0 pd=0 as=5022 ps=490 
M2516 diff_3511_2267# diff_2584_2299# diff_3607_2272# GND efet w=82 l=17
+ ad=0 pd=0 as=4566 ps=478 
M2517 diff_3715_2267# diff_2584_2299# diff_3811_2272# GND efet w=83 l=19
+ ad=0 pd=0 as=4677 ps=484 
M2518 diff_3919_2267# diff_2584_2299# diff_4015_2272# GND efet w=82 l=17
+ ad=0 pd=0 as=4566 ps=478 
M2519 diff_4123_2270# diff_2584_2299# diff_4219_2272# GND efet w=82 l=19
+ ad=0 pd=0 as=4677 ps=484 
M2520 diff_4330_2267# diff_2584_2299# diff_4426_2269# GND efet w=80 l=17
+ ad=0 pd=0 as=4794 ps=484 
M2521 diff_4534_2270# diff_2584_2299# diff_4630_2269# GND efet w=80 l=17
+ ad=0 pd=0 as=4905 ps=490 
M2522 diff_4735_2267# diff_2584_2299# diff_4831_2269# GND efet w=82 l=19
+ ad=0 pd=0 as=4794 ps=484 
M2523 diff_4939_2270# diff_2584_2299# diff_5035_2269# GND efet w=82 l=19
+ ad=0 pd=0 as=4905 ps=490 
M2524 diff_5143_2267# diff_2584_2299# diff_5239_2269# GND efet w=82 l=19
+ ad=0 pd=0 as=4794 ps=484 
M2525 diff_5347_2270# diff_2584_2299# diff_5443_2269# GND efet w=82 l=19
+ ad=0 pd=0 as=4905 ps=490 
M2526 diff_5554_2267# diff_2584_2299# diff_5650_2269# GND efet w=79 l=19
+ ad=0 pd=0 as=4647 ps=478 
M2527 diff_1030_2168# diff_1030_2168# diff_1030_2168# GND efet w=1 l=1
+ ad=0 pd=0 as=0 ps=0 
M2528 diff_2500_2240# diff_2584_2299# diff_2593_2260# GND efet w=70 l=13
+ ad=0 pd=0 as=4752 ps=478 
M2529 diff_2695_2267# diff_2488_3064# diff_2687_2066# GND efet w=74 l=14
+ ad=0 pd=0 as=4074 ps=466 
M2530 diff_2899_2270# diff_2488_3064# diff_2891_2072# GND efet w=76 l=14
+ ad=0 pd=0 as=4206 ps=466 
M2531 diff_3100_2267# diff_2488_3064# diff_3095_2072# GND efet w=76 l=14
+ ad=0 pd=0 as=4170 ps=466 
M2532 diff_3304_2261# diff_2488_3064# diff_3299_2072# GND efet w=83 l=13
+ ad=0 pd=0 as=4374 ps=472 
M2533 diff_3511_2267# diff_2488_3064# diff_3503_2072# GND efet w=76 l=14
+ ad=0 pd=0 as=3807 ps=460 
M2534 diff_3715_2267# diff_2488_3064# diff_3707_2072# GND efet w=79 l=13
+ ad=0 pd=0 as=3966 ps=460 
M2535 diff_3919_2267# diff_2488_3064# diff_3911_2072# GND efet w=76 l=14
+ ad=0 pd=0 as=3807 ps=460 
M2536 diff_4123_2270# diff_2488_3064# diff_4115_2072# GND efet w=76 l=14
+ ad=0 pd=0 as=3987 ps=460 
M2537 diff_4330_2267# diff_2488_3064# diff_4319_2072# GND efet w=73 l=13
+ ad=0 pd=0 as=4041 ps=466 
M2538 diff_4534_2270# diff_2488_3064# diff_4523_2072# GND efet w=74 l=14
+ ad=0 pd=0 as=4218 ps=466 
M2539 diff_2500_2240# diff_2488_3064# diff_2494_2092# GND efet w=94 l=10
+ ad=0 pd=0 as=5093 ps=486 
M2540 diff_4735_2267# diff_2488_3064# diff_4727_2072# GND efet w=74 l=14
+ ad=0 pd=0 as=4038 ps=466 
M2541 diff_4939_2270# diff_2488_3064# diff_4931_2072# GND efet w=76 l=14
+ ad=0 pd=0 as=4206 ps=466 
M2542 diff_5143_2267# diff_2488_3064# diff_5135_2072# GND efet w=74 l=14
+ ad=0 pd=0 as=4038 ps=466 
M2543 diff_5347_2270# diff_2488_3064# diff_5339_2072# GND efet w=76 l=14
+ ad=0 pd=0 as=4206 ps=466 
M2544 diff_5554_2267# diff_2488_3064# diff_5543_2072# GND efet w=70 l=13
+ ad=0 pd=0 as=3921 ps=454 
M2545 diff_2582_2126# diff_2563_2125# GND GND efet w=114 l=15
+ ad=2399 pd=264 as=0 ps=0 
M2546 diff_1030_2168# diff_1030_2168# diff_1030_2168# GND efet w=0 l=1
+ ad=0 pd=0 as=0 ps=0 
M2547 GND diff_1120_1930# diff_475_2011# GND efet w=226 l=16
+ ad=0 pd=0 as=31376 ps=2928 
M2548 diff_475_2011# diff_1054_1822# Vdd GND efet w=206 l=14
+ ad=0 pd=0 as=0 ps=0 
M2549 diff_1394_1915# diff_1024_1190# diff_1342_1942# GND efet w=88 l=16
+ ad=5408 pd=562 as=5237 ps=548 
M2550 diff_1342_1942# diff_850_1331# diff_1243_1996# GND efet w=97 l=16
+ ad=0 pd=0 as=3614 ps=378 
M2551 GND diff_2521_1937# diff_2494_2092# GND efet w=70 l=13
+ ad=0 pd=0 as=0 ps=0 
M2552 diff_2500_2240# diff_2623_2116# diff_2582_2126# GND efet w=76 l=13
+ ad=0 pd=0 as=0 ps=0 
M2553 GND diff_2725_1937# diff_2686_2320# GND efet w=86 l=16
+ ad=0 pd=0 as=0 ps=0 
M2554 diff_2789_2123# diff_2776_1937# GND GND efet w=88 l=16
+ ad=2159 pd=234 as=0 ps=0 
M2555 diff_2695_2267# diff_2623_2116# diff_2789_2123# GND efet w=73 l=13
+ ad=0 pd=0 as=0 ps=0 
M2556 GND diff_2929_1937# diff_2890_2320# GND efet w=86 l=16
+ ad=0 pd=0 as=0 ps=0 
M2557 diff_2993_2123# diff_2980_1937# GND GND efet w=88 l=16
+ ad=2159 pd=234 as=0 ps=0 
M2558 diff_2899_2270# diff_2623_2116# diff_2993_2123# GND efet w=73 l=13
+ ad=0 pd=0 as=0 ps=0 
M2559 GND diff_3133_1937# diff_3091_2317# GND efet w=86 l=16
+ ad=0 pd=0 as=0 ps=0 
M2560 diff_3197_2123# diff_3184_1937# GND GND efet w=88 l=16
+ ad=2159 pd=234 as=0 ps=0 
M2561 diff_3100_2267# diff_2623_2116# diff_3197_2123# GND efet w=73 l=13
+ ad=0 pd=0 as=0 ps=0 
M2562 GND diff_3337_1937# diff_3295_2317# GND efet w=86 l=16
+ ad=0 pd=0 as=0 ps=0 
M2563 diff_3401_2123# diff_3388_1937# GND GND efet w=88 l=16
+ ad=2159 pd=234 as=0 ps=0 
M2564 diff_3304_2261# diff_2623_2116# diff_3401_2123# GND efet w=73 l=13
+ ad=0 pd=0 as=0 ps=0 
M2565 GND diff_3541_1937# diff_3502_2323# GND efet w=86 l=16
+ ad=0 pd=0 as=0 ps=0 
M2566 diff_3605_2123# diff_3592_1937# GND GND efet w=88 l=16
+ ad=2159 pd=234 as=0 ps=0 
M2567 diff_3511_2267# diff_2623_2116# diff_3605_2123# GND efet w=73 l=13
+ ad=0 pd=0 as=0 ps=0 
M2568 GND diff_3745_1937# diff_3706_2323# GND efet w=86 l=16
+ ad=0 pd=0 as=0 ps=0 
M2569 diff_3809_2123# diff_3796_1937# GND GND efet w=88 l=16
+ ad=2159 pd=234 as=0 ps=0 
M2570 diff_3715_2267# diff_2623_2116# diff_3809_2123# GND efet w=73 l=13
+ ad=0 pd=0 as=0 ps=0 
M2571 GND diff_3949_1937# diff_3910_2323# GND efet w=86 l=16
+ ad=0 pd=0 as=0 ps=0 
M2572 diff_4013_2123# diff_4000_1937# GND GND efet w=88 l=16
+ ad=2159 pd=234 as=0 ps=0 
M2573 diff_3919_2267# diff_2623_2116# diff_4013_2123# GND efet w=73 l=13
+ ad=0 pd=0 as=0 ps=0 
M2574 GND diff_4153_1937# diff_4114_2323# GND efet w=86 l=16
+ ad=0 pd=0 as=0 ps=0 
M2575 diff_4217_2123# diff_4204_1937# GND GND efet w=88 l=16
+ ad=2159 pd=234 as=0 ps=0 
M2576 diff_4123_2270# diff_2623_2116# diff_4217_2123# GND efet w=73 l=13
+ ad=0 pd=0 as=0 ps=0 
M2577 GND diff_4357_1937# diff_4321_2320# GND efet w=86 l=16
+ ad=0 pd=0 as=0 ps=0 
M2578 diff_4421_2123# diff_4408_1937# GND GND efet w=88 l=16
+ ad=2159 pd=234 as=0 ps=0 
M2579 diff_4330_2267# diff_2623_2116# diff_4421_2123# GND efet w=73 l=13
+ ad=0 pd=0 as=0 ps=0 
M2580 GND diff_4561_1937# diff_4525_2320# GND efet w=86 l=16
+ ad=0 pd=0 as=0 ps=0 
M2581 diff_4625_2123# diff_4612_1937# GND GND efet w=88 l=16
+ ad=2159 pd=234 as=0 ps=0 
M2582 diff_4534_2270# diff_2623_2116# diff_4625_2123# GND efet w=73 l=13
+ ad=0 pd=0 as=0 ps=0 
M2583 GND diff_4765_1937# diff_4726_2320# GND efet w=86 l=16
+ ad=0 pd=0 as=0 ps=0 
M2584 diff_4829_2123# diff_4816_1937# GND GND efet w=88 l=16
+ ad=2159 pd=234 as=0 ps=0 
M2585 diff_4735_2267# diff_2623_2116# diff_4829_2123# GND efet w=73 l=13
+ ad=0 pd=0 as=0 ps=0 
M2586 GND diff_4969_1937# diff_4930_2320# GND efet w=86 l=16
+ ad=0 pd=0 as=0 ps=0 
M2587 diff_5033_2123# diff_5020_1937# GND GND efet w=88 l=16
+ ad=2159 pd=234 as=0 ps=0 
M2588 diff_4939_2270# diff_2623_2116# diff_5033_2123# GND efet w=73 l=13
+ ad=0 pd=0 as=0 ps=0 
M2589 GND diff_5173_1937# diff_5134_2320# GND efet w=86 l=16
+ ad=0 pd=0 as=0 ps=0 
M2590 diff_5237_2123# diff_5224_1937# GND GND efet w=88 l=16
+ ad=2159 pd=234 as=0 ps=0 
M2591 diff_5143_2267# diff_2623_2116# diff_5237_2123# GND efet w=73 l=13
+ ad=0 pd=0 as=0 ps=0 
M2592 GND diff_5377_1937# diff_5338_2320# GND efet w=86 l=16
+ ad=0 pd=0 as=0 ps=0 
M2593 diff_5441_2123# diff_5428_1937# GND GND efet w=88 l=16
+ ad=2159 pd=234 as=0 ps=0 
M2594 diff_5347_2270# diff_2623_2116# diff_5441_2123# GND efet w=73 l=13
+ ad=0 pd=0 as=0 ps=0 
M2595 GND diff_5581_1937# diff_5545_2320# GND efet w=86 l=16
+ ad=0 pd=0 as=0 ps=0 
M2596 diff_5645_2123# diff_5632_1937# GND GND efet w=88 l=16
+ ad=2159 pd=234 as=0 ps=0 
M2597 diff_5554_2267# diff_2623_2116# diff_5645_2123# GND efet w=73 l=13
+ ad=0 pd=0 as=0 ps=0 
M2598 diff_6479_3832# Vdd Vdd GND efet w=31 l=16
+ ad=961 pd=136 as=0 ps=0 
M2599 diff_6479_3832# diff_6479_3832# diff_6479_3832# GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M2600 diff_6479_3832# diff_6479_3832# diff_6479_3832# GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M2601 Vdd Vdd Vdd GND efet w=0 l=1
+ ad=0 pd=0 as=0 ps=0 
M2602 GND diff_6919_3958# diff_6625_3799# GND efet w=199 l=13
+ ad=0 pd=0 as=8083 ps=630 
M2603 Vdd Vdd diff_6625_3799# GND efet w=19 l=40
+ ad=0 pd=0 as=0 ps=0 
M2604 Vdd Vdd Vdd GND efet w=0 l=1
+ ad=0 pd=0 as=0 ps=0 
M2605 GND d2 diff_7033_2509# GND efet w=487 l=13
+ ad=0 pd=0 as=12827 ps=986 
M2606 diff_7033_2509# Vdd Vdd GND efet w=19 l=40
+ ad=0 pd=0 as=0 ps=0 
M2607 diff_6625_3799# clk1 diff_6922_3853# GND efet w=31 l=13
+ ad=0 pd=0 as=1001 ps=130 
M2608 Vdd Vdd diff_7033_2836# GND efet w=19 l=40
+ ad=0 pd=0 as=6521 ps=570 
M2609 diff_6922_3853# diff_6922_3853# diff_6922_3853# GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M2610 GND diff_6922_3853# diff_6778_3391# GND efet w=109 l=13
+ ad=0 pd=0 as=0 ps=0 
M2611 Vdd Vdd diff_6778_3391# GND efet w=22 l=46
+ ad=0 pd=0 as=0 ps=0 
M2612 Vdd Vdd Vdd GND efet w=5 l=9
+ ad=0 pd=0 as=0 ps=0 
M2613 Vdd Vdd Vdd GND efet w=4 l=5
+ ad=0 pd=0 as=0 ps=0 
M2614 diff_6778_3391# clk2 diff_6922_3745# GND efet w=28 l=13
+ ad=0 pd=0 as=818 ps=116 
M2615 diff_2509_4258# diff_6473_3661# Vdd GND efet w=37 l=13
+ ad=24308 pd=1836 as=0 ps=0 
M2616 GND diff_6625_3571# diff_2509_4258# GND efet w=739 l=13
+ ad=0 pd=0 as=0 ps=0 
M2617 diff_2509_4258# diff_6473_3661# diff_2509_4258# GND efet w=99 l=11
+ ad=0 pd=0 as=0 ps=0 
M2618 diff_6473_3661# Vdd Vdd GND efet w=28 l=13
+ ad=1051 pd=142 as=0 ps=0 
M2619 diff_6473_3661# diff_6473_3661# diff_6473_3661# GND efet w=2 l=9
+ ad=0 pd=0 as=0 ps=0 
M2620 diff_6473_3661# diff_6473_3661# diff_6473_3661# GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M2621 diff_6922_3745# diff_6922_3745# diff_6922_3745# GND efet w=2 l=3
+ ad=0 pd=0 as=0 ps=0 
M2622 GND diff_6922_3745# diff_6661_3556# GND efet w=109 l=16
+ ad=0 pd=0 as=9289 ps=844 
M2623 Vdd Vdd diff_6661_3556# GND efet w=19 l=43
+ ad=0 pd=0 as=0 ps=0 
M2624 Vdd Vdd Vdd GND efet w=0 l=1
+ ad=0 pd=0 as=0 ps=0 
M2625 GND diff_7033_2509# diff_7033_2836# GND efet w=109 l=13
+ ad=0 pd=0 as=0 ps=0 
M2626 diff_6661_3556# clk1 diff_6919_3643# GND efet w=34 l=13
+ ad=0 pd=0 as=984 ps=128 
M2627 GND diff_6919_3643# diff_6808_2113# GND efet w=109 l=13
+ ad=0 pd=0 as=6797 ps=564 
M2628 Vdd Vdd diff_6808_2113# GND efet w=19 l=40
+ ad=0 pd=0 as=0 ps=0 
M2629 Vdd Vdd Vdd GND efet w=1 l=1
+ ad=0 pd=0 as=0 ps=0 
M2630 Vdd Vdd Vdd GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M2631 GND diff_6661_3556# diff_6566_3529# GND efet w=31 l=13
+ ad=0 pd=0 as=2765 ps=348 
M2632 diff_6566_3529# Vdd Vdd GND efet w=16 l=88
+ ad=0 pd=0 as=0 ps=0 
M2633 diff_6514_3431# Vdd Vdd GND efet w=16 l=43
+ ad=4373 pd=438 as=0 ps=0 
M2634 diff_6770_3481# diff_6661_3556# diff_6505_3421# GND efet w=37 l=13
+ ad=1691 pd=222 as=3084 ps=334 
M2635 diff_6514_3431# diff_6505_3421# GND GND efet w=151 l=13
+ ad=0 pd=0 as=0 ps=0 
M2636 diff_6505_3421# diff_6505_3421# diff_6505_3421# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M2637 diff_6505_3421# diff_6505_3421# diff_6505_3421# GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M2638 diff_6770_3481# diff_6535_4298# diff_6778_3391# GND efet w=31 l=13
+ ad=0 pd=0 as=0 ps=0 
M2639 diff_6505_3421# diff_6566_3529# GND GND efet w=28 l=13
+ ad=0 pd=0 as=0 ps=0 
M2640 diff_6845_3187# diff_6778_3391# diff_6316_3109# GND efet w=49 l=13
+ ad=3509 pd=338 as=1746 ps=170 
M2641 diff_6935_3271# clk2 diff_6845_3187# GND efet w=49 l=13
+ ad=6109 pd=412 as=0 ps=0 
M2642 GND diff_6421_3205# diff_2812_2884# GND efet w=349 l=13
+ ad=0 pd=0 as=11987 ps=986 
M2643 diff_6845_3187# diff_6808_2113# diff_6421_3205# GND efet w=46 l=13
+ ad=0 pd=0 as=1500 ps=158 
M2644 GND diff_1030_2168# diff_1342_1942# GND efet w=65 l=17
+ ad=0 pd=0 as=0 ps=0 
M2645 diff_1394_1915# diff_1411_1187# GND GND efet w=91 l=16
+ ad=0 pd=0 as=0 ps=0 
M2646 GND diff_1561_1187# diff_1394_1915# GND efet w=88 l=16
+ ad=0 pd=0 as=0 ps=0 
M2647 diff_2065_1957# d3 GND GND efet w=89 l=14
+ ad=5404 pd=528 as=0 ps=0 
M2648 GND diff_1751_1699# diff_1741_1957# GND efet w=52 l=16
+ ad=0 pd=0 as=2078 ps=204 
M2649 GND diff_1741_1957# diff_388_2056# GND efet w=40 l=16
+ ad=0 pd=0 as=12920 ps=1838 
M2650 diff_2039_1969# clk2 diff_1751_1699# GND efet w=25 l=16
+ ad=650 pd=102 as=2006 ps=264 
M2651 Vdd diff_2065_1957# diff_2039_1969# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M2652 diff_2065_1957# Vdd Vdd GND efet w=16 l=82
+ ad=0 pd=0 as=0 ps=0 
M2653 GND diff_1738_1391# diff_2065_1957# GND efet w=43 l=16
+ ad=0 pd=0 as=0 ps=0 
M2654 GND diff_2299_1054# diff_2065_1957# GND efet w=43 l=16
+ ad=0 pd=0 as=0 ps=0 
M2655 GND diff_2623_1937# diff_2593_2260# GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2656 diff_2687_2066# diff_2674_1937# GND GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2657 GND diff_2827_1937# diff_2791_2269# GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2658 diff_2891_2072# diff_2878_1937# GND GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2659 GND diff_3031_1937# diff_2995_2269# GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2660 diff_3095_2072# diff_3082_1937# GND GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2661 GND diff_3235_1937# diff_3196_2266# GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2662 diff_3299_2072# diff_3286_1937# GND GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2663 GND diff_3439_1937# diff_3400_2266# GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2664 diff_3503_2072# diff_3490_1937# GND GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2665 GND diff_3643_1937# diff_3607_2272# GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2666 diff_3707_2072# diff_3694_1937# GND GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2667 GND diff_3847_1937# diff_3811_2272# GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2668 diff_3911_2072# diff_3898_1937# GND GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2669 GND diff_4051_1937# diff_4015_2272# GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2670 diff_4115_2072# diff_4102_1937# GND GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2671 GND diff_4255_1937# diff_4219_2272# GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2672 diff_4319_2072# diff_4306_1937# GND GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2673 GND diff_4459_1937# diff_4426_2269# GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2674 diff_4523_2072# diff_4510_1937# GND GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2675 GND diff_4663_1937# diff_4630_2269# GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2676 diff_4727_2072# diff_4714_1937# GND GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2677 GND diff_4867_1937# diff_4831_2269# GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2678 diff_4931_2072# diff_4918_1937# GND GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2679 GND diff_5071_1937# diff_5035_2269# GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2680 diff_5135_2072# diff_5122_1937# GND GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2681 GND diff_5275_1937# diff_5239_2269# GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2682 diff_5339_2072# diff_5326_1937# GND GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2683 GND diff_5479_1937# diff_5443_2269# GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2684 diff_5543_2072# diff_5530_1937# GND GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2685 GND diff_5683_1937# diff_5650_2269# GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2686 diff_5747_2072# diff_5734_1937# GND GND efet w=97 l=13
+ ad=0 pd=0 as=0 ps=0 
M2687 GND diff_1202_2005# diff_1246_1787# GND efet w=119 l=14
+ ad=0 pd=0 as=2449 ps=316 
M2688 diff_1246_1787# diff_1018_1732# diff_1054_1822# GND efet w=25 l=13
+ ad=0 pd=0 as=1755 ps=248 
M2689 diff_1246_1787# Vdd Vdd GND efet w=16 l=37
+ ad=0 pd=0 as=0 ps=0 
M2690 Vdd Vdd Vdd GND efet w=2 l=9
+ ad=0 pd=0 as=0 ps=0 
M2691 Vdd Vdd Vdd GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M2692 Vdd Vdd diff_1243_1996# GND efet w=16 l=166
+ ad=0 pd=0 as=0 ps=0 
M2693 Vdd Vdd Vdd GND efet w=3 l=7
+ ad=0 pd=0 as=0 ps=0 
M2694 Vdd Vdd Vdd GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M2695 diff_652_1966# Vdd Vdd GND efet w=22 l=43
+ ad=5891 pd=534 as=0 ps=0 
M2696 diff_1018_1732# diff_1199_1537# Vdd GND efet w=19 l=19
+ ad=6271 pd=596 as=0 ps=0 
M2697 diff_1018_1732# diff_1199_1537# diff_1018_1732# GND efet w=112 l=57
+ ad=0 pd=0 as=0 ps=0 
M2698 diff_1199_1537# Vdd Vdd GND efet w=19 l=16
+ ad=1023 pd=140 as=0 ps=0 
M2699 Vdd Vdd diff_850_1331# GND efet w=19 l=43
+ ad=0 pd=0 as=8720 ps=732 
M2700 diff_652_1966# diff_850_1331# GND GND efet w=214 l=16
+ ad=0 pd=0 as=0 ps=0 
M2701 reset GND reset GND efet w=457 l=277
+ ad=22005 pd=2188 as=0 ps=0 
M2702 GND clk2 diff_1018_1732# GND efet w=112 l=16
+ ad=0 pd=0 as=0 ps=0 
M2703 Vdd Vdd Vdd GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M2704 diff_850_1331# reset GND GND efet w=359 l=14
+ ad=0 pd=0 as=0 ps=0 
M2705 sync clk2 diff_712_1165# GND efet w=28 l=16
+ ad=0 pd=0 as=1108 ps=146 
M2706 diff_712_1165# diff_712_1165# diff_712_1165# GND efet w=5 l=8
+ ad=0 pd=0 as=0 ps=0 
M2707 diff_712_1165# diff_712_1165# diff_712_1165# GND efet w=2 l=9
+ ad=0 pd=0 as=0 ps=0 
M2708 GND diff_712_1165# diff_724_1144# GND efet w=98 l=14
+ ad=0 pd=0 as=6514 ps=742 
M2709 Vdd Vdd Vdd GND efet w=3 l=4
+ ad=0 pd=0 as=0 ps=0 
M2710 Vdd Vdd Vdd GND efet w=0 l=1
+ ad=0 pd=0 as=0 ps=0 
M2711 Vdd Vdd diff_1024_1190# GND efet w=20 l=86
+ ad=0 pd=0 as=2297 ps=252 
M2712 Vdd Vdd diff_1226_1252# GND efet w=19 l=160
+ ad=0 pd=0 as=2569 ps=250 
M2713 diff_388_2056# diff_1738_1906# GND GND efet w=40 l=16
+ ad=0 pd=0 as=0 ps=0 
M2714 diff_388_2056# Vdd Vdd GND efet w=16 l=82
+ ad=0 pd=0 as=0 ps=0 
M2715 Vdd Vdd Vdd GND efet w=2 l=6
+ ad=0 pd=0 as=0 ps=0 
M2716 Vdd Vdd Vdd GND efet w=1 l=3
+ ad=0 pd=0 as=0 ps=0 
M2717 diff_1741_1957# Vdd Vdd GND efet w=16 l=124
+ ad=0 pd=0 as=0 ps=0 
M2718 diff_1751_1699# diff_847_938# GND GND efet w=28 l=16
+ ad=0 pd=0 as=0 ps=0 
M2719 diff_1751_1699# diff_1751_1699# diff_1751_1699# GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M2720 diff_1751_1699# diff_1751_1699# diff_1751_1699# GND efet w=1 l=2
+ ad=0 pd=0 as=0 ps=0 
M2721 diff_2261_1924# Vdd Vdd GND efet w=16 l=127
+ ad=3392 pd=438 as=0 ps=0 
M2722 GND d3 diff_2261_1924# GND efet w=70 l=14
+ ad=0 pd=0 as=0 ps=0 
M2723 diff_2521_1937# diff_2512_1924# diff_2521_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2724 diff_2563_2125# diff_2512_1924# diff_2572_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2725 diff_2623_1937# diff_2512_1924# diff_2623_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2726 diff_2674_1937# diff_2512_1924# diff_2674_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2727 diff_2725_1937# diff_2512_1924# diff_2725_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2728 diff_2776_1937# diff_2512_1924# diff_2776_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2729 diff_2827_1937# diff_2512_1924# diff_2827_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2730 diff_2878_1937# diff_2512_1924# diff_2878_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2731 diff_2929_1937# diff_2512_1924# diff_2929_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2732 diff_2980_1937# diff_2512_1924# diff_2980_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2733 diff_3031_1937# diff_2512_1924# diff_3031_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2734 diff_3082_1937# diff_2512_1924# diff_3082_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2735 diff_3133_1937# diff_2512_1924# diff_3133_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2736 diff_3184_1937# diff_2512_1924# diff_3184_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2737 diff_3235_1937# diff_2512_1924# diff_3235_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2738 diff_3286_1937# diff_2512_1924# diff_3286_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2739 diff_3337_1937# diff_2512_1924# diff_3337_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2740 diff_3388_1937# diff_2512_1924# diff_3388_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2741 diff_3439_1937# diff_2512_1924# diff_3439_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2742 diff_3490_1937# diff_2512_1924# diff_3490_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2743 diff_3541_1937# diff_2512_1924# diff_3541_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2744 diff_3592_1937# diff_2512_1924# diff_3592_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2745 diff_3643_1937# diff_2512_1924# diff_3643_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2746 diff_3694_1937# diff_2512_1924# diff_3694_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2747 diff_3745_1937# diff_2512_1924# diff_3745_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2748 diff_3796_1937# diff_2512_1924# diff_3796_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2749 diff_3847_1937# diff_2512_1924# diff_3847_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2750 diff_3898_1937# diff_2512_1924# diff_3898_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2751 diff_3949_1937# diff_2512_1924# diff_3949_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2752 diff_4000_1937# diff_2512_1924# diff_4000_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2753 diff_4051_1937# diff_2512_1924# diff_4051_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2754 diff_4102_1937# diff_2512_1924# diff_4102_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2755 diff_4153_1937# diff_2512_1924# diff_4153_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2756 diff_4204_1937# diff_2512_1924# diff_4204_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2757 diff_4255_1937# diff_2512_1924# diff_4255_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2758 diff_4306_1937# diff_2512_1924# diff_4306_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2759 diff_4357_1937# diff_2512_1924# diff_4357_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2760 diff_4408_1937# diff_2512_1924# diff_4408_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2761 diff_4459_1937# diff_2512_1924# diff_4459_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2762 diff_4510_1937# diff_2512_1924# diff_4510_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2763 diff_4561_1937# diff_2512_1924# diff_4561_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2764 diff_4612_1937# diff_2512_1924# diff_4612_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2765 diff_4663_1937# diff_2512_1924# diff_4663_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2766 diff_4714_1937# diff_2512_1924# diff_4714_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2767 diff_4765_1937# diff_2512_1924# diff_4765_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2768 diff_4816_1937# diff_2512_1924# diff_4816_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2769 diff_4867_1937# diff_2512_1924# diff_4867_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2770 diff_4918_1937# diff_2512_1924# diff_4918_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2771 diff_4969_1937# diff_2512_1924# diff_4969_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2772 diff_5020_1937# diff_2512_1924# diff_5020_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2773 diff_5071_1937# diff_2512_1924# diff_5071_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2774 diff_5122_1937# diff_2512_1924# diff_5122_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2775 diff_5173_1937# diff_2512_1924# diff_5173_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2776 diff_5224_1937# diff_2512_1924# diff_5224_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2777 diff_5275_1937# diff_2512_1924# diff_5275_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2778 diff_5326_1937# diff_2512_1924# diff_5326_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2779 diff_5377_1937# diff_2512_1924# diff_5377_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2780 diff_5428_1937# diff_2512_1924# diff_5428_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2781 diff_5479_1937# diff_2512_1924# diff_5479_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2782 diff_5530_1937# diff_2512_1924# diff_5530_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2783 diff_5581_1937# diff_2512_1924# diff_5581_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2784 diff_5632_1937# diff_2512_1924# diff_5632_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2785 diff_5683_1937# diff_2512_1924# diff_5683_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2786 diff_5734_1937# diff_2512_1924# diff_5734_1880# GND efet w=25 l=16
+ ad=657 pd=104 as=1025 ps=132 
M2787 GND diff_6316_3109# diff_6079_2449# GND efet w=304 l=13
+ ad=0 pd=0 as=10427 ps=828 
M2788 Vdd Vdd diff_2812_2884# GND efet w=16 l=34
+ ad=0 pd=0 as=0 ps=0 
M2789 Vdd Vdd diff_6079_2449# GND efet w=16 l=34
+ ad=0 pd=0 as=0 ps=0 
M2790 diff_6845_3073# diff_6808_2113# diff_6328_3004# GND efet w=46 l=13
+ ad=3632 pd=344 as=1638 ps=164 
M2791 Vdd Vdd diff_2812_2410# GND efet w=16 l=34
+ ad=0 pd=0 as=10937 ps=804 
M2792 diff_2812_2410# diff_6328_3004# GND GND efet w=304 l=13
+ ad=0 pd=0 as=0 ps=0 
M2793 GND diff_6328_2947# diff_5905_1069# GND efet w=304 l=13
+ ad=0 pd=0 as=12326 ps=828 
M2794 Vdd Vdd diff_5905_1069# GND efet w=16 l=34
+ ad=0 pd=0 as=0 ps=0 
M2795 Vdd Vdd diff_5962_1069# GND efet w=16 l=34
+ ad=0 pd=0 as=12266 ps=816 
M2796 diff_6935_3271# Vdd Vdd GND efet w=19 l=82
+ ad=0 pd=0 as=0 ps=0 
M2797 diff_7046_3232# diff_7033_2836# diff_6935_3271# GND efet w=88 l=13
+ ad=2288 pd=228 as=0 ps=0 
M2798 GND diff_7072_3184# diff_7046_3232# GND efet w=88 l=13
+ ad=0 pd=0 as=0 ps=0 
M2799 Vdd Vdd Vdd GND efet w=2 l=3
+ ad=0 pd=0 as=0 ps=0 
M2800 Vdd Vdd Vdd GND efet w=2 l=3
+ ad=0 pd=0 as=0 ps=0 
M2801 Vdd Vdd diff_6935_2974# GND efet w=19 l=82
+ ad=0 pd=0 as=7172 ps=524 
M2802 diff_6845_3073# diff_6778_3391# diff_6328_2947# GND efet w=52 l=13
+ ad=0 pd=0 as=2010 ps=182 
M2803 diff_6935_2974# clk2 diff_6845_3073# GND efet w=52 l=13
+ ad=0 pd=0 as=0 ps=0 
M2804 diff_7103_3070# diff_7072_3184# diff_6935_2974# GND efet w=85 l=13
+ ad=2210 pd=222 as=0 ps=0 
M2805 GND diff_7033_2509# diff_7103_3070# GND efet w=85 l=13
+ ad=0 pd=0 as=0 ps=0 
M2806 GND diff_7072_2716# diff_7046_2842# GND efet w=88 l=13
+ ad=0 pd=0 as=6036 ps=490 
M2807 diff_6845_2788# diff_6778_3391# diff_6328_2833# GND efet w=46 l=13
+ ad=3485 pd=338 as=1638 ps=164 
M2808 diff_6935_2884# clk2 diff_6845_2788# GND efet w=46 l=13
+ ad=5518 pd=388 as=0 ps=0 
M2809 diff_5962_1069# diff_6328_2833# GND GND efet w=304 l=13
+ ad=0 pd=0 as=0 ps=0 
M2810 GND diff_6331_2779# diff_2530_2884# GND efet w=304 l=13
+ ad=0 pd=0 as=11588 ps=810 
M2811 diff_6845_2788# diff_6808_2113# diff_6331_2779# GND efet w=49 l=13
+ ad=0 pd=0 as=1746 ps=170 
M2812 Vdd Vdd diff_2530_2884# GND efet w=16 l=34
+ ad=0 pd=0 as=0 ps=0 
M2813 diff_6845_2695# diff_6808_2113# diff_6328_2647# GND efet w=46 l=13
+ ad=3386 pd=332 as=1638 ps=164 
M2814 Vdd Vdd diff_2536_2407# GND efet w=16 l=34
+ ad=0 pd=0 as=11768 ps=810 
M2815 diff_2536_2407# diff_6328_2647# GND GND efet w=304 l=13
+ ad=0 pd=0 as=0 ps=0 
M2816 GND diff_6328_2590# diff_6034_2491# GND efet w=304 l=13
+ ad=0 pd=0 as=11975 ps=810 
M2817 Vdd Vdd diff_6034_2491# GND efet w=16 l=34
+ ad=0 pd=0 as=0 ps=0 
M2818 Vdd Vdd diff_6175_2281# GND efet w=16 l=34
+ ad=0 pd=0 as=12023 ps=816 
M2819 diff_6175_2281# diff_6328_2479# GND GND efet w=304 l=13
+ ad=0 pd=0 as=0 ps=0 
M2820 GND diff_6328_2422# diff_2584_2299# GND efet w=304 l=13
+ ad=0 pd=0 as=11396 ps=816 
M2821 diff_6935_2884# Vdd Vdd GND efet w=16 l=82
+ ad=0 pd=0 as=0 ps=0 
M2822 diff_7046_2842# diff_7033_2836# diff_6935_2884# GND efet w=88 l=13
+ ad=0 pd=0 as=0 ps=0 
M2823 diff_7163_2812# diff_7033_2509# diff_6935_2602# GND efet w=91 l=13
+ ad=2639 pd=240 as=7190 ps=536 
M2824 GND diff_7072_2716# diff_7163_2812# GND efet w=91 l=13
+ ad=0 pd=0 as=0 ps=0 
M2825 Vdd Vdd Vdd GND efet w=3 l=7
+ ad=0 pd=0 as=0 ps=0 
M2826 Vdd Vdd Vdd GND efet w=3 l=7
+ ad=0 pd=0 as=0 ps=0 
M2827 Vdd Vdd diff_6935_2602# GND efet w=16 l=82
+ ad=0 pd=0 as=0 ps=0 
M2828 diff_6845_2695# diff_6778_3391# diff_6328_2590# GND efet w=46 l=13
+ ad=0 pd=0 as=1638 ps=164 
M2829 diff_6935_2602# clk2 diff_6845_2695# GND efet w=46 l=13
+ ad=0 pd=0 as=0 ps=0 
M2830 diff_6845_2413# diff_6778_3391# diff_6328_2479# GND efet w=49 l=13
+ ad=3608 pd=344 as=1746 ps=170 
M2831 diff_6935_2506# clk2 diff_6845_2413# GND efet w=49 l=13
+ ad=7211 pd=536 as=0 ps=0 
M2832 d1 GND d1 GND efet w=445 l=274
+ ad=0 pd=0 as=0 ps=0 
M2833 GND diff_7072_2716# diff_7081_2687# GND efet w=157 l=13
+ ad=0 pd=0 as=4082 ps=366 
M2834 diff_7081_2687# diff_7033_2509# diff_7081_2641# GND efet w=157 l=13
+ ad=0 pd=0 as=11895 ps=868 
M2835 diff_2299_1054# diff_7033_2509# diff_7123_2480# GND efet w=115 l=13
+ ad=16636 pd=1484 as=2990 ps=282 
M2836 diff_6845_2413# diff_6808_2113# diff_6328_2422# GND efet w=49 l=13
+ ad=0 pd=0 as=1746 ps=170 
M2837 Vdd Vdd diff_2584_2299# GND efet w=13 l=34
+ ad=0 pd=0 as=0 ps=0 
M2838 Vdd Vdd diff_2659_2353# GND efet w=13 l=34
+ ad=0 pd=0 as=10847 ps=810 
M2839 diff_6845_2317# diff_6808_2113# diff_6325_2290# GND efet w=52 l=13
+ ad=3707 pd=350 as=1854 ps=176 
M2840 diff_2659_2353# diff_6325_2290# GND GND efet w=301 l=13
+ ad=0 pd=0 as=0 ps=0 
M2841 GND diff_6325_2236# diff_6130_2449# GND efet w=301 l=13
+ ad=0 pd=0 as=12101 ps=810 
M2842 Vdd Vdd diff_6130_2449# GND efet w=19 l=34
+ ad=0 pd=0 as=0 ps=0 
M2843 Vdd Vdd Vdd GND efet w=13 l=11
+ ad=0 pd=0 as=0 ps=0 
M2844 diff_2521_1880# diff_2512_1867# diff_2521_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2845 diff_2572_1880# diff_2512_1867# diff_2572_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2846 diff_2623_1880# diff_2512_1867# diff_2623_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2847 diff_2674_1880# diff_2512_1867# diff_2674_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2848 diff_2725_1880# diff_2512_1867# diff_2725_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2849 diff_2776_1880# diff_2512_1867# diff_2776_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2850 diff_2827_1880# diff_2512_1867# diff_2827_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2851 diff_2878_1880# diff_2512_1867# diff_2878_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2852 diff_2929_1880# diff_2512_1867# diff_2929_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2853 diff_2980_1880# diff_2512_1867# diff_2980_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2854 diff_3031_1880# diff_2512_1867# diff_3031_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2855 diff_3082_1880# diff_2512_1867# diff_3082_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2856 diff_3133_1880# diff_2512_1867# diff_3133_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2857 diff_3184_1880# diff_2512_1867# diff_3184_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2858 diff_3235_1880# diff_2512_1867# diff_3235_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2859 diff_3286_1880# diff_2512_1867# diff_3286_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2860 diff_3337_1880# diff_2512_1867# diff_3337_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2861 diff_3388_1880# diff_2512_1867# diff_3388_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2862 diff_3439_1880# diff_2512_1867# diff_3439_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2863 diff_3490_1880# diff_2512_1867# diff_3490_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2864 diff_3541_1880# diff_2512_1867# diff_3541_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2865 diff_3592_1880# diff_2512_1867# diff_3592_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2866 diff_3643_1880# diff_2512_1867# diff_3643_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2867 diff_3694_1880# diff_2512_1867# diff_3694_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2868 diff_3745_1880# diff_2512_1867# diff_3745_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2869 diff_3796_1880# diff_2512_1867# diff_3796_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2870 diff_3847_1880# diff_2512_1867# diff_3847_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2871 diff_3898_1880# diff_2512_1867# diff_3898_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2872 diff_3949_1880# diff_2512_1867# diff_3949_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2873 diff_4000_1880# diff_2512_1867# diff_4000_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2874 diff_4051_1880# diff_2512_1867# diff_4051_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2875 diff_4102_1880# diff_2512_1867# diff_4102_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2876 diff_4153_1880# diff_2512_1867# diff_4153_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2877 diff_4204_1880# diff_2512_1867# diff_4204_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2878 diff_4255_1880# diff_2512_1867# diff_4255_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2879 diff_4306_1880# diff_2512_1867# diff_4306_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2880 diff_4357_1880# diff_2512_1867# diff_4357_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2881 diff_4408_1880# diff_2512_1867# diff_4408_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2882 diff_4459_1880# diff_2512_1867# diff_4459_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2883 diff_4510_1880# diff_2512_1867# diff_4510_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2884 diff_4561_1880# diff_2512_1867# diff_4561_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2885 diff_4612_1880# diff_2512_1867# diff_4612_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2886 diff_4663_1880# diff_2512_1867# diff_4663_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2887 diff_4714_1880# diff_2512_1867# diff_4714_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2888 diff_4765_1880# diff_2512_1867# diff_4765_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2889 diff_4816_1880# diff_2512_1867# diff_4816_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2890 diff_4867_1880# diff_2512_1867# diff_4867_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2891 diff_4918_1880# diff_2512_1867# diff_4918_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2892 diff_4969_1880# diff_2512_1867# diff_4969_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2893 diff_5020_1880# diff_2512_1867# diff_5020_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2894 diff_5071_1880# diff_2512_1867# diff_5071_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2895 diff_5122_1880# diff_2512_1867# diff_5122_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2896 diff_5173_1880# diff_2512_1867# diff_5173_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2897 diff_5224_1880# diff_2512_1867# diff_5224_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2898 diff_5275_1880# diff_2512_1867# diff_5275_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2899 diff_5326_1880# diff_2512_1867# diff_5326_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2900 diff_5377_1880# diff_2512_1867# diff_5377_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2901 diff_5428_1880# diff_2512_1867# diff_5428_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2902 diff_5479_1880# diff_2512_1867# diff_5479_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2903 diff_5530_1880# diff_2512_1867# diff_5530_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2904 diff_5581_1880# diff_2512_1867# diff_5581_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2905 diff_5632_1880# diff_2512_1867# diff_5632_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2906 diff_5683_1880# diff_2512_1867# diff_5683_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2907 diff_5734_1880# diff_2512_1867# diff_5734_1826# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2908 diff_2512_1924# Vdd Vdd GND efet w=13 l=31
+ ad=5625 pd=646 as=0 ps=0 
M2909 Vdd Vdd Vdd GND efet w=5 l=12
+ ad=0 pd=0 as=0 ps=0 
M2910 Vdd Vdd Vdd GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M2911 diff_2165_1729# Vdd Vdd GND efet w=16 l=124
+ ad=3699 pd=368 as=0 ps=0 
M2912 diff_1030_2168# diff_2101_938# GND GND efet w=52 l=13
+ ad=0 pd=0 as=0 ps=0 
M2913 GND diff_2165_1729# diff_1030_2168# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2914 diff_2521_1826# diff_2512_1813# diff_2521_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2915 diff_2572_1826# diff_2512_1813# diff_2572_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2916 diff_2623_1826# diff_2512_1813# diff_2623_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2917 diff_2674_1826# diff_2512_1813# diff_2674_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2918 diff_2725_1826# diff_2512_1813# diff_2725_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2919 diff_2776_1826# diff_2512_1813# diff_2776_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2920 diff_2827_1826# diff_2512_1813# diff_2827_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2921 diff_2878_1826# diff_2512_1813# diff_2878_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2922 diff_2929_1826# diff_2512_1813# diff_2929_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2923 diff_2980_1826# diff_2512_1813# diff_2980_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2924 diff_3031_1826# diff_2512_1813# diff_3031_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2925 diff_3082_1826# diff_2512_1813# diff_3082_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2926 diff_3133_1826# diff_2512_1813# diff_3133_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2927 diff_3184_1826# diff_2512_1813# diff_3184_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2928 diff_3235_1826# diff_2512_1813# diff_3235_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2929 diff_3286_1826# diff_2512_1813# diff_3286_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2930 diff_3337_1826# diff_2512_1813# diff_3337_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2931 diff_3388_1826# diff_2512_1813# diff_3388_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2932 diff_3439_1826# diff_2512_1813# diff_3439_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2933 diff_3490_1826# diff_2512_1813# diff_3490_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2934 diff_3541_1826# diff_2512_1813# diff_3541_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2935 diff_3592_1826# diff_2512_1813# diff_3592_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2936 diff_3643_1826# diff_2512_1813# diff_3643_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2937 diff_3694_1826# diff_2512_1813# diff_3694_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2938 diff_3745_1826# diff_2512_1813# diff_3745_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2939 diff_3796_1826# diff_2512_1813# diff_3796_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2940 diff_3847_1826# diff_2512_1813# diff_3847_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2941 diff_3898_1826# diff_2512_1813# diff_3898_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2942 diff_3949_1826# diff_2512_1813# diff_3949_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2943 diff_4000_1826# diff_2512_1813# diff_4000_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2944 diff_4051_1826# diff_2512_1813# diff_4051_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2945 diff_4102_1826# diff_2512_1813# diff_4102_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2946 diff_4153_1826# diff_2512_1813# diff_4153_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2947 diff_4204_1826# diff_2512_1813# diff_4204_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2948 diff_4255_1826# diff_2512_1813# diff_4255_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2949 diff_4306_1826# diff_2512_1813# diff_4306_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2950 diff_4357_1826# diff_2512_1813# diff_4357_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2951 diff_4408_1826# diff_2512_1813# diff_4408_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2952 diff_4459_1826# diff_2512_1813# diff_4459_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2953 diff_4510_1826# diff_2512_1813# diff_4510_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2954 diff_4561_1826# diff_2512_1813# diff_4561_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2955 diff_4612_1826# diff_2512_1813# diff_4612_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2956 diff_4663_1826# diff_2512_1813# diff_4663_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2957 diff_4714_1826# diff_2512_1813# diff_4714_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2958 diff_4765_1826# diff_2512_1813# diff_4765_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2959 diff_4816_1826# diff_2512_1813# diff_4816_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2960 diff_4867_1826# diff_2512_1813# diff_4867_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2961 diff_4918_1826# diff_2512_1813# diff_4918_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2962 diff_4969_1826# diff_2512_1813# diff_4969_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2963 diff_5020_1826# diff_2512_1813# diff_5020_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2964 diff_5071_1826# diff_2512_1813# diff_5071_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2965 diff_5122_1826# diff_2512_1813# diff_5122_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2966 diff_5173_1826# diff_2512_1813# diff_5173_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2967 diff_5224_1826# diff_2512_1813# diff_5224_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2968 diff_5275_1826# diff_2512_1813# diff_5275_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2969 diff_5326_1826# diff_2512_1813# diff_5326_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2970 diff_5377_1826# diff_2512_1813# diff_5377_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2971 diff_5428_1826# diff_2512_1813# diff_5428_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2972 diff_5479_1826# diff_2512_1813# diff_5479_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2973 diff_5530_1826# diff_2512_1813# diff_5530_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2974 diff_5581_1826# diff_2512_1813# diff_5581_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2975 diff_5632_1826# diff_2512_1813# diff_5632_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2976 diff_5683_1826# diff_2512_1813# diff_5683_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2977 diff_5734_1826# diff_2512_1813# diff_5734_1769# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M2978 Vdd Vdd diff_2512_1756# GND efet w=13 l=28
+ ad=0 pd=0 as=5342 ps=570 
M2979 diff_5918_1741# diff_5905_1069# diff_2512_1756# GND efet w=214 l=13
+ ad=23356 pd=1814 as=0 ps=0 
M2980 diff_2165_1729# diff_2165_1729# diff_2165_1729# GND efet w=3 l=4
+ ad=0 pd=0 as=0 ps=0 
M2981 diff_2165_1729# diff_2165_1729# diff_2165_1729# GND efet w=4 l=4
+ ad=0 pd=0 as=0 ps=0 
M2982 GND diff_2261_1642# diff_2165_1729# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M2983 diff_2521_1769# diff_2512_1756# diff_2521_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2984 diff_2572_1769# diff_2512_1756# diff_2572_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2985 diff_2623_1769# diff_2512_1756# diff_2623_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2986 diff_2674_1769# diff_2512_1756# diff_2674_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2987 diff_2725_1769# diff_2512_1756# diff_2725_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2988 diff_2776_1769# diff_2512_1756# diff_2776_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2989 diff_2827_1769# diff_2512_1756# diff_2827_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2990 diff_2878_1769# diff_2512_1756# diff_2878_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2991 diff_2929_1769# diff_2512_1756# diff_2929_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2992 diff_2980_1769# diff_2512_1756# diff_2980_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2993 diff_3031_1769# diff_2512_1756# diff_3031_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2994 diff_3082_1769# diff_2512_1756# diff_3082_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2995 diff_3133_1769# diff_2512_1756# diff_3133_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2996 diff_3184_1769# diff_2512_1756# diff_3184_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2997 diff_3235_1769# diff_2512_1756# diff_3235_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2998 diff_3286_1769# diff_2512_1756# diff_3286_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M2999 diff_3337_1769# diff_2512_1756# diff_3337_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3000 diff_3388_1769# diff_2512_1756# diff_3388_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3001 diff_3439_1769# diff_2512_1756# diff_3439_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3002 diff_3490_1769# diff_2512_1756# diff_3490_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3003 diff_3541_1769# diff_2512_1756# diff_3541_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3004 diff_3592_1769# diff_2512_1756# diff_3592_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3005 diff_3643_1769# diff_2512_1756# diff_3643_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3006 diff_3694_1769# diff_2512_1756# diff_3694_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3007 diff_3745_1769# diff_2512_1756# diff_3745_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3008 diff_3796_1769# diff_2512_1756# diff_3796_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3009 diff_3847_1769# diff_2512_1756# diff_3847_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3010 diff_3898_1769# diff_2512_1756# diff_3898_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3011 diff_3949_1769# diff_2512_1756# diff_3949_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3012 diff_4000_1769# diff_2512_1756# diff_4000_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3013 diff_4051_1769# diff_2512_1756# diff_4051_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3014 diff_4102_1769# diff_2512_1756# diff_4102_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3015 diff_4153_1769# diff_2512_1756# diff_4153_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3016 diff_4204_1769# diff_2512_1756# diff_4204_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3017 diff_4255_1769# diff_2512_1756# diff_4255_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3018 diff_4306_1769# diff_2512_1756# diff_4306_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3019 diff_4357_1769# diff_2512_1756# diff_4357_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3020 diff_4408_1769# diff_2512_1756# diff_4408_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3021 diff_4459_1769# diff_2512_1756# diff_4459_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3022 diff_4510_1769# diff_2512_1756# diff_4510_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3023 diff_4561_1769# diff_2512_1756# diff_4561_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3024 diff_4612_1769# diff_2512_1756# diff_4612_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3025 diff_4663_1769# diff_2512_1756# diff_4663_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3026 diff_4714_1769# diff_2512_1756# diff_4714_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3027 diff_4765_1769# diff_2512_1756# diff_4765_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3028 diff_4816_1769# diff_2512_1756# diff_4816_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3029 diff_4867_1769# diff_2512_1756# diff_4867_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3030 diff_4918_1769# diff_2512_1756# diff_4918_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3031 diff_4969_1769# diff_2512_1756# diff_4969_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3032 diff_5020_1769# diff_2512_1756# diff_5020_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3033 diff_5071_1769# diff_2512_1756# diff_5071_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3034 diff_5122_1769# diff_2512_1756# diff_5122_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3035 diff_5173_1769# diff_2512_1756# diff_5173_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3036 diff_5224_1769# diff_2512_1756# diff_5224_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3037 diff_5275_1769# diff_2512_1756# diff_5275_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3038 diff_5326_1769# diff_2512_1756# diff_5326_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3039 diff_5377_1769# diff_2512_1756# diff_5377_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3040 diff_5428_1769# diff_2512_1756# diff_5428_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3041 diff_5479_1769# diff_2512_1756# diff_5479_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3042 diff_5530_1769# diff_2512_1756# diff_5530_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3043 diff_5581_1769# diff_2512_1756# diff_5581_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3044 diff_5632_1769# diff_2512_1756# diff_5632_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3045 diff_5683_1769# diff_2512_1756# diff_5683_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3046 diff_5734_1769# diff_2512_1756# diff_5734_1715# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3047 diff_2512_1924# diff_5962_1069# diff_5918_1741# GND efet w=184 l=13
+ ad=0 pd=0 as=0 ps=0 
M3048 diff_2512_1867# Vdd Vdd GND efet w=16 l=31
+ ad=6288 pd=616 as=0 ps=0 
M3049 Vdd Vdd diff_2512_1813# GND efet w=16 l=25
+ ad=0 pd=0 as=6479 ps=564 
M3050 diff_5918_1741# diff_6034_2491# diff_2512_1813# GND efet w=211 l=13
+ ad=0 pd=0 as=0 ps=0 
M3051 diff_2521_1715# diff_2512_1702# diff_2521_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3052 diff_2572_1715# diff_2512_1702# diff_2572_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3053 diff_2623_1715# diff_2512_1702# diff_2623_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3054 diff_2674_1715# diff_2512_1702# diff_2674_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3055 diff_2725_1715# diff_2512_1702# diff_2725_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3056 diff_2776_1715# diff_2512_1702# diff_2776_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3057 diff_2827_1715# diff_2512_1702# diff_2827_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3058 diff_2878_1715# diff_2512_1702# diff_2878_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3059 diff_2929_1715# diff_2512_1702# diff_2929_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3060 diff_2980_1715# diff_2512_1702# diff_2980_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3061 diff_3031_1715# diff_2512_1702# diff_3031_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3062 diff_3082_1715# diff_2512_1702# diff_3082_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3063 diff_3133_1715# diff_2512_1702# diff_3133_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3064 diff_3184_1715# diff_2512_1702# diff_3184_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3065 diff_3235_1715# diff_2512_1702# diff_3235_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3066 diff_3286_1715# diff_2512_1702# diff_3286_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3067 diff_3337_1715# diff_2512_1702# diff_3337_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3068 diff_3388_1715# diff_2512_1702# diff_3388_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3069 diff_3439_1715# diff_2512_1702# diff_3439_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3070 diff_3490_1715# diff_2512_1702# diff_3490_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3071 diff_3541_1715# diff_2512_1702# diff_3541_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3072 diff_3592_1715# diff_2512_1702# diff_3592_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3073 diff_3643_1715# diff_2512_1702# diff_3643_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3074 diff_3694_1715# diff_2512_1702# diff_3694_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3075 diff_3745_1715# diff_2512_1702# diff_3745_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3076 diff_3796_1715# diff_2512_1702# diff_3796_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3077 diff_3847_1715# diff_2512_1702# diff_3847_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3078 diff_3898_1715# diff_2512_1702# diff_3898_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3079 diff_3949_1715# diff_2512_1702# diff_3949_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3080 diff_4000_1715# diff_2512_1702# diff_4000_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3081 diff_4051_1715# diff_2512_1702# diff_4051_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3082 diff_4102_1715# diff_2512_1702# diff_4102_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3083 diff_4153_1715# diff_2512_1702# diff_4153_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3084 diff_4204_1715# diff_2512_1702# diff_4204_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3085 diff_4255_1715# diff_2512_1702# diff_4255_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3086 diff_4306_1715# diff_2512_1702# diff_4306_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3087 diff_4357_1715# diff_2512_1702# diff_4357_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3088 diff_4408_1715# diff_2512_1702# diff_4408_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3089 diff_4459_1715# diff_2512_1702# diff_4459_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3090 diff_4510_1715# diff_2512_1702# diff_4510_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3091 diff_4561_1715# diff_2512_1702# diff_4561_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3092 diff_4612_1715# diff_2512_1702# diff_4612_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3093 diff_4663_1715# diff_2512_1702# diff_4663_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3094 diff_4714_1715# diff_2512_1702# diff_4714_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3095 diff_4765_1715# diff_2512_1702# diff_4765_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3096 diff_4816_1715# diff_2512_1702# diff_4816_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3097 diff_4867_1715# diff_2512_1702# diff_4867_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3098 diff_4918_1715# diff_2512_1702# diff_4918_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3099 diff_4969_1715# diff_2512_1702# diff_4969_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3100 diff_5020_1715# diff_2512_1702# diff_5020_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3101 diff_5071_1715# diff_2512_1702# diff_5071_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3102 diff_5122_1715# diff_2512_1702# diff_5122_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3103 diff_5173_1715# diff_2512_1702# diff_5173_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3104 diff_5224_1715# diff_2512_1702# diff_5224_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3105 diff_5275_1715# diff_2512_1702# diff_5275_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3106 diff_5326_1715# diff_2512_1702# diff_5326_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3107 diff_5377_1715# diff_2512_1702# diff_5377_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3108 diff_5428_1715# diff_2512_1702# diff_5428_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3109 diff_5479_1715# diff_2512_1702# diff_5479_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3110 diff_5530_1715# diff_2512_1702# diff_5530_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3111 diff_5581_1715# diff_2512_1702# diff_5581_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3112 diff_5632_1715# diff_2512_1702# diff_5632_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3113 diff_5683_1715# diff_2512_1702# diff_5683_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3114 diff_5734_1715# diff_2512_1702# diff_5734_1658# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3115 diff_2512_1867# diff_6079_2449# diff_5918_1741# GND efet w=196 l=13
+ ad=0 pd=0 as=0 ps=0 
M3116 diff_5918_1519# diff_5905_1069# diff_2512_1534# GND efet w=218 l=16
+ ad=25921 pd=1796 as=5198 ps=570 
M3117 diff_2228_1642# clk2 Vdd GND efet w=28 l=16
+ ad=476 pd=90 as=0 ps=0 
M3118 diff_2261_1642# diff_2245_1597# diff_2228_1642# GND efet w=28 l=16
+ ad=2744 pd=252 as=0 ps=0 
M3119 GND diff_847_938# diff_2261_1642# GND efet w=28 l=16
+ ad=0 pd=0 as=0 ps=0 
M3120 diff_2521_1658# diff_2512_1645# diff_2521_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3121 diff_2572_1658# diff_2512_1645# diff_2572_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3122 diff_2623_1658# diff_2512_1645# diff_2623_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3123 diff_2674_1658# diff_2512_1645# diff_2674_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3124 diff_2725_1658# diff_2512_1645# diff_2725_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3125 diff_2776_1658# diff_2512_1645# diff_2776_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3126 diff_2827_1658# diff_2512_1645# diff_2827_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3127 diff_2878_1658# diff_2512_1645# diff_2878_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3128 diff_2929_1658# diff_2512_1645# diff_2929_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3129 diff_2980_1658# diff_2512_1645# diff_2980_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3130 diff_3031_1658# diff_2512_1645# diff_3031_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3131 diff_3082_1658# diff_2512_1645# diff_3082_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3132 diff_3133_1658# diff_2512_1645# diff_3133_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3133 diff_3184_1658# diff_2512_1645# diff_3184_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3134 diff_3235_1658# diff_2512_1645# diff_3235_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3135 diff_3286_1658# diff_2512_1645# diff_3286_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3136 diff_3337_1658# diff_2512_1645# diff_3337_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3137 diff_3388_1658# diff_2512_1645# diff_3388_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3138 diff_3439_1658# diff_2512_1645# diff_3439_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3139 diff_3490_1658# diff_2512_1645# diff_3490_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3140 diff_3541_1658# diff_2512_1645# diff_3541_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3141 diff_3592_1658# diff_2512_1645# diff_3592_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3142 diff_3643_1658# diff_2512_1645# diff_3643_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3143 diff_3694_1658# diff_2512_1645# diff_3694_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3144 diff_3745_1658# diff_2512_1645# diff_3745_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3145 diff_3796_1658# diff_2512_1645# diff_3796_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3146 diff_3847_1658# diff_2512_1645# diff_3847_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3147 diff_3898_1658# diff_2512_1645# diff_3898_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3148 diff_3949_1658# diff_2512_1645# diff_3949_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3149 diff_4000_1658# diff_2512_1645# diff_4000_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3150 diff_4051_1658# diff_2512_1645# diff_4051_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3151 diff_4102_1658# diff_2512_1645# diff_4102_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3152 diff_4153_1658# diff_2512_1645# diff_4153_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3153 diff_4204_1658# diff_2512_1645# diff_4204_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3154 diff_4255_1658# diff_2512_1645# diff_4255_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3155 diff_4306_1658# diff_2512_1645# diff_4306_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3156 diff_4357_1658# diff_2512_1645# diff_4357_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3157 diff_4408_1658# diff_2512_1645# diff_4408_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3158 diff_4459_1658# diff_2512_1645# diff_4459_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3159 diff_4510_1658# diff_2512_1645# diff_4510_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3160 diff_4561_1658# diff_2512_1645# diff_4561_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3161 diff_4612_1658# diff_2512_1645# diff_4612_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3162 diff_4663_1658# diff_2512_1645# diff_4663_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3163 diff_4714_1658# diff_2512_1645# diff_4714_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3164 diff_4765_1658# diff_2512_1645# diff_4765_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3165 diff_4816_1658# diff_2512_1645# diff_4816_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3166 diff_4867_1658# diff_2512_1645# diff_4867_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3167 diff_4918_1658# diff_2512_1645# diff_4918_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3168 diff_4969_1658# diff_2512_1645# diff_4969_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3169 diff_5020_1658# diff_2512_1645# diff_5020_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3170 diff_5071_1658# diff_2512_1645# diff_5071_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3171 diff_5122_1658# diff_2512_1645# diff_5122_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3172 diff_5173_1658# diff_2512_1645# diff_5173_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3173 diff_5224_1658# diff_2512_1645# diff_5224_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3174 diff_5275_1658# diff_2512_1645# diff_5275_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3175 diff_5326_1658# diff_2512_1645# diff_5326_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3176 diff_5377_1658# diff_2512_1645# diff_5377_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3177 diff_5428_1658# diff_2512_1645# diff_5428_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3178 diff_5479_1658# diff_2512_1645# diff_5479_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3179 diff_5530_1658# diff_2512_1645# diff_5530_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3180 diff_5581_1658# diff_2512_1645# diff_5581_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3181 diff_5632_1658# diff_2512_1645# diff_5632_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3182 diff_5683_1658# diff_2512_1645# diff_5683_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3183 diff_5734_1658# diff_2512_1645# diff_5734_1604# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3184 diff_2512_1702# Vdd Vdd GND efet w=13 l=31
+ ad=5625 pd=646 as=0 ps=0 
M3185 diff_1738_1906# diff_1867_1564# GND GND efet w=28 l=16
+ ad=1466 pd=174 as=0 ps=0 
M3186 Vdd Vdd diff_1738_1906# GND efet w=17 l=125
+ ad=0 pd=0 as=0 ps=0 
M3187 diff_1411_1187# diff_1411_1187# diff_1411_1187# GND efet w=5 l=7
+ ad=6736 pd=626 as=0 ps=0 
M3188 diff_1411_1187# diff_1411_1187# diff_1411_1187# GND efet w=5 l=8
+ ad=0 pd=0 as=0 ps=0 
M3189 Vdd Vdd diff_1411_1187# GND efet w=22 l=40
+ ad=0 pd=0 as=0 ps=0 
M3190 diff_2521_1604# diff_2512_1591# diff_2521_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3191 diff_2572_1604# diff_2512_1591# diff_2572_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3192 diff_2623_1604# diff_2512_1591# diff_2623_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3193 diff_2674_1604# diff_2512_1591# diff_2674_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3194 diff_2725_1604# diff_2512_1591# diff_2725_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3195 diff_2776_1604# diff_2512_1591# diff_2776_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3196 diff_2827_1604# diff_2512_1591# diff_2827_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3197 diff_2878_1604# diff_2512_1591# diff_2878_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3198 diff_2929_1604# diff_2512_1591# diff_2929_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3199 diff_2980_1604# diff_2512_1591# diff_2980_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3200 diff_3031_1604# diff_2512_1591# diff_3031_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3201 diff_3082_1604# diff_2512_1591# diff_3082_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3202 diff_3133_1604# diff_2512_1591# diff_3133_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3203 diff_3184_1604# diff_2512_1591# diff_3184_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3204 diff_3235_1604# diff_2512_1591# diff_3235_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3205 diff_3286_1604# diff_2512_1591# diff_3286_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3206 diff_3337_1604# diff_2512_1591# diff_3337_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3207 diff_3388_1604# diff_2512_1591# diff_3388_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3208 diff_3439_1604# diff_2512_1591# diff_3439_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3209 diff_3490_1604# diff_2512_1591# diff_3490_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3210 diff_3541_1604# diff_2512_1591# diff_3541_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3211 diff_3592_1604# diff_2512_1591# diff_3592_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3212 diff_3643_1604# diff_2512_1591# diff_3643_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3213 diff_3694_1604# diff_2512_1591# diff_3694_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3214 diff_3745_1604# diff_2512_1591# diff_3745_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3215 diff_3796_1604# diff_2512_1591# diff_3796_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3216 diff_3847_1604# diff_2512_1591# diff_3847_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3217 diff_3898_1604# diff_2512_1591# diff_3898_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3218 diff_3949_1604# diff_2512_1591# diff_3949_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3219 diff_4000_1604# diff_2512_1591# diff_4000_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3220 diff_4051_1604# diff_2512_1591# diff_4051_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3221 diff_4102_1604# diff_2512_1591# diff_4102_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3222 diff_4153_1604# diff_2512_1591# diff_4153_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3223 diff_4204_1604# diff_2512_1591# diff_4204_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3224 diff_4255_1604# diff_2512_1591# diff_4255_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3225 diff_4306_1604# diff_2512_1591# diff_4306_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3226 diff_4357_1604# diff_2512_1591# diff_4357_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3227 diff_4408_1604# diff_2512_1591# diff_4408_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3228 diff_4459_1604# diff_2512_1591# diff_4459_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3229 diff_4510_1604# diff_2512_1591# diff_4510_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3230 diff_4561_1604# diff_2512_1591# diff_4561_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3231 diff_4612_1604# diff_2512_1591# diff_4612_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3232 diff_4663_1604# diff_2512_1591# diff_4663_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3233 diff_4714_1604# diff_2512_1591# diff_4714_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3234 diff_4765_1604# diff_2512_1591# diff_4765_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3235 diff_4816_1604# diff_2512_1591# diff_4816_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3236 diff_4867_1604# diff_2512_1591# diff_4867_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3237 diff_4918_1604# diff_2512_1591# diff_4918_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3238 diff_4969_1604# diff_2512_1591# diff_4969_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3239 diff_5020_1604# diff_2512_1591# diff_5020_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3240 diff_5071_1604# diff_2512_1591# diff_5071_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3241 diff_5122_1604# diff_2512_1591# diff_5122_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3242 diff_5173_1604# diff_2512_1591# diff_5173_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3243 diff_5224_1604# diff_2512_1591# diff_5224_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3244 diff_5275_1604# diff_2512_1591# diff_5275_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3245 diff_5326_1604# diff_2512_1591# diff_5326_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3246 diff_5377_1604# diff_2512_1591# diff_5377_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3247 diff_5428_1604# diff_2512_1591# diff_5428_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3248 diff_5479_1604# diff_2512_1591# diff_5479_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3249 diff_5530_1604# diff_2512_1591# diff_5530_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3250 diff_5581_1604# diff_2512_1591# diff_5581_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3251 diff_5632_1604# diff_2512_1591# diff_5632_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3252 diff_5683_1604# diff_2512_1591# diff_5683_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3253 diff_5734_1604# diff_2512_1591# diff_5734_1547# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3254 Vdd Vdd diff_2512_1534# GND efet w=13 l=28
+ ad=0 pd=0 as=0 ps=0 
M3255 Vdd Vdd diff_1561_1187# GND efet w=22 l=40
+ ad=0 pd=0 as=5121 ps=466 
M3256 Vdd Vdd Vdd GND efet w=8 l=8
+ ad=0 pd=0 as=0 ps=0 
M3257 Vdd Vdd diff_1738_1391# GND efet w=16 l=157
+ ad=0 pd=0 as=5285 ps=522 
M3258 diff_1738_1391# cm diff_1738_1232# GND efet w=193 l=16
+ ad=0 pd=0 as=4568 ps=432 
M3259 diff_1012_1177# diff_847_938# Vdd GND efet w=31 l=13
+ ad=1550 pd=162 as=0 ps=0 
M3260 diff_1187_1252# clk2 diff_1012_1177# GND efet w=31 l=16
+ ad=713 pd=108 as=0 ps=0 
M3261 diff_1226_1252# diff_1198_1177# diff_1187_1252# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M3262 Vdd Vdd diff_1729_1219# GND efet w=19 l=124
+ ad=0 pd=0 as=6029 ps=552 
M3263 Vdd Vdd diff_1891_1138# GND efet w=16 l=124
+ ad=0 pd=0 as=2808 ps=316 
M3264 Vdd Vdd Vdd GND efet w=8 l=8
+ ad=0 pd=0 as=0 ps=0 
M3265 diff_2245_1597# Vdd Vdd GND efet w=16 l=85
+ ad=3895 pd=408 as=0 ps=0 
M3266 GND diff_1738_1391# diff_2245_1597# GND efet w=43 l=16
+ ad=0 pd=0 as=0 ps=0 
M3267 diff_2245_1597# diff_2261_1924# GND GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M3268 GND diff_2299_1054# diff_2245_1597# GND efet w=43 l=16
+ ad=0 pd=0 as=0 ps=0 
M3269 diff_2521_1547# diff_2512_1534# diff_2521_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3270 diff_2572_1547# diff_2512_1534# diff_2572_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3271 diff_2623_1547# diff_2512_1534# diff_2623_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3272 diff_2674_1547# diff_2512_1534# diff_2674_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3273 diff_2725_1547# diff_2512_1534# diff_2725_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3274 diff_2776_1547# diff_2512_1534# diff_2776_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3275 diff_2827_1547# diff_2512_1534# diff_2827_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3276 diff_2878_1547# diff_2512_1534# diff_2878_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3277 diff_2929_1547# diff_2512_1534# diff_2929_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3278 diff_2980_1547# diff_2512_1534# diff_2980_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3279 diff_3031_1547# diff_2512_1534# diff_3031_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3280 diff_3082_1547# diff_2512_1534# diff_3082_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3281 diff_3133_1547# diff_2512_1534# diff_3133_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3282 diff_3184_1547# diff_2512_1534# diff_3184_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3283 diff_3235_1547# diff_2512_1534# diff_3235_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3284 diff_3286_1547# diff_2512_1534# diff_3286_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3285 diff_3337_1547# diff_2512_1534# diff_3337_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3286 diff_3388_1547# diff_2512_1534# diff_3388_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3287 diff_3439_1547# diff_2512_1534# diff_3439_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3288 diff_3490_1547# diff_2512_1534# diff_3490_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3289 diff_3541_1547# diff_2512_1534# diff_3541_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3290 diff_3592_1547# diff_2512_1534# diff_3592_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3291 diff_3643_1547# diff_2512_1534# diff_3643_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3292 diff_3694_1547# diff_2512_1534# diff_3694_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3293 diff_3745_1547# diff_2512_1534# diff_3745_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3294 diff_3796_1547# diff_2512_1534# diff_3796_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3295 diff_3847_1547# diff_2512_1534# diff_3847_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3296 diff_3898_1547# diff_2512_1534# diff_3898_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3297 diff_3949_1547# diff_2512_1534# diff_3949_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3298 diff_4000_1547# diff_2512_1534# diff_4000_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3299 diff_4051_1547# diff_2512_1534# diff_4051_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3300 diff_4102_1547# diff_2512_1534# diff_4102_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3301 diff_4153_1547# diff_2512_1534# diff_4153_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3302 diff_4204_1547# diff_2512_1534# diff_4204_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3303 diff_4255_1547# diff_2512_1534# diff_4255_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3304 diff_4306_1547# diff_2512_1534# diff_4306_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3305 diff_4357_1547# diff_2512_1534# diff_4357_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3306 diff_4408_1547# diff_2512_1534# diff_4408_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3307 diff_4459_1547# diff_2512_1534# diff_4459_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3308 diff_4510_1547# diff_2512_1534# diff_4510_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3309 diff_4561_1547# diff_2512_1534# diff_4561_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3310 diff_4612_1547# diff_2512_1534# diff_4612_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3311 diff_4663_1547# diff_2512_1534# diff_4663_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3312 diff_4714_1547# diff_2512_1534# diff_4714_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3313 diff_4765_1547# diff_2512_1534# diff_4765_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3314 diff_4816_1547# diff_2512_1534# diff_4816_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3315 diff_4867_1547# diff_2512_1534# diff_4867_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3316 diff_4918_1547# diff_2512_1534# diff_4918_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3317 diff_4969_1547# diff_2512_1534# diff_4969_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3318 diff_5020_1547# diff_2512_1534# diff_5020_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3319 diff_5071_1547# diff_2512_1534# diff_5071_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3320 diff_5122_1547# diff_2512_1534# diff_5122_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3321 diff_5173_1547# diff_2512_1534# diff_5173_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3322 diff_5224_1547# diff_2512_1534# diff_5224_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3323 diff_5275_1547# diff_2512_1534# diff_5275_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3324 diff_5326_1547# diff_2512_1534# diff_5326_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3325 diff_5377_1547# diff_2512_1534# diff_5377_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3326 diff_5428_1547# diff_2512_1534# diff_5428_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3327 diff_5479_1547# diff_2512_1534# diff_5479_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3328 diff_5530_1547# diff_2512_1534# diff_5530_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3329 diff_5581_1547# diff_2512_1534# diff_5581_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3330 diff_5632_1547# diff_2512_1534# diff_5632_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3331 diff_5683_1547# diff_2512_1534# diff_5683_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3332 diff_5734_1547# diff_2512_1534# diff_5734_1493# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3333 Vdd Vdd diff_2026_1276# GND efet w=16 l=127
+ ad=0 pd=0 as=3683 ps=432 
M3334 diff_2512_1702# diff_5962_1069# diff_5918_1519# GND efet w=184 l=13
+ ad=0 pd=0 as=0 ps=0 
M3335 diff_2512_1645# Vdd Vdd GND efet w=16 l=28
+ ad=6288 pd=616 as=0 ps=0 
M3336 Vdd Vdd diff_2512_1591# GND efet w=16 l=25
+ ad=0 pd=0 as=6512 ps=564 
M3337 diff_5918_1519# diff_6034_2491# diff_2512_1591# GND efet w=208 l=13
+ ad=0 pd=0 as=0 ps=0 
M3338 diff_2521_1493# diff_2512_1480# diff_2521_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3339 diff_2572_1493# diff_2512_1480# diff_2572_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3340 diff_2623_1493# diff_2512_1480# diff_2623_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3341 diff_2674_1493# diff_2512_1480# diff_2674_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3342 diff_2725_1493# diff_2512_1480# diff_2725_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3343 diff_2776_1493# diff_2512_1480# diff_2776_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3344 diff_2827_1493# diff_2512_1480# diff_2827_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3345 diff_2878_1493# diff_2512_1480# diff_2878_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3346 diff_2929_1493# diff_2512_1480# diff_2929_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3347 diff_2980_1493# diff_2512_1480# diff_2980_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3348 diff_3031_1493# diff_2512_1480# diff_3031_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3349 diff_3082_1493# diff_2512_1480# diff_3082_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3350 diff_3133_1493# diff_2512_1480# diff_3133_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3351 diff_3184_1493# diff_2512_1480# diff_3184_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3352 diff_3235_1493# diff_2512_1480# diff_3235_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3353 diff_3286_1493# diff_2512_1480# diff_3286_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3354 diff_3337_1493# diff_2512_1480# diff_3337_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3355 diff_3388_1493# diff_2512_1480# diff_3388_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3356 diff_3439_1493# diff_2512_1480# diff_3439_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3357 diff_3490_1493# diff_2512_1480# diff_3490_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3358 diff_3541_1493# diff_2512_1480# diff_3541_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3359 diff_3592_1493# diff_2512_1480# diff_3592_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3360 diff_3643_1493# diff_2512_1480# diff_3643_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3361 diff_3694_1493# diff_2512_1480# diff_3694_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3362 diff_3745_1493# diff_2512_1480# diff_3745_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3363 diff_3796_1493# diff_2512_1480# diff_3796_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3364 diff_3847_1493# diff_2512_1480# diff_3847_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3365 diff_3898_1493# diff_2512_1480# diff_3898_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3366 diff_3949_1493# diff_2512_1480# diff_3949_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3367 diff_4000_1493# diff_2512_1480# diff_4000_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3368 diff_4051_1493# diff_2512_1480# diff_4051_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3369 diff_4102_1493# diff_2512_1480# diff_4102_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3370 diff_4153_1493# diff_2512_1480# diff_4153_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3371 diff_4204_1493# diff_2512_1480# diff_4204_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3372 diff_4255_1493# diff_2512_1480# diff_4255_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3373 diff_4306_1493# diff_2512_1480# diff_4306_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3374 diff_4357_1493# diff_2512_1480# diff_4357_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3375 diff_4408_1493# diff_2512_1480# diff_4408_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3376 diff_4459_1493# diff_2512_1480# diff_4459_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3377 diff_4510_1493# diff_2512_1480# diff_4510_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3378 diff_4561_1493# diff_2512_1480# diff_4561_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3379 diff_4612_1493# diff_2512_1480# diff_4612_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3380 diff_4663_1493# diff_2512_1480# diff_4663_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3381 diff_4714_1493# diff_2512_1480# diff_4714_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3382 diff_4765_1493# diff_2512_1480# diff_4765_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3383 diff_4816_1493# diff_2512_1480# diff_4816_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3384 diff_4867_1493# diff_2512_1480# diff_4867_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3385 diff_4918_1493# diff_2512_1480# diff_4918_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3386 diff_4969_1493# diff_2512_1480# diff_4969_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3387 diff_5020_1493# diff_2512_1480# diff_5020_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3388 diff_5071_1493# diff_2512_1480# diff_5071_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3389 diff_5122_1493# diff_2512_1480# diff_5122_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3390 diff_5173_1493# diff_2512_1480# diff_5173_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3391 diff_5224_1493# diff_2512_1480# diff_5224_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3392 diff_5275_1493# diff_2512_1480# diff_5275_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3393 diff_5326_1493# diff_2512_1480# diff_5326_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3394 diff_5377_1493# diff_2512_1480# diff_5377_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3395 diff_5428_1493# diff_2512_1480# diff_5428_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3396 diff_5479_1493# diff_2512_1480# diff_5479_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3397 diff_5530_1493# diff_2512_1480# diff_5530_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3398 diff_5581_1493# diff_2512_1480# diff_5581_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3399 diff_5632_1493# diff_2512_1480# diff_5632_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3400 diff_5683_1493# diff_2512_1480# diff_5683_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3401 diff_5734_1493# diff_2512_1480# diff_5734_1436# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3402 diff_2512_1645# diff_6079_2449# diff_5918_1519# GND efet w=196 l=13
+ ad=0 pd=0 as=0 ps=0 
M3403 diff_6269_1078# diff_6130_2449# diff_5918_1741# GND efet w=385 l=16
+ ad=46744 pd=2806 as=0 ps=0 
M3404 diff_5918_1519# diff_6175_2281# diff_6269_1078# GND efet w=385 l=16
+ ad=0 pd=0 as=0 ps=0 
M3405 diff_5918_1300# diff_5905_1069# diff_2512_1312# GND efet w=217 l=14
+ ad=23338 pd=1820 as=4874 ps=558 
M3406 diff_2521_1436# diff_2512_1423# diff_2521_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3407 diff_2572_1436# diff_2512_1423# diff_2572_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3408 diff_2623_1436# diff_2512_1423# diff_2623_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3409 diff_2674_1436# diff_2512_1423# diff_2674_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3410 diff_2725_1436# diff_2512_1423# diff_2725_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3411 diff_2776_1436# diff_2512_1423# diff_2776_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3412 diff_2827_1436# diff_2512_1423# diff_2827_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3413 diff_2878_1436# diff_2512_1423# diff_2878_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3414 diff_2929_1436# diff_2512_1423# diff_2929_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3415 diff_2980_1436# diff_2512_1423# diff_2980_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3416 diff_3031_1436# diff_2512_1423# diff_3031_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3417 diff_3082_1436# diff_2512_1423# diff_3082_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3418 diff_3133_1436# diff_2512_1423# diff_3133_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3419 diff_3184_1436# diff_2512_1423# diff_3184_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3420 diff_3235_1436# diff_2512_1423# diff_3235_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3421 diff_3286_1436# diff_2512_1423# diff_3286_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3422 diff_3337_1436# diff_2512_1423# diff_3337_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3423 diff_3388_1436# diff_2512_1423# diff_3388_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3424 diff_3439_1436# diff_2512_1423# diff_3439_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3425 diff_3490_1436# diff_2512_1423# diff_3490_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3426 diff_3541_1436# diff_2512_1423# diff_3541_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3427 diff_3592_1436# diff_2512_1423# diff_3592_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3428 diff_3643_1436# diff_2512_1423# diff_3643_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3429 diff_3694_1436# diff_2512_1423# diff_3694_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3430 diff_3745_1436# diff_2512_1423# diff_3745_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3431 diff_3796_1436# diff_2512_1423# diff_3796_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3432 diff_3847_1436# diff_2512_1423# diff_3847_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3433 diff_3898_1436# diff_2512_1423# diff_3898_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3434 diff_3949_1436# diff_2512_1423# diff_3949_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3435 diff_4000_1436# diff_2512_1423# diff_4000_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3436 diff_4051_1436# diff_2512_1423# diff_4051_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3437 diff_4102_1436# diff_2512_1423# diff_4102_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3438 diff_4153_1436# diff_2512_1423# diff_4153_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3439 diff_4204_1436# diff_2512_1423# diff_4204_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3440 diff_4255_1436# diff_2512_1423# diff_4255_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3441 diff_4306_1436# diff_2512_1423# diff_4306_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3442 diff_4357_1436# diff_2512_1423# diff_4357_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3443 diff_4408_1436# diff_2512_1423# diff_4408_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3444 diff_4459_1436# diff_2512_1423# diff_4459_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3445 diff_4510_1436# diff_2512_1423# diff_4510_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3446 diff_4561_1436# diff_2512_1423# diff_4561_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3447 diff_4612_1436# diff_2512_1423# diff_4612_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3448 diff_4663_1436# diff_2512_1423# diff_4663_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3449 diff_4714_1436# diff_2512_1423# diff_4714_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3450 diff_4765_1436# diff_2512_1423# diff_4765_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3451 diff_4816_1436# diff_2512_1423# diff_4816_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3452 diff_4867_1436# diff_2512_1423# diff_4867_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3453 diff_4918_1436# diff_2512_1423# diff_4918_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3454 diff_4969_1436# diff_2512_1423# diff_4969_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3455 diff_5020_1436# diff_2512_1423# diff_5020_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3456 diff_5071_1436# diff_2512_1423# diff_5071_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3457 diff_5122_1436# diff_2512_1423# diff_5122_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3458 diff_5173_1436# diff_2512_1423# diff_5173_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3459 diff_5224_1436# diff_2512_1423# diff_5224_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3460 diff_5275_1436# diff_2512_1423# diff_5275_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3461 diff_5326_1436# diff_2512_1423# diff_5326_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3462 diff_5377_1436# diff_2512_1423# diff_5377_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3463 diff_5428_1436# diff_2512_1423# diff_5428_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3464 diff_5479_1436# diff_2512_1423# diff_5479_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3465 diff_5530_1436# diff_2512_1423# diff_5530_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3466 diff_5581_1436# diff_2512_1423# diff_5581_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3467 diff_5632_1436# diff_2512_1423# diff_5632_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3468 diff_5683_1436# diff_2512_1423# diff_5683_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3469 diff_5734_1436# diff_2512_1423# diff_5734_1382# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3470 diff_2512_1480# Vdd Vdd GND efet w=13 l=31
+ ad=5625 pd=646 as=0 ps=0 
M3471 diff_1942_1222# Vdd Vdd GND efet w=17 l=215
+ ad=2172 pd=266 as=0 ps=0 
M3472 diff_2521_1382# diff_2512_1369# diff_2521_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3473 diff_2572_1382# diff_2512_1369# diff_2572_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3474 diff_2623_1382# diff_2512_1369# diff_2623_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3475 diff_2674_1382# diff_2512_1369# diff_2674_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3476 diff_2725_1382# diff_2512_1369# diff_2725_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3477 diff_2776_1382# diff_2512_1369# diff_2776_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3478 diff_2827_1382# diff_2512_1369# diff_2827_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3479 diff_2878_1382# diff_2512_1369# diff_2878_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3480 diff_2929_1382# diff_2512_1369# diff_2929_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3481 diff_2980_1382# diff_2512_1369# diff_2980_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3482 diff_3031_1382# diff_2512_1369# diff_3031_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3483 diff_3082_1382# diff_2512_1369# diff_3082_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3484 diff_3133_1382# diff_2512_1369# diff_3133_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3485 diff_3184_1382# diff_2512_1369# diff_3184_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3486 diff_3235_1382# diff_2512_1369# diff_3235_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3487 diff_3286_1382# diff_2512_1369# diff_3286_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3488 diff_3337_1382# diff_2512_1369# diff_3337_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3489 diff_3388_1382# diff_2512_1369# diff_3388_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3490 diff_3439_1382# diff_2512_1369# diff_3439_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3491 diff_3490_1382# diff_2512_1369# diff_3490_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3492 diff_3541_1382# diff_2512_1369# diff_3541_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3493 diff_3592_1382# diff_2512_1369# diff_3592_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3494 diff_3643_1382# diff_2512_1369# diff_3643_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3495 diff_3694_1382# diff_2512_1369# diff_3694_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3496 diff_3745_1382# diff_2512_1369# diff_3745_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3497 diff_3796_1382# diff_2512_1369# diff_3796_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3498 diff_3847_1382# diff_2512_1369# diff_3847_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3499 diff_3898_1382# diff_2512_1369# diff_3898_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3500 diff_3949_1382# diff_2512_1369# diff_3949_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3501 diff_4000_1382# diff_2512_1369# diff_4000_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3502 diff_4051_1382# diff_2512_1369# diff_4051_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3503 diff_4102_1382# diff_2512_1369# diff_4102_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3504 diff_4153_1382# diff_2512_1369# diff_4153_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3505 diff_4204_1382# diff_2512_1369# diff_4204_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3506 diff_4255_1382# diff_2512_1369# diff_4255_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3507 diff_4306_1382# diff_2512_1369# diff_4306_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3508 diff_4357_1382# diff_2512_1369# diff_4357_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3509 diff_4408_1382# diff_2512_1369# diff_4408_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3510 diff_4459_1382# diff_2512_1369# diff_4459_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3511 diff_4510_1382# diff_2512_1369# diff_4510_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3512 diff_4561_1382# diff_2512_1369# diff_4561_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3513 diff_4612_1382# diff_2512_1369# diff_4612_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3514 diff_4663_1382# diff_2512_1369# diff_4663_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3515 diff_4714_1382# diff_2512_1369# diff_4714_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3516 diff_4765_1382# diff_2512_1369# diff_4765_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3517 diff_4816_1382# diff_2512_1369# diff_4816_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3518 diff_4867_1382# diff_2512_1369# diff_4867_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3519 diff_4918_1382# diff_2512_1369# diff_4918_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3520 diff_4969_1382# diff_2512_1369# diff_4969_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3521 diff_5020_1382# diff_2512_1369# diff_5020_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3522 diff_5071_1382# diff_2512_1369# diff_5071_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3523 diff_5122_1382# diff_2512_1369# diff_5122_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3524 diff_5173_1382# diff_2512_1369# diff_5173_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3525 diff_5224_1382# diff_2512_1369# diff_5224_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3526 diff_5275_1382# diff_2512_1369# diff_5275_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3527 diff_5326_1382# diff_2512_1369# diff_5326_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3528 diff_5377_1382# diff_2512_1369# diff_5377_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3529 diff_5428_1382# diff_2512_1369# diff_5428_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3530 diff_5479_1382# diff_2512_1369# diff_5479_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3531 diff_5530_1382# diff_2512_1369# diff_5530_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3532 diff_5581_1382# diff_2512_1369# diff_5581_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3533 diff_5632_1382# diff_2512_1369# diff_5632_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3534 diff_5683_1382# diff_2512_1369# diff_5683_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3535 diff_5734_1382# diff_2512_1369# diff_5734_1325# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3536 diff_1024_1190# diff_1012_1177# GND GND efet w=79 l=16
+ ad=0 pd=0 as=0 ps=0 
M3537 diff_1226_1252# diff_1243_1231# diff_1252_1199# GND efet w=46 l=16
+ ad=0 pd=0 as=1973 ps=222 
M3538 diff_1951_1117# diff_1942_1222# diff_1729_1219# GND efet w=31 l=16
+ ad=5172 pd=488 as=0 ps=0 
M3539 diff_1243_1231# diff_2026_1276# diff_1951_1117# GND efet w=31 l=16
+ ad=6143 pd=596 as=0 ps=0 
M3540 diff_1252_1199# cm GND GND efet w=82 l=16
+ ad=0 pd=0 as=0 ps=0 
M3541 diff_1738_1232# diff_1729_1219# diff_1738_1196# GND efet w=73 l=16
+ ad=0 pd=0 as=1559 ps=210 
M3542 diff_1729_1219# diff_1729_1219# diff_1729_1219# GND efet w=1 l=1
+ ad=0 pd=0 as=0 ps=0 
M3543 diff_1729_1219# diff_1729_1219# diff_1729_1219# GND efet w=3 l=4
+ ad=0 pd=0 as=0 ps=0 
M3544 diff_1738_1196# diff_1729_1183# GND GND efet w=85 l=14
+ ad=0 pd=0 as=0 ps=0 
M3545 diff_1411_1187# diff_1378_1138# GND GND efet w=112 l=16
+ ad=0 pd=0 as=0 ps=0 
M3546 diff_1561_1187# diff_1555_1174# GND GND efet w=112 l=16
+ ad=0 pd=0 as=0 ps=0 
M3547 diff_847_938# diff_803_997# GND GND efet w=49 l=16
+ ad=5215 pd=514 as=0 ps=0 
M3548 diff_958_938# diff_917_997# GND GND efet w=46 l=16
+ ad=4384 pd=484 as=0 ps=0 
M3549 diff_1075_938# diff_1034_997# GND GND efet w=49 l=16
+ ad=4006 pd=472 as=0 ps=0 
M3550 diff_803_997# clk1 diff_724_1144# GND efet w=25 l=16
+ ad=844 pd=130 as=0 ps=0 
M3551 diff_803_997# diff_803_997# diff_803_997# GND efet w=2 l=10
+ ad=0 pd=0 as=0 ps=0 
M3552 diff_803_997# diff_803_997# diff_803_997# GND efet w=2 l=4
+ ad=0 pd=0 as=0 ps=0 
M3553 diff_917_997# clk2 diff_847_938# GND efet w=28 l=16
+ ad=889 pd=124 as=0 ps=0 
M3554 diff_917_997# diff_917_997# diff_917_997# GND efet w=2 l=4
+ ad=0 pd=0 as=0 ps=0 
M3555 diff_917_997# diff_917_997# diff_917_997# GND efet w=0 l=1
+ ad=0 pd=0 as=0 ps=0 
M3556 diff_1034_997# clk1 diff_958_938# GND efet w=28 l=16
+ ad=871 pd=130 as=0 ps=0 
M3557 diff_1034_997# diff_1034_997# diff_1034_997# GND efet w=5 l=8
+ ad=0 pd=0 as=0 ps=0 
M3558 GND diff_1891_1138# diff_1729_1219# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M3559 diff_1186_938# diff_1148_997# GND GND efet w=46 l=16
+ ad=4330 pd=484 as=0 ps=0 
M3560 diff_1198_1177# diff_1265_997# GND GND efet w=49 l=16
+ ad=5026 pd=532 as=0 ps=0 
M3561 diff_1378_1138# diff_1376_997# GND GND efet w=46 l=16
+ ad=5119 pd=532 as=0 ps=0 
M3562 diff_1534_938# diff_1493_997# GND GND efet w=49 l=16
+ ad=4006 pd=472 as=0 ps=0 
M3563 diff_1555_1174# diff_1607_997# GND GND efet w=46 l=16
+ ad=4993 pd=532 as=0 ps=0 
M3564 diff_1891_1138# diff_1951_1117# GND GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M3565 diff_1942_1222# diff_1942_1222# diff_1942_1222# GND efet w=0 l=1
+ ad=0 pd=0 as=0 ps=0 
M3566 diff_2026_1276# diff_1942_1222# GND GND efet w=28 l=16
+ ad=0 pd=0 as=0 ps=0 
M3567 diff_1942_1222# diff_1942_1222# diff_1942_1222# GND efet w=1 l=1
+ ad=0 pd=0 as=0 ps=0 
M3568 diff_1951_1117# diff_1951_1117# diff_1951_1117# GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M3569 diff_1951_1117# diff_1951_1117# diff_1951_1117# GND efet w=2 l=7
+ ad=0 pd=0 as=0 ps=0 
M3570 diff_2261_1162# clk2 diff_1942_1222# GND efet w=55 l=16
+ ad=1865 pd=198 as=0 ps=0 
M3571 diff_2306_1147# diff_1867_1564# diff_2261_1162# GND efet w=70 l=16
+ ad=5792 pd=498 as=0 ps=0 
M3572 Vdd Vdd diff_2512_1312# GND efet w=13 l=31
+ ad=0 pd=0 as=0 ps=0 
M3573 diff_2521_1325# diff_2512_1312# diff_2521_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3574 diff_2572_1325# diff_2512_1312# diff_2572_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3575 diff_2623_1325# diff_2512_1312# diff_2623_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3576 diff_2674_1325# diff_2512_1312# diff_2674_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3577 diff_2725_1325# diff_2512_1312# diff_2725_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3578 diff_2776_1325# diff_2512_1312# diff_2776_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3579 diff_2827_1325# diff_2512_1312# diff_2827_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3580 diff_2878_1325# diff_2512_1312# diff_2878_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3581 diff_2929_1325# diff_2512_1312# diff_2929_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3582 diff_2980_1325# diff_2512_1312# diff_2980_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3583 diff_3031_1325# diff_2512_1312# diff_3031_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3584 diff_3082_1325# diff_2512_1312# diff_3082_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3585 diff_3133_1325# diff_2512_1312# diff_3133_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3586 diff_3184_1325# diff_2512_1312# diff_3184_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3587 diff_3235_1325# diff_2512_1312# diff_3235_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3588 diff_3286_1325# diff_2512_1312# diff_3286_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3589 diff_3337_1325# diff_2512_1312# diff_3337_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3590 diff_3388_1325# diff_2512_1312# diff_3388_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3591 diff_3439_1325# diff_2512_1312# diff_3439_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3592 diff_3490_1325# diff_2512_1312# diff_3490_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3593 diff_3541_1325# diff_2512_1312# diff_3541_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3594 diff_3592_1325# diff_2512_1312# diff_3592_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3595 diff_3643_1325# diff_2512_1312# diff_3643_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3596 diff_3694_1325# diff_2512_1312# diff_3694_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3597 diff_3745_1325# diff_2512_1312# diff_3745_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3598 diff_3796_1325# diff_2512_1312# diff_3796_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3599 diff_3847_1325# diff_2512_1312# diff_3847_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3600 diff_3898_1325# diff_2512_1312# diff_3898_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3601 diff_3949_1325# diff_2512_1312# diff_3949_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3602 diff_4000_1325# diff_2512_1312# diff_4000_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3603 diff_4051_1325# diff_2512_1312# diff_4051_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3604 diff_4102_1325# diff_2512_1312# diff_4102_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3605 diff_4153_1325# diff_2512_1312# diff_4153_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3606 diff_4204_1325# diff_2512_1312# diff_4204_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3607 diff_4255_1325# diff_2512_1312# diff_4255_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3608 diff_4306_1325# diff_2512_1312# diff_4306_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3609 diff_4357_1325# diff_2512_1312# diff_4357_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3610 diff_4408_1325# diff_2512_1312# diff_4408_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3611 diff_4459_1325# diff_2512_1312# diff_4459_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3612 diff_4510_1325# diff_2512_1312# diff_4510_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3613 diff_4561_1325# diff_2512_1312# diff_4561_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3614 diff_4612_1325# diff_2512_1312# diff_4612_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3615 diff_4663_1325# diff_2512_1312# diff_4663_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3616 diff_4714_1325# diff_2512_1312# diff_4714_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3617 diff_4765_1325# diff_2512_1312# diff_4765_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3618 diff_4816_1325# diff_2512_1312# diff_4816_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3619 diff_4867_1325# diff_2512_1312# diff_4867_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3620 diff_4918_1325# diff_2512_1312# diff_4918_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3621 diff_4969_1325# diff_2512_1312# diff_4969_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3622 diff_5020_1325# diff_2512_1312# diff_5020_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3623 diff_5071_1325# diff_2512_1312# diff_5071_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3624 diff_5122_1325# diff_2512_1312# diff_5122_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3625 diff_5173_1325# diff_2512_1312# diff_5173_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3626 diff_5224_1325# diff_2512_1312# diff_5224_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3627 diff_5275_1325# diff_2512_1312# diff_5275_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3628 diff_5326_1325# diff_2512_1312# diff_5326_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3629 diff_5377_1325# diff_2512_1312# diff_5377_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3630 diff_5428_1325# diff_2512_1312# diff_5428_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3631 diff_5479_1325# diff_2512_1312# diff_5479_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3632 diff_5530_1325# diff_2512_1312# diff_5530_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3633 diff_5581_1325# diff_2512_1312# diff_5581_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3634 diff_5632_1325# diff_2512_1312# diff_5632_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3635 diff_5683_1325# diff_2512_1312# diff_5683_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3636 diff_5734_1325# diff_2512_1312# diff_5734_1271# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3637 diff_2512_1480# diff_5962_1069# diff_5918_1300# GND efet w=184 l=13
+ ad=0 pd=0 as=0 ps=0 
M3638 diff_2512_1423# Vdd Vdd GND efet w=16 l=31
+ ad=6288 pd=616 as=0 ps=0 
M3639 Vdd Vdd diff_2512_1369# GND efet w=16 l=34
+ ad=0 pd=0 as=6332 ps=552 
M3640 diff_5918_1300# diff_6034_2491# diff_2512_1369# GND efet w=209 l=14
+ ad=0 pd=0 as=0 ps=0 
M3641 diff_2521_1271# diff_2512_1258# diff_2521_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3642 diff_2572_1271# diff_2512_1258# diff_2572_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3643 diff_2623_1271# diff_2512_1258# diff_2623_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3644 diff_2674_1271# diff_2512_1258# diff_2674_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3645 diff_2725_1271# diff_2512_1258# diff_2725_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3646 diff_2776_1271# diff_2512_1258# diff_2776_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3647 diff_2827_1271# diff_2512_1258# diff_2827_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3648 diff_2878_1271# diff_2512_1258# diff_2878_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3649 diff_2929_1271# diff_2512_1258# diff_2929_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3650 diff_2980_1271# diff_2512_1258# diff_2980_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3651 diff_3031_1271# diff_2512_1258# diff_3031_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3652 diff_3082_1271# diff_2512_1258# diff_3082_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3653 diff_3133_1271# diff_2512_1258# diff_3133_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3654 diff_3184_1271# diff_2512_1258# diff_3184_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3655 diff_3235_1271# diff_2512_1258# diff_3235_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3656 diff_3286_1271# diff_2512_1258# diff_3286_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3657 diff_3337_1271# diff_2512_1258# diff_3337_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3658 diff_3388_1271# diff_2512_1258# diff_3388_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3659 diff_3439_1271# diff_2512_1258# diff_3439_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3660 diff_3490_1271# diff_2512_1258# diff_3490_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3661 diff_3541_1271# diff_2512_1258# diff_3541_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3662 diff_3592_1271# diff_2512_1258# diff_3592_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3663 diff_3643_1271# diff_2512_1258# diff_3643_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3664 diff_3694_1271# diff_2512_1258# diff_3694_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3665 diff_3745_1271# diff_2512_1258# diff_3745_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3666 diff_3796_1271# diff_2512_1258# diff_3796_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3667 diff_3847_1271# diff_2512_1258# diff_3847_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3668 diff_3898_1271# diff_2512_1258# diff_3898_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3669 diff_3949_1271# diff_2512_1258# diff_3949_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3670 diff_4000_1271# diff_2512_1258# diff_4000_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3671 diff_4051_1271# diff_2512_1258# diff_4051_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3672 diff_4102_1271# diff_2512_1258# diff_4102_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3673 diff_4153_1271# diff_2512_1258# diff_4153_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3674 diff_4204_1271# diff_2512_1258# diff_4204_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3675 diff_4255_1271# diff_2512_1258# diff_4255_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3676 diff_4306_1271# diff_2512_1258# diff_4306_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3677 diff_4357_1271# diff_2512_1258# diff_4357_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3678 diff_4408_1271# diff_2512_1258# diff_4408_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3679 diff_4459_1271# diff_2512_1258# diff_4459_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3680 diff_4510_1271# diff_2512_1258# diff_4510_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3681 diff_4561_1271# diff_2512_1258# diff_4561_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3682 diff_4612_1271# diff_2512_1258# diff_4612_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3683 diff_4663_1271# diff_2512_1258# diff_4663_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3684 diff_4714_1271# diff_2512_1258# diff_4714_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3685 diff_4765_1271# diff_2512_1258# diff_4765_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3686 diff_4816_1271# diff_2512_1258# diff_4816_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3687 diff_4867_1271# diff_2512_1258# diff_4867_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3688 diff_4918_1271# diff_2512_1258# diff_4918_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3689 diff_4969_1271# diff_2512_1258# diff_4969_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3690 diff_5020_1271# diff_2512_1258# diff_5020_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3691 diff_5071_1271# diff_2512_1258# diff_5071_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3692 diff_5122_1271# diff_2512_1258# diff_5122_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3693 diff_5173_1271# diff_2512_1258# diff_5173_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3694 diff_5224_1271# diff_2512_1258# diff_5224_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3695 diff_5275_1271# diff_2512_1258# diff_5275_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3696 diff_5326_1271# diff_2512_1258# diff_5326_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3697 diff_5377_1271# diff_2512_1258# diff_5377_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3698 diff_5428_1271# diff_2512_1258# diff_5428_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3699 diff_5479_1271# diff_2512_1258# diff_5479_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3700 diff_5530_1271# diff_2512_1258# diff_5530_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3701 diff_5581_1271# diff_2512_1258# diff_5581_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3702 diff_5632_1271# diff_2512_1258# diff_5632_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3703 diff_5683_1271# diff_2512_1258# diff_5683_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3704 diff_5734_1271# diff_2512_1258# diff_5734_1214# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3705 diff_2512_1423# diff_6079_2449# diff_5918_1300# GND efet w=196 l=13
+ ad=0 pd=0 as=0 ps=0 
M3706 Vdd Vdd Vdd GND efet w=11 l=17
+ ad=0 pd=0 as=0 ps=0 
M3707 Vdd Vdd diff_6223_2134# GND efet w=16 l=34
+ ad=0 pd=0 as=14777 ps=1056 
M3708 diff_6935_2506# Vdd Vdd GND efet w=16 l=79
+ ad=0 pd=0 as=0 ps=0 
M3709 diff_7123_2480# diff_6949_1216# diff_7123_2441# GND efet w=115 l=13
+ ad=0 pd=0 as=2990 ps=282 
M3710 Vdd Vdd Vdd GND efet w=5 l=9
+ ad=0 pd=0 as=0 ps=0 
M3711 Vdd Vdd Vdd GND efet w=3 l=7
+ ad=0 pd=0 as=0 ps=0 
M3712 Vdd Vdd diff_6935_2224# GND efet w=16 l=79
+ ad=0 pd=0 as=6025 ps=406 
M3713 diff_7123_2441# diff_6832_1375# GND GND efet w=115 l=13
+ ad=0 pd=0 as=0 ps=0 
M3714 diff_6845_2317# diff_6778_3391# diff_6325_2236# GND efet w=49 l=13
+ ad=0 pd=0 as=1893 ps=176 
M3715 diff_6935_2224# clk2 diff_6845_2317# GND efet w=49 l=13
+ ad=0 pd=0 as=0 ps=0 
M3716 diff_7046_2224# diff_6845_1381# diff_6935_2224# GND efet w=91 l=13
+ ad=5871 pd=490 as=0 ps=0 
M3717 diff_6845_2035# diff_6778_3391# diff_6496_1642# GND efet w=49 l=13
+ ad=3608 pd=344 as=1746 ps=170 
M3718 diff_6935_2131# clk2 diff_6845_2035# GND efet w=49 l=13
+ ad=7013 pd=524 as=0 ps=0 
M3719 Vdd Vdd diff_2623_2116# GND efet w=16 l=31
+ ad=0 pd=0 as=11162 ps=810 
M3720 Vdd Vdd diff_2488_3064# GND efet w=16 l=31
+ ad=0 pd=0 as=13004 ps=822 
M3721 Vdd Vdd diff_6265_2299# GND efet w=19 l=31
+ ad=0 pd=0 as=12278 ps=816 
M3722 diff_6845_2035# diff_6808_2113# diff_6544_1975# GND efet w=49 l=13
+ ad=0 pd=0 as=1746 ps=170 
M3723 GND diff_6496_1642# diff_6223_2134# GND efet w=307 l=13
+ ad=0 pd=0 as=0 ps=0 
M3724 diff_2623_2116# diff_6544_1975# GND GND efet w=307 l=13
+ ad=0 pd=0 as=0 ps=0 
M3725 GND diff_6664_1975# diff_2488_3064# GND efet w=307 l=13
+ ad=0 pd=0 as=0 ps=0 
M3726 diff_6265_2299# diff_6718_1975# GND GND efet w=307 l=13
+ ad=0 pd=0 as=0 ps=0 
M3727 diff_6845_1942# diff_6808_2113# diff_6664_1975# GND efet w=49 l=13
+ ad=3731 pd=350 as=1746 ps=170 
M3728 diff_6935_2131# Vdd Vdd GND efet w=16 l=82
+ ad=0 pd=0 as=0 ps=0 
M3729 Vdd Vdd Vdd GND efet w=6 l=13
+ ad=0 pd=0 as=0 ps=0 
M3730 Vdd Vdd Vdd GND efet w=2 l=9
+ ad=0 pd=0 as=0 ps=0 
M3731 Vdd Vdd diff_6935_1846# GND efet w=16 l=79
+ ad=0 pd=0 as=6271 ps=406 
M3732 diff_7163_2251# diff_6832_1375# diff_6935_2506# GND efet w=94 l=13
+ ad=2444 pd=240 as=0 ps=0 
M3733 GND diff_6880_1132# diff_7163_2251# GND efet w=94 l=13
+ ad=0 pd=0 as=0 ps=0 
M3734 d0 GND d0 GND efet w=449 l=275
+ ad=0 pd=0 as=0 ps=0 
M3735 GND diff_6880_1132# diff_7046_2224# GND efet w=88 l=13
+ ad=0 pd=0 as=0 ps=0 
M3736 diff_7103_1999# diff_6949_1216# diff_6935_2131# GND efet w=88 l=13
+ ad=2288 pd=228 as=0 ps=0 
M3737 GND diff_6832_1375# diff_7103_1999# GND efet w=88 l=13
+ ad=0 pd=0 as=0 ps=0 
M3738 diff_6845_1942# diff_6778_3391# diff_6718_1975# GND efet w=52 l=13
+ ad=0 pd=0 as=1992 ps=182 
M3739 diff_6935_1846# clk2 diff_6845_1942# GND efet w=52 l=13
+ ad=0 pd=0 as=0 ps=0 
M3740 diff_7046_1846# diff_6845_1381# diff_6935_1846# GND efet w=94 l=13
+ ad=2444 pd=240 as=0 ps=0 
M3741 GND diff_6949_1216# diff_7046_1846# GND efet w=94 l=13
+ ad=0 pd=0 as=0 ps=0 
M3742 Vdd Vdd Vdd GND efet w=5 l=8
+ ad=0 pd=0 as=0 ps=0 
M3743 Vdd Vdd Vdd GND efet w=5 l=9
+ ad=0 pd=0 as=0 ps=0 
M3744 diff_6832_1375# Vdd Vdd GND efet w=25 l=40
+ ad=10925 pd=846 as=0 ps=0 
M3745 GND diff_6085_4357# diff_6269_1078# GND efet w=751 l=13
+ ad=0 pd=0 as=0 ps=0 
M3746 diff_5918_1078# diff_5905_1069# diff_2512_1090# GND efet w=221 l=16
+ ad=24382 pd=1728 as=5294 ps=570 
M3747 diff_2521_1214# diff_2512_1201# diff_2521_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3748 diff_2572_1214# diff_2512_1201# diff_2572_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3749 diff_2623_1214# diff_2512_1201# diff_2623_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3750 diff_2674_1214# diff_2512_1201# diff_2674_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3751 diff_2725_1214# diff_2512_1201# diff_2725_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3752 diff_2776_1214# diff_2512_1201# diff_2776_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3753 diff_2827_1214# diff_2512_1201# diff_2827_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3754 diff_2878_1214# diff_2512_1201# diff_2878_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3755 diff_2929_1214# diff_2512_1201# diff_2929_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3756 diff_2980_1214# diff_2512_1201# diff_2980_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3757 diff_3031_1214# diff_2512_1201# diff_3031_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3758 diff_3082_1214# diff_2512_1201# diff_3082_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3759 diff_3133_1214# diff_2512_1201# diff_3133_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3760 diff_3184_1214# diff_2512_1201# diff_3184_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3761 diff_3235_1214# diff_2512_1201# diff_3235_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3762 diff_3286_1214# diff_2512_1201# diff_3286_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3763 diff_3337_1214# diff_2512_1201# diff_3337_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3764 diff_3388_1214# diff_2512_1201# diff_3388_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3765 diff_3439_1214# diff_2512_1201# diff_3439_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3766 diff_3490_1214# diff_2512_1201# diff_3490_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3767 diff_3541_1214# diff_2512_1201# diff_3541_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3768 diff_3592_1214# diff_2512_1201# diff_3592_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3769 diff_3643_1214# diff_2512_1201# diff_3643_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3770 diff_3694_1214# diff_2512_1201# diff_3694_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3771 diff_3745_1214# diff_2512_1201# diff_3745_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3772 diff_3796_1214# diff_2512_1201# diff_3796_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3773 diff_3847_1214# diff_2512_1201# diff_3847_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3774 diff_3898_1214# diff_2512_1201# diff_3898_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3775 diff_3949_1214# diff_2512_1201# diff_3949_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3776 diff_4000_1214# diff_2512_1201# diff_4000_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3777 diff_4051_1214# diff_2512_1201# diff_4051_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3778 diff_4102_1214# diff_2512_1201# diff_4102_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3779 diff_4153_1214# diff_2512_1201# diff_4153_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3780 diff_4204_1214# diff_2512_1201# diff_4204_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3781 diff_4255_1214# diff_2512_1201# diff_4255_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3782 diff_4306_1214# diff_2512_1201# diff_4306_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3783 diff_4357_1214# diff_2512_1201# diff_4357_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3784 diff_4408_1214# diff_2512_1201# diff_4408_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3785 diff_4459_1214# diff_2512_1201# diff_4459_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3786 diff_4510_1214# diff_2512_1201# diff_4510_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3787 diff_4561_1214# diff_2512_1201# diff_4561_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3788 diff_4612_1214# diff_2512_1201# diff_4612_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3789 diff_4663_1214# diff_2512_1201# diff_4663_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3790 diff_4714_1214# diff_2512_1201# diff_4714_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3791 diff_4765_1214# diff_2512_1201# diff_4765_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3792 diff_4816_1214# diff_2512_1201# diff_4816_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3793 diff_4867_1214# diff_2512_1201# diff_4867_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3794 diff_4918_1214# diff_2512_1201# diff_4918_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3795 diff_4969_1214# diff_2512_1201# diff_4969_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3796 diff_5020_1214# diff_2512_1201# diff_5020_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3797 diff_5071_1214# diff_2512_1201# diff_5071_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3798 diff_5122_1214# diff_2512_1201# diff_5122_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3799 diff_5173_1214# diff_2512_1201# diff_5173_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3800 diff_5224_1214# diff_2512_1201# diff_5224_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3801 diff_5275_1214# diff_2512_1201# diff_5275_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3802 diff_5326_1214# diff_2512_1201# diff_5326_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3803 diff_5377_1214# diff_2512_1201# diff_5377_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3804 diff_5428_1214# diff_2512_1201# diff_5428_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3805 diff_5479_1214# diff_2512_1201# diff_5479_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3806 diff_5530_1214# diff_2512_1201# diff_5530_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3807 diff_5581_1214# diff_2512_1201# diff_5581_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3808 diff_5632_1214# diff_2512_1201# diff_5632_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3809 diff_5683_1214# diff_2512_1201# diff_5683_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3810 diff_5734_1214# diff_2512_1201# diff_5734_1160# GND efet w=25 l=16
+ ad=0 pd=0 as=950 ps=126 
M3811 diff_2512_1258# Vdd Vdd GND efet w=13 l=28
+ ad=5625 pd=646 as=0 ps=0 
M3812 GND cm diff_2306_1147# GND efet w=166 l=16
+ ad=0 pd=0 as=0 ps=0 
M3813 diff_1729_1183# diff_1724_997# GND GND efet w=49 l=16
+ ad=4867 pd=520 as=0 ps=0 
M3814 diff_1873_938# diff_1832_997# GND GND efet w=46 l=16
+ ad=4384 pd=484 as=0 ps=0 
M3815 diff_1990_938# diff_1949_997# GND GND efet w=49 l=16
+ ad=4006 pd=472 as=0 ps=0 
M3816 diff_1034_997# diff_1034_997# diff_1034_997# GND efet w=1 l=2
+ ad=0 pd=0 as=0 ps=0 
M3817 diff_1148_997# clk2 diff_1075_938# GND efet w=28 l=16
+ ad=818 pd=116 as=0 ps=0 
M3818 diff_1148_997# diff_1148_997# diff_1148_997# GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M3819 diff_1265_997# clk1 diff_1186_938# GND efet w=28 l=16
+ ad=787 pd=124 as=0 ps=0 
M3820 diff_1265_997# diff_1265_997# diff_1265_997# GND efet w=5 l=8
+ ad=0 pd=0 as=0 ps=0 
M3821 diff_1265_997# diff_1265_997# diff_1265_997# GND efet w=1 l=2
+ ad=0 pd=0 as=0 ps=0 
M3822 diff_1376_997# clk2 diff_1198_1177# GND efet w=28 l=16
+ ad=889 pd=124 as=0 ps=0 
M3823 diff_1376_997# diff_1376_997# diff_1376_997# GND efet w=2 l=4
+ ad=0 pd=0 as=0 ps=0 
M3824 diff_1376_997# diff_1376_997# diff_1376_997# GND efet w=0 l=1
+ ad=0 pd=0 as=0 ps=0 
M3825 diff_1493_997# clk1 diff_1378_1138# GND efet w=28 l=16
+ ad=871 pd=130 as=0 ps=0 
M3826 diff_1493_997# diff_1493_997# diff_1493_997# GND efet w=5 l=8
+ ad=0 pd=0 as=0 ps=0 
M3827 diff_1493_997# diff_1493_997# diff_1493_997# GND efet w=1 l=2
+ ad=0 pd=0 as=0 ps=0 
M3828 diff_1607_997# clk2 diff_1534_938# GND efet w=28 l=16
+ ad=818 pd=116 as=0 ps=0 
M3829 diff_1607_997# diff_1607_997# diff_1607_997# GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M3830 diff_1724_997# clk1 diff_1555_1174# GND efet w=28 l=16
+ ad=763 pd=130 as=0 ps=0 
M3831 diff_1724_997# diff_1724_997# diff_1724_997# GND efet w=5 l=10
+ ad=0 pd=0 as=0 ps=0 
M3832 diff_1724_997# diff_1724_997# diff_1724_997# GND efet w=2 l=4
+ ad=0 pd=0 as=0 ps=0 
M3833 diff_1832_997# clk2 diff_1729_1183# GND efet w=28 l=16
+ ad=889 pd=124 as=0 ps=0 
M3834 diff_1832_997# diff_1832_997# diff_1832_997# GND efet w=2 l=4
+ ad=0 pd=0 as=0 ps=0 
M3835 diff_1832_997# diff_1832_997# diff_1832_997# GND efet w=0 l=1
+ ad=0 pd=0 as=0 ps=0 
M3836 diff_1949_997# clk1 diff_1873_938# GND efet w=28 l=16
+ ad=871 pd=130 as=0 ps=0 
M3837 diff_1949_997# diff_1949_997# diff_1949_997# GND efet w=5 l=8
+ ad=0 pd=0 as=0 ps=0 
M3838 diff_2101_938# diff_2063_997# GND GND efet w=46 l=16
+ ad=4846 pd=526 as=0 ps=0 
M3839 diff_1867_1564# diff_2180_997# GND GND efet w=49 l=13
+ ad=4352 pd=498 as=0 ps=0 
M3840 diff_2521_1160# diff_2512_1147# diff_2521_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3841 diff_2572_1160# diff_2512_1147# diff_2572_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3842 diff_2623_1160# diff_2512_1147# diff_2623_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3843 diff_2674_1160# diff_2512_1147# diff_2674_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3844 diff_2725_1160# diff_2512_1147# diff_2725_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3845 diff_2776_1160# diff_2512_1147# diff_2776_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3846 diff_2827_1160# diff_2512_1147# diff_2827_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3847 diff_2878_1160# diff_2512_1147# diff_2878_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3848 diff_2929_1160# diff_2512_1147# diff_2929_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3849 diff_2980_1160# diff_2512_1147# diff_2980_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3850 diff_3031_1160# diff_2512_1147# diff_3031_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3851 diff_3082_1160# diff_2512_1147# diff_3082_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3852 diff_3133_1160# diff_2512_1147# diff_3133_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3853 diff_3184_1160# diff_2512_1147# diff_3184_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3854 diff_3235_1160# diff_2512_1147# diff_3235_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3855 diff_3286_1160# diff_2512_1147# diff_3286_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3856 diff_3337_1160# diff_2512_1147# diff_3337_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3857 diff_3388_1160# diff_2512_1147# diff_3388_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3858 diff_3439_1160# diff_2512_1147# diff_3439_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3859 diff_3490_1160# diff_2512_1147# diff_3490_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3860 diff_3541_1160# diff_2512_1147# diff_3541_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3861 diff_3592_1160# diff_2512_1147# diff_3592_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3862 diff_3643_1160# diff_2512_1147# diff_3643_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3863 diff_3694_1160# diff_2512_1147# diff_3694_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3864 diff_3745_1160# diff_2512_1147# diff_3745_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3865 diff_3796_1160# diff_2512_1147# diff_3796_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3866 diff_3847_1160# diff_2512_1147# diff_3847_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3867 diff_3898_1160# diff_2512_1147# diff_3898_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3868 diff_3949_1160# diff_2512_1147# diff_3949_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3869 diff_4000_1160# diff_2512_1147# diff_4000_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3870 diff_4051_1160# diff_2512_1147# diff_4051_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3871 diff_4102_1160# diff_2512_1147# diff_4102_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3872 diff_4153_1160# diff_2512_1147# diff_4153_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3873 diff_4204_1160# diff_2512_1147# diff_4204_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3874 diff_4255_1160# diff_2512_1147# diff_4255_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3875 diff_4306_1160# diff_2512_1147# diff_4306_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3876 diff_4357_1160# diff_2512_1147# diff_4357_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3877 diff_4408_1160# diff_2512_1147# diff_4408_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3878 diff_4459_1160# diff_2512_1147# diff_4459_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3879 diff_4510_1160# diff_2512_1147# diff_4510_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3880 diff_4561_1160# diff_2512_1147# diff_4561_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3881 diff_4612_1160# diff_2512_1147# diff_4612_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3882 diff_4663_1160# diff_2512_1147# diff_4663_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3883 diff_4714_1160# diff_2512_1147# diff_4714_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3884 diff_4765_1160# diff_2512_1147# diff_4765_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3885 diff_4816_1160# diff_2512_1147# diff_4816_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3886 diff_4867_1160# diff_2512_1147# diff_4867_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3887 diff_4918_1160# diff_2512_1147# diff_4918_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3888 diff_4969_1160# diff_2512_1147# diff_4969_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3889 diff_5020_1160# diff_2512_1147# diff_5020_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3890 diff_5071_1160# diff_2512_1147# diff_5071_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3891 diff_5122_1160# diff_2512_1147# diff_5122_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3892 diff_5173_1160# diff_2512_1147# diff_5173_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3893 diff_5224_1160# diff_2512_1147# diff_5224_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3894 diff_5275_1160# diff_2512_1147# diff_5275_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3895 diff_5326_1160# diff_2512_1147# diff_5326_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3896 diff_5377_1160# diff_2512_1147# diff_5377_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3897 diff_5428_1160# diff_2512_1147# diff_5428_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3898 diff_5479_1160# diff_2512_1147# diff_5479_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3899 diff_5530_1160# diff_2512_1147# diff_5530_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3900 diff_5581_1160# diff_2512_1147# diff_5581_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3901 diff_5632_1160# diff_2512_1147# diff_5632_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3902 diff_5683_1160# diff_2512_1147# diff_5683_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3903 diff_5734_1160# diff_2512_1147# diff_5734_1103# GND efet w=25 l=16
+ ad=0 pd=0 as=1025 ps=132 
M3904 diff_1949_997# diff_1949_997# diff_1949_997# GND efet w=1 l=2
+ ad=0 pd=0 as=0 ps=0 
M3905 diff_2063_997# clk2 diff_1990_938# GND efet w=28 l=16
+ ad=818 pd=116 as=0 ps=0 
M3906 diff_2063_997# diff_2063_997# diff_2063_997# GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M3907 diff_2180_997# clk1 diff_2101_938# GND efet w=28 l=16
+ ad=799 pd=126 as=0 ps=0 
M3908 diff_2180_997# diff_2180_997# diff_2180_997# GND efet w=4 l=5
+ ad=0 pd=0 as=0 ps=0 
M3909 diff_2180_997# diff_2180_997# diff_2180_997# GND efet w=1 l=2
+ ad=0 pd=0 as=0 ps=0 
M3910 Vdd Vdd diff_724_1144# GND efet w=17 l=86
+ ad=0 pd=0 as=0 ps=0 
M3911 diff_847_938# Vdd Vdd GND efet w=16 l=85
+ ad=0 pd=0 as=0 ps=0 
M3912 Vdd Vdd diff_958_938# GND efet w=17 l=89
+ ad=0 pd=0 as=0 ps=0 
M3913 diff_1075_938# Vdd Vdd GND efet w=16 l=82
+ ad=0 pd=0 as=0 ps=0 
M3914 Vdd Vdd diff_1186_938# GND efet w=17 l=92
+ ad=0 pd=0 as=0 ps=0 
M3915 diff_1198_1177# Vdd Vdd GND efet w=16 l=82
+ ad=0 pd=0 as=0 ps=0 
M3916 Vdd Vdd diff_1378_1138# GND efet w=17 l=89
+ ad=0 pd=0 as=0 ps=0 
M3917 diff_1534_938# Vdd Vdd GND efet w=16 l=82
+ ad=0 pd=0 as=0 ps=0 
M3918 Vdd Vdd diff_1555_1174# GND efet w=17 l=92
+ ad=0 pd=0 as=0 ps=0 
M3919 diff_1729_1183# Vdd Vdd GND efet w=16 l=85
+ ad=0 pd=0 as=0 ps=0 
M3920 Vdd Vdd diff_1873_938# GND efet w=17 l=89
+ ad=0 pd=0 as=0 ps=0 
M3921 diff_1990_938# Vdd Vdd GND efet w=16 l=82
+ ad=0 pd=0 as=0 ps=0 
M3922 Vdd Vdd diff_2101_938# GND efet w=17 l=92
+ ad=0 pd=0 as=0 ps=0 
M3923 diff_1867_1564# Vdd Vdd GND efet w=16 l=82
+ ad=0 pd=0 as=0 ps=0 
M3924 cl GND GND GND efet w=244 l=16
+ ad=23611 pd=2414 as=0 ps=0 
M3925 Vdd Vdd diff_2512_1090# GND efet w=13 l=28
+ ad=0 pd=0 as=0 ps=0 
M3926 diff_2521_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=124138 ps=7198 
M3927 diff_2572_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3928 diff_2623_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3929 diff_2674_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3930 diff_2725_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3931 diff_2776_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3932 diff_2827_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3933 diff_2878_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3934 diff_2929_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3935 diff_2980_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3936 diff_3031_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3937 diff_3082_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3938 diff_3133_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3939 diff_3184_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3940 diff_3235_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3941 diff_3286_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3942 diff_3337_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3943 diff_3388_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3944 diff_3439_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3945 diff_3490_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3946 diff_3541_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3947 diff_3592_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3948 diff_3643_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3949 diff_3694_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3950 diff_3745_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3951 diff_3796_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3952 diff_3847_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3953 diff_3898_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3954 diff_3949_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3955 diff_4000_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3956 diff_4051_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3957 diff_4102_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3958 diff_4153_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3959 diff_4204_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3960 diff_4255_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3961 diff_4306_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3962 diff_4357_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3963 diff_4408_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3964 diff_4459_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3965 diff_4510_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3966 diff_4561_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3967 diff_4612_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3968 diff_4663_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3969 diff_4714_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3970 diff_4765_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3971 diff_4816_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3972 diff_4867_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3973 diff_4918_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3974 diff_4969_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3975 diff_5020_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3976 diff_5071_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3977 diff_5122_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3978 diff_5173_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3979 diff_5224_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3980 diff_5275_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3981 diff_5326_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3982 diff_5377_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3983 diff_5428_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3984 diff_5479_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3985 diff_5530_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3986 diff_5581_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3987 diff_5632_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3988 diff_5683_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3989 diff_5734_1103# diff_2512_1090# diff_2521_1046# GND efet w=25 l=16
+ ad=0 pd=0 as=0 ps=0 
M3990 diff_2512_1258# diff_5962_1069# diff_5918_1078# GND efet w=184 l=13
+ ad=0 pd=0 as=0 ps=0 
M3991 diff_2512_1201# Vdd Vdd GND efet w=16 l=28
+ ad=6288 pd=616 as=0 ps=0 
M3992 Vdd Vdd diff_2512_1147# GND efet w=16 l=28
+ ad=0 pd=0 as=6050 ps=552 
M3993 diff_5918_1078# diff_6034_2491# diff_2512_1147# GND efet w=205 l=16
+ ad=0 pd=0 as=0 ps=0 
M3994 diff_2512_1201# diff_6079_2449# diff_5918_1078# GND efet w=196 l=13
+ ad=0 pd=0 as=0 ps=0 
M3995 diff_6269_1078# diff_6223_2134# diff_5918_1300# GND efet w=385 l=16
+ ad=0 pd=0 as=0 ps=0 
M3996 diff_5918_1078# diff_6265_2299# diff_6269_1078# GND efet w=403 l=16
+ ad=0 pd=0 as=0 ps=0 
M3997 diff_6832_1375# d0 GND GND efet w=427 l=13
+ ad=0 pd=0 as=0 ps=0 
M3998 diff_7148_1529# diff_6832_1375# diff_2380_1093# GND efet w=205 l=13
+ ad=5555 pd=468 as=19372 ps=1742 
M3999 diff_7081_2641# diff_6880_1132# diff_7148_1529# GND efet w=208 l=13
+ ad=0 pd=0 as=0 ps=0 
M4000 diff_6845_1381# diff_6832_1375# GND GND efet w=109 l=13
+ ad=4367 pd=388 as=0 ps=0 
M4001 diff_6845_1381# Vdd Vdd GND efet w=16 l=40
+ ad=0 pd=0 as=0 ps=0 
M4002 diff_6949_1216# Vdd Vdd GND efet w=22 l=40
+ ad=3581 pd=312 as=0 ps=0 
M4003 Vdd Vdd diff_6880_1132# GND efet w=16 l=43
+ ad=0 pd=0 as=13050 ps=1292 
M4004 GND diff_6880_1132# diff_6949_1216# GND efet w=109 l=13
+ ad=0 pd=0 as=0 ps=0 
M4005 diff_6880_1132# d1 GND GND efet w=427 l=13
+ ad=0 pd=0 as=0 ps=0 
M4006 GND diff_2380_1093# diff_1243_1231# GND efet w=46 l=16
+ ad=0 pd=0 as=0 ps=0 
M4007 diff_2521_1046# diff_2509_4258# GND GND efet w=1546 l=16
+ ad=0 pd=0 as=0 ps=0 
M4008 diff_2521_1046# diff_4144_4258# Vdd GND efet w=1606 l=16
+ ad=0 pd=0 as=0 ps=0 
M4009 Vdd Vdd Vdd GND efet w=6 l=10
+ ad=0 pd=0 as=0 ps=0 
M4010 Vdd Vdd Vdd GND efet w=5 l=13
+ ad=0 pd=0 as=0 ps=0 
M4011 Vdd Vdd diff_1243_1231# GND efet w=19 l=82
+ ad=0 pd=0 as=0 ps=0 
M4012 Vdd Vdd Vdd GND efet w=0 l=1
+ ad=0 pd=0 as=0 ps=0 
M4013 Vdd Vdd Vdd GND efet w=4 l=5
+ ad=0 pd=0 as=0 ps=0 
M4014 diff_2299_1054# Vdd Vdd GND efet w=17 l=101
+ ad=0 pd=0 as=0 ps=0 
M4015 Vdd Vdd diff_2380_1093# GND efet w=20 l=83
+ ad=0 pd=0 as=0 ps=0 
M4016 cm GND GND GND efet w=247 l=16
+ ad=20469 pd=1930 as=0 ps=0 
C0 metal_4573_463# gnd! 30.0fF ;**FLOATING
C1 metal_4528_472# gnd! 37.9fF ;**FLOATING
C2 metal_4273_391# gnd! 33.8fF ;**FLOATING
C3 metal_4258_391# gnd! 14.1fF ;**FLOATING
C4 metal_4324_448# gnd! 105.3fF ;**FLOATING
C5 metal_4144_418# gnd! 39.8fF ;**FLOATING
C6 metal_4258_469# gnd! 2.1fF ;**FLOATING
C7 metal_4486_394# gnd! 54.7fF ;**FLOATING
C8 metal_4459_463# gnd! 30.0fF ;**FLOATING
C9 metal_4123_409# gnd! 92.1fF ;**FLOATING
C10 metal_1030_409# gnd! 106.5fF ;**FLOATING
C11 metal_904_427# gnd! 224.7fF ;**FLOATING
C12 metal_781_433# gnd! 236.3fF ;**FLOATING
C13 metal_664_454# gnd! 216.0fF ;**FLOATING
C14 diff_6556_175# gnd! 18188.5fF ;**FLOATING
C15 diff_7148_1529# gnd! 602.3fF
C16 diff_2521_1046# gnd! 16143.9fF
C17 diff_2380_1093# gnd! 5445.9fF
C18 diff_5734_1103# gnd! 137.9fF
C19 diff_5683_1103# gnd! 137.9fF
C20 diff_5632_1103# gnd! 137.9fF
C21 diff_5581_1103# gnd! 137.9fF
C22 diff_5530_1103# gnd! 137.9fF
C23 diff_5479_1103# gnd! 137.9fF
C24 diff_5428_1103# gnd! 137.9fF
C25 diff_5377_1103# gnd! 137.9fF
C26 diff_5326_1103# gnd! 137.9fF
C27 diff_5275_1103# gnd! 137.9fF
C28 diff_5224_1103# gnd! 137.9fF
C29 diff_5173_1103# gnd! 137.9fF
C30 diff_5122_1103# gnd! 137.9fF
C31 diff_5071_1103# gnd! 137.9fF
C32 diff_5020_1103# gnd! 137.9fF
C33 diff_4969_1103# gnd! 137.9fF
C34 diff_4918_1103# gnd! 137.9fF
C35 diff_4867_1103# gnd! 137.9fF
C36 diff_4816_1103# gnd! 137.9fF
C37 diff_4765_1103# gnd! 137.9fF
C38 diff_4714_1103# gnd! 137.9fF
C39 diff_4663_1103# gnd! 137.9fF
C40 diff_4612_1103# gnd! 137.9fF
C41 diff_4561_1103# gnd! 137.9fF
C42 diff_4510_1103# gnd! 137.9fF
C43 diff_4459_1103# gnd! 137.9fF
C44 diff_4408_1103# gnd! 137.9fF
C45 diff_4357_1103# gnd! 137.9fF
C46 diff_4306_1103# gnd! 137.9fF
C47 diff_4255_1103# gnd! 137.9fF
C48 diff_4204_1103# gnd! 137.9fF
C49 diff_4153_1103# gnd! 137.9fF
C50 diff_4102_1103# gnd! 137.9fF
C51 diff_4051_1103# gnd! 137.9fF
C52 diff_4000_1103# gnd! 137.9fF
C53 diff_3949_1103# gnd! 137.9fF
C54 diff_3898_1103# gnd! 137.9fF
C55 diff_3847_1103# gnd! 137.9fF
C56 diff_3796_1103# gnd! 137.9fF
C57 diff_3745_1103# gnd! 137.9fF
C58 diff_3694_1103# gnd! 137.9fF
C59 diff_3643_1103# gnd! 137.9fF
C60 diff_3592_1103# gnd! 137.9fF
C61 diff_3541_1103# gnd! 137.9fF
C62 diff_3490_1103# gnd! 137.9fF
C63 diff_3439_1103# gnd! 137.9fF
C64 diff_3388_1103# gnd! 137.9fF
C65 diff_3337_1103# gnd! 137.9fF
C66 diff_3286_1103# gnd! 137.9fF
C67 diff_3235_1103# gnd! 137.9fF
C68 diff_3184_1103# gnd! 137.9fF
C69 diff_3133_1103# gnd! 137.9fF
C70 diff_3082_1103# gnd! 137.9fF
C71 diff_3031_1103# gnd! 137.9fF
C72 diff_2980_1103# gnd! 137.9fF
C73 diff_2929_1103# gnd! 137.9fF
C74 diff_2878_1103# gnd! 137.9fF
C75 diff_2827_1103# gnd! 137.9fF
C76 diff_2776_1103# gnd! 137.9fF
C77 diff_2725_1103# gnd! 137.9fF
C78 diff_2674_1103# gnd! 137.9fF
C79 diff_2623_1103# gnd! 137.9fF
C80 diff_2572_1103# gnd! 137.9fF
C81 diff_2521_1103# gnd! 137.9fF
C82 diff_2512_1147# gnd! 3500.1fF
C83 diff_5734_1160# gnd! 129.8fF
C84 diff_5683_1160# gnd! 129.8fF
C85 diff_5632_1160# gnd! 129.8fF
C86 diff_5581_1160# gnd! 129.8fF
C87 diff_5530_1160# gnd! 129.8fF
C88 diff_5479_1160# gnd! 129.8fF
C89 diff_5428_1160# gnd! 129.8fF
C90 diff_5377_1160# gnd! 129.8fF
C91 diff_5326_1160# gnd! 129.8fF
C92 diff_5275_1160# gnd! 129.8fF
C93 diff_5224_1160# gnd! 129.8fF
C94 diff_5173_1160# gnd! 129.8fF
C95 diff_5122_1160# gnd! 129.8fF
C96 diff_5071_1160# gnd! 129.8fF
C97 diff_5020_1160# gnd! 129.8fF
C98 diff_4969_1160# gnd! 129.8fF
C99 diff_4918_1160# gnd! 129.8fF
C100 diff_4867_1160# gnd! 129.8fF
C101 diff_4816_1160# gnd! 129.8fF
C102 diff_4765_1160# gnd! 129.8fF
C103 diff_4714_1160# gnd! 129.8fF
C104 diff_4663_1160# gnd! 129.8fF
C105 diff_4612_1160# gnd! 129.8fF
C106 diff_4561_1160# gnd! 129.8fF
C107 diff_4510_1160# gnd! 129.8fF
C108 diff_4459_1160# gnd! 129.8fF
C109 diff_4408_1160# gnd! 129.8fF
C110 diff_4357_1160# gnd! 129.8fF
C111 diff_4306_1160# gnd! 129.8fF
C112 diff_4255_1160# gnd! 129.8fF
C113 diff_4204_1160# gnd! 129.8fF
C114 diff_4153_1160# gnd! 129.8fF
C115 diff_4102_1160# gnd! 129.8fF
C116 diff_4051_1160# gnd! 129.8fF
C117 diff_4000_1160# gnd! 129.8fF
C118 diff_3949_1160# gnd! 129.8fF
C119 diff_3898_1160# gnd! 129.8fF
C120 diff_3847_1160# gnd! 129.8fF
C121 diff_3796_1160# gnd! 129.8fF
C122 diff_3745_1160# gnd! 129.8fF
C123 diff_3694_1160# gnd! 129.8fF
C124 diff_3643_1160# gnd! 129.8fF
C125 diff_3592_1160# gnd! 129.8fF
C126 diff_3541_1160# gnd! 129.8fF
C127 diff_3490_1160# gnd! 129.8fF
C128 diff_3439_1160# gnd! 129.8fF
C129 diff_3388_1160# gnd! 129.8fF
C130 diff_3337_1160# gnd! 129.8fF
C131 diff_3286_1160# gnd! 129.8fF
C132 diff_3235_1160# gnd! 129.8fF
C133 diff_3184_1160# gnd! 129.8fF
C134 diff_3133_1160# gnd! 129.8fF
C135 diff_3082_1160# gnd! 129.8fF
C136 diff_3031_1160# gnd! 129.8fF
C137 diff_2980_1160# gnd! 129.8fF
C138 diff_2929_1160# gnd! 129.8fF
C139 diff_2878_1160# gnd! 129.8fF
C140 diff_2827_1160# gnd! 129.8fF
C141 diff_2776_1160# gnd! 129.8fF
C142 diff_2725_1160# gnd! 129.8fF
C143 diff_2674_1160# gnd! 129.8fF
C144 diff_2623_1160# gnd! 129.8fF
C145 diff_2572_1160# gnd! 129.8fF
C146 diff_2180_997# gnd! 197.5fF
C147 diff_1990_938# gnd! 447.8fF
C148 diff_1873_938# gnd! 486.8fF
C149 diff_2063_997# gnd! 220.3fF
C150 diff_1949_997# gnd! 224.2fF
C151 diff_1832_997# gnd! 225.7fF
C152 diff_2521_1160# gnd! 129.8fF
C153 diff_2512_1201# gnd! 3605.4fF
C154 diff_5734_1214# gnd! 137.9fF
C155 diff_5683_1214# gnd! 137.9fF
C156 diff_5632_1214# gnd! 137.9fF
C157 diff_5581_1214# gnd! 137.9fF
C158 diff_5530_1214# gnd! 137.9fF
C159 diff_5479_1214# gnd! 137.9fF
C160 diff_5428_1214# gnd! 137.9fF
C161 diff_5377_1214# gnd! 137.9fF
C162 diff_5326_1214# gnd! 137.9fF
C163 diff_5275_1214# gnd! 137.9fF
C164 diff_5224_1214# gnd! 137.9fF
C165 diff_5173_1214# gnd! 137.9fF
C166 diff_5122_1214# gnd! 137.9fF
C167 diff_5071_1214# gnd! 137.9fF
C168 diff_5020_1214# gnd! 137.9fF
C169 diff_4969_1214# gnd! 137.9fF
C170 diff_4918_1214# gnd! 137.9fF
C171 diff_4867_1214# gnd! 137.9fF
C172 diff_4816_1214# gnd! 137.9fF
C173 diff_4765_1214# gnd! 137.9fF
C174 diff_4714_1214# gnd! 137.9fF
C175 diff_4663_1214# gnd! 137.9fF
C176 diff_4612_1214# gnd! 137.9fF
C177 diff_4561_1214# gnd! 137.9fF
C178 diff_4510_1214# gnd! 137.9fF
C179 diff_4459_1214# gnd! 137.9fF
C180 diff_4408_1214# gnd! 137.9fF
C181 diff_4357_1214# gnd! 137.9fF
C182 diff_4306_1214# gnd! 137.9fF
C183 diff_4255_1214# gnd! 137.9fF
C184 diff_4204_1214# gnd! 137.9fF
C185 diff_4153_1214# gnd! 137.9fF
C186 diff_4102_1214# gnd! 137.9fF
C187 diff_4051_1214# gnd! 137.9fF
C188 diff_4000_1214# gnd! 137.9fF
C189 diff_3949_1214# gnd! 137.9fF
C190 diff_3898_1214# gnd! 137.9fF
C191 diff_3847_1214# gnd! 137.9fF
C192 diff_3796_1214# gnd! 137.9fF
C193 diff_3745_1214# gnd! 137.9fF
C194 diff_3694_1214# gnd! 137.9fF
C195 diff_3643_1214# gnd! 137.9fF
C196 diff_3592_1214# gnd! 137.9fF
C197 diff_3541_1214# gnd! 137.9fF
C198 diff_3490_1214# gnd! 137.9fF
C199 diff_3439_1214# gnd! 137.9fF
C200 diff_3388_1214# gnd! 137.9fF
C201 diff_3337_1214# gnd! 137.9fF
C202 diff_3286_1214# gnd! 137.9fF
C203 diff_3235_1214# gnd! 137.9fF
C204 diff_3184_1214# gnd! 137.9fF
C205 diff_3133_1214# gnd! 137.9fF
C206 diff_3082_1214# gnd! 137.9fF
C207 diff_3031_1214# gnd! 137.9fF
C208 diff_2980_1214# gnd! 137.9fF
C209 diff_2929_1214# gnd! 137.9fF
C210 diff_2878_1214# gnd! 137.9fF
C211 diff_2827_1214# gnd! 137.9fF
C212 diff_2776_1214# gnd! 137.9fF
C213 diff_2725_1214# gnd! 137.9fF
C214 diff_2674_1214# gnd! 137.9fF
C215 diff_2623_1214# gnd! 137.9fF
C216 diff_2572_1214# gnd! 137.9fF
C217 diff_2521_1214# gnd! 137.9fF
C218 diff_5918_1078# gnd! 3009.8fF
C219 diff_2512_1090# gnd! 3302.5fF
C220 diff_7046_1846# gnd! 268.4fF
C221 diff_6935_1846# gnd! 667.7fF
C222 diff_7103_1999# gnd! 251.6fF
C223 diff_7163_2251# gnd! 268.4fF
C224 diff_6845_1942# gnd! 508.4fF
C225 diff_6718_1975# gnd! 619.1fF
C226 diff_6664_1975# gnd! 601.1fF
C227 diff_6544_1975# gnd! 667.7fF
C228 diff_6935_2131# gnd! 911.1fF
C229 diff_6845_2035# gnd! 493.8fF
C230 diff_6496_1642# gnd! 756.4fF
C231 diff_7046_2224# gnd! 805.2fF
C232 diff_6935_2224# gnd! 643.1fF
C233 diff_6845_1381# gnd! 1189.5fF
C234 diff_6880_1132# gnd! 2948.9fF
C235 diff_6832_1375# gnd! 2542.7fF
C236 diff_7123_2441# gnd! 327.2fF
C237 diff_6949_1216# gnd! 1808.1fF
C238 diff_7123_2480# gnd! 327.2fF
C239 diff_2512_1258# gnd! 3419.8fF
C240 diff_5734_1271# gnd! 129.8fF
C241 diff_5683_1271# gnd! 129.8fF
C242 diff_5632_1271# gnd! 129.8fF
C243 diff_5581_1271# gnd! 129.8fF
C244 diff_5530_1271# gnd! 129.8fF
C245 diff_5479_1271# gnd! 129.8fF
C246 diff_5428_1271# gnd! 129.8fF
C247 diff_5377_1271# gnd! 129.8fF
C248 diff_5326_1271# gnd! 129.8fF
C249 diff_5275_1271# gnd! 129.8fF
C250 diff_5224_1271# gnd! 129.8fF
C251 diff_5173_1271# gnd! 129.8fF
C252 diff_5122_1271# gnd! 129.8fF
C253 diff_5071_1271# gnd! 129.8fF
C254 diff_5020_1271# gnd! 129.8fF
C255 diff_4969_1271# gnd! 129.8fF
C256 diff_4918_1271# gnd! 129.8fF
C257 diff_4867_1271# gnd! 129.8fF
C258 diff_4816_1271# gnd! 129.8fF
C259 diff_4765_1271# gnd! 129.8fF
C260 diff_4714_1271# gnd! 129.8fF
C261 diff_4663_1271# gnd! 129.8fF
C262 diff_4612_1271# gnd! 129.8fF
C263 diff_4561_1271# gnd! 129.8fF
C264 diff_4510_1271# gnd! 129.8fF
C265 diff_4459_1271# gnd! 129.8fF
C266 diff_4408_1271# gnd! 129.8fF
C267 diff_4357_1271# gnd! 129.8fF
C268 diff_4306_1271# gnd! 129.8fF
C269 diff_4255_1271# gnd! 129.8fF
C270 diff_4204_1271# gnd! 129.8fF
C271 diff_4153_1271# gnd! 129.8fF
C272 diff_4102_1271# gnd! 129.8fF
C273 diff_4051_1271# gnd! 129.8fF
C274 diff_4000_1271# gnd! 129.8fF
C275 diff_3949_1271# gnd! 129.8fF
C276 diff_3898_1271# gnd! 129.8fF
C277 diff_3847_1271# gnd! 129.8fF
C278 diff_3796_1271# gnd! 129.8fF
C279 diff_3745_1271# gnd! 129.8fF
C280 diff_3694_1271# gnd! 129.8fF
C281 diff_3643_1271# gnd! 129.8fF
C282 diff_3592_1271# gnd! 129.8fF
C283 diff_3541_1271# gnd! 129.8fF
C284 diff_3490_1271# gnd! 129.8fF
C285 diff_3439_1271# gnd! 129.8fF
C286 diff_3388_1271# gnd! 129.8fF
C287 diff_3337_1271# gnd! 129.8fF
C288 diff_3286_1271# gnd! 129.8fF
C289 diff_3235_1271# gnd! 129.8fF
C290 diff_3184_1271# gnd! 129.8fF
C291 diff_3133_1271# gnd! 129.8fF
C292 diff_3082_1271# gnd! 129.8fF
C293 diff_3031_1271# gnd! 129.8fF
C294 diff_2980_1271# gnd! 129.8fF
C295 diff_2929_1271# gnd! 129.8fF
C296 diff_2878_1271# gnd! 129.8fF
C297 diff_2827_1271# gnd! 129.8fF
C298 diff_2776_1271# gnd! 129.8fF
C299 diff_2725_1271# gnd! 129.8fF
C300 diff_2674_1271# gnd! 129.8fF
C301 diff_2623_1271# gnd! 129.8fF
C302 diff_2572_1271# gnd! 129.8fF
C303 diff_2521_1271# gnd! 129.8fF
C304 diff_5734_1325# gnd! 137.9fF
C305 diff_5683_1325# gnd! 137.9fF
C306 diff_5632_1325# gnd! 137.9fF
C307 diff_5581_1325# gnd! 137.9fF
C308 diff_5530_1325# gnd! 137.9fF
C309 diff_5479_1325# gnd! 137.9fF
C310 diff_5428_1325# gnd! 137.9fF
C311 diff_5377_1325# gnd! 137.9fF
C312 diff_5326_1325# gnd! 137.9fF
C313 diff_5275_1325# gnd! 137.9fF
C314 diff_5224_1325# gnd! 137.9fF
C315 diff_5173_1325# gnd! 137.9fF
C316 diff_5122_1325# gnd! 137.9fF
C317 diff_5071_1325# gnd! 137.9fF
C318 diff_5020_1325# gnd! 137.9fF
C319 diff_4969_1325# gnd! 137.9fF
C320 diff_4918_1325# gnd! 137.9fF
C321 diff_4867_1325# gnd! 137.9fF
C322 diff_4816_1325# gnd! 137.9fF
C323 diff_4765_1325# gnd! 137.9fF
C324 diff_4714_1325# gnd! 137.9fF
C325 diff_4663_1325# gnd! 137.9fF
C326 diff_4612_1325# gnd! 137.9fF
C327 diff_4561_1325# gnd! 137.9fF
C328 diff_4510_1325# gnd! 137.9fF
C329 diff_4459_1325# gnd! 137.9fF
C330 diff_4408_1325# gnd! 137.9fF
C331 diff_4357_1325# gnd! 137.9fF
C332 diff_4306_1325# gnd! 137.9fF
C333 diff_4255_1325# gnd! 137.9fF
C334 diff_4204_1325# gnd! 137.9fF
C335 diff_4153_1325# gnd! 137.9fF
C336 diff_4102_1325# gnd! 137.9fF
C337 diff_4051_1325# gnd! 137.9fF
C338 diff_4000_1325# gnd! 137.9fF
C339 diff_3949_1325# gnd! 137.9fF
C340 diff_3898_1325# gnd! 137.9fF
C341 diff_3847_1325# gnd! 137.9fF
C342 diff_3796_1325# gnd! 137.9fF
C343 diff_3745_1325# gnd! 137.9fF
C344 diff_3694_1325# gnd! 137.9fF
C345 diff_3643_1325# gnd! 137.9fF
C346 diff_3592_1325# gnd! 137.9fF
C347 diff_3541_1325# gnd! 137.9fF
C348 diff_3490_1325# gnd! 137.9fF
C349 diff_3439_1325# gnd! 137.9fF
C350 diff_3388_1325# gnd! 137.9fF
C351 diff_3337_1325# gnd! 137.9fF
C352 diff_3286_1325# gnd! 137.9fF
C353 diff_3235_1325# gnd! 137.9fF
C354 diff_3184_1325# gnd! 137.9fF
C355 diff_3133_1325# gnd! 137.9fF
C356 diff_3082_1325# gnd! 137.9fF
C357 diff_3031_1325# gnd! 137.9fF
C358 diff_2980_1325# gnd! 137.9fF
C359 diff_2929_1325# gnd! 137.9fF
C360 diff_2878_1325# gnd! 137.9fF
C361 diff_2827_1325# gnd! 137.9fF
C362 diff_2776_1325# gnd! 137.9fF
C363 diff_2725_1325# gnd! 137.9fF
C364 diff_2674_1325# gnd! 137.9fF
C365 diff_2623_1325# gnd! 137.9fF
C366 diff_2572_1325# gnd! 137.9fF
C367 diff_2306_1147# gnd! 629.0fF
C368 diff_2261_1162# gnd! 206.3fF
C369 diff_1724_997# gnd! 208.6fF
C370 diff_1534_938# gnd! 447.8fF
C371 diff_1607_997# gnd! 222.6fF
C372 diff_1493_997# gnd! 221.9fF
C373 diff_1186_938# gnd! 481.4fF
C374 diff_1376_997# gnd! 227.9fF
C375 diff_1265_997# gnd! 212.9fF
C376 diff_1148_997# gnd! 222.6fF
C377 diff_1075_938# gnd! 447.8fF
C378 diff_958_938# gnd! 486.8fF
C379 diff_1034_997# gnd! 221.9fF
C380 diff_917_997# gnd! 227.9fF
C381 diff_803_997# gnd! 216.7fF
C382 diff_1555_1174# gnd! 768.6fF
C383 diff_1378_1138# gnd! 815.9fF
C384 diff_1729_1183# gnd! 731.5fF
C385 diff_1738_1196# gnd! 176.9fF
C386 diff_1252_1199# gnd! 219.5fF
C387 diff_1951_1117# gnd! 749.4fF
C388 diff_724_1144# gnd! 725.6fF
C389 diff_2026_1276# gnd! 560.8fF
C390 diff_2521_1325# gnd! 137.9fF
C391 diff_2512_1369# gnd! 3532.4fF
C392 diff_5734_1382# gnd! 129.8fF
C393 diff_5683_1382# gnd! 129.8fF
C394 diff_5632_1382# gnd! 129.8fF
C395 diff_5581_1382# gnd! 129.8fF
C396 diff_5530_1382# gnd! 129.8fF
C397 diff_5479_1382# gnd! 129.8fF
C398 diff_5428_1382# gnd! 129.8fF
C399 diff_5377_1382# gnd! 129.8fF
C400 diff_5326_1382# gnd! 129.8fF
C401 diff_5275_1382# gnd! 129.8fF
C402 diff_5224_1382# gnd! 129.8fF
C403 diff_5173_1382# gnd! 129.8fF
C404 diff_5122_1382# gnd! 129.8fF
C405 diff_5071_1382# gnd! 129.8fF
C406 diff_5020_1382# gnd! 129.8fF
C407 diff_4969_1382# gnd! 129.8fF
C408 diff_4918_1382# gnd! 129.8fF
C409 diff_4867_1382# gnd! 129.8fF
C410 diff_4816_1382# gnd! 129.8fF
C411 diff_4765_1382# gnd! 129.8fF
C412 diff_4714_1382# gnd! 129.8fF
C413 diff_4663_1382# gnd! 129.8fF
C414 diff_4612_1382# gnd! 129.8fF
C415 diff_4561_1382# gnd! 129.8fF
C416 diff_4510_1382# gnd! 129.8fF
C417 diff_4459_1382# gnd! 129.8fF
C418 diff_4408_1382# gnd! 129.8fF
C419 diff_4357_1382# gnd! 129.8fF
C420 diff_4306_1382# gnd! 129.8fF
C421 diff_4255_1382# gnd! 129.8fF
C422 diff_4204_1382# gnd! 129.8fF
C423 diff_4153_1382# gnd! 129.8fF
C424 diff_4102_1382# gnd! 129.8fF
C425 diff_4051_1382# gnd! 129.8fF
C426 diff_4000_1382# gnd! 129.8fF
C427 diff_3949_1382# gnd! 129.8fF
C428 diff_3898_1382# gnd! 129.8fF
C429 diff_3847_1382# gnd! 129.8fF
C430 diff_3796_1382# gnd! 129.8fF
C431 diff_3745_1382# gnd! 129.8fF
C432 diff_3694_1382# gnd! 129.8fF
C433 diff_3643_1382# gnd! 129.8fF
C434 diff_3592_1382# gnd! 129.8fF
C435 diff_3541_1382# gnd! 129.8fF
C436 diff_3490_1382# gnd! 129.8fF
C437 diff_3439_1382# gnd! 129.8fF
C438 diff_3388_1382# gnd! 129.8fF
C439 diff_3337_1382# gnd! 129.8fF
C440 diff_3286_1382# gnd! 129.8fF
C441 diff_3235_1382# gnd! 129.8fF
C442 diff_3184_1382# gnd! 129.8fF
C443 diff_3133_1382# gnd! 129.8fF
C444 diff_3082_1382# gnd! 129.8fF
C445 diff_3031_1382# gnd! 129.8fF
C446 diff_2980_1382# gnd! 129.8fF
C447 diff_2929_1382# gnd! 129.8fF
C448 diff_2878_1382# gnd! 129.8fF
C449 diff_2827_1382# gnd! 129.8fF
C450 diff_2776_1382# gnd! 129.8fF
C451 diff_2725_1382# gnd! 129.8fF
C452 diff_2674_1382# gnd! 129.8fF
C453 diff_2623_1382# gnd! 129.8fF
C454 diff_2572_1382# gnd! 129.8fF
C455 diff_2521_1382# gnd! 129.8fF
C456 diff_2512_1423# gnd! 3599.4fF
C457 diff_5734_1436# gnd! 137.9fF
C458 diff_5683_1436# gnd! 137.9fF
C459 diff_5632_1436# gnd! 137.9fF
C460 diff_5581_1436# gnd! 137.9fF
C461 diff_5530_1436# gnd! 137.9fF
C462 diff_5479_1436# gnd! 137.9fF
C463 diff_5428_1436# gnd! 137.9fF
C464 diff_5377_1436# gnd! 137.9fF
C465 diff_5326_1436# gnd! 137.9fF
C466 diff_5275_1436# gnd! 137.9fF
C467 diff_5224_1436# gnd! 137.9fF
C468 diff_5173_1436# gnd! 137.9fF
C469 diff_5122_1436# gnd! 137.9fF
C470 diff_5071_1436# gnd! 137.9fF
C471 diff_5020_1436# gnd! 137.9fF
C472 diff_4969_1436# gnd! 137.9fF
C473 diff_4918_1436# gnd! 137.9fF
C474 diff_4867_1436# gnd! 137.9fF
C475 diff_4816_1436# gnd! 137.9fF
C476 diff_4765_1436# gnd! 137.9fF
C477 diff_4714_1436# gnd! 137.9fF
C478 diff_4663_1436# gnd! 137.9fF
C479 diff_4612_1436# gnd! 137.9fF
C480 diff_4561_1436# gnd! 137.9fF
C481 diff_4510_1436# gnd! 137.9fF
C482 diff_4459_1436# gnd! 137.9fF
C483 diff_4408_1436# gnd! 137.9fF
C484 diff_4357_1436# gnd! 137.9fF
C485 diff_4306_1436# gnd! 137.9fF
C486 diff_4255_1436# gnd! 137.9fF
C487 diff_4204_1436# gnd! 137.9fF
C488 diff_4153_1436# gnd! 137.9fF
C489 diff_4102_1436# gnd! 137.9fF
C490 diff_4051_1436# gnd! 137.9fF
C491 diff_4000_1436# gnd! 137.9fF
C492 diff_3949_1436# gnd! 137.9fF
C493 diff_3898_1436# gnd! 137.9fF
C494 diff_3847_1436# gnd! 137.9fF
C495 diff_3796_1436# gnd! 137.9fF
C496 diff_3745_1436# gnd! 137.9fF
C497 diff_3694_1436# gnd! 137.9fF
C498 diff_3643_1436# gnd! 137.9fF
C499 diff_3592_1436# gnd! 137.9fF
C500 diff_3541_1436# gnd! 137.9fF
C501 diff_3490_1436# gnd! 137.9fF
C502 diff_3439_1436# gnd! 137.9fF
C503 diff_3388_1436# gnd! 137.9fF
C504 diff_3337_1436# gnd! 137.9fF
C505 diff_3286_1436# gnd! 137.9fF
C506 diff_3235_1436# gnd! 137.9fF
C507 diff_3184_1436# gnd! 137.9fF
C508 diff_3133_1436# gnd! 137.9fF
C509 diff_3082_1436# gnd! 137.9fF
C510 diff_3031_1436# gnd! 137.9fF
C511 diff_2980_1436# gnd! 137.9fF
C512 diff_2929_1436# gnd! 137.9fF
C513 diff_2878_1436# gnd! 137.9fF
C514 diff_2827_1436# gnd! 137.9fF
C515 diff_2776_1436# gnd! 137.9fF
C516 diff_2725_1436# gnd! 137.9fF
C517 diff_2674_1436# gnd! 137.9fF
C518 diff_2623_1436# gnd! 137.9fF
C519 diff_2572_1436# gnd! 137.9fF
C520 diff_2521_1436# gnd! 137.9fF
C521 diff_5918_1300# gnd! 2770.8fF
C522 diff_2512_1312# gnd! 3268.1fF
C523 diff_6269_1078# gnd! 5769.5fF
C524 diff_2512_1480# gnd! 3414.0fF
C525 diff_5734_1493# gnd! 129.8fF
C526 diff_5683_1493# gnd! 129.8fF
C527 diff_5632_1493# gnd! 129.8fF
C528 diff_5581_1493# gnd! 129.8fF
C529 diff_5530_1493# gnd! 129.8fF
C530 diff_5479_1493# gnd! 129.8fF
C531 diff_5428_1493# gnd! 129.8fF
C532 diff_5377_1493# gnd! 129.8fF
C533 diff_5326_1493# gnd! 129.8fF
C534 diff_5275_1493# gnd! 129.8fF
C535 diff_5224_1493# gnd! 129.8fF
C536 diff_5173_1493# gnd! 129.8fF
C537 diff_5122_1493# gnd! 129.8fF
C538 diff_5071_1493# gnd! 129.8fF
C539 diff_5020_1493# gnd! 129.8fF
C540 diff_4969_1493# gnd! 129.8fF
C541 diff_4918_1493# gnd! 129.8fF
C542 diff_4867_1493# gnd! 129.8fF
C543 diff_4816_1493# gnd! 129.8fF
C544 diff_4765_1493# gnd! 129.8fF
C545 diff_4714_1493# gnd! 129.8fF
C546 diff_4663_1493# gnd! 129.8fF
C547 diff_4612_1493# gnd! 129.8fF
C548 diff_4561_1493# gnd! 129.8fF
C549 diff_4510_1493# gnd! 129.8fF
C550 diff_4459_1493# gnd! 129.8fF
C551 diff_4408_1493# gnd! 129.8fF
C552 diff_4357_1493# gnd! 129.8fF
C553 diff_4306_1493# gnd! 129.8fF
C554 diff_4255_1493# gnd! 129.8fF
C555 diff_4204_1493# gnd! 129.8fF
C556 diff_4153_1493# gnd! 129.8fF
C557 diff_4102_1493# gnd! 129.8fF
C558 diff_4051_1493# gnd! 129.8fF
C559 diff_4000_1493# gnd! 129.8fF
C560 diff_3949_1493# gnd! 129.8fF
C561 diff_3898_1493# gnd! 129.8fF
C562 diff_3847_1493# gnd! 129.8fF
C563 diff_3796_1493# gnd! 129.8fF
C564 diff_3745_1493# gnd! 129.8fF
C565 diff_3694_1493# gnd! 129.8fF
C566 diff_3643_1493# gnd! 129.8fF
C567 diff_3592_1493# gnd! 129.8fF
C568 diff_3541_1493# gnd! 129.8fF
C569 diff_3490_1493# gnd! 129.8fF
C570 diff_3439_1493# gnd! 129.8fF
C571 diff_3388_1493# gnd! 129.8fF
C572 diff_3337_1493# gnd! 129.8fF
C573 diff_3286_1493# gnd! 129.8fF
C574 diff_3235_1493# gnd! 129.8fF
C575 diff_3184_1493# gnd! 129.8fF
C576 diff_3133_1493# gnd! 129.8fF
C577 diff_3082_1493# gnd! 129.8fF
C578 diff_3031_1493# gnd! 129.8fF
C579 diff_2980_1493# gnd! 129.8fF
C580 diff_2929_1493# gnd! 129.8fF
C581 diff_2878_1493# gnd! 129.8fF
C582 diff_2827_1493# gnd! 129.8fF
C583 diff_2776_1493# gnd! 129.8fF
C584 diff_2725_1493# gnd! 129.8fF
C585 diff_2674_1493# gnd! 129.8fF
C586 diff_2623_1493# gnd! 129.8fF
C587 diff_2572_1493# gnd! 129.8fF
C588 diff_1942_1222# gnd! 573.4fF
C589 diff_1729_1219# gnd! 784.6fF
C590 diff_1891_1138# gnd! 554.3fF
C591 diff_2521_1493# gnd! 129.8fF
C592 diff_1738_1232# gnd! 500.0fF
C593 diff_1187_1252# gnd! 82.1fF
C594 diff_1012_1177# gnd! 370.1fF
C595 diff_1226_1252# gnd! 281.9fF
C596 diff_1198_1177# gnd! 799.5fF
C597 diff_1243_1231# gnd! 1948.6fF
C598 cm gnd! 7433.1fF
C599 diff_5918_1519# gnd! 3153.4fF
C600 diff_5734_1547# gnd! 137.9fF
C601 diff_5683_1547# gnd! 137.9fF
C602 diff_5632_1547# gnd! 137.9fF
C603 diff_5581_1547# gnd! 137.9fF
C604 diff_5530_1547# gnd! 137.9fF
C605 diff_5479_1547# gnd! 137.9fF
C606 diff_5428_1547# gnd! 137.9fF
C607 diff_5377_1547# gnd! 137.9fF
C608 diff_5326_1547# gnd! 137.9fF
C609 diff_5275_1547# gnd! 137.9fF
C610 diff_5224_1547# gnd! 137.9fF
C611 diff_5173_1547# gnd! 137.9fF
C612 diff_5122_1547# gnd! 137.9fF
C613 diff_5071_1547# gnd! 137.9fF
C614 diff_5020_1547# gnd! 137.9fF
C615 diff_4969_1547# gnd! 137.9fF
C616 diff_4918_1547# gnd! 137.9fF
C617 diff_4867_1547# gnd! 137.9fF
C618 diff_4816_1547# gnd! 137.9fF
C619 diff_4765_1547# gnd! 137.9fF
C620 diff_4714_1547# gnd! 137.9fF
C621 diff_4663_1547# gnd! 137.9fF
C622 diff_4612_1547# gnd! 137.9fF
C623 diff_4561_1547# gnd! 137.9fF
C624 diff_4510_1547# gnd! 137.9fF
C625 diff_4459_1547# gnd! 137.9fF
C626 diff_4408_1547# gnd! 137.9fF
C627 diff_4357_1547# gnd! 137.9fF
C628 diff_4306_1547# gnd! 137.9fF
C629 diff_4255_1547# gnd! 137.9fF
C630 diff_4204_1547# gnd! 137.9fF
C631 diff_4153_1547# gnd! 137.9fF
C632 diff_4102_1547# gnd! 137.9fF
C633 diff_4051_1547# gnd! 137.9fF
C634 diff_4000_1547# gnd! 137.9fF
C635 diff_3949_1547# gnd! 137.9fF
C636 diff_3898_1547# gnd! 137.9fF
C637 diff_3847_1547# gnd! 137.9fF
C638 diff_3796_1547# gnd! 137.9fF
C639 diff_3745_1547# gnd! 137.9fF
C640 diff_3694_1547# gnd! 137.9fF
C641 diff_3643_1547# gnd! 137.9fF
C642 diff_3592_1547# gnd! 137.9fF
C643 diff_3541_1547# gnd! 137.9fF
C644 diff_3490_1547# gnd! 137.9fF
C645 diff_3439_1547# gnd! 137.9fF
C646 diff_3388_1547# gnd! 137.9fF
C647 diff_3337_1547# gnd! 137.9fF
C648 diff_3286_1547# gnd! 137.9fF
C649 diff_3235_1547# gnd! 137.9fF
C650 diff_3184_1547# gnd! 137.9fF
C651 diff_3133_1547# gnd! 137.9fF
C652 diff_3082_1547# gnd! 137.9fF
C653 diff_3031_1547# gnd! 137.9fF
C654 diff_2980_1547# gnd! 137.9fF
C655 diff_2929_1547# gnd! 137.9fF
C656 diff_2878_1547# gnd! 137.9fF
C657 diff_2827_1547# gnd! 137.9fF
C658 diff_2776_1547# gnd! 137.9fF
C659 diff_2725_1547# gnd! 137.9fF
C660 diff_2674_1547# gnd! 137.9fF
C661 diff_2623_1547# gnd! 137.9fF
C662 diff_2572_1547# gnd! 137.9fF
C663 diff_2521_1547# gnd! 137.9fF
C664 diff_2512_1591# gnd! 3555.8fF
C665 diff_5734_1604# gnd! 129.8fF
C666 diff_5683_1604# gnd! 129.8fF
C667 diff_5632_1604# gnd! 129.8fF
C668 diff_5581_1604# gnd! 129.8fF
C669 diff_5530_1604# gnd! 129.8fF
C670 diff_5479_1604# gnd! 129.8fF
C671 diff_5428_1604# gnd! 129.8fF
C672 diff_5377_1604# gnd! 129.8fF
C673 diff_5326_1604# gnd! 129.8fF
C674 diff_5275_1604# gnd! 129.8fF
C675 diff_5224_1604# gnd! 129.8fF
C676 diff_5173_1604# gnd! 129.8fF
C677 diff_5122_1604# gnd! 129.8fF
C678 diff_5071_1604# gnd! 129.8fF
C679 diff_5020_1604# gnd! 129.8fF
C680 diff_4969_1604# gnd! 129.8fF
C681 diff_4918_1604# gnd! 129.8fF
C682 diff_4867_1604# gnd! 129.8fF
C683 diff_4816_1604# gnd! 129.8fF
C684 diff_4765_1604# gnd! 129.8fF
C685 diff_4714_1604# gnd! 129.8fF
C686 diff_4663_1604# gnd! 129.8fF
C687 diff_4612_1604# gnd! 129.8fF
C688 diff_4561_1604# gnd! 129.8fF
C689 diff_4510_1604# gnd! 129.8fF
C690 diff_4459_1604# gnd! 129.8fF
C691 diff_4408_1604# gnd! 129.8fF
C692 diff_4357_1604# gnd! 129.8fF
C693 diff_4306_1604# gnd! 129.8fF
C694 diff_4255_1604# gnd! 129.8fF
C695 diff_4204_1604# gnd! 129.8fF
C696 diff_4153_1604# gnd! 129.8fF
C697 diff_4102_1604# gnd! 129.8fF
C698 diff_4051_1604# gnd! 129.8fF
C699 diff_4000_1604# gnd! 129.8fF
C700 diff_3949_1604# gnd! 129.8fF
C701 diff_3898_1604# gnd! 129.8fF
C702 diff_3847_1604# gnd! 129.8fF
C703 diff_3796_1604# gnd! 129.8fF
C704 diff_3745_1604# gnd! 129.8fF
C705 diff_3694_1604# gnd! 129.8fF
C706 diff_3643_1604# gnd! 129.8fF
C707 diff_3592_1604# gnd! 129.8fF
C708 diff_3541_1604# gnd! 129.8fF
C709 diff_3490_1604# gnd! 129.8fF
C710 diff_3439_1604# gnd! 129.8fF
C711 diff_3388_1604# gnd! 129.8fF
C712 diff_3337_1604# gnd! 129.8fF
C713 diff_3286_1604# gnd! 129.8fF
C714 diff_3235_1604# gnd! 129.8fF
C715 diff_3184_1604# gnd! 129.8fF
C716 diff_3133_1604# gnd! 129.8fF
C717 diff_3082_1604# gnd! 129.8fF
C718 diff_3031_1604# gnd! 129.8fF
C719 diff_2980_1604# gnd! 129.8fF
C720 diff_2929_1604# gnd! 129.8fF
C721 diff_2878_1604# gnd! 129.8fF
C722 diff_2827_1604# gnd! 129.8fF
C723 diff_2776_1604# gnd! 129.8fF
C724 diff_2725_1604# gnd! 129.8fF
C725 diff_2674_1604# gnd! 129.8fF
C726 diff_2623_1604# gnd! 129.8fF
C727 diff_2572_1604# gnd! 129.8fF
C728 diff_2521_1604# gnd! 129.8fF
C729 diff_1867_1564# gnd! 1273.0fF
C730 diff_2512_1645# gnd! 3604.0fF
C731 diff_5734_1658# gnd! 137.9fF
C732 diff_5683_1658# gnd! 137.9fF
C733 diff_5632_1658# gnd! 137.9fF
C734 diff_5581_1658# gnd! 137.9fF
C735 diff_5530_1658# gnd! 137.9fF
C736 diff_5479_1658# gnd! 137.9fF
C737 diff_5428_1658# gnd! 137.9fF
C738 diff_5377_1658# gnd! 137.9fF
C739 diff_5326_1658# gnd! 137.9fF
C740 diff_5275_1658# gnd! 137.9fF
C741 diff_5224_1658# gnd! 137.9fF
C742 diff_5173_1658# gnd! 137.9fF
C743 diff_5122_1658# gnd! 137.9fF
C744 diff_5071_1658# gnd! 137.9fF
C745 diff_5020_1658# gnd! 137.9fF
C746 diff_4969_1658# gnd! 137.9fF
C747 diff_4918_1658# gnd! 137.9fF
C748 diff_4867_1658# gnd! 137.9fF
C749 diff_4816_1658# gnd! 137.9fF
C750 diff_4765_1658# gnd! 137.9fF
C751 diff_4714_1658# gnd! 137.9fF
C752 diff_4663_1658# gnd! 137.9fF
C753 diff_4612_1658# gnd! 137.9fF
C754 diff_4561_1658# gnd! 137.9fF
C755 diff_4510_1658# gnd! 137.9fF
C756 diff_4459_1658# gnd! 137.9fF
C757 diff_4408_1658# gnd! 137.9fF
C758 diff_4357_1658# gnd! 137.9fF
C759 diff_4306_1658# gnd! 137.9fF
C760 diff_4255_1658# gnd! 137.9fF
C761 diff_4204_1658# gnd! 137.9fF
C762 diff_4153_1658# gnd! 137.9fF
C763 diff_4102_1658# gnd! 137.9fF
C764 diff_4051_1658# gnd! 137.9fF
C765 diff_4000_1658# gnd! 137.9fF
C766 diff_3949_1658# gnd! 137.9fF
C767 diff_3898_1658# gnd! 137.9fF
C768 diff_3847_1658# gnd! 137.9fF
C769 diff_3796_1658# gnd! 137.9fF
C770 diff_3745_1658# gnd! 137.9fF
C771 diff_3694_1658# gnd! 137.9fF
C772 diff_3643_1658# gnd! 137.9fF
C773 diff_3592_1658# gnd! 137.9fF
C774 diff_3541_1658# gnd! 137.9fF
C775 diff_3490_1658# gnd! 137.9fF
C776 diff_3439_1658# gnd! 137.9fF
C777 diff_3388_1658# gnd! 137.9fF
C778 diff_3337_1658# gnd! 137.9fF
C779 diff_3286_1658# gnd! 137.9fF
C780 diff_3235_1658# gnd! 137.9fF
C781 diff_3184_1658# gnd! 137.9fF
C782 diff_3133_1658# gnd! 137.9fF
C783 diff_3082_1658# gnd! 137.9fF
C784 diff_3031_1658# gnd! 137.9fF
C785 diff_2980_1658# gnd! 137.9fF
C786 diff_2929_1658# gnd! 137.9fF
C787 diff_2878_1658# gnd! 137.9fF
C788 diff_2827_1658# gnd! 137.9fF
C789 diff_2776_1658# gnd! 137.9fF
C790 diff_2725_1658# gnd! 137.9fF
C791 diff_2674_1658# gnd! 137.9fF
C792 diff_2623_1658# gnd! 137.9fF
C793 diff_2572_1658# gnd! 137.9fF
C794 diff_2228_1642# gnd! 56.6fF
C795 diff_2245_1597# gnd! 678.1fF
C796 diff_2521_1658# gnd! 137.9fF
C797 diff_2512_1534# gnd! 3299.3fF
C798 diff_2512_1702# gnd! 3420.2fF
C799 diff_5734_1715# gnd! 129.8fF
C800 diff_5683_1715# gnd! 129.8fF
C801 diff_5632_1715# gnd! 129.8fF
C802 diff_5581_1715# gnd! 129.8fF
C803 diff_5530_1715# gnd! 129.8fF
C804 diff_5479_1715# gnd! 129.8fF
C805 diff_5428_1715# gnd! 129.8fF
C806 diff_5377_1715# gnd! 129.8fF
C807 diff_5326_1715# gnd! 129.8fF
C808 diff_5275_1715# gnd! 129.8fF
C809 diff_5224_1715# gnd! 129.8fF
C810 diff_5173_1715# gnd! 129.8fF
C811 diff_5122_1715# gnd! 129.8fF
C812 diff_5071_1715# gnd! 129.8fF
C813 diff_5020_1715# gnd! 129.8fF
C814 diff_4969_1715# gnd! 129.8fF
C815 diff_4918_1715# gnd! 129.8fF
C816 diff_4867_1715# gnd! 129.8fF
C817 diff_4816_1715# gnd! 129.8fF
C818 diff_4765_1715# gnd! 129.8fF
C819 diff_4714_1715# gnd! 129.8fF
C820 diff_4663_1715# gnd! 129.8fF
C821 diff_4612_1715# gnd! 129.8fF
C822 diff_4561_1715# gnd! 129.8fF
C823 diff_4510_1715# gnd! 129.8fF
C824 diff_4459_1715# gnd! 129.8fF
C825 diff_4408_1715# gnd! 129.8fF
C826 diff_4357_1715# gnd! 129.8fF
C827 diff_4306_1715# gnd! 129.8fF
C828 diff_4255_1715# gnd! 129.8fF
C829 diff_4204_1715# gnd! 129.8fF
C830 diff_4153_1715# gnd! 129.8fF
C831 diff_4102_1715# gnd! 129.8fF
C832 diff_4051_1715# gnd! 129.8fF
C833 diff_4000_1715# gnd! 129.8fF
C834 diff_3949_1715# gnd! 129.8fF
C835 diff_3898_1715# gnd! 129.8fF
C836 diff_3847_1715# gnd! 129.8fF
C837 diff_3796_1715# gnd! 129.8fF
C838 diff_3745_1715# gnd! 129.8fF
C839 diff_3694_1715# gnd! 129.8fF
C840 diff_3643_1715# gnd! 129.8fF
C841 diff_3592_1715# gnd! 129.8fF
C842 diff_3541_1715# gnd! 129.8fF
C843 diff_3490_1715# gnd! 129.8fF
C844 diff_3439_1715# gnd! 129.8fF
C845 diff_3388_1715# gnd! 129.8fF
C846 diff_3337_1715# gnd! 129.8fF
C847 diff_3286_1715# gnd! 129.8fF
C848 diff_3235_1715# gnd! 129.8fF
C849 diff_3184_1715# gnd! 129.8fF
C850 diff_3133_1715# gnd! 129.8fF
C851 diff_3082_1715# gnd! 129.8fF
C852 diff_3031_1715# gnd! 129.8fF
C853 diff_2980_1715# gnd! 129.8fF
C854 diff_2929_1715# gnd! 129.8fF
C855 diff_2878_1715# gnd! 129.8fF
C856 diff_2827_1715# gnd! 129.8fF
C857 diff_2776_1715# gnd! 129.8fF
C858 diff_2725_1715# gnd! 129.8fF
C859 diff_2674_1715# gnd! 129.8fF
C860 diff_2623_1715# gnd! 129.8fF
C861 diff_2572_1715# gnd! 129.8fF
C862 diff_2521_1715# gnd! 129.8fF
C863 diff_5918_1741# gnd! 2761.9fF
C864 diff_5734_1769# gnd! 137.9fF
C865 diff_5683_1769# gnd! 137.9fF
C866 diff_5632_1769# gnd! 137.9fF
C867 diff_5581_1769# gnd! 137.9fF
C868 diff_5530_1769# gnd! 137.9fF
C869 diff_5479_1769# gnd! 137.9fF
C870 diff_5428_1769# gnd! 137.9fF
C871 diff_5377_1769# gnd! 137.9fF
C872 diff_5326_1769# gnd! 137.9fF
C873 diff_5275_1769# gnd! 137.9fF
C874 diff_5224_1769# gnd! 137.9fF
C875 diff_5173_1769# gnd! 137.9fF
C876 diff_5122_1769# gnd! 137.9fF
C877 diff_5071_1769# gnd! 137.9fF
C878 diff_5020_1769# gnd! 137.9fF
C879 diff_4969_1769# gnd! 137.9fF
C880 diff_4918_1769# gnd! 137.9fF
C881 diff_4867_1769# gnd! 137.9fF
C882 diff_4816_1769# gnd! 137.9fF
C883 diff_4765_1769# gnd! 137.9fF
C884 diff_4714_1769# gnd! 137.9fF
C885 diff_4663_1769# gnd! 137.9fF
C886 diff_4612_1769# gnd! 137.9fF
C887 diff_4561_1769# gnd! 137.9fF
C888 diff_4510_1769# gnd! 137.9fF
C889 diff_4459_1769# gnd! 137.9fF
C890 diff_4408_1769# gnd! 137.9fF
C891 diff_4357_1769# gnd! 137.9fF
C892 diff_4306_1769# gnd! 137.9fF
C893 diff_4255_1769# gnd! 137.9fF
C894 diff_4204_1769# gnd! 137.9fF
C895 diff_4153_1769# gnd! 137.9fF
C896 diff_4102_1769# gnd! 137.9fF
C897 diff_4051_1769# gnd! 137.9fF
C898 diff_4000_1769# gnd! 137.9fF
C899 diff_3949_1769# gnd! 137.9fF
C900 diff_3898_1769# gnd! 137.9fF
C901 diff_3847_1769# gnd! 137.9fF
C902 diff_3796_1769# gnd! 137.9fF
C903 diff_3745_1769# gnd! 137.9fF
C904 diff_3694_1769# gnd! 137.9fF
C905 diff_3643_1769# gnd! 137.9fF
C906 diff_3592_1769# gnd! 137.9fF
C907 diff_3541_1769# gnd! 137.9fF
C908 diff_3490_1769# gnd! 137.9fF
C909 diff_3439_1769# gnd! 137.9fF
C910 diff_3388_1769# gnd! 137.9fF
C911 diff_3337_1769# gnd! 137.9fF
C912 diff_3286_1769# gnd! 137.9fF
C913 diff_3235_1769# gnd! 137.9fF
C914 diff_3184_1769# gnd! 137.9fF
C915 diff_3133_1769# gnd! 137.9fF
C916 diff_3082_1769# gnd! 137.9fF
C917 diff_3031_1769# gnd! 137.9fF
C918 diff_2980_1769# gnd! 137.9fF
C919 diff_2929_1769# gnd! 137.9fF
C920 diff_2878_1769# gnd! 137.9fF
C921 diff_2827_1769# gnd! 137.9fF
C922 diff_2776_1769# gnd! 137.9fF
C923 diff_2725_1769# gnd! 137.9fF
C924 diff_2674_1769# gnd! 137.9fF
C925 diff_2623_1769# gnd! 137.9fF
C926 diff_2572_1769# gnd! 137.9fF
C927 diff_2261_1642# gnd! 420.7fF
C928 diff_2521_1769# gnd! 137.9fF
C929 diff_2512_1813# gnd! 3548.7fF
C930 diff_5734_1826# gnd! 129.8fF
C931 diff_5683_1826# gnd! 129.8fF
C932 diff_5632_1826# gnd! 129.8fF
C933 diff_5581_1826# gnd! 129.8fF
C934 diff_5530_1826# gnd! 129.8fF
C935 diff_5479_1826# gnd! 129.8fF
C936 diff_5428_1826# gnd! 129.8fF
C937 diff_5377_1826# gnd! 129.8fF
C938 diff_5326_1826# gnd! 129.8fF
C939 diff_5275_1826# gnd! 129.8fF
C940 diff_5224_1826# gnd! 129.8fF
C941 diff_5173_1826# gnd! 129.8fF
C942 diff_5122_1826# gnd! 129.8fF
C943 diff_5071_1826# gnd! 129.8fF
C944 diff_5020_1826# gnd! 129.8fF
C945 diff_4969_1826# gnd! 129.8fF
C946 diff_4918_1826# gnd! 129.8fF
C947 diff_4867_1826# gnd! 129.8fF
C948 diff_4816_1826# gnd! 129.8fF
C949 diff_4765_1826# gnd! 129.8fF
C950 diff_4714_1826# gnd! 129.8fF
C951 diff_4663_1826# gnd! 129.8fF
C952 diff_4612_1826# gnd! 129.8fF
C953 diff_4561_1826# gnd! 129.8fF
C954 diff_4510_1826# gnd! 129.8fF
C955 diff_4459_1826# gnd! 129.8fF
C956 diff_4408_1826# gnd! 129.8fF
C957 diff_4357_1826# gnd! 129.8fF
C958 diff_4306_1826# gnd! 129.8fF
C959 diff_4255_1826# gnd! 129.8fF
C960 diff_4204_1826# gnd! 129.8fF
C961 diff_4153_1826# gnd! 129.8fF
C962 diff_4102_1826# gnd! 129.8fF
C963 diff_4051_1826# gnd! 129.8fF
C964 diff_4000_1826# gnd! 129.8fF
C965 diff_3949_1826# gnd! 129.8fF
C966 diff_3898_1826# gnd! 129.8fF
C967 diff_3847_1826# gnd! 129.8fF
C968 diff_3796_1826# gnd! 129.8fF
C969 diff_3745_1826# gnd! 129.8fF
C970 diff_3694_1826# gnd! 129.8fF
C971 diff_3643_1826# gnd! 129.8fF
C972 diff_3592_1826# gnd! 129.8fF
C973 diff_3541_1826# gnd! 129.8fF
C974 diff_3490_1826# gnd! 129.8fF
C975 diff_3439_1826# gnd! 129.8fF
C976 diff_3388_1826# gnd! 129.8fF
C977 diff_3337_1826# gnd! 129.8fF
C978 diff_3286_1826# gnd! 129.8fF
C979 diff_3235_1826# gnd! 129.8fF
C980 diff_3184_1826# gnd! 129.8fF
C981 diff_3133_1826# gnd! 129.8fF
C982 diff_3082_1826# gnd! 129.8fF
C983 diff_3031_1826# gnd! 129.8fF
C984 diff_2980_1826# gnd! 129.8fF
C985 diff_2929_1826# gnd! 129.8fF
C986 diff_2878_1826# gnd! 129.8fF
C987 diff_2827_1826# gnd! 129.8fF
C988 diff_2776_1826# gnd! 129.8fF
C989 diff_2725_1826# gnd! 129.8fF
C990 diff_2674_1826# gnd! 129.8fF
C991 diff_2623_1826# gnd! 129.8fF
C992 diff_2572_1826# gnd! 129.8fF
C993 diff_2521_1826# gnd! 129.8fF
C994 diff_2512_1867# gnd! 3604.0fF
C995 diff_5734_1880# gnd! 137.9fF
C996 diff_5683_1880# gnd! 137.9fF
C997 diff_5632_1880# gnd! 137.9fF
C998 diff_5581_1880# gnd! 137.9fF
C999 diff_5530_1880# gnd! 137.9fF
C1000 diff_5479_1880# gnd! 137.9fF
C1001 diff_5428_1880# gnd! 137.9fF
C1002 diff_5377_1880# gnd! 137.9fF
C1003 diff_5326_1880# gnd! 137.9fF
C1004 diff_5275_1880# gnd! 137.9fF
C1005 diff_5224_1880# gnd! 137.9fF
C1006 diff_5173_1880# gnd! 137.9fF
C1007 diff_5122_1880# gnd! 137.9fF
C1008 diff_5071_1880# gnd! 137.9fF
C1009 diff_5020_1880# gnd! 137.9fF
C1010 diff_4969_1880# gnd! 137.9fF
C1011 diff_4918_1880# gnd! 137.9fF
C1012 diff_4867_1880# gnd! 137.9fF
C1013 diff_4816_1880# gnd! 137.9fF
C1014 diff_4765_1880# gnd! 137.9fF
C1015 diff_4714_1880# gnd! 137.9fF
C1016 diff_4663_1880# gnd! 137.9fF
C1017 diff_4612_1880# gnd! 137.9fF
C1018 diff_4561_1880# gnd! 137.9fF
C1019 diff_4510_1880# gnd! 137.9fF
C1020 diff_4459_1880# gnd! 137.9fF
C1021 diff_4408_1880# gnd! 137.9fF
C1022 diff_4357_1880# gnd! 137.9fF
C1023 diff_4306_1880# gnd! 137.9fF
C1024 diff_4255_1880# gnd! 137.9fF
C1025 diff_4204_1880# gnd! 137.9fF
C1026 diff_4153_1880# gnd! 137.9fF
C1027 diff_4102_1880# gnd! 137.9fF
C1028 diff_4051_1880# gnd! 137.9fF
C1029 diff_4000_1880# gnd! 137.9fF
C1030 diff_3949_1880# gnd! 137.9fF
C1031 diff_3898_1880# gnd! 137.9fF
C1032 diff_3847_1880# gnd! 137.9fF
C1033 diff_3796_1880# gnd! 137.9fF
C1034 diff_3745_1880# gnd! 137.9fF
C1035 diff_3694_1880# gnd! 137.9fF
C1036 diff_3643_1880# gnd! 137.9fF
C1037 diff_3592_1880# gnd! 137.9fF
C1038 diff_3541_1880# gnd! 137.9fF
C1039 diff_3490_1880# gnd! 137.9fF
C1040 diff_3439_1880# gnd! 137.9fF
C1041 diff_3388_1880# gnd! 137.9fF
C1042 diff_3337_1880# gnd! 137.9fF
C1043 diff_3286_1880# gnd! 137.9fF
C1044 diff_3235_1880# gnd! 137.9fF
C1045 diff_3184_1880# gnd! 137.9fF
C1046 diff_3133_1880# gnd! 137.9fF
C1047 diff_3082_1880# gnd! 137.9fF
C1048 diff_3031_1880# gnd! 137.9fF
C1049 diff_2980_1880# gnd! 137.9fF
C1050 diff_2929_1880# gnd! 137.9fF
C1051 diff_2878_1880# gnd! 137.9fF
C1052 diff_2827_1880# gnd! 137.9fF
C1053 diff_2776_1880# gnd! 137.9fF
C1054 diff_2725_1880# gnd! 137.9fF
C1055 diff_2674_1880# gnd! 137.9fF
C1056 diff_2623_1880# gnd! 137.9fF
C1057 diff_2572_1880# gnd! 137.9fF
C1058 diff_2521_1880# gnd! 137.9fF
C1059 diff_2165_1729# gnd! 522.8fF
C1060 diff_2101_938# gnd! 1139.8fF
C1061 diff_2512_1756# gnd! 3314.0fF
C1062 diff_6325_2236# gnd! 585.5fF
C1063 diff_6845_2317# gnd! 504.0fF
C1064 diff_6325_2290# gnd! 578.6fF
C1065 diff_7081_2641# gnd! 2106.1fF
C1066 diff_7081_2687# gnd! 444.8fF
C1067 diff_6935_2506# gnd! 1031.1fF
C1068 diff_6845_2413# gnd! 509.0fF
C1069 diff_7163_2812# gnd! 287.9fF
C1070 diff_6935_2602# gnd! 1011.4fF
C1071 diff_6328_2422# gnd! 550.5fF
C1072 diff_6328_2479# gnd! 596.2fF
C1073 diff_6328_2590# gnd! 567.5fF
C1074 diff_6845_2695# gnd! 474.4fF
C1075 diff_6328_2647# gnd! 562.2fF
C1076 diff_6331_2779# gnd! 551.7fF
C1077 diff_6935_2884# gnd! 590.6fF
C1078 diff_6845_2788# gnd! 469.3fF
C1079 diff_6328_2833# gnd! 591.2fF
C1080 diff_7046_2842# gnd! 820.8fF
C1081 diff_7103_3070# gnd! 243.2fF
C1082 diff_6935_2974# gnd! 917.7fF
C1083 diff_7046_3232# gnd! 251.6fF
C1084 diff_6328_2947# gnd! 621.0fF
C1085 diff_6845_3073# gnd! 500.7fF
C1086 diff_6328_3004# gnd! 580.8fF
C1087 diff_2512_1924# gnd! 3420.2fF
C1088 diff_2261_1924# gnd! 676.6fF
C1089 diff_712_1165# gnd! 317.0fF
C1090 diff_847_938# gnd! 2358.1fF
C1091 reset gnd! 5796.5fF
C1092 diff_1199_1537# gnd! 517.8fF
C1093 diff_1246_1787# gnd! 276.5fF
C1094 diff_1738_1906# gnd! 740.4fF
C1095 diff_5734_1937# gnd! 214.1fF
C1096 diff_5683_1937# gnd! 217.4fF
C1097 diff_5530_1937# gnd! 214.1fF
C1098 diff_5479_1937# gnd! 217.4fF
C1099 diff_5326_1937# gnd! 214.1fF
C1100 diff_5275_1937# gnd! 217.4fF
C1101 diff_5122_1937# gnd! 214.1fF
C1102 diff_5071_1937# gnd! 217.4fF
C1103 diff_4918_1937# gnd! 214.1fF
C1104 diff_4867_1937# gnd! 217.4fF
C1105 diff_4714_1937# gnd! 214.1fF
C1106 diff_4663_1937# gnd! 217.4fF
C1107 diff_4510_1937# gnd! 214.1fF
C1108 diff_4459_1937# gnd! 217.4fF
C1109 diff_4306_1937# gnd! 214.1fF
C1110 diff_4255_1937# gnd! 217.4fF
C1111 diff_4102_1937# gnd! 214.1fF
C1112 diff_4051_1937# gnd! 217.4fF
C1113 diff_3898_1937# gnd! 214.1fF
C1114 diff_3847_1937# gnd! 217.4fF
C1115 diff_3694_1937# gnd! 214.1fF
C1116 diff_3643_1937# gnd! 217.4fF
C1117 diff_3490_1937# gnd! 214.1fF
C1118 diff_3439_1937# gnd! 217.4fF
C1119 diff_3286_1937# gnd! 214.1fF
C1120 diff_3235_1937# gnd! 217.4fF
C1121 diff_3082_1937# gnd! 214.1fF
C1122 diff_3031_1937# gnd! 217.4fF
C1123 diff_2878_1937# gnd! 214.1fF
C1124 diff_2827_1937# gnd! 217.4fF
C1125 diff_2674_1937# gnd! 207.6fF
C1126 diff_2623_1937# gnd! 212.3fF
C1127 diff_2039_1969# gnd! 75.2fF
C1128 diff_1741_1957# gnd! 378.9fF
C1129 diff_1751_1699# gnd! 795.0fF
C1130 diff_1738_1391# gnd! 1464.3fF
C1131 diff_2299_1054# gnd! 6704.5fF
C1132 diff_2065_1957# gnd! 912.8fF
C1133 diff_6935_3271# gnd! 652.1fF
C1134 diff_6845_3187# gnd! 491.1fF
C1135 diff_6316_3109# gnd! 775.7fF
C1136 diff_6421_3205# gnd! 472.4fF
C1137 diff_6770_3481# gnd! 191.3fF
C1138 diff_6514_3431# gnd! 500.5fF
C1139 diff_6505_3421# gnd! 519.2fF
C1140 diff_6566_3529# gnd! 469.1fF
C1141 diff_6808_2113# gnd! 1968.5fF
C1142 diff_6919_3643# gnd! 263.9fF
C1143 diff_6473_3661# gnd! 439.2fF
C1144 diff_7033_2836# gnd! 1643.0fF
C1145 diff_6922_3745# gnd! 267.2fF
C1146 diff_6922_3853# gnd! 256.7fF
C1147 diff_5632_1937# gnd! 277.2fF
C1148 diff_5581_1937# gnd! 276.8fF
C1149 diff_5645_2123# gnd! 239.3fF
C1150 diff_5428_1937# gnd! 277.2fF
C1151 diff_5377_1937# gnd! 276.8fF
C1152 diff_5441_2123# gnd! 239.3fF
C1153 diff_5224_1937# gnd! 277.2fF
C1154 diff_5173_1937# gnd! 276.8fF
C1155 diff_5237_2123# gnd! 239.3fF
C1156 diff_5020_1937# gnd! 277.2fF
C1157 diff_4969_1937# gnd! 276.8fF
C1158 diff_5033_2123# gnd! 239.3fF
C1159 diff_4816_1937# gnd! 277.2fF
C1160 diff_4765_1937# gnd! 276.8fF
C1161 diff_4829_2123# gnd! 239.3fF
C1162 diff_4612_1937# gnd! 277.2fF
C1163 diff_4561_1937# gnd! 276.8fF
C1164 diff_4625_2123# gnd! 239.3fF
C1165 diff_4408_1937# gnd! 277.2fF
C1166 diff_4357_1937# gnd! 276.8fF
C1167 diff_4421_2123# gnd! 239.3fF
C1168 diff_4204_1937# gnd! 277.2fF
C1169 diff_4153_1937# gnd! 276.8fF
C1170 diff_4217_2123# gnd! 239.3fF
C1171 diff_4000_1937# gnd! 277.2fF
C1172 diff_3949_1937# gnd! 276.8fF
C1173 diff_4013_2123# gnd! 239.3fF
C1174 diff_3796_1937# gnd! 277.2fF
C1175 diff_3745_1937# gnd! 276.8fF
C1176 diff_3809_2123# gnd! 239.3fF
C1177 diff_3592_1937# gnd! 277.2fF
C1178 diff_3541_1937# gnd! 276.8fF
C1179 diff_3605_2123# gnd! 239.3fF
C1180 diff_3388_1937# gnd! 277.2fF
C1181 diff_3337_1937# gnd! 276.8fF
C1182 diff_3401_2123# gnd! 239.3fF
C1183 diff_3184_1937# gnd! 277.2fF
C1184 diff_3133_1937# gnd! 276.8fF
C1185 diff_3197_2123# gnd! 239.3fF
C1186 diff_2980_1937# gnd! 277.2fF
C1187 diff_2929_1937# gnd! 276.8fF
C1188 diff_2993_2123# gnd! 239.3fF
C1189 diff_2776_1937# gnd! 277.2fF
C1190 diff_2725_1937# gnd! 276.8fF
C1191 diff_2789_2123# gnd! 239.3fF
C1192 diff_1394_1915# gnd! 750.9fF
C1193 diff_1054_1822# gnd! 517.7fF
C1194 diff_1342_1942# gnd! 697.7fF
C1195 diff_850_1331# gnd! 2193.0fF
C1196 diff_1024_1190# gnd! 1153.4fF
C1197 diff_2521_1937# gnd! 249.9fF
C1198 diff_2582_2126# gnd! 266.3fF
C1199 diff_2563_2125# gnd! 288.9fF
C1200 diff_5543_2072# gnd! 589.1fF
C1201 diff_5339_2072# gnd! 618.8fF
C1202 diff_5135_2072# gnd! 602.0fF
C1203 diff_5650_2269# gnd! 665.0fF
C1204 diff_5443_2269# gnd! 692.0fF
C1205 diff_4931_2072# gnd! 618.8fF
C1206 diff_4727_2072# gnd! 602.0fF
C1207 diff_5239_2269# gnd! 680.3fF
C1208 diff_5035_2269# gnd! 692.0fF
C1209 diff_4523_2072# gnd! 620.0fF
C1210 diff_4319_2072# gnd! 602.3fF
C1211 diff_2494_2092# gnd! 557.9fF
C1212 diff_4831_2269# gnd! 680.3fF
C1213 diff_4630_2269# gnd! 692.0fF
C1214 diff_4115_2072# gnd! 596.3fF
C1215 diff_3911_2072# gnd! 578.3fF
C1216 diff_4426_2269# gnd! 680.3fF
C1217 diff_4219_2272# gnd! 668.6fF
C1218 diff_3707_2072# gnd! 594.2fF
C1219 diff_3503_2072# gnd! 578.3fF
C1220 diff_4015_2272# gnd! 656.9fF
C1221 diff_3811_2272# gnd! 668.6fF
C1222 diff_3299_2072# gnd! 636.2fF
C1223 diff_3095_2072# gnd! 615.2fF
C1224 diff_3607_2272# gnd! 656.9fF
C1225 diff_2891_2072# gnd! 618.8fF
C1226 diff_2687_2066# gnd! 605.6fF
C1227 diff_3196_2266# gnd! 703.7fF
C1228 diff_2995_2269# gnd! 692.0fF
C1229 diff_3400_2266# gnd! 716.9fF
C1230 diff_2791_2269# gnd! 681.8fF
C1231 diff_2593_2260# gnd! 675.5fF
C1232 diff_5545_2320# gnd! 606.7fF
C1233 diff_5338_2320# gnd! 617.2fF
C1234 diff_5134_2320# gnd! 613.6fF
C1235 diff_4930_2320# gnd! 617.2fF
C1236 diff_4726_2320# gnd! 613.6fF
C1237 diff_4525_2320# gnd! 617.2fF
C1238 diff_4321_2320# gnd! 613.6fF
C1239 diff_4114_2323# gnd! 593.8fF
C1240 diff_3910_2323# gnd! 590.2fF
C1241 diff_3706_2323# gnd! 593.8fF
C1242 diff_3502_2323# gnd! 590.2fF
C1243 diff_3295_2317# gnd! 640.6fF
C1244 diff_3091_2317# gnd! 637.0fF
C1245 diff_2890_2320# gnd! 617.2fF
C1246 diff_1120_1930# gnd! 420.9fF
C1247 diff_1243_1996# gnd! 738.8fF
C1248 diff_2246_2221# gnd! 613.0fF
C1249 diff_2686_2320# gnd! 613.6fF
C1250 diff_5747_2072# gnd! 727.6fF
C1251 diff_5143_2267# gnd! 1420.5fF
C1252 diff_5554_2267# gnd! 1447.7fF
C1253 diff_4735_2267# gnd! 1423.1fF
C1254 diff_5347_2270# gnd! 1564.2fF
C1255 diff_4330_2267# gnd! 1427.0fF
C1256 diff_4939_2270# gnd! 1555.3fF
C1257 diff_3919_2267# gnd! 1453.1fF
C1258 diff_4534_2270# gnd! 1570.2fF
C1259 diff_3511_2267# gnd! 1445.2fF
C1260 diff_3100_2267# gnd! 1369.8fF
C1261 diff_2695_2267# gnd! 1411.6fF
C1262 diff_2500_2240# gnd! 1717.0fF
C1263 diff_2812_2410# gnd! 4156.6fF
C1264 diff_4123_2270# gnd! 1566.0fF
C1265 diff_3715_2267# gnd! 1589.2fF
C1266 diff_3304_2261# gnd! 1542.2fF
C1267 diff_2899_2270# gnd! 1528.6fF
C1268 diff_2003_2221# gnd! 607.5fF
C1269 diff_1202_2005# gnd! 822.1fF
C1270 diff_2536_2407# gnd! 4547.1fF
C1271 diff_4993_2519# gnd! 1612.3fF
C1272 diff_4177_2519# gnd! 1809.0fF
C1273 diff_1561_1187# gnd! 4731.5fF
C1274 diff_3361_2519# gnd! 1578.3fF
C1275 diff_2500_2719# gnd! 1440.7fF
C1276 diff_1616_2221# gnd! 613.0fF
C1277 diff_1420_2140# gnd! 560.6fF
C1278 diff_1030_2134# gnd! 308.9fF
C1279 diff_1235_2224# gnd! 607.5fF
C1280 diff_2072_2599# gnd! 2151.9fF
C1281 diff_2008_2417# gnd! 681.8fF
C1282 diff_2417_2710# gnd! 597.8fF
C1283 diff_2254_2420# gnd! 992.0fF
C1284 diff_5401_2462# gnd! 2610.2fF
C1285 diff_4993_2459# gnd! 3084.8fF
C1286 diff_1411_1187# gnd! 5455.3fF
C1287 diff_4588_2459# gnd! 2939.6fF
C1288 diff_4177_2459# gnd! 2946.8fF
C1289 diff_3769_2459# gnd! 3188.5fF
C1290 diff_3358_2806# gnd! 3030.7fF
C1291 diff_2953_2462# gnd! 2796.7fF
C1292 diff_1030_2168# gnd! 3706.4fF
C1293 diff_1706_2587# gnd! 2282.0fF
C1294 diff_1621_2417# gnd! 634.1fF
C1295 diff_1358_2545# gnd! 3118.5fF
C1296 diff_1243_2417# gnd! 592.1fF
C1297 io0 gnd! 16366.9fF
C1298 diff_1117_2257# gnd! 2408.4fF
C1299 diff_1018_1732# gnd! 3298.7fF
C1300 io1 gnd! 15856.8fF
C1301 io2 gnd! 14955.2fF
C1302 io3 gnd! 14371.8fF
C1303 diff_2542_2420# gnd! 2948.6fF
C1304 diff_2530_2884# gnd! 4412.0fF
C1305 diff_2008_2719# gnd! 1208.3fF
C1306 diff_2659_2353# gnd! 6340.9fF
C1307 diff_1621_2719# gnd! 1205.9fF
C1308 diff_1234_2719# gnd! 1173.1fF
C1309 diff_844_2719# gnd! 1173.8fF
C1310 diff_2584_2299# gnd! 6851.6fF
C1311 diff_2488_3064# gnd! 7476.2fF
C1312 diff_5554_3016# gnd! 1472.4fF
C1313 diff_5645_3164# gnd! 236.9fF
C1314 diff_5347_3019# gnd! 1596.5fF
C1315 diff_5545_2951# gnd! 565.3fF
C1316 diff_5441_3164# gnd! 236.9fF
C1317 diff_5143_3019# gnd! 1409.8fF
C1318 diff_5338_2951# gnd! 574.0fF
C1319 diff_5237_3164# gnd! 236.9fF
C1320 diff_4939_3019# gnd! 1581.0fF
C1321 diff_5134_2951# gnd! 571.3fF
C1322 diff_5033_3164# gnd! 236.9fF
C1323 diff_4735_3019# gnd! 1409.8fF
C1324 diff_4930_2951# gnd! 574.0fF
C1325 diff_4829_3164# gnd! 236.9fF
C1326 diff_4534_3019# gnd! 1571.5fF
C1327 diff_4726_2951# gnd! 571.3fF
C1328 diff_4625_3164# gnd! 236.9fF
C1329 diff_4330_3019# gnd! 1412.8fF
C1330 diff_4525_2951# gnd! 574.0fF
C1331 diff_4421_3164# gnd! 236.9fF
C1332 diff_4123_3016# gnd! 1584.7fF
C1333 diff_4321_2951# gnd! 571.3fF
C1334 diff_4217_3164# gnd! 236.9fF
C1335 diff_3919_3016# gnd! 1444.9fF
C1336 diff_4114_2951# gnd! 550.6fF
C1337 diff_4013_3164# gnd! 236.9fF
C1338 diff_3715_3016# gnd! 1609.3fF
C1339 diff_3910_2951# gnd! 547.9fF
C1340 diff_3809_3164# gnd! 236.9fF
C1341 diff_3511_3016# gnd! 1444.9fF
C1342 diff_3706_2951# gnd! 550.6fF
C1343 diff_3605_3164# gnd! 236.9fF
C1344 diff_3304_3022# gnd! 1572.7fF
C1345 diff_3502_2951# gnd! 547.9fF
C1346 diff_3401_3164# gnd! 236.9fF
C1347 diff_3100_3022# gnd! 1365.6fF
C1348 diff_3295_2951# gnd! 579.3fF
C1349 diff_3197_3164# gnd! 236.9fF
C1350 diff_2899_3019# gnd! 1545.1fF
C1351 diff_3091_2951# gnd! 594.7fF
C1352 diff_2993_3164# gnd! 236.9fF
C1353 diff_2695_3019# gnd! 1411.6fF
C1354 diff_2890_2951# gnd! 574.0fF
C1355 diff_2789_3164# gnd! 236.9fF
C1356 diff_2500_3043# gnd! 1703.1fF
C1357 diff_2582_3167# gnd! 268.4fF
C1358 diff_2686_2951# gnd! 571.3fF
C1359 diff_2623_2116# gnd! 8781.3fF
C1360 diff_5747_3211# gnd! 695.2fF
C1361 diff_5650_3005# gnd! 635.5fF
C1362 diff_5543_3211# gnd! 549.3fF
C1363 diff_5443_3005# gnd! 662.4fF
C1364 diff_5339_3211# gnd! 583.1fF
C1365 diff_5239_3005# gnd! 649.6fF
C1366 diff_5135_3211# gnd! 561.3fF
C1367 diff_5035_3005# gnd! 662.4fF
C1368 diff_4931_3211# gnd! 583.1fF
C1369 diff_4831_3005# gnd! 649.6fF
C1370 diff_4727_3211# gnd! 561.3fF
C1371 diff_4630_3005# gnd! 662.4fF
C1372 diff_4523_3211# gnd! 584.4fF
C1373 diff_4426_3005# gnd! 649.6fF
C1374 diff_4319_3211# gnd! 561.6fF
C1375 diff_4219_3005# gnd! 639.0fF
C1376 diff_4115_3211# gnd! 560.6fF
C1377 diff_4015_3005# gnd! 626.2fF
C1378 diff_3911_3211# gnd! 537.6fF
C1379 diff_3811_3005# gnd! 639.0fF
C1380 diff_3707_3211# gnd! 556.6fF
C1381 diff_3607_3005# gnd! 626.2fF
C1382 diff_3503_3211# gnd! 537.6fF
C1383 diff_3400_3002# gnd! 687.3fF
C1384 diff_3299_3211# gnd! 601.1fF
C1385 diff_3196_3005# gnd! 673.0fF
C1386 diff_3095_3211# gnd! 574.5fF
C1387 diff_2995_3005# gnd! 662.4fF
C1388 diff_2891_3211# gnd! 585.1fF
C1389 diff_2791_3002# gnd! 651.1fF
C1390 diff_2687_3211# gnd! 564.9fF
C1391 diff_2593_3005# gnd! 646.6fF
C1392 diff_2812_2884# gnd! 4317.3fF
C1393 diff_652_1966# gnd! 3711.4fF
C1394 cl gnd! 9643.8fF
C1395 diff_2494_3091# gnd! 529.4fF
C1396 diff_2053_3250# gnd! 1084.8fF
C1397 diff_2341_3208# gnd! 138.2fF ;**FLOATING
C1398 diff_1666_3250# gnd! 1066.4fF
C1399 diff_2005_2926# gnd! 1683.8fF
C1400 diff_5734_3205# gnd! 222.2fF
C1401 diff_5683_3304# gnd! 225.5fF
C1402 diff_5632_3157# gnd! 285.3fF
C1403 diff_5581_3304# gnd! 284.9fF
C1404 diff_5530_3205# gnd! 222.2fF
C1405 diff_5479_3304# gnd! 225.5fF
C1406 diff_5428_3157# gnd! 285.3fF
C1407 diff_5377_3304# gnd! 284.9fF
C1408 diff_5326_3205# gnd! 222.2fF
C1409 diff_5275_3304# gnd! 225.5fF
C1410 diff_5224_3157# gnd! 285.3fF
C1411 diff_5173_3304# gnd! 284.9fF
C1412 diff_5122_3205# gnd! 222.2fF
C1413 diff_5071_3304# gnd! 225.5fF
C1414 diff_5020_3157# gnd! 285.3fF
C1415 diff_4969_3304# gnd! 284.9fF
C1416 diff_4918_3205# gnd! 222.2fF
C1417 diff_4867_3304# gnd! 225.5fF
C1418 diff_4816_3157# gnd! 285.3fF
C1419 diff_4765_3304# gnd! 284.9fF
C1420 diff_4714_3205# gnd! 222.2fF
C1421 diff_4663_3304# gnd! 225.5fF
C1422 diff_4612_3157# gnd! 285.3fF
C1423 diff_4561_3304# gnd! 284.9fF
C1424 diff_4510_3205# gnd! 222.2fF
C1425 diff_4459_3304# gnd! 225.5fF
C1426 diff_4408_3157# gnd! 285.3fF
C1427 diff_4357_3304# gnd! 284.9fF
C1428 diff_4306_3205# gnd! 222.2fF
C1429 diff_4255_3304# gnd! 225.5fF
C1430 diff_4204_3157# gnd! 285.3fF
C1431 diff_4153_3304# gnd! 284.9fF
C1432 diff_4102_3205# gnd! 222.2fF
C1433 diff_4051_3304# gnd! 225.5fF
C1434 diff_4000_3157# gnd! 285.3fF
C1435 diff_3949_3304# gnd! 284.9fF
C1436 diff_3898_3205# gnd! 222.2fF
C1437 diff_3847_3304# gnd! 225.5fF
C1438 diff_3796_3157# gnd! 285.3fF
C1439 diff_3745_3304# gnd! 284.9fF
C1440 diff_3694_3205# gnd! 222.2fF
C1441 diff_3643_3304# gnd! 225.5fF
C1442 diff_3592_3157# gnd! 285.3fF
C1443 diff_3541_3304# gnd! 284.9fF
C1444 diff_3490_3205# gnd! 222.2fF
C1445 diff_3439_3304# gnd! 225.5fF
C1446 diff_3388_3157# gnd! 285.3fF
C1447 diff_3337_3304# gnd! 284.9fF
C1448 diff_3286_3205# gnd! 222.2fF
C1449 diff_3235_3304# gnd! 225.5fF
C1450 diff_3184_3157# gnd! 285.3fF
C1451 diff_3133_3304# gnd! 284.9fF
C1452 diff_3082_3205# gnd! 222.2fF
C1453 diff_3031_3304# gnd! 225.5fF
C1454 diff_2980_3157# gnd! 285.3fF
C1455 diff_2929_3304# gnd! 284.9fF
C1456 diff_2878_3205# gnd! 222.2fF
C1457 diff_2827_3304# gnd! 225.5fF
C1458 diff_2776_3157# gnd! 285.3fF
C1459 diff_2725_3304# gnd! 284.9fF
C1460 diff_2674_3205# gnd! 215.7fF
C1461 diff_2623_3307# gnd! 220.4fF
C1462 diff_2563_3160# gnd! 297.0fF
C1463 diff_1999_3193# gnd! 1691.5fF
C1464 diff_1273_3250# gnd! 1088.6fF
C1465 diff_1618_2926# gnd! 1743.6fF
C1466 diff_1612_3193# gnd! 1686.0fF
C1467 diff_889_3250# gnd! 1089.4fF
C1468 diff_1231_2926# gnd! 1679.1fF
C1469 diff_1222_3193# gnd! 1645.7fF
C1470 diff_841_2926# gnd! 1687.5fF
C1471 diff_835_3196# gnd! 1678.6fF
C1472 diff_701_3292# gnd! 1535.3fF
C1473 diff_2521_3301# gnd! 263.6fF
C1474 diff_2512_3367# gnd! 3364.9fF
C1475 diff_5734_3380# gnd! 137.9fF
C1476 diff_5683_3380# gnd! 137.9fF
C1477 diff_5632_3380# gnd! 137.9fF
C1478 diff_5581_3380# gnd! 137.9fF
C1479 diff_5530_3380# gnd! 137.9fF
C1480 diff_5479_3380# gnd! 137.9fF
C1481 diff_5428_3380# gnd! 137.9fF
C1482 diff_5377_3380# gnd! 137.9fF
C1483 diff_5326_3380# gnd! 137.9fF
C1484 diff_5275_3380# gnd! 137.9fF
C1485 diff_5224_3380# gnd! 137.9fF
C1486 diff_5173_3380# gnd! 137.9fF
C1487 diff_5122_3380# gnd! 137.9fF
C1488 diff_5071_3380# gnd! 137.9fF
C1489 diff_5020_3380# gnd! 137.9fF
C1490 diff_4969_3380# gnd! 137.9fF
C1491 diff_4918_3380# gnd! 137.9fF
C1492 diff_4867_3380# gnd! 137.9fF
C1493 diff_4816_3380# gnd! 137.9fF
C1494 diff_4765_3380# gnd! 137.9fF
C1495 diff_4714_3380# gnd! 137.9fF
C1496 diff_4663_3380# gnd! 137.9fF
C1497 diff_4612_3380# gnd! 137.9fF
C1498 diff_4561_3380# gnd! 137.9fF
C1499 diff_4510_3380# gnd! 137.9fF
C1500 diff_4459_3380# gnd! 137.9fF
C1501 diff_4408_3380# gnd! 137.9fF
C1502 diff_4357_3380# gnd! 137.9fF
C1503 diff_4306_3380# gnd! 137.9fF
C1504 diff_4255_3380# gnd! 137.9fF
C1505 diff_4204_3380# gnd! 137.9fF
C1506 diff_4153_3380# gnd! 137.9fF
C1507 diff_4102_3380# gnd! 137.9fF
C1508 diff_4051_3380# gnd! 137.9fF
C1509 diff_4000_3380# gnd! 137.9fF
C1510 diff_3949_3380# gnd! 137.9fF
C1511 diff_3898_3380# gnd! 137.9fF
C1512 diff_3847_3380# gnd! 137.9fF
C1513 diff_3796_3380# gnd! 137.9fF
C1514 diff_3745_3380# gnd! 137.9fF
C1515 diff_3694_3380# gnd! 137.9fF
C1516 diff_3643_3380# gnd! 137.9fF
C1517 diff_3592_3380# gnd! 137.9fF
C1518 diff_3541_3380# gnd! 137.9fF
C1519 diff_3490_3380# gnd! 137.9fF
C1520 diff_3439_3380# gnd! 137.9fF
C1521 diff_3388_3380# gnd! 137.9fF
C1522 diff_3337_3380# gnd! 137.9fF
C1523 diff_3286_3380# gnd! 137.9fF
C1524 diff_3235_3380# gnd! 137.9fF
C1525 diff_3184_3380# gnd! 137.9fF
C1526 diff_3133_3380# gnd! 137.9fF
C1527 diff_3082_3380# gnd! 137.9fF
C1528 diff_3031_3380# gnd! 137.9fF
C1529 diff_2980_3380# gnd! 137.9fF
C1530 diff_2929_3380# gnd! 137.9fF
C1531 diff_2878_3380# gnd! 137.9fF
C1532 diff_2827_3380# gnd! 137.9fF
C1533 diff_2776_3380# gnd! 137.9fF
C1534 diff_2725_3380# gnd! 137.9fF
C1535 diff_2674_3380# gnd! 137.9fF
C1536 diff_2623_3380# gnd! 137.9fF
C1537 diff_2572_3380# gnd! 137.9fF
C1538 diff_1999_3365# gnd! 74.6fF
C1539 diff_1612_3365# gnd! 74.6fF
C1540 diff_1222_3365# gnd! 74.6fF
C1541 diff_835_3365# gnd! 74.6fF
C1542 diff_388_2056# gnd! 4204.9fF
C1543 diff_2521_3380# gnd! 137.9fF
C1544 diff_2512_3424# gnd! 3555.5fF
C1545 diff_5734_3437# gnd! 129.8fF
C1546 diff_5683_3437# gnd! 129.8fF
C1547 diff_5632_3437# gnd! 129.8fF
C1548 diff_5581_3437# gnd! 129.8fF
C1549 diff_5530_3437# gnd! 129.8fF
C1550 diff_5479_3437# gnd! 129.8fF
C1551 diff_5428_3437# gnd! 129.8fF
C1552 diff_5377_3437# gnd! 129.8fF
C1553 diff_5326_3437# gnd! 129.8fF
C1554 diff_5275_3437# gnd! 129.8fF
C1555 diff_5224_3437# gnd! 129.8fF
C1556 diff_5173_3437# gnd! 129.8fF
C1557 diff_5122_3437# gnd! 129.8fF
C1558 diff_5071_3437# gnd! 129.8fF
C1559 diff_5020_3437# gnd! 129.8fF
C1560 diff_4969_3437# gnd! 129.8fF
C1561 diff_4918_3437# gnd! 129.8fF
C1562 diff_4867_3437# gnd! 129.8fF
C1563 diff_4816_3437# gnd! 129.8fF
C1564 diff_4765_3437# gnd! 129.8fF
C1565 diff_4714_3437# gnd! 129.8fF
C1566 diff_4663_3437# gnd! 129.8fF
C1567 diff_4612_3437# gnd! 129.8fF
C1568 diff_4561_3437# gnd! 129.8fF
C1569 diff_4510_3437# gnd! 129.8fF
C1570 diff_4459_3437# gnd! 129.8fF
C1571 diff_4408_3437# gnd! 129.8fF
C1572 diff_4357_3437# gnd! 129.8fF
C1573 diff_4306_3437# gnd! 129.8fF
C1574 diff_4255_3437# gnd! 129.8fF
C1575 diff_4204_3437# gnd! 129.8fF
C1576 diff_4153_3437# gnd! 129.8fF
C1577 diff_4102_3437# gnd! 129.8fF
C1578 diff_4051_3437# gnd! 129.8fF
C1579 diff_4000_3437# gnd! 129.8fF
C1580 diff_3949_3437# gnd! 129.8fF
C1581 diff_3898_3437# gnd! 129.8fF
C1582 diff_3847_3437# gnd! 129.8fF
C1583 diff_3796_3437# gnd! 129.8fF
C1584 diff_3745_3437# gnd! 129.8fF
C1585 diff_3694_3437# gnd! 129.8fF
C1586 diff_3643_3437# gnd! 129.8fF
C1587 diff_3592_3437# gnd! 129.8fF
C1588 diff_3541_3437# gnd! 129.8fF
C1589 diff_3490_3437# gnd! 129.8fF
C1590 diff_3439_3437# gnd! 129.8fF
C1591 diff_3388_3437# gnd! 129.8fF
C1592 diff_3337_3437# gnd! 129.8fF
C1593 diff_3286_3437# gnd! 129.8fF
C1594 diff_3235_3437# gnd! 129.8fF
C1595 diff_3184_3437# gnd! 129.8fF
C1596 diff_3133_3437# gnd! 129.8fF
C1597 diff_3082_3437# gnd! 129.8fF
C1598 diff_3031_3437# gnd! 129.8fF
C1599 diff_2980_3437# gnd! 129.8fF
C1600 diff_2929_3437# gnd! 129.8fF
C1601 diff_2878_3437# gnd! 129.8fF
C1602 diff_2827_3437# gnd! 129.8fF
C1603 diff_2776_3437# gnd! 129.8fF
C1604 diff_2725_3437# gnd! 129.8fF
C1605 diff_2674_3437# gnd! 129.8fF
C1606 diff_2623_3437# gnd! 129.8fF
C1607 diff_2572_3437# gnd! 129.8fF
C1608 diff_2521_3437# gnd! 129.8fF
C1609 diff_2512_3478# gnd! 3608.6fF
C1610 diff_5918_3518# gnd! 2880.8fF
C1611 diff_5734_3491# gnd! 137.9fF
C1612 diff_5683_3491# gnd! 137.9fF
C1613 diff_5632_3491# gnd! 137.9fF
C1614 diff_5581_3491# gnd! 137.9fF
C1615 diff_5530_3491# gnd! 137.9fF
C1616 diff_5479_3491# gnd! 137.9fF
C1617 diff_5428_3491# gnd! 137.9fF
C1618 diff_5377_3491# gnd! 137.9fF
C1619 diff_5326_3491# gnd! 137.9fF
C1620 diff_5275_3491# gnd! 137.9fF
C1621 diff_5224_3491# gnd! 137.9fF
C1622 diff_5173_3491# gnd! 137.9fF
C1623 diff_5122_3491# gnd! 137.9fF
C1624 diff_5071_3491# gnd! 137.9fF
C1625 diff_5020_3491# gnd! 137.9fF
C1626 diff_4969_3491# gnd! 137.9fF
C1627 diff_4918_3491# gnd! 137.9fF
C1628 diff_4867_3491# gnd! 137.9fF
C1629 diff_4816_3491# gnd! 137.9fF
C1630 diff_4765_3491# gnd! 137.9fF
C1631 diff_4714_3491# gnd! 137.9fF
C1632 diff_4663_3491# gnd! 137.9fF
C1633 diff_4612_3491# gnd! 137.9fF
C1634 diff_4561_3491# gnd! 137.9fF
C1635 diff_4510_3491# gnd! 137.9fF
C1636 diff_4459_3491# gnd! 137.9fF
C1637 diff_4408_3491# gnd! 137.9fF
C1638 diff_4357_3491# gnd! 137.9fF
C1639 diff_4306_3491# gnd! 137.9fF
C1640 diff_4255_3491# gnd! 137.9fF
C1641 diff_4204_3491# gnd! 137.9fF
C1642 diff_4153_3491# gnd! 137.9fF
C1643 diff_4102_3491# gnd! 137.9fF
C1644 diff_4051_3491# gnd! 137.9fF
C1645 diff_4000_3491# gnd! 137.9fF
C1646 diff_3949_3491# gnd! 137.9fF
C1647 diff_3898_3491# gnd! 137.9fF
C1648 diff_3847_3491# gnd! 137.9fF
C1649 diff_3796_3491# gnd! 137.9fF
C1650 diff_3745_3491# gnd! 137.9fF
C1651 diff_3694_3491# gnd! 137.9fF
C1652 diff_3643_3491# gnd! 137.9fF
C1653 diff_3592_3491# gnd! 137.9fF
C1654 diff_3541_3491# gnd! 137.9fF
C1655 diff_3490_3491# gnd! 137.9fF
C1656 diff_3439_3491# gnd! 137.9fF
C1657 diff_3388_3491# gnd! 137.9fF
C1658 diff_3337_3491# gnd! 137.9fF
C1659 diff_3286_3491# gnd! 137.9fF
C1660 diff_3235_3491# gnd! 137.9fF
C1661 diff_3184_3491# gnd! 137.9fF
C1662 diff_3133_3491# gnd! 137.9fF
C1663 diff_3082_3491# gnd! 137.9fF
C1664 diff_3031_3491# gnd! 137.9fF
C1665 diff_2980_3491# gnd! 137.9fF
C1666 diff_2929_3491# gnd! 137.9fF
C1667 diff_2878_3491# gnd! 137.9fF
C1668 diff_2827_3491# gnd! 137.9fF
C1669 diff_2776_3491# gnd! 137.9fF
C1670 diff_2725_3491# gnd! 137.9fF
C1671 diff_2674_3491# gnd! 137.9fF
C1672 diff_2623_3491# gnd! 137.9fF
C1673 diff_2572_3491# gnd! 137.9fF
C1674 diff_2521_3491# gnd! 137.9fF
C1675 diff_2512_3535# gnd! 3369.2fF
C1676 diff_5734_3548# gnd! 129.8fF
C1677 diff_5683_3548# gnd! 129.8fF
C1678 diff_5632_3548# gnd! 129.8fF
C1679 diff_5581_3548# gnd! 129.8fF
C1680 diff_5530_3548# gnd! 129.8fF
C1681 diff_5479_3548# gnd! 129.8fF
C1682 diff_5428_3548# gnd! 129.8fF
C1683 diff_5377_3548# gnd! 129.8fF
C1684 diff_5326_3548# gnd! 129.8fF
C1685 diff_5275_3548# gnd! 129.8fF
C1686 diff_5224_3548# gnd! 129.8fF
C1687 diff_5173_3548# gnd! 129.8fF
C1688 diff_5122_3548# gnd! 129.8fF
C1689 diff_5071_3548# gnd! 129.8fF
C1690 diff_5020_3548# gnd! 129.8fF
C1691 diff_4969_3548# gnd! 129.8fF
C1692 diff_4918_3548# gnd! 129.8fF
C1693 diff_4867_3548# gnd! 129.8fF
C1694 diff_4816_3548# gnd! 129.8fF
C1695 diff_4765_3548# gnd! 129.8fF
C1696 diff_4714_3548# gnd! 129.8fF
C1697 diff_4663_3548# gnd! 129.8fF
C1698 diff_4612_3548# gnd! 129.8fF
C1699 diff_4561_3548# gnd! 129.8fF
C1700 diff_4510_3548# gnd! 129.8fF
C1701 diff_4459_3548# gnd! 129.8fF
C1702 diff_4408_3548# gnd! 129.8fF
C1703 diff_4357_3548# gnd! 129.8fF
C1704 diff_4306_3548# gnd! 129.8fF
C1705 diff_4255_3548# gnd! 129.8fF
C1706 diff_4204_3548# gnd! 129.8fF
C1707 diff_4153_3548# gnd! 129.8fF
C1708 diff_4102_3548# gnd! 129.8fF
C1709 diff_4051_3548# gnd! 129.8fF
C1710 diff_4000_3548# gnd! 129.8fF
C1711 diff_3949_3548# gnd! 129.8fF
C1712 diff_3898_3548# gnd! 129.8fF
C1713 diff_3847_3548# gnd! 129.8fF
C1714 diff_3796_3548# gnd! 129.8fF
C1715 diff_3745_3548# gnd! 129.8fF
C1716 diff_3694_3548# gnd! 129.8fF
C1717 diff_3643_3548# gnd! 129.8fF
C1718 diff_3592_3548# gnd! 129.8fF
C1719 diff_3541_3548# gnd! 129.8fF
C1720 diff_3490_3548# gnd! 129.8fF
C1721 diff_3439_3548# gnd! 129.8fF
C1722 diff_3388_3548# gnd! 129.8fF
C1723 diff_3337_3548# gnd! 129.8fF
C1724 diff_3286_3548# gnd! 129.8fF
C1725 diff_3235_3548# gnd! 129.8fF
C1726 diff_3184_3548# gnd! 129.8fF
C1727 diff_3133_3548# gnd! 129.8fF
C1728 diff_3082_3548# gnd! 129.8fF
C1729 diff_3031_3548# gnd! 129.8fF
C1730 diff_2980_3548# gnd! 129.8fF
C1731 diff_2929_3548# gnd! 129.8fF
C1732 diff_2878_3548# gnd! 129.8fF
C1733 diff_2827_3548# gnd! 129.8fF
C1734 diff_2776_3548# gnd! 129.8fF
C1735 diff_2725_3548# gnd! 129.8fF
C1736 diff_2674_3548# gnd! 129.8fF
C1737 diff_2623_3548# gnd! 129.8fF
C1738 diff_2572_3548# gnd! 129.8fF
C1739 diff_2521_3548# gnd! 129.8fF
C1740 diff_2512_3589# gnd! 3368.9fF
C1741 diff_5734_3602# gnd! 137.9fF
C1742 diff_5683_3602# gnd! 137.9fF
C1743 diff_5632_3602# gnd! 137.9fF
C1744 diff_5581_3602# gnd! 137.9fF
C1745 diff_5530_3602# gnd! 137.9fF
C1746 diff_5479_3602# gnd! 137.9fF
C1747 diff_5428_3602# gnd! 137.9fF
C1748 diff_5377_3602# gnd! 137.9fF
C1749 diff_5326_3602# gnd! 137.9fF
C1750 diff_5275_3602# gnd! 137.9fF
C1751 diff_5224_3602# gnd! 137.9fF
C1752 diff_5173_3602# gnd! 137.9fF
C1753 diff_5122_3602# gnd! 137.9fF
C1754 diff_5071_3602# gnd! 137.9fF
C1755 diff_5020_3602# gnd! 137.9fF
C1756 diff_4969_3602# gnd! 137.9fF
C1757 diff_4918_3602# gnd! 137.9fF
C1758 diff_4867_3602# gnd! 137.9fF
C1759 diff_4816_3602# gnd! 137.9fF
C1760 diff_4765_3602# gnd! 137.9fF
C1761 diff_4714_3602# gnd! 137.9fF
C1762 diff_4663_3602# gnd! 137.9fF
C1763 diff_4612_3602# gnd! 137.9fF
C1764 diff_4561_3602# gnd! 137.9fF
C1765 diff_4510_3602# gnd! 137.9fF
C1766 diff_4459_3602# gnd! 137.9fF
C1767 diff_4408_3602# gnd! 137.9fF
C1768 diff_4357_3602# gnd! 137.9fF
C1769 diff_4306_3602# gnd! 137.9fF
C1770 diff_4255_3602# gnd! 137.9fF
C1771 diff_4204_3602# gnd! 137.9fF
C1772 diff_4153_3602# gnd! 137.9fF
C1773 diff_4102_3602# gnd! 137.9fF
C1774 diff_4051_3602# gnd! 137.9fF
C1775 diff_4000_3602# gnd! 137.9fF
C1776 diff_3949_3602# gnd! 137.9fF
C1777 diff_3898_3602# gnd! 137.9fF
C1778 diff_3847_3602# gnd! 137.9fF
C1779 diff_3796_3602# gnd! 137.9fF
C1780 diff_3745_3602# gnd! 137.9fF
C1781 diff_3694_3602# gnd! 137.9fF
C1782 diff_3643_3602# gnd! 137.9fF
C1783 diff_3592_3602# gnd! 137.9fF
C1784 diff_3541_3602# gnd! 137.9fF
C1785 diff_3490_3602# gnd! 137.9fF
C1786 diff_3439_3602# gnd! 137.9fF
C1787 diff_3388_3602# gnd! 137.9fF
C1788 diff_3337_3602# gnd! 137.9fF
C1789 diff_3286_3602# gnd! 137.9fF
C1790 diff_3235_3602# gnd! 137.9fF
C1791 diff_3184_3602# gnd! 137.9fF
C1792 diff_3133_3602# gnd! 137.9fF
C1793 diff_3082_3602# gnd! 137.9fF
C1794 diff_3031_3602# gnd! 137.9fF
C1795 diff_2980_3602# gnd! 137.9fF
C1796 diff_2929_3602# gnd! 137.9fF
C1797 diff_2878_3602# gnd! 137.9fF
C1798 diff_2827_3602# gnd! 137.9fF
C1799 diff_2776_3602# gnd! 137.9fF
C1800 diff_2725_3602# gnd! 137.9fF
C1801 diff_2674_3602# gnd! 137.9fF
C1802 diff_2623_3602# gnd! 137.9fF
C1803 diff_2572_3602# gnd! 137.9fF
C1804 diff_2521_3602# gnd! 137.9fF
C1805 diff_2512_3646# gnd! 3562.6fF
C1806 diff_5734_3659# gnd! 129.8fF
C1807 diff_5683_3659# gnd! 129.8fF
C1808 diff_5632_3659# gnd! 129.8fF
C1809 diff_5581_3659# gnd! 129.8fF
C1810 diff_5530_3659# gnd! 129.8fF
C1811 diff_5479_3659# gnd! 129.8fF
C1812 diff_5428_3659# gnd! 129.8fF
C1813 diff_5377_3659# gnd! 129.8fF
C1814 diff_5326_3659# gnd! 129.8fF
C1815 diff_5275_3659# gnd! 129.8fF
C1816 diff_5224_3659# gnd! 129.8fF
C1817 diff_5173_3659# gnd! 129.8fF
C1818 diff_5122_3659# gnd! 129.8fF
C1819 diff_5071_3659# gnd! 129.8fF
C1820 diff_5020_3659# gnd! 129.8fF
C1821 diff_4969_3659# gnd! 129.8fF
C1822 diff_4918_3659# gnd! 129.8fF
C1823 diff_4867_3659# gnd! 129.8fF
C1824 diff_4816_3659# gnd! 129.8fF
C1825 diff_4765_3659# gnd! 129.8fF
C1826 diff_4714_3659# gnd! 129.8fF
C1827 diff_4663_3659# gnd! 129.8fF
C1828 diff_4612_3659# gnd! 129.8fF
C1829 diff_4561_3659# gnd! 129.8fF
C1830 diff_4510_3659# gnd! 129.8fF
C1831 diff_4459_3659# gnd! 129.8fF
C1832 diff_4408_3659# gnd! 129.8fF
C1833 diff_4357_3659# gnd! 129.8fF
C1834 diff_4306_3659# gnd! 129.8fF
C1835 diff_4255_3659# gnd! 129.8fF
C1836 diff_4204_3659# gnd! 129.8fF
C1837 diff_4153_3659# gnd! 129.8fF
C1838 diff_4102_3659# gnd! 129.8fF
C1839 diff_4051_3659# gnd! 129.8fF
C1840 diff_4000_3659# gnd! 129.8fF
C1841 diff_3949_3659# gnd! 129.8fF
C1842 diff_3898_3659# gnd! 129.8fF
C1843 diff_3847_3659# gnd! 129.8fF
C1844 diff_3796_3659# gnd! 129.8fF
C1845 diff_3745_3659# gnd! 129.8fF
C1846 diff_3694_3659# gnd! 129.8fF
C1847 diff_3643_3659# gnd! 129.8fF
C1848 diff_3592_3659# gnd! 129.8fF
C1849 diff_3541_3659# gnd! 129.8fF
C1850 diff_3490_3659# gnd! 129.8fF
C1851 diff_3439_3659# gnd! 129.8fF
C1852 diff_3388_3659# gnd! 129.8fF
C1853 diff_3337_3659# gnd! 129.8fF
C1854 diff_3286_3659# gnd! 129.8fF
C1855 diff_3235_3659# gnd! 129.8fF
C1856 diff_3184_3659# gnd! 129.8fF
C1857 diff_3133_3659# gnd! 129.8fF
C1858 diff_3082_3659# gnd! 129.8fF
C1859 diff_3031_3659# gnd! 129.8fF
C1860 diff_2980_3659# gnd! 129.8fF
C1861 diff_2929_3659# gnd! 129.8fF
C1862 diff_2878_3659# gnd! 129.8fF
C1863 diff_2827_3659# gnd! 129.8fF
C1864 diff_2776_3659# gnd! 129.8fF
C1865 diff_2725_3659# gnd! 129.8fF
C1866 diff_2674_3659# gnd! 129.8fF
C1867 diff_2623_3659# gnd! 129.8fF
C1868 diff_2572_3659# gnd! 129.8fF
C1869 diff_2521_3659# gnd! 129.8fF
C1870 diff_2512_3700# gnd! 3612.3fF
C1871 diff_6130_2449# gnd! 3489.4fF
C1872 diff_6175_2281# gnd! 3568.3fF
C1873 diff_6479_3832# gnd! 438.8fF
C1874 diff_7033_2509# gnd! 3700.5fF
C1875 diff_6919_3958# gnd! 286.4fF
C1876 diff_6778_3391# gnd! 2894.5fF
C1877 diff_7072_3184# gnd! 1705.9fF
C1878 diff_7072_2716# gnd! 3180.7fF
C1879 diff_6706_4228# gnd! 286.1fF
C1880 diff_6625_3799# gnd! 2109.7fF
C1881 diff_6859_4258# gnd! 314.6fF
C1882 diff_6661_3556# gnd! 1796.4fF
C1883 diff_6859_4286# gnd! 285.2fF
C1884 diff_6661_4216# gnd! 811.7fF
C1885 diff_5918_3734# gnd! 3054.9fF
C1886 diff_5734_3713# gnd! 137.9fF
C1887 diff_5683_3713# gnd! 137.9fF
C1888 diff_5632_3713# gnd! 137.9fF
C1889 diff_5581_3713# gnd! 137.9fF
C1890 diff_5530_3713# gnd! 137.9fF
C1891 diff_5479_3713# gnd! 137.9fF
C1892 diff_5428_3713# gnd! 137.9fF
C1893 diff_5377_3713# gnd! 137.9fF
C1894 diff_5326_3713# gnd! 137.9fF
C1895 diff_5275_3713# gnd! 137.9fF
C1896 diff_5224_3713# gnd! 137.9fF
C1897 diff_5173_3713# gnd! 137.9fF
C1898 diff_5122_3713# gnd! 137.9fF
C1899 diff_5071_3713# gnd! 137.9fF
C1900 diff_5020_3713# gnd! 137.9fF
C1901 diff_4969_3713# gnd! 137.9fF
C1902 diff_4918_3713# gnd! 137.9fF
C1903 diff_4867_3713# gnd! 137.9fF
C1904 diff_4816_3713# gnd! 137.9fF
C1905 diff_4765_3713# gnd! 137.9fF
C1906 diff_4714_3713# gnd! 137.9fF
C1907 diff_4663_3713# gnd! 137.9fF
C1908 diff_4612_3713# gnd! 137.9fF
C1909 diff_4561_3713# gnd! 137.9fF
C1910 diff_4510_3713# gnd! 137.9fF
C1911 diff_4459_3713# gnd! 137.9fF
C1912 diff_4408_3713# gnd! 137.9fF
C1913 diff_4357_3713# gnd! 137.9fF
C1914 diff_4306_3713# gnd! 137.9fF
C1915 diff_4255_3713# gnd! 137.9fF
C1916 diff_4204_3713# gnd! 137.9fF
C1917 diff_4153_3713# gnd! 137.9fF
C1918 diff_4102_3713# gnd! 137.9fF
C1919 diff_4051_3713# gnd! 137.9fF
C1920 diff_4000_3713# gnd! 137.9fF
C1921 diff_3949_3713# gnd! 137.9fF
C1922 diff_3898_3713# gnd! 137.9fF
C1923 diff_3847_3713# gnd! 137.9fF
C1924 diff_3796_3713# gnd! 137.9fF
C1925 diff_3745_3713# gnd! 137.9fF
C1926 diff_3694_3713# gnd! 137.9fF
C1927 diff_3643_3713# gnd! 137.9fF
C1928 diff_3592_3713# gnd! 137.9fF
C1929 diff_3541_3713# gnd! 137.9fF
C1930 diff_3490_3713# gnd! 137.9fF
C1931 diff_3439_3713# gnd! 137.9fF
C1932 diff_3388_3713# gnd! 137.9fF
C1933 diff_3337_3713# gnd! 137.9fF
C1934 diff_3286_3713# gnd! 137.9fF
C1935 diff_3235_3713# gnd! 137.9fF
C1936 diff_3184_3713# gnd! 137.9fF
C1937 diff_3133_3713# gnd! 137.9fF
C1938 diff_3082_3713# gnd! 137.9fF
C1939 diff_3031_3713# gnd! 137.9fF
C1940 diff_2980_3713# gnd! 137.9fF
C1941 diff_2929_3713# gnd! 137.9fF
C1942 diff_2878_3713# gnd! 137.9fF
C1943 diff_2827_3713# gnd! 137.9fF
C1944 diff_2776_3713# gnd! 137.9fF
C1945 diff_2725_3713# gnd! 137.9fF
C1946 diff_2674_3713# gnd! 137.9fF
C1947 diff_2623_3713# gnd! 137.9fF
C1948 diff_2572_3713# gnd! 137.9fF
C1949 diff_2185_3622# gnd! 1306.1fF
C1950 diff_2521_3713# gnd! 137.9fF
C1951 diff_1798_3622# gnd! 1671.9fF
C1952 diff_2512_3757# gnd! 3354.4fF
C1953 diff_5734_3770# gnd! 129.8fF
C1954 diff_5683_3770# gnd! 129.8fF
C1955 diff_5632_3770# gnd! 129.8fF
C1956 diff_5581_3770# gnd! 129.8fF
C1957 diff_5530_3770# gnd! 129.8fF
C1958 diff_5479_3770# gnd! 129.8fF
C1959 diff_5428_3770# gnd! 129.8fF
C1960 diff_5377_3770# gnd! 129.8fF
C1961 diff_5326_3770# gnd! 129.8fF
C1962 diff_5275_3770# gnd! 129.8fF
C1963 diff_5224_3770# gnd! 129.8fF
C1964 diff_5173_3770# gnd! 129.8fF
C1965 diff_5122_3770# gnd! 129.8fF
C1966 diff_5071_3770# gnd! 129.8fF
C1967 diff_5020_3770# gnd! 129.8fF
C1968 diff_4969_3770# gnd! 129.8fF
C1969 diff_4918_3770# gnd! 129.8fF
C1970 diff_4867_3770# gnd! 129.8fF
C1971 diff_4816_3770# gnd! 129.8fF
C1972 diff_4765_3770# gnd! 129.8fF
C1973 diff_4714_3770# gnd! 129.8fF
C1974 diff_4663_3770# gnd! 129.8fF
C1975 diff_4612_3770# gnd! 129.8fF
C1976 diff_4561_3770# gnd! 129.8fF
C1977 diff_4510_3770# gnd! 129.8fF
C1978 diff_4459_3770# gnd! 129.8fF
C1979 diff_4408_3770# gnd! 129.8fF
C1980 diff_4357_3770# gnd! 129.8fF
C1981 diff_4306_3770# gnd! 129.8fF
C1982 diff_4255_3770# gnd! 129.8fF
C1983 diff_4204_3770# gnd! 129.8fF
C1984 diff_4153_3770# gnd! 129.8fF
C1985 diff_4102_3770# gnd! 129.8fF
C1986 diff_4051_3770# gnd! 129.8fF
C1987 diff_4000_3770# gnd! 129.8fF
C1988 diff_3949_3770# gnd! 129.8fF
C1989 diff_3898_3770# gnd! 129.8fF
C1990 diff_3847_3770# gnd! 129.8fF
C1991 diff_3796_3770# gnd! 129.8fF
C1992 diff_3745_3770# gnd! 129.8fF
C1993 diff_3694_3770# gnd! 129.8fF
C1994 diff_3643_3770# gnd! 129.8fF
C1995 diff_3592_3770# gnd! 129.8fF
C1996 diff_3541_3770# gnd! 129.8fF
C1997 diff_3490_3770# gnd! 129.8fF
C1998 diff_3439_3770# gnd! 129.8fF
C1999 diff_3388_3770# gnd! 129.8fF
C2000 diff_3337_3770# gnd! 129.8fF
C2001 diff_3286_3770# gnd! 129.8fF
C2002 diff_3235_3770# gnd! 129.8fF
C2003 diff_3184_3770# gnd! 129.8fF
C2004 diff_3133_3770# gnd! 129.8fF
C2005 diff_3082_3770# gnd! 129.8fF
C2006 diff_3031_3770# gnd! 129.8fF
C2007 diff_2980_3770# gnd! 129.8fF
C2008 diff_2929_3770# gnd! 129.8fF
C2009 diff_2878_3770# gnd! 129.8fF
C2010 diff_2827_3770# gnd! 129.8fF
C2011 diff_2776_3770# gnd! 129.8fF
C2012 diff_2725_3770# gnd! 129.8fF
C2013 diff_2674_3770# gnd! 129.8fF
C2014 diff_2623_3770# gnd! 129.8fF
C2015 diff_2572_3770# gnd! 129.8fF
C2016 diff_2521_3770# gnd! 129.8fF
C2017 diff_2512_3811# gnd! 3370.3fF
C2018 diff_5734_3824# gnd! 137.9fF
C2019 diff_5683_3824# gnd! 137.9fF
C2020 diff_5632_3824# gnd! 137.9fF
C2021 diff_5581_3824# gnd! 137.9fF
C2022 diff_5530_3824# gnd! 137.9fF
C2023 diff_5479_3824# gnd! 137.9fF
C2024 diff_5428_3824# gnd! 137.9fF
C2025 diff_5377_3824# gnd! 137.9fF
C2026 diff_5326_3824# gnd! 137.9fF
C2027 diff_5275_3824# gnd! 137.9fF
C2028 diff_5224_3824# gnd! 137.9fF
C2029 diff_5173_3824# gnd! 137.9fF
C2030 diff_5122_3824# gnd! 137.9fF
C2031 diff_5071_3824# gnd! 137.9fF
C2032 diff_5020_3824# gnd! 137.9fF
C2033 diff_4969_3824# gnd! 137.9fF
C2034 diff_4918_3824# gnd! 137.9fF
C2035 diff_4867_3824# gnd! 137.9fF
C2036 diff_4816_3824# gnd! 137.9fF
C2037 diff_4765_3824# gnd! 137.9fF
C2038 diff_4714_3824# gnd! 137.9fF
C2039 diff_4663_3824# gnd! 137.9fF
C2040 diff_4612_3824# gnd! 137.9fF
C2041 diff_4561_3824# gnd! 137.9fF
C2042 diff_4510_3824# gnd! 137.9fF
C2043 diff_4459_3824# gnd! 137.9fF
C2044 diff_4408_3824# gnd! 137.9fF
C2045 diff_4357_3824# gnd! 137.9fF
C2046 diff_4306_3824# gnd! 137.9fF
C2047 diff_4255_3824# gnd! 137.9fF
C2048 diff_4204_3824# gnd! 137.9fF
C2049 diff_4153_3824# gnd! 137.9fF
C2050 diff_4102_3824# gnd! 137.9fF
C2051 diff_4051_3824# gnd! 137.9fF
C2052 diff_4000_3824# gnd! 137.9fF
C2053 diff_3949_3824# gnd! 137.9fF
C2054 diff_3898_3824# gnd! 137.9fF
C2055 diff_3847_3824# gnd! 137.9fF
C2056 diff_3796_3824# gnd! 137.9fF
C2057 diff_3745_3824# gnd! 137.9fF
C2058 diff_3694_3824# gnd! 137.9fF
C2059 diff_3643_3824# gnd! 137.9fF
C2060 diff_3592_3824# gnd! 137.9fF
C2061 diff_3541_3824# gnd! 137.9fF
C2062 diff_3490_3824# gnd! 137.9fF
C2063 diff_3439_3824# gnd! 137.9fF
C2064 diff_3388_3824# gnd! 137.9fF
C2065 diff_3337_3824# gnd! 137.9fF
C2066 diff_3286_3824# gnd! 137.9fF
C2067 diff_3235_3824# gnd! 137.9fF
C2068 diff_3184_3824# gnd! 137.9fF
C2069 diff_3133_3824# gnd! 137.9fF
C2070 diff_3082_3824# gnd! 137.9fF
C2071 diff_3031_3824# gnd! 137.9fF
C2072 diff_2980_3824# gnd! 137.9fF
C2073 diff_2929_3824# gnd! 137.9fF
C2074 diff_2878_3824# gnd! 137.9fF
C2075 diff_2827_3824# gnd! 137.9fF
C2076 diff_2776_3824# gnd! 137.9fF
C2077 diff_2725_3824# gnd! 137.9fF
C2078 diff_2674_3824# gnd! 137.9fF
C2079 diff_2623_3824# gnd! 137.9fF
C2080 diff_2572_3824# gnd! 137.9fF
C2081 diff_2521_3824# gnd! 137.9fF
C2082 diff_2512_3868# gnd! 3558.9fF
C2083 diff_5734_3881# gnd! 129.8fF
C2084 diff_5683_3881# gnd! 129.8fF
C2085 diff_5632_3881# gnd! 129.8fF
C2086 diff_5581_3881# gnd! 129.8fF
C2087 diff_5530_3881# gnd! 129.8fF
C2088 diff_5479_3881# gnd! 129.8fF
C2089 diff_5428_3881# gnd! 129.8fF
C2090 diff_5377_3881# gnd! 129.8fF
C2091 diff_5326_3881# gnd! 129.8fF
C2092 diff_5275_3881# gnd! 129.8fF
C2093 diff_5224_3881# gnd! 129.8fF
C2094 diff_5173_3881# gnd! 129.8fF
C2095 diff_5122_3881# gnd! 129.8fF
C2096 diff_5071_3881# gnd! 129.8fF
C2097 diff_5020_3881# gnd! 129.8fF
C2098 diff_4969_3881# gnd! 129.8fF
C2099 diff_4918_3881# gnd! 129.8fF
C2100 diff_4867_3881# gnd! 129.8fF
C2101 diff_4816_3881# gnd! 129.8fF
C2102 diff_4765_3881# gnd! 129.8fF
C2103 diff_4714_3881# gnd! 129.8fF
C2104 diff_4663_3881# gnd! 129.8fF
C2105 diff_4612_3881# gnd! 129.8fF
C2106 diff_4561_3881# gnd! 129.8fF
C2107 diff_4510_3881# gnd! 129.8fF
C2108 diff_4459_3881# gnd! 129.8fF
C2109 diff_4408_3881# gnd! 129.8fF
C2110 diff_4357_3881# gnd! 129.8fF
C2111 diff_4306_3881# gnd! 129.8fF
C2112 diff_4255_3881# gnd! 129.8fF
C2113 diff_4204_3881# gnd! 129.8fF
C2114 diff_4153_3881# gnd! 129.8fF
C2115 diff_4102_3881# gnd! 129.8fF
C2116 diff_4051_3881# gnd! 129.8fF
C2117 diff_4000_3881# gnd! 129.8fF
C2118 diff_3949_3881# gnd! 129.8fF
C2119 diff_3898_3881# gnd! 129.8fF
C2120 diff_3847_3881# gnd! 129.8fF
C2121 diff_3796_3881# gnd! 129.8fF
C2122 diff_3745_3881# gnd! 129.8fF
C2123 diff_3694_3881# gnd! 129.8fF
C2124 diff_3643_3881# gnd! 129.8fF
C2125 diff_3592_3881# gnd! 129.8fF
C2126 diff_3541_3881# gnd! 129.8fF
C2127 diff_3490_3881# gnd! 129.8fF
C2128 diff_3439_3881# gnd! 129.8fF
C2129 diff_3388_3881# gnd! 129.8fF
C2130 diff_3337_3881# gnd! 129.8fF
C2131 diff_3286_3881# gnd! 129.8fF
C2132 diff_3235_3881# gnd! 129.8fF
C2133 diff_3184_3881# gnd! 129.8fF
C2134 diff_3133_3881# gnd! 129.8fF
C2135 diff_3082_3881# gnd! 129.8fF
C2136 diff_3031_3881# gnd! 129.8fF
C2137 diff_2980_3881# gnd! 129.8fF
C2138 diff_2929_3881# gnd! 129.8fF
C2139 diff_2878_3881# gnd! 129.8fF
C2140 diff_2827_3881# gnd! 129.8fF
C2141 diff_2776_3881# gnd! 129.8fF
C2142 diff_2725_3881# gnd! 129.8fF
C2143 diff_2674_3881# gnd! 129.8fF
C2144 diff_2623_3881# gnd! 129.8fF
C2145 diff_2572_3881# gnd! 129.8fF
C2146 diff_2521_3881# gnd! 129.8fF
C2147 diff_1408_3622# gnd! 1748.7fF
C2148 diff_1021_3622# gnd! 1905.9fF
C2149 diff_2512_3922# gnd! 3591.9fF
C2150 diff_5918_3962# gnd! 2908.3fF
C2151 diff_5734_3935# gnd! 137.9fF
C2152 diff_5683_3935# gnd! 137.9fF
C2153 diff_5632_3935# gnd! 137.9fF
C2154 diff_5581_3935# gnd! 137.9fF
C2155 diff_5530_3935# gnd! 137.9fF
C2156 diff_5479_3935# gnd! 137.9fF
C2157 diff_5428_3935# gnd! 137.9fF
C2158 diff_5377_3935# gnd! 137.9fF
C2159 diff_5326_3935# gnd! 137.9fF
C2160 diff_5275_3935# gnd! 137.9fF
C2161 diff_5224_3935# gnd! 137.9fF
C2162 diff_5173_3935# gnd! 137.9fF
C2163 diff_5122_3935# gnd! 137.9fF
C2164 diff_5071_3935# gnd! 137.9fF
C2165 diff_5020_3935# gnd! 137.9fF
C2166 diff_4969_3935# gnd! 137.9fF
C2167 diff_4918_3935# gnd! 137.9fF
C2168 diff_4867_3935# gnd! 137.9fF
C2169 diff_4816_3935# gnd! 137.9fF
C2170 diff_4765_3935# gnd! 137.9fF
C2171 diff_4714_3935# gnd! 137.9fF
C2172 diff_4663_3935# gnd! 137.9fF
C2173 diff_4612_3935# gnd! 137.9fF
C2174 diff_4561_3935# gnd! 137.9fF
C2175 diff_4510_3935# gnd! 137.9fF
C2176 diff_4459_3935# gnd! 137.9fF
C2177 diff_4408_3935# gnd! 137.9fF
C2178 diff_4357_3935# gnd! 137.9fF
C2179 diff_4306_3935# gnd! 137.9fF
C2180 diff_4255_3935# gnd! 137.9fF
C2181 diff_4204_3935# gnd! 137.9fF
C2182 diff_4153_3935# gnd! 137.9fF
C2183 diff_4102_3935# gnd! 137.9fF
C2184 diff_4051_3935# gnd! 137.9fF
C2185 diff_4000_3935# gnd! 137.9fF
C2186 diff_3949_3935# gnd! 137.9fF
C2187 diff_3898_3935# gnd! 137.9fF
C2188 diff_3847_3935# gnd! 137.9fF
C2189 diff_3796_3935# gnd! 137.9fF
C2190 diff_3745_3935# gnd! 137.9fF
C2191 diff_3694_3935# gnd! 137.9fF
C2192 diff_3643_3935# gnd! 137.9fF
C2193 diff_3592_3935# gnd! 137.9fF
C2194 diff_3541_3935# gnd! 137.9fF
C2195 diff_3490_3935# gnd! 137.9fF
C2196 diff_3439_3935# gnd! 137.9fF
C2197 diff_3388_3935# gnd! 137.9fF
C2198 diff_3337_3935# gnd! 137.9fF
C2199 diff_3286_3935# gnd! 137.9fF
C2200 diff_3235_3935# gnd! 137.9fF
C2201 diff_3184_3935# gnd! 137.9fF
C2202 diff_3133_3935# gnd! 137.9fF
C2203 diff_3082_3935# gnd! 137.9fF
C2204 diff_3031_3935# gnd! 137.9fF
C2205 diff_2980_3935# gnd! 137.9fF
C2206 diff_2929_3935# gnd! 137.9fF
C2207 diff_2878_3935# gnd! 137.9fF
C2208 diff_2827_3935# gnd! 137.9fF
C2209 diff_2776_3935# gnd! 137.9fF
C2210 diff_2725_3935# gnd! 137.9fF
C2211 diff_2674_3935# gnd! 137.9fF
C2212 diff_2623_3935# gnd! 137.9fF
C2213 diff_2572_3935# gnd! 137.9fF
C2214 diff_2521_3935# gnd! 137.9fF
C2215 diff_2512_3979# gnd! 3320.1fF
C2216 diff_5734_3992# gnd! 129.8fF
C2217 diff_5683_3992# gnd! 129.8fF
C2218 diff_5632_3992# gnd! 129.8fF
C2219 diff_5581_3992# gnd! 129.8fF
C2220 diff_5530_3992# gnd! 129.8fF
C2221 diff_5479_3992# gnd! 129.8fF
C2222 diff_5428_3992# gnd! 129.8fF
C2223 diff_5377_3992# gnd! 129.8fF
C2224 diff_5326_3992# gnd! 129.8fF
C2225 diff_5275_3992# gnd! 129.8fF
C2226 diff_5224_3992# gnd! 129.8fF
C2227 diff_5173_3992# gnd! 129.8fF
C2228 diff_5122_3992# gnd! 129.8fF
C2229 diff_5071_3992# gnd! 129.8fF
C2230 diff_5020_3992# gnd! 129.8fF
C2231 diff_4969_3992# gnd! 129.8fF
C2232 diff_4918_3992# gnd! 129.8fF
C2233 diff_4867_3992# gnd! 129.8fF
C2234 diff_4816_3992# gnd! 129.8fF
C2235 diff_4765_3992# gnd! 129.8fF
C2236 diff_4714_3992# gnd! 129.8fF
C2237 diff_4663_3992# gnd! 129.8fF
C2238 diff_4612_3992# gnd! 129.8fF
C2239 diff_4561_3992# gnd! 129.8fF
C2240 diff_4510_3992# gnd! 129.8fF
C2241 diff_4459_3992# gnd! 129.8fF
C2242 diff_4408_3992# gnd! 129.8fF
C2243 diff_4357_3992# gnd! 129.8fF
C2244 diff_4306_3992# gnd! 129.8fF
C2245 diff_4255_3992# gnd! 129.8fF
C2246 diff_4204_3992# gnd! 129.8fF
C2247 diff_4153_3992# gnd! 129.8fF
C2248 diff_4102_3992# gnd! 129.8fF
C2249 diff_4051_3992# gnd! 129.8fF
C2250 diff_4000_3992# gnd! 129.8fF
C2251 diff_3949_3992# gnd! 129.8fF
C2252 diff_3898_3992# gnd! 129.8fF
C2253 diff_3847_3992# gnd! 129.8fF
C2254 diff_3796_3992# gnd! 129.8fF
C2255 diff_3745_3992# gnd! 129.8fF
C2256 diff_3694_3992# gnd! 129.8fF
C2257 diff_3643_3992# gnd! 129.8fF
C2258 diff_3592_3992# gnd! 129.8fF
C2259 diff_3541_3992# gnd! 129.8fF
C2260 diff_3490_3992# gnd! 129.8fF
C2261 diff_3439_3992# gnd! 129.8fF
C2262 diff_3388_3992# gnd! 129.8fF
C2263 diff_3337_3992# gnd! 129.8fF
C2264 diff_3286_3992# gnd! 129.8fF
C2265 diff_3235_3992# gnd! 129.8fF
C2266 diff_3184_3992# gnd! 129.8fF
C2267 diff_3133_3992# gnd! 129.8fF
C2268 diff_3082_3992# gnd! 129.8fF
C2269 diff_3031_3992# gnd! 129.8fF
C2270 diff_2980_3992# gnd! 129.8fF
C2271 diff_2929_3992# gnd! 129.8fF
C2272 diff_2878_3992# gnd! 129.8fF
C2273 diff_2827_3992# gnd! 129.8fF
C2274 diff_2776_3992# gnd! 129.8fF
C2275 diff_2725_3992# gnd! 129.8fF
C2276 diff_2674_3992# gnd! 129.8fF
C2277 diff_2623_3992# gnd! 129.8fF
C2278 diff_2572_3992# gnd! 129.8fF
C2279 diff_2521_3992# gnd! 129.8fF
C2280 diff_2512_4033# gnd! 3361.6fF
C2281 diff_5734_4046# gnd! 137.9fF
C2282 diff_5683_4046# gnd! 137.9fF
C2283 diff_5632_4046# gnd! 137.9fF
C2284 diff_5581_4046# gnd! 137.9fF
C2285 diff_5530_4046# gnd! 137.9fF
C2286 diff_5479_4046# gnd! 137.9fF
C2287 diff_5428_4046# gnd! 137.9fF
C2288 diff_5377_4046# gnd! 137.9fF
C2289 diff_5326_4046# gnd! 137.9fF
C2290 diff_5275_4046# gnd! 137.9fF
C2291 diff_5224_4046# gnd! 137.9fF
C2292 diff_5173_4046# gnd! 137.9fF
C2293 diff_5122_4046# gnd! 137.9fF
C2294 diff_5071_4046# gnd! 137.9fF
C2295 diff_5020_4046# gnd! 137.9fF
C2296 diff_4969_4046# gnd! 137.9fF
C2297 diff_4918_4046# gnd! 137.9fF
C2298 diff_4867_4046# gnd! 137.9fF
C2299 diff_4816_4046# gnd! 137.9fF
C2300 diff_4765_4046# gnd! 137.9fF
C2301 diff_4714_4046# gnd! 137.9fF
C2302 diff_4663_4046# gnd! 137.9fF
C2303 diff_4612_4046# gnd! 137.9fF
C2304 diff_4561_4046# gnd! 137.9fF
C2305 diff_4510_4046# gnd! 137.9fF
C2306 diff_4459_4046# gnd! 137.9fF
C2307 diff_4408_4046# gnd! 137.9fF
C2308 diff_4357_4046# gnd! 137.9fF
C2309 diff_4306_4046# gnd! 137.9fF
C2310 diff_4255_4046# gnd! 137.9fF
C2311 diff_4204_4046# gnd! 137.9fF
C2312 diff_4153_4046# gnd! 137.9fF
C2313 diff_4102_4046# gnd! 137.9fF
C2314 diff_4051_4046# gnd! 137.9fF
C2315 diff_4000_4046# gnd! 137.9fF
C2316 diff_3949_4046# gnd! 137.9fF
C2317 diff_3898_4046# gnd! 137.9fF
C2318 diff_3847_4046# gnd! 137.9fF
C2319 diff_3796_4046# gnd! 137.9fF
C2320 diff_3745_4046# gnd! 137.9fF
C2321 diff_3694_4046# gnd! 137.9fF
C2322 diff_3643_4046# gnd! 137.9fF
C2323 diff_3592_4046# gnd! 137.9fF
C2324 diff_3541_4046# gnd! 137.9fF
C2325 diff_3490_4046# gnd! 137.9fF
C2326 diff_3439_4046# gnd! 137.9fF
C2327 diff_3388_4046# gnd! 137.9fF
C2328 diff_3337_4046# gnd! 137.9fF
C2329 diff_3286_4046# gnd! 137.9fF
C2330 diff_3235_4046# gnd! 137.9fF
C2331 diff_3184_4046# gnd! 137.9fF
C2332 diff_3133_4046# gnd! 137.9fF
C2333 diff_3082_4046# gnd! 137.9fF
C2334 diff_3031_4046# gnd! 137.9fF
C2335 diff_2980_4046# gnd! 137.9fF
C2336 diff_2929_4046# gnd! 137.9fF
C2337 diff_2878_4046# gnd! 137.9fF
C2338 diff_2827_4046# gnd! 137.9fF
C2339 diff_2776_4046# gnd! 137.9fF
C2340 diff_2725_4046# gnd! 137.9fF
C2341 diff_2674_4046# gnd! 137.9fF
C2342 diff_2623_4046# gnd! 137.9fF
C2343 diff_2572_4046# gnd! 137.9fF
C2344 diff_2521_4046# gnd! 137.9fF
C2345 diff_2512_4090# gnd! 3554.3fF
C2346 diff_5734_4103# gnd! 129.8fF
C2347 diff_5683_4103# gnd! 129.8fF
C2348 diff_5632_4103# gnd! 129.8fF
C2349 diff_5581_4103# gnd! 129.8fF
C2350 diff_5530_4103# gnd! 129.8fF
C2351 diff_5479_4103# gnd! 129.8fF
C2352 diff_5428_4103# gnd! 129.8fF
C2353 diff_5377_4103# gnd! 129.8fF
C2354 diff_5326_4103# gnd! 129.8fF
C2355 diff_5275_4103# gnd! 129.8fF
C2356 diff_5224_4103# gnd! 129.8fF
C2357 diff_5173_4103# gnd! 129.8fF
C2358 diff_5122_4103# gnd! 129.8fF
C2359 diff_5071_4103# gnd! 129.8fF
C2360 diff_5020_4103# gnd! 129.8fF
C2361 diff_4969_4103# gnd! 129.8fF
C2362 diff_4918_4103# gnd! 129.8fF
C2363 diff_4867_4103# gnd! 129.8fF
C2364 diff_4816_4103# gnd! 129.8fF
C2365 diff_4765_4103# gnd! 129.8fF
C2366 diff_4714_4103# gnd! 129.8fF
C2367 diff_4663_4103# gnd! 129.8fF
C2368 diff_4612_4103# gnd! 129.8fF
C2369 diff_4561_4103# gnd! 129.8fF
C2370 diff_4510_4103# gnd! 129.8fF
C2371 diff_4459_4103# gnd! 129.8fF
C2372 diff_4408_4103# gnd! 129.8fF
C2373 diff_4357_4103# gnd! 129.8fF
C2374 diff_4306_4103# gnd! 129.8fF
C2375 diff_4255_4103# gnd! 129.8fF
C2376 diff_4204_4103# gnd! 129.8fF
C2377 diff_4153_4103# gnd! 129.8fF
C2378 diff_4102_4103# gnd! 129.8fF
C2379 diff_4051_4103# gnd! 129.8fF
C2380 diff_4000_4103# gnd! 129.8fF
C2381 diff_3949_4103# gnd! 129.8fF
C2382 diff_3898_4103# gnd! 129.8fF
C2383 diff_3847_4103# gnd! 129.8fF
C2384 diff_3796_4103# gnd! 129.8fF
C2385 diff_3745_4103# gnd! 129.8fF
C2386 diff_3694_4103# gnd! 129.8fF
C2387 diff_3643_4103# gnd! 129.8fF
C2388 diff_3592_4103# gnd! 129.8fF
C2389 diff_3541_4103# gnd! 129.8fF
C2390 diff_3490_4103# gnd! 129.8fF
C2391 diff_3439_4103# gnd! 129.8fF
C2392 diff_3388_4103# gnd! 129.8fF
C2393 diff_3337_4103# gnd! 129.8fF
C2394 diff_3286_4103# gnd! 129.8fF
C2395 diff_3235_4103# gnd! 129.8fF
C2396 diff_3184_4103# gnd! 129.8fF
C2397 diff_3133_4103# gnd! 129.8fF
C2398 diff_3082_4103# gnd! 129.8fF
C2399 diff_3031_4103# gnd! 129.8fF
C2400 diff_2980_4103# gnd! 129.8fF
C2401 diff_2929_4103# gnd! 129.8fF
C2402 diff_2878_4103# gnd! 129.8fF
C2403 diff_2827_4103# gnd! 129.8fF
C2404 diff_2776_4103# gnd! 129.8fF
C2405 diff_2725_4103# gnd! 129.8fF
C2406 diff_2674_4103# gnd! 129.8fF
C2407 diff_2623_4103# gnd! 129.8fF
C2408 diff_2572_4103# gnd! 129.8fF
C2409 diff_2521_4103# gnd! 129.8fF
C2410 diff_2218_3868# gnd! 493.6fF
C2411 diff_2080_3763# gnd! 504.6fF
C2412 diff_2053_3415# gnd! 3443.7fF
C2413 diff_1846_3766# gnd! 494.1fF
C2414 diff_1684_3766# gnd! 546.2fF
C2415 diff_1663_3415# gnd! 3390.2fF
C2416 diff_475_2011# gnd! 10359.2fF
C2417 diff_1459_3766# gnd! 528.7fF
C2418 diff_1303_3760# gnd! 499.0fF
C2419 diff_1276_3418# gnd! 3459.4fF
C2420 diff_1072_3769# gnd! 508.1fF
C2421 diff_916_3763# gnd! 527.7fF
C2422 diff_2512_4144# gnd! 3564.6fF
C2423 diff_6265_2299# gnd! 4706.6fF
C2424 diff_6223_2134# gnd! 4741.4fF
C2425 diff_5918_4184# gnd! 2889.6fF
C2426 diff_5734_4157# gnd! 137.9fF
C2427 diff_5683_4157# gnd! 137.9fF
C2428 diff_5632_4157# gnd! 137.9fF
C2429 diff_5581_4157# gnd! 137.9fF
C2430 diff_5530_4157# gnd! 137.9fF
C2431 diff_5479_4157# gnd! 137.9fF
C2432 diff_5428_4157# gnd! 137.9fF
C2433 diff_5377_4157# gnd! 137.9fF
C2434 diff_5326_4157# gnd! 137.9fF
C2435 diff_5275_4157# gnd! 137.9fF
C2436 diff_5224_4157# gnd! 137.9fF
C2437 diff_5173_4157# gnd! 137.9fF
C2438 diff_5122_4157# gnd! 137.9fF
C2439 diff_5071_4157# gnd! 137.9fF
C2440 diff_5020_4157# gnd! 137.9fF
C2441 diff_4969_4157# gnd! 137.9fF
C2442 diff_4918_4157# gnd! 137.9fF
C2443 diff_4867_4157# gnd! 137.9fF
C2444 diff_4816_4157# gnd! 137.9fF
C2445 diff_4765_4157# gnd! 137.9fF
C2446 diff_4714_4157# gnd! 137.9fF
C2447 diff_4663_4157# gnd! 137.9fF
C2448 diff_4612_4157# gnd! 137.9fF
C2449 diff_4561_4157# gnd! 137.9fF
C2450 diff_4510_4157# gnd! 137.9fF
C2451 diff_4459_4157# gnd! 137.9fF
C2452 diff_4408_4157# gnd! 137.9fF
C2453 diff_4357_4157# gnd! 137.9fF
C2454 diff_4306_4157# gnd! 137.9fF
C2455 diff_4255_4157# gnd! 137.9fF
C2456 diff_4204_4157# gnd! 137.9fF
C2457 diff_4153_4157# gnd! 137.9fF
C2458 diff_4102_4157# gnd! 137.9fF
C2459 diff_4051_4157# gnd! 137.9fF
C2460 diff_4000_4157# gnd! 137.9fF
C2461 diff_3949_4157# gnd! 137.9fF
C2462 diff_3898_4157# gnd! 137.9fF
C2463 diff_3847_4157# gnd! 137.9fF
C2464 diff_3796_4157# gnd! 137.9fF
C2465 diff_3745_4157# gnd! 137.9fF
C2466 diff_3694_4157# gnd! 137.9fF
C2467 diff_3643_4157# gnd! 137.9fF
C2468 diff_3592_4157# gnd! 137.9fF
C2469 diff_3541_4157# gnd! 137.9fF
C2470 diff_3490_4157# gnd! 137.9fF
C2471 diff_3439_4157# gnd! 137.9fF
C2472 diff_3388_4157# gnd! 137.9fF
C2473 diff_3337_4157# gnd! 137.9fF
C2474 diff_3286_4157# gnd! 137.9fF
C2475 diff_3235_4157# gnd! 137.9fF
C2476 diff_3184_4157# gnd! 137.9fF
C2477 diff_3133_4157# gnd! 137.9fF
C2478 diff_3082_4157# gnd! 137.9fF
C2479 diff_3031_4157# gnd! 137.9fF
C2480 diff_2980_4157# gnd! 137.9fF
C2481 diff_2929_4157# gnd! 137.9fF
C2482 diff_2878_4157# gnd! 137.9fF
C2483 diff_2827_4157# gnd! 137.9fF
C2484 diff_2776_4157# gnd! 137.9fF
C2485 diff_2725_4157# gnd! 137.9fF
C2486 diff_2674_4157# gnd! 137.9fF
C2487 diff_2623_4157# gnd! 137.9fF
C2488 diff_2572_4157# gnd! 137.9fF
C2489 diff_2521_4157# gnd! 137.9fF
C2490 diff_2512_4201# gnd! 3359.1fF
C2491 diff_6079_2449# gnd! 3869.4fF
C2492 diff_6034_2491# gnd! 4113.3fF
C2493 diff_5962_1069# gnd! 4001.8fF
C2494 diff_5905_1069# gnd! 4136.2fF
C2495 diff_2521_4214# gnd! 16118.7fF
C2496 diff_4144_4258# gnd! 9958.6fF
C2497 diff_6625_3571# gnd! 1578.2fF
C2498 diff_6535_4298# gnd! 1307.2fF
C2499 diff_6094_4246# gnd! 6836.5fF
C2500 diff_2509_4258# gnd! 11197.3fF
C2501 diff_6085_4357# gnd! 6368.1fF
C2502 diff_6880_4216# gnd! 671.7fF
C2503 diff_7004_4333# gnd! 510.7fF
C2504 diff_2011_4156# gnd! 5454.2fF
C2505 diff_1624_4156# gnd! 5461.2fF
C2506 Vdd gnd! 108985.0fF
C2507 diff_889_3418# gnd! 3458.4fF
C2508 diff_1237_4156# gnd! 5524.8fF
C2509 diff_847_4156# gnd! 5521.2fF
C2510 d0 gnd! 19333.9fF
C2511 d1 gnd! 19994.5fF
C2512 d3 gnd! 23806.3fF
C2513 sync gnd! 15164.1fF
C2514 d2 gnd! 19672.6fF
C2515 clk1 gnd! 14866.5fF
C2516 clk2 gnd! 19579.0fF
