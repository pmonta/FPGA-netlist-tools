* SPICE3 file created from 4004.ext - technology: 4004-nmos-buried-stacked

.option scale=0.001u

M1000 GND N0770 N0385 GND efet w=89900 l=11600
M1001 GND GND TEST_PAD GND efet w=119625 l=15225
M1002 POC_PAD GND GND GND efet w=118175 l=15225
M1003 GND N0754 N0761 GND efet w=26100 l=13050
M1004 GND PC0.11 N0785 GND efet w=30450 l=12325
M1005 N0785 N0406 N0770 GND efet w=26100 l=13050
M1006 GND N0301 N0754 GND efet w=21750 l=11600
M1007 N0761 N0301 N0753 GND efet w=78300 l=11600
M1008 N0754 VDD VDD GND efet w=7250 l=69600
M1009 N0754 N0289 GND GND efet w=23925 l=13775
M1010 VDD VDD N0761 GND efet w=8700 l=30450
M1011 N0753 N0289 GND GND efet w=136300 l=20300
M1012 D3 RADB1 N0386 GND efet w=44225 l=13775
M1013 N0385 RADB2 D3 GND efet w=49300 l=12325
M1014 N0770 WADB2 N0761 GND efet w=14500 l=13050
M1015 GND N0289 N0311 GND efet w=15225 l=12325
M1016 VDD N0325 N0301 GND efet w=9425 l=13775
M1017 N0289 M12+M22+CLK1~(M11+M12) D3 GND efet w=21025 l=12325
M1018 N0387 RADB0 D3 GND efet w=44950 l=10875
M1019 N0290 M12+M22+CLK1~(M11+M12) D2 GND efet w=20300 l=11600
M1020 N0311 N0290 N0312 GND efet w=14500 l=12325
M1021 N0301 N0290 N0302 GND efet w=26100 l=11600
M1022 GND N0290 N0755 GND efet w=123250 l=11600
M1023 GND N0740 SYNC GND efet w=1224525 l=10875
M1025 VDD VDD S00531 GND efet w=5800 l=13050
M1026 VDD S00531 N0740 GND efet w=10150 l=13050
M1028 VDD S00536 N0738 GND efet w=11600 l=11600
M1029 VDD VDD S00536 GND efet w=6525 l=13775
M1030 SYNC N0738 VDD GND efet w=679325 l=13050
M1031 N0388 RADB0 D2 GND efet w=42050 l=11600
M1032 VDD N0325 N0298 GND efet w=13050 l=14500
M1033 N0762 N0298 N0755 GND efet w=68150 l=11600
M1034 GND N0290 N0756 GND efet w=23200 l=10150
M1035 N0756 VDD VDD GND efet w=7250 l=68150
M1036 VDD VDD N0762 GND efet w=7250 l=27550
M1037 N0756 N0298 GND GND efet w=23925 l=12325
M1038 N0762 N0756 GND GND efet w=26100 l=11600
M1039 GND N0758 N0763 GND efet w=26100 l=11600
M1040 GND N0293 N0758 GND efet w=23925 l=11600
M1041 N0763 N0293 N0757 GND efet w=70325 l=12325
M1042 N0758 VDD VDD GND efet w=7975 l=67425
M1043 N0758 N0291 GND GND efet w=23200 l=11600
M1044 VDD VDD N0763 GND efet w=7975 l=29725
M1045 N0757 N0291 GND GND efet w=125425 l=12325
M1046 N0298 N0291 N0299 GND efet w=23200 l=18850
M1047 N0312 N0291 N0313 GND efet w=13050 l=11600
M1048 N0302 N0291 N0303 GND efet w=23200 l=11600
M1049 VDD N0325 N0293 GND efet w=9425 l=13775
M1050 N0291 M12+M22+CLK1~(M11+M12) D1 GND efet w=20300 l=11600
M1051 N0761 WADB1 N0774 GND efet w=14500 l=13775
M1052 N0778 WADB0 N0761 GND efet w=14500 l=11600
M1053 N0779 WADB0 N0762 GND efet w=17400 l=10150
M1054 N0762 WADB1 N0775 GND efet w=15950 l=13050
M1055 D2 RADB1 N0389 GND efet w=44225 l=12325
M1056 N0390 RADB2 D2 GND efet w=47125 l=10875
M1057 D1 RADB1 N0392 GND efet w=44225 l=14500
M1058 N0391 RADB2 D1 GND efet w=53650 l=10150
M1059 N0393 RADB0 D1 GND efet w=43500 l=11600
M1060 N0313 N0292 N0305 GND efet w=13050 l=11600
M1061 N0303 N0292 N0294 GND efet w=23200 l=11600
M1062 N0299 N0292 N0294 GND efet w=17400 l=11600
M1063 N0293 N0292 N0294 GND efet w=8700 l=11600
M1064 N0292 M12+M22+CLK1~(M11+M12) D0 GND efet w=23200 l=12325
M1065 GND N0292 N0759 GND efet w=125425 l=12325
M1066 N0305 N0325 VDD GND efet w=7975 l=12325
M1067 N0394 RADB0 D0 GND efet w=43500 l=13775
M1068 VDD N0325 N0752 GND efet w=10875 l=14500
M1069 N0764 N0752 N0759 GND efet w=69600 l=11600
M1070 GND N0292 N0760 GND efet w=29000 l=11600
M1071 N0760 VDD VDD GND efet w=7975 l=67425
M1072 VDD VDD N0764 GND efet w=7250 l=27550
M1073 GND N0307 N0294 GND efet w=31900 l=13050
M1074 N0760 N0752 GND GND efet w=21750 l=10150
M1075 N0752 N0307 GND GND efet w=14500 l=11600
M1076 N0764 N0760 GND GND efet w=27550 l=10150
M1077 GND N0738 N0740 GND efet w=101500 l=13050
M1078 N0305 N0307 N0306 GND efet w=14500 l=11600
M1079 GND N0295 N0738 GND efet w=112375 l=13775
M1080 GND PC2.11 N0821 GND efet w=26100 l=14500
M1081 N0806 PC1.11 GND GND efet w=19575 l=10875
M1082 N0770 N0424 N0806 GND efet w=26825 l=12325
M1083 N0821 N0434 N0770 GND efet w=26100 l=12325
M1084 N0770 N0444 N0834 GND efet w=28275 l=12325
M1085 N0834 PC3.11 GND GND efet w=23200 l=11600
M1086 N0386 N0774 GND GND efet w=72500 l=16675
M1087 N0385 N0381 PC0.11 GND efet w=6525 l=12325
M1088 PC1.11 N0410 N0385 GND efet w=7975 l=10875
M1089 N0386 N0381 PC0.7 GND efet w=6525 l=12325
M1090 PC1.7 N0410 N0386 GND efet w=5800 l=10150
M1091 N0786 N0406 N0774 GND efet w=27550 l=11600
M1092 GND PC0.7 N0786 GND efet w=25375 l=15225
M1093 N0385 N0426 PC2.11 GND efet w=6525 l=12325
M1094 PC3.11 N0439 N0385 GND efet w=5800 l=11600
M1095 N0386 N0426 PC2.7 GND efet w=6525 l=12325
M1096 GND N0778 N0387 GND efet w=72500 l=13775
M1097 N0787 N0406 N0778 GND efet w=24650 l=10875
M1098 GND PC0.3 N0787 GND efet w=24650 l=15225
M1099 N0807 PC1.7 GND GND efet w=22475 l=13775
M1100 N0774 N0424 N0807 GND efet w=27550 l=11600
M1101 N0822 N0434 N0774 GND efet w=26825 l=10875
M1102 GND PC2.7 N0822 GND efet w=23925 l=12325
M1103 N0388 N0779 GND GND efet w=71050 l=13775
M1104 N0387 N0381 PC0.3 GND efet w=7975 l=12325
M1105 N0808 PC1.3 GND GND efet w=23925 l=15225
M1106 PC3.7 N0439 N0386 GND efet w=5800 l=13050
M1107 VDD (~INH)(X11+X31)CLK1 N0770 GND efet w=8700 l=11600
M1108 D0 M12+M22+CLK1~(M11+M12) N0497 GND efet w=14500 l=13050
M1109 N0862 WRAB1 N0866 GND efet w=17400 l=13050
M1110 GND N0866 N0531 GND efet w=63800 l=11600
M1111 VDD VDD N0385 GND efet w=6525 l=31175
M1112 GND N0497 N0862 GND efet w=109475 l=12325
M1113 VDD VDD N0386 GND efet w=7250 l=30450
M1114 GND PC2.3 N0823 GND efet w=25375 l=12325
M1115 N0778 N0424 N0808 GND efet w=25375 l=11600
M1116 N0823 N0434 N0778 GND efet w=26825 l=10875
M1117 N0835 PC3.7 GND GND efet w=23925 l=13775
M1118 N0774 N0444 N0835 GND efet w=26825 l=10875
M1119 VDD (~INH)(X11+X31)CLK1 N0774 GND efet w=9425 l=13050
M1120 D0 RRAB1 N0531 GND efet w=46400 l=11600
M1121 N0532 RRAB0 D0 GND efet w=45675 l=13050
M1122 N0862 VDD VDD GND efet w=7975 l=22475
M1123 N0836 PC3.3 GND GND efet w=23925 l=13775
M1124 N0778 N0444 N0836 GND efet w=28275 l=10875
M1125 PC1.3 N0410 N0387 GND efet w=6525 l=10150
M1126 N0388 N0381 PC0.2 GND efet w=5800 l=10150
M1127 PC1.2 N0410 N0388 GND efet w=5800 l=10150
M1128 N0788 N0406 N0779 GND efet w=28275 l=10875
M1129 GND PC0.2 N0788 GND efet w=24650 l=13050
M1130 N0387 N0426 PC2.3 GND efet w=6525 l=12325
M1131 VDD (~INH)(X11+X31)CLK1 N0778 GND efet w=9425 l=13775
M1132 N0863 VDD VDD GND efet w=7975 l=21025
M1133 PC3.3 N0439 N0387 GND efet w=5800 l=11600
M1134 N0388 N0426 PC2.2 GND efet w=6525 l=10150
M1135 PC3.2 N0439 N0388 GND efet w=5800 l=11600
M1136 GND N0775 N0389 GND efet w=63800 l=11600
M1137 GND N0771 N0390 GND efet w=68875 l=13775
M1138 N0771 WADB2 N0762 GND efet w=13050 l=11600
M1139 N0789 N0406 N0775 GND efet w=24650 l=10875
M1140 GND PC0.6 N0789 GND efet w=24650 l=14500
M1141 N0809 PC1.2 GND GND efet w=23925 l=13775
M1142 N0779 N0424 N0809 GND efet w=26100 l=11600
M1143 N0824 N0434 N0779 GND efet w=26825 l=10875
M1144 GND PC2.2 N0824 GND efet w=24650 l=11600
M1145 GND N0498 N0863 GND efet w=114550 l=11600
M1146 VDD VDD N0387 GND efet w=7250 l=31900
M1147 VDD VDD N0388 GND efet w=7975 l=29725
M1148 N0837 PC3.2 GND GND efet w=23925 l=18125
M1149 N0810 PC1.6 GND GND efet w=22475 l=15225
M1150 GND PC2.6 N0825 GND efet w=23925 l=12325
M1151 N0775 N0424 N0810 GND efet w=26825 l=10875
M1152 N0825 N0434 N0775 GND efet w=25375 l=10875
M1153 N0779 N0444 N0837 GND efet w=26100 l=11600
M1154 VDD (~INH)(X11+X31)CLK1 N0779 GND efet w=8700 l=13050
M1155 D1 RRAB1 N0534 GND efet w=44950 l=11600
M1156 N0533 RRAB0 D1 GND efet w=46400 l=11600
M1157 N0880 WRAB0 N0862 GND efet w=13775 l=13050
M1158 N0532 N0880 GND GND efet w=59450 l=11600
M1159 N0903 N0543 N0866 GND efet w=24650 l=13050
M1160 GND R1.0 N0903 GND efet w=26100 l=14500
M1161 N0920 R3.0 GND GND efet w=24650 l=14500
M1162 N0866 N0565 N0920 GND efet w=24650 l=13050
M1163 N0929 N0581 N0866 GND efet w=26100 l=13050
M1164 GND R5.0 N0929 GND efet w=23925 l=13775
M1165 N0947 R7.0 GND GND efet w=25375 l=16675
M1166 N0866 N0591 N0947 GND efet w=24650 l=13775
M1167 N0956 N0616 N0866 GND efet w=26100 l=14500
M1168 GND R9.0 N0956 GND efet w=26825 l=19575
M1169 N0966 R11.0 GND GND efet w=25375 l=13775
M1170 N0531 N0529 R1.0 GND efet w=5800 l=11600
M1171 R3.0 N0544 N0531 GND efet w=5800 l=11600
M1172 N0531 N0569 R5.0 GND efet w=6525 l=12325
M1173 N0532 N0529 R0.0 GND efet w=5800 l=11600
M1174 R2.0 N0544 N0532 GND efet w=5800 l=11600
M1175 N0904 N0543 N0880 GND efet w=27550 l=13050
M1176 GND R0.0 N0904 GND efet w=24650 l=12325
M1177 R7.0 N0583 N0531 GND efet w=5800 l=11600
M1178 GND R0.1 N0905 GND efet w=23925 l=13775
M1179 N0498 M12+M22+CLK1~(M11+M12) D1 GND efet w=13050 l=11600
M1180 N0838 PC3.6 GND GND efet w=24650 l=16675
M1181 N0775 N0444 N0838 GND efet w=25375 l=10875
M1182 N0389 N0381 PC0.6 GND efet w=7975 l=12325
M1183 PC1.6 N0410 N0389 GND efet w=5800 l=12325
M1184 N0390 N0381 PC0.10 GND efet w=5800 l=10150
M1185 PC1.10 N0410 N0390 GND efet w=5800 l=10150
M1186 N0790 N0406 N0771 GND efet w=27550 l=10875
M1187 GND PC0.10 N0790 GND efet w=23925 l=12325
M1188 N0389 N0426 PC2.6 GND efet w=6525 l=10875
M1189 PC3.6 N0439 N0389 GND efet w=5800 l=10150
M1190 N0390 N0426 PC2.10 GND efet w=5800 l=10150
M1191 PC3.10 N0439 N0390 GND efet w=5800 l=10150
M1192 GND N0772 N0391 GND efet w=73225 l=12325
M1193 N0772 WADB2 N0763 GND efet w=14500 l=10875
M1194 N0763 WADB1 N0776 GND efet w=14500 l=13050
M1195 N0791 N0406 N0772 GND efet w=26825 l=10875
M1196 GND PC0.9 N0791 GND efet w=24650 l=13050
M1197 N0811 PC1.10 GND GND efet w=23200 l=14500
M1198 N0771 N0424 N0811 GND efet w=27550 l=11600
M1199 N0826 N0434 N0771 GND efet w=27550 l=11600
M1200 GND PC2.10 N0826 GND efet w=24650 l=11600
M1201 VDD (~INH)(X11+X31)CLK1 N0775 GND efet w=8700 l=11600
M1202 N0499 M12+M22+CLK1~(M11+M12) D2 GND efet w=14500 l=13050
M1203 N0780 WADB0 N0763 GND efet w=14500 l=13050
M1204 N0781 WADB0 N0764 GND efet w=15225 l=12325
M1205 N0392 N0776 GND GND efet w=65975 l=10875
M1206 N0391 N0381 PC0.9 GND efet w=6525 l=13050
M1207 N0812 PC1.9 GND GND efet w=23200 l=14500
M1208 GND PC2.9 N0827 GND efet w=26100 l=13050
M1209 N0772 N0424 N0812 GND efet w=25375 l=12325
M1210 N0827 N0434 N0772 GND efet w=26100 l=11600
M1211 N0839 PC3.10 GND GND efet w=24650 l=13050
M1212 N0771 N0444 N0839 GND efet w=26100 l=11600
M1213 VDD VDD N0389 GND efet w=6525 l=29725
M1214 D2 RRAB1 N0535 GND efet w=44225 l=12325
M1215 GND N0499 N0864 GND efet w=109475 l=10875
M1216 VDD VDD N0390 GND efet w=7975 l=28275
M1217 VDD (~INH)(X11+X31)CLK1 N0771 GND efet w=10150 l=11600
M1218 N0881 WRAB0 N0863 GND efet w=13050 l=13050
M1219 N0863 WRAB1 N0867 GND efet w=13050 l=11600
M1220 N0864 WRAB1 N0868 GND efet w=13050 l=11600
M1221 N0840 PC3.9 GND GND efet w=25375 l=13775
M1222 PC1.9 N0410 N0391 GND efet w=5800 l=11600
M1223 PC1.5 N0410 N0392 GND efet w=5800 l=13050
M1224 N0392 N0381 PC0.5 GND efet w=5800 l=11600
M1225 N0792 N0406 N0776 GND efet w=28275 l=10875
M1226 GND PC0.5 N0792 GND efet w=23925 l=12325
M1227 N0391 N0426 PC2.9 GND efet w=5800 l=10150
M1228 N0772 N0444 N0840 GND efet w=25375 l=12325
M1229 PC3.9 N0439 N0391 GND efet w=5800 l=10150
M1230 N0392 N0426 PC2.5 GND efet w=5800 l=10150
M1231 N0813 PC1.5 GND GND efet w=23925 l=12325
M1232 GND PC0.1 N0793 GND efet w=25375 l=13775
M1233 GND N0780 N0393 GND efet w=69600 l=11600
M1234 N0793 N0406 N0780 GND efet w=25375 l=10875
M1235 N0776 N0424 N0813 GND efet w=26825 l=10875
M1236 N0828 N0434 N0776 GND efet w=26100 l=11600
M1237 GND PC2.5 N0828 GND efet w=26100 l=11600
M1238 PC3.5 N0439 N0392 GND efet w=5800 l=11600
M1239 N0841 PC3.5 GND GND efet w=23925 l=13775
M1240 N0776 N0444 N0841 GND efet w=24650 l=11600
M1241 N0394 N0781 GND GND efet w=68150 l=13050
M1242 N0393 N0381 PC0.1 GND efet w=5800 l=11600
M1243 N0814 PC1.1 GND GND efet w=24650 l=13050
M1244 GND PC2.1 N0829 GND efet w=23925 l=12325
M1245 N0780 N0424 N0814 GND efet w=26100 l=11600
M1246 N0829 N0434 N0780 GND efet w=26100 l=11600
M1247 N0864 VDD VDD GND efet w=7250 l=20300
M1248 VDD (~INH)(X11+X31)CLK1 N0772 GND efet w=9425 l=13775
M1249 VDD VDD N0391 GND efet w=7975 l=28275
M1250 N0865 VDD VDD GND efet w=7975 l=20300
M1251 GND N0500 N0865 GND efet w=114550 l=13050
M1252 N0536 RRAB0 D2 GND efet w=44950 l=11600
M1253 GND N0881 N0533 GND efet w=59450 l=11600
M1254 N0534 N0867 GND GND efet w=60175 l=10875
M1255 N0905 N0543 N0881 GND efet w=26100 l=11600
M1256 N0921 R2.0 GND GND efet w=29000 l=14500
M1257 N0880 N0565 N0921 GND efet w=27550 l=11600
M1258 N0930 N0581 N0880 GND efet w=26100 l=13050
M1259 N0532 N0569 R4.0 GND efet w=5800 l=11600
M1260 GND R4.0 N0930 GND efet w=21750 l=13050
M1261 N0922 R2.1 GND GND efet w=26825 l=15225
M1262 N0533 N0529 R0.1 GND efet w=5800 l=11600
M1263 R6.0 N0583 N0532 GND efet w=5800 l=11600
M1264 N0948 R6.0 GND GND efet w=24650 l=15950
M1265 N0866 N0632 N0966 GND efet w=30450 l=13050
M1266 N0975 N0645 N0866 GND efet w=27550 l=13050
M1267 GND R13.0 N0975 GND efet w=26825 l=18850
M1268 N0984 R15.0 GND GND efet w=27550 l=13050
M1269 N0866 N0657 N0984 GND efet w=29000 l=13775
M1270 N0880 N0591 N0948 GND efet w=26825 l=13775
M1271 N0531 N0598 R9.0 GND efet w=5800 l=13050
M1272 R11.0 N0619 N0531 GND efet w=7975 l=12325
M1273 N0532 N0598 R8.0 GND efet w=7250 l=13050
M1274 GND R8.0 N0957 GND efet w=21750 l=14500
M1275 R10.0 N0619 N0532 GND efet w=6525 l=12325
M1276 N0957 N0616 N0880 GND efet w=24650 l=11600
M1277 GND R4.1 N0931 GND efet w=23200 l=15225
M1278 N0881 N0565 N0922 GND efet w=28275 l=10875
M1279 N0931 N0581 N0881 GND efet w=25375 l=10875
M1280 N0531 N0634 R13.0 GND efet w=5800 l=13050
M1281 R15.0 N0647 N0531 GND efet w=5800 l=14500
M1282 N0532 N0634 R12.0 GND efet w=7250 l=13775
M1283 N0949 R6.1 GND GND efet w=25375 l=16675
M1284 N0881 N0591 N0949 GND efet w=27550 l=13050
M1285 R2.1 N0544 N0533 GND efet w=5800 l=11600
M1286 N0534 N0529 R1.1 GND efet w=5800 l=11600
M1287 R3.1 N0544 N0534 GND efet w=5800 l=11600
M1288 N0906 N0543 N0867 GND efet w=27550 l=11600
M1289 GND R1.1 N0906 GND efet w=23200 l=13050
M1290 N0533 N0569 R4.1 GND efet w=6525 l=10875
M1291 N0958 N0616 N0881 GND efet w=25375 l=13050
M1292 GND R8.1 N0958 GND efet w=22475 l=13775
M1293 N0967 R10.0 GND GND efet w=26825 l=13775
M1294 N0880 N0632 N0967 GND efet w=25375 l=12325
M1295 N0976 N0645 N0880 GND efet w=25375 l=12325
M1296 GND R12.0 N0976 GND efet w=20300 l=13050
M1297 R14.0 N0647 N0532 GND efet w=7975 l=15225
M1298 N0968 R10.1 GND GND efet w=26100 l=13050
M1299 N0881 N0632 N0968 GND efet w=26100 l=12325
M1300 N0985 R14.0 GND GND efet w=26100 l=13050
M1301 N0880 N0657 N0985 GND efet w=26100 l=14500
M1302 R6.1 N0583 N0533 GND efet w=5800 l=11600
M1303 N0534 N0569 R5.1 GND efet w=5800 l=10875
M1304 R7.1 N0583 N0534 GND efet w=5800 l=11600
M1305 N0923 R3.1 GND GND efet w=24650 l=13050
M1306 GND R1.2 N0907 GND efet w=23925 l=13775
M1307 GND N0868 N0535 GND efet w=58725 l=12325
M1308 N0907 N0543 N0868 GND efet w=25375 l=12325
M1309 N0867 N0565 N0923 GND efet w=29000 l=10875
M1310 N0932 N0581 N0867 GND efet w=26100 l=11600
M1311 GND R5.1 N0932 GND efet w=23200 l=13050
M1312 N0533 N0598 R8.1 GND efet w=5800 l=13050
M1313 N0977 N0645 N0881 GND efet w=24650 l=11600
M1314 GND R12.1 N0977 GND efet w=21025 l=13775
M1315 VDD SC(A22+M22)CLK2 N0866 GND efet w=11600 l=14500
M1316 VDD VDD N0531 GND efet w=8700 l=33350
M1317 VDD VDD N0532 GND efet w=8700 l=33350
M1318 VDD SC(A22+M22)CLK2 N0880 GND efet w=13050 l=11600
M1319 N0986 R14.1 GND GND efet w=26100 l=13050
M1320 R10.1 N0619 N0533 GND efet w=5800 l=11600
M1321 N0534 N0598 R9.1 GND efet w=5800 l=14500
M1322 N0536 N0882 GND GND efet w=62350 l=11600
M1323 N0882 WRAB0 N0864 GND efet w=13050 l=11600
M1324 N0924 R3.2 GND GND efet w=23200 l=13050
M1325 N0868 N0565 N0924 GND efet w=27550 l=11600
M1326 N0933 N0581 N0868 GND efet w=24650 l=11600
M1327 GND R5.2 N0933 GND efet w=23200 l=13050
M1328 N0950 R7.1 GND GND efet w=23925 l=13775
M1329 N0867 N0591 N0950 GND efet w=27550 l=11600
M1330 N0959 N0616 N0867 GND efet w=26100 l=11600
M1331 GND R9.1 N0959 GND efet w=23200 l=14500
M1332 R11.1 N0619 N0534 GND efet w=7250 l=13050
M1333 N0533 N0634 R12.1 GND efet w=5800 l=13050
M1334 N0881 N0657 N0986 GND efet w=26100 l=14500
M1335 R14.1 N0647 N0533 GND efet w=6525 l=13775
M1336 N0534 N0634 R13.1 GND efet w=7250 l=13050
M1337 N0969 R11.1 GND GND efet w=23200 l=13775
M1338 N0867 N0632 N0969 GND efet w=25375 l=13775
M1339 N0978 N0645 N0867 GND efet w=24650 l=12325
M1340 GND R13.1 N0978 GND efet w=20300 l=11600
M1341 N0951 R7.2 GND GND efet w=23200 l=14500
M1342 N0535 N0529 R1.2 GND efet w=5800 l=12325
M1343 R3.2 N0544 N0535 GND efet w=6525 l=12325
M1344 N0536 N0529 R0.2 GND efet w=7975 l=10875
M1345 R2.2 N0544 N0536 GND efet w=5800 l=11600
M1346 N0908 N0543 N0882 GND efet w=24650 l=11600
M1347 GND R0.2 N0908 GND efet w=23200 l=13050
M1348 N0868 N0591 N0951 GND efet w=24650 l=11600
M1349 N0960 N0616 N0868 GND efet w=24650 l=11600
M1350 GND R9.2 N0960 GND efet w=23925 l=16675
M1351 R15.1 N0647 N0534 GND efet w=7975 l=15225
M1352 N0987 R15.1 GND GND efet w=27550 l=14500
M1353 N0970 R11.2 GND GND efet w=23200 l=14500
M1354 N0535 N0569 R5.2 GND efet w=5800 l=13050
M1355 R7.2 N0583 N0535 GND efet w=7250 l=10875
M1356 N0536 N0569 R4.2 GND efet w=5800 l=11600
M1357 GND R0.3 N0909 GND efet w=23925 l=13775
M1358 VDD VDD N0392 GND efet w=7250 l=29000
M1359 VDD (~INH)(X11+X31)CLK1 N0776 GND efet w=10875 l=11600
M1360 N0500 M12+M22+CLK1~(M11+M12) D3 GND efet w=13050 l=11600
M1361 D3 RRAB1 N0538 GND efet w=46400 l=11600
M1362 N0537 RRAB0 D3 GND efet w=44950 l=11600
M1363 N0842 PC3.1 GND GND efet w=23925 l=15225
M1364 PC1.1 N0410 N0393 GND efet w=5800 l=11600
M1365 N0780 N0444 N0842 GND efet w=25375 l=11600
M1366 N0393 N0426 PC2.1 GND efet w=5800 l=10150
M1367 PC3.1 N0439 N0393 GND efet w=5800 l=10150
M1368 N0394 N0381 PC0.0 GND efet w=5800 l=11600
M1369 N0794 N0406 N0781 GND efet w=27550 l=10875
M1370 GND PC0.0 N0794 GND efet w=23925 l=12325
M1371 PC1.0 N0410 N0394 GND efet w=5800 l=11600
M1372 N0815 PC1.0 GND GND efet w=23925 l=13775
M1373 N0394 N0426 PC2.0 GND efet w=5800 l=10150
M1374 GND N0777 N0395 GND efet w=68150 l=11600
M1375 GND PC0.4 N0795 GND efet w=24650 l=14500
M1376 N0764 WADB1 N0777 GND efet w=14500 l=11600
M1377 D0 RADB1 N0395 GND efet w=43500 l=11600
M1378 N0396 RADB2 D0 GND efet w=48575 l=10875
M1379 VDD N0325 N0306 GND efet w=7250 l=11600
M1380 N0314 N0306 GND GND efet w=29000 l=11600
M1381 N0795 N0406 N0777 GND efet w=26100 l=11600
M1382 N0781 N0424 N0815 GND efet w=25375 l=10875
M1383 N0830 N0434 N0781 GND efet w=26100 l=11600
M1384 GND PC2.0 N0830 GND efet w=23925 l=13050
M1385 PC3.0 N0439 N0394 GND efet w=5800 l=10875
M1386 N0843 PC3.0 GND GND efet w=22475 l=15225
M1387 N0816 PC1.4 GND GND efet w=21750 l=14500
M1388 N0777 N0424 N0816 GND efet w=25375 l=10875
M1389 GND N0773 N0396 GND efet w=68875 l=13775
M1390 N0773 WADB2 N0764 GND efet w=13050 l=11600
M1391 N0395 N0381 PC0.4 GND efet w=6525 l=13775
M1392 N0831 N0434 N0777 GND efet w=24650 l=11600
M1393 GND PC2.4 N0831 GND efet w=23200 l=14500
M1394 N0781 N0444 N0843 GND efet w=24650 l=11600
M1395 VDD (~INH)(X11+X31)CLK1 N0780 GND efet w=8700 l=13050
M1396 N0883 WRAB0 N0865 GND efet w=13050 l=11600
M1397 N0865 WRAB1 N0869 GND efet w=15225 l=10150
M1398 GND N0883 N0537 GND efet w=59450 l=11600
M1399 N0909 N0543 N0883 GND efet w=24650 l=11600
M1400 N0925 R2.2 GND GND efet w=23925 l=13775
M1401 N0882 N0565 N0925 GND efet w=24650 l=11600
M1402 N0934 N0581 N0882 GND efet w=24650 l=13050
M1403 GND R4.2 N0934 GND efet w=25375 l=12325
M1404 N0926 R2.3 GND GND efet w=23200 l=13050
M1405 R6.2 N0583 N0536 GND efet w=5800 l=11600
M1406 N0868 N0632 N0970 GND efet w=25375 l=12325
M1407 N0979 N0645 N0868 GND efet w=27550 l=11600
M1408 GND R13.2 N0979 GND efet w=20300 l=11600
M1409 N0535 N0598 R9.2 GND efet w=5800 l=11600
M1410 R11.2 N0619 N0535 GND efet w=6525 l=13050
M1411 N0867 N0657 N0987 GND efet w=25375 l=12325
M1412 VDD SC(A22+M22)CLK2 N0881 GND efet w=11600 l=14500
M1413 VDD VDD N0533 GND efet w=7250 l=37700
M1414 VDD VDD N0534 GND efet w=7975 l=35525
M1415 VDD SC(A22+M22)CLK2 N0867 GND efet w=12325 l=13775
M1416 N0988 R15.2 GND GND efet w=27550 l=14500
M1417 N0868 N0657 N0988 GND efet w=26100 l=12325
M1418 N0536 N0598 R8.2 GND efet w=5800 l=11600
M1419 N0538 N0869 GND GND efet w=59450 l=11600
M1420 N0883 N0565 N0926 GND efet w=24650 l=11600
M1421 N0935 N0581 N0883 GND efet w=24650 l=11600
M1422 GND R4.3 N0935 GND efet w=26825 l=13050
M1423 N0952 R6.2 GND GND efet w=23925 l=15225
M1424 N0882 N0591 N0952 GND efet w=28275 l=10875
M1425 N0961 N0616 N0882 GND efet w=29725 l=10875
M1426 GND R8.2 N0961 GND efet w=25375 l=13775
M1427 R10.2 N0619 N0536 GND efet w=5800 l=11600
M1428 N0535 N0634 R13.2 GND efet w=5800 l=12325
M1429 R15.2 N0647 N0535 GND efet w=6525 l=13775
M1430 N0536 N0634 R12.2 GND efet w=6525 l=13775
M1431 R14.2 N0647 N0536 GND efet w=6525 l=15225
M1432 N0971 R10.2 GND GND efet w=24650 l=13050
M1433 N0882 N0632 N0971 GND efet w=26825 l=12325
M1434 N0980 N0645 N0882 GND efet w=29000 l=11600
M1435 N0953 R6.3 GND GND efet w=23200 l=13775
M1436 N0537 N0529 R0.3 GND efet w=6525 l=13775
M1437 R2.3 N0544 N0537 GND efet w=4350 l=12325
M1438 N0538 N0529 R1.3 GND efet w=7250 l=11600
M1439 R3.3 N0544 N0538 GND efet w=5800 l=11600
M1440 N0910 N0543 N0869 GND efet w=24650 l=13775
M1441 GND R1.3 N0910 GND efet w=23200 l=13050
M1442 N0537 N0569 R4.3 GND efet w=7250 l=11600
M1443 N0883 N0591 N0953 GND efet w=26825 l=11600
M1444 N0962 N0616 N0883 GND efet w=26825 l=12325
M1445 GND R8.3 N0962 GND efet w=26100 l=15950
M1446 GND R12.2 N0980 GND efet w=21025 l=15225
M1447 N0972 R10.3 GND GND efet w=24650 l=14500
M1448 R6.3 N0583 N0537 GND efet w=6525 l=13775
M1449 N0538 N0569 R5.3 GND efet w=5800 l=11600
M1450 VDD VDD N0393 GND efet w=5800 l=30450
M1451 GND N0461 N0469 GND efet w=13050 l=13050
M1452 N0469 VDD VDD GND efet w=8700 l=65250
M1453 N0461 N0469 GND GND efet w=11600 l=11600
M1454 N0927 R3.3 GND GND efet w=23925 l=13775
M1455 N0869 N0565 N0927 GND efet w=27550 l=11600
M1456 N0936 N0581 N0869 GND efet w=27550 l=13050
M1457 GND R5.3 N0936 GND efet w=27550 l=13050
M1458 R7.3 N0583 N0538 GND efet w=5800 l=11600
M1459 N0883 N0632 N0972 GND efet w=26100 l=13050
M1460 N0981 N0645 N0883 GND efet w=31175 l=13775
M1461 GND R12.3 N0981 GND efet w=22475 l=17400
M1462 N0989 R14.2 GND GND efet w=29725 l=15225
M1463 N0882 N0657 N0989 GND efet w=27550 l=13050
M1464 VDD SC(A22+M22)CLK2 N0868 GND efet w=14500 l=14500
M1465 VDD VDD N0535 GND efet w=8700 l=34075
M1466 VDD VDD N0536 GND efet w=7975 l=32625
M1467 VDD SC(A22+M22)CLK2 N0882 GND efet w=11600 l=13050
M1468 N0990 R14.3 GND GND efet w=29000 l=13050
M1469 N0883 N0657 N0990 GND efet w=29000 l=11600
M1470 N0537 N0598 R8.3 GND efet w=5800 l=11600
M1471 R10.3 N0619 N0537 GND efet w=5800 l=13775
M1472 N0538 N0598 R9.3 GND efet w=5800 l=11600
M1473 N0954 R7.3 GND GND efet w=23925 l=13775
M1474 N0869 N0591 N0954 GND efet w=27550 l=11600
M1475 N0963 N0616 N0869 GND efet w=27550 l=11600
M1476 GND R9.3 N0963 GND efet w=25375 l=13775
M1477 R11.3 N0619 N0538 GND efet w=5800 l=11600
M1478 N0973 R11.3 GND GND efet w=26825 l=14500
M1479 N0537 N0634 R12.3 GND efet w=5800 l=11600
M1480 VDD SC(A22+M22)CLK2 N0883 GND efet w=11600 l=13050
M1481 R14.3 N0647 N0537 GND efet w=5800 l=13050
M1482 N0538 N0634 R13.3 GND efet w=5800 l=13050
M1483 R15.3 N0647 N0538 GND efet w=7250 l=14500
M1484 N0869 N0632 N0973 GND efet w=26100 l=12325
M1485 N0982 N0645 N0869 GND efet w=26100 l=13050
M1486 GND R13.3 N0982 GND efet w=27550 l=15950
M1487 VDD VDD N0537 GND efet w=8700 l=34075
M1488 GND GND CLK2 GND efet w=118175 l=13775
M1489 GND GND CLK1 GND efet w=113100 l=13050
M1490 VDD VDD N0538 GND efet w=8700 l=34075
M1491 N0991 R15.3 GND GND efet w=26100 l=15950
M1492 N0869 N0657 N0991 GND efet w=26825 l=12325
M1493 VDD SC(A22+M22)CLK2 N0869 GND efet w=11600 l=14500
M1494 VDD VDD N0394 GND efet w=5800 l=29000
M1495 VDD VDD N0461 GND efet w=5800 l=65250
M1496 ADDR-RFSH.1 VDD VDD GND efet w=8700 l=66700
M1497 GND N0461 ADDR-RFSH.1 GND efet w=15225 l=10875
M1498 N0453 N0469 GND GND efet w=14500 l=11600
M1499 GND N0902 N0543 GND efet w=14500 l=11600
M1500 GND N0902 N0529 GND efet w=11600 l=11600
M1501 GND N0919 N0544 GND efet w=11600 l=11600
M1502 GND N0919 N0565 GND efet w=14500 l=11600
M1503 VDD VDD N0453 GND efet w=9425 l=65975
M1504 VDD (~INH)(X11+X31)CLK1 N0781 GND efet w=9425 l=10875
M1505 N0902 VDD VDD GND efet w=6525 l=61625
M1506 N0543 N0530 (~POC)&CLK2&SC(A32+X12) GND efet w=16675 l=10875
M1507 N0529 N0530 CLK2&SC(A12+M12) GND efet w=13775 l=13050
M1508 N0544 N0545 CLK2&SC(A12+M12) GND efet w=12325 l=10875
M1509 N0565 N0545 (~POC)&CLK2&SC(A32+X12) GND efet w=16675 l=12325
M1510 N0844 PC3.4 GND GND efet w=22475 l=18125
M1511 ADDR-RFSH.1 N0455 N0489 GND efet w=8700 l=10150
M1512 N0453 N0455 N0454 GND efet w=8700 l=13050
M1513 PC1.4 N0410 N0395 GND efet w=6525 l=12325
M1514 N0396 N0381 PC0.8 GND efet w=5800 l=11600
M1515 N0796 N0406 N0773 GND efet w=27550 l=13050
M1516 VDD VDD N0314 GND efet w=7250 l=65250
M1517 GND A32 N0712 GND efet w=24650 l=11600
M1518 N0314 CLK2 N0315 GND efet w=13050 l=14500
M1519 CMROM N0717 VDD GND efet w=417600 l=11600
M1520 GND N0737 CMROM GND efet w=607550 l=10875
M1521 N0712 A22 GND GND efet w=26825 l=12325
M1522 N0325 VDD CLK1 GND efet w=34800 l=11600
M1523 VDD VDD WADB1 GND efet w=5800 l=27550
M1524 GND A12 N0711 GND efet w=13050 l=12325
M1525 N0316 N0315 GND GND efet w=20300 l=11600
M1526 WADB0 VDD VDD GND efet w=7250 l=27550
M1527 GND N0300 WADB0 GND efet w=29000 l=13050
M1528 VDD VDD N0316 GND efet w=6525 l=51475
M1529 N0711 VDD VDD GND efet w=6525 l=67425
M1530 N0317 CLK1 N0316 GND efet w=8700 l=11600
M1531 GND N0326 WADB0 GND efet w=36250 l=11600
M1532 GND PC0.8 N0796 GND efet w=23925 l=12325
M1533 PC1.8 N0410 N0396 GND efet w=5800 l=11600
M1534 N0777 N0444 N0844 GND efet w=24650 l=11600
M1535 N0395 N0426 PC2.4 GND efet w=6525 l=10875
M1536 PC3.4 N0439 N0395 GND efet w=5800 l=10150
M1537 N0396 N0426 PC2.8 GND efet w=5800 l=10150
M1538 PC3.8 N0439 N0396 GND efet w=5800 l=10150
M1539 N0817 PC1.8 GND GND efet w=26100 l=13050
M1540 N0773 N0424 N0817 GND efet w=27550 l=13050
M1541 N0832 N0434 N0773 GND efet w=25375 l=12325
M1542 WADB2 VDD VDD GND efet w=7975 l=31175
M1543 GND PC2.8 N0832 GND efet w=25375 l=13050
M1544 N0845 PC3.8 GND GND efet w=23925 l=15225
M1545 N0773 N0444 N0845 GND efet w=26825 l=13775
M1546 VDD (~INH)(X11+X31)CLK1 N0777 GND efet w=8700 l=11600
M1547 N0488 N0463 N0469 GND efet w=21750 l=12325
M1548 VDD VDD N0395 GND efet w=6525 l=32625
M1549 GND N0489 N0488 GND efet w=34075 l=11600
M1550 N0462 N0454 GND GND efet w=34800 l=11600
M1551 N0461 N0463 N0462 GND efet w=20300 l=11600
M1552 VDD VDD N0396 GND efet w=6525 l=31175
M1553 GND N0928 N0581 GND efet w=14500 l=10150
M1554 GND N0928 N0569 GND efet w=11600 l=10150
M1555 GND N0938 N0583 GND efet w=13050 l=10150
M1556 GND N0938 N0591 GND efet w=15950 l=10150
M1557 GND N0955 N0616 GND efet w=13775 l=10875
M1558 N0581 N0570 (~POC)&CLK2&SC(A32+X12) GND efet w=14500 l=11600
M1559 N0569 N0570 CLK2&SC(A12+M12) GND efet w=12325 l=12325
M1560 N0583 N0584 CLK2&SC(A12+M12) GND efet w=13050 l=11600
M1561 N0591 N0584 (~POC)&CLK2&SC(A32+X12) GND efet w=14500 l=13050
M1562 GND N0530 N0902 GND efet w=11600 l=13050
M1563 N0919 N0545 GND GND efet w=10150 l=11600
M1564 GND N0570 N0928 GND efet w=10875 l=12325
M1565 N0938 N0584 GND GND efet w=10150 l=13050
M1566 GND N0955 N0598 GND efet w=13050 l=10875
M1567 GND N0965 N0619 GND efet w=11600 l=11600
M1568 GND N0965 N0632 GND efet w=13050 l=12325
M1569 N0616 N0599 (~POC)&CLK2&SC(A32+X12) GND efet w=14500 l=10875
M1570 CLK2&SC(A12+M12) N0599 N0598 GND efet w=12325 l=10875
M1571 N0619 N0620 CLK2&SC(A12+M12) GND efet w=12325 l=10875
M1572 N0632 N0620 (~POC)&CLK2&SC(A32+X12) GND efet w=13050 l=10150
M1573 GND N0599 N0955 GND efet w=12325 l=12325
M1575 RRAB1 S00557 VDD GND efet w=10150 l=23200
M1576 S00557 VDD VDD GND efet w=6525 l=13775
M1577 VDD (~INH)(X11+X31)CLK1 N0773 GND efet w=10150 l=11600
M1578 N0463 VDD VDD GND efet w=6525 l=71775
M1579 GND N0455 N0463 GND efet w=11600 l=11600
M1580 N0455 N0463 GND GND efet w=13050 l=11600
M1581 N0919 VDD VDD GND efet w=6525 l=45675
M1582 VDD VDD N0928 GND efet w=7975 l=51475
M1583 N0965 N0620 GND GND efet w=11600 l=13050
M1584 GND N0974 N0645 GND efet w=14500 l=11600
M1585 GND N0974 N0634 GND efet w=11600 l=11600
M1586 GND N0983 N0647 GND efet w=11600 l=11600
M1587 GND N0983 N0657 GND efet w=14500 l=11600
M1588 N0645 N0635 (~POC)&CLK2&SC(A32+X12) GND efet w=15225 l=10875
M1589 N0634 N0635 CLK2&SC(A12+M12) GND efet w=12325 l=10875
M1590 N0647 N0648 CLK2&SC(A12+M12) GND efet w=12325 l=10875
M1591 N0657 N0648 (~POC)&CLK2&SC(A32+X12) GND efet w=14500 l=11600
M1592 N0938 VDD VDD GND efet w=5800 l=47850
M1593 VDD VDD N0955 GND efet w=6525 l=52925
M1594 GND N0635 N0974 GND efet w=10150 l=13050
M1595 N0983 N0648 GND GND efet w=10150 l=13050
M1596 VDD VDD N0613 GND efet w=13050 l=45675
M1597 N0965 VDD VDD GND efet w=6525 l=48575
M1598 VDD VDD N0974 GND efet w=5800 l=47850
M1599 N0983 VDD VDD GND efet w=5800 l=47850
M1600 N0539 N0540 GND GND efet w=27550 l=13050
M1601 VDD VDD N0540 GND efet w=7250 l=29000
M1602 VDD VDD N0455 GND efet w=6525 l=68875
M1603 ADDR-RFSH.0 VDD VDD GND efet w=9425 l=73950
M1604 GND N0455 ADDR-RFSH.0 GND efet w=13775 l=10875
M1605 N0503 N0463 GND GND efet w=13050 l=11600
M1606 VDD VDD N0503 GND efet w=8700 l=66700
M1607 S00564 VDD VDD GND efet w=6525 l=13775
M1609 RRAB0 S00564 VDD GND efet w=7250 l=21750
M1610 WADB1 N0318 GND GND efet w=27550 l=11600
M1611 GND N0304 WADB2 GND efet w=29000 l=13050
M1612 GND N0300 WADB1 GND efet w=27550 l=12325
M1613 WADB2 N0300 GND GND efet w=29725 l=10875
M1614 GND N0783 N0406 GND efet w=15950 l=10150
M1615 GND N0783 N0381 GND efet w=11600 l=10150
M1616 GND N0804 N0410 GND efet w=11600 l=11600
M1617 GND N0804 N0424 GND efet w=15950 l=10150
M1618 N0406 N0382 (~POC)CLK2(X12+X32)~INH GND efet w=15950 l=11600
M1619 N0381 N0382 ((~SC)(JIN+FIN))CLK1(M11+X21~INH) GND efet w=10150 l=11600
M1620 N0410 N0411 ((~SC)(JIN+FIN))CLK1(M11+X21~INH) GND efet w=12325 l=12325
M1621 N0424 N0411 (~POC)CLK2(X12+X32)~INH GND efet w=15950 l=11600
M1622 N0737 VDD VDD GND efet w=9425 l=13775
M1623 N0711 N0732 N0712 GND efet w=23200 l=10150
M1624 GND N0820 N0434 GND efet w=15950 l=10150
M1625 N0426 N0820 GND GND efet w=11600 l=11600
M1626 GND N0833 N0439 GND efet w=11600 l=11600
M1627 N0444 N0833 GND GND efet w=15950 l=13050
M1628 ADDR-RFSH.0 CLK1 N0519 GND efet w=7250 l=11600
M1629 N0545 N0540 GND GND efet w=14500 l=10150
M1630 N0570 N0540 GND GND efet w=14500 l=11600
M1631 N0584 N0540 GND GND efet w=13775 l=14500
M1632 N0599 N0613 GND GND efet w=13775 l=13775
M1633 GND N0613 N0540 GND efet w=32625 l=10875
M1634 N0620 N0613 GND GND efet w=15225 l=12325
M1635 N0635 N0613 GND GND efet w=13775 l=13775
M1636 N0648 N0613 GND GND efet w=16675 l=13050
M1637 N0613 N0646 GND GND efet w=52925 l=15225
M1638 N0539 N0541 GND GND efet w=27550 l=10150
M1639 N0545 N0541 GND GND efet w=14500 l=10875
M1640 GND N0541 N0599 GND efet w=13775 l=12325
M1641 GND N0541 N0620 GND efet w=13775 l=10875
M1642 N0570 N0577 GND GND efet w=13775 l=13775
M1643 GND N0542 N0539 GND efet w=29000 l=11600
M1644 N0584 N0577 GND GND efet w=13775 l=13775
M1645 N0503 CLK1 N0504 GND efet w=7250 l=13050
M1646 N0635 N0577 GND GND efet w=13050 l=10150
M1647 N0648 N0577 GND GND efet w=15950 l=15950
M1648 VDD VDD N0541 GND efet w=9425 l=38425
M1649 N0570 N0542 GND GND efet w=14500 l=15950
M1650 N0434 N0427 (~POC)CLK2(X12+X32)~INH GND efet w=15950 l=11600
M1651 N0426 N0427 ((~SC)(JIN+FIN))CLK1(M11+X21~INH) GND efet w=10875 l=13775
M1652 N0439 N0440 ((~SC)(JIN+FIN))CLK1(M11+X21~INH) GND efet w=11600 l=11600
M1653 N0444 N0440 (~POC)CLK2(X12+X32)~INH GND efet w=18125 l=12325
M1654 GND N0519 N0518 GND efet w=40600 l=11600
M1655 GND N0382 N0783 GND efet w=12325 l=12325
M1656 N0804 N0411 GND GND efet w=11600 l=11600
M1657 N0518 (~INH)&X32&CLK2 N0463 GND efet w=21750 l=13050
M1658 N0508 N0504 GND GND efet w=38425 l=12325
M1659 GND N0542 N0599 GND efet w=14500 l=13050
M1660 GND N0542 N0635 GND efet w=13050 l=10150
M1661 N0541 N0577 GND GND efet w=26100 l=11600
M1662 N0577 N0617 GND GND efet w=52200 l=13050
M1663 N0455 (~INH)&X32&CLK2 N0508 GND efet w=19575 l=13050
M1664 N0539 ~(FIN&X12) N0530 GND efet w=41325 l=12325
M1665 N0561 VDD VDD GND efet w=8700 l=40600
M1666 GND ~(FIN&X12) N0561 GND efet w=29000 l=11600
M1667 VDD VDD N0833 GND efet w=5800 l=60900
M1668 GND N0427 N0820 GND efet w=11600 l=10875
M1669 N0833 N0440 GND GND efet w=11600 l=11600
M1670 N0732 N0317 GND GND efet w=19575 l=12325
M1671 VDD VDD N0732 GND efet w=8700 l=65250
M1672 GND N0711 N0307 GND efet w=13775 l=11600
M1673 GND N0416 RADB0 GND efet w=43500 l=13050
M1674 RADB2 VDD VDD GND efet w=7975 l=23200
M1675 N0300 CLK2 GND GND efet w=26100 l=13050
M1676 N0307 VDD VDD GND efet w=10150 l=50750
M1677 GND CLK1 N0307 GND efet w=15950 l=10150
M1678 VDD VDD N0300 GND efet w=6525 l=29725
M1679 GND N0717 N0737 GND efet w=94250 l=13050
M1680 M12+M22+CLK1~(M11+M12) N0710 VDD GND efet w=23925 l=15225
M1681 GND N0708 M12+M22+CLK1~(M11+M12) GND efet w=20300 l=13775
M1683 S00609 VDD VDD GND efet w=7250 l=11600
M1684 GND N0708 N0710 GND efet w=14500 l=11600
M1685 N0402 VDD VDD GND efet w=7975 l=60900
M1686 GND X32 N0402 GND efet w=15950 l=10150
M1687 RADB1 VDD VDD GND efet w=7975 l=26825
M1688 RADB0 VDD VDD GND efet w=8700 l=21750
M1689 RADB1 CLK2 GND GND efet w=50750 l=11600
M1690 GND N0384 RADB1 GND efet w=42775 l=13775
M1691 RADB2 CLK2 GND GND efet w=53650 l=13050
M1692 GND N0374 RADB2 GND efet w=50025 l=11600
M1693 VDD VDD N0783 GND efet w=5800 l=62350
M1694 VDD VDD N0804 GND efet w=6525 l=50025
M1695 N0820 VDD VDD GND efet w=5800 l=52200
M1696 N0400 N0409 GND GND efet w=23925 l=10875
M1697 GND N0560 N0545 GND efet w=15225 l=10875
M1698 N0584 N0560 GND GND efet w=14500 l=11600
M1699 N0620 N0560 GND GND efet w=14500 l=10150
M1700 N0648 N0560 GND GND efet w=14500 l=12325
M1701 N0545 N0561 GND GND efet w=14500 l=13775
M1702 N0570 N0561 GND GND efet w=15225 l=13775
M1703 N0584 N0561 GND GND efet w=15225 l=12325
M1704 N0599 N0561 GND GND efet w=16675 l=11600
M1705 N0620 N0561 GND GND efet w=15225 l=10875
M1706 N0635 N0561 GND GND efet w=14500 l=11600
M1707 N0648 N0561 GND GND efet w=14500 l=13050
M1709 VDD VDD N0400 GND efet w=8700 l=65250
M1711 N0427 N0400 GND GND efet w=11600 l=13050
M1712 N0475 VDD VDD GND efet w=7250 l=65250
M1713 GND N0464 N0475 GND efet w=14500 l=13050
M1714 ADDR-PTR.1 VDD VDD GND efet w=8700 l=68150
M1715 GND N0464 ADDR-PTR.1 GND efet w=15225 l=13050
M1716 N0464 N0475 GND GND efet w=13050 l=11600
M1717 VDD VDD N0464 GND efet w=6525 l=67425
M1718 N0457 N0475 GND GND efet w=14500 l=13050
M1719 VDD VDD N0457 GND efet w=8700 l=66700
M1720 N0440 N0409 GND GND efet w=19575 l=12325
M1721 ADDR-PTR.1 N0459 N0492 GND efet w=8700 l=11600
M1722 N0457 N0459 N0458 GND efet w=9425 l=12325
M1723 N0402 CLK2 N0416 GND efet w=7250 l=13050
M1724 N0384 CLK2 N0379 GND efet w=7250 l=11600
M1725 N0374 CLK2 N0365 GND efet w=7975 l=13775
M1726 N0710 S00609 VDD GND efet w=7975 l=37700
M1727 N0379 A12 GND GND efet w=14500 l=11600
M1728 GND A22 N0365 GND efet w=15950 l=10150
M1729 VDD VDD N0365 GND efet w=9425 l=55825
M1730 VDD VDD N0708 GND efet w=8700 l=34800
M1731 N0708 CLK1 N0709 GND efet w=48575 l=15225
M1732 N0709 N0278 GND GND efet w=44225 l=12325
M1733 VDD VDD N0279 GND efet w=6525 l=41325
M1734 GND M12 N0708 GND efet w=22475 l=13050
M1735 N0708 M22 GND GND efet w=23200 l=8700
M1736 VDD VDD N0379 GND efet w=6525 l=52925
M1737 N0278 CLK2 N0279 GND efet w=14500 l=11600
M1738 GND M12 N0279 GND efet w=21025 l=12325
M1739 RADB0 CLK2 GND GND efet w=43500 l=11600
M1740 N0382 N0400 GND GND efet w=13050 l=10150
M1741 N0411 N0409 GND GND efet w=20300 l=10150
M1742 N0382 N0401 GND GND efet w=12325 l=10150
M1743 N0411 N0401 GND GND efet w=13050 l=11600
M1744 GND N0420 N0427 GND efet w=20300 l=10150
M1745 N0440 N0420 GND GND efet w=20300 l=13050
M1747 GND A32 N0279 GND efet w=23200 l=11600
M1748 VDD VDD N0304 GND efet w=7250 l=69600
M1749 N0382 S00598 VDD GND efet w=7250 l=56550
M1752 GND N0492 N0491 GND efet w=39150 l=11600
M1754 N0411 S00599 VDD GND efet w=7250 l=55100
M1755 N0427 S00600 VDD GND efet w=7250 l=56550
M1756 N0401 N0420 GND GND efet w=24650 l=11600
M1757 VDD VDD N0401 GND efet w=8700 l=66700
M1758 N0491 N0466 N0475 GND efet w=21750 l=14500
M1759 N0465 N0458 GND GND efet w=39150 l=13050
M1760 N0464 N0466 N0465 GND efet w=19575 l=13775
M1761 N0530 S00578 VDD GND efet w=10150 l=55825
M1763 N0545 S00579 VDD GND efet w=7975 l=60175
M1764 N0570 S00580 VDD GND efet w=7250 l=56550
M1769 N0584 S00581 VDD GND efet w=7250 l=56550
M1770 N0599 S00582 VDD GND efet w=8700 l=59450
M1771 N0620 S00583 VDD GND efet w=9425 l=54375
M1772 N0635 S00584 VDD GND efet w=9425 l=55825
M1773 VDD VDD N0577 GND efet w=8700 l=37700
M1774 VDD VDD N0542 GND efet w=11600 l=42775
M1776 N0542 N0560 GND GND efet w=26100 l=10150
M1777 N0560 N0582 GND GND efet w=48575 l=10875
M1778 VDD VDD N0560 GND efet w=10150 l=44225
M1779 N0648 S00585 VDD GND efet w=7250 l=53650
M1780 D1 SC&M22&CLK2 N0582 GND efet w=8700 l=13050
M1781 D2 SC&M22&CLK2 N0617 GND efet w=7250 l=13050
M1782 S00578 VDD VDD GND efet w=8700 l=11600
M1783 S00579 VDD VDD GND efet w=8700 l=12325
M1784 S00580 VDD VDD GND efet w=10150 l=10150
M1785 S00581 VDD VDD GND efet w=10150 l=10150
M1786 S00582 VDD VDD GND efet w=8700 l=10150
M1787 S00583 VDD VDD GND efet w=9425 l=10875
M1788 S00584 VDD VDD GND efet w=10875 l=14500
M1789 S00585 VDD VDD GND efet w=10150 l=11600
M1790 VDD VDD N0571 GND efet w=5800 l=68875
M1791 VDD VDD N0574 GND efet w=6525 l=65975
M1792 VDD VDD N0573 GND efet w=5800 l=66700
M1793 VDD VDD N0600 GND efet w=5800 l=63800
M1794 N0582 SC&A22 REG-RFSH.0 GND efet w=8700 l=11600
M1795 VDD VDD REG-RFSH.0 GND efet w=5800 l=33350
M1796 VDD VDD N0610 GND efet w=5800 l=72500
M1797 VDD VDD N0609 GND efet w=5800 l=63800
M1798 VDD VDD REG-RFSH.1 GND efet w=6525 l=41325
M1799 N0617 SC&A22 REG-RFSH.1 GND efet w=10875 l=10875
M1800 N0440 S00601 VDD GND efet w=7250 l=53650
M1801 N0409 X12 ADDR-RFSH.1 GND efet w=8700 l=11600
M1802 ADDR-PTR.1 X32 N0409 GND efet w=8700 l=11600
M1803 N0420 X12 ADDR-RFSH.0 GND efet w=8700 l=11600
M1804 ADDR-PTR.0 X32 N0420 GND efet w=7975 l=13050
M1806 VDD VDD N0450 GND efet w=7250 l=59450
M1807 S00598 VDD VDD GND efet w=10150 l=11600
M1808 S00599 VDD VDD GND efet w=11600 l=10150
M1809 S00600 VDD VDD GND efet w=10875 l=10150
M1810 S00601 VDD VDD GND efet w=11600 l=11600
M1811 (~POC)CLK2(X12+X32)~INH N0449 VDD GND efet w=41325 l=21025
M1812 VDD VDD S00613 GND efet w=7975 l=12325
M1813 GND JUN+JMS N0309 GND efet w=34075 l=13775
M1814 VDD S00613 N0449 GND efet w=5800 l=43500
M1815 GND N0450 (~POC)CLK2(X12+X32)~INH GND efet w=29725 l=12325
M1816 VDD VDD N0318 GND efet w=6525 l=68875
M1817 N0308 X22 N0304 GND efet w=30450 l=11600
M1818 N0309 N0310 N0308 GND efet w=30450 l=11600
M1819 N0323 M12 GND GND efet w=32625 l=12325
M1820 N0304 A32 GND GND efet w=13050 l=11600
M1821 N0323 JUN+JMS N0324 GND efet w=36975 l=20300
M1822 N0320 SC GND GND efet w=30450 l=13050
M1823 N0319 JIN+FIN N0320 GND efet w=29000 l=13050
M1824 N0318 X22 N0319 GND efet w=30450 l=11600
M1825 N0324 N0310 N0318 GND efet w=29000 l=11600
M1826 N0321 JCN+ISZ N0323 GND efet w=30450 l=11600
M1827 N0318 N0322 N0321 GND efet w=31175 l=12325
M1828 N0450 N0449 GND GND efet w=13050 l=14500
M1829 VDD VDD N0437 GND efet w=8700 l=51475
M1830 GND N0437 ((~SC)(JIN+FIN))CLK1(M11+X21~INH) GND efet w=20300 l=10150
M1831 VDD S00612 N0436 GND efet w=7250 l=40600
M1832 VDD VDD S00612 GND efet w=5800 l=10150
M1833 S00628 VDD VDD GND efet w=5800 l=11600
M1834 VDD S00628 (~INH)(X11+X31)CLK1 GND efet w=7975 l=18125
M1836 VDD N0436 ((~SC)(JIN+FIN))CLK1(M11+X21~INH) GND efet w=21025 l=12325
M1837 GND N0436 N0437 GND efet w=13775 l=13775
M1839 (~INH)(X11+X31)CLK1 N0517 GND GND efet w=35525 l=12325
M1840 GND INH (~INH)(X11+X31)CLK1 GND efet w=36250 l=11600
M1841 GND N0522 (~INH)(X11+X31)CLK1 GND efet w=34800 l=11600
M1842 VDD VDD N0451 GND efet w=5800 l=50750
M1843 N0449 INH GND GND efet w=13775 l=10875
M1844 N0436 N0443 GND GND efet w=13775 l=10875
M1845 N0436 N0435 N0441 GND efet w=29725 l=10875
M1846 N0449 POC GND GND efet w=15225 l=12325
M1847 GND N0447 N0449 GND efet w=14500 l=12325
M1848 N0449 N0451 GND GND efet w=14500 l=11600
M1849 N0441 JIN+FIN GND GND efet w=29725 l=10875
M1850 GND N0438 N0436 GND efet w=15225 l=10875
M1851 GND A22 N0318 GND efet w=18125 l=13775
M1852 N0451 CLK2 GND GND efet w=14500 l=10150
M1853 GND ~CN N0322 GND efet w=34075 l=13775
M1854 N0322 SC GND GND efet w=26825 l=13775
M1855 N0333 SC N0326 GND efet w=32625 l=10150
M1856 N0326 A12 GND GND efet w=12325 l=10875
M1857 N0334 JIN+FIN N0333 GND efet w=31900 l=10150
M1858 GND X32 N0334 GND efet w=30450 l=10150
M1859 VDD VDD N0326 GND efet w=7975 l=64525
M1860 N0341 N0310 N0339 GND efet w=36250 l=11600
M1861 N0326 JUN+JMS N0341 GND efet w=38425 l=10875
M1862 N0338 JCN+ISZ N0326 GND efet w=33350 l=11600
M1863 N0339 N0322 N0338 GND efet w=33350 l=11600
M1864 GND M22 N0339 GND efet w=34800 l=10150
M1865 GND SC N0310 GND efet w=27550 l=10875
M1866 N0310 VDD VDD GND efet w=5800 l=27550
M1867 N0322 VDD VDD GND efet w=6525 l=28275
M1868 N0344 S00654 VDD GND efet w=6525 l=28275
M1869 VDD N0344 SC GND efet w=37700 l=11600
M1870 VDD VDD S00654 GND efet w=6525 l=13050
M1871 GND X12 N0447 GND efet w=15225 l=12325
M1872 GND X32 N0447 GND efet w=12325 l=12325
M1873 VDD VDD N0443 GND efet w=6525 l=51475
M1874 N0447 VDD VDD GND efet w=5800 l=66700
M1875 N0443 CLK1 GND GND efet w=14500 l=10150
M1876 VDD VDD ~INH GND efet w=5800 l=27550
M1877 VDD VDD INH GND efet w=5800 l=29000
M1878 N0511 VDD VDD GND efet w=7975 l=54375
M1879 N0517 CLK2 N0511 GND efet w=9425 l=15225
M1880 N0466 VDD VDD GND efet w=6525 l=73225
M1881 GND N0459 N0466 GND efet w=11600 l=11600
M1882 GND N0459 ADDR-PTR.0 GND efet w=18850 l=10150
M1883 ADDR-PTR.0 VDD VDD GND efet w=7975 l=68875
M1884 N0459 N0466 GND GND efet w=13050 l=11600
M1885 VDD VDD N0459 GND efet w=6525 l=65250
M1886 N0505 N0466 GND GND efet w=14500 l=11600
M1887 VDD VDD N0505 GND efet w=9425 l=76125
M1888 N0521 CLK1 ADDR-PTR.0 GND efet w=8700 l=10875
M1889 N0505 CLK1 N0506 GND efet w=7250 l=10150
M1890 REG-RFSH.0 CLK1 N0566 GND efet w=7975 l=15225
M1891 N0571 SC&A12&CLK2 N0572 GND efet w=24650 l=12325
M1892 N0572 N0566 GND GND efet w=34075 l=12325
M1893 GND N0574 REG-RFSH.0 GND efet w=21750 l=11600
M1894 GND N0574 N0571 GND efet w=12325 l=12325
M1895 N0586 CLK1 N0573 GND efet w=7975 l=13775
M1896 N0573 N0571 GND GND efet w=12325 l=12325
M1897 N0574 N0571 GND GND efet w=12325 l=12325
M1898 REG-RFSH.1 N0571 N0593 GND efet w=10150 l=12325
M1899 GND N0521 N0520 GND efet w=39150 l=13050
M1900 VDD VDD N0494 GND efet w=7250 l=65250
M1901 (~INH)&X32&CLK2 VDD VDD GND efet w=6525 l=28275
M1902 N0520 CLK2(JMS&DC&M22+BBL(M22+X12+X22)) N0466 GND efet w=19575 l=14500
M1903 N0509 N0506 GND GND efet w=39150 l=11600
M1904 N0459 CLK2(JMS&DC&M22+BBL(M22+X12+X22)) N0509 GND efet w=20300 l=13050
M1905 GND N0592 RRAB1 GND efet w=40600 l=12325
M1906 GND N0494 (~INH)&X32&CLK2 GND efet w=26100 l=11600
M1907 VDD VDD N0522 GND efet w=5800 l=36250
M1908 CLK2(JMS&DC&M22+BBL(M22+X12+X22)) N0467 GND GND efet w=26825 l=13050
M1909 GND DC RRAB1 GND efet w=31175 l=15225
M1910 N0574 SC&A12&CLK2 N0585 GND efet w=21025 l=12325
M1911 N0625 N0571 N0609 GND efet w=8700 l=13050
M1912 GND N0600 N0609 GND efet w=13050 l=12325
M1913 N0600 N0574 N0601 GND efet w=21750 l=13050
M1914 GND N0610 REG-RFSH.1 GND efet w=21750 l=10150
M1915 N0600 N0610 GND GND efet w=11600 l=10150
M1916 N0585 N0586 GND GND efet w=35525 l=13050
M1917 N0601 N0593 GND GND efet w=33350 l=11600
M1918 RRAB1 CLK2 GND GND efet w=29000 l=13050
M1919 VDD VDD CLK2(JMS&DC&M22+BBL(M22+X12+X22)) GND efet w=9425 l=30450
M1920 GND CLK2 N0496 GND efet w=29725 l=15225
M1921 N0496 X32 N0495 GND efet w=31175 l=12325
M1922 GND INH ~INH GND efet w=26100 l=13775
M1923 GND N0524 INH GND efet w=26100 l=11600
M1924 GND M22 N0511 GND efet w=18850 l=11600
M1925 N0522 CLK1 GND GND efet w=23200 l=11600
M1926 N0495 ~INH N0494 GND efet w=29000 l=11600
M1927 N0429 X12 GND GND efet w=21750 l=13050
M1928 N0438 CLK2 N0428 GND efet w=7975 l=12325
M1929 N0428 ~INH N0429 GND efet w=21750 l=11600
M1930 N0435 SC GND GND efet w=14500 l=10875
M1931 VDD VDD N0528 GND efet w=5800 l=52200
M1932 N0428 VDD VDD GND efet w=5800 l=65250
M1933 N0428 A32 GND GND efet w=14500 l=10875
M1934 N0435 VDD VDD GND efet w=7250 l=47850
M1935 GND X22 N0511 GND efet w=15225 l=12325
M1936 GND DC N0526 GND efet w=29725 l=12325
M1937 GND ~CN N0528 GND efet w=16675 l=11600
M1938 GND SC N0525 GND efet w=21750 l=11600
M1939 N0525 JIN+FIN N0524 GND efet w=25375 l=10875
M1940 N0526 N0528 N0527 GND efet w=29725 l=12325
M1941 VDD VDD N0467 GND efet w=5800 l=63800
M1942 N0485 JMS GND GND efet w=30450 l=11600
M1943 N0484 M22 N0485 GND efet w=31900 l=11600
M1944 N0467 DC N0484 GND efet w=30450 l=11600
M1945 VDD VDD N0460 GND efet w=5800 l=33350
M1946 VDD VDD N0588 GND efet w=5800 l=70325
M1947 N0592 CLK2 N0588 GND efet w=13050 l=13050
M1948 GND CLK2 N0460 GND efet w=21750 l=11600
M1949 N0610 N0600 GND GND efet w=12325 l=10875
M1950 N0610 N0574 N0624 GND efet w=21750 l=13050
M1951 N0624 N0625 GND GND efet w=36250 l=11600
M1952 D3 SC&M22&CLK2 N0646 GND efet w=10150 l=13050
M1953 VDD VDD N0637 GND efet w=5800 l=65250
M1954 VDD VDD N0642 GND efet w=6525 l=67425
M1955 VDD VDD N0641 GND efet w=7250 l=69600
M1956 N0646 SC&A22 REG-RFSH.2 GND efet w=7250 l=11600
M1957 VDD VDD REG-RFSH.2 GND efet w=5075 l=34075
M1958 REG-RFSH.2 N0600 N0633 GND efet w=7975 l=12325
M1959 N0637 N0610 N0638 GND efet w=21025 l=12325
M1960 GND N0642 REG-RFSH.2 GND efet w=21750 l=11600
M1961 N0637 N0642 GND GND efet w=13050 l=11600
M1962 N0638 N0633 GND GND efet w=36250 l=11600
M1963 N0653 N0600 N0641 GND efet w=10875 l=15225
M1964 N0641 N0637 GND GND efet w=11600 l=10150
M1965 N0642 N0637 GND GND efet w=13050 l=11600
M1966 VDD VDD ~(FIN&X12) GND efet w=5800 l=51475
M1967 GND N0578 WRAB1 GND efet w=24650 l=11600
M1968 GND N0649 SC&A12&CLK2 GND efet w=21025 l=12325
M1970 RRAB0 DC GND GND efet w=39150 l=14500
M1971 VDD VDD N0608 GND efet w=5800 l=71050
M1972 GND N0615 RRAB0 GND efet w=36975 l=14500
M1973 GND N0460 CLK2(JMS&DC&M22+BBL(M22+X12+X22)) GND efet w=29725 l=12325
M1974 N0608 CLK2 N0615 GND efet w=16675 l=10875
M1975 N0589 X22 GND GND efet w=22475 l=12325
M1976 N0594 N0580 N0588 GND efet w=32625 l=13775
M1977 N0588 FIN+FIM+SRC+JIN N0589 GND efet w=21750 l=12325
M1978 N0595 X12 N0594 GND efet w=29725 l=13775
M1979 N0468 BBL GND GND efet w=23925 l=12325
M1980 N0527 JCN+ISZ N0524 GND efet w=29000 l=11600
M1981 N0524 JUN+JMS N0526 GND efet w=21750 l=11600
M1982 N0468 M22 N0467 GND efet w=25375 l=13775
M1983 N0467 X22 N0468 GND efet w=23200 l=11600
M1984 N0467 X12 N0468 GND efet w=21750 l=13050
M1985 GND INC+ISZ+ADD+SUB+XCH+LD N0595 GND efet w=30450 l=13050
M1986 GND CLK2 RRAB0 GND efet w=34800 l=15950
M1987 N0608 X12 N0602 GND efet w=31175 l=15225
M1988 ~(FIN&X12) X12 N0639 GND efet w=42775 l=13775
M1989 VDD VDD DC GND efet w=8700 l=24650
M1990 WRAB1 VDD VDD GND efet w=5800 l=33350
M1991 N0547 VDD VDD GND efet w=5800 l=69600
M1992 VDD VDD WRAB0 GND efet w=7250 l=29000
M1993 SC&A12&CLK2 VDD VDD GND efet w=5800 l=36250
M1994 SC(A22+M22)CLK2 S00624 VDD GND efet w=10150 l=27550
M1995 SC(A22+M22)CLK2 N0655 GND GND efet w=37700 l=14500
M1996 N0642 N0610 N0652 GND efet w=24650 l=15950
M1997 N0652 N0653 GND GND efet w=33350 l=11600
M1998 GND N0622 N0621 GND efet w=12325 l=12325
M2000 VDD S00620 N0621 GND efet w=6525 l=54375
M2001 GND N0622 CLK2&SC(A12+M12) GND efet w=20300 l=11600
M2002 GND N0626 N0627 GND efet w=11600 l=11600
M2004 CLK2&SC(A12+M12) N0621 VDD GND efet w=18850 l=11600
M2005 (~POC)&CLK2&SC(A32+X12) N0627 GND GND efet w=24650 l=11600
M2006 S00624 VDD VDD GND efet w=6525 l=10875
M2007 WRAB0 N0547 GND GND efet w=33350 l=13775
M2008 N0602 ~OPA.0 N0614 GND efet w=52925 l=12325
M2009 N0640 ~OPA.0 N0639 GND efet w=80475 l=13050
M2010 GND N0636 N0640 GND efet w=42775 l=13775
M2011 GND INC+ISZ+ADD+SUB+XCH+LD N0614 GND efet w=29725 l=12325
M2012 GND SC N0612 GND efet w=29725 l=13775
M2013 DC SC GND GND efet w=60175 l=13050
M2014 GND FIN+FIM+SRC+JIN N0602 GND efet w=21750 l=10150
M2015 N0580 ~OPA.0 GND GND efet w=55100 l=11600
M2016 GND DC N0597 GND efet w=30450 l=11600
M2017 N0597 FIN+FIM+SRC+JIN N0596 GND efet w=31175 l=10875
M2018 N0649 VDD VDD GND efet w=5800 l=71050
M2019 VDD VDD N0655 GND efet w=5800 l=71050
M2020 S00620 VDD VDD GND efet w=7250 l=11600
M2021 N0655 CLK2 N0656 GND efet w=30450 l=10150
M2022 N0649 CLK2 N0650 GND efet w=30450 l=11600
M2023 N0626 S00627 VDD GND efet w=5800 l=52200
M2024 N0612 X32 N0611 GND efet w=36975 l=12325
M2025 N0564 N0590 GND GND efet w=29725 l=14500
M2026 N0524 VDD VDD GND efet w=5800 l=60900
M2027 GND ~OPR.3 IO GND efet w=31900 l=12325
M2028 OPE ~OPR.3 GND GND efet w=32625 l=10875
M2029 GND DC INC/ISZ GND efet w=24650 l=11600
M2030 N0580 VDD VDD GND efet w=5800 l=27550
M2031 GND N0603 N0568 GND efet w=28275 l=14500
M2032 N0596 ~OPA.0 N0590 GND efet w=54375 l=12325
M2033 N0568 VDD VDD GND efet w=5800 l=27550
M2034 N0563 N0564 N0562 GND efet w=34075 l=15950
M2035 GND M12 N0563 GND efet w=34075 l=13050
M2036 N0576 M22 GND GND efet w=31175 l=13775
M2037 N0575 N0564 N0576 GND efet w=30450 l=13050
M2038 N0562 CLK2 N0547 GND efet w=34075 l=12325
M2039 N0567 ~OPA.0 N0562 GND efet w=53650 l=13775
M2040 N0603 INC+ISZ+XCH N0611 GND efet w=31175 l=12325
M2041 VDD VDD N0603 GND efet w=6525 l=64525
M2042 N0564 VDD VDD GND efet w=5800 l=27550
M2043 N0579 N0568 GND GND efet w=31175 l=13775
M2044 GND N0568 N0567 GND efet w=30450 l=13050
M2045 N0575 N0580 N0579 GND efet w=30450 l=13050
M2046 N0654 SC N0656 GND efet w=32625 l=15225
M2047 N0651 A12 N0650 GND efet w=32625 l=13775
M2048 GND SC N0651 GND efet w=30450 l=14500
M2049 GND M22 N0654 GND efet w=31175 l=15225
M2050 VDD VDD N0622 GND efet w=7250 l=68150
M2051 S00627 VDD VDD GND efet w=6525 l=10875
M2052 VDD VDD N0627 GND efet w=5800 l=52200
M2053 N0622 CLK2 N0623 GND efet w=36975 l=10875
M2054 GND M12 N0618 GND efet w=30450 l=11600
M2055 N0682 X12 N0683 GND efet w=84825 l=16675
M2056 N0618 A12 GND GND efet w=36250 l=15225
M2057 GND A22 N0654 GND efet w=29725 l=13775
M2058 N0578 CLK2 N0575 GND efet w=31900 l=13050
M2059 VDD VDD N0578 GND efet w=7975 l=67425
M2060 N0590 VDD VDD GND efet w=5800 l=65250
M2061 N0618 SC N0623 GND efet w=34075 l=15225
M2062 GND POC N0683 GND efet w=86275 l=12325
M2063 VDD VDD SC&A22 GND efet w=5800 l=34800
M2064 (~POC)&CLK2&SC(A32+X12) N0626 VDD GND efet w=21750 l=10150
M2065 VDD VDD N0679 GND efet w=9425 l=65975
M2066 VDD VDD SC&M22&CLK2 GND efet w=7975 l=25375
M2067 SC&M22&CLK2 N0679 GND GND efet w=37700 l=14500
M2068 N0626 N0630 GND GND efet w=13775 l=10875
M2069 GND POC N0626 GND efet w=16675 l=12325
M2070 N0679 M22 N0680 GND efet w=32625 l=12325
M2071 GND N0643 SC&A22 GND efet w=25375 l=15225
M2072 N0703 CLK2 N0682 GND efet w=14500 l=13050
M2073 N0681 CLK2 N0680 GND efet w=30450 l=11600
M2074 N0681 SC GND GND efet w=30450 l=11600
M2075 N0629 X12 GND GND efet w=31175 l=12325
M2076 XCH ~OPR.3 GND GND efet w=30450 l=15225
M2077 GND ~OPR.3 BBL GND efet w=30450 l=13050
M2078 N0628 ~OPR.3 GND GND efet w=53650 l=11600
M2079 INC+ISZ+XCH ~OPR.3 N0587 GND efet w=47850 l=11600
M2080 LD ~OPR.3 GND GND efet w=31175 l=11600
M2081 SUB ~OPR.3 GND GND efet w=30450 l=10875
M2082 ADD ~OPR.3 GND GND efet w=31175 l=13050
M2083 JCN+ISZ OPR.3 GND GND efet w=50025 l=11600
M2084 GND OPR.3 JCN GND efet w=25375 l=13050
M2085 FIN+FIM OPR.3 GND GND efet w=23925 l=13775
M2086 N0361 VDD VDD GND efet w=6525 l=35525
M2088 GND N0343 SC GND efet w=30450 l=11600
M2089 N0344 N0343 GND GND efet w=29000 l=11600
M2090 GND OPR.3 ISZ GND efet w=24650 l=11600
M2091 GND OPR.3 FIM+SRC GND efet w=23925 l=12325
M2092 GND OPR.3 JIN+FIN GND efet w=44950 l=11600
M2093 JUN+JMS OPR.3 GND GND efet w=44225 l=11600
M2094 GND OPR.3 INC/ISZ GND efet w=23200 l=13050
M2095 ISZ ~OPR.2 GND GND efet w=31175 l=11600
M2096 IO ~OPR.2 GND GND efet w=29725 l=12325
M2097 OPE ~OPR.2 GND GND efet w=31175 l=11600
M2098 JUN+JMS ~OPR.2 GND GND efet w=55825 l=13775
M2099 GND OPR.3 JMS GND efet w=24650 l=11600
M2100 GND OPR.3 N0636 GND efet w=23200 l=11600
M2101 LDM/BBL ~OPR.3 GND GND efet w=31900 l=13050
M2102 GND A32 N0629 GND efet w=29725 l=13775
M2103 N0629 SC N0631 GND efet w=34075 l=13775
M2104 GND IOR N0683 GND efet w=81925 l=12325
M2105 GND A32 N0682 GND efet w=51475 l=15225
M2106 N0682 M12 GND GND efet w=36975 l=13775
M2107 GND N0703 L GND efet w=52925 l=13775
M2108 L N0703 GND GND efet w=60900 l=14500
M2109 N0631 CLK2 N0630 GND efet w=30450 l=8700
M2110 GND M12 N0662 GND efet w=29725 l=10875
M2111 N0662 SC N0661 GND efet w=29725 l=10875
M2112 N0644 A22 N0643 GND efet w=23925 l=9425
M2113 GND SC N0644 GND efet w=23200 l=11600
M2114 N0661 CLK2 N0660 GND efet w=30450 l=10150
M2115 N0682 VDD VDD GND efet w=9425 l=35525
M2116 VDD VDD N0630 GND efet w=6525 l=64525
M2117 INC+ISZ+ADD+SUB+XCH+LD OPR.3 N0628 GND efet w=47850 l=13050
M2118 N0587 OPR.3 GND GND efet w=39875 l=13775
M2119 GND ~OPR.2 N0523 GND efet w=92075 l=10875
M2120 INC/ISZ ~OPR.2 GND GND efet w=30450 l=12325
M2121 BBL ~OPR.2 GND GND efet w=30450 l=12325
M2122 N0373 JCN+ISZ N0372 GND efet w=36250 l=15950
M2123 N0372 FIN+FIM N0373 GND efet w=33350 l=14500
M2124 JMS ~OPR.2 GND GND efet w=31900 l=11600
M2125 GND OPR.3 FIN+FIM+SRC+JIN GND efet w=24650 l=11600
M2126 GND OPR.3 JUN2+JMS2 GND efet w=24650 l=11600
M2127 N0628 ~OPR.2 INC+ISZ+ADD+SUB+XCH+LD GND efet w=56550 l=11600
M2128 N0587 ~OPR.2 GND GND efet w=46400 l=13775
M2129 LDM/BBL ~OPR.2 GND GND efet w=32625 l=12325
M2130 N0523 OPR.2 JCN+ISZ GND efet w=98600 l=11600
M2131 GND OPR.2 FIN+FIM GND efet w=23200 l=11600
M2132 GND OPR.2 JCN GND efet w=23925 l=13775
M2133 FIM+SRC OPR.2 GND GND efet w=23200 l=11600
M2134 JUN2+JMS2 ~OPR.2 GND GND efet w=32625 l=12325
M2135 GND OPR.2 JIN+FIN GND efet w=44950 l=10150
M2136 FIN+FIM ~OPR.1 GND GND efet w=31175 l=12325
M2137 ISZ ~OPR.1 GND GND efet w=31900 l=13050
M2138 GND OPR.2 XCH GND efet w=23200 l=11600
M2139 GND OPR.2 N0636 GND efet w=23925 l=12325
M2140 N0628 OPR.2 GND GND efet w=46400 l=15950
M2141 OPR.2 N0995 VDD GND efet w=47850 l=20300
M2142 VDD N0994 ~OPR.2 GND efet w=33350 l=15950
M2143 N0587 OPR.2 INC+ISZ+XCH GND efet w=40600 l=13050
M2144 GND OPR.2 FIN+FIM+SRC+JIN GND efet w=25375 l=12325
M2145 FIM+SRC ~OPR.1 GND GND efet w=29725 l=11600
M2146 IO ~OPR.1 GND GND efet w=29725 l=11600
M2147 OPE ~OPR.1 GND GND efet w=30450 l=12325
M2148 JIN+FIN ~OPR.1 GND GND efet w=53650 l=11600
M2149 INC/ISZ ~OPR.1 GND GND efet w=29725 l=10875
M2150 N0523 ~OPR.1 GND GND efet w=89175 l=13050
M2151 XCH ~OPR.1 GND GND efet w=30450 l=12325
M2152 GND OPR.2 LD GND efet w=24650 l=11600
M2153 GND OPR.2 SUB GND efet w=23200 l=12325
M2154 GND OPR.2 ADD GND efet w=23200 l=11600
M2155 N0628 ~OPR.1 INC+ISZ+ADD+SUB+XCH+LD GND efet w=57275 l=14500
M2156 GND ~OPR.1 N0587 GND efet w=45675 l=11600
M2157 N0361 CLK1 N0343 GND efet w=14500 l=13050
M2158 N0372 X32 GND GND efet w=37700 l=13050
M2159 N0352 VDD VDD GND efet w=7975 l=64525
M2160 GND N0362 N0361 GND efet w=22475 l=10875
M2161 N0373 JUN+JMS N0372 GND efet w=31900 l=13050
M2162 N0368 SC N0373 GND efet w=34800 l=11600
M2163 GND OPR.1 JCN GND efet w=23925 l=12325
M2164 GND OPR.1 JUN+JMS GND efet w=46400 l=13050
M2165 N0636 ~OPR.1 GND GND efet w=23200 l=10150
M2166 N0523 OPR.1 JCN+ISZ GND efet w=96425 l=14500
M2167 GND OPR.1 BBL GND efet w=23200 l=11600
M2168 GND OPR.1 JMS GND efet w=26100 l=11600
M2169 INC+ISZ+XCH ~OPR.1 N0587 GND efet w=46400 l=13050
M2170 FIN+FIM+SRC+JIN ~OPR.1 GND GND efet w=30450 l=12325
M2171 LD ~OPR.1 GND GND efet w=31900 l=11600
M2172 GND N0995 ~OPR.2 GND efet w=32625 l=13775
M2173 OPR.2 N0994 GND GND efet w=29725 l=13775
M2174 L VDD VDD GND efet w=10150 l=14500
M2175 OPR.3 N0993 VDD GND efet w=39150 l=14500
M2176 VDD N0992 ~OPR.3 GND efet w=20300 l=14500
M2177 VDD VDD N0643 GND efet w=7250 l=60900
M2178 N0660 VDD VDD GND efet w=6525 l=63075
M2179 GND N0660 SC&M12&CLK2 GND efet w=36975 l=9425
M2180 SC&M12&CLK2 VDD VDD GND efet w=6525 l=26100
M2181 D0 SC&M12&CLK2 N1011 GND efet w=11600 l=12325
M2182 D2 SC&M12&CLK2 N1009 GND efet w=10875 l=11600
M2183 OPR.3 N0992 GND GND efet w=29725 l=15225
M2184 GND N0993 ~OPR.3 GND efet w=20300 l=11600
M2185 N0998 VDD VDD GND efet w=8700 l=30450
M2186 N0994 VDD VDD GND efet w=10150 l=32625
M2187 GND N1011 N0998 GND efet w=58725 l=13775
M2188 GND N1008 N0992 GND efet w=62350 l=11600
M2189 D1 SC&M12&CLK2 N1010 GND efet w=10875 l=12325
M2190 N0996 VDD VDD GND efet w=12325 l=29000
M2191 GND N1009 N0994 GND efet w=61625 l=12325
M2192 N0992 VDD VDD GND efet w=8700 l=33350
M2193 GND OPR.1 SUB GND efet w=23925 l=10875
M2194 GND OPR.1 ADD GND efet w=23925 l=10875
M2195 LDM/BBL OPR.1 GND GND efet w=23925 l=12325
M2196 ISZ ~OPR.0 GND GND efet w=31900 l=13050
M2197 JCN ~OPR.0 GND GND efet w=31175 l=12325
M2198 OPE ~OPR.0 GND GND efet w=30450 l=12325
M2199 JIN+FIN ~OPR.0 GND GND efet w=52200 l=10875
M2200 GND X32 N0352 GND efet w=12325 l=12325
M2201 N0367 N0352 GND GND efet w=21750 l=11600
M2202 N0368 N0343 N0367 GND efet w=21750 l=11600
M2203 N0362 CLK2 N0368 GND efet w=8700 l=11600
M2204 VDD VDD N0368 GND efet w=6525 l=67425
M2205 XCH ~OPR.0 GND GND efet w=29725 l=10875
M2206 GND ~OPR.0 JCN+ISZ GND efet w=53650 l=11600
M2207 JMS ~OPR.0 GND GND efet w=31175 l=10150
M2208 GND OPR.1 JUN2+JMS2 GND efet w=24650 l=11600
M2209 INC+ISZ+XCH ~OPR.0 N0587 GND efet w=52200 l=13050
M2210 N0636 ~OPR.0 GND GND efet w=23925 l=12325
M2211 SUB ~OPR.0 GND GND efet w=31175 l=12325
M2212 VDD N0998 ~OPR.0 GND efet w=39875 l=21750
M2213 GND OPA.0 FIN+FIM GND efet w=21750 l=14500
M2214 GND OPR.0 FIM+SRC GND efet w=25375 l=15225
M2215 GND OPR.0 IO GND efet w=23200 l=11600
M2216 VDD VDD N0769 GND efet w=6525 l=39875
M2217 POC VDD VDD GND efet w=7975 l=22475
M2218 ~CN VDD VDD GND efet w=10150 l=28275
M2219 N0769 A12 GND GND efet w=18125 l=12325
M2220 FIN+FIM VDD VDD GND efet w=5800 l=59450
M2221 GND OPR.0 BBL GND efet w=23200 l=11600
M2222 OPR.0 N0999 VDD GND efet w=20300 l=17400
M2223 GND OPR.0 LD GND efet w=24650 l=10150
M2224 GND OPR.0 ADD GND efet w=23200 l=12325
M2225 ISZ VDD VDD GND efet w=7250 l=63800
M2226 JCN VDD VDD GND efet w=5800 l=62350
M2227 FIM+SRC VDD VDD GND efet w=5800 l=63075
M2228 IO VDD VDD GND efet w=9425 l=73225
M2229 N0493 VDD VDD GND efet w=7250 l=72500
M2230 VDD VDD OPE GND efet w=7250 l=56550
M2231 JIN+FIN VDD VDD GND efet w=7250 l=36975
M2232 VDD VDD N0510 GND efet w=7250 l=50750
M2233 JUN+JMS VDD VDD GND efet w=8700 l=39150
M2234 JCN+ISZ VDD VDD GND efet w=8700 l=34800
M2235 INC/ISZ VDD VDD GND efet w=7250 l=55100
M2236 VDD VDD DCL GND efet w=5800 l=63800
M2237 GND OPA.0 N0516 GND efet w=38425 l=10875
M2238 N0516 FIM+SRC ~SRC GND efet w=23200 l=13050
M2239 GND SC N0417 GND efet w=33350 l=10150
M2240 GND POC_PAD N0327 GND efet w=35525 l=12325
M2241 GND N0397 ~CN GND efet w=57275 l=13050
M2242 GND N0327 N0769 GND efet w=19575 l=12325
M2243 POC N0327 GND GND efet w=55825 l=12325
M2244 N0412 N0397 GND GND efet w=21750 l=13050
M2245 N0399 X32 GND GND efet w=13775 l=12325
M2246 N0417 X32 N0418 GND efet w=34075 l=10875
M2247 GND IO N0493 GND efet w=13775 l=11600
M2248 N0510 OPE GND GND efet w=15225 l=12325
M2249 VDD N0510 ~OPE GND efet w=29000 l=11600
M2250 GND IO ~I/O GND efet w=34800 l=11600
M2251 ~I/O N0493 VDD GND efet w=13775 l=12325
M2252 GND ISZ N0456 GND efet w=13050 l=11600
M2253 GND JCN N0476 GND efet w=13775 l=12325
M2254 ~OPE OPE GND GND efet w=29725 l=12325
M2255 VDD VDD O-IB GND efet w=7250 l=53650
M2256 VDD VDD KBP GND efet w=5800 l=65975
M2257 VDD VDD TCS GND efet w=8700 l=43500
M2258 VDD VDD DAA GND efet w=8700 l=43500
M2259 XCH VDD VDD GND efet w=5800 l=57275
M2260 BBL VDD VDD GND efet w=6525 l=57275
M2261 JMS VDD VDD GND efet w=7250 l=55100
M2262 N0636 VDD VDD GND efet w=6525 l=60900
M2263 INC+ISZ+ADD+SUB+XCH+LD VDD VDD GND efet w=10150 l=65250
M2264 VDD VDD IOW GND efet w=5800 l=56550
M2265 VDD VDD RAR GND efet w=7250 l=55100
M2266 RAL VDD VDD GND efet w=6525 l=55100
M2267 CMA VDD VDD GND efet w=6525 l=55825
M2268 VDD VDD TCC GND efet w=7250 l=56550
M2269 STC VDD VDD GND efet w=5800 l=61625
M2270 INC+ISZ+XCH VDD VDD GND efet w=5800 l=65250
M2271 LD VDD VDD GND efet w=6525 l=67425
M2272 FIN+FIM+SRC+JIN VDD VDD GND efet w=7250 l=50750
M2273 IOW ~I/O GND GND efet w=38425 l=10875
M2274 VDD VDD CMC GND efet w=7250 l=53650
M2275 VDD VDD DAC GND efet w=6525 l=52925
M2276 VDD VDD IAC GND efet w=5800 l=56550
M2277 VDD VDD CLC GND efet w=7250 l=63075
M2278 SUB VDD VDD GND efet w=7250 l=60900
M2279 ADD VDD VDD GND efet w=7250 l=59450
M2280 LDM/BBL VDD VDD GND efet w=7975 l=58725
M2281 JUN2+JMS2 VDD VDD GND efet w=7250 l=63800
M2282 VDD VDD CLB GND efet w=7975 l=65250
M2283 VDD VDD SBM GND efet w=7250 l=56550
M2284 ADM VDD VDD GND efet w=5800 l=56550
M2285 OPR.0 N0998 GND GND efet w=21025 l=12325
M2286 GND N0999 ~OPR.0 GND efet w=29725 l=12325
M2287 ~OPR.1 N0996 VDD GND efet w=38425 l=15950
M2288 VDD N0997 OPR.1 GND efet w=24650 l=13050
M2289 N0999 N0998 GND GND efet w=27550 l=11600
M2290 GND N1010 N0996 GND efet w=58000 l=11600
M2291 N0995 N0994 GND GND efet w=29000 l=11600
M2292 N0997 N0996 GND GND efet w=29000 l=10150
M2293 D3 SC&M12&CLK2 N1008 GND efet w=10150 l=12325
M2294 N0993 N0992 GND GND efet w=26825 l=10875
M2295 N0999 VDD VDD GND efet w=13050 l=42050
M2296 ~OPR.1 N0997 GND GND efet w=34075 l=13050
M2297 GND N0996 OPR.1 GND efet w=24650 l=11600
M2298 N0995 VDD VDD GND efet w=14500 l=43500
M2299 N0997 VDD VDD GND efet w=9425 l=36975
M2300 N0993 VDD VDD GND efet w=15950 l=38425
M2301 D3 OPA-IB OPA.3 GND efet w=58725 l=13775
M2302 VDD VDD IOR GND efet w=10875 l=41325
M2303 SBM ~I/O GND GND efet w=31900 l=13050
M2304 ADM ~I/O GND GND efet w=31900 l=12325
M2305 VDD VDD N0477 GND efet w=5800 l=49300
M2306 GND ~(X31&~CLK2) N0480 GND efet w=13775 l=12325
M2307 N0480 VDD VDD GND efet w=7250 l=67425
M2308 N0482 N0480 N0477 GND efet w=27550 l=11600
M2309 N0479 VDD VDD GND efet w=7250 l=77575
M2310 N0482 N0479 GND GND efet w=26825 l=10875
M2311 N0479 IOR GND GND efet w=12325 l=10150
M2312 N0412 N0399 N0413 GND efet w=20300 l=11600
M2313 N0418 N0419 N0413 GND efet w=30450 l=10150
M2314 GND N0769 N0327 GND efet w=33350 l=11600
M2315 N0297 CLK2 GND GND efet w=26100 l=11600
M2317 X22 CLK2 N0280 GND efet w=13775 l=12325
M2318 VDD S00678 N0297 GND efet w=7975 l=32625
M2319 VDD VDD S00678 GND efet w=5800 l=13050
M2320 N0295 N0297 N0296 GND efet w=27550 l=11600
M2321 N0296 N0280 GND GND efet w=62350 l=13050
M2322 VDD VDD N0296 GND efet w=7975 l=21025
M2323 N0739 CLK1 N0296 GND efet w=11600 l=11600
M2324 N0404 CLK1 N0397 GND efet w=14500 l=11600
M2325 GND N0405 N0404 GND efet w=26825 l=12325
M2326 N0413 CLK2 N0405 GND efet w=8700 l=11600
M2327 VDD VDD N0399 GND efet w=7250 l=84100
M2328 GND TEST_PAD N0432 GND efet w=36250 l=10150
M2329 VDD VDD N0432 GND efet w=7250 l=55100
M2330 N0327 VDD VDD GND efet w=5800 l=26100
M2331 VDD VDD N0404 GND efet w=7250 l=36250
M2332 VDD VDD N0784 GND efet w=5800 l=50750
M2333 N0741 N0739 GND GND efet w=31900 l=10875
M2334 VDD VDD N0329 GND efet w=8700 l=20300
M2335 N0413 VDD VDD GND efet w=6525 l=63075
M2336 N0456 VDD VDD GND efet w=10875 l=65975
M2337 GND N0476 N0478 GND efet w=23200 l=11600
M2338 GND ~OPE DCL GND efet w=23200 l=11600
M2339 O-IB ~OPE GND GND efet w=23200 l=12325
M2340 GND ~OPE KBP GND efet w=23925 l=12325
M2341 GND ~OPE TCS GND efet w=38425 l=10875
M2342 DAA ~OPE GND GND efet w=34075 l=12325
M2343 RAR ~OPE GND GND efet w=23925 l=10875
M2344 GND ~OPE RAL GND efet w=23925 l=10875
M2345 GND ~OPE CMA GND efet w=25375 l=10875
M2346 N0478 N0487 N0481 GND efet w=44225 l=15225
M2347 N0478 ~OPA.3 N0481 GND efet w=63800 l=13050
M2348 N0478 N0456 N0419 GND efet w=41325 l=13775
M2349 GND ~I/O N0329 GND efet w=59450 l=11600
M2350 N0476 VDD VDD GND efet w=5800 l=58000
M2351 N0478 ADD_0 N0419 GND efet w=47125 l=13050
M2352 N0419 VDD VDD GND efet w=5800 l=50025
M2353 VDD VDD ~SRC GND efet w=5800 l=68875
M2354 DCL ~OPA.3 GND GND efet w=30450 l=10875
M2355 KBP ~OPA.3 GND GND efet w=30450 l=11600
M2356 TCS ~OPA.3 GND GND efet w=40600 l=11600
M2357 DAA ~OPA.3 GND GND efet w=40600 l=13775
M2358 GND N0486 N0481 GND efet w=50750 l=14500
M2359 GND OPA.3 N0481 GND efet w=75400 l=13050
M2360 GND ~OPE TCC GND efet w=23200 l=11600
M2361 STC ~OPE GND GND efet w=23925 l=12325
M2362 GND ~OPE CMC GND efet w=23925 l=12325
M2363 GND ~OPE DAC GND efet w=23200 l=13050
M2364 GND ~OPE IAC GND efet w=23925 l=12325
M2365 GND ~I/O IOR GND efet w=39875 l=10875
M2366 N0477 A12 N0483 GND efet w=31900 l=11600
M2367 D2 OPA-IB OPA.2 GND efet w=61625 l=16675
M2368 GND IOR N0483 GND efet w=31175 l=15225
M2369 GND ~OPE CLC GND efet w=23200 l=10150
M2370 CLB ~OPE GND GND efet w=23200 l=11600
M2371 STC ~OPA.3 GND GND efet w=31175 l=13050
M2372 DAC ~OPA.3 GND GND efet w=30450 l=10875
M2373 SBM ~OPA.3 GND GND efet w=32625 l=11600
M2374 ADM ~OPA.3 GND GND efet w=30450 l=13775
M2375 IOR ~OPA.3 GND GND efet w=44950 l=11600
M2376 GND N1001 ~OPA.3 GND efet w=29725 l=11600
M2377 OPA.3 N1000 GND GND efet w=57275 l=12325
M2378 GND OPA.3 O-IB GND efet w=23200 l=12325
M2379 GND OPA.3 IOW GND efet w=31900 l=10150
M2380 GND OPA.3 RAR GND efet w=24650 l=10150
M2381 GND OPA.3 RAL GND efet w=23925 l=10875
M2382 GND OPA.3 CMA GND efet w=23200 l=10150
M2383 GND OPA.3 TCC GND efet w=23200 l=10150
M2384 GND OPA.3 CMC GND efet w=24650 l=11600
M2385 GND OPA.3 IAC GND efet w=23925 l=10875
M2386 GND N0486 N0487 GND efet w=13050 l=11600
M2387 DCL ~OPA.2 GND GND efet w=30450 l=10875
M2388 GND OPA.2 N0501 GND efet w=44950 l=14500
M2389 N0501 ACC_0 N0486 GND efet w=29000 l=10875
M2390 N0487 VDD VDD GND efet w=5800 l=50750
M2391 VDD VDD N0398 GND efet w=6525 l=26100
M2392 KBP ~OPA.2 GND GND efet w=30450 l=10875
M2393 RAR ~OPA.2 GND GND efet w=31900 l=12325
M2394 RAL ~OPA.2 GND GND efet w=31175 l=13050
M2395 GND OPA.3 CLC GND efet w=23200 l=11600
M2396 GND OPA.3 CLB GND efet w=24650 l=11600
M2397 CMA ~OPA.2 GND GND efet w=30450 l=11600
M2398 TCC ~OPA.2 GND GND efet w=31175 l=11600
M2399 N0486 VDD VDD GND efet w=5800 l=47850
M2400 GND OPA.2 TCS GND efet w=34075 l=13775
M2401 GND OPA.2 DAA GND efet w=34800 l=11600
M2402 GND N1003 ~OPA.2 GND efet w=36975 l=15225
M2403 OPA.2 N1002 GND GND efet w=54375 l=15950
M2404 VDD N1000 ~OPA.3 GND efet w=22475 l=10875
M2405 OPA.3 N1001 VDD GND efet w=25375 l=9425
M2406 GND OPA.2 STC GND efet w=23200 l=10150
M2407 GND OPA.2 CMC GND efet w=24650 l=10150
M2408 GND OPA.2 DAC GND efet w=23925 l=11600
M2409 GND OPA.2 IAC GND efet w=27550 l=10150
M2410 GND OPA.2 CLC GND efet w=27550 l=10150
M2411 CLB OPA.2 GND GND efet w=23200 l=13050
M2412 DAA ~OPA.1 GND GND efet w=43500 l=10875
M2413 GND CLK2 N0398 GND efet w=47850 l=10150
M2414 VDD VDD N0799 GND efet w=6525 l=67425
M2416 VDD S00690 N0741 GND efet w=6525 l=26825
M2417 VDD VDD S00690 GND efet w=5800 l=13050
M2418 X32 N0739 GND GND efet w=31900 l=11600
M2419 GND N0782 N0784 GND efet w=14500 l=11600
M2420 VDD N0741 X32 GND efet w=36250 l=12325
M2421 N0414 CLK2 A22 GND efet w=8700 l=11600
M2422 N0799 ~SRC GND GND efet w=13050 l=13050
M2423 N0407 N0414 GND GND efet w=14500 l=11600
M2424 N0407 N0398 N0408 GND efet w=8700 l=13050
M2425 VDD VDD S00685 GND efet w=6525 l=11600
M2426 VDD S00685 N0415 GND efet w=5800 l=16675
M2428 N0507 CY_1 N0486 GND efet w=27550 l=11600
M2429 RAR ~OPA.1 GND GND efet w=31175 l=10150
M2430 TCC ~OPA.1 GND GND efet w=30450 l=11600
M2431 GND OPA.1 N0507 GND efet w=45675 l=13050
M2432 STC ~OPA.1 GND GND efet w=31900 l=11600
M2433 CMC ~OPA.1 GND GND efet w=31175 l=12325
M2434 IAC ~OPA.1 GND GND efet w=31900 l=11600
M2435 GND OPA.2 SBM GND efet w=28275 l=10875
M2436 GND OPA.2 ADM GND efet w=26100 l=11600
M2437 ADM ~OPA.1 GND GND efet w=29725 l=12325
M2438 ~COM N0782 VDD GND efet w=20300 l=11600
M2439 GND N0784 ~COM GND efet w=20300 l=11600
M2440 N0800 N0801 N0782 GND efet w=30450 l=10150
M2441 GND N0329 N0800 GND efet w=27550 l=11600
M2442 N0798 N0805 GND GND efet w=27550 l=11600
M2443 N0782 N0799 N0798 GND efet w=29725 l=12325
M2444 GND N0797 N0782 GND efet w=15225 l=12325
M2445 GND CLK2 N0375 GND efet w=16675 l=12325
M2446 N0797 N0408 GND GND efet w=20300 l=12325
M2447 VDD VDD N0797 GND efet w=7975 l=55100
M2448 VDD N0742 X22 GND efet w=39150 l=13050
M2449 X22 N0719 GND GND efet w=36975 l=12325
M2450 GND X22 N0288 GND efet w=25375 l=13775
M2451 N0742 N0719 GND GND efet w=30450 l=11600
M2453 VDD VDD S00710 GND efet w=6525 l=13775
M2454 VDD S00710 N0742 GND efet w=7250 l=27550
M2455 N0718 N0281 GND GND efet w=26825 l=10875
M2456 N0281 CLK2 X12 GND efet w=13050 l=13775
M2457 N0719 CLK1 N0718 GND efet w=14500 l=11600
M2458 VDD VDD N0718 GND efet w=8700 l=37700
M2459 N0383 X22 GND GND efet w=14500 l=11600
M2461 N0288 X12 GND GND efet w=21750 l=13775
M2462 VDD N0743 X12 GND efet w=35525 l=12325
M2463 X12 N0721 GND GND efet w=36975 l=12325
M2465 N0743 N0721 GND GND efet w=26100 l=10875
M2466 VDD VDD S00725 GND efet w=5800 l=11600
M2467 VDD S00725 N0743 GND efet w=7975 l=26825
M2468 VDD S00699 N0782 GND efet w=5800 l=39875
M2469 N0380 CLK2 N0383 GND efet w=8700 l=11600
M2470 VDD VDD N0407 GND efet w=5800 l=49300
M2471 GND OPA.1 DCL GND efet w=24650 l=13050
M2472 GND OPA.1 KBP GND efet w=29000 l=11600
M2473 GND OPA.1 TCS GND efet w=33350 l=11600
M2474 GND OPA.1 RAL GND efet w=23925 l=12325
M2475 GND OPA.1 CMA GND efet w=24650 l=10875
M2476 GND OPA.1 DAC GND efet w=23200 l=10150
M2477 GND OPA.1 CLC GND efet w=23200 l=10150
M2478 GND OPA.1 CLB GND efet w=24650 l=13050
M2479 GND OPA.1 SBM GND efet w=23925 l=13050
M2480 N0512 N0432 N0486 GND efet w=27550 l=11600
M2481 GND OPA.0 N0512 GND efet w=49300 l=14500
M2482 DCL ~OPA.0 GND GND efet w=30450 l=11600
M2483 TCS ~OPA.0 GND GND efet w=42050 l=10875
M2484 DAA ~OPA.0 GND GND efet w=41325 l=11600
M2485 RAL ~OPA.0 GND GND efet w=31175 l=13775
M2486 TCC ~OPA.0 GND GND efet w=30450 l=11600
M2487 CMC ~OPA.0 GND GND efet w=31900 l=11600
M2488 CLC ~OPA.0 GND GND efet w=31175 l=10150
M2489 ADM ~OPA.0 GND GND efet w=29725 l=11600
M2490 GND OPA.0 KBP GND efet w=24650 l=10150
M2491 GND OPA.0 RAR GND efet w=24650 l=11600
M2492 GND OPA.0 DAC GND efet w=26100 l=13050
M2493 VDD N1002 ~OPA.2 GND efet w=14500 l=11600
M2494 OPA.1 N1004 GND GND efet w=68875 l=12325
M2495 GND OPA.0 CMA GND efet w=23200 l=11600
M2496 GND OPA.0 STC GND efet w=23200 l=10875
M2497 GND OPA.0 IAC GND efet w=23200 l=10150
M2498 GND OPA.0 CLB GND efet w=24650 l=11600
M2499 GND OPA.0 SBM GND efet w=24650 l=10150
M2500 GND ~OPE N0415 GND efet w=44225 l=10875
M2501 GND N0353 N0351 GND efet w=22475 l=10875
M2502 N0351 ~(X21&~CLK2) GND GND efet w=20300 l=11600
M2503 GND DCL N0353 GND efet w=14500 l=10150
M2504 WRITE_ACC(1) KBP GND GND efet w=14500 l=10150
M2505 N0415 ~(X21&~CLK2) GND GND efet w=44225 l=10875
M2506 VDD VDD N0383 GND efet w=5800 l=47850
M2507 N0375 N0380 GND GND efet w=21750 l=13775
M2508 VDD VDD ~(X31&~CLK2) GND efet w=5800 l=15950
M2509 N0353 VDD VDD GND efet w=6525 l=64525
M2510 GND TCS WRITE_ACC(1) GND efet w=13050 l=11600
M2511 WRITE_ACC(1) DAA GND GND efet w=13050 l=11600
M2512 S00699 VDD VDD GND efet w=5800 l=11600
M2513 VDD VDD ~(X21&~CLK2) GND efet w=6525 l=18850
M2514 ~(X31&~CLK2) N0375 GND GND efet w=65250 l=11600
M2515 N0375 VDD VDD GND efet w=5800 l=36250
M2516 N0369 VDD VDD GND efet w=5800 l=56550
M2517 N0337 VDD VDD GND efet w=5800 l=29000
M2518 VDD VDD N0328 GND efet w=6525 l=64525
M2519 N0720 N0282 GND GND efet w=26825 l=10875
M2520 N0282 CLK2 M22 GND efet w=15950 l=11600
M2521 N0721 CLK1 N0720 GND efet w=14500 l=11600
M2522 VDD VDD N0720 GND efet w=7250 l=30450
M2523 N0337 N0360 GND GND efet w=34800 l=12325
M2524 GND CLK2 N0337 GND efet w=28275 l=12325
M2525 ~(X21&~CLK2) N0337 GND GND efet w=53650 l=11600
M2526 GND N0329 N0328 GND efet w=13775 l=12325
M2527 N0328 POC GND GND efet w=11600 l=11600
M2528 N0330 X22 N0331 GND efet w=29000 l=13050
M2529 GND CLK2 N0330 GND efet w=29725 l=13775
M2530 N0369 X12 GND GND efet w=15225 l=12325
M2531 N0360 CLK2 N0369 GND efet w=9425 l=12325
M2532 N0335 CLK1 GND GND efet w=31175 l=12325
M2533 N0336 N0337 N0335 GND efet w=31175 l=10875
M2534 N0332 N0328 N0336 GND efet w=29725 l=12325
M2535 N0331 N0329 N0332 GND efet w=30450 l=10875
M2536 GND CLK2 N0423 GND efet w=21750 l=13050
M2537 N0332 POC N0331 GND efet w=29000 l=11600
M2538 N0351 VDD VDD GND efet w=7250 l=43500
M2539 GND INC/ISZ N0442 GND efet w=15950 l=10150
M2540 N0442 VDD VDD GND efet w=6525 l=58725
M2541 GND TCS WRITE_CARRY(2) GND efet w=11600 l=11600
M2542 GND TCS ADD_GROUP(4) GND efet w=12325 l=12325
M2543 READ_ACC(3) DAA GND GND efet w=13050 l=11600
M2544 GND N0446 N0448 GND efet w=76125 l=10875
M2545 N0342 N0332 VDD GND efet w=21025 l=11600
M2546 VDD VDD N0423 GND efet w=6525 l=31175
M2547 GND M22 N0288 GND efet w=22475 l=13775
M2548 VDD N0744 M22 GND efet w=40600 l=11600
M2549 M22 N0723 GND GND efet w=34800 l=11600
M2551 N0744 N0723 GND GND efet w=27550 l=13050
M2552 VDD VDD S00740 GND efet w=5800 l=11600
M2553 VDD S00740 N0744 GND efet w=4350 l=31175
M2554 VDD VDD N0430 GND efet w=5800 l=49300
M2555 N0340 VDD VDD GND efet w=7250 l=72500
M2556 N0430 N0423 N0431 GND efet w=10150 l=10875
M2557 N0722 N0283 GND GND efet w=26825 l=10875
M2558 N0283 CLK2 M12 GND efet w=13775 l=15225
M2559 N0723 CLK1 N0722 GND efet w=14500 l=11600
M2560 M12 CLK2 N0433 GND efet w=8700 l=12325
M2561 N0342 N0340 GND GND efet w=20300 l=13050
M2562 GND N0332 N0340 GND efet w=11600 l=11600
M2563 VDD S00731 N0332 GND efet w=6525 l=52925
M2564 S00731 VDD VDD GND efet w=6525 l=12325
M2566 VDD VDD N0805 GND efet w=11600 l=54375
M2567 N0853 VDD VDD GND efet w=7975 l=67425
M2568 X12 CLK2 N0425 GND efet w=7975 l=13050
M2569 N0421 VDD VDD GND efet w=5800 l=56550
M2570 N0421 N0423 N0422 GND efet w=10875 l=10875
M2571 GND N0422 N0805 GND efet w=31175 l=10150
M2572 N0853 X12 GND GND efet w=13050 l=11600
M2573 GND N0433 N0430 GND efet w=15225 l=12325
M2574 GND N0425 N0421 GND efet w=15225 l=10875
M2575 N0801 VDD VDD GND efet w=6525 l=51475
M2576 VDD VDD N0722 GND efet w=7975 l=38425
M2577 GND N0431 N0801 GND efet w=23925 l=13775
M2578 N0288 M12 GND GND efet w=21750 l=13050
M2579 VDD N0745 M12 GND efet w=39150 l=21750
M2580 GND N0803 N0403 GND efet w=24650 l=10150
M2581 M12 N0725 GND GND efet w=38425 l=12325
M2583 GND POC N0717 GND efet w=70325 l=12325
M2584 N0717 S00757 VDD GND efet w=10150 l=15950
M2586 N0403 N0802 GND GND efet w=21750 l=11600
M2587 GND ~(X21&~CLK2) N0448 GND efet w=73950 l=11600
M2588 GND XCH WRITE_ACC(1) GND efet w=13050 l=11600
M2589 WRITE_ACC(1) POC GND GND efet w=13050 l=11600
M2590 INC_GROUP(5) INC/ISZ GND GND efet w=11600 l=12325
M2591 WRITE_CARRY(2) POC GND GND efet w=15950 l=13050
M2592 GND CMA WRITE_ACC(1) GND efet w=13050 l=11600
M2593 WRITE_ACC(1) TCC GND GND efet w=13775 l=10875
M2594 GND DAC WRITE_ACC(1) GND efet w=11600 l=10150
M2595 WRITE_ACC(1) IAC GND GND efet w=11600 l=10150
M2596 GND N1005 ~OPA.1 GND efet w=34075 l=15225
M2597 WRITE_ACC(1) CLB GND GND efet w=12325 l=10875
M2598 VDD N1004 ~OPA.1 GND efet w=30450 l=26100
M2599 OPA.1 N1005 VDD GND efet w=26825 l=16675
M2600 GND LD WRITE_ACC(1) GND efet w=14500 l=11600
M2601 WRITE_ACC(1) SUB GND GND efet w=15225 l=10875
M2602 GND ADD WRITE_ACC(1) GND efet w=13775 l=10875
M2603 WRITE_ACC(1) LDM/BBL GND GND efet w=13775 l=10875
M2604 WRITE_CARRY(2) SUB GND GND efet w=16675 l=13775
M2605 WRITE_CARRY(2) TCC GND GND efet w=13050 l=11600
M2606 GND STC WRITE_CARRY(2) GND efet w=13050 l=11600
M2607 WRITE_CARRY(2) CMC GND GND efet w=13050 l=11600
M2608 GND DAC WRITE_CARRY(2) GND efet w=13775 l=11600
M2609 WRITE_CARRY(2) IAC GND GND efet w=15225 l=10875
M2610 GND CLC WRITE_CARRY(2) GND efet w=13050 l=11600
M2611 WRITE_CARRY(2) CLB GND GND efet w=13775 l=12325
M2612 GND SBM WRITE_CARRY(2) GND efet w=13050 l=10150
M2613 WRITE_CARRY(2) ADM GND GND efet w=13775 l=10150
M2614 GND RAR READ_ACC(3) GND efet w=13050 l=11600
M2615 READ_ACC(3) RAL GND GND efet w=13050 l=11600
M2616 N0448 N0445 ACB-IB GND efet w=74675 l=10875
M2617 ACB-IB ~(X31&~CLK2) N0448 GND efet w=76125 l=10875
M2618 GND N0442 ADD-IB GND efet w=39150 l=12325
M2619 GND XCH N0445 GND efet w=21750 l=11600
M2620 GND N0446 CY-IB GND efet w=14500 l=11600
M2621 GND IOW N0446 GND efet w=21750 l=11600
M2622 ADD_GROUP(4) TCC GND GND efet w=13050 l=13050
M2623 READ_ACC(3) IAC GND GND efet w=12325 l=14500
M2624 GND DAC READ_ACC(3) GND efet w=12325 l=10875
M2625 GND SBM READ_ACC(3) GND efet w=11600 l=10150
M2627 GND STC INC_GROUP(5) GND efet w=11600 l=11600
M2628 N0502 RAL GND GND efet w=15225 l=10875
M2629 CY-IB ~(X31&~CLK2) GND GND efet w=15950 l=12325
M2630 SUB_GROUP(6) CMC GND GND efet w=23925 l=15225
M2631 SUB_GROUP(6) S00709 VDD GND efet w=5800 l=40600
M2632 INC_GROUP(5) IAC GND GND efet w=14500 l=13050
M2633 INC_GROUP(5) VDD VDD GND efet w=7250 l=66700
M2634 READ_ACC(3) VDD VDD GND efet w=7250 l=69600
M2635 GND RAR N0490 GND efet w=15225 l=15225
M2636 GND ~(X31&~CLK2) ADSL GND efet w=17400 l=10875
M2637 GND ~(X31&~CLK2) ADD-IB GND efet w=38425 l=10875
M2639 ADD-IB S00729 VDD GND efet w=8700 l=24650
M2641 N0445 VDD VDD GND efet w=8700 l=41325
M2642 GND N0502 ADSL GND efet w=13050 l=13050
M2643 CY-IB VDD VDD GND efet w=7975 l=70325
M2644 N0446 VDD VDD GND efet w=8700 l=43500
M2645 GND ~(X31&~CLK2) ADSR GND efet w=14500 l=11600
M2646 ADSR N0490 GND GND efet w=15950 l=14500
M2647 GND CMA N0515 GND efet w=11600 l=11600
M2648 VDD VDD S00709 GND efet w=6525 l=13775
M2649 ACB-IB S00724 VDD GND efet w=10875 l=29725
M2650 VDD VDD ADSL GND efet w=8700 l=65250
M2651 N0502 VDD VDD GND efet w=5800 l=60900
M2652 VDD VDD N0490 GND efet w=7975 l=84825
M2653 ADSR VDD VDD GND efet w=7250 l=65250
M2654 ACC-ADAC N0515 GND GND efet w=13775 l=11600
M2655 GND N0342 ACC-ADAC GND efet w=13050 l=13050
M2656 WRITE_CARRY(2) VDD VDD GND efet w=6525 l=63800
M2657 N0515 VDD VDD GND efet w=7250 l=84100
M2658 GND N0853 N0854 GND efet w=19575 l=13775
M2659 READ_ACC(3) ADM GND GND efet w=13050 l=13050
M2660 ADD_GROUP(4) ADM GND GND efet w=12325 l=16675
M2661 GND SBM SUB_GROUP(6) GND efet w=21750 l=13050
M2662 ADD_GROUP(4) VDD VDD GND efet w=6525 l=60175
M2663 GND ADD WRITE_CARRY(2) GND efet w=13050 l=11600
M2664 READ_ACC(3) SUB GND GND efet w=13050 l=13050
M2665 GND IOR WRITE_ACC(1) GND efet w=13050 l=11600
M2666 GND ADD READ_ACC(3) GND efet w=13775 l=12325
M2667 GND ADD ADD_GROUP(4) GND efet w=13050 l=11600
M2668 SUB_GROUP(6) SUB GND GND efet w=23200 l=11600
M2669 VDD VDD N1001 GND efet w=13050 l=37700
M2670 OPA.2 N1003 VDD GND efet w=32625 l=25375
M2671 N1001 N1000 GND GND efet w=27550 l=14500
M2672 VDD VDD N1005 GND efet w=13050 l=33350
M2673 D1 OPA-IB OPA.1 GND efet w=58725 l=18125
M2674 GND CLK2 N0702 GND efet w=54375 l=12325
M2676 S00676 VDD VDD GND efet w=8700 l=15950
M2677 VDD VDD N0671 GND efet w=13050 l=33350
M2678 D0 OPA-IB OPA.0 GND efet w=65250 l=13050
M2679 GND N1007 ~OPA.0 GND efet w=37700 l=14500
M2680 OPA.0 N1006 GND GND efet w=70325 l=12325
M2681 N0702 S00676 VDD GND efet w=13050 l=15950
M2682 N0671 N0702 N0688 GND efet w=27550 l=13775
M2683 N0671 D3 GND GND efet w=53650 l=13050
M2684 VDD N1006 ~OPA.0 GND efet w=52925 l=25375
M2685 OPA.0 N1007 VDD GND efet w=29000 l=15225
M2686 VDD VDD N1003 GND efet w=12325 l=35525
M2687 N1005 N1004 GND GND efet w=26825 l=14500
M2688 GND N1012 N1000 GND efet w=56550 l=13050
M2689 GND N1014 N1004 GND efet w=55825 l=12325
M2690 GND JUN2+JMS2 N0658 GND efet w=15225 l=12325
M2691 N1003 N1002 GND GND efet w=26100 l=15225
M2692 VDD VDD N1007 GND efet w=9425 l=35525
M2693 N1007 N1006 GND GND efet w=34800 l=12325
M2694 GND N1013 N1002 GND efet w=57275 l=12325
M2695 GND N1015 N1006 GND efet w=64525 l=12325
M2696 VDD VDD S00689 GND efet w=8700 l=11600
M2697 S00687 VDD VDD GND efet w=8700 l=17400
M2699 N0687 S00687 VDD GND efet w=10150 l=14500
M2700 VDD S00689 N0689 GND efet w=10150 l=11600
M2702 VDD N0659 D0 GND efet w=47125 l=18125
M2703 N0687 N0700 GND GND efet w=253750 l=11600
M2704 GND N0700 N0689 GND efet w=228375 l=10875
M2705 N0687 N0688 GND GND efet w=98600 l=11600
M2706 GND N0687 N0689 GND efet w=74675 l=5800
M2707 D0 SC&M22&CLK2 N1015 GND efet w=10150 l=13050
M2708 VDD N0659 D2 GND efet w=47125 l=16675
M2709 N1000 VDD VDD GND efet w=19575 l=42050
M2710 N0658 LDM/BBL GND GND efet w=14500 l=10875
M2711 WRITE_ACC(1) VDD VDD GND efet w=6525 l=71775
M2712 N1004 VDD VDD GND efet w=11600 l=30450
M2713 N1002 VDD VDD GND efet w=19575 l=42050
M2714 N1006 VDD VDD GND efet w=20300 l=40600
M2715 D2 SC&M22&CLK2 N1013 GND efet w=10875 l=13775
M2716 GND N0689 D3_PAD GND efet w=1246275 l=6525
M2717 GND N0658 OPA-IB GND efet w=42050 l=15950
M2718 VDD VDD N0658 GND efet w=7250 l=69600
M2719 OPA-IB ~(X21&~CLK2) GND GND efet w=41325 l=10875
M2720 D1 SC&M22&CLK2 N1014 GND efet w=10875 l=13775
M2721 D3_PAD N0687 VDD GND efet w=657575 l=10875
M2723 D3 SC&M22&CLK2 N1012 GND efet w=10150 l=11600
M2724 VDD S00716 OPA-IB GND efet w=8700 l=20300
M2725 D1 N0659 VDD GND efet w=46400 l=13050
M2726 D3 N0659 VDD GND efet w=39875 l=12325
M2727 VDD VDD S00716 GND efet w=7250 l=11600
M2728 N0675 VDD VDD GND efet w=7975 l=36250
M2729 N0659 VDD VDD GND efet w=11600 l=21025
M2730 N0659 N0675 GND GND efet w=53650 l=10150
M2731 VDD VDD N0678 GND efet w=11600 l=37700
M2732 GND INC_GROUP(5) N0546 GND efet w=11600 l=12325
M2733 N0701 VDD VDD GND efet w=7250 l=20300
M2734 GND L N0686 GND efet w=57275 l=15225
M2735 GND L N0701 GND efet w=42775 l=10875
M2736 VDD VDD N0546 GND efet w=13050 l=87000
M2737 N0546 N0342 GND GND efet w=12325 l=14500
M2738 GND SUB_GROUP(6) CY-ADAC GND efet w=14500 l=11600
M2739 GND ADD_GROUP(4) CY-ADA GND efet w=11600 l=10875
M2740 VDD VDD N0677 GND efet w=8700 l=34075
M2741 N0685 CLK1 N0701 GND efet w=21025 l=18850
M2742 CY_1 ADSR N0513 GND efet w=14500 l=11600
M2743 S00729 VDD VDD GND efet w=5800 l=11600
M2744 S00724 VDD VDD GND efet w=6525 l=15225
M2745 CY N0415 N0860 GND efet w=15950 l=10150
M2746 N0860 N0403 VDD GND efet w=13775 l=13050
M2748 CY M12 N0470 GND efet w=7975 l=12325
M2749 N0550 CY-ADA N0470 GND efet w=14500 l=11600
M2750 N0470 VDD VDD GND efet w=10150 l=34800
M2751 N0470 N0855 GND GND efet w=41325 l=11600
M2752 N0513 ADSL CY GND efet w=14500 l=11600
M2753 D0 CY-IB CY_1 GND efet w=57275 l=10150
M2754 GND N0342 CY-ADAC GND efet w=13775 l=13775
M2756 N0861 ADC-CY CY GND efet w=10150 l=13050
M2757 GND CY N0855 GND efet w=59450 l=11600
M2758 N0855 VDD VDD GND efet w=10150 l=33350
M2759 N0846 ADSR CY GND efet w=7250 l=11600
M2760 CY-ADAC S00732 VDD GND efet w=6525 l=48575
M2761 GND N0342 CY-ADA GND efet w=13050 l=11600
M2762 GND READ_ACC(3) ACC-ADA GND efet w=14500 l=11600
M2763 GND N0342 ACC-ADA GND efet w=15225 l=14500
M2764 GND WRITE_CARRY(2) ADC-CY GND efet w=13775 l=10875
M2765 GND WRITE_ACC(1) ADD-ACC GND efet w=15225 l=11600
M2766 N0678 CLK1 GND GND efet w=22475 l=12325
M2767 N0686 CLK1 N0675 GND efet w=46400 l=11600
M2768 GND N0678 N0677 GND efet w=29000 l=15950
M2769 GND N0699 N0678 GND efet w=24650 l=14500
M2770 N0701 N0702 N0699 GND efet w=10150 l=11600
M2771 N0676 N0677 VDD GND efet w=41325 l=14500
M2772 N0678 N0685 GND GND efet w=23200 l=11600
M2773 GND N0678 N0676 GND efet w=45675 l=12325
M2774 GND N0477 ADC-CY GND efet w=13050 l=13050
M2775 GND N0477 ADD-ACC GND efet w=14500 l=13050
M2776 ADD-ACC VDD VDD GND efet w=10150 l=65250
M2777 VDD S00734 CY-ADA GND efet w=5800 l=58000
M2778 ADC-CY VDD VDD GND efet w=8700 l=79750
M2779 S00734 VDD VDD GND efet w=7250 l=11600
M2780 S00732 VDD VDD GND efet w=7975 l=10150
M2781 L CLK1 N0707 GND efet w=10875 l=13050
M2782 N0675 CLK2 N0684 GND efet w=44950 l=15950
M2783 N0684 N0685 GND GND efet w=56550 l=8700
M2784 N0705 N0707 GND GND efet w=59450 l=9425
M2785 N0705 L N0706 GND efet w=126150 l=13050
M2786 GND POC N0705 GND efet w=60175 l=11600
M2787 N0706 N0702 GND GND efet w=96425 l=10875
M2788 N0705 VDD VDD GND efet w=15225 l=27550
M2789 GND N0705 N0704 GND efet w=37700 l=15950
M2790 GND M12 N0550 GND efet w=10150 l=10150
M2791 N0550 N0546 VDD GND efet w=9425 l=15225
M2792 GND N0452 CY_1 GND efet w=53650 l=10150
M2793 CY_1 VDD VDD GND efet w=6525 l=29000
M2794 N0855 N0854 N0452 GND efet w=8700 l=10150
M2795 N0550 CY-ADAC N0855 GND efet w=15950 l=13050
M2796 GND SUB_GROUP(6) N0937 GND efet w=13050 l=11600
M2797 N0937 M12 GND GND efet w=18125 l=9425
M2798 N0704 VDD VDD GND efet w=9425 l=38425
M2799 N0700 N0704 VDD GND efet w=65975 l=12325
M2800 GND M12 SUB_GROUP(6) GND efet w=13775 l=11600
M2801 N0886 N0550 N0894 GND efet w=59450 l=11600
M2802 N0548 N0550 N0549 GND efet w=61625 l=10875
M2803 GND N0878 N0846 GND efet w=60900 l=11600
M2804 VDD VDD N0350 GND efet w=7250 l=50750
M2805 GND N0849 N0346 GND efet w=58725 l=12325
M2806 N0856 N0854 N0849 GND efet w=7975 l=12325
M2807 N0346 VDD VDD GND efet w=6525 l=32625
M2808 N0870 ACC-ADAC N0856 GND efet w=14500 l=13050
M2809 N0846 N0874 VDD GND efet w=13050 l=10150
M2810 N0894 N0870 GND GND efet w=44225 l=10875
M2811 GND CY_1 N0803 GND efet w=14500 l=17400
M2812 N0745 N0725 GND GND efet w=29000 l=13050
M2813 VDD VDD S00761 GND efet w=6525 l=11600
M2814 S00757 VDD VDD GND efet w=8700 l=13050
M2815 GND ~COM N0717 GND efet w=77575 l=10875
M2816 VDD S00761 N0745 GND efet w=5800 l=27550
M2817 N0725 CLK1 N0724 GND efet w=15950 l=10150
M2818 N0724 N0284 GND GND efet w=27550 l=13050
M2819 N0284 CLK2 A32 GND efet w=14500 l=11600
M2820 VDD VDD N0724 GND efet w=8700 l=40600
M2821 N0288 A32 GND GND efet w=23200 l=12325
M2822 GND DAA N0802 GND efet w=13050 l=11600
M2823 N0818 N0803 GND GND efet w=28275 l=11600
M2824 N0378 DAA N0818 GND efet w=29000 l=11600
M2825 GND O-IB N0378 GND efet w=15225 l=10875
M2826 N0350 KBP GND GND efet w=17400 l=11600
M2827 N0856 VDD VDD GND efet w=10150 l=37700
M2828 N0803 N0356 N0819 GND efet w=28275 l=10150
M2829 VDD N0746 A32 GND efet w=38425 l=12325
M2830 A32 N0727 GND GND efet w=39150 l=13050
M2832 N0746 N0727 GND GND efet w=34800 l=13050
M2833 VDD VDD S00778 GND efet w=5800 l=13050
M2834 VDD S00778 N0746 GND efet w=7250 l=26100
M2835 VDD VDD N0766 GND efet w=8700 l=43500
M2836 VDD VDD N0751 GND efet w=7975 l=45675
M2837 DCL.0 VDD VDD GND efet w=7250 l=44950
M2838 GND N0348 N0819 GND efet w=34800 l=10875
M2839 N0819 N0347 GND GND efet w=37700 l=11600
M2840 N0803 VDD VDD GND efet w=5800 l=50750
M2841 N0403 VDD VDD GND efet w=6525 l=33350
M2842 N0802 VDD VDD GND efet w=6525 l=70325
M2843 N0354 VDD VDD GND efet w=7250 l=46400
M2844 N0363 VDD VDD GND efet w=9425 l=50025
M2845 N0370 VDD VDD GND efet w=7975 l=42775
M2846 VDD VDD N0345 GND efet w=7975 l=51475
M2847 N0378 VDD VDD GND efet w=7250 l=47850
M2848 N0377 N0378 N0376 GND efet w=34075 l=12325
M2849 GND N0346 ACC_0 GND efet w=21750 l=11600
M2850 CY_1 ADSL ACC.0 GND efet w=7250 l=12325
M2851 GND ACC.0 N0856 GND efet w=61625 l=11600
M2852 GND M12 N0870 GND efet w=13050 l=12325
M2853 N0471 VDD VDD GND efet w=9425 l=36975
M2854 N0346 ACB-IB D0 GND efet w=43500 l=10875
M2855 ACC_0 VDD VDD GND efet w=8700 l=44950
M2856 GND N0846 ADD_0 GND efet w=42775 l=10875
M2857 ACC.0 M12 N0471 GND efet w=7250 l=11600
M2858 N0846 ADD-ACC ACC.0 GND efet w=10150 l=11600
M2859 GND N0878 N0874 GND efet w=12325 l=13775
M2860 N0878 N0887 N0886 GND efet w=60900 l=12325
M2861 N0548 N0870 GND GND efet w=62350 l=11600
M2862 N0549 N0887 GND GND efet w=50025 l=10875
M2863 GND N0856 N0471 GND efet w=36250 l=11600
M2864 N0874 VDD VDD GND efet w=5800 l=59450
M2865 N0549 N0870 N0911 GND efet w=68875 l=17400
M2866 N0911 N0887 N0548 GND efet w=55825 l=12325
M2867 ~TMP.0 N0940 GND GND efet w=22475 l=12325
M2868 GND N0705 N0700 GND efet w=95700 l=8700
M2869 ~TMP.0 N0937 N0887 GND efet w=13775 l=10875
M2870 VDD N0939 ~TMP.0 GND efet w=14500 l=11600
M2871 VDD VDD N0911 GND efet w=5800 l=66700
M2872 N0847 ADSR ACC.0 GND efet w=10150 l=11600
M2873 N0878 VDD VDD GND efet w=7250 l=53650
M2874 N0898 N0553 N0878 GND efet w=36250 l=13050
M2875 GND N0870 N0898 GND efet w=35525 l=13775
M2876 N0898 N0550 GND GND efet w=43500 l=13050
M2877 GND N0887 N0898 GND efet w=35525 l=12325
M2878 N0915 N0911 GND GND efet w=11600 l=11600
M2879 VDD VDD N0915 GND efet w=7250 l=63075
M2880 D0 ADD-IB N0846 GND efet w=40600 l=11600
M2881 N0870 ACC-ADA N0471 GND efet w=14500 l=13050
M2882 N0940 VDD VDD GND efet w=6525 l=45675
M2883 GND N0939 N0940 GND efet w=15225 l=12325
M2884 TMP.0 SUB_GROUP(6) N0887 GND efet w=15225 l=12325
M2885 TMP.0 N0940 VDD GND efet w=13050 l=11600
M2886 GND N0939 TMP.0 GND efet w=23200 l=10875
M2887 VDD M12 N0604 GND efet w=7250 l=11600
M2888 N0553 N0915 GND GND efet w=20300 l=10150
M2889 D0 N0964 N0604 GND efet w=12325 l=12325
M2890 GND N0604 N0939 GND efet w=42050 l=13775
M2892 N0939 S00762 VDD GND efet w=5800 l=47850
M2893 VDD N0911 N0553 GND efet w=14500 l=11600
M2894 GND N0884 N0847 GND efet w=63075 l=13775
M2895 VDD S00764 ACC-ADAC GND efet w=5800 l=45675
M2897 ADD_0 VDD VDD GND efet w=8700 l=46400
M2898 VDD VDD N0377 GND efet w=8700 l=43500
M2899 GND DCL.0 N0751 GND efet w=35525 l=10150
M2900 N0766 N0351 GND GND efet w=22475 l=13050
M2901 GND DCL.0 N0716 GND efet w=47850 l=10150
M2902 N0751 N0766 N0767 GND efet w=12325 l=12325
M2903 DCL.0 POC GND GND efet w=23200 l=11600
M2904 GND N0350 N0376 GND efet w=37700 l=13050
M2905 GND N0767 DCL.0 GND efet w=50750 l=10150
M2906 N0345 N0350 GND GND efet w=17400 l=13050
M2907 N0354 N0350 GND GND efet w=14500 l=11600
M2908 GND N0350 N0363 GND efet w=17400 l=13050
M2909 N0370 N0350 GND GND efet w=18125 l=13775
M2910 VDD VDD N0371 GND efet w=5800 l=59450
M2911 GND N0847 ADD_0 GND efet w=39875 l=10875
M2912 N0847 ADD-IB D1 GND efet w=39875 l=11600
M2913 VDD VDD S00764 GND efet w=5800 l=11600
M2914 N0847 N0875 VDD GND efet w=15950 l=13050
M2915 VDD VDD S00767 GND efet w=9425 l=10875
M2916 D1 ACB-IB N0347 GND efet w=39875 l=11600
M2917 N0871 ACC-ADAC N0472 GND efet w=14500 l=13050
M2918 N0888 N0553 N0895 GND efet w=57275 l=10875
M2919 N0895 N0871 GND GND efet w=58000 l=11600
M2920 N0875 N0889 N0888 GND efet w=60175 l=11600
M2921 GND N0347 ACC_0 GND efet w=23200 l=10150
M2922 N0472 VDD VDD GND efet w=10875 l=35525
M2923 N0472 M12 ACC.1 GND efet w=8700 l=11600
M2924 N0472 N0857 GND GND efet w=36975 l=11600
M2925 N0846 ADSL ACC.1 GND efet w=8700 l=12325
M2926 GND N0875 N0884 GND efet w=12325 l=10875
M2927 N0551 N0553 N0552 GND efet w=60900 l=10150
M2928 N0551 N0871 GND GND efet w=65975 l=12325
M2929 N0552 N0889 GND GND efet w=48575 l=10875
M2930 N0370 N0371 GND GND efet w=17400 l=11600
M2931 N0371 N0346 GND GND efet w=14500 l=10150
M2932 VDD VDD N0364 GND efet w=6525 l=68875
M2933 N0726 N0285 GND GND efet w=27550 l=11600
M2934 N0285 CLK2 A22 GND efet w=13775 l=12325
M2935 N0727 CLK1 N0726 GND efet w=14500 l=11600
M2936 VDD VDD N0726 GND efet w=7975 l=37700
M2937 GND DCL.1 N0716 GND efet w=49300 l=11600
M2938 N0371 N0351 N0767 GND efet w=12325 l=10150
M2939 N0912 N0889 N0551 GND efet w=57275 l=13775
M2940 N0552 N0871 N0912 GND efet w=67425 l=15225
M2942 S00762 VDD VDD GND efet w=8700 l=11600
M2943 GND N0342 N0964 GND efet w=23925 l=13775
M2944 N0964 VDD VDD GND efet w=10875 l=35525
M2945 GND N0871 N0899 GND efet w=34800 l=14500
M2946 GND ACC.1 N0857 GND efet w=59450 l=11600
M2947 N0847 ADD-ACC ACC.1 GND efet w=8700 l=11600
M2948 N0884 VDD VDD GND efet w=10150 l=47125
M2949 N0857 VDD VDD GND efet w=10150 l=33350
M2950 N0848 ADSR ACC.1 GND efet w=7975 l=13775
M2951 N0347 VDD VDD GND efet w=7250 l=33350
M2952 GND N0850 N0347 GND efet w=58000 l=11600
M2953 N0857 N0854 N0850 GND efet w=8700 l=11600
M2954 VDD M12 N0871 GND efet w=13050 l=11600
M2955 N0875 VDD VDD GND efet w=8700 l=65250
M2956 N0899 N0556 N0875 GND efet w=35525 l=12325
M2957 N0899 N0553 GND GND efet w=43500 l=13050
M2958 GND N0889 N0899 GND efet w=36250 l=10150
M2959 N0871 ACC-ADA N0857 GND efet w=15950 l=12325
M2960 N0345 N0346 GND GND efet w=18125 l=12325
M2961 GND N0346 N0354 GND efet w=14500 l=10150
M2962 GND N0346 N0363 GND efet w=19575 l=10875
M2963 N0288 A22 GND GND efet w=23200 l=13050
M2964 GND N0765 DCL.1 GND efet w=39150 l=11600
M2965 GND N0346 N0376 GND efet w=36250 l=11600
M2966 GND N0879 N0848 GND efet w=60900 l=10150
M2967 VDD S00767 N0912 GND efet w=5800 l=51475
M2968 TMP.1 N0937 N0889 GND efet w=14500 l=11600
M2969 ~TMP.1 N0942 GND GND efet w=20300 l=11600
M2970 N0672 D2 GND GND efet w=57275 l=12325
M2971 D2_PAD POC GND GND efet w=29725 l=13775
M2972 VDD VDD N0672 GND efet w=10875 l=40600
M2973 S00765 VDD VDD GND efet w=7250 l=15950
M2974 S00766 VDD VDD GND efet w=7250 l=15225
M2976 VDD S00766 N0692 GND efet w=10150 l=12325
M2977 N0690 S00765 VDD GND efet w=12325 l=18125
M2978 VDD N0941 ~TMP.1 GND efet w=13775 l=12325
M2979 N0691 N0702 N0672 GND efet w=27550 l=12325
M2980 N0942 VDD VDD GND efet w=6525 l=47125
M2981 N0916 N0912 GND GND efet w=13050 l=10150
M2982 VDD VDD N0916 GND efet w=7250 l=63075
M2983 GND N0941 N0942 GND efet w=13050 l=11600
M2985 VDD M12 N0605 GND efet w=7975 l=10150
M2986 TMP.1 N0942 VDD GND efet w=14500 l=11600
M2987 ~TMP.1 SUB_GROUP(6) N0889 GND efet w=18125 l=12325
M2988 GND N0941 TMP.1 GND efet w=20300 l=11600
M2989 N0690 N0700 GND GND efet w=262450 l=13050
M2990 D1 N0964 N0605 GND efet w=12325 l=13775
M2991 N0556 N0916 GND GND efet w=20300 l=10150
M2992 N0692 N0700 GND GND efet w=228375 l=10150
M2993 GND N0605 N0941 GND efet w=41325 l=18125
M2994 VDD N0912 N0556 GND efet w=14500 l=10150
M2996 N0941 S00781 VDD GND efet w=5800 l=43500
M2997 GND N0851 N0348 GND efet w=56550 l=11600
M2998 N0858 N0854 N0851 GND efet w=7250 l=13050
M2999 N0348 VDD VDD GND efet w=8700 l=29000
M3000 VDD N0747 A22 GND efet w=41325 l=10875
M3001 A22 N0729 GND GND efet w=37700 l=11600
M3002 GND POC DCL.1 GND efet w=23200 l=11600
M3003 DCL.1 VDD VDD GND efet w=7250 l=49300
M3004 N0364 N0351 N0765 GND efet w=12325 l=15225
M3005 GND N0364 N0363 GND efet w=17400 l=10150
M3006 GND N0347 N0345 GND efet w=24650 l=12325
M3007 N0354 N0347 GND GND efet w=13775 l=12325
M3008 N0364 N0347 GND GND efet w=14500 l=10150
M3009 N0872 ACC-ADAC N0858 GND efet w=15225 l=12325
M3010 N0848 N0876 VDD GND efet w=13775 l=15225
M3011 N0858 VDD VDD GND efet w=10150 l=41325
M3012 GND N0347 N0370 GND efet w=18850 l=10150
M3013 GND N0347 N0376 GND efet w=36250 l=10150
M3014 GND DCL.1 N0750 GND efet w=23200 l=11600
M3015 N0750 VDD VDD GND efet w=7250 l=52200
M3017 N0747 N0729 GND GND efet w=32625 l=15225
M3018 VDD VDD S00800 GND efet w=6525 l=13775
M3019 VDD S00800 N0747 GND efet w=5800 l=24650
M3020 N0750 N0766 N0765 GND efet w=10150 l=11600
M3021 VDD VDD N0355 GND efet w=6525 l=73225
M3022 N0355 N0351 N0768 GND efet w=10150 l=10150
M3023 N0354 N0355 GND GND efet w=13050 l=11600
M3024 N0355 N0348 GND GND efet w=15225 l=10875
M3025 GND N0348 ACC_0 GND efet w=23200 l=11600
M3026 N0847 ADSL ACC.2 GND efet w=7250 l=14500
M3027 GND ACC.2 N0858 GND efet w=64525 l=11600
M3028 N0473 VDD VDD GND efet w=12325 l=36975
M3029 GND N0848 ADD_0 GND efet w=42775 l=10875
M3030 N0348 ACB-IB D2 GND efet w=39150 l=13775
M3031 N0848 ADD-ACC ACC.2 GND efet w=7975 l=11600
M3032 ACC.2 M12 N0473 GND efet w=7975 l=12325
M3033 GND N0858 N0473 GND efet w=36250 l=11600
M3034 N0890 N0556 N0896 GND efet w=59450 l=11600
M3035 N0896 N0872 GND GND efet w=60900 l=10150
M3036 N0879 N0891 N0890 GND efet w=65250 l=10875
M3037 N0554 N0872 GND GND efet w=64525 l=10875
M3038 GND N0879 N0876 GND efet w=10150 l=12325
M3039 GND M12 N0872 GND efet w=15225 l=10875
M3040 N0514 ADSR ACC.2 GND efet w=9425 l=12325
M3041 N0555 N0891 GND GND efet w=52925 l=10875
M3042 N0555 N0872 N0913 GND efet w=68150 l=14500
M3043 N0913 N0891 N0554 GND efet w=56550 l=11600
M3044 N0876 VDD VDD GND efet w=8700 l=65975
M3045 D2 ADD-IB N0848 GND efet w=42775 l=11600
M3046 N0872 ACC-ADA N0473 GND efet w=14500 l=11600
M3047 N0879 VDD VDD GND efet w=9425 l=57275
M3048 GND DCL.2 N0716 GND efet w=43500 l=10150
M3049 N0728 N0286 GND GND efet w=27550 l=11600
M3050 N0729 CLK1 N0728 GND efet w=13775 l=12325
M3051 N0286 CLK2 A12 GND efet w=15950 l=11600
M3052 GND N0768 DCL.2 GND efet w=42050 l=10150
M3053 GND N0348 N0345 GND efet w=18850 l=11600
M3054 GND N0348 N0363 GND efet w=20300 l=11600
M3055 GND N0348 N0370 GND efet w=19575 l=10875
M3056 GND N0348 N0376 GND efet w=36250 l=10150
M3057 N0900 N0559 N0879 GND efet w=34800 l=12325
M3058 GND N0872 N0900 GND efet w=36250 l=10150
M3059 N0900 N0556 GND GND efet w=43500 l=11600
M3060 GND N0891 N0900 GND efet w=40600 l=13050
M3062 N0554 N0556 N0555 GND efet w=60900 l=11600
M3063 GND N0691 N0690 GND efet w=97875 l=9425
M3064 D2 N0964 N0606 GND efet w=19575 l=17400
M3065 GND N0690 N0692 GND efet w=73950 l=11600
M3066 S00781 VDD VDD GND efet w=9425 l=12325
M3067 VDD VDD N0913 GND efet w=5800 l=58000
M3068 ~TMP.2 N0944 GND GND efet w=22475 l=11600
M3069 ~TMP.2 N0937 N0891 GND efet w=15950 l=10875
M3070 VDD N0943 ~TMP.2 GND efet w=14500 l=13050
M3071 GND N0692 D2_PAD GND efet w=1202775 l=7250
M3072 N0606 M12 VDD GND efet w=8700 l=11600
M3073 N0665 N0676 GND GND efet w=26100 l=13050
M3074 N0917 N0913 GND GND efet w=13050 l=10875
M3075 VDD VDD N0917 GND efet w=5800 l=63800
M3076 N0559 N0917 GND GND efet w=20300 l=11600
M3077 VDD N0913 N0559 GND efet w=15225 l=10875
M3078 VDD VDD S00804 GND efet w=5800 l=11600
M3079 N0944 VDD VDD GND efet w=7975 l=44225
M3080 GND N0943 N0944 GND efet w=13775 l=15225
M3081 TMP.2 N0944 VDD GND efet w=15950 l=13775
M3082 GND N0943 TMP.2 GND efet w=19575 l=13775
M3083 TMP.2 SUB_GROUP(6) N0891 GND efet w=15225 l=12325
M3084 D2_PAD N0690 VDD GND efet w=640175 l=13775
M3085 VDD VDD N0665 GND efet w=11600 l=52200
M3086 N0665 N0666 GND GND efet w=14500 l=13050
M3087 N0943 S00801 VDD GND efet w=8700 l=53650
M3088 VDD VDD N0349 GND efet w=6525 l=61625
M3089 VDD S00803 ACC-ADA GND efet w=6525 l=45675
M3090 VDD VDD N0728 GND efet w=7250 l=38425
M3091 N0288 A12 GND GND efet w=22475 l=11600
M3092 DCL.2 VDD VDD GND efet w=8700 l=43500
M3093 N0749 VDD VDD GND efet w=7250 l=43500
M3094 VDD N0748 A12 GND efet w=39150 l=13050
M3095 GND POC DCL.2 GND efet w=26100 l=10875
M3096 GND DCL.2 N0749 GND efet w=23200 l=11600
M3097 A12 N0731 GND GND efet w=38425 l=12325
M3099 N0748 N0731 GND GND efet w=27550 l=11600
M3100 VDD VDD S00814 GND efet w=5800 l=12325
M3101 N0768 N0766 N0749 GND efet w=9425 l=13775
M3102 GND N0349 N0345 GND efet w=19575 l=13050
M3103 N0354 N0356 GND GND efet w=15225 l=10875
M3104 N0349 N0356 GND GND efet w=11600 l=10150
M3105 GND N0514 ADD_0 GND efet w=41325 l=10875
M3106 GND N0356 N0363 GND efet w=17400 l=10150
M3107 GND N0356 N0370 GND efet w=19575 l=15225
M3108 GND N0356 N0376 GND efet w=33350 l=10150
M3109 VDD S00814 N0748 GND efet w=5800 l=26100
M3110 N0514 ADD-IB D3 GND efet w=40600 l=11600
M3111 VDD VDD S00803 GND efet w=5800 l=10150
M3112 N0514 N0877 VDD GND efet w=19575 l=12325
M3113 D3 ACB-IB N0356 GND efet w=40600 l=11600
M3114 N0873 ACC-ADAC N0474 GND efet w=15950 l=13775
M3115 GND N0377 N0358 GND efet w=64525 l=13775
M3116 GND N0345 N0358 GND efet w=72500 l=11600
M3117 N0358 N0354 GND GND efet w=66700 l=11600
M3118 GND N0363 N0358 GND efet w=74675 l=12325
M3119 N0358 N0370 GND GND efet w=60175 l=10875
M3120 N0358 VDD VDD GND efet w=6525 l=65975
M3122 N0714 N0749 GND GND efet w=45675 l=12325
M3123 N0731 CLK1 N0730 GND efet w=13775 l=10150
M3124 N0730 N0287 GND GND efet w=29000 l=12325
M3125 VDD VDD N0730 GND efet w=7975 l=39150
M3126 N0287 CLK2 N0288 GND efet w=13050 l=11600
M3127 GND ~COM N0714 GND efet w=45675 l=10875
M3128 VDD VDD S00818 GND efet w=7975 l=12325
M3129 VDD S00818 N0714 GND efet w=10150 l=24650
M3130 N0366 VDD VDD GND efet w=5800 l=66700
M3131 VDD VDD N0288 GND efet w=8700 l=34800
M3133 N0715 N0750 GND GND efet w=44950 l=11600
M3134 VDD N0714 CMRAM3 GND efet w=142100 l=11600
M3135 N0734 N0714 GND GND efet w=47850 l=18850
M3136 GND ~COM N0715 GND efet w=43500 l=10150
M3137 N0366 N0354 GND GND efet w=61625 l=10875
M3138 GND N0363 N0366 GND efet w=59450 l=11600
M3139 N0366 N0370 GND GND efet w=60900 l=10875
M3140 GND N0377 N0366 GND efet w=59450 l=11600
M3141 GND N0403 N0358 GND efet w=60900 l=10150
M3142 GND N0356 ACC_0 GND efet w=23200 l=11600
M3143 N0474 VDD VDD GND efet w=10875 l=35525
M3144 N0356 N0852 GND GND efet w=53650 l=13050
M3145 N0356 VDD VDD GND efet w=8700 l=34800
M3146 N0366 TCS GND GND efet w=60175 l=10875
M3147 VDD VDD S00825 GND efet w=7975 l=12325
M3148 VDD N0715 CMRAM2 GND efet w=141375 l=12325
M3149 VDD VDD N0734 GND efet w=8700 l=20300
M3150 VDD VDD N0735 GND efet w=9425 l=19575
M3151 GND N0715 N0735 GND efet w=40600 l=13050
M3152 VDD S00825 N0715 GND efet w=10150 l=24650
M3153 N0359 VDD VDD GND efet w=6525 l=61625
M3154 GND N0345 N0359 GND efet w=61625 l=10875
M3155 N0357 VDD VDD GND efet w=6525 l=68150
M3157 CMRAM2 N0735 GND GND efet w=263900 l=14500
M3158 CMRAM3 N0734 GND GND efet w=263900 l=11600
M3159 GND ~COM N0713 GND efet w=43500 l=13050
M3160 N0716 ~COM GND GND efet w=59450 l=11600
M3162 S00834 VDD VDD GND efet w=7975 l=12325
M3163 N0713 N0751 GND GND efet w=47125 l=10875
M3164 N0359 N0370 GND GND efet w=65975 l=12325
M3165 GND N0377 N0359 GND efet w=60175 l=12325
M3166 D2 N0415 N0366 GND efet w=49300 l=11600
M3167 D3 N0415 N0358 GND efet w=49300 l=14500
M3168 N0359 TCS GND GND efet w=59450 l=11600
M3169 VDD VDD S00833 GND efet w=7975 l=12325
M3170 VDD S00833 N0716 GND efet w=10875 l=23925
M3171 N0713 S00834 VDD GND efet w=9425 l=22475
M3172 GND N0345 N0357 GND efet w=62350 l=13775
M3173 GND N0363 N0357 GND efet w=63800 l=15950
M3174 GND N0377 N0357 GND efet w=60175 l=12325
M3175 D1 N0415 N0359 GND efet w=50750 l=11600
M3176 D0 N0415 N0357 GND efet w=55825 l=11600
M3177 N0474 M12 ACC.3 GND efet w=8700 l=11600
M3178 N0474 N0859 GND GND efet w=36250 l=11600
M3179 N0848 ADSL ACC.3 GND efet w=8700 l=11600
M3180 GND N0885 N0514 GND efet w=65975 l=10875
M3181 GND N0606 N0943 GND efet w=41325 l=13775
M3182 N0897 N0873 GND GND efet w=60175 l=10875
M3183 GND N0877 N0885 GND efet w=13775 l=10150
M3184 N0892 N0559 N0897 GND efet w=56550 l=11600
M3185 N0877 N0893 N0892 GND efet w=65250 l=10150
M3186 N0557 N0873 GND GND efet w=76125 l=19575
M3187 GND N0893 N0558 GND efet w=61625 l=28275
M3188 GND ACC.3 N0859 GND efet w=58725 l=13775
M3189 N0514 ADD-ACC ACC.3 GND efet w=9425 l=10875
M3190 N0859 VDD VDD GND efet w=9425 l=35525
M3191 N0514 ADSL N0513 GND efet w=15225 l=12325
M3192 N0859 N0854 N0852 GND efet w=7250 l=13050
M3193 N0513 ADSR ACC.3 GND efet w=13050 l=13775
M3194 N0914 N0893 N0557 GND efet w=55825 l=12325
M3195 GND N0873 N0901 GND efet w=35525 l=12325
M3196 N0885 VDD VDD GND efet w=9425 l=54375
M3197 VDD M12 N0873 GND efet w=13775 l=12325
M3198 N0901 N0861 N0877 GND efet w=37700 l=10150
M3199 N0877 VDD VDD GND efet w=7975 l=64525
M3200 N0873 ACC-ADA N0859 GND efet w=15950 l=10875
M3201 N0558 N0873 N0914 GND efet w=65975 l=16675
M3202 N0901 N0559 GND GND efet w=43500 l=10150
M3203 GND N0893 N0901 GND efet w=37700 l=11600
M3204 N0557 N0559 N0558 GND efet w=58000 l=10150
M3207 S00801 VDD VDD GND efet w=12325 l=13050
M3208 D2 N0666 GND GND efet w=49300 l=13775
M3209 VDD N0665 D2 GND efet w=39875 l=15225
M3210 VDD S00804 N0914 GND efet w=5075 l=52200
M3211 VDD VDD N0666 GND efet w=10150 l=39150
M3212 ~TMP.3 N0946 GND GND efet w=21025 l=13050
M3213 N0666 D2_PAD GND GND efet w=71050 l=12325
M3214 ~TMP.3 SUB_GROUP(6) N0893 GND efet w=14500 l=11600
M3215 N0666 N0676 GND GND efet w=44950 l=12325
M3216 VDD N0945 ~TMP.3 GND efet w=13775 l=12325
M3217 N0918 N0914 GND GND efet w=12325 l=12325
M3218 VDD VDD N0918 GND efet w=5800 l=63800
M3219 N0861 N0918 GND GND efet w=18850 l=11600
M3220 N0946 VDD VDD GND efet w=8700 l=43500
M3221 GND N0945 N0946 GND efet w=13050 l=11600
M3222 VDD M12 N0607 GND efet w=9425 l=8700
M3223 TMP.3 N0937 N0893 GND efet w=15225 l=12325
M3224 TMP.3 N0946 VDD GND efet w=13775 l=12325
M3225 VDD N0914 N0861 GND efet w=13050 l=11600
M3226 VDD VDD S00817 GND efet w=6525 l=9425
M3227 GND N0945 TMP.3 GND efet w=20300 l=11600
M3228 D3 N0964 N0607 GND efet w=14500 l=14500
M3230 GND N0607 N0945 GND efet w=38425 l=13775
M3231 D0_PAD GND GND GND efet w=116000 l=13050
M3233 GND N0403 N0357 GND efet w=60175 l=13775
M3234 VDD VDD S00819 GND efet w=7250 l=9425
M3235 N0945 S00817 VDD GND efet w=5800 l=40600
M3237 N0670 D0_PAD GND GND efet w=71775 l=12325
M3238 GND N0670 D0 GND efet w=49300 l=11600
M3239 GND N0670 N0669 GND efet w=13775 l=11600
M3240 D1_PAD GND GND GND efet w=114550 l=14500
M3241 N0854 S00828 VDD GND efet w=7250 l=52200
M3242 VDD VDD S00828 GND efet w=8700 l=13050
M3243 N0670 N0676 GND GND efet w=51475 l=13775
M3244 GND N0676 N0669 GND efet w=25375 l=11600
M3245 D0 N0669 VDD GND efet w=38425 l=13050
M3246 N0670 VDD VDD GND efet w=10150 l=36975
M3247 N0669 VDD VDD GND efet w=5800 l=50750
M3248 GND D0 N0674 GND efet w=57275 l=12325
M3249 N0674 VDD VDD GND efet w=13050 l=39150
M3250 N0674 N0702 N0697 GND efet w=27550 l=11600
M3251 GND N0697 N0696 GND efet w=99325 l=10875
M3252 D0_PAD N0696 VDD GND efet w=666275 l=10875
M3253 N0733 N0713 GND GND efet w=55100 l=14500
M3254 VDD N0713 CMRAM1 GND efet w=142100 l=11600
M3255 VDD N0716 CMRAM0 GND efet w=142100 l=11600
M3256 VDD VDD N0733 GND efet w=7250 l=23200
M3257 VDD VDD N0736 GND efet w=8700 l=21750
M3258 GND N0716 N0736 GND efet w=43500 l=11600
M3259 CMRAM1 N0733 GND GND efet w=261725 l=12325
M3260 CMRAM0 N0736 GND GND efet w=256650 l=11600
M3261 GND N0698 D0_PAD GND efet w=1218725 l=6525
M3262 N0696 N0700 GND GND efet w=247950 l=11600
M3263 VDD VDD S00835 GND efet w=9425 l=12325
M3264 VDD S00835 N0696 GND efet w=10875 l=13775
M3266 GND N0696 N0698 GND efet w=81925 l=12325
M3267 N0698 N0700 GND GND efet w=229100 l=11600
M3268 VDD S00839 N0698 GND efet w=10150 l=11600
M3270 VDD VDD S00839 GND efet w=10150 l=13050
M3271 N0668 D1_PAD GND GND efet w=66700 l=13050
M3272 N0937 S00819 VDD GND efet w=6525 l=33350
M3273 GND GND D2_PAD GND efet w=99325 l=15225
M3274 GND N0668 D1 GND efet w=49300 l=11600
M3275 N0667 N0668 GND GND efet w=16675 l=10875
M3276 GND N0676 N0667 GND efet w=26825 l=12325
M3277 N0668 N0676 GND GND efet w=44225 l=13775
M3278 VDD VDD N0667 GND efet w=6525 l=55825
M3279 D1 N0667 VDD GND efet w=39150 l=11600
M3280 N0668 VDD VDD GND efet w=8700 l=35525
M3281 GND D1 N0673 GND efet w=50750 l=10875
M3282 N0673 N0702 N0694 GND efet w=27550 l=12325
M3283 N0673 VDD VDD GND efet w=10875 l=36975
M3284 D3 N0664 GND GND efet w=49300 l=12325
M3285 VDD N0663 D3 GND efet w=39875 l=12325
M3286 GND POC D3_PAD GND efet w=29000 l=14500
M3287 VDD N0693 D1_PAD GND efet w=681500 l=11600
M3288 D0_PAD POC GND GND efet w=33350 l=11600
M3289 GND N0694 N0693 GND efet w=99325 l=10875
M3290 N0693 N0700 GND GND efet w=257375 l=19575
M3291 VDD VDD S00836 GND efet w=7250 l=11600
M3292 VDD S00836 N0693 GND efet w=9425 l=13775
M3293 GND N0695 D1_PAD GND efet w=1217275 l=6525
M3295 VDD VDD N0663 GND efet w=9425 l=49300
M3296 VDD VDD N0664 GND efet w=8700 l=36250
M3297 GND N0676 N0664 GND efet w=56550 l=14500
M3298 GND N0693 N0695 GND efet w=75400 l=13050
M3299 N0695 N0700 GND GND efet w=229825 l=10875
M3300 VDD S00840 N0695 GND efet w=10150 l=14500
M3302 VDD VDD S00840 GND efet w=7250 l=13775
M3303 GND N0664 N0663 GND efet w=23200 l=15950
M3304 N0663 N0676 GND GND efet w=23925 l=11600
M3305 GND D3_PAD N0664 GND efet w=86275 l=15225
M3306 D3_PAD GND GND GND efet w=124700 l=13050
M3307 D1_PAD POC GND GND efet w=30450 l=10875
