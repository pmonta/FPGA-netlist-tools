* SPICE3 file created from 6800.ext - technology: 6800-nmos

.option scale=0.001u

M1000 diff_82000_3097000# diff_82000_3097000# diff_82000_3097000# GND efet w=500 l=8000
+ ad=-1.55338e+09 pd=3.46428e+08 as=0 ps=0 
M1001 diff_616000_6169000# diff_82000_3097000# diff_82000_3097000# GND efet w=84000 l=14000
+ ad=1.43813e+09 pd=3.178e+06 as=0 ps=0 
M1002 diff_1119000_5759000# diff_1277000_5967000# diff_82000_3097000# GND efet w=164500 l=10500
+ ad=8.64033e+08 pd=644000 as=0 ps=0 
M1003 diff_82000_3097000# diff_1277000_5967000# diff_1129000_5768000# GND efet w=327500 l=10500
+ ad=0 pd=0 as=-8.60706e+08 ps=4.128e+06 
M1004 diff_82000_3097000# diff_1277000_5967000# diff_1129000_5768000# GND efet w=328500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1005 diff_1119000_5759000# diff_1277000_5967000# diff_82000_3097000# GND efet w=164500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1006 diff_1277000_5967000# diff_1585000_6056000# diff_82000_3097000# GND efet w=306500 l=10500
+ ad=-7.82967e+08 pd=434000 as=0 ps=0 
M1007 diff_82000_3097000# diff_1277000_5967000# diff_1129000_5768000# GND efet w=328500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1008 diff_1119000_5759000# diff_1277000_5967000# diff_82000_3097000# GND efet w=154500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M1009 diff_82000_3097000# diff_1277000_5967000# diff_1129000_5768000# GND efet w=328000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1010 diff_94000_5193000# diff_1119000_5759000# diff_1119000_5759000# GND efet w=41000 l=11000
+ ad=-1.3245e+09 pd=1.23898e+08 as=0 ps=0 
M1011 diff_1277000_5967000# diff_1277000_5967000# diff_94000_5193000# GND efet w=29000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1012 diff_513000_5775000# diff_743000_5833000# diff_82000_3097000# GND efet w=122500 l=10500
+ ad=-5.97967e+08 pd=678000 as=0 ps=0 
M1013 diff_773000_5784000# diff_67000_5287000# diff_743000_5833000# GND efet w=15000 l=13000
+ ad=4.08e+08 pd=84000 as=-6.61967e+08 ps=552000 
M1014 diff_513000_5775000# diff_67000_5287000# diff_508000_5592000# GND efet w=22000 l=14000
+ ad=0 pd=0 as=3.15e+08 ps=110000 
M1015 diff_82000_3097000# diff_773000_5784000# diff_513000_5775000# GND efet w=113500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1016 diff_743000_5833000# diff_513000_5775000# diff_82000_3097000# GND efet w=98000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1017 diff_82000_3097000# diff_835000_5745000# diff_743000_5833000# GND efet w=116500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1018 diff_895000_5770000# diff_71000_4514000# diff_773000_5784000# GND efet w=15000 l=13000
+ ad=1.876e+09 pd=330000 as=0 ps=0 
M1019 diff_835000_5745000# diff_67000_5287000# diff_82000_3097000# GND efet w=67000 l=11000
+ ad=1.397e+09 pd=308000 as=0 ps=0 
M1020 diff_82000_3097000# diff_895000_5770000# diff_835000_5745000# GND efet w=70000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1021 diff_234000_3316000# diff_508000_5592000# diff_82000_3097000# GND efet w=132500 l=10500
+ ad=-1.81297e+09 pd=404000 as=0 ps=0 
M1022 diff_94000_5193000# diff_234000_3316000# diff_234000_3316000# GND efet w=15000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M1023 diff_513000_5775000# diff_513000_5775000# diff_94000_5193000# GND efet w=15000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M1024 diff_743000_5833000# diff_743000_5833000# diff_94000_5193000# GND efet w=14000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M1025 diff_82000_3097000# diff_968000_5799000# diff_895000_5770000# GND efet w=85000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1026 diff_895000_5770000# diff_895000_5770000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M1027 diff_82000_3097000# diff_616000_6169000# diff_968000_5799000# GND efet w=128000 l=12000
+ ad=0 pd=0 as=1.585e+09 ps=348000 
M1028 diff_94000_5193000# diff_616000_6169000# diff_616000_6169000# GND efet w=72000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1029 diff_1129000_5768000# diff_1119000_5759000# diff_94000_5193000# GND efet w=268000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1030 diff_1129000_5768000# diff_1119000_5759000# diff_94000_5193000# GND efet w=262000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1031 diff_1129000_5768000# diff_1119000_5759000# diff_94000_5193000# GND efet w=229000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1032 diff_1129000_5768000# diff_1119000_5759000# diff_94000_5193000# GND efet w=228500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1033 diff_1129000_5768000# diff_1119000_5759000# diff_94000_5193000# GND efet w=230000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1034 diff_1129000_5768000# diff_1119000_5759000# diff_94000_5193000# GND efet w=230000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1035 diff_1129000_5768000# diff_1119000_5759000# diff_94000_5193000# GND efet w=230000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1036 diff_835000_5745000# diff_835000_5745000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M1037 diff_1585000_6056000# diff_1585000_5875000# diff_82000_3097000# GND efet w=262000 l=11000
+ ad=3.98065e+08 pd=1.294e+06 as=0 ps=0 
M1038 diff_82000_3097000# diff_87000_5399000# diff_1585000_6056000# GND efet w=230000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1039 diff_1585000_6056000# diff_1647000_5846000# diff_82000_3097000# GND efet w=229000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1040 diff_82000_3097000# diff_196000_5469000# diff_1585000_6056000# GND efet w=229000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1041 diff_1585000_6056000# diff_1585000_6056000# diff_94000_5193000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1042 diff_968000_5799000# diff_968000_5799000# diff_94000_5193000# GND efet w=15000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M1043 diff_1747000_6169000# diff_82000_3097000# diff_82000_3097000# GND efet w=95500 l=15500
+ ad=-1.25684e+09 pd=3.486e+06 as=0 ps=0 
M1044 diff_82000_3097000# diff_94000_5193000# diff_2048000_5822000# GND efet w=72000 l=12000
+ ad=0 pd=0 as=1.524e+09 ps=320000 
M1045 diff_82000_3097000# diff_1747000_6169000# diff_300000_4193000# GND efet w=127000 l=12000
+ ad=0 pd=0 as=5.60327e+07 ps=836000 
M1046 diff_94000_5193000# diff_300000_4193000# diff_300000_4193000# GND efet w=16000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M1047 diff_572000_4609000# diff_67000_5287000# diff_1585000_5875000# GND efet w=17000 l=13000
+ ad=-6.04967e+08 pd=700000 as=2.82e+08 ps=100000 
M1048 diff_82000_3097000# diff_475000_5142000# diff_505000_5536000# GND efet w=97500 l=11500
+ ad=0 pd=0 as=-5.47935e+08 ps=1.086e+06 
M1049 diff_134000_5506000# diff_90000_5336000# diff_82000_3097000# GND efet w=215000 l=10000
+ ad=-1.54293e+09 pd=970000 as=0 ps=0 
M1050 diff_505000_5536000# diff_475000_5142000# diff_82000_3097000# GND efet w=96500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1051 diff_82000_3097000# diff_475000_5142000# diff_505000_5536000# GND efet w=107000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1052 diff_82000_3097000# diff_90000_5336000# diff_134000_5506000# GND efet w=78000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1053 diff_505000_5536000# diff_505000_5536000# diff_94000_5193000# GND efet w=30000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1054 diff_94000_5193000# diff_834000_5620000# diff_834000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=2.39033e+08 ps=916000 
M1055 diff_94000_5193000# diff_893000_5620000# diff_893000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=2.52033e+08 ps=920000 
M1056 diff_94000_5193000# diff_952000_5620000# diff_952000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=4.73033e+08 ps=936000 
M1057 diff_94000_5193000# diff_1011000_5620000# diff_1011000_5620000# GND efet w=13000 l=49000
+ ad=0 pd=0 as=1.12033e+08 ps=914000 
M1058 diff_94000_5193000# diff_760000_5560000# diff_760000_5560000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-8.39673e+07 ps=836000 
M1059 diff_796000_5586000# diff_796000_5586000# diff_94000_5193000# GND efet w=15000 l=49000
+ ad=-3.08967e+08 pd=806000 as=0 ps=0 
M1060 diff_94000_5193000# diff_854000_5586000# diff_854000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-5.48967e+08 ps=784000 
M1061 diff_94000_5193000# diff_913000_5586000# diff_913000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-4.12967e+08 ps=796000 
M1062 diff_94000_5193000# diff_972000_5586000# diff_972000_5586000# GND efet w=16000 l=49000
+ ad=0 pd=0 as=-3.47967e+08 ps=802000 
M1063 diff_94000_5193000# diff_1031000_5586000# diff_1031000_5586000# GND efet w=16000 l=49000
+ ad=0 pd=0 as=-9.79673e+07 ps=826000 
M1064 diff_94000_5193000# diff_1109000_5620000# diff_1109000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=2.76033e+08 ps=918000 
M1065 diff_94000_5193000# diff_1168000_5620000# diff_1168000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=4.68033e+08 ps=934000 
M1066 diff_94000_5193000# diff_1227000_5620000# diff_1227000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=1.50033e+08 ps=912000 
M1067 diff_94000_5193000# diff_1285000_5620000# diff_1285000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=3.23033e+08 ps=922000 
M1068 diff_94000_5193000# diff_1345000_5620000# diff_1345000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=1.27033e+08 ps=910000 
M1069 diff_94000_5193000# diff_1403000_5620000# diff_1403000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=2.54033e+08 ps=916000 
M1070 diff_1463000_5620000# diff_1463000_5620000# diff_94000_5193000# GND efet w=14000 l=49000
+ ad=3.49033e+08 pd=930000 as=0 ps=0 
M1071 diff_94000_5193000# diff_1521000_5620000# diff_1521000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=5.98033e+08 ps=948000 
M1072 diff_94000_5193000# diff_1129000_5586000# diff_1129000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-4.16967e+08 ps=796000 
M1073 diff_94000_5193000# diff_1187000_5586000# diff_1187000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-4.30967e+08 ps=794000 
M1074 diff_94000_5193000# diff_1247000_5586000# diff_1247000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-3.91967e+08 ps=798000 
M1075 diff_94000_5193000# diff_1305000_5586000# diff_1305000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-3.75967e+08 ps=800000 
M1076 diff_94000_5193000# diff_1365000_5586000# diff_1365000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-1.45967e+08 ps=822000 
M1077 diff_94000_5193000# diff_1423000_5586000# diff_1423000_5586000# GND efet w=16000 l=49000
+ ad=0 pd=0 as=-1.78967e+08 ps=818000 
M1078 diff_94000_5193000# diff_1483000_5586000# diff_1483000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-4.51967e+08 ps=792000 
M1079 diff_94000_5193000# diff_1541000_5586000# diff_1541000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-4.78967e+08 ps=792000 
M1080 diff_94000_5193000# diff_1618000_5620000# diff_1618000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=2.52033e+08 ps=922000 
M1081 diff_94000_5193000# diff_1677000_5620000# diff_1677000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=4.19033e+08 ps=932000 
M1082 diff_94000_5193000# diff_1736000_5620000# diff_1736000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=1.57033e+08 ps=912000 
M1083 diff_94000_5193000# diff_1794000_5620000# diff_1794000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=3.62033e+08 ps=926000 
M1084 diff_2072000_5822000# diff_71000_4514000# diff_2048000_5822000# GND efet w=14000 l=13000
+ ad=1.12e+08 pd=44000 as=0 ps=0 
M1085 diff_2093000_5822000# diff_67000_5287000# diff_2072000_5822000# GND efet w=14000 l=13000
+ ad=4.77e+08 pd=108000 as=0 ps=0 
M1086 diff_2093000_5822000# diff_1747000_6169000# diff_1747000_6169000# GND efet w=12000 l=76000
+ ad=0 pd=0 as=0 ps=0 
M1087 diff_82000_3097000# diff_82000_3097000# diff_82000_3097000# GND efet w=2000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1088 diff_82000_3097000# diff_82000_3097000# diff_67000_5287000# GND efet w=80000 l=15000
+ ad=0 pd=0 as=-1.23493e+09 ps=712000 
M1089 diff_2158000_5725000# diff_2048000_5822000# diff_1747000_6169000# GND efet w=14000 l=13000
+ ad=1.82e+08 pd=54000 as=0 ps=0 
M1090 diff_2195000_5725000# diff_82000_3097000# diff_2158000_5725000# GND efet w=14000 l=24000
+ ad=1.93013e+09 pd=3.34e+06 as=0 ps=0 
M1091 diff_82000_3097000# diff_82000_3097000# diff_2195000_5725000# GND efet w=82000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M1092 diff_2522000_5769000# diff_2195000_5725000# diff_82000_3097000# GND efet w=139000 l=12000
+ ad=-1.83597e+09 pd=462000 as=0 ps=0 
M1093 diff_2622000_5835000# diff_2612000_5826000# diff_82000_3097000# GND efet w=126000 l=10000
+ ad=1.945e+09 pd=438000 as=0 ps=0 
M1094 diff_82000_3097000# diff_1580000_4324000# diff_2747000_5771000# GND efet w=71500 l=10500
+ ad=0 pd=0 as=1.558e+09 ps=348000 
M1095 diff_2622000_5835000# diff_2622000_5835000# diff_94000_5193000# GND efet w=14000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M1096 diff_2612000_5826000# diff_67000_5287000# diff_2522000_5769000# GND efet w=14000 l=13000
+ ad=3.4e+08 pd=104000 as=0 ps=0 
M1097 diff_2522000_5769000# diff_2522000_5769000# diff_94000_5193000# GND efet w=15000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M1098 diff_82000_3097000# diff_2622000_5835000# diff_2747000_5771000# GND efet w=66000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1099 diff_2840000_5927000# diff_2834000_5760000# diff_82000_3097000# GND efet w=114000 l=11000
+ ad=-1.01967e+08 pd=804000 as=0 ps=0 
M1100 diff_82000_3097000# diff_93000_3550000# diff_2840000_5927000# GND efet w=111000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1101 diff_2840000_5927000# diff_2878000_5744000# diff_82000_3097000# GND efet w=113500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1102 diff_2878000_5744000# diff_2840000_5927000# diff_82000_3097000# GND efet w=128000 l=10000
+ ad=6.87033e+08 pd=918000 as=0 ps=0 
M1103 diff_2878000_5744000# diff_2984000_5745000# diff_82000_3097000# GND efet w=135500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M1104 diff_196000_5469000# diff_3100000_5786000# diff_82000_3097000# GND efet w=427500 l=9500
+ ad=1.44307e+09 pd=1.708e+06 as=0 ps=0 
M1105 diff_2747000_5771000# diff_2747000_5771000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M1106 diff_2834000_5760000# diff_71000_4514000# diff_2622000_5835000# GND efet w=15000 l=13000
+ ad=6.09e+08 pd=138000 as=0 ps=0 
M1107 diff_2840000_5927000# diff_2840000_5927000# diff_94000_5193000# GND efet w=16000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M1108 diff_2878000_5744000# diff_67000_5287000# diff_2834000_5760000# GND efet w=16000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M1109 diff_3100000_5786000# diff_67000_5287000# diff_2878000_5744000# GND efet w=36000 l=13000
+ ad=4.8e+08 pd=132000 as=0 ps=0 
M1110 diff_2747000_5771000# diff_71000_4514000# diff_2984000_5745000# GND efet w=14500 l=14500
+ ad=0 pd=0 as=8.03e+08 ps=162000 
M1111 diff_2984000_5745000# diff_67000_5287000# diff_2840000_5927000# GND efet w=15000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M1112 diff_196000_5469000# diff_93000_3550000# diff_82000_3097000# GND efet w=332000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1113 diff_3582000_5809000# diff_3504000_5808000# diff_82000_3097000# GND efet w=124500 l=10500
+ ad=-1.60897e+09 pd=504000 as=0 ps=0 
M1114 diff_196000_5469000# diff_93000_3550000# diff_82000_3097000# GND efet w=26000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1115 diff_196000_5469000# diff_93000_3550000# diff_82000_3097000# GND efet w=64000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1116 diff_93000_3550000# diff_3504000_5808000# diff_94000_5193000# GND efet w=27000 l=9000
+ ad=7.44033e+08 pd=726000 as=0 ps=0 
M1117 diff_2878000_5744000# diff_2878000_5744000# diff_94000_5193000# GND efet w=14000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M1118 diff_94000_5193000# diff_196000_5469000# diff_196000_5469000# GND efet w=27000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1119 diff_93000_3550000# diff_3504000_5808000# diff_94000_5193000# GND efet w=202500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M1120 diff_94000_5193000# diff_1943000_5620000# diff_1943000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=2.25033e+08 ps=918000 
M1121 diff_94000_5193000# diff_2001000_5620000# diff_2001000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=2.20033e+08 ps=912000 
M1122 diff_94000_5193000# diff_2060000_5620000# diff_2060000_5620000# GND efet w=13000 l=49000
+ ad=0 pd=0 as=2.80033e+08 ps=930000 
M1123 diff_94000_5193000# diff_2118000_5620000# diff_2118000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=5.11033e+08 ps=940000 
M1124 diff_94000_5193000# diff_1638000_5586000# diff_1638000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-5.02967e+08 ps=788000 
M1125 diff_94000_5193000# diff_1697000_5586000# diff_1697000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-1.49967e+08 ps=822000 
M1126 diff_94000_5193000# diff_1756000_5586000# diff_1756000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-2.23967e+08 ps=816000 
M1127 diff_94000_5193000# diff_1814000_5586000# diff_1814000_5586000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=-4.49967e+08 ps=794000 
M1128 diff_94000_5193000# diff_1963000_5586000# diff_1963000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-3.74967e+08 ps=802000 
M1129 diff_94000_5193000# diff_2021000_5586000# diff_2021000_5586000# GND efet w=16000 l=49000
+ ad=0 pd=0 as=-3.92967e+08 ps=798000 
M1130 diff_94000_5193000# diff_2080000_5586000# diff_2080000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-4.47967e+08 ps=794000 
M1131 diff_94000_5193000# diff_2138000_5586000# diff_2138000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-2.93967e+08 ps=808000 
M1132 diff_94000_5193000# diff_2217000_5620000# diff_2217000_5620000# GND efet w=16000 l=49000
+ ad=0 pd=0 as=3.62033e+08 ps=920000 
M1133 diff_94000_5193000# diff_2275000_5620000# diff_2275000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=6.29033e+08 ps=952000 
M1134 diff_94000_5193000# diff_2334000_5620000# diff_2334000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=3.11033e+08 ps=926000 
M1135 diff_94000_5193000# diff_2393000_5620000# diff_2393000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=2.63033e+08 ps=916000 
M1136 diff_93000_3550000# diff_3582000_5809000# diff_82000_3097000# GND efet w=368500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M1137 diff_1647000_5846000# diff_3694000_5840000# diff_3676000_5838000# GND efet w=108500 l=9500
+ ad=-1.89597e+09 pd=400000 as=1.70033e+08 ps=900000 
M1138 diff_3676000_5838000# diff_3694000_5840000# diff_1647000_5846000# GND efet w=161000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1139 diff_82000_3097000# diff_3756000_5781000# diff_3676000_5838000# GND efet w=151000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1140 diff_82000_3097000# diff_3756000_5781000# diff_3504000_5808000# GND efet w=184500 l=10500
+ ad=0 pd=0 as=2.139e+09 ps=426000 
M1141 diff_3582000_5809000# diff_3504000_5808000# diff_82000_3097000# GND efet w=34000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1142 diff_94000_5193000# diff_3582000_5809000# diff_3582000_5809000# GND efet w=14000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1143 diff_1647000_5846000# diff_1647000_5846000# diff_94000_5193000# GND efet w=14000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M1144 diff_1647000_5846000# diff_1647000_5846000# diff_1647000_5846000# GND efet w=500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M1145 diff_3676000_5838000# diff_3756000_5781000# diff_82000_3097000# GND efet w=101000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1146 diff_82000_3097000# diff_3883000_5843000# diff_3871000_5818000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=3.94033e+08 ps=870000 
M1147 diff_3902000_5736000# diff_3871000_5818000# diff_82000_3097000# GND efet w=57000 l=10000
+ ad=-1.38097e+09 pd=508000 as=0 ps=0 
M1148 diff_82000_3097000# diff_3883000_5843000# diff_3871000_5818000# GND efet w=81000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1149 diff_82000_3097000# diff_3961000_5823000# diff_3902000_5736000# GND efet w=121000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1150 diff_82000_3097000# diff_3961000_5823000# diff_3883000_5843000# GND efet w=70500 l=10500
+ ad=0 pd=0 as=-1.99897e+09 ps=416000 
M1151 diff_3902000_5736000# diff_3871000_5818000# diff_82000_3097000# GND efet w=61500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M1152 diff_82000_3097000# diff_67000_5287000# diff_3883000_5843000# GND efet w=77000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1153 diff_3871000_5818000# diff_3902000_5736000# diff_82000_3097000# GND efet w=117000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1154 diff_3883000_5843000# diff_3883000_5843000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M1155 diff_3961000_5823000# diff_67000_5287000# diff_3871000_5818000# GND efet w=30000 l=14000
+ ad=9.66e+08 pd=236000 as=0 ps=0 
M1156 diff_82000_3097000# diff_4197000_5802000# diff_3694000_5840000# GND efet w=104500 l=10500
+ ad=0 pd=0 as=-2.05897e+09 ps=470000 
M1157 diff_3504000_5808000# diff_3504000_5808000# diff_94000_5193000# GND efet w=14000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M1158 diff_3871000_5818000# diff_67000_5287000# diff_3756000_5781000# GND efet w=29000 l=13000
+ ad=0 pd=0 as=3.71e+08 ps=114000 
M1159 diff_3902000_5736000# diff_3902000_5736000# diff_94000_5193000# GND efet w=15000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M1160 diff_3694000_5840000# diff_71000_4514000# diff_3961000_5823000# GND efet w=22000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M1161 diff_82000_3097000# diff_4055000_6170000# diff_4197000_5802000# GND efet w=130500 l=12500
+ ad=0 pd=0 as=1.555e+09 ps=328000 
M1162 diff_4426000_5700000# diff_4355000_5716000# diff_82000_3097000# GND efet w=180500 l=11500
+ ad=1.642e+09 pd=280000 as=0 ps=0 
M1163 diff_94000_5193000# diff_3871000_5818000# diff_3871000_5818000# GND efet w=15000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M1164 diff_3694000_5840000# diff_3694000_5840000# diff_3694000_5840000# GND efet w=1000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1165 diff_3694000_5840000# diff_3694000_5840000# diff_94000_5193000# GND efet w=14000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M1166 diff_4055000_6170000# diff_82000_3097000# diff_82000_3097000# GND efet w=81000 l=14000
+ ad=-1.40687e+09 pd=2.734e+06 as=0 ps=0 
M1167 diff_87000_5399000# diff_4355000_5716000# diff_82000_3097000# GND efet w=190500 l=11500
+ ad=2.09803e+09 pd=930000 as=0 ps=0 
M1168 diff_87000_5399000# diff_4355000_5716000# diff_82000_3097000# GND efet w=230500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1169 diff_94000_5193000# diff_4426000_5700000# diff_87000_5399000# GND efet w=321500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1170 diff_4197000_5802000# diff_4197000_5802000# diff_94000_5193000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M1171 diff_4055000_6170000# diff_4055000_6170000# diff_94000_5193000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M1172 diff_94000_5193000# diff_4426000_5700000# diff_87000_5399000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1173 diff_4426000_5700000# diff_4426000_5700000# diff_94000_5193000# GND efet w=13000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1174 diff_4355000_5716000# diff_4355000_5716000# diff_94000_5193000# GND efet w=14000 l=14000
+ ad=1.697e+09 pd=324000 as=0 ps=0 
M1175 diff_82000_3097000# diff_4397000_6170000# diff_4355000_5716000# GND efet w=135500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M1176 diff_4397000_6170000# diff_82000_3097000# diff_82000_3097000# GND efet w=82000 l=14000
+ ad=-2.49869e+08 pd=2.83e+06 as=0 ps=0 
M1177 diff_82000_3097000# diff_82000_3097000# diff_82000_3097000# GND efet w=1000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1178 diff_5256000_3172000# diff_5405000_5991000# diff_82000_3097000# GND efet w=701000 l=10000
+ ad=-7.98692e+07 pd=1.994e+06 as=0 ps=0 
M1179 diff_5256000_3172000# diff_5405000_5991000# diff_82000_3097000# GND efet w=170000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1180 diff_82000_3097000# diff_5771000_6154000# diff_5760000_6139000# GND efet w=405500 l=10500
+ ad=0 pd=0 as=1.33907e+09 ps=1.49e+06 
M1181 diff_5429000_5897000# diff_5452000_5801000# diff_82000_3097000# GND efet w=206000 l=11000
+ ad=1.607e+09 pd=282000 as=0 ps=0 
M1182 diff_82000_3097000# diff_5405000_5991000# diff_5256000_3172000# GND efet w=77500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M1183 diff_82000_3097000# diff_5405000_5991000# diff_5256000_3172000# GND efet w=15000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1184 diff_82000_3097000# diff_134000_5506000# diff_5760000_6139000# GND efet w=383500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1185 diff_5429000_5897000# diff_5429000_5897000# diff_94000_5193000# GND efet w=14000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1186 diff_5771000_6154000# diff_67000_5287000# diff_5508000_5788000# GND efet w=36000 l=15000
+ ad=4.29e+08 pd=124000 as=-1.10697e+09 ps=698000 
M1187 diff_5405000_5991000# diff_5172000_5734000# diff_82000_3097000# GND efet w=74500 l=11500
+ ad=1.63e+09 pd=342000 as=0 ps=0 
M1188 diff_5258000_5769000# diff_5429000_5897000# diff_5405000_5991000# GND efet w=76500 l=11500
+ ad=-1.89593e+09 pd=914000 as=0 ps=0 
M1189 diff_94000_5193000# diff_2482000_5620000# diff_2482000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=4.07033e+08 ps=936000 
M1190 diff_94000_5193000# diff_2540000_5620000# diff_2540000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=3.21033e+08 ps=922000 
M1191 diff_94000_5193000# diff_2599000_5620000# diff_2599000_5620000# GND efet w=13000 l=49000
+ ad=0 pd=0 as=1.72033e+08 ps=912000 
M1192 diff_94000_5193000# diff_2658000_5620000# diff_2658000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=3.61033e+08 ps=926000 
M1193 diff_94000_5193000# diff_2237000_5586000# diff_2237000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-3.03967e+08 ps=808000 
M1194 diff_94000_5193000# diff_2295000_5586000# diff_2295000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-5.12967e+08 ps=786000 
M1195 diff_94000_5193000# diff_2354000_5586000# diff_2354000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-1.83967e+08 ps=818000 
M1196 diff_94000_5193000# diff_2413000_5586000# diff_2413000_5586000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=-4.40967e+08 ps=794000 
M1197 diff_94000_5193000# diff_2502000_5586000# diff_2502000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-1.55967e+08 ps=820000 
M1198 diff_94000_5193000# diff_2560000_5586000# diff_2560000_5586000# GND efet w=16000 l=49000
+ ad=0 pd=0 as=-3.34967e+08 ps=804000 
M1199 diff_94000_5193000# diff_2619000_5586000# diff_2619000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-2.25967e+08 ps=814000 
M1200 diff_94000_5193000# diff_2678000_5586000# diff_2678000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-2.87967e+08 ps=808000 
M1201 diff_94000_5193000# diff_2756000_5620000# diff_2756000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=2.61033e+08 ps=916000 
M1202 diff_94000_5193000# diff_2814000_5620000# diff_2814000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=4.00033e+08 ps=930000 
M1203 diff_94000_5193000# diff_2873000_5620000# diff_2873000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=3.25033e+08 ps=928000 
M1204 diff_94000_5193000# diff_2932000_5620000# diff_2932000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=3.25033e+08 ps=922000 
M1205 diff_2991000_5620000# diff_2991000_5620000# diff_94000_5193000# GND efet w=13000 l=49000
+ ad=1.29033e+08 pd=916000 as=0 ps=0 
M1206 diff_3050000_5620000# diff_3050000_5620000# diff_94000_5193000# GND efet w=14000 l=49000
+ ad=4.08033e+08 pd=936000 as=0 ps=0 
M1207 diff_94000_5193000# diff_3109000_5620000# diff_3109000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=1.82033e+08 ps=910000 
M1208 diff_94000_5193000# diff_2776000_5586000# diff_2776000_5586000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=-4.15967e+08 ps=798000 
M1209 diff_94000_5193000# diff_2834000_5586000# diff_2834000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-2.59967e+08 ps=812000 
M1210 diff_94000_5193000# diff_2893000_5586000# diff_2893000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-2.01967e+08 ps=816000 
M1211 diff_94000_5193000# diff_2952000_5586000# diff_2952000_5586000# GND efet w=16000 l=49000
+ ad=0 pd=0 as=-3.25967e+08 ps=804000 
M1212 diff_94000_5193000# diff_3011000_5586000# diff_3011000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-2.07967e+08 ps=816000 
M1213 diff_94000_5193000# diff_3168000_5620000# diff_3168000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=2.28033e+08 ps=918000 
M1214 diff_94000_5193000# diff_3070000_5586000# diff_3070000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-3.25967e+08 ps=804000 
M1215 diff_94000_5193000# diff_3129000_5586000# diff_3129000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-1.22967e+08 ps=826000 
M1216 diff_94000_5193000# diff_3188000_5586000# diff_3188000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-2.94967e+08 ps=808000 
M1217 diff_94000_5193000# diff_3265000_5620000# diff_3265000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=4.39033e+08 ps=934000 
M1218 diff_3323000_5620000# diff_3323000_5620000# diff_94000_5193000# GND efet w=14000 l=49000
+ ad=2.85033e+08 pd=924000 as=0 ps=0 
M1219 diff_94000_5193000# diff_3382000_5620000# diff_3382000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=3.54033e+08 ps=932000 
M1220 diff_94000_5193000# diff_3441000_5620000# diff_3441000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=2.51033e+08 ps=916000 
M1221 diff_94000_5193000# diff_3500000_5620000# diff_3500000_5620000# GND efet w=13000 l=49000
+ ad=0 pd=0 as=1.29033e+08 ps=916000 
M1222 diff_94000_5193000# diff_3559000_5620000# diff_3559000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=5.37033e+08 ps=942000 
M1223 diff_94000_5193000# diff_3285000_5586000# diff_3285000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-4.19967e+08 ps=796000 
M1224 diff_94000_5193000# diff_3343000_5586000# diff_3343000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-3.39967e+08 ps=804000 
M1225 diff_94000_5193000# diff_3402000_5586000# diff_3402000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-4.68967e+08 ps=792000 
M1226 diff_94000_5193000# diff_3461000_5586000# diff_3461000_5586000# GND efet w=16000 l=49000
+ ad=0 pd=0 as=-2.82967e+08 ps=810000 
M1227 diff_94000_5193000# diff_3618000_5620000# diff_3618000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=2.32033e+08 ps=914000 
M1228 diff_94000_5193000# diff_3677000_5620000# diff_3677000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=5.33033e+08 ps=942000 
M1229 diff_94000_5193000# diff_3520000_5586000# diff_3520000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-4.48967e+08 ps=794000 
M1230 diff_94000_5193000# diff_3579000_5586000# diff_3579000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-2.08967e+08 ps=816000 
M1231 diff_94000_5193000# diff_3638000_5586000# diff_3638000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-1.66967e+08 ps=820000 
M1232 diff_94000_5193000# diff_3697000_5586000# diff_3697000_5586000# GND efet w=16000 l=49000
+ ad=0 pd=0 as=-4.79967e+08 ps=788000 
M1233 diff_94000_5193000# diff_3775000_5620000# diff_3775000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=2.93033e+08 ps=920000 
M1234 diff_94000_5193000# diff_3833000_5620000# diff_3833000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=4.83033e+08 ps=938000 
M1235 diff_94000_5193000# diff_3892000_5620000# diff_3892000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=3.11033e+08 ps=928000 
M1236 diff_94000_5193000# diff_3951000_5620000# diff_3951000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=3.82033e+08 ps=928000 
M1237 diff_4010000_5620000# diff_4010000_5620000# diff_94000_5193000# GND efet w=13000 l=49000
+ ad=2.97033e+08 pd=932000 as=0 ps=0 
M1238 diff_94000_5193000# diff_4069000_5620000# diff_4069000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=4.51033e+08 ps=940000 
M1239 diff_94000_5193000# diff_4128000_5620000# diff_4128000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=3.66033e+08 ps=928000 
M1240 diff_94000_5193000# diff_3795000_5586000# diff_3795000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-2.52967e+08 ps=812000 
M1241 diff_94000_5193000# diff_3853000_5586000# diff_3853000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-3.85967e+08 ps=800000 
M1242 diff_94000_5193000# diff_3912000_5586000# diff_3912000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-3.94967e+08 ps=798000 
M1243 diff_94000_5193000# diff_3971000_5586000# diff_3971000_5586000# GND efet w=16000 l=49000
+ ad=0 pd=0 as=-3.78967e+08 ps=800000 
M1244 diff_94000_5193000# diff_4030000_5586000# diff_4030000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-3.50967e+08 ps=802000 
M1245 diff_94000_5193000# diff_4187000_5620000# diff_4187000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=1.19033e+08 ps=908000 
M1246 diff_94000_5193000# diff_4089000_5586000# diff_4089000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-5.48967e+08 ps=784000 
M1247 diff_94000_5193000# diff_4148000_5586000# diff_4148000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-2.19967e+08 ps=816000 
M1248 diff_94000_5193000# diff_4207000_5586000# diff_4207000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-2.33967e+08 ps=814000 
M1249 diff_94000_5193000# diff_4287000_5620000# diff_4287000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=3.48033e+08 ps=930000 
M1250 diff_94000_5193000# diff_4345000_5620000# diff_4345000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=1.82033e+08 ps=916000 
M1251 diff_94000_5193000# diff_4404000_5620000# diff_4404000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=2.47033e+08 ps=920000 
M1252 diff_94000_5193000# diff_4306000_5586000# diff_4306000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-3.94967e+08 ps=798000 
M1253 diff_94000_5193000# diff_4463000_5620000# diff_4463000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=2.07033e+08 ps=912000 
M1254 diff_94000_5193000# diff_4522000_5620000# diff_4522000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=4.22033e+08 ps=938000 
M1255 diff_4581000_5620000# diff_4581000_5620000# diff_94000_5193000# GND efet w=14000 l=49000
+ ad=2.91033e+08 pd=926000 as=0 ps=0 
M1256 diff_82000_3097000# diff_82000_3097000# diff_71000_4514000# GND efet w=82000 l=15000
+ ad=0 pd=0 as=1.20803e+09 ps=524000 
M1257 diff_5066000_5899000# diff_82000_3097000# diff_82000_3097000# GND efet w=83000 l=15000
+ ad=-2.12869e+08 pd=2.772e+06 as=0 ps=0 
M1258 diff_82000_3097000# diff_5066000_5899000# diff_5172000_5734000# GND efet w=312500 l=10500
+ ad=0 pd=0 as=7.77033e+08 ps=816000 
M1259 diff_82000_3097000# diff_5172000_5734000# diff_5258000_5769000# GND efet w=381500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1260 diff_94000_5193000# diff_5172000_5734000# diff_5172000_5734000# GND efet w=26000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1261 diff_5403000_5746000# diff_5258000_5769000# diff_82000_3097000# GND efet w=249500 l=11500
+ ad=1.66e+09 pd=360000 as=0 ps=0 
M1262 diff_5256000_3172000# diff_5403000_5746000# diff_94000_5193000# GND efet w=115000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M1263 diff_5256000_3172000# diff_5403000_5746000# diff_94000_5193000# GND efet w=22000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M1264 diff_94000_5193000# diff_5403000_5746000# diff_5256000_3172000# GND efet w=277000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1265 diff_94000_5193000# diff_67000_5287000# diff_94000_5193000# GND efet w=12500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M1266 diff_5927000_6129000# diff_5760000_6139000# diff_82000_3097000# GND efet w=840000 l=10000
+ ad=1.44229e+08 pd=4.164e+06 as=0 ps=0 
M1267 diff_5927000_6129000# diff_5760000_6139000# diff_82000_3097000# GND efet w=599000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1268 diff_5774000_5846000# diff_5774000_5846000# diff_5774000_5846000# GND efet w=500 l=2500
+ ad=2.00307e+09 pd=1.592e+06 as=0 ps=0 
M1269 diff_5927000_6129000# diff_5774000_5846000# diff_94000_5193000# GND efet w=483000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1270 diff_94000_5193000# diff_5760000_6139000# diff_5760000_6139000# GND efet w=37000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1271 diff_94000_5193000# diff_5774000_5846000# diff_5774000_5846000# GND efet w=43000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1272 diff_5774000_5846000# diff_5760000_6139000# diff_82000_3097000# GND efet w=495000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1273 diff_94000_5193000# diff_5774000_5846000# diff_5927000_6129000# GND efet w=240500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1274 diff_5774000_5846000# diff_134000_5506000# diff_82000_3097000# GND efet w=127000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1275 diff_94000_5193000# diff_5774000_5846000# diff_5927000_6129000# GND efet w=242500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M1276 diff_5774000_5846000# diff_134000_5506000# diff_82000_3097000# GND efet w=271000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1277 diff_5927000_6129000# diff_5774000_5846000# diff_94000_5193000# GND efet w=681000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1278 diff_5488000_5788000# diff_5403000_5746000# diff_5452000_5801000# GND efet w=37000 l=14000
+ ad=2.59e+08 pd=88000 as=5.88e+08 ps=132000 
M1279 diff_5508000_5788000# diff_67000_5287000# diff_5488000_5788000# GND efet w=37000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M1280 diff_5403000_5746000# diff_5403000_5746000# diff_94000_5193000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1281 diff_5258000_5769000# diff_5258000_5769000# diff_94000_5193000# GND efet w=36000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1282 diff_4477000_4816000# diff_71000_4514000# diff_6104000_5744000# GND efet w=22000 l=14000
+ ad=1.43703e+09 pd=1.008e+06 as=3.54e+08 ps=120000 
M1283 diff_94000_5193000# diff_5508000_5788000# diff_5508000_5788000# GND efet w=15000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1284 diff_5508000_5788000# diff_6104000_5744000# diff_82000_3097000# GND efet w=161000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1285 diff_94000_5193000# diff_4729000_5620000# diff_4729000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=4.14033e+08 ps=938000 
M1286 diff_94000_5193000# diff_4787000_5620000# diff_4787000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=1.30033e+08 ps=910000 
M1287 diff_94000_5193000# diff_4846000_5620000# diff_4846000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=3.72033e+08 ps=934000 
M1288 diff_94000_5193000# diff_4365000_5586000# diff_4365000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-4.97967e+08 ps=788000 
M1289 diff_94000_5193000# diff_4424000_5586000# diff_4424000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-3.22967e+08 ps=806000 
M1290 diff_94000_5193000# diff_4483000_5586000# diff_4483000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-3.05967e+08 ps=808000 
M1291 diff_94000_5193000# diff_4542000_5586000# diff_4542000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-4.78967e+08 ps=790000 
M1292 diff_94000_5193000# diff_4601000_5586000# diff_4601000_5586000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=-4.03967e+08 ps=798000 
M1293 diff_94000_5193000# diff_4749000_5586000# diff_4749000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-3.94967e+08 ps=798000 
M1294 diff_4905000_5620000# diff_4905000_5620000# diff_94000_5193000# GND efet w=14000 l=49000
+ ad=3.36033e+08 pd=930000 as=0 ps=0 
M1295 diff_94000_5193000# diff_4807000_5586000# diff_4807000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-3.31967e+08 ps=804000 
M1296 diff_94000_5193000# diff_4866000_5586000# diff_4866000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-2.79967e+08 ps=808000 
M1297 diff_94000_5193000# diff_4925000_5586000# diff_4925000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-3.26967e+08 ps=804000 
M1298 diff_94000_5193000# diff_5003000_5620000# diff_5003000_5620000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=2.49033e+08 ps=916000 
M1299 diff_94000_5193000# diff_5061000_5620000# diff_5061000_5620000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=1.81033e+08 ps=916000 
M1300 diff_774000_5478000# diff_774000_5478000# diff_94000_5193000# GND efet w=16000 l=10000
+ ad=6.40033e+08 pd=954000 as=0 ps=0 
M1301 diff_774000_5478000# diff_5251000_5061000# diff_82000_3097000# GND efet w=184000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1302 diff_774000_5478000# diff_5500000_5677000# diff_82000_3097000# GND efet w=191000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1303 diff_82000_3097000# diff_5501000_5645000# diff_5500000_5677000# GND efet w=103500 l=9500
+ ad=0 pd=0 as=-1.22697e+09 ps=710000 
M1304 diff_5500000_5677000# diff_5500000_5677000# diff_5500000_5677000# GND efet w=500 l=1500
+ ad=0 pd=0 as=0 ps=0 
M1305 diff_82000_3097000# diff_5251000_5061000# diff_774000_5447000# GND efet w=181500 l=10500
+ ad=0 pd=0 as=2.13903e+09 ps=954000 
M1306 diff_774000_5447000# diff_5501000_5645000# diff_82000_3097000# GND efet w=181000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1307 diff_94000_5193000# diff_5023000_5586000# diff_5023000_5586000# GND efet w=15000 l=49000
+ ad=0 pd=0 as=-4.82967e+08 ps=790000 
M1308 diff_94000_5193000# diff_774000_5447000# diff_774000_5447000# GND efet w=15000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1309 diff_94000_5193000# diff_5081000_5586000# diff_5081000_5586000# GND efet w=14000 l=49000
+ ad=0 pd=0 as=-6.10967e+08 ps=776000 
M1310 diff_134000_5506000# diff_134000_5506000# diff_94000_5193000# GND efet w=27000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1311 diff_505000_5536000# diff_401000_4712000# diff_82000_3097000# GND efet w=142000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1312 diff_760000_5560000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1313 diff_796000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1314 diff_834000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1315 diff_854000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1316 diff_893000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1317 diff_913000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1318 diff_952000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1319 diff_972000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1320 diff_1011000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1321 diff_1031000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1322 diff_1109000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1323 diff_1129000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1324 diff_1168000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1325 diff_1187000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1326 diff_1227000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1327 diff_1247000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1328 diff_1285000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1329 diff_1305000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1330 diff_1345000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1331 diff_1365000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1332 diff_1403000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1333 diff_1423000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1334 diff_1463000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1335 diff_1483000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1336 diff_1521000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1337 diff_1541000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1338 diff_1618000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1339 diff_1638000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1340 diff_1677000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1341 diff_1697000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1342 diff_1736000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1343 diff_1756000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1344 diff_1794000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1345 diff_1814000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1346 diff_1943000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1347 diff_1963000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1348 diff_2001000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1349 diff_2021000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1350 diff_2060000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1351 diff_2080000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1352 diff_2118000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1353 diff_2138000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1354 diff_2217000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1355 diff_2237000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1356 diff_2275000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1357 diff_2295000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1358 diff_2334000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1359 diff_2354000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1360 diff_2393000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1361 diff_2413000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1362 diff_2482000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1363 diff_2502000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1364 diff_2540000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1365 diff_2560000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1366 diff_2599000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1367 diff_2619000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1368 diff_2658000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1369 diff_2678000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1370 diff_2756000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1371 diff_2776000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1372 diff_2814000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1373 diff_2834000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1374 diff_2873000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1375 diff_2893000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1376 diff_2932000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1377 diff_2952000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1378 diff_2991000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1379 diff_3011000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1380 diff_3050000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1381 diff_3070000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1382 diff_3109000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1383 diff_3129000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1384 diff_3168000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1385 diff_3188000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1386 diff_3265000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1387 diff_3285000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1388 diff_3323000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1389 diff_3343000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1390 diff_3382000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1391 diff_3402000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1392 diff_3441000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1393 diff_3461000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1394 diff_3500000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1395 diff_3520000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1396 diff_3559000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1397 diff_3579000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1398 diff_3618000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1399 diff_3638000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1400 diff_3677000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1401 diff_3697000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1402 diff_3775000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1403 diff_3795000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1404 diff_3833000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1405 diff_3853000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1406 diff_3892000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1407 diff_3912000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1408 diff_3951000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1409 diff_3971000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1410 diff_4010000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1411 diff_4030000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1412 diff_4069000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1413 diff_4089000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1414 diff_4128000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1415 diff_4148000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1416 diff_4187000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1417 diff_4207000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1418 diff_4287000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1419 diff_4306000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1420 diff_4345000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1421 diff_4365000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1422 diff_4404000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1423 diff_4424000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1424 diff_4463000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1425 diff_4483000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1426 diff_4522000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1427 diff_4542000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1428 diff_4581000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1429 diff_4601000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1430 diff_4729000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1431 diff_4749000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1432 diff_4787000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1433 diff_4807000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1434 diff_4846000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1435 diff_4866000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1436 diff_4905000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1437 diff_4925000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1438 diff_5003000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1439 diff_5023000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1440 diff_5061000_5620000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1441 diff_5081000_5586000# diff_475000_5142000# diff_94000_5193000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1442 diff_90000_5336000# diff_196000_5469000# diff_82000_3097000# GND efet w=234000 l=11000
+ ad=1.5181e+09 pd=1.804e+06 as=0 ps=0 
M1443 diff_94000_5193000# diff_90000_5336000# diff_90000_5336000# GND efet w=45000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1444 diff_82000_3097000# diff_401000_4712000# diff_505000_5536000# GND efet w=142000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1445 diff_82000_3097000# diff_774000_5478000# diff_760000_5560000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1446 diff_82000_3097000# diff_774000_5478000# diff_893000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1447 diff_82000_3097000# diff_774000_5478000# diff_972000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1448 diff_82000_3097000# diff_774000_5478000# diff_1031000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1449 diff_82000_3097000# diff_774000_5478000# diff_1168000_5620000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1450 diff_82000_3097000# diff_774000_5478000# diff_1227000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1451 diff_82000_3097000# diff_774000_5478000# diff_1365000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1452 diff_82000_3097000# diff_774000_5478000# diff_1423000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1453 diff_82000_3097000# diff_774000_5478000# diff_1521000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1454 diff_82000_3097000# diff_774000_5478000# diff_1677000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1455 diff_82000_3097000# diff_774000_5478000# diff_2118000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1456 diff_82000_3097000# diff_774000_5478000# diff_2275000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1457 diff_82000_3097000# diff_774000_5478000# diff_2354000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1458 diff_82000_3097000# diff_774000_5478000# diff_2502000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1459 diff_82000_3097000# diff_774000_5478000# diff_2678000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1460 diff_82000_3097000# diff_774000_5478000# diff_2893000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1461 diff_82000_3097000# diff_774000_5478000# diff_3011000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1462 diff_82000_3097000# diff_774000_5478000# diff_3070000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1463 diff_82000_3097000# diff_774000_5478000# diff_3129000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1464 diff_82000_3097000# diff_774000_5478000# diff_3168000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1465 diff_82000_3097000# diff_774000_5478000# diff_3265000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1466 diff_82000_3097000# diff_774000_5478000# diff_3559000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1467 diff_82000_3097000# diff_774000_5478000# diff_3579000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1468 diff_82000_3097000# diff_774000_5478000# diff_3638000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1469 diff_82000_3097000# diff_774000_5478000# diff_3892000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1470 diff_82000_3097000# diff_774000_5478000# diff_3912000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1471 diff_82000_3097000# diff_774000_5478000# diff_4010000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1472 diff_82000_3097000# diff_774000_5478000# diff_4306000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1473 diff_82000_3097000# diff_774000_5478000# diff_4807000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1474 diff_5500000_5677000# diff_5500000_5677000# diff_94000_5193000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M1475 diff_82000_3097000# diff_5699000_5645000# diff_5501000_5645000# GND efet w=103000 l=10000
+ ad=0 pd=0 as=-9.80967e+08 ps=624000 
M1476 diff_5500000_5677000# diff_5953000_5146000# diff_5699000_5645000# GND efet w=15000 l=13000
+ ad=0 pd=0 as=6.15e+08 ps=148000 
M1477 diff_5953000_5146000# diff_5953000_5146000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=1.327e+09 pd=320000 as=0 ps=0 
M1478 diff_5953000_5146000# diff_475000_5142000# diff_82000_3097000# GND efet w=66000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1479 diff_94000_5193000# diff_5501000_5645000# diff_5501000_5645000# GND efet w=15000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M1480 diff_5501000_5645000# diff_5501000_5645000# diff_5501000_5645000# GND efet w=1000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1481 diff_5699000_5645000# diff_475000_5142000# diff_5971000_5631000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=-1.72997e+09 ps=524000 
M1482 diff_5971000_5631000# diff_5971000_5631000# diff_94000_5193000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M1483 diff_82000_3097000# diff_6061000_5631000# diff_5971000_5631000# GND efet w=117500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1484 diff_82000_3097000# diff_774000_5478000# diff_5003000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1485 diff_82000_3097000# diff_87000_5399000# diff_90000_5336000# GND efet w=85000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1486 diff_82000_3097000# diff_87000_5399000# diff_90000_5336000# GND efet w=114000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1487 diff_90000_5336000# diff_196000_5469000# diff_82000_3097000# GND efet w=51500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1488 diff_90000_5336000# diff_87000_5399000# diff_82000_3097000# GND efet w=85000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1489 diff_401000_4712000# diff_401000_4712000# diff_94000_5193000# GND efet w=18000 l=14000
+ ad=4.26033e+08 pd=812000 as=0 ps=0 
M1490 diff_774000_5420000# diff_774000_5420000# diff_94000_5193000# GND efet w=16000 l=10000
+ ad=-1.55193e+09 pd=1.394e+06 as=0 ps=0 
M1491 diff_774000_5420000# diff_5251000_5061000# diff_82000_3097000# GND efet w=184000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1492 diff_774000_5420000# diff_5500000_5602000# diff_82000_3097000# GND efet w=191000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1493 diff_82000_3097000# diff_5501000_5570000# diff_5500000_5602000# GND efet w=103500 l=9500
+ ad=0 pd=0 as=-1.22697e+09 ps=710000 
M1494 diff_5500000_5602000# diff_5500000_5602000# diff_5500000_5602000# GND efet w=500 l=1500
+ ad=0 pd=0 as=0 ps=0 
M1495 diff_82000_3097000# diff_5251000_5061000# diff_774000_5389000# GND efet w=181500 l=10500
+ ad=0 pd=0 as=2.13903e+09 ps=954000 
M1496 diff_774000_5389000# diff_5501000_5570000# diff_82000_3097000# GND efet w=181000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1497 diff_94000_5193000# diff_774000_5389000# diff_774000_5389000# GND efet w=15000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1498 diff_5500000_5602000# diff_5500000_5602000# diff_94000_5193000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M1499 diff_82000_3097000# diff_5699000_5570000# diff_5501000_5570000# GND efet w=103000 l=10000
+ ad=0 pd=0 as=-9.80967e+08 ps=624000 
M1500 diff_5500000_5602000# diff_5953000_5146000# diff_5699000_5570000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=6e+08 ps=146000 
M1501 diff_5971000_5631000# diff_6021000_5609000# diff_82000_3097000# GND efet w=103000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1502 diff_6175000_5603000# diff_71000_4514000# diff_6021000_5609000# GND efet w=22000 l=14000
+ ad=-1.45397e+09 pd=588000 as=3.41e+08 ps=96000 
M1503 diff_6175000_5603000# diff_6175000_5603000# diff_6175000_5603000# GND efet w=2000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M1504 diff_94000_5193000# diff_6175000_5603000# diff_6175000_5603000# GND efet w=14000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M1505 diff_6175000_5603000# diff_5618000_2892000# diff_82000_3097000# GND efet w=128000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1506 diff_94000_5193000# diff_5501000_5570000# diff_5501000_5570000# GND efet w=15000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M1507 diff_5501000_5570000# diff_5501000_5570000# diff_5501000_5570000# GND efet w=1000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1508 diff_5699000_5570000# diff_475000_5142000# diff_5971000_5556000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=1.875e+09 ps=416000 
M1509 diff_94000_5193000# diff_5971000_5556000# diff_5971000_5556000# GND efet w=15000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M1510 diff_82000_3097000# diff_5618000_2171000# diff_6195000_5552000# GND efet w=130000 l=12000
+ ad=0 pd=0 as=-1.94997e+09 ps=540000 
M1511 diff_82000_3097000# diff_93000_3550000# diff_401000_4712000# GND efet w=79000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1512 diff_796000_5586000# diff_774000_5447000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1513 diff_1463000_5620000# diff_774000_5447000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1514 diff_1697000_5586000# diff_774000_5447000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1515 diff_2060000_5620000# diff_774000_5447000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1516 diff_2873000_5620000# diff_774000_5447000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1517 diff_3188000_5586000# diff_774000_5447000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1518 diff_3323000_5620000# diff_774000_5447000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1519 diff_3343000_5586000# diff_774000_5447000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1520 diff_3677000_5620000# diff_774000_5447000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1521 diff_3795000_5586000# diff_774000_5447000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1522 diff_3833000_5620000# diff_774000_5447000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1523 diff_4030000_5586000# diff_774000_5447000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1524 diff_4069000_5620000# diff_774000_5447000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1525 diff_4128000_5620000# diff_774000_5447000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1526 diff_4207000_5586000# diff_774000_5447000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1527 diff_4483000_5586000# diff_774000_5447000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1528 diff_6195000_5552000# diff_71000_4514000# diff_6015000_5534000# GND efet w=23000 l=14000
+ ad=0 pd=0 as=3.44e+08 ps=96000 
M1529 diff_82000_3097000# diff_6061000_5631000# diff_6195000_5552000# GND efet w=123500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1530 diff_82000_3097000# diff_6015000_5534000# diff_5971000_5556000# GND efet w=106000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1531 diff_90000_5336000# diff_87000_5399000# diff_82000_3097000# GND efet w=101000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1532 diff_90000_5336000# diff_196000_5469000# diff_82000_3097000# GND efet w=53500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M1533 diff_401000_4712000# diff_93000_3550000# diff_82000_3097000# GND efet w=71000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1534 diff_760000_5560000# diff_774000_5420000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1535 diff_893000_5620000# diff_774000_5420000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1536 diff_1011000_5620000# diff_774000_5420000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1537 diff_82000_3097000# diff_774000_5420000# diff_1129000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1538 diff_82000_3097000# diff_774000_5420000# diff_1463000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1539 diff_82000_3097000# diff_774000_5420000# diff_1677000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1540 diff_82000_3097000# diff_774000_5420000# diff_1697000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1541 diff_82000_3097000# diff_774000_5420000# diff_2060000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1542 diff_82000_3097000# diff_774000_5420000# diff_2560000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1543 diff_82000_3097000# diff_774000_5420000# diff_2776000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1544 diff_82000_3097000# diff_774000_5420000# diff_2834000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1545 diff_2873000_5620000# diff_774000_5420000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1546 diff_82000_3097000# diff_774000_5420000# diff_2893000_5586000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1547 diff_82000_3097000# diff_774000_5420000# diff_2932000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1548 diff_82000_3097000# diff_774000_5420000# diff_3011000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1549 diff_82000_3097000# diff_774000_5420000# diff_3050000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1550 diff_3070000_5586000# diff_774000_5420000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1551 diff_3129000_5586000# diff_774000_5420000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1552 diff_82000_3097000# diff_774000_5420000# diff_3323000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1553 diff_3559000_5620000# diff_774000_5420000# diff_82000_3097000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1554 diff_82000_3097000# diff_774000_5420000# diff_3579000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1555 diff_82000_3097000# diff_774000_5420000# diff_3638000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1556 diff_3677000_5620000# diff_774000_5420000# diff_82000_3097000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1557 diff_82000_3097000# diff_774000_5420000# diff_3697000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1558 diff_3833000_5620000# diff_774000_5420000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1559 diff_82000_3097000# diff_774000_5420000# diff_3892000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1560 diff_82000_3097000# diff_774000_5420000# diff_3951000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1561 diff_82000_3097000# diff_774000_5420000# diff_4010000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1562 diff_82000_3097000# diff_774000_5420000# diff_4030000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1563 diff_4069000_5620000# diff_774000_5420000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1564 diff_82000_3097000# diff_774000_5420000# diff_4128000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1565 diff_82000_3097000# diff_774000_5420000# diff_4581000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1566 diff_82000_3097000# diff_774000_5420000# diff_4846000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1567 diff_82000_3097000# diff_774000_5420000# diff_4866000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1568 diff_82000_3097000# diff_774000_5420000# diff_4905000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1569 diff_82000_3097000# diff_774000_5420000# diff_5081000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1570 diff_82000_3097000# diff_196000_5469000# diff_401000_4712000# GND efet w=132000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1571 diff_774000_5363000# diff_774000_5363000# diff_94000_5193000# GND efet w=16000 l=11000
+ ad=-1.84993e+09 pd=1.382e+06 as=0 ps=0 
M1572 diff_774000_5363000# diff_5251000_5061000# diff_82000_3097000# GND efet w=184000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1573 diff_774000_5363000# diff_5500000_5527000# diff_82000_3097000# GND efet w=191000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1574 diff_5500000_5527000# diff_5500000_5527000# diff_5500000_5527000# GND efet w=1000 l=2000
+ ad=-1.12597e+09 pd=710000 as=0 ps=0 
M1575 diff_82000_3097000# diff_5501000_5495000# diff_5500000_5527000# GND efet w=103000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1576 diff_82000_3097000# diff_5251000_5061000# diff_774000_5332000# GND efet w=181500 l=10500
+ ad=0 pd=0 as=2.11703e+09 ps=956000 
M1577 diff_774000_5332000# diff_5501000_5495000# diff_82000_3097000# GND efet w=181000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1578 diff_94000_5193000# diff_774000_5332000# diff_774000_5332000# GND efet w=15000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1579 diff_5500000_5527000# diff_5500000_5527000# diff_94000_5193000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M1580 diff_82000_3097000# diff_5699000_5495000# diff_5501000_5495000# GND efet w=103000 l=10000
+ ad=0 pd=0 as=-7.47967e+08 ps=626000 
M1581 diff_5500000_5527000# diff_5953000_5146000# diff_5699000_5495000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=6.3e+08 ps=144000 
M1582 diff_94000_5193000# diff_5501000_5495000# diff_5501000_5495000# GND efet w=15000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M1583 diff_82000_3097000# diff_6016000_5509000# diff_5971000_5481000# GND efet w=105000 l=11000
+ ad=0 pd=0 as=-2.10997e+09 ps=426000 
M1584 diff_5501000_5495000# diff_5501000_5495000# diff_5501000_5495000# GND efet w=1000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1585 diff_5699000_5495000# diff_475000_5142000# diff_5971000_5481000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M1586 diff_6195000_5552000# diff_6195000_5552000# diff_94000_5193000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M1587 diff_94000_5193000# diff_5971000_5481000# diff_5971000_5481000# GND efet w=14000 l=18000
+ ad=0 pd=0 as=0 ps=0 
M1588 diff_6195000_5480000# diff_71000_4514000# diff_6016000_5509000# GND efet w=21000 l=14000
+ ad=-1.94097e+09 pd=532000 as=3.01e+08 ps=92000 
M1589 diff_94000_5193000# diff_6195000_5480000# diff_6195000_5480000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M1590 diff_82000_3097000# diff_6061000_5631000# diff_6195000_5480000# GND efet w=124000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1591 diff_82000_3097000# diff_6039000_2950000# diff_6195000_5480000# GND efet w=132000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1592 diff_82000_3097000# diff_74000_5300000# diff_90000_5336000# GND efet w=225500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1593 diff_952000_5620000# diff_774000_5389000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1594 diff_1031000_5586000# diff_774000_5389000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1595 diff_1109000_5620000# diff_774000_5389000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1596 diff_1168000_5620000# diff_774000_5389000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1597 diff_1365000_5586000# diff_774000_5389000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1598 diff_1423000_5586000# diff_774000_5389000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1599 diff_1521000_5620000# diff_774000_5389000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1600 diff_1756000_5586000# diff_774000_5389000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1601 diff_2118000_5620000# diff_774000_5389000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1602 diff_2138000_5586000# diff_774000_5389000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1603 diff_2275000_5620000# diff_774000_5389000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1604 diff_2354000_5586000# diff_774000_5389000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1605 diff_2482000_5620000# diff_774000_5389000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1606 diff_2502000_5586000# diff_774000_5389000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1607 diff_2619000_5586000# diff_774000_5389000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1608 diff_2658000_5620000# diff_774000_5389000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1609 diff_3188000_5586000# diff_774000_5389000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1610 diff_3265000_5620000# diff_774000_5389000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1611 diff_3285000_5586000# diff_774000_5389000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1612 diff_3343000_5586000# diff_774000_5389000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1613 diff_3382000_5620000# diff_774000_5389000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1614 diff_3795000_5586000# diff_774000_5389000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1615 diff_3912000_5586000# diff_774000_5389000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1616 diff_4148000_5586000# diff_774000_5389000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1617 diff_4207000_5586000# diff_774000_5389000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1618 diff_4287000_5620000# diff_774000_5389000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1619 diff_4522000_5620000# diff_774000_5389000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1620 diff_4729000_5620000# diff_774000_5389000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1621 diff_4925000_5586000# diff_774000_5389000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1622 diff_401000_4712000# diff_472000_5334000# diff_82000_3097000# GND efet w=157500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1623 diff_90000_5336000# diff_196000_5469000# diff_82000_3097000# GND efet w=51500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1624 diff_90000_5336000# diff_74000_5300000# diff_82000_3097000# GND efet w=189000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1625 diff_90000_5336000# diff_196000_5469000# diff_82000_3097000# GND efet w=51500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1626 diff_82000_3097000# diff_774000_5363000# diff_760000_5560000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1627 diff_796000_5586000# diff_774000_5363000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1628 diff_82000_3097000# diff_774000_5363000# diff_893000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1629 diff_82000_3097000# diff_774000_5363000# diff_913000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1630 diff_1031000_5586000# diff_774000_5363000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1631 diff_82000_3097000# diff_774000_5363000# diff_1129000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1632 diff_1168000_5620000# diff_774000_5363000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1633 diff_82000_3097000# diff_774000_5363000# diff_1365000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1634 diff_1423000_5586000# diff_774000_5363000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1635 diff_82000_3097000# diff_774000_5363000# diff_1463000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1636 diff_82000_3097000# diff_774000_5363000# diff_1521000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1637 diff_82000_3097000# diff_774000_5363000# diff_1677000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1638 diff_82000_3097000# diff_774000_5363000# diff_1697000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1639 diff_82000_3097000# diff_774000_5363000# diff_2060000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1640 diff_2118000_5620000# diff_774000_5363000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1641 diff_82000_3097000# diff_774000_5363000# diff_2237000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1642 diff_82000_3097000# diff_774000_5363000# diff_2275000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1643 diff_82000_3097000# diff_774000_5363000# diff_2334000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1644 diff_82000_3097000# diff_774000_5363000# diff_2502000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1645 diff_82000_3097000# diff_774000_5363000# diff_2560000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1646 diff_82000_3097000# diff_774000_5363000# diff_2599000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1647 diff_82000_3097000# diff_774000_5363000# diff_2678000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1648 diff_82000_3097000# diff_774000_5363000# diff_2776000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1649 diff_82000_3097000# diff_774000_5363000# diff_2814000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1650 diff_2834000_5586000# diff_774000_5363000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1651 diff_2873000_5620000# diff_774000_5363000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1652 diff_82000_3097000# diff_774000_5363000# diff_2932000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1653 diff_2952000_5586000# diff_774000_5363000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1654 diff_82000_3097000# diff_774000_5363000# diff_3011000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1655 diff_82000_3097000# diff_774000_5363000# diff_3050000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1656 diff_3070000_5586000# diff_774000_5363000# diff_82000_3097000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1657 diff_82000_3097000# diff_774000_5363000# diff_3129000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1658 diff_82000_3097000# diff_774000_5363000# diff_3188000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1659 diff_82000_3097000# diff_774000_5363000# diff_3461000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1660 diff_3500000_5620000# diff_774000_5363000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1661 diff_82000_3097000# diff_774000_5363000# diff_3559000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1662 diff_82000_3097000# diff_774000_5363000# diff_3579000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1663 diff_82000_3097000# diff_774000_5363000# diff_3638000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1664 diff_82000_3097000# diff_774000_5363000# diff_3677000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1665 diff_82000_3097000# diff_774000_5363000# diff_3697000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1666 diff_82000_3097000# diff_774000_5363000# diff_3795000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1667 diff_82000_3097000# diff_774000_5363000# diff_3833000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1668 diff_3951000_5620000# diff_774000_5363000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1669 diff_82000_3097000# diff_774000_5363000# diff_4010000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1670 diff_82000_3097000# diff_774000_5363000# diff_4030000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1671 diff_82000_3097000# diff_774000_5363000# diff_4069000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1672 diff_82000_3097000# diff_774000_5363000# diff_4207000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1673 diff_82000_3097000# diff_774000_5363000# diff_4404000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1674 diff_82000_3097000# diff_774000_5363000# diff_4424000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1675 diff_82000_3097000# diff_774000_5363000# diff_4542000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1676 diff_82000_3097000# diff_774000_5363000# diff_4581000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1677 diff_82000_3097000# diff_774000_5363000# diff_4601000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1678 diff_82000_3097000# diff_774000_5363000# diff_4749000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1679 diff_82000_3097000# diff_774000_5363000# diff_4866000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1680 diff_4925000_5586000# diff_774000_5363000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1681 diff_5061000_5620000# diff_774000_5363000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1682 diff_774000_5305000# diff_774000_5305000# diff_94000_5193000# GND efet w=16000 l=11000
+ ad=-1.12093e+09 pd=1.468e+06 as=0 ps=0 
M1683 diff_774000_5305000# diff_5251000_5061000# diff_82000_3097000# GND efet w=184000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1684 diff_774000_5305000# diff_5500000_5452000# diff_82000_3097000# GND efet w=189500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1685 diff_5500000_5452000# diff_5500000_5452000# diff_5500000_5452000# GND efet w=1000 l=2000
+ ad=-9.99967e+08 pd=706000 as=0 ps=0 
M1686 diff_82000_3097000# diff_5501000_5420000# diff_5500000_5452000# GND efet w=103000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1687 diff_82000_3097000# diff_5251000_5061000# diff_774000_5274000# GND efet w=180000 l=10000
+ ad=0 pd=0 as=2.05903e+09 ps=950000 
M1688 diff_774000_5274000# diff_5501000_5420000# diff_82000_3097000# GND efet w=179500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1689 diff_82000_3097000# diff_492000_5342000# diff_498000_5333000# GND efet w=140000 l=10000
+ ad=0 pd=0 as=1.522e+09 ps=386000 
M1690 diff_94000_5193000# diff_774000_5274000# diff_774000_5274000# GND efet w=16000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1691 diff_5500000_5452000# diff_5500000_5452000# diff_94000_5193000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M1692 diff_82000_3097000# diff_5699000_5420000# diff_5501000_5420000# GND efet w=103000 l=11000
+ ad=0 pd=0 as=-8.51967e+08 ps=624000 
M1693 diff_5500000_5452000# diff_5953000_5146000# diff_5699000_5420000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=6.3e+08 ps=144000 
M1694 diff_94000_5193000# diff_5971000_5405000# diff_5971000_5405000# GND efet w=14000 l=18000
+ ad=0 pd=0 as=1.999e+09 ps=454000 
M1695 diff_94000_5193000# diff_5501000_5420000# diff_5501000_5420000# GND efet w=15000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M1696 diff_82000_3097000# diff_5999000_2952000# diff_6171000_5415000# GND efet w=132000 l=12000
+ ad=0 pd=0 as=-1.55097e+09 ps=580000 
M1697 diff_82000_3097000# diff_6016000_5421000# diff_5971000_5405000# GND efet w=106500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1698 diff_5501000_5420000# diff_5501000_5420000# diff_5501000_5420000# GND efet w=1000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1699 diff_5699000_5420000# diff_475000_5142000# diff_5971000_5405000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M1700 diff_6171000_5415000# diff_71000_4514000# diff_6016000_5421000# GND efet w=23000 l=14000
+ ad=0 pd=0 as=3.27e+08 ps=98000 
M1701 diff_82000_3097000# diff_6061000_5631000# diff_6171000_5415000# GND efet w=123500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M1702 diff_82000_3097000# diff_196000_5469000# diff_82000_3097000# GND efet w=8000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1703 diff_74000_5300000# diff_67000_5287000# diff_63000_4638000# GND efet w=30000 l=13000
+ ad=3.73e+08 pd=112000 as=7.10033e+08 ps=828000 
M1704 diff_472000_5334000# diff_67000_5287000# diff_464000_5279000# GND efet w=13000 l=13000
+ ad=2.04e+08 pd=96000 as=-1.55497e+09 ps=390000 
M1705 diff_498000_5333000# diff_501000_5321000# diff_464000_5279000# GND efet w=149500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1706 diff_464000_5279000# diff_464000_5279000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M1707 diff_94000_5193000# diff_84000_5212000# diff_94000_5159000# GND efet w=236500 l=9500
+ ad=0 pd=0 as=-7.26771e+08 ps=2.98e+06 
M1708 diff_501000_5321000# diff_71000_4514000# diff_99000_3991000# GND efet w=15000 l=13000
+ ad=2.54e+08 pd=102000 as=-3.49967e+08 ps=796000 
M1709 diff_952000_5620000# diff_774000_5332000# diff_82000_3097000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1710 diff_972000_5586000# diff_774000_5332000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1711 diff_1011000_5620000# diff_774000_5332000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1712 diff_1756000_5586000# diff_774000_5332000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1713 diff_2138000_5586000# diff_774000_5332000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1714 diff_2354000_5586000# diff_774000_5332000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1715 diff_2482000_5620000# diff_774000_5332000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1716 diff_2619000_5586000# diff_774000_5332000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1717 diff_2658000_5620000# diff_774000_5332000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1718 diff_2756000_5620000# diff_774000_5332000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1719 diff_2893000_5586000# diff_774000_5332000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1720 diff_3168000_5620000# diff_774000_5332000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1721 diff_3265000_5620000# diff_774000_5332000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1722 diff_3285000_5586000# diff_774000_5332000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1723 diff_3323000_5620000# diff_774000_5332000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1724 diff_3343000_5586000# diff_774000_5332000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1725 diff_3382000_5620000# diff_774000_5332000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1726 diff_3892000_5620000# diff_774000_5332000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1727 diff_4128000_5620000# diff_774000_5332000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1728 diff_4148000_5586000# diff_774000_5332000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1729 diff_4187000_5620000# diff_774000_5332000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1730 diff_4287000_5620000# diff_774000_5332000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1731 diff_4365000_5586000# diff_774000_5332000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1732 diff_4483000_5586000# diff_774000_5332000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1733 diff_4522000_5620000# diff_774000_5332000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1734 diff_4729000_5620000# diff_774000_5332000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1735 diff_4807000_5586000# diff_774000_5332000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1736 diff_4846000_5620000# diff_774000_5332000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1737 diff_4905000_5620000# diff_774000_5332000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1738 diff_82000_3097000# diff_774000_5305000# diff_796000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1739 diff_82000_3097000# diff_774000_5305000# diff_913000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1740 diff_82000_3097000# diff_774000_5305000# diff_952000_5620000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1741 diff_82000_3097000# diff_774000_5305000# diff_972000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1742 diff_82000_3097000# diff_774000_5305000# diff_1031000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1743 diff_82000_3097000# diff_774000_5305000# diff_1168000_5620000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1744 diff_82000_3097000# diff_774000_5305000# diff_1365000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1745 diff_82000_3097000# diff_774000_5305000# diff_1423000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1746 diff_82000_3097000# diff_774000_5305000# diff_1463000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1747 diff_82000_3097000# diff_774000_5305000# diff_1521000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1748 diff_82000_3097000# diff_774000_5305000# diff_1697000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1749 diff_82000_3097000# diff_774000_5305000# diff_1756000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1750 diff_82000_3097000# diff_774000_5305000# diff_2060000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1751 diff_82000_3097000# diff_774000_5305000# diff_2118000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1752 diff_82000_3097000# diff_774000_5305000# diff_2138000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1753 diff_82000_3097000# diff_774000_5305000# diff_2237000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1754 diff_82000_3097000# diff_774000_5305000# diff_2275000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1755 diff_82000_3097000# diff_774000_5305000# diff_2354000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1756 diff_82000_3097000# diff_774000_5305000# diff_2482000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1757 diff_82000_3097000# diff_774000_5305000# diff_2560000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1758 diff_82000_3097000# diff_774000_5305000# diff_2599000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1759 diff_82000_3097000# diff_774000_5305000# diff_2619000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1760 diff_82000_3097000# diff_774000_5305000# diff_2658000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1761 diff_82000_3097000# diff_774000_5305000# diff_2678000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1762 diff_82000_3097000# diff_774000_5305000# diff_2756000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1763 diff_82000_3097000# diff_774000_5305000# diff_2814000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1764 diff_82000_3097000# diff_774000_5305000# diff_2834000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1765 diff_82000_3097000# diff_774000_5305000# diff_2893000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1766 diff_82000_3097000# diff_774000_5305000# diff_2932000_5620000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1767 diff_82000_3097000# diff_774000_5305000# diff_2952000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1768 diff_82000_3097000# diff_774000_5305000# diff_3011000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1769 diff_82000_3097000# diff_774000_5305000# diff_3168000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1770 diff_82000_3097000# diff_774000_5305000# diff_3188000_5586000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1771 diff_82000_3097000# diff_774000_5305000# diff_3265000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1772 diff_82000_3097000# diff_774000_5305000# diff_3382000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1773 diff_82000_3097000# diff_774000_5305000# diff_3461000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1774 diff_82000_3097000# diff_774000_5305000# diff_3638000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1775 diff_82000_3097000# diff_774000_5305000# diff_3677000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1776 diff_82000_3097000# diff_774000_5305000# diff_3795000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1777 diff_82000_3097000# diff_774000_5305000# diff_4148000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1778 diff_82000_3097000# diff_774000_5305000# diff_4207000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1779 diff_82000_3097000# diff_774000_5305000# diff_4287000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1780 diff_82000_3097000# diff_774000_5305000# diff_4306000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1781 diff_82000_3097000# diff_774000_5305000# diff_4404000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1782 diff_82000_3097000# diff_774000_5305000# diff_4424000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1783 diff_82000_3097000# diff_774000_5305000# diff_4483000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1784 diff_82000_3097000# diff_774000_5305000# diff_4522000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1785 diff_82000_3097000# diff_774000_5305000# diff_4581000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1786 diff_82000_3097000# diff_774000_5305000# diff_4729000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1787 diff_82000_3097000# diff_774000_5305000# diff_4807000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1788 diff_82000_3097000# diff_774000_5305000# diff_4846000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1789 diff_82000_3097000# diff_774000_5305000# diff_4866000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1790 diff_82000_3097000# diff_774000_5305000# diff_4905000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1791 diff_82000_3097000# diff_774000_5305000# diff_4925000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1792 diff_82000_3097000# diff_774000_5305000# diff_5023000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1793 diff_774000_5248000# diff_774000_5248000# diff_94000_5193000# GND efet w=16000 l=10000
+ ad=-2.08693e+09 pd=1.336e+06 as=0 ps=0 
M1794 diff_774000_5248000# diff_5251000_5061000# diff_82000_3097000# GND efet w=182500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1795 diff_774000_5248000# diff_5500000_5376000# diff_82000_3097000# GND efet w=190500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1796 diff_5500000_5376000# diff_5500000_5376000# diff_5500000_5376000# GND efet w=500 l=1500
+ ad=-1.30697e+09 pd=664000 as=0 ps=0 
M1797 diff_82000_3097000# diff_5501000_5345000# diff_5500000_5376000# GND efet w=103000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1798 diff_82000_3097000# diff_5251000_5061000# diff_774000_5217000# GND efet w=180500 l=10500
+ ad=0 pd=0 as=1.93903e+09 ps=952000 
M1799 diff_774000_5217000# diff_5501000_5345000# diff_82000_3097000# GND efet w=181000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1800 diff_760000_5560000# diff_774000_5274000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1801 diff_834000_5620000# diff_774000_5274000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1802 diff_893000_5620000# diff_774000_5274000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1803 diff_1011000_5620000# diff_774000_5274000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1804 diff_1109000_5620000# diff_774000_5274000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1805 diff_1129000_5586000# diff_774000_5274000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1806 diff_2502000_5586000# diff_774000_5274000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1807 diff_2873000_5620000# diff_774000_5274000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1808 diff_3050000_5620000# diff_774000_5274000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1809 diff_3129000_5586000# diff_774000_5274000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1810 diff_3285000_5586000# diff_774000_5274000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1811 diff_3323000_5620000# diff_774000_5274000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1812 diff_3343000_5586000# diff_774000_5274000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1813 diff_3520000_5586000# diff_774000_5274000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1814 diff_3559000_5620000# diff_774000_5274000# diff_82000_3097000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1815 diff_3579000_5586000# diff_774000_5274000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1816 diff_3833000_5620000# diff_774000_5274000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1817 diff_3892000_5620000# diff_774000_5274000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1818 diff_3912000_5586000# diff_774000_5274000# diff_82000_3097000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1819 diff_3951000_5620000# diff_774000_5274000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1820 diff_4010000_5620000# diff_774000_5274000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1821 diff_4030000_5586000# diff_774000_5274000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1822 diff_4069000_5620000# diff_774000_5274000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1823 diff_4128000_5620000# diff_774000_5274000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1824 diff_4187000_5620000# diff_774000_5274000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1825 diff_4365000_5586000# diff_774000_5274000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1826 diff_4542000_5586000# diff_774000_5274000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1827 diff_4601000_5586000# diff_774000_5274000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1828 diff_4749000_5586000# diff_774000_5274000# diff_82000_3097000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1829 diff_94000_5193000# diff_774000_5217000# diff_774000_5217000# GND efet w=15000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1830 diff_5500000_5376000# diff_5500000_5376000# diff_94000_5193000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M1831 diff_82000_3097000# diff_5699000_5344000# diff_5501000_5345000# GND efet w=103000 l=11000
+ ad=0 pd=0 as=-8.52967e+08 ps=624000 
M1832 diff_5500000_5376000# diff_5953000_5146000# diff_5699000_5344000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=6.21e+08 ps=146000 
M1833 diff_6171000_5415000# diff_6171000_5415000# diff_94000_5193000# GND efet w=15000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M1834 diff_82000_3097000# diff_6011000_5359000# diff_5971000_5330000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=-2.04497e+09 ps=420000 
M1835 diff_94000_5193000# diff_5501000_5345000# diff_5501000_5345000# GND efet w=15000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M1836 diff_5501000_5345000# diff_5501000_5345000# diff_5501000_5345000# GND efet w=1000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1837 diff_5699000_5344000# diff_475000_5142000# diff_5971000_5330000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M1838 diff_94000_5193000# diff_5971000_5330000# diff_5971000_5330000# GND efet w=14000 l=18000
+ ad=0 pd=0 as=0 ps=0 
M1839 diff_6171000_5341000# diff_71000_4514000# diff_6011000_5359000# GND efet w=24000 l=14000
+ ad=-1.60697e+09 pd=588000 as=3.53e+08 ps=100000 
M1840 diff_94000_5193000# diff_6171000_5341000# diff_6171000_5341000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M1841 diff_82000_3097000# diff_6061000_5631000# diff_6171000_5341000# GND efet w=124000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1842 diff_82000_3097000# diff_5970000_2952000# diff_6171000_5341000# GND efet w=130000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1843 diff_492000_5342000# diff_71000_4514000# diff_513000_5203000# GND efet w=13500 l=14500
+ ad=3.86e+08 pd=112000 as=1.683e+09 ps=318000 
M1844 diff_82000_3097000# diff_774000_5248000# diff_1187000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1845 diff_82000_3097000# diff_774000_5248000# diff_1247000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1846 diff_82000_3097000# diff_774000_5248000# diff_1285000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1847 diff_82000_3097000# diff_774000_5248000# diff_1305000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1848 diff_82000_3097000# diff_774000_5248000# diff_1345000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1849 diff_82000_3097000# diff_774000_5248000# diff_1794000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1850 diff_82000_3097000# diff_774000_5248000# diff_1943000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1851 diff_82000_3097000# diff_774000_5248000# diff_2334000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1852 diff_82000_3097000# diff_774000_5248000# diff_2393000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1853 diff_82000_3097000# diff_774000_5248000# diff_2502000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1854 diff_82000_3097000# diff_774000_5248000# diff_2619000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1855 diff_82000_3097000# diff_774000_5248000# diff_2893000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1856 diff_82000_3097000# diff_774000_5248000# diff_3050000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1857 diff_82000_3097000# diff_774000_5248000# diff_3441000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1858 diff_82000_3097000# diff_774000_5248000# diff_3559000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1859 diff_82000_3097000# diff_774000_5248000# diff_3618000_5620000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1860 diff_82000_3097000# diff_774000_5248000# diff_3833000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1861 diff_82000_3097000# diff_774000_5248000# diff_3853000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1862 diff_82000_3097000# diff_774000_5248000# diff_4069000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1863 diff_82000_3097000# diff_774000_5248000# diff_4148000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1864 diff_82000_3097000# diff_774000_5248000# diff_4846000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1865 diff_774000_5191000# diff_774000_5191000# diff_94000_5193000# GND efet w=16000 l=10000
+ ad=1.77203e+09 pd=1.23e+06 as=0 ps=0 
M1866 diff_774000_5191000# diff_5251000_5061000# diff_82000_3097000# GND efet w=182500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1867 diff_94000_5159000# diff_84000_5212000# diff_94000_5193000# GND efet w=243000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1868 diff_94000_5193000# diff_84000_5212000# diff_94000_5159000# GND efet w=243000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1869 diff_513000_5203000# diff_513000_5203000# diff_94000_5193000# GND efet w=15000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M1870 diff_82000_3097000# diff_196000_5469000# diff_513000_5203000# GND efet w=84000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1871 diff_82000_3097000# diff_76000_4826000# diff_94000_5159000# GND efet w=222000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1872 diff_94000_5159000# diff_76000_4826000# diff_82000_3097000# GND efet w=222000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1873 diff_82000_3097000# diff_76000_4826000# diff_94000_5159000# GND efet w=222000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1874 diff_94000_5159000# diff_76000_4826000# diff_82000_3097000# GND efet w=222000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1875 diff_82000_3097000# diff_76000_4826000# diff_94000_5159000# GND efet w=222000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1876 diff_94000_5159000# diff_76000_4826000# diff_82000_3097000# GND efet w=222000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1877 diff_82000_3097000# diff_76000_4826000# diff_84000_5212000# GND efet w=254500 l=10500
+ ad=0 pd=0 as=-5.40967e+08 ps=548000 
M1878 diff_94000_5193000# diff_84000_5212000# diff_94000_5159000# GND efet w=271500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1879 diff_475000_5142000# diff_464000_5068000# diff_82000_3097000# GND efet w=195000 l=10000
+ ad=4.07033e+08 pd=810000 as=0 ps=0 
M1880 diff_475000_5142000# diff_464000_5068000# diff_82000_3097000# GND efet w=164000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1881 diff_82000_3097000# diff_486000_5097000# diff_464000_5068000# GND efet w=132000 l=11000
+ ad=0 pd=0 as=-2.04897e+09 ps=360000 
M1882 diff_464000_5068000# diff_464000_5068000# diff_94000_5193000# GND efet w=14000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1883 diff_94000_5193000# diff_486000_5097000# diff_475000_5142000# GND efet w=147000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1884 diff_774000_5191000# diff_5500000_5301000# diff_82000_3097000# GND efet w=189500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1885 diff_5500000_5301000# diff_5500000_5301000# diff_5500000_5301000# GND efet w=500 l=1500
+ ad=-1.30597e+09 pd=666000 as=0 ps=0 
M1886 diff_82000_3097000# diff_5501000_5269000# diff_5500000_5301000# GND efet w=103000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1887 diff_82000_3097000# diff_5251000_5061000# diff_774000_5159000# GND efet w=180500 l=10500
+ ad=0 pd=0 as=1.83203e+09 ps=938000 
M1888 diff_774000_5159000# diff_5501000_5269000# diff_82000_3097000# GND efet w=180500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1889 diff_5500000_5301000# diff_5500000_5301000# diff_94000_5193000# GND efet w=14000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M1890 diff_94000_5193000# diff_774000_5159000# diff_774000_5159000# GND efet w=15000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1891 diff_952000_5620000# diff_774000_5217000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1892 diff_1168000_5620000# diff_774000_5217000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1893 diff_1403000_5620000# diff_774000_5217000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1894 diff_1483000_5586000# diff_774000_5217000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1895 diff_1521000_5620000# diff_774000_5217000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1896 diff_1638000_5586000# diff_774000_5217000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1897 diff_1756000_5586000# diff_774000_5217000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1898 diff_1814000_5586000# diff_774000_5217000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1899 diff_1963000_5586000# diff_774000_5217000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1900 diff_2021000_5586000# diff_774000_5217000# diff_82000_3097000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1901 diff_2080000_5586000# diff_774000_5217000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1902 diff_2138000_5586000# diff_774000_5217000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1903 diff_2275000_5620000# diff_774000_5217000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1904 diff_2295000_5586000# diff_774000_5217000# diff_82000_3097000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1905 diff_2354000_5586000# diff_774000_5217000# diff_82000_3097000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1906 diff_2413000_5586000# diff_774000_5217000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1907 diff_2482000_5620000# diff_774000_5217000# diff_82000_3097000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1908 diff_2540000_5620000# diff_774000_5217000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1909 diff_2873000_5620000# diff_774000_5217000# diff_82000_3097000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1910 diff_3129000_5586000# diff_774000_5217000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1911 diff_3382000_5620000# diff_774000_5217000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1912 diff_3951000_5620000# diff_774000_5217000# diff_82000_3097000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1913 diff_3971000_5586000# diff_774000_5217000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1914 diff_4345000_5620000# diff_774000_5217000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1915 diff_4787000_5620000# diff_774000_5217000# diff_82000_3097000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1916 diff_4866000_5586000# diff_774000_5217000# diff_82000_3097000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1917 diff_4905000_5620000# diff_774000_5217000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1918 diff_4925000_5586000# diff_774000_5217000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1919 diff_82000_3097000# diff_5699000_5269000# diff_5501000_5269000# GND efet w=103000 l=11000
+ ad=0 pd=0 as=-9.49967e+08 ps=628000 
M1920 diff_5500000_5301000# diff_5953000_5146000# diff_5699000_5269000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=6.13e+08 ps=146000 
M1921 diff_5971000_5255000# diff_5971000_5255000# diff_94000_5193000# GND efet w=14000 l=17000
+ ad=1.951e+09 pd=440000 as=0 ps=0 
M1922 diff_94000_5193000# diff_5501000_5269000# diff_5501000_5269000# GND efet w=15000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M1923 diff_82000_3097000# diff_6011000_5271000# diff_5971000_5255000# GND efet w=105000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1924 diff_5501000_5269000# diff_5501000_5269000# diff_5501000_5269000# GND efet w=1000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1925 diff_5699000_5269000# diff_475000_5142000# diff_5971000_5255000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M1926 diff_6171000_5281000# diff_71000_4514000# diff_6011000_5271000# GND efet w=23000 l=13000
+ ad=-7.89967e+08 pd=656000 as=3.64e+08 ps=100000 
M1927 diff_82000_3097000# diff_774000_5191000# diff_1031000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1928 diff_82000_3097000# diff_774000_5191000# diff_1187000_5586000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1929 diff_82000_3097000# diff_774000_5191000# diff_1247000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1930 diff_82000_3097000# diff_774000_5191000# diff_1403000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1931 diff_82000_3097000# diff_774000_5191000# diff_1483000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1932 diff_82000_3097000# diff_774000_5191000# diff_1618000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1933 diff_82000_3097000# diff_774000_5191000# diff_1697000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1934 diff_82000_3097000# diff_774000_5191000# diff_1814000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1935 diff_82000_3097000# diff_774000_5191000# diff_1943000_5620000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1936 diff_82000_3097000# diff_774000_5191000# diff_2080000_5586000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1937 diff_82000_3097000# diff_774000_5191000# diff_2217000_5620000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1938 diff_82000_3097000# diff_774000_5191000# diff_2295000_5586000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1939 diff_82000_3097000# diff_774000_5191000# diff_2334000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1940 diff_82000_3097000# diff_774000_5191000# diff_2393000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1941 diff_82000_3097000# diff_774000_5191000# diff_2413000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1942 diff_82000_3097000# diff_774000_5191000# diff_2502000_5586000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1943 diff_82000_3097000# diff_774000_5191000# diff_2540000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1944 diff_82000_3097000# diff_774000_5191000# diff_2619000_5586000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1945 diff_82000_3097000# diff_774000_5191000# diff_2893000_5586000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1946 diff_82000_3097000# diff_774000_5191000# diff_2991000_5620000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1947 diff_82000_3097000# diff_774000_5191000# diff_3050000_5620000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1948 diff_82000_3097000# diff_774000_5191000# diff_3559000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1949 diff_82000_3097000# diff_774000_5191000# diff_4069000_5620000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1950 diff_774000_5133000# diff_774000_5133000# diff_94000_5193000# GND efet w=16000 l=10000
+ ad=-2.01393e+09 pd=1.286e+06 as=0 ps=0 
M1951 diff_82000_3097000# diff_5251000_5061000# diff_774000_5133000# GND efet w=182000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1952 diff_774000_5133000# diff_5500000_5226000# diff_82000_3097000# GND efet w=188500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M1953 diff_82000_3097000# diff_5501000_5194000# diff_5500000_5226000# GND efet w=103000 l=10000
+ ad=0 pd=0 as=-1.30497e+09 ps=664000 
M1954 diff_5500000_5226000# diff_5500000_5226000# diff_5500000_5226000# GND efet w=500 l=1500
+ ad=0 pd=0 as=0 ps=0 
M1955 diff_952000_5620000# diff_774000_5159000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1956 diff_1285000_5620000# diff_774000_5159000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1957 diff_1305000_5586000# diff_774000_5159000# diff_82000_3097000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1958 diff_1521000_5620000# diff_774000_5159000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1959 diff_1736000_5620000# diff_774000_5159000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1960 diff_1756000_5586000# diff_774000_5159000# diff_82000_3097000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1961 diff_1794000_5620000# diff_774000_5159000# diff_82000_3097000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1962 diff_1963000_5586000# diff_774000_5159000# diff_82000_3097000# GND efet w=24000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1963 diff_2001000_5620000# diff_774000_5159000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1964 diff_2021000_5586000# diff_774000_5159000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1965 diff_2138000_5586000# diff_774000_5159000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1966 diff_2275000_5620000# diff_774000_5159000# diff_82000_3097000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1967 diff_2354000_5586000# diff_774000_5159000# diff_82000_3097000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1968 diff_2482000_5620000# diff_774000_5159000# diff_82000_3097000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1969 diff_2873000_5620000# diff_774000_5159000# diff_82000_3097000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1970 diff_3129000_5586000# diff_774000_5159000# diff_82000_3097000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1971 diff_3382000_5620000# diff_774000_5159000# diff_82000_3097000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1972 diff_3441000_5620000# diff_774000_5159000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1973 diff_3618000_5620000# diff_774000_5159000# diff_82000_3097000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1974 diff_3833000_5620000# diff_774000_5159000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1975 diff_3853000_5586000# diff_774000_5159000# diff_82000_3097000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1976 diff_3951000_5620000# diff_774000_5159000# diff_82000_3097000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1977 diff_3971000_5586000# diff_774000_5159000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1978 diff_4030000_5586000# diff_774000_5159000# diff_82000_3097000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1979 diff_4148000_5586000# diff_774000_5159000# diff_82000_3097000# GND efet w=24000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1980 diff_4345000_5620000# diff_774000_5159000# diff_82000_3097000# GND efet w=24000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1981 diff_4463000_5620000# diff_774000_5159000# diff_82000_3097000# GND efet w=24000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1982 diff_4787000_5620000# diff_774000_5159000# diff_82000_3097000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1983 diff_4846000_5620000# diff_774000_5159000# diff_82000_3097000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1984 diff_4866000_5586000# diff_774000_5159000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1985 diff_4905000_5620000# diff_774000_5159000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1986 diff_4925000_5586000# diff_774000_5159000# diff_82000_3097000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1987 diff_82000_3097000# diff_5251000_5061000# diff_774000_5102000# GND efet w=180000 l=11000
+ ad=0 pd=0 as=1.78903e+09 ps=952000 
M1988 diff_774000_5102000# diff_5501000_5194000# diff_82000_3097000# GND efet w=181000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1989 diff_5500000_5226000# diff_5500000_5226000# diff_94000_5193000# GND efet w=14000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M1990 diff_94000_5193000# diff_774000_5102000# diff_774000_5102000# GND efet w=15000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1991 diff_5501000_5194000# diff_5699000_5194000# diff_82000_3097000# GND efet w=103000 l=11000
+ ad=-9.71967e+08 pd=630000 as=0 ps=0 
M1992 diff_5500000_5226000# diff_5953000_5146000# diff_5699000_5194000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=6.02e+08 ps=146000 
M1993 diff_94000_5193000# diff_6171000_5281000# diff_6171000_5281000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M1994 diff_82000_3097000# diff_5599000_574000# diff_6171000_5281000# GND efet w=129500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M1995 diff_82000_3097000# diff_6061000_5631000# diff_5971000_5180000# GND efet w=105000 l=10000
+ ad=0 pd=0 as=-1.93197e+09 ps=534000 
M1996 diff_82000_3097000# diff_6061000_5631000# diff_6171000_5281000# GND efet w=123000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1997 diff_94000_5193000# diff_5501000_5194000# diff_5501000_5194000# GND efet w=15000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M1998 diff_5501000_5194000# diff_5501000_5194000# diff_5501000_5194000# GND efet w=1000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1999 diff_5699000_5194000# diff_475000_5142000# diff_5971000_5180000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M2000 diff_82000_3097000# diff_6073000_5194000# diff_5971000_5180000# GND efet w=106000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2001 diff_5971000_5180000# diff_5971000_5180000# diff_94000_5193000# GND efet w=14000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M2002 diff_6227000_5190000# diff_71000_4514000# diff_6073000_5194000# GND efet w=21000 l=13000
+ ad=-1.50497e+09 pd=584000 as=3.22e+08 ps=94000 
M2003 diff_82000_3097000# diff_774000_5133000# diff_1031000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2004 diff_1463000_5620000# diff_774000_5133000# diff_82000_3097000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2005 diff_82000_3097000# diff_774000_5133000# diff_1618000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2006 diff_82000_3097000# diff_774000_5133000# diff_1697000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2007 diff_82000_3097000# diff_774000_5133000# diff_2060000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2008 diff_82000_3097000# diff_774000_5133000# diff_2217000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2009 diff_82000_3097000# diff_774000_5133000# diff_2678000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2010 diff_82000_3097000# diff_774000_5133000# diff_2991000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2011 diff_82000_3097000# diff_774000_5133000# diff_3500000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2012 diff_82000_3097000# diff_774000_5133000# diff_3520000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2013 diff_82000_3097000# diff_774000_5133000# diff_3579000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2014 diff_3638000_5586000# diff_774000_5133000# diff_82000_3097000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2015 diff_82000_3097000# diff_774000_5133000# diff_3677000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2016 diff_82000_3097000# diff_774000_5133000# diff_3775000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2017 diff_82000_3097000# diff_774000_5133000# diff_3853000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2018 diff_82000_3097000# diff_774000_5133000# diff_3971000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2019 diff_4287000_5620000# diff_774000_5133000# diff_82000_3097000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2020 diff_82000_3097000# diff_774000_5133000# diff_4522000_5620000# GND efet w=24000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2021 diff_82000_3097000# diff_774000_5133000# diff_4601000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2022 diff_4729000_5620000# diff_774000_5133000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2023 diff_82000_3097000# diff_774000_5133000# diff_4749000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2024 diff_774000_5075000# diff_774000_5075000# diff_94000_5193000# GND efet w=16000 l=10000
+ ad=2.12003e+09 pd=1.23e+06 as=0 ps=0 
M2025 diff_774000_5075000# diff_5251000_5061000# diff_82000_3097000# GND efet w=182500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2026 diff_774000_5075000# diff_5500000_5151000# diff_82000_3097000# GND efet w=189500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2027 diff_82000_3097000# diff_6073000_5170000# diff_5971000_5105000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=-1.67597e+09 ps=580000 
M2028 diff_82000_3097000# diff_5501000_5119000# diff_5500000_5151000# GND efet w=103000 l=10000
+ ad=0 pd=0 as=-1.29697e+09 ps=680000 
M2029 diff_5500000_5151000# diff_5500000_5151000# diff_5500000_5151000# GND efet w=500 l=1500
+ ad=0 pd=0 as=0 ps=0 
M2030 diff_952000_5620000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2031 diff_1247000_5586000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2032 diff_1403000_5620000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2033 diff_1756000_5586000# diff_774000_5102000# diff_82000_3097000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2034 diff_1814000_5586000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2035 diff_2080000_5586000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2036 diff_2138000_5586000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2037 diff_2295000_5586000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2038 diff_2334000_5620000# diff_774000_5102000# diff_82000_3097000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2039 diff_2354000_5586000# diff_774000_5102000# diff_82000_3097000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2040 diff_2482000_5620000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2041 diff_2502000_5586000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2042 diff_2619000_5586000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2043 diff_2834000_5586000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2044 diff_2873000_5620000# diff_774000_5102000# diff_82000_3097000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2045 diff_2893000_5586000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2046 diff_3050000_5620000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2047 diff_3109000_5620000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2048 diff_3129000_5586000# diff_774000_5102000# diff_82000_3097000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2049 diff_3382000_5620000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2050 diff_3402000_5586000# diff_774000_5102000# diff_82000_3097000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2051 diff_3441000_5620000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2052 diff_3559000_5620000# diff_774000_5102000# diff_82000_3097000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2053 diff_3833000_5620000# diff_774000_5102000# diff_82000_3097000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2054 diff_3951000_5620000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2055 diff_4010000_5620000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2056 diff_4030000_5586000# diff_774000_5102000# diff_82000_3097000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2057 diff_4069000_5620000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2058 diff_4148000_5586000# diff_774000_5102000# diff_82000_3097000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2059 diff_4345000_5620000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2060 diff_4787000_5620000# diff_774000_5102000# diff_82000_3097000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2061 diff_4846000_5620000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2062 diff_4866000_5586000# diff_774000_5102000# diff_82000_3097000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2063 diff_4905000_5620000# diff_774000_5102000# diff_82000_3097000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2064 diff_4925000_5586000# diff_774000_5102000# diff_82000_3097000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2065 diff_82000_3097000# diff_5251000_5061000# diff_777000_5045000# GND efet w=181000 l=11000
+ ad=0 pd=0 as=-2.12493e+09 ps=956000 
M2066 diff_777000_5045000# diff_5501000_5119000# diff_82000_3097000# GND efet w=180000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2067 diff_5500000_5151000# diff_5500000_5151000# diff_94000_5193000# GND efet w=14000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M2068 diff_82000_3097000# diff_774000_5075000# diff_760000_5560000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2069 diff_82000_3097000# diff_774000_5075000# diff_796000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2070 diff_82000_3097000# diff_774000_5075000# diff_1168000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2071 diff_82000_3097000# diff_774000_5075000# diff_1285000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2072 diff_82000_3097000# diff_774000_5075000# diff_1305000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2073 diff_82000_3097000# diff_774000_5075000# diff_1365000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2074 diff_82000_3097000# diff_774000_5075000# diff_1423000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2075 diff_82000_3097000# diff_774000_5075000# diff_1521000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2076 diff_82000_3097000# diff_774000_5075000# diff_1638000_5586000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2077 diff_82000_3097000# diff_774000_5075000# diff_1677000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2078 diff_82000_3097000# diff_774000_5075000# diff_1794000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2079 diff_82000_3097000# diff_774000_5075000# diff_1943000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2080 diff_82000_3097000# diff_774000_5075000# diff_1963000_5586000# GND efet w=24000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2081 diff_82000_3097000# diff_774000_5075000# diff_2021000_5586000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2082 diff_82000_3097000# diff_774000_5075000# diff_2118000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2083 diff_82000_3097000# diff_774000_5075000# diff_2237000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2084 diff_82000_3097000# diff_774000_5075000# diff_2275000_5620000# GND efet w=24000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2085 diff_82000_3097000# diff_774000_5075000# diff_2540000_5620000# GND efet w=24000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2086 diff_82000_3097000# diff_774000_5075000# diff_2814000_5620000# GND efet w=24000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2087 diff_82000_3097000# diff_774000_5075000# diff_2834000_5586000# GND efet w=24000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2088 diff_82000_3097000# diff_774000_5075000# diff_2952000_5586000# GND efet w=24000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2089 diff_82000_3097000# diff_774000_5075000# diff_3011000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2090 diff_82000_3097000# diff_774000_5075000# diff_3070000_5586000# GND efet w=24000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2091 diff_82000_3097000# diff_774000_5075000# diff_3323000_5620000# GND efet w=24000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2092 diff_82000_3097000# diff_774000_5075000# diff_3402000_5586000# GND efet w=24000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2093 diff_82000_3097000# diff_774000_5075000# diff_3461000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2094 diff_82000_3097000# diff_774000_5075000# diff_3579000_5586000# GND efet w=24000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2095 diff_82000_3097000# diff_774000_5075000# diff_3638000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2096 diff_82000_3097000# diff_774000_5075000# diff_3677000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2097 diff_82000_3097000# diff_774000_5075000# diff_3775000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2098 diff_82000_3097000# diff_774000_5075000# diff_3795000_5586000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2099 diff_82000_3097000# diff_774000_5075000# diff_4010000_5620000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2100 diff_82000_3097000# diff_774000_5075000# diff_4207000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2101 diff_82000_3097000# diff_774000_5075000# diff_4404000_5620000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2102 diff_82000_3097000# diff_774000_5075000# diff_4424000_5586000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2103 diff_82000_3097000# diff_774000_5075000# diff_4483000_5586000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2104 diff_82000_3097000# diff_774000_5075000# diff_4807000_5586000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2105 diff_486000_5097000# diff_486000_5097000# diff_94000_5193000# GND efet w=15000 l=16000
+ ad=1.811e+09 pd=380000 as=0 ps=0 
M2106 diff_377000_4962000# diff_67000_5287000# diff_94000_5193000# GND efet w=173500 l=11500
+ ad=1.40103e+09 pd=956000 as=0 ps=0 
M2107 diff_94000_5193000# diff_377000_4962000# diff_377000_4962000# GND efet w=13000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M2108 diff_486000_5097000# diff_377000_4962000# diff_82000_3097000# GND efet w=98500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2109 diff_82000_3097000# diff_445000_4909000# diff_377000_4962000# GND efet w=257500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2110 diff_475000_5142000# diff_486000_5097000# diff_94000_5193000# GND efet w=37000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2111 diff_94000_5193000# diff_777000_5045000# diff_777000_5045000# GND efet w=16000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2112 diff_5501000_5119000# diff_5699000_5119000# diff_82000_3097000# GND efet w=103000 l=11000
+ ad=-9.75967e+08 pd=628000 as=0 ps=0 
M2113 diff_5500000_5151000# diff_5953000_5146000# diff_5699000_5119000# GND efet w=15000 l=15000
+ ad=0 pd=0 as=5.86e+08 ps=144000 
M2114 diff_94000_5193000# diff_5971000_5105000# diff_5971000_5105000# GND efet w=13000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M2115 diff_6227000_5160000# diff_71000_4514000# diff_6073000_5170000# GND efet w=22000 l=13000
+ ad=-8.84967e+08 pd=628000 as=3.48e+08 ps=96000 
M2116 diff_6227000_5190000# diff_6227000_5190000# diff_94000_5193000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M2117 diff_82000_3097000# diff_6061000_5631000# diff_5971000_5105000# GND efet w=115500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2118 diff_94000_5193000# diff_5501000_5119000# diff_5501000_5119000# GND efet w=15000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M2119 diff_5501000_5119000# diff_5501000_5119000# diff_5501000_5119000# GND efet w=1000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2120 diff_5699000_5119000# diff_475000_5142000# diff_5971000_5105000# GND efet w=14000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M2121 diff_6061000_5631000# diff_71000_4514000# diff_666000_3268000# GND efet w=57000 l=14000
+ ad=5.1e+08 pd=164000 as=6.71033e+08 ps=1.026e+06 
M2122 diff_82000_3097000# diff_5595000_413000# diff_6227000_5190000# GND efet w=151000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2123 diff_94000_5193000# diff_6227000_5160000# diff_6227000_5160000# GND efet w=14000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M2124 diff_82000_3097000# diff_4953000_397000# diff_6227000_5160000# GND efet w=150500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M2125 diff_5251000_5061000# diff_5251000_5061000# diff_94000_5193000# GND efet w=19000 l=10000
+ ad=-1.42797e+09 pd=600000 as=0 ps=0 
M2126 diff_82000_3097000# diff_377000_4962000# diff_5251000_5061000# GND efet w=210500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M2127 diff_854000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2128 diff_952000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2129 diff_1031000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2130 diff_1247000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2131 diff_1403000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2132 diff_1463000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2133 diff_1541000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2134 diff_1618000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2135 diff_1697000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2136 diff_1736000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2137 diff_1756000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2138 diff_1814000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2139 diff_2001000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2140 diff_2060000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2141 diff_2080000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2142 diff_2138000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2143 diff_2217000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2144 diff_2295000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2145 diff_2334000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2146 diff_2354000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2147 diff_2482000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2148 diff_2502000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2149 diff_2619000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2150 diff_2678000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2151 diff_2873000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2152 diff_2893000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2153 diff_2991000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2154 diff_3050000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2155 diff_3109000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2156 diff_3129000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2157 diff_3382000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2158 diff_3441000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2159 diff_3500000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2160 diff_3520000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2161 diff_3559000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2162 diff_3618000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2163 diff_3833000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2164 diff_3853000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2165 diff_3951000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2166 diff_3971000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2167 diff_4030000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2168 diff_4069000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2169 diff_4089000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2170 diff_4148000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2171 diff_4287000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2172 diff_4345000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2173 diff_4463000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2174 diff_4522000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2175 diff_4601000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2176 diff_4729000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2177 diff_4749000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2178 diff_4787000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2179 diff_4846000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2180 diff_4866000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2181 diff_4905000_5620000# diff_777000_5045000# diff_82000_3097000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2182 diff_4925000_5586000# diff_777000_5045000# diff_82000_3097000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2183 diff_82000_3097000# diff_505000_5536000# diff_952000_5620000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2184 diff_82000_3097000# diff_505000_5536000# diff_1187000_5586000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2185 diff_82000_3097000# diff_505000_5536000# diff_1247000_5586000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2186 diff_82000_3097000# diff_505000_5536000# diff_1285000_5620000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2187 diff_82000_3097000# diff_505000_5536000# diff_1305000_5586000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2188 diff_82000_3097000# diff_505000_5536000# diff_1483000_5586000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2189 diff_82000_3097000# diff_505000_5536000# diff_1521000_5620000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2190 diff_82000_3097000# diff_505000_5536000# diff_1736000_5620000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2191 diff_82000_3097000# diff_505000_5536000# diff_1794000_5620000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2192 diff_82000_3097000# diff_505000_5536000# diff_2001000_5620000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2193 diff_82000_3097000# diff_505000_5536000# diff_2021000_5586000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2194 diff_82000_3097000# diff_505000_5536000# diff_2334000_5620000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2195 diff_82000_3097000# diff_505000_5536000# diff_2354000_5586000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2196 diff_82000_3097000# diff_505000_5536000# diff_2413000_5586000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2197 diff_82000_3097000# diff_505000_5536000# diff_2482000_5620000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2198 diff_82000_3097000# diff_505000_5536000# diff_2502000_5586000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2199 diff_82000_3097000# diff_505000_5536000# diff_2873000_5620000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2200 diff_82000_3097000# diff_505000_5536000# diff_3050000_5620000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2201 diff_82000_3097000# diff_505000_5536000# diff_3129000_5586000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2202 diff_82000_3097000# diff_505000_5536000# diff_3559000_5620000# GND efet w=23000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2203 diff_82000_3097000# diff_505000_5536000# diff_4069000_5620000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2204 diff_82000_3097000# diff_505000_5536000# diff_4866000_5586000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2205 diff_377000_4962000# diff_67000_5287000# diff_94000_5193000# GND efet w=36000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2206 diff_377000_4962000# diff_445000_4909000# diff_82000_3097000# GND efet w=184000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2207 diff_84000_5212000# diff_84000_5212000# diff_94000_5193000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2208 diff_82000_3097000# diff_67000_5287000# diff_445000_4909000# GND efet w=174000 l=11000
+ ad=0 pd=0 as=1.38803e+09 ps=954000 
M2209 diff_760000_5560000# diff_377000_4962000# diff_699000_4693000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.35e+08 ps=96000 
M2210 diff_796000_5586000# diff_377000_4962000# diff_667000_4503000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2211 diff_834000_5620000# diff_377000_4962000# diff_763000_4720000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2212 diff_854000_5586000# diff_377000_4962000# diff_830000_4715000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.12e+08 ps=74000 
M2213 diff_893000_5620000# diff_377000_4962000# diff_860000_4715000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2214 diff_913000_5586000# diff_377000_4962000# diff_887000_4705000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.12e+08 ps=74000 
M2215 diff_952000_5620000# diff_377000_4962000# diff_885000_3952000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2216 diff_972000_5586000# diff_377000_4962000# diff_987000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2217 diff_1011000_5620000# diff_377000_4962000# diff_1017000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.24e+08 ps=94000 
M2218 diff_1031000_5586000# diff_377000_4962000# diff_983000_4376000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2219 diff_1109000_5620000# diff_377000_4962000# diff_1037000_4589000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.13e+08 ps=76000 
M2220 diff_1129000_5586000# diff_377000_4962000# diff_1145000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.32e+08 ps=94000 
M2221 diff_1168000_5620000# diff_377000_4962000# diff_1144000_4573000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2222 diff_1187000_5586000# diff_377000_4962000# diff_1203000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2223 diff_1227000_5620000# diff_377000_4962000# diff_1232000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.35e+08 ps=96000 
M2224 diff_1247000_5586000# diff_377000_4962000# diff_1262000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2225 diff_1285000_5620000# diff_377000_4962000# diff_1291000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.23e+08 ps=94000 
M2226 diff_1305000_5586000# diff_377000_4962000# diff_1321000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.32e+08 ps=92000 
M2227 diff_1345000_5620000# diff_377000_4962000# diff_1350000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.55e+08 ps=96000 
M2228 diff_1365000_5586000# diff_377000_4962000# diff_1380000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.55e+08 ps=94000 
M2229 diff_1403000_5620000# diff_377000_4962000# diff_1409000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.32e+08 ps=94000 
M2230 diff_1423000_5586000# diff_377000_4962000# diff_1439000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.32e+08 ps=94000 
M2231 diff_1463000_5620000# diff_377000_4962000# diff_1468000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2232 diff_1483000_5586000# diff_377000_4962000# diff_1498000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.55e+08 ps=96000 
M2233 diff_1521000_5620000# diff_377000_4962000# diff_1527000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2234 diff_1541000_5586000# diff_377000_4962000# diff_1556000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.55e+08 ps=96000 
M2235 diff_1618000_5620000# diff_377000_4962000# diff_1624000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2236 diff_1638000_5586000# diff_377000_4962000# diff_1654000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.32e+08 ps=94000 
M2237 diff_1677000_5620000# diff_377000_4962000# diff_1682000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2238 diff_1697000_5586000# diff_377000_4962000# diff_1712000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.12e+08 ps=94000 
M2239 diff_1736000_5620000# diff_377000_4962000# diff_1741000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2240 diff_1756000_5586000# diff_377000_4962000# diff_1771000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2241 diff_1794000_5620000# diff_377000_4962000# diff_1800000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2242 diff_1814000_5586000# diff_377000_4962000# diff_1830000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2243 diff_445000_4909000# diff_196000_5469000# diff_82000_3097000# GND efet w=175000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2244 diff_94000_5193000# diff_76000_4826000# diff_76000_4826000# GND efet w=36000 l=10000
+ ad=0 pd=0 as=1.30033e+08 ps=750000 
M2245 diff_82000_3097000# diff_77000_4694000# diff_76000_4826000# GND efet w=324500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2246 diff_445000_4909000# diff_410000_4782000# diff_82000_3097000# GND efet w=180000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2247 diff_82000_3097000# diff_87000_5399000# diff_77000_4694000# GND efet w=184000 l=10000
+ ad=0 pd=0 as=1.81003e+09 ps=1.066e+06 
M2248 diff_94000_5193000# diff_77000_4694000# diff_77000_4694000# GND efet w=14500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2249 diff_82000_3097000# diff_200000_4773000# diff_77000_4694000# GND efet w=180000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2250 diff_82000_3097000# diff_84000_4682000# diff_77000_4694000# GND efet w=180000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2251 diff_230000_4714000# diff_204000_4723000# diff_82000_3097000# GND efet w=77500 l=10500
+ ad=1.336e+09 pd=278000 as=0 ps=0 
M2252 diff_410000_4782000# diff_99000_3991000# diff_82000_3097000# GND efet w=70000 l=10000
+ ad=1.18e+09 pd=226000 as=0 ps=0 
M2253 diff_94000_5193000# diff_410000_4782000# diff_410000_4782000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2254 diff_94000_5193000# diff_445000_4909000# diff_445000_4909000# GND efet w=15500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M2255 diff_200000_4773000# diff_71000_4514000# diff_230000_4714000# GND efet w=19000 l=13000
+ ad=3.66e+08 pd=108000 as=0 ps=0 
M2256 diff_204000_4723000# diff_67000_5287000# diff_120000_4668000# GND efet w=15000 l=13000
+ ad=2.42e+08 pd=82000 as=1.896e+09 ps=330000 
M2257 diff_230000_4714000# diff_230000_4714000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2258 diff_82000_3097000# diff_84000_4682000# diff_120000_4668000# GND efet w=66000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2259 diff_94000_5193000# diff_120000_4668000# diff_120000_4668000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2260 diff_84000_4682000# diff_84000_4682000# diff_94000_5193000# GND efet w=15000 l=16000
+ ad=-7.26967e+08 pd=644000 as=0 ps=0 
M2261 diff_84000_4682000# diff_63000_4638000# diff_82000_3097000# GND efet w=107000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2262 diff_84000_4682000# diff_196000_5469000# diff_82000_3097000# GND efet w=108000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2263 diff_63000_4638000# diff_229000_4600000# diff_82000_3097000# GND efet w=109500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2264 diff_82000_3097000# diff_80000_4528000# diff_63000_4638000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2265 diff_94000_5193000# diff_63000_4638000# diff_63000_4638000# GND efet w=15000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M2266 diff_82000_3097000# diff_105000_4535000# diff_63000_4638000# GND efet w=116000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2267 diff_82000_3097000# diff_215000_4573000# diff_63000_4638000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2268 diff_154000_4529000# diff_168000_4544000# diff_82000_3097000# GND efet w=105500 l=10500
+ ad=1.734e+09 pd=310000 as=0 ps=0 
M2269 diff_154000_4529000# diff_71000_4514000# diff_105000_4535000# GND efet w=14000 l=13000
+ ad=0 pd=0 as=2.42e+08 ps=74000 
M2270 diff_80000_4528000# diff_71000_4514000# diff_73000_3121000# GND efet w=23000 l=14000
+ ad=3.86e+08 pd=112000 as=-1.93797e+09 ps=468000 
M2271 diff_154000_4529000# diff_154000_4529000# diff_94000_5193000# GND efet w=16000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M2272 diff_215000_4573000# diff_71000_4514000# diff_336000_4527000# GND efet w=15000 l=14000
+ ad=2.29e+08 pd=72000 as=-1.18297e+09 ps=634000 
M2273 diff_572000_4609000# diff_558000_4357000# diff_82000_3097000# GND efet w=199500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2274 diff_82000_3097000# diff_699000_4693000# diff_641000_4582000# GND efet w=44000 l=10000
+ ad=0 pd=0 as=1.598e+09 ps=320000 
M2275 diff_82000_3097000# diff_64000_4219000# diff_82000_4447000# GND efet w=67000 l=10000
+ ad=0 pd=0 as=-1.98797e+09 ps=432000 
M2276 diff_82000_3097000# diff_166000_4460000# diff_82000_4447000# GND efet w=66000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2277 diff_82000_4447000# diff_71000_4514000# diff_80000_4320000# GND efet w=20000 l=14000
+ ad=0 pd=0 as=1.081e+09 ps=284000 
M2278 diff_94000_5193000# diff_82000_4447000# diff_82000_4447000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2279 diff_82000_3097000# diff_80000_4320000# diff_108000_4358000# GND efet w=77000 l=10000
+ ad=0 pd=0 as=1.123e+09 ps=238000 
M2280 diff_80000_4320000# diff_80000_4320000# diff_80000_4320000# GND efet w=500 l=1500
+ ad=0 pd=0 as=0 ps=0 
M2281 diff_94000_5193000# diff_108000_4358000# diff_108000_4358000# GND efet w=13000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2282 diff_82000_3097000# diff_108000_4358000# diff_87000_4248000# GND efet w=66500 l=11500
+ ad=0 pd=0 as=1.294e+09 ps=284000 
M2283 diff_87000_4248000# diff_67000_5287000# diff_80000_4320000# GND efet w=20000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M2284 diff_94000_5193000# diff_87000_4248000# diff_87000_4248000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2285 diff_94000_5193000# diff_479000_4479000# diff_479000_4479000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=-1.13897e+09 ps=536000 
M2286 diff_82000_3097000# diff_530000_4621000# diff_521000_4361000# GND efet w=131000 l=9000
+ ad=0 pd=0 as=-1.42397e+09 ps=628000 
M2287 diff_572000_4609000# diff_572000_4609000# diff_94000_5193000# GND efet w=14000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2288 diff_97000_4259000# diff_87000_4248000# diff_77000_4234000# GND efet w=105500 l=10500
+ ad=1.895e+09 pd=478000 as=5.17033e+08 ps=784000 
M2289 diff_82000_3097000# diff_105000_4267000# diff_97000_4259000# GND efet w=208000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2290 diff_315000_4257000# diff_315000_4257000# diff_94000_5193000# GND efet w=14000 l=16000
+ ad=2.055e+09 pd=392000 as=0 ps=0 
M2291 diff_77000_4234000# diff_87000_4248000# diff_97000_4259000# GND efet w=123000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2292 diff_315000_4257000# diff_71000_4514000# diff_105000_4267000# GND efet w=27000 l=13000
+ ad=0 pd=0 as=4.13e+08 ps=122000 
M2293 diff_82000_3097000# diff_100000_4085000# diff_77000_4234000# GND efet w=133500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M2294 diff_94000_5193000# diff_77000_4234000# diff_77000_4234000# GND efet w=14000 l=18000
+ ad=0 pd=0 as=0 ps=0 
M2295 diff_166000_4460000# diff_166000_4460000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=-1.39597e+09 pd=538000 as=0 ps=0 
M2296 diff_82000_3097000# diff_353000_4246000# diff_315000_4257000# GND efet w=110000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2297 diff_521000_4361000# diff_511000_4351000# diff_479000_4479000# GND efet w=135500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2298 diff_82000_3097000# diff_529000_4371000# diff_521000_4361000# GND efet w=149000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2299 diff_641000_4582000# diff_641000_4582000# diff_94000_5193000# GND efet w=15000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M2300 diff_82000_3097000# diff_667000_4503000# diff_641000_4582000# GND efet w=45000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2301 diff_577000_4446000# diff_577000_4446000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=1.631e+09 pd=320000 as=0 ps=0 
M2302 diff_82000_3097000# diff_582000_4389000# diff_577000_4446000# GND efet w=69500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2303 diff_740000_4507000# diff_724000_4489000# diff_685000_4520000# GND efet w=216500 l=9500
+ ad=1.95503e+09 pd=1.084e+06 as=-9.13967e+08 ps=688000 
M2304 diff_781000_4736000# diff_781000_4736000# diff_94000_5193000# GND efet w=13000 l=38000
+ ad=1.123e+09 pd=260000 as=0 ps=0 
M2305 diff_82000_3097000# diff_830000_4715000# diff_781000_4736000# GND efet w=45000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2306 diff_860000_4691000# diff_860000_4715000# diff_82000_3097000# GND efet w=45000 l=10000
+ ad=1.393e+09 pd=278000 as=0 ps=0 
M2307 diff_1015000_4729000# diff_987000_4961000# diff_82000_3097000# GND efet w=141500 l=10500
+ ad=2.21033e+08 pd=734000 as=0 ps=0 
M2308 diff_82000_3097000# diff_887000_4705000# diff_860000_4691000# GND efet w=43000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2309 diff_94000_5193000# diff_685000_4520000# diff_685000_4520000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2310 diff_653000_4323000# diff_71000_4514000# diff_624000_4564000# GND efet w=14000 l=13000
+ ad=4.99e+08 pd=146000 as=-1.97297e+09 ps=498000 
M2311 diff_860000_4691000# diff_860000_4691000# diff_94000_5193000# GND efet w=15000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M2312 diff_794000_4432000# diff_763000_4720000# diff_724000_4489000# GND efet w=134000 l=10000
+ ad=9.41e+08 pd=282000 as=1.30033e+08 ps=794000 
M2313 diff_82000_3097000# diff_529000_4371000# diff_794000_4432000# GND efet w=134000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2314 diff_837000_4492000# diff_781000_4736000# diff_82000_3097000# GND efet w=208500 l=9500
+ ad=1.554e+09 pd=432000 as=0 ps=0 
M2315 diff_854000_4511000# diff_790000_4021000# diff_837000_4492000# GND efet w=209500 l=10500
+ ad=1.548e+09 pd=432000 as=0 ps=0 
M2316 diff_724000_4489000# diff_860000_4691000# diff_854000_4511000# GND efet w=208500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2317 diff_1015000_4729000# diff_596000_3012000# diff_935000_4585000# GND efet w=131000 l=10000
+ ad=0 pd=0 as=2.014e+09 ps=480000 
M2318 diff_82000_3097000# diff_1017000_4961000# diff_1015000_4729000# GND efet w=132000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2319 diff_935000_4585000# diff_935000_4585000# diff_94000_5193000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2320 diff_94000_5193000# diff_724000_4489000# diff_724000_4489000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M2321 diff_582000_4389000# diff_71000_4514000# diff_479000_4479000# GND efet w=14000 l=13000
+ ad=2.96e+08 pd=102000 as=0 ps=0 
M2322 diff_82000_3097000# diff_577000_4446000# diff_558000_4357000# GND efet w=67000 l=10000
+ ad=0 pd=0 as=-2.08893e+09 ps=1.172e+06 
M2323 diff_558000_4357000# diff_653000_4323000# diff_82000_3097000# GND efet w=79000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2324 diff_166000_4460000# diff_300000_4193000# diff_82000_3097000# GND efet w=69000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2325 diff_223000_4164000# diff_67000_5287000# diff_100000_4085000# GND efet w=16000 l=12000
+ ad=3.62e+08 pd=112000 as=-1.00997e+09 ps=706000 
M2326 diff_82000_3097000# diff_223000_4164000# diff_166000_4460000# GND efet w=75000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2327 diff_82000_3097000# diff_127000_4096000# diff_100000_4085000# GND efet w=120500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2328 diff_353000_4246000# diff_67000_5287000# diff_127000_4096000# GND efet w=21000 l=14000
+ ad=3.71e+08 pd=82000 as=2.008e+09 ps=408000 
M2329 diff_82000_3097000# diff_679000_4313000# diff_558000_4357000# GND efet w=62000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2330 diff_94000_5193000# diff_100000_4085000# diff_100000_4085000# GND efet w=14500 l=17500
+ ad=0 pd=0 as=0 ps=0 
M2331 diff_100000_4085000# diff_77000_4234000# diff_82000_3097000# GND efet w=106000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2332 diff_281000_4043000# diff_281000_4043000# diff_94000_5193000# GND efet w=14000 l=17000
+ ad=2.089e+09 pd=384000 as=0 ps=0 
M2333 diff_281000_4043000# diff_168000_4544000# diff_82000_3097000# GND efet w=93000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2334 diff_281000_4043000# diff_168000_4544000# diff_82000_3097000# GND efet w=17000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2335 diff_82000_3097000# diff_281000_4043000# diff_129000_3948000# GND efet w=117000 l=10000
+ ad=0 pd=0 as=1.896e+09 ps=366000 
M2336 diff_82000_3097000# diff_99000_3991000# diff_105000_3784000# GND efet w=109500 l=9500
+ ad=0 pd=0 as=-2.02097e+09 ps=388000 
M2337 diff_94000_5193000# diff_105000_3784000# diff_105000_3784000# GND efet w=13000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M2338 diff_129000_3948000# diff_129000_3948000# diff_94000_5193000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M2339 diff_82000_3097000# diff_129000_3948000# diff_105000_3784000# GND efet w=118000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M2340 diff_129000_3948000# diff_229000_4600000# diff_82000_3097000# GND efet w=102000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2341 diff_100000_4085000# diff_67000_5287000# diff_131000_3834000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.66e+08 ps=100000 
M2342 diff_336000_4527000# diff_233000_3859000# diff_82000_3097000# GND efet w=112500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2343 diff_140000_3843000# diff_131000_3834000# diff_82000_3097000# GND efet w=160000 l=10000
+ ad=-1.94297e+09 pd=542000 as=0 ps=0 
M2344 diff_233000_3859000# diff_233000_3859000# diff_94000_5193000# GND efet w=13000 l=23000
+ ad=1.761e+09 pd=374000 as=0 ps=0 
M2345 diff_233000_3859000# diff_93000_3752000# diff_140000_3843000# GND efet w=171500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2346 diff_336000_4527000# diff_336000_4527000# diff_94000_5193000# GND efet w=14000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M2347 diff_140000_3843000# diff_73000_3121000# diff_82000_3097000# GND efet w=27000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2348 diff_140000_3843000# diff_73000_3121000# diff_82000_3097000# GND efet w=106000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2349 diff_726000_4203000# diff_641000_4582000# diff_82000_3097000# GND efet w=202500 l=9500
+ ad=2.80033e+08 pd=976000 as=0 ps=0 
M2350 diff_740000_4507000# diff_667000_4503000# diff_726000_4203000# GND efet w=200500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2351 diff_726000_4203000# diff_756000_4474000# diff_740000_4507000# GND efet w=203000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2352 diff_94000_5193000# diff_558000_4357000# diff_558000_4357000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2353 diff_82000_3097000# diff_636000_4099000# diff_558000_4357000# GND efet w=79500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2354 diff_558000_4357000# diff_658000_4116000# diff_82000_3097000# GND efet w=77000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2355 diff_82000_3097000# diff_690000_4134000# diff_558000_4357000# GND efet w=66000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2356 diff_82000_3097000# diff_772000_4077000# diff_726000_4203000# GND efet w=201500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2357 diff_1025000_4535000# diff_518000_3031000# diff_82000_3097000# GND efet w=159500 l=10500
+ ad=-1.26967e+08 pd=780000 as=0 ps=0 
M2358 diff_1075000_4556000# diff_1075000_4556000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=2.059e+09 pd=498000 as=0 ps=0 
M2359 diff_1159000_4672000# diff_518000_3031000# diff_1075000_4556000# GND efet w=132000 l=10000
+ ad=1.056e+09 pd=280000 as=0 ps=0 
M2360 diff_82000_3097000# diff_1145000_4961000# diff_1159000_4672000# GND efet w=132000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2361 diff_1176000_4477000# diff_1144000_4573000# diff_82000_3097000# GND efet w=44000 l=10000
+ ad=1.183e+09 pd=228000 as=0 ps=0 
M2362 diff_992000_4387000# diff_983000_4376000# diff_974000_4363000# GND efet w=147500 l=9500
+ ad=1.171e+09 pd=312000 as=-1.82997e+09 ps=564000 
M2363 diff_82000_3097000# diff_1000000_4393000# diff_992000_4387000# GND efet w=147500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2364 diff_1025000_4535000# diff_596000_3012000# diff_82000_3097000# GND efet w=164500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2365 diff_1052000_4266000# diff_1037000_4589000# diff_1025000_4535000# GND efet w=151500 l=10500
+ ad=-1.56697e+09 pd=570000 as=0 ps=0 
M2366 diff_530000_4621000# diff_71000_4514000# diff_1125000_4458000# GND efet w=13000 l=12000
+ ad=-8.74935e+08 pd=1.132e+06 as=3.01e+08 ps=112000 
M2367 diff_82000_3097000# diff_105000_3784000# diff_93000_3752000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=-9.67967e+08 ps=624000 
M2368 diff_94000_5193000# diff_93000_3752000# diff_93000_3752000# GND efet w=15000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M2369 diff_82000_3097000# diff_91000_3713000# diff_93000_3752000# GND efet w=110000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2370 diff_93000_3752000# diff_196000_5469000# diff_82000_3097000# GND efet w=106500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2371 diff_82000_3097000# diff_117000_3657000# diff_91000_3713000# GND efet w=197000 l=10000
+ ad=0 pd=0 as=-2.11693e+09 ps=1.12e+06 
M2372 diff_91000_3713000# diff_93000_3550000# diff_82000_3097000# GND efet w=175500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2373 diff_186000_3711000# diff_67000_5287000# diff_117000_3657000# GND efet w=14000 l=13000
+ ad=1.225e+09 pd=250000 as=2.29e+08 ps=74000 
M2374 diff_94000_5193000# diff_186000_3711000# diff_186000_3711000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2375 diff_186000_3711000# diff_181000_3690000# diff_82000_3097000# GND efet w=74000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2376 diff_196000_5469000# diff_71000_4514000# diff_181000_3690000# GND efet w=15000 l=13000
+ ad=0 pd=0 as=2.42e+08 ps=90000 
M2377 diff_82000_3097000# diff_196000_5469000# diff_91000_3713000# GND efet w=65000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2378 diff_91000_3713000# diff_196000_5469000# diff_82000_3097000# GND efet w=103500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M2379 diff_91000_3713000# diff_91000_3713000# diff_94000_5193000# GND efet w=14000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2380 diff_651000_3858000# diff_607000_3764000# diff_82000_3097000# GND efet w=141500 l=10500
+ ad=1.016e+09 pd=298000 as=0 ps=0 
M2381 diff_634000_3799000# diff_659000_3852000# diff_651000_3858000# GND efet w=141500 l=10500
+ ad=1.36903e+09 pd=954000 as=0 ps=0 
M2382 diff_659000_3852000# diff_71000_4514000# diff_731000_3737000# GND efet w=16000 l=15000
+ ad=2.49e+08 pd=86000 as=-1.05697e+09 ps=564000 
M2383 diff_696000_3857000# diff_686000_3825000# diff_634000_3799000# GND efet w=132000 l=10000
+ ad=9.24e+08 pd=278000 as=0 ps=0 
M2384 diff_82000_3097000# diff_229000_4600000# diff_696000_3857000# GND efet w=132000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2385 diff_731000_3737000# diff_229000_4600000# diff_82000_3097000# GND efet w=99500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M2386 diff_82000_3097000# diff_751000_3796000# diff_731000_3737000# GND efet w=66000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2387 diff_634000_3799000# diff_634000_3799000# diff_94000_5193000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2388 diff_686000_3825000# diff_71000_4514000# diff_168000_4544000# GND efet w=14000 l=13000
+ ad=5.06e+08 pd=142000 as=-1.42097e+09 ps=596000 
M2389 diff_607000_3764000# diff_71000_4514000# diff_336000_4527000# GND efet w=13000 l=13000
+ ad=8.35e+08 pd=216000 as=0 ps=0 
M2390 diff_100000_3536000# diff_93000_3550000# diff_82000_3097000# GND efet w=123500 l=10500
+ ad=-4.78967e+08 pd=644000 as=0 ps=0 
M2391 diff_94000_5193000# diff_100000_3536000# diff_100000_3536000# GND efet w=15000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M2392 diff_810000_3855000# diff_569000_3596000# diff_791000_3824000# GND efet w=144500 l=9500
+ ad=1.173e+09 pd=304000 as=-7.27967e+08 ps=708000 
M2393 diff_82000_3097000# diff_659000_3852000# diff_810000_3855000# GND efet w=144000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2394 diff_974000_4363000# diff_974000_4363000# diff_94000_5193000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2395 diff_1052000_4266000# diff_1052000_4266000# diff_94000_5193000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2396 diff_1176000_4477000# diff_1176000_4477000# diff_94000_5193000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M2397 diff_1943000_5620000# diff_377000_4962000# diff_1948000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2398 diff_1963000_5586000# diff_377000_4962000# diff_1978000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.32e+08 ps=94000 
M2399 diff_2001000_5620000# diff_377000_4962000# diff_2006000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2400 diff_2021000_5586000# diff_377000_4962000# diff_2036000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2401 diff_2060000_5620000# diff_377000_4962000# diff_2066000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2402 diff_2080000_5586000# diff_377000_4962000# diff_2096000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.23e+08 ps=94000 
M2403 diff_2118000_5620000# diff_377000_4962000# diff_2124000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.32e+08 ps=94000 
M2404 diff_2138000_5586000# diff_377000_4962000# diff_2154000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.12e+08 ps=94000 
M2405 diff_2217000_5620000# diff_377000_4962000# diff_2222000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.35e+08 ps=96000 
M2406 diff_2237000_5586000# diff_377000_4962000# diff_2252000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2407 diff_2275000_5620000# diff_377000_4962000# diff_2281000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2408 diff_2295000_5586000# diff_377000_4962000# diff_2311000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2409 diff_2334000_5620000# diff_377000_4962000# diff_2340000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2410 diff_2354000_5586000# diff_377000_4962000# diff_2370000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2411 diff_2393000_5620000# diff_377000_4962000# diff_2398000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2412 diff_2413000_5586000# diff_377000_4962000# diff_2428000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2413 diff_2482000_5620000# diff_377000_4962000# diff_2487000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2414 diff_2502000_5586000# diff_377000_4962000# diff_2517000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2415 diff_2540000_5620000# diff_377000_4962000# diff_2546000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2416 diff_2560000_5586000# diff_377000_4962000# diff_2576000_4948000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.02e+08 ps=76000 
M2417 diff_2599000_5620000# diff_377000_4962000# diff_2605000_4946000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.12e+08 ps=74000 
M2418 diff_2619000_5586000# diff_377000_4962000# diff_2635000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2419 diff_2658000_5620000# diff_377000_4962000# diff_2663000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.36e+08 ps=98000 
M2420 diff_2678000_5586000# diff_377000_4962000# diff_2693000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2421 diff_2756000_5620000# diff_377000_4962000# diff_2761000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2422 diff_2776000_5586000# diff_377000_4962000# diff_2791000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.55e+08 ps=96000 
M2423 diff_2814000_5620000# diff_377000_4962000# diff_2820000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2424 diff_2834000_5586000# diff_377000_4962000# diff_2850000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=1.385e+09 ps=362000 
M2425 diff_2873000_5620000# diff_377000_4962000# diff_2879000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2426 diff_2893000_5586000# diff_377000_4962000# diff_2909000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.32e+08 ps=94000 
M2427 diff_2932000_5620000# diff_377000_4962000# diff_2848000_2985000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.35e+08 ps=96000 
M2428 diff_2952000_5586000# diff_377000_4962000# diff_2967000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2429 diff_2991000_5620000# diff_377000_4962000# diff_2997000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2430 diff_3011000_5586000# diff_377000_4962000# diff_3027000_4946000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.13e+08 ps=76000 
M2431 diff_3050000_5620000# diff_377000_4962000# diff_3055000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.35e+08 ps=96000 
M2432 diff_3070000_5586000# diff_377000_4962000# diff_3085000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2433 diff_3109000_5620000# diff_377000_4962000# diff_3115000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2434 diff_3129000_5586000# diff_377000_4962000# diff_3105000_3437000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=74000 
M2435 diff_3168000_5620000# diff_377000_4962000# diff_3173000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.55e+08 ps=96000 
M2436 diff_3188000_5586000# diff_377000_4962000# diff_3203000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.55e+08 ps=96000 
M2437 diff_3265000_5620000# diff_377000_4962000# diff_3270000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.55e+08 ps=96000 
M2438 diff_3285000_5586000# diff_377000_4962000# diff_3300000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2439 diff_3323000_5620000# diff_377000_4962000# diff_3329000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2440 diff_3343000_5586000# diff_377000_4962000# diff_3359000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.32e+08 ps=94000 
M2441 diff_3382000_5620000# diff_377000_4962000# diff_3388000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.32e+08 ps=94000 
M2442 diff_3402000_5586000# diff_377000_4962000# diff_3418000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.02e+08 ps=96000 
M2443 diff_3441000_5620000# diff_377000_4962000# diff_3446000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.37e+08 ps=98000 
M2444 diff_3461000_5586000# diff_377000_4962000# diff_3476000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2445 diff_3500000_5620000# diff_377000_4962000# diff_3506000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2446 diff_3520000_5586000# diff_377000_4962000# diff_3536000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.13e+08 ps=96000 
M2447 diff_3559000_5620000# diff_377000_4962000# diff_3564000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.35e+08 ps=98000 
M2448 diff_3579000_5586000# diff_377000_4962000# diff_3594000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.36e+08 ps=98000 
M2449 diff_3618000_5620000# diff_377000_4962000# diff_3624000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2450 diff_3638000_5586000# diff_377000_4962000# diff_3653000_3514000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2451 diff_3677000_5620000# diff_377000_4962000# diff_3682000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.55e+08 ps=96000 
M2452 diff_3697000_5586000# diff_377000_4962000# diff_3712000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.46e+08 ps=98000 
M2453 diff_3775000_5620000# diff_377000_4962000# diff_3780000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.35e+08 ps=96000 
M2454 diff_3795000_5586000# diff_377000_4962000# diff_3810000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2455 diff_3833000_5620000# diff_377000_4962000# diff_3839000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2456 diff_3853000_5586000# diff_377000_4962000# diff_3869000_4933000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.12e+08 ps=74000 
M2457 diff_3892000_5620000# diff_377000_4962000# diff_3898000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.12e+08 ps=96000 
M2458 diff_3912000_5586000# diff_377000_4962000# diff_3928000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2459 diff_3951000_5620000# diff_377000_4962000# diff_3956000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.25e+08 ps=98000 
M2460 diff_3971000_5586000# diff_377000_4962000# diff_3986000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.55e+08 ps=96000 
M2461 diff_4010000_5620000# diff_377000_4962000# diff_4016000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.12e+08 ps=96000 
M2462 diff_4030000_5586000# diff_377000_4962000# diff_4046000_4929000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.03e+08 ps=76000 
M2463 diff_4069000_5620000# diff_377000_4962000# diff_4074000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.35e+08 ps=96000 
M2464 diff_4089000_5586000# diff_377000_4962000# diff_4104000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.26e+08 ps=98000 
M2465 diff_4128000_5620000# diff_377000_4962000# diff_4134000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.32e+08 ps=94000 
M2466 diff_4148000_5586000# diff_377000_4962000# diff_4164000_4928000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.13e+08 ps=76000 
M2467 diff_4187000_5620000# diff_377000_4962000# diff_4192000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.36e+08 ps=98000 
M2468 diff_4207000_5586000# diff_377000_4962000# diff_4222000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.35e+08 ps=98000 
M2469 diff_4287000_5620000# diff_377000_4962000# diff_4292000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.12e+08 ps=96000 
M2470 diff_4306000_5586000# diff_377000_4962000# diff_4322000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.12e+08 ps=96000 
M2471 diff_4345000_5620000# diff_377000_4962000# diff_4350000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.35e+08 ps=96000 
M2472 diff_4365000_5586000# diff_377000_4962000# diff_4380000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2473 diff_4404000_5620000# diff_377000_4962000# diff_4410000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.23e+08 ps=96000 
M2474 diff_4424000_5586000# diff_377000_4962000# diff_4318000_4838000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.12e+08 ps=96000 
M2475 diff_4463000_5620000# diff_377000_4962000# diff_4468000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.24e+08 ps=98000 
M2476 diff_4483000_5586000# diff_377000_4962000# diff_4498000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.46e+08 ps=98000 
M2477 diff_4522000_5620000# diff_377000_4962000# diff_4528000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=8e+08 ps=310000 
M2478 diff_4542000_5586000# diff_377000_4962000# diff_4558000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2479 diff_4581000_5620000# diff_377000_4962000# diff_4586000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.35e+08 ps=98000 
M2480 diff_4601000_5586000# diff_377000_4962000# diff_4616000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.36e+08 ps=98000 
M2481 diff_4729000_5620000# diff_377000_4962000# diff_4734000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.35e+08 ps=96000 
M2482 diff_4749000_5586000# diff_377000_4962000# diff_4427000_3812000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.35e+08 ps=98000 
M2483 diff_4787000_5620000# diff_377000_4962000# diff_4769000_4457000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2484 diff_4807000_5586000# diff_377000_4962000# diff_4823000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M2485 diff_4846000_5620000# diff_377000_4962000# diff_4842000_4667000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.13e+08 ps=96000 
M2486 diff_4866000_5586000# diff_377000_4962000# diff_4882000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=4.71e+08 ps=164000 
M2487 diff_4905000_5620000# diff_377000_4962000# diff_4901000_4753000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=4.72e+08 ps=184000 
M2488 diff_4925000_5586000# diff_377000_4962000# diff_4919000_4771000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=1.452e+09 ps=378000 
M2489 diff_5003000_5620000# diff_377000_4962000# diff_5008000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.25e+08 ps=98000 
M2490 diff_5023000_5586000# diff_377000_4962000# diff_5038000_4961000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.36e+08 ps=98000 
M2491 diff_5061000_5620000# diff_377000_4962000# diff_5067000_4961000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.12e+08 ps=96000 
M2492 diff_5081000_5586000# diff_377000_4962000# diff_5097000_4893000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.12e+08 ps=74000 
M2493 diff_82000_3097000# diff_1232000_4961000# diff_93000_3157000# GND efet w=66000 l=10000
+ ad=0 pd=0 as=1.333e+09 ps=268000 
M2494 diff_806000_3039000# diff_1262000_4961000# diff_82000_3097000# GND efet w=66000 l=10000
+ ad=1.669e+09 pd=312000 as=0 ps=0 
M2495 diff_82000_3097000# diff_1291000_4961000# diff_990000_3075000# GND efet w=102000 l=9000
+ ad=0 pd=0 as=-1.71497e+09 ps=442000 
M2496 diff_93000_3157000# diff_93000_3157000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2497 diff_806000_3039000# diff_806000_3039000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2498 diff_1196000_3118000# diff_71000_4514000# diff_1199000_4479000# GND efet w=15000 l=14000
+ ad=-1.37967e+08 pd=822000 as=2.69e+08 ps=108000 
M2499 diff_1150000_4300000# diff_1125000_4458000# diff_82000_3097000# GND efet w=133000 l=10000
+ ad=1.541e+09 pd=320000 as=0 ps=0 
M2500 diff_1162000_4604000# diff_1144000_4573000# diff_1150000_4300000# GND efet w=132000 l=10000
+ ad=-5.01967e+08 pd=702000 as=0 ps=0 
M2501 diff_1196000_4347000# diff_1176000_4477000# diff_1162000_4604000# GND efet w=137000 l=10000
+ ad=1.105e+09 pd=292000 as=0 ps=0 
M2502 diff_82000_3097000# diff_1199000_4479000# diff_1196000_4347000# GND efet w=138000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2503 diff_1263000_4412000# diff_1252000_4406000# diff_1234000_4460000# GND efet w=133000 l=11000
+ ad=7.98e+08 pd=278000 as=-1.29397e+09 ps=590000 
M2504 diff_82000_3097000# diff_1203000_4961000# diff_1263000_4412000# GND efet w=133000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2505 diff_1447000_4597000# diff_1321000_4961000# diff_82000_3097000# GND efet w=66000 l=11000
+ ad=1.561e+09 pd=314000 as=0 ps=0 
M2506 diff_990000_3075000# diff_990000_3075000# diff_94000_5193000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M2507 diff_1234000_4460000# diff_1234000_4460000# diff_94000_5193000# GND efet w=15000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2508 diff_1447000_4597000# diff_1447000_4597000# diff_94000_5193000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2509 diff_94000_5193000# diff_1179000_3098000# diff_1179000_3098000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=1.377e+09 ps=366000 
M2510 diff_996000_3890000# diff_67000_5287000# diff_679000_4313000# GND efet w=15000 l=15000
+ ad=2.52e+08 pd=102000 as=-1.65497e+09 ps=576000 
M2511 diff_872000_3937000# diff_71000_4514000# diff_928000_3955000# GND efet w=16000 l=13000
+ ad=7.27033e+08 pd=860000 as=2.84e+08 ps=100000 
M2512 diff_791000_3824000# diff_67000_5287000# diff_751000_3796000# GND efet w=14000 l=13000
+ ad=0 pd=0 as=2.14e+08 ps=86000 
M2513 diff_731000_3737000# diff_731000_3737000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2514 diff_94000_5193000# diff_791000_3824000# diff_791000_3824000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2515 diff_82000_3097000# diff_123000_3548000# diff_100000_3536000# GND efet w=113000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2516 diff_82000_3097000# diff_607000_3764000# diff_569000_3596000# GND efet w=83000 l=10000
+ ad=0 pd=0 as=-6.98967e+08 ps=660000 
M2517 diff_82000_3097000# diff_93000_3550000# diff_634000_3799000# GND efet w=66000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2518 diff_94000_5193000# diff_229000_4600000# diff_229000_4600000# GND efet w=13000 l=24000
+ ad=0 pd=0 as=1.409e+09 ps=286000 
M2519 diff_100000_3536000# diff_87000_3356000# diff_82000_3097000# GND efet w=104000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2520 diff_100000_3536000# diff_71000_4514000# diff_103000_3495000# GND efet w=21000 l=15000
+ ad=0 pd=0 as=3.33e+08 ps=104000 
M2521 diff_123000_3548000# diff_71000_4514000# diff_103000_3449000# GND efet w=22000 l=15000
+ ad=2.96e+08 pd=108000 as=-1.23597e+09 ps=564000 
M2522 diff_103000_3449000# diff_103000_3495000# diff_82000_3097000# GND efet w=107500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2523 diff_82000_3097000# diff_110000_3413000# diff_103000_3449000# GND efet w=128500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2524 diff_94000_5193000# diff_103000_3449000# diff_103000_3449000# GND efet w=15000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M2525 diff_73000_3121000# diff_103000_3449000# diff_82000_3097000# GND efet w=117000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2526 diff_94000_5193000# diff_73000_3121000# diff_73000_3121000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M2527 diff_82000_3097000# diff_93000_3550000# diff_569000_3596000# GND efet w=81000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2528 diff_791000_3824000# diff_786000_3668000# diff_82000_3097000# GND efet w=71000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2529 diff_1162000_4604000# diff_1162000_4604000# diff_94000_5193000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2530 diff_82000_3097000# diff_885000_3952000# diff_872000_3937000# GND efet w=42000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2531 diff_679000_4313000# diff_928000_3955000# diff_82000_3097000# GND efet w=72000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2532 diff_935000_4585000# diff_71000_4514000# diff_1054000_3958000# GND efet w=16000 l=14000
+ ad=0 pd=0 as=2.83e+08 ps=102000 
M2533 diff_974000_4363000# diff_71000_4514000# diff_1078000_3957000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.52e+08 ps=102000 
M2534 diff_986000_3873000# diff_996000_3890000# diff_82000_3097000# GND efet w=67000 l=11000
+ ad=1.374e+09 pd=294000 as=0 ps=0 
M2535 diff_1030000_3948000# diff_71000_4514000# diff_986000_3873000# GND efet w=16000 l=13000
+ ad=4.25e+08 pd=124000 as=0 ps=0 
M2536 diff_1052000_4266000# diff_71000_4514000# diff_1133000_3806000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=3.25e+08 ps=100000 
M2537 diff_1075000_4556000# diff_71000_4514000# diff_1151000_3808000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.58e+08 ps=90000 
M2538 diff_872000_3937000# diff_872000_3937000# diff_94000_5193000# GND efet w=14000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M2539 diff_986000_3873000# diff_986000_3873000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2540 diff_679000_4313000# diff_679000_4313000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2541 diff_786000_3668000# diff_71000_4514000# diff_783000_3632000# GND efet w=14000 l=14000
+ ad=2.48e+08 pd=86000 as=7.30033e+08 ps=818000 
M2542 diff_791000_3824000# diff_67000_5287000# diff_730000_3543000# GND efet w=15000 l=15000
+ ad=0 pd=0 as=2.76e+08 ps=100000 
M2543 diff_82000_3097000# diff_93000_3157000# diff_229000_4600000# GND efet w=69000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2544 diff_1049000_3791000# diff_1030000_3948000# diff_690000_4134000# GND efet w=133000 l=10000
+ ad=1.064e+09 pd=282000 as=-1.96497e+09 ps=444000 
M2545 diff_82000_3097000# diff_1054000_3958000# diff_1049000_3791000# GND efet w=133000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2546 diff_636000_4099000# diff_1078000_3957000# diff_82000_3097000# GND efet w=66000 l=10000
+ ad=1.836e+09 pd=346000 as=0 ps=0 
M2547 diff_636000_4099000# diff_636000_4099000# diff_94000_5193000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2548 diff_1143000_3813000# diff_1133000_3806000# diff_658000_4116000# GND efet w=134000 l=10000
+ ad=1.072e+09 pd=284000 as=-1.24797e+09 ps=614000 
M2549 diff_82000_3097000# diff_1151000_3808000# diff_1143000_3813000# GND efet w=134000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2550 diff_658000_4116000# diff_658000_4116000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2551 diff_94000_5193000# diff_690000_4134000# diff_690000_4134000# GND efet w=13000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2552 diff_634000_3799000# diff_67000_5287000# diff_905000_3510000# GND efet w=22000 l=14000
+ ad=0 pd=0 as=3.22e+08 ps=114000 
M2553 diff_110000_3413000# diff_67000_5287000# diff_110000_3357000# GND efet w=23000 l=14000
+ ad=3.17e+08 pd=104000 as=-1.64967e+08 ps=646000 
M2554 diff_127000_3342000# diff_205000_3371000# diff_82000_3097000# GND efet w=86500 l=10500
+ ad=1.128e+09 pd=224000 as=0 ps=0 
M2555 diff_234000_3316000# diff_71000_4514000# diff_205000_3371000# GND efet w=16000 l=14000
+ ad=0 pd=0 as=2.59e+08 ps=88000 
M2556 diff_82000_3097000# diff_127000_3342000# diff_110000_3357000# GND efet w=112000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2557 diff_94000_5193000# diff_127000_3342000# diff_127000_3342000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2558 diff_94000_5193000# diff_110000_3357000# diff_110000_3357000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M2559 diff_110000_3357000# diff_87000_3356000# diff_82000_3097000# GND efet w=105000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2560 diff_110000_3357000# diff_234000_3316000# diff_82000_3097000# GND efet w=102000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2561 diff_82000_3097000# diff_730000_3543000# diff_168000_4544000# GND efet w=128000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2562 diff_94000_5193000# diff_64000_4219000# diff_64000_4219000# GND efet w=18000 l=10000
+ ad=0 pd=0 as=1.24303e+09 ps=1.084e+06 
M2563 diff_64000_4219000# diff_905000_3510000# diff_82000_3097000# GND efet w=257000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2564 diff_1580000_4324000# diff_859000_2986000# diff_82000_3097000# GND efet w=118000 l=10000
+ ad=-1.1989e+09 pd=1.93e+06 as=0 ps=0 
M2565 diff_82000_3097000# diff_1409000_4961000# diff_1540000_4609000# GND efet w=43000 l=12000
+ ad=0 pd=0 as=-1.55197e+09 ps=424000 
M2566 diff_1540000_4609000# diff_1439000_4961000# diff_82000_3097000# GND efet w=43000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2567 diff_82000_3097000# diff_1468000_4961000# diff_1540000_4609000# GND efet w=46000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2568 diff_82000_3097000# diff_1673000_4605000# diff_1580000_4324000# GND efet w=102000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2569 diff_1540000_4609000# diff_1540000_4609000# diff_94000_5193000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M2570 diff_82000_3097000# diff_1447000_4597000# diff_1179000_3098000# GND efet w=72000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2571 diff_168000_4544000# diff_168000_4544000# diff_94000_5193000# GND efet w=13000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M2572 diff_569000_3596000# diff_569000_3596000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2573 diff_87000_3356000# diff_67000_5287000# diff_89000_3264000# GND efet w=16000 l=14000
+ ad=2.71e+08 pd=92000 as=2.089e+09 ps=400000 
M2574 diff_89000_3264000# diff_110000_3253000# diff_82000_3097000# GND efet w=87000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2575 diff_94000_5193000# diff_89000_3264000# diff_89000_3264000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2576 diff_103000_3168000# diff_71000_4514000# diff_110000_3253000# GND efet w=14000 l=13000
+ ad=-1.08297e+09 pd=572000 as=2.88e+08 ps=94000 
M2577 diff_103000_3168000# diff_93000_3157000# diff_82000_3149000# GND efet w=215500 l=10500
+ ad=0 pd=0 as=2.007e+09 ps=490000 
M2578 diff_94000_5193000# diff_103000_3168000# diff_103000_3168000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2579 diff_82000_3149000# diff_64000_4219000# diff_82000_3132000# GND efet w=200000 l=10000
+ ad=0 pd=0 as=1.4e+09 ps=414000 
M2580 diff_82000_3132000# diff_73000_3121000# diff_82000_3097000# GND efet w=200000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2581 diff_82000_3097000# diff_533000_2988000# diff_518000_3031000# GND efet w=144000 l=10000
+ ad=0 pd=0 as=-1.32497e+09 ps=760000 
M2582 diff_518000_3031000# diff_518000_3031000# diff_94000_5193000# GND efet w=14000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M2583 diff_558000_2987000# diff_67000_5287000# diff_533000_2988000# GND efet w=15000 l=13000
+ ad=-1.63997e+09 pd=478000 as=5.72e+08 ps=154000 
M2584 diff_94000_5193000# diff_1594000_4501000# diff_1594000_4501000# GND efet w=15000 l=38000
+ ad=0 pd=0 as=1.332e+09 ps=254000 
M2585 diff_1550000_4376000# diff_1522000_4350000# diff_82000_3097000# GND efet w=105500 l=10500
+ ad=7.39e+08 pd=224000 as=0 ps=0 
M2586 diff_857000_3300000# diff_1380000_4961000# diff_1550000_4376000# GND efet w=105500 l=10500
+ ad=-1.37597e+09 pd=528000 as=0 ps=0 
M2587 diff_1594000_4501000# diff_1540000_4609000# diff_82000_3097000# GND efet w=62500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2588 diff_1741000_4512000# diff_1691000_4496000# diff_82000_3097000# GND efet w=201500 l=9500
+ ad=1.664e+09 pd=432000 as=0 ps=0 
M2589 diff_999000_2989000# diff_67000_5287000# diff_1691000_4496000# GND efet w=15000 l=12000
+ ad=-1.69793e+09 pd=1.38e+06 as=3.2e+08 ps=104000 
M2590 diff_82000_3097000# diff_639000_3021000# diff_558000_2987000# GND efet w=77000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2591 diff_666000_3268000# diff_668000_2929000# diff_82000_3097000# GND efet w=200000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2592 diff_82000_3097000# diff_686000_3100000# diff_666000_3268000# GND efet w=220500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2593 diff_1522000_4350000# diff_71000_4514000# diff_1476000_3931000# GND efet w=14000 l=14000
+ ad=3.92e+08 pd=110000 as=-1.84297e+09 ps=528000 
M2594 diff_1580000_4324000# diff_1580000_4324000# diff_94000_5193000# GND efet w=15000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M2595 diff_1405000_3518000# diff_71000_4514000# diff_530000_4621000# GND efet w=15000 l=13000
+ ad=1.359e+09 pd=348000 as=0 ps=0 
M2596 diff_1420000_3777000# diff_1350000_4961000# diff_82000_3097000# GND efet w=149000 l=10000
+ ad=1.151e+09 pd=314000 as=0 ps=0 
M2597 diff_1437000_3777000# diff_1405000_3518000# diff_1420000_3777000# GND efet w=150000 l=10000
+ ad=-2.04197e+09 pd=508000 as=0 ps=0 
M2598 diff_94000_5193000# diff_857000_3300000# diff_857000_3300000# GND efet w=13000 l=29000
+ ad=0 pd=0 as=0 ps=0 
M2599 diff_1580000_4324000# diff_1468000_4961000# diff_1741000_4512000# GND efet w=206000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2600 diff_1692000_4258000# diff_1594000_4501000# diff_82000_3097000# GND efet w=225500 l=10500
+ ad=2.046e+09 pd=466000 as=0 ps=0 
M2601 diff_1509000_3891000# diff_1236000_3460000# diff_1476000_3931000# GND efet w=103000 l=10000
+ ad=6.69e+08 pd=218000 as=0 ps=0 
M2602 diff_82000_3097000# diff_1515000_3899000# diff_1509000_3891000# GND efet w=102500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M2603 diff_1339000_3494000# diff_71000_4514000# diff_1234000_4460000# GND efet w=13000 l=13000
+ ad=4.73e+08 pd=138000 as=0 ps=0 
M2604 diff_686000_3100000# diff_99000_3991000# diff_82000_3097000# GND efet w=94500 l=10500
+ ad=-1.89497e+09 pd=432000 as=0 ps=0 
M2605 diff_999000_2989000# diff_67000_5287000# diff_1271000_3499000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.89e+08 ps=106000 
M2606 diff_1236000_3460000# diff_1271000_3499000# diff_82000_3097000# GND efet w=49000 l=10000
+ ad=1.274e+09 pd=256000 as=0 ps=0 
M2607 diff_857000_3300000# diff_67000_5287000# diff_822000_3288000# GND efet w=15000 l=13000
+ ad=0 pd=0 as=3.91e+08 ps=122000 
M2608 diff_1236000_3460000# diff_1236000_3460000# diff_94000_5193000# GND efet w=13000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M2609 diff_94000_5193000# diff_999000_2989000# diff_999000_2989000# GND efet w=13000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M2610 diff_999000_2989000# diff_1339000_3494000# diff_82000_3097000# GND efet w=147000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2611 diff_94000_5193000# diff_1437000_3777000# diff_1437000_3777000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2612 diff_596000_3012000# diff_93000_3550000# diff_82000_3097000# GND efet w=164000 l=10000
+ ad=8.47033e+08 pd=908000 as=0 ps=0 
M2613 diff_639000_3021000# diff_71000_4514000# diff_596000_3012000# GND efet w=14000 l=13000
+ ad=3.39e+08 pd=100000 as=0 ps=0 
M2614 diff_94000_5193000# diff_558000_2987000# diff_558000_2987000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2615 diff_82000_3097000# diff_93000_3157000# diff_742000_2973000# GND efet w=85000 l=10000
+ ad=0 pd=0 as=1.581e+09 ps=304000 
M2616 diff_686000_3100000# diff_686000_3100000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2617 diff_816000_3049000# diff_806000_3039000# diff_596000_3012000# GND efet w=338500 l=10500
+ ad=-1.70397e+09 pd=692000 as=0 ps=0 
M2618 diff_82000_3097000# diff_822000_3288000# diff_816000_3049000# GND efet w=338500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2619 diff_1476000_3931000# diff_1476000_3931000# diff_94000_5193000# GND efet w=15000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M2620 diff_1580000_4324000# diff_1482000_3489000# diff_1692000_4258000# GND efet w=218500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2621 diff_82000_3097000# diff_1275000_3286000# diff_624000_4564000# GND efet w=135500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M2622 diff_1965000_4583000# diff_1712000_4961000# diff_82000_3097000# GND efet w=44000 l=11000
+ ad=1.239e+09 pd=262000 as=0 ps=0 
M2623 diff_82000_3097000# diff_1741000_4961000# diff_2004000_4583000# GND efet w=69500 l=10500
+ ad=0 pd=0 as=1.064e+09 ps=260000 
M2624 diff_1673000_4605000# diff_2004000_4583000# diff_82000_3097000# GND efet w=70000 l=10000
+ ad=1.568e+09 pd=310000 as=0 ps=0 
M2625 diff_82000_3097000# diff_1771000_4961000# diff_1673000_4605000# GND efet w=67000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2626 diff_624000_4564000# diff_624000_4564000# diff_94000_5193000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M2627 diff_1965000_4583000# diff_1965000_4583000# diff_94000_5193000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M2628 diff_2004000_4583000# diff_2004000_4583000# diff_94000_5193000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2629 diff_82000_3097000# diff_685000_4520000# diff_1580000_4324000# GND efet w=99000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2630 diff_1515000_3899000# diff_1498000_4961000# diff_82000_3097000# GND efet w=69000 l=10000
+ ad=1.2e+09 pd=276000 as=0 ps=0 
M2631 diff_82000_3097000# diff_1527000_4961000# diff_1515000_3899000# GND efet w=78500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2632 diff_1515000_3899000# diff_1515000_3899000# diff_94000_5193000# GND efet w=13000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2633 diff_1162000_4604000# diff_67000_5287000# diff_1588000_4011000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.98e+08 ps=104000 
M2634 diff_1096000_3118000# diff_1588000_4011000# diff_82000_3097000# GND efet w=114000 l=10000
+ ad=2.093e+09 pd=490000 as=0 ps=0 
M2635 diff_82000_3097000# diff_93000_3550000# diff_1096000_3118000# GND efet w=116500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M2636 diff_1196000_3118000# diff_1515000_3899000# diff_82000_3097000# GND efet w=223000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2637 diff_1580000_4324000# diff_71000_4514000# diff_1740000_3999000# GND efet w=16000 l=12000
+ ad=0 pd=0 as=2.64e+08 ps=102000 
M2638 diff_1096000_3118000# diff_1096000_3118000# diff_94000_5193000# GND efet w=15000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M2639 diff_82000_3097000# diff_1712000_3884000# diff_1647000_3413000# GND efet w=112000 l=10000
+ ad=0 pd=0 as=4.93033e+08 ps=874000 
M2640 diff_1712000_3884000# diff_1740000_3999000# diff_82000_3097000# GND efet w=66000 l=11000
+ ad=1.547e+09 pd=336000 as=0 ps=0 
M2641 diff_82000_3097000# diff_93000_3550000# diff_1712000_3884000# GND efet w=84000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2642 diff_1437000_3777000# diff_67000_5287000# diff_1458000_3631000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.55e+08 ps=94000 
M2643 diff_94000_5193000# diff_945000_3262000# diff_945000_3262000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=-1.81697e+09 ps=568000 
M2644 diff_945000_3262000# diff_1458000_3631000# diff_82000_3097000# GND efet w=107500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M2645 diff_1196000_3118000# diff_1196000_3118000# diff_94000_5193000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2646 diff_82000_3097000# diff_93000_3550000# diff_1405000_3518000# GND efet w=70000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M2647 diff_94000_5193000# diff_1560000_3638000# diff_1560000_3638000# GND efet w=13000 l=37000
+ ad=0 pd=0 as=1.653e+09 ps=314000 
M2648 diff_1712000_3884000# diff_1712000_3884000# diff_94000_5193000# GND efet w=15000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M2649 diff_1096000_3118000# diff_71000_4514000# diff_1538000_3466000# GND efet w=14000 l=13000
+ ad=0 pd=0 as=1.045e+09 ps=254000 
M2650 diff_94000_5193000# diff_99000_3991000# diff_99000_3991000# GND efet w=17000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2651 diff_1647000_3413000# diff_91000_3713000# diff_82000_3097000# GND efet w=102000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2652 diff_94000_5193000# diff_1482000_3489000# diff_1482000_3489000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=1.533e+09 ps=274000 
M2653 diff_82000_3097000# diff_1538000_3466000# diff_1560000_3638000# GND efet w=48000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2654 diff_1560000_3638000# diff_67000_5287000# diff_1474000_3479000# GND efet w=14000 l=13000
+ ad=0 pd=0 as=3.15e+08 ps=104000 
M2655 diff_1482000_3489000# diff_1474000_3479000# diff_82000_3097000# GND efet w=71000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2656 diff_82000_3097000# diff_1621000_3413000# diff_99000_3991000# GND efet w=213500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2657 diff_1673000_4605000# diff_1673000_4605000# diff_94000_5193000# GND efet w=16000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2658 diff_999000_2989000# diff_67000_5287000# diff_2059000_4466000# GND efet w=15000 l=15000
+ ad=0 pd=0 as=2.35e+08 ps=96000 
M2659 diff_82000_3097000# diff_1800000_4961000# diff_2062000_4303000# GND efet w=65000 l=10000
+ ad=0 pd=0 as=-1.67997e+09 ps=562000 
M2660 diff_82000_3097000# diff_2186000_4494000# diff_790000_4021000# GND efet w=309000 l=10000
+ ad=0 pd=0 as=-2.94902e+08 ps=2.462e+06 
M2661 diff_82000_3097000# diff_2006000_4961000# diff_2186000_4494000# GND efet w=112000 l=11000
+ ad=0 pd=0 as=2.11303e+09 ps=1.122e+06 
M2662 diff_2186000_4494000# diff_2036000_4961000# diff_82000_3097000# GND efet w=115000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2663 diff_790000_4021000# diff_2066000_4961000# diff_82000_3097000# GND efet w=317000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2664 diff_82000_3097000# diff_2096000_4961000# diff_790000_4021000# GND efet w=317000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2665 diff_790000_4021000# diff_2124000_4961000# diff_82000_3097000# GND efet w=324500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2666 diff_82000_3097000# diff_93000_3550000# diff_790000_4021000# GND efet w=327000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2667 diff_2062000_4303000# diff_2059000_4466000# diff_82000_3097000# GND efet w=68000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2668 diff_82000_3097000# diff_1482000_3489000# diff_2062000_4303000# GND efet w=68000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2669 diff_2062000_4303000# diff_2062000_4303000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2670 diff_1903000_3916000# diff_1654000_4961000# diff_82000_3097000# GND efet w=133000 l=10000
+ ad=1.064e+09 pd=282000 as=0 ps=0 
M2671 diff_1275000_3286000# diff_530000_4621000# diff_1903000_3916000# GND efet w=133000 l=10000
+ ad=1.94907e+09 pd=1.798e+06 as=0 ps=0 
M2672 diff_2186000_4494000# diff_2193000_4239000# diff_82000_3097000# GND efet w=110000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2673 diff_2172000_3037000# diff_2134000_4720000# diff_82000_3097000# GND efet w=68500 l=10500
+ ad=1.72033e+08 pd=814000 as=0 ps=0 
M2674 diff_2172000_3037000# diff_2370000_4961000# diff_82000_3097000# GND efet w=66500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M2675 diff_790000_4021000# diff_790000_4021000# diff_94000_5193000# GND efet w=28000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2676 diff_82000_3097000# diff_2154000_4961000# diff_2404000_4386000# GND efet w=46500 l=10500
+ ad=0 pd=0 as=-1.98597e+09 ps=526000 
M2677 diff_2565000_3499000# diff_2487000_4961000# diff_82000_3097000# GND efet w=80000 l=10000
+ ad=-2.39967e+08 pd=754000 as=0 ps=0 
M2678 diff_82000_3097000# diff_2517000_4961000# diff_2565000_3499000# GND efet w=67000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2679 diff_2172000_3037000# diff_2340000_4961000# diff_82000_3097000# GND efet w=68500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2680 diff_2197000_2999000# diff_2281000_4961000# diff_82000_3097000# GND efet w=71000 l=11000
+ ad=1.182e+09 pd=272000 as=0 ps=0 
M2681 diff_2404000_4386000# diff_2222000_4961000# diff_82000_3097000# GND efet w=45000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2682 diff_82000_3097000# diff_2252000_4961000# diff_2404000_4386000# GND efet w=46500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2683 diff_82000_3097000# diff_2311000_4961000# diff_2197000_2999000# GND efet w=71000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2684 diff_2186000_4494000# diff_2186000_4494000# diff_94000_5193000# GND efet w=15000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M2685 diff_1977000_3920000# diff_1952000_3749000# diff_82000_3097000# GND efet w=198000 l=11000
+ ad=1.386e+09 pd=410000 as=0 ps=0 
M2686 diff_1994000_3920000# diff_1624000_4961000# diff_1977000_3920000# GND efet w=198000 l=10000
+ ad=1.386e+09 pd=410000 as=0 ps=0 
M2687 diff_1464000_3203000# diff_1965000_4583000# diff_1994000_3920000# GND efet w=198000 l=11000
+ ad=1.06503e+09 pd=1.012e+06 as=0 ps=0 
M2688 diff_1647000_3413000# diff_1647000_3413000# diff_94000_5193000# GND efet w=15000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M2689 diff_1275000_3286000# diff_1275000_3286000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2690 diff_94000_5193000# diff_511000_4351000# diff_511000_4351000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=2.057e+09 ps=454000 
M2691 diff_1945000_3755000# diff_1682000_4961000# diff_1275000_3286000# GND efet w=145500 l=10500
+ ad=1.022e+09 pd=306000 as=0 ps=0 
M2692 diff_82000_3097000# diff_1952000_3749000# diff_1945000_3755000# GND efet w=146000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2693 diff_2094000_3974000# diff_1482000_3489000# diff_82000_3097000# GND efet w=213000 l=10000
+ ad=1.632e+09 pd=440000 as=0 ps=0 
M2694 diff_2112000_3993000# diff_1830000_4961000# diff_2094000_3974000# GND efet w=212000 l=10000
+ ad=1.574e+09 pd=440000 as=0 ps=0 
M2695 diff_2130000_4010000# diff_2119000_4000000# diff_2112000_3993000# GND efet w=212500 l=10500
+ ad=2.07403e+09 pd=1.088e+06 as=0 ps=0 
M2696 diff_2193000_4239000# diff_67000_5287000# diff_2221000_4171000# GND efet w=22000 l=14000
+ ad=3.7e+08 pd=98000 as=-1.87297e+09 ps=452000 
M2697 diff_2155000_3996000# diff_530000_4621000# diff_2130000_4010000# GND efet w=149500 l=10500
+ ad=-2.70967e+08 pd=638000 as=0 ps=0 
M2698 diff_82000_3097000# diff_1948000_4961000# diff_2155000_3996000# GND efet w=133000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2699 diff_2155000_3996000# diff_1978000_4961000# diff_82000_3097000# GND efet w=148000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2700 diff_772000_4077000# diff_1000000_4393000# diff_82000_3097000# GND efet w=65000 l=10000
+ ad=1.501e+09 pd=338000 as=0 ps=0 
M2701 diff_2404000_4386000# diff_2404000_4386000# diff_94000_5193000# GND efet w=15000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M2702 diff_2197000_2999000# diff_2197000_2999000# diff_94000_5193000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2703 diff_2569000_4387000# diff_2398000_4961000# diff_2172000_3037000# GND efet w=133000 l=11000
+ ad=9.31e+08 pd=280000 as=0 ps=0 
M2704 diff_82000_3097000# diff_530000_4621000# diff_2569000_4387000# GND efet w=133000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2705 diff_772000_4077000# diff_772000_4077000# diff_94000_5193000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2706 diff_2062000_4303000# diff_71000_4514000# diff_2255000_3931000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.45e+08 ps=96000 
M2707 diff_790000_4021000# diff_71000_4514000# diff_2336000_4017000# GND efet w=16000 l=14000
+ ad=0 pd=0 as=3.64e+08 ps=112000 
M2708 diff_94000_5193000# diff_2172000_3037000# diff_2172000_3037000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2709 diff_82000_3097000# diff_2255000_3931000# diff_2221000_4171000# GND efet w=80000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2710 diff_82000_3097000# diff_2062000_4303000# diff_1952000_3749000# GND efet w=70000 l=10000
+ ad=0 pd=0 as=-1.77397e+09 ps=454000 
M2711 diff_2323000_3767000# diff_2336000_4017000# diff_82000_3097000# GND efet w=66500 l=10500
+ ad=1.916e+09 pd=408000 as=0 ps=0 
M2712 diff_2072000_3805000# diff_67000_5287000# diff_2049000_3806000# GND efet w=14000 l=13000
+ ad=5.23e+08 pd=144000 as=-1.34897e+09 ps=550000 
M2713 diff_1464000_3203000# diff_1464000_3203000# diff_94000_5193000# GND efet w=15000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M2714 diff_82000_3097000# diff_1556000_4961000# diff_511000_4351000# GND efet w=66000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2715 diff_82000_3097000# diff_93000_3550000# diff_1538000_3466000# GND efet w=28000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M2716 diff_945000_3262000# diff_71000_4514000# diff_945000_3224000# GND efet w=16000 l=14000
+ ad=0 pd=0 as=3.65e+08 ps=116000 
M2717 diff_905000_3225000# diff_71000_4514000# diff_916000_3185000# GND efet w=15000 l=14000
+ ad=-6.71967e+08 pd=734000 as=2.72e+08 ps=96000 
M2718 diff_1835000_3560000# diff_790000_4021000# diff_82000_3097000# GND efet w=132000 l=10000
+ ad=9.24e+08 pd=278000 as=0 ps=0 
M2719 diff_1275000_3286000# diff_1624000_4961000# diff_1835000_3560000# GND efet w=132000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2720 diff_1275000_3286000# diff_1096000_3118000# diff_82000_3097000# GND efet w=65000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2721 diff_82000_3097000# diff_1196000_3118000# diff_1275000_3286000# GND efet w=64000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2722 diff_82000_3097000# diff_874000_3124000# diff_859000_2986000# GND efet w=124500 l=11500
+ ad=0 pd=0 as=-9.06967e+08 ps=584000 
M2723 diff_94000_5193000# diff_666000_3268000# diff_666000_3268000# GND efet w=18000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2724 diff_742000_2973000# diff_742000_2973000# diff_94000_5193000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2725 diff_596000_3012000# diff_596000_3012000# diff_94000_5193000# GND efet w=15000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2726 diff_913000_3047000# diff_916000_3185000# diff_82000_3097000# GND efet w=87500 l=10500
+ ad=-1.70897e+09 pd=500000 as=0 ps=0 
M2727 diff_963000_3081000# diff_945000_3224000# diff_913000_3047000# GND efet w=133000 l=10000
+ ad=1.064e+09 pd=282000 as=0 ps=0 
M2728 diff_82000_3097000# diff_511000_4351000# diff_963000_3081000# GND efet w=133000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2729 diff_966000_2988000# diff_990000_3075000# diff_82000_3097000# GND efet w=95500 l=10500
+ ad=-1.11897e+09 pd=510000 as=0 ps=0 
M2730 diff_913000_3047000# diff_67000_5287000# diff_874000_3124000# GND efet w=15000 l=13000
+ ad=0 pd=0 as=3.02e+08 ps=82000 
M2731 diff_859000_2986000# diff_859000_2986000# diff_94000_5193000# GND efet w=15000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M2732 diff_94000_5193000# diff_668000_2929000# diff_668000_2929000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=1.703e+09 ps=320000 
M2733 diff_668000_2929000# diff_336000_4527000# diff_82000_3097000# GND efet w=129500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2734 diff_913000_3047000# diff_913000_3047000# diff_94000_5193000# GND efet w=15000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M2735 diff_82000_3097000# diff_1047000_3118000# diff_1027000_3007000# GND efet w=78000 l=11000
+ ad=0 pd=0 as=-1.55497e+09 ps=564000 
M2736 diff_82000_3097000# diff_1096000_3118000# diff_1047000_3118000# GND efet w=102000 l=10000
+ ad=0 pd=0 as=4.27065e+08 ps=1.514e+06 
M2737 diff_1047000_3118000# diff_64000_4219000# diff_82000_3097000# GND efet w=97000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2738 diff_82000_3097000# diff_1147000_3108000# diff_1047000_3118000# GND efet w=119500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M2739 diff_1027000_3007000# diff_1027000_3007000# diff_94000_5193000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M2740 diff_966000_2988000# diff_966000_2988000# diff_94000_5193000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2741 diff_82000_3097000# diff_966000_2988000# diff_1047000_3118000# GND efet w=102000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2742 diff_1189000_3106000# diff_1179000_3098000# diff_82000_3097000# GND efet w=67000 l=10000
+ ad=2.07033e+08 pd=748000 as=0 ps=0 
M2743 diff_82000_3097000# diff_1196000_3118000# diff_1189000_3106000# GND efet w=95000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2744 diff_1275000_3286000# diff_71000_4514000# diff_1275000_3248000# GND efet w=16000 l=14000
+ ad=0 pd=0 as=2.84e+08 ps=100000 
M2745 diff_1647000_3413000# diff_67000_5287000# diff_1621000_3413000# GND efet w=21000 l=13000
+ ad=0 pd=0 as=7.5e+08 ps=176000 
M2746 diff_82000_3097000# diff_168000_4544000# diff_1275000_3286000# GND efet w=67000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2747 diff_1978000_3618000# diff_1501000_2924000# diff_1555000_2818000# GND efet w=223000 l=10000
+ ad=1.653e+09 pd=492000 as=-1.08397e+09 ps=580000 
M2748 diff_82000_3097000# diff_1658000_2819000# diff_1978000_3618000# GND efet w=220000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2749 diff_2130000_4010000# diff_2130000_4010000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2750 diff_2221000_4171000# diff_2221000_4171000# diff_94000_5193000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2751 diff_2183000_3680000# diff_2173000_3676000# diff_2130000_4010000# GND efet w=132000 l=10000
+ ad=5.33033e+08 pd=790000 as=0 ps=0 
M2752 diff_2323000_3767000# diff_2323000_3767000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2753 diff_1952000_3749000# diff_1952000_3749000# diff_94000_5193000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M2754 diff_2173000_3676000# diff_2173000_3676000# diff_94000_5193000# GND efet w=14000 l=39000
+ ad=-2.01297e+09 pd=418000 as=0 ps=0 
M2755 diff_2648000_4396000# diff_2428000_4961000# diff_82000_3097000# GND efet w=133000 l=10000
+ ad=1.064e+09 pd=282000 as=0 ps=0 
M2756 diff_2565000_3499000# diff_1252000_4406000# diff_2648000_4396000# GND efet w=133000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2757 diff_2641000_3474000# diff_2635000_4961000# diff_82000_3097000# GND efet w=44000 l=11000
+ ad=1.102e+09 pd=224000 as=0 ps=0 
M2758 diff_2641000_3474000# diff_2641000_3474000# diff_94000_5193000# GND efet w=14000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M2759 diff_2688000_4367000# diff_2546000_4961000# diff_2565000_3499000# GND efet w=135500 l=10500
+ ad=9.34e+08 pd=284000 as=0 ps=0 
M2760 diff_82000_3097000# diff_530000_4621000# diff_2688000_4367000# GND efet w=134500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2761 diff_772000_4077000# diff_71000_4514000# diff_2470000_3861000# GND efet w=15000 l=15000
+ ad=0 pd=0 as=2.61e+08 ps=100000 
M2762 diff_2404000_4386000# diff_71000_4514000# diff_2489000_3878000# GND efet w=15000 l=15000
+ ad=0 pd=0 as=5.34e+08 ps=130000 
M2763 diff_2565000_3499000# diff_2565000_3499000# diff_94000_5193000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2764 diff_2049000_3806000# diff_2470000_3861000# diff_82000_3097000# GND efet w=68000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2765 diff_82000_3097000# diff_2489000_3878000# diff_2049000_3806000# GND efet w=80000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2766 diff_2134000_4720000# diff_2508000_3808000# diff_82000_3097000# GND efet w=76000 l=10000
+ ad=-2.03897e+09 pd=400000 as=0 ps=0 
M2767 diff_2916000_4681000# diff_2905000_4657000# diff_2877000_4621000# GND efet w=88000 l=11000
+ ad=5.28e+08 pd=188000 as=-1.80497e+09 ps=544000 
M2768 diff_82000_3097000# diff_2761000_4961000# diff_2916000_4681000# GND efet w=88000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2769 diff_2930000_4556000# diff_2791000_4961000# diff_82000_3097000# GND efet w=66000 l=9000
+ ad=-1.36397e+09 pd=556000 as=0 ps=0 
M2770 diff_82000_3097000# diff_2820000_4961000# diff_2930000_4556000# GND efet w=68500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2771 diff_2877000_4621000# diff_2877000_4621000# diff_94000_5193000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M2772 diff_94000_5193000# diff_2859000_4569000# diff_2859000_4569000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=1.436e+09 ps=326000 
M2773 diff_82000_3097000# diff_2970000_4655000# diff_2930000_4556000# GND efet w=70000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2774 diff_94000_5193000# diff_2930000_4556000# diff_2930000_4556000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2775 diff_3008000_4522000# diff_2879000_4961000# diff_82000_3097000# GND efet w=72500 l=10500
+ ad=-1.47597e+09 pd=606000 as=0 ps=0 
M2776 diff_3063000_4309000# diff_2909000_4961000# diff_3008000_4522000# GND efet w=136500 l=10500
+ ad=-8.08967e+08 pd=604000 as=0 ps=0 
M2777 diff_82000_3097000# diff_2876000_4436000# diff_2859000_4569000# GND efet w=87000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2778 diff_2876000_4436000# diff_71000_4514000# diff_2912000_4303000# GND efet w=14000 l=13000
+ ad=2.67e+08 pd=88000 as=-1.83597e+09 ps=472000 
M2779 diff_94000_5193000# diff_3008000_4522000# diff_3008000_4522000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2780 diff_2905000_4657000# diff_71000_4514000# diff_529000_4371000# GND efet w=15000 l=11000
+ ad=2.058e+09 pd=396000 as=8.91033e+08 ps=992000 
M2781 diff_2896000_4349000# diff_2693000_4961000# diff_82000_3097000# GND efet w=110500 l=10500
+ ad=8.69e+08 pd=236000 as=0 ps=0 
M2782 diff_2912000_4303000# diff_1000000_4393000# diff_2896000_4349000# GND efet w=89000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2783 diff_82000_3097000# diff_93000_3550000# diff_2905000_4657000# GND efet w=74000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M2784 diff_82000_3097000# diff_2569000_3911000# diff_2558000_3888000# GND efet w=148500 l=10500
+ ad=0 pd=0 as=-1.44693e+09 ps=1.318e+06 
M2785 diff_2558000_3888000# diff_945000_3262000# diff_82000_3097000# GND efet w=130500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M2786 diff_82000_3097000# diff_530000_4621000# diff_2558000_3888000# GND efet w=147500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2787 diff_2558000_3888000# diff_529000_4371000# diff_82000_3097000# GND efet w=141000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2788 diff_2912000_4303000# diff_2912000_4303000# diff_94000_5193000# GND efet w=13000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M2789 diff_82000_3097000# diff_2850000_4961000# diff_3011000_4153000# GND efet w=132000 l=11000
+ ad=0 pd=0 as=-8.75967e+08 ps=630000 
M2790 diff_3063000_4309000# diff_529000_4371000# diff_82000_3097000# GND efet w=131000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2791 diff_3228000_4781000# diff_3055000_4961000# diff_82000_3097000# GND efet w=68000 l=11000
+ ad=1.94603e+09 pd=1.206e+06 as=0 ps=0 
M2792 diff_3228000_4781000# diff_2134000_4720000# diff_82000_3097000# GND efet w=82000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2793 diff_3034000_4153000# diff_790000_4021000# diff_3011000_4153000# GND efet w=133000 l=11000
+ ad=-1.88297e+09 pd=454000 as=0 ps=0 
M2794 diff_1252000_4406000# diff_3115000_4961000# diff_82000_3097000# GND efet w=69500 l=10500
+ ad=1.911e+09 pd=370000 as=0 ps=0 
M2795 diff_1252000_4406000# diff_1252000_4406000# diff_94000_5193000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M2796 diff_82000_3097000# diff_2997000_4961000# diff_3183000_4335000# GND efet w=132000 l=10000
+ ad=0 pd=0 as=-6.67967e+08 ps=780000 
M2797 diff_3183000_4335000# diff_3027000_4946000# diff_82000_3097000# GND efet w=178500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2798 diff_3228000_4781000# diff_1000000_4393000# diff_3183000_4335000# GND efet w=154500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2799 diff_3358000_4500000# diff_3203000_4961000# diff_82000_3097000# GND efet w=84000 l=11000
+ ad=8.89065e+08 pd=1.796e+06 as=0 ps=0 
M2800 diff_82000_3097000# diff_3300000_4961000# diff_3358000_4500000# GND efet w=67000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2801 diff_3431000_4646000# diff_3420000_4637000# diff_3358000_4500000# GND efet w=147500 l=10500
+ ad=1.107e+09 pd=310000 as=0 ps=0 
M2802 diff_82000_3097000# diff_3329000_4961000# diff_3431000_4646000# GND efet w=149500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2803 diff_94000_5193000# diff_3358000_4500000# diff_3358000_4500000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2804 diff_3273000_4384000# diff_3085000_4961000# diff_3228000_4781000# GND efet w=151000 l=10000
+ ad=1.283e+09 pd=330000 as=0 ps=0 
M2805 diff_82000_3097000# diff_790000_4021000# diff_3273000_4384000# GND efet w=157000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2806 diff_3487000_4661000# diff_3487000_4661000# diff_94000_5193000# GND efet w=14000 l=38000
+ ad=1.529e+09 pd=376000 as=0 ps=0 
M2807 diff_3540000_4682000# diff_3388000_4961000# diff_3487000_4661000# GND efet w=89000 l=10000
+ ad=7.12e+08 pd=194000 as=0 ps=0 
M2808 diff_82000_3097000# diff_1000000_4393000# diff_3540000_4682000# GND efet w=89000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2809 diff_3701000_4747000# diff_2569000_3911000# diff_82000_3097000# GND efet w=44000 l=10000
+ ad=-1.80297e+09 pd=478000 as=0 ps=0 
M2810 diff_82000_3097000# diff_3564000_4961000# diff_3701000_4747000# GND efet w=44000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2811 diff_3755000_4643000# diff_3594000_4961000# diff_82000_3097000# GND efet w=87000 l=11000
+ ad=-1.94997e+09 pd=430000 as=0 ps=0 
M2812 diff_2798000_4039000# diff_2798000_4039000# diff_94000_5193000# GND efet w=14000 l=37000
+ ad=-9.99967e+08 pd=526000 as=0 ps=0 
M2813 diff_2798000_4039000# diff_2663000_4961000# diff_2852000_4057000# GND efet w=88000 l=11000
+ ad=0 pd=0 as=6.16e+08 ps=190000 
M2814 diff_2852000_4057000# diff_518000_3031000# diff_82000_3097000# GND efet w=88000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2815 diff_2798000_4039000# diff_71000_4514000# diff_2911000_3917000# GND efet w=16000 l=12000
+ ad=0 pd=0 as=5.8e+08 ps=148000 
M2816 diff_94000_5193000# diff_1000000_4393000# diff_1000000_4393000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=-1.07797e+09 ps=518000 
M2817 diff_2049000_3806000# diff_93000_3550000# diff_82000_3097000# GND efet w=66000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2818 diff_2134000_4720000# diff_2134000_4720000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2819 diff_2323000_3767000# diff_67000_5287000# diff_2339000_3696000# GND efet w=21000 l=12000
+ ad=0 pd=0 as=3.18e+08 ps=106000 
M2820 diff_2027000_3554000# diff_2027000_3554000# diff_94000_5193000# GND efet w=15000 l=23000
+ ad=1.648e+09 pd=274000 as=0 ps=0 
M2821 diff_756000_4474000# diff_756000_4474000# diff_94000_5193000# GND efet w=14000 l=16000
+ ad=1.825e+09 pd=342000 as=0 ps=0 
M2822 diff_1189000_3106000# diff_99000_3991000# diff_82000_3097000# GND efet w=68500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2823 diff_82000_3097000# diff_1250000_3050000# diff_1189000_3106000# GND efet w=81000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2824 diff_1280000_3070000# diff_1275000_3248000# diff_82000_3097000# GND efet w=44000 l=10000
+ ad=2.71033e+08 pd=736000 as=0 ps=0 
M2825 diff_1329000_3050000# diff_668000_2929000# diff_82000_3097000# GND efet w=247000 l=11000
+ ad=-1.17197e+09 pd=792000 as=0 ps=0 
M2826 diff_82000_3097000# diff_686000_3100000# diff_1329000_3050000# GND efet w=206500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2827 diff_1280000_3070000# diff_67000_5287000# diff_1410000_3065000# GND efet w=15000 l=13000
+ ad=0 pd=0 as=3.02e+08 ps=98000 
M2828 diff_1047000_3118000# diff_859000_2986000# diff_82000_3097000# GND efet w=115500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2829 diff_1189000_3106000# diff_1189000_3106000# diff_94000_5193000# GND efet w=16000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2830 diff_1280000_3070000# diff_1280000_3070000# diff_94000_5193000# GND efet w=16000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M2831 diff_1333000_2957000# diff_1339000_3007000# diff_1329000_3050000# GND efet w=239000 l=10000
+ ad=2.101e+09 pd=408000 as=0 ps=0 
M2832 diff_1147000_3108000# diff_67000_5287000# diff_999000_2989000# GND efet w=15000 l=13000
+ ad=2.45e+08 pd=86000 as=0 ps=0 
M2833 diff_1047000_3118000# diff_1047000_3118000# diff_94000_5193000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M2834 diff_1250000_3050000# diff_67000_5287000# diff_999000_2989000# GND efet w=14000 l=12000
+ ad=2.5e+08 pd=90000 as=0 ps=0 
M2835 diff_1481000_3102000# diff_71000_4514000# diff_1464000_3203000# GND efet w=15000 l=13000
+ ad=6.12e+08 pd=160000 as=0 ps=0 
M2836 diff_1339000_3007000# diff_1410000_3065000# diff_82000_3097000# GND efet w=120500 l=10500
+ ad=-7.54967e+08 pd=652000 as=0 ps=0 
M2837 diff_82000_3097000# diff_196000_5469000# diff_1339000_3007000# GND efet w=123500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2838 diff_1458000_2942000# diff_1481000_3102000# diff_82000_3097000# GND efet w=58000 l=10000
+ ad=-1.69497e+09 pd=486000 as=0 ps=0 
M2839 diff_133000_2383000# diff_122000_2594000# diff_94000_5193000# GND efet w=862000 l=11000
+ ad=-2.11974e+09 pd=4.28e+06 as=0 ps=0 
M2840 diff_82000_3097000# diff_552000_1210000# diff_122000_2594000# GND efet w=415500 l=10500
+ ad=0 pd=0 as=-1.5979e+09 ps=1.364e+06 
M2841 diff_94000_5193000# diff_122000_2594000# diff_133000_2383000# GND efet w=344000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2842 diff_82000_3097000# diff_122000_2373000# diff_122000_2594000# GND efet w=271000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2843 diff_94000_5193000# diff_122000_2594000# diff_133000_2383000# GND efet w=240500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M2844 diff_82000_3097000# diff_122000_2373000# diff_122000_2594000# GND efet w=183000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2845 diff_94000_5193000# diff_122000_2594000# diff_133000_2383000# GND efet w=240500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2846 diff_122000_2594000# diff_122000_2594000# diff_94000_5193000# GND efet w=43000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2847 diff_855000_2599000# diff_90000_5336000# diff_82000_3097000# GND efet w=306500 l=10500
+ ad=9.88033e+08 pd=634000 as=0 ps=0 
M2848 diff_133000_2383000# diff_122000_2373000# diff_82000_3097000# GND efet w=881000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2849 diff_82000_3097000# diff_122000_2373000# diff_133000_2383000# GND efet w=242000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2850 diff_94000_5193000# diff_122000_2373000# diff_122000_2373000# GND efet w=37000 l=10000
+ ad=0 pd=0 as=1.27607e+09 ps=1.28e+06 
M2851 diff_718000_2539000# diff_679000_1018000# diff_581000_2471000# GND efet w=36000 l=13000
+ ad=1.054e+09 pd=210000 as=5.75e+08 ps=112000 
M2852 diff_82000_3097000# diff_581000_2471000# diff_122000_2373000# GND efet w=414500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2853 diff_886000_2526000# diff_90000_5336000# diff_855000_2599000# GND efet w=297000 l=11000
+ ad=1.64503e+09 pd=634000 as=0 ps=0 
M2854 diff_916000_2526000# diff_90000_5336000# diff_886000_2526000# GND efet w=297000 l=10000
+ ad=-1.9179e+09 pd=1.194e+06 as=0 ps=0 
M2855 diff_947000_2557000# diff_937000_2547000# diff_916000_2526000# GND efet w=36000 l=10000
+ ad=1.77803e+09 pd=620000 as=0 ps=0 
M2856 diff_937000_2547000# diff_937000_2547000# diff_947000_2557000# GND efet w=28000 l=9000
+ ad=-1.28097e+09 pd=568000 as=0 ps=0 
M2857 diff_964000_2516000# diff_90000_5336000# diff_937000_2547000# GND efet w=262500 l=10500
+ ad=5.09065e+08 pd=842000 as=0 ps=0 
M2858 diff_947000_2557000# diff_937000_2547000# diff_916000_2526000# GND efet w=303000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2859 diff_1333000_2957000# diff_1333000_2957000# diff_94000_5193000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M2860 diff_82000_3097000# diff_1404000_2968000# diff_1339000_3007000# GND efet w=130500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M2861 diff_1658000_2819000# diff_2027000_3554000# diff_82000_3097000# GND efet w=101500 l=9500
+ ad=4.19033e+08 pd=854000 as=0 ps=0 
M2862 diff_1555000_2818000# diff_1555000_2818000# diff_94000_5193000# GND efet w=15000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M2863 diff_82000_3097000# diff_2072000_3805000# diff_756000_4474000# GND efet w=102000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2864 diff_82000_3097000# diff_2130000_4010000# diff_2027000_3554000# GND efet w=65000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2865 diff_2183000_3680000# diff_685000_4520000# diff_82000_3097000# GND efet w=134000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2866 diff_82000_3097000# diff_1673000_4605000# diff_2183000_3680000# GND efet w=134500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M2867 diff_82000_3097000# diff_1978000_4961000# diff_2173000_3676000# GND efet w=44000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2868 diff_1000000_4393000# diff_2339000_3696000# diff_82000_3097000# GND efet w=280500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M2869 diff_94000_5193000# diff_2049000_3806000# diff_2049000_3806000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2870 diff_2508000_3808000# diff_2576000_4948000# diff_2558000_3888000# GND efet w=151500 l=10500
+ ad=2.005e+09 pd=462000 as=0 ps=0 
M2871 diff_2558000_3888000# diff_783000_3632000# diff_82000_3097000# GND efet w=148000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2872 diff_2698000_3826000# diff_518000_3031000# diff_2508000_3808000# GND efet w=132500 l=11500
+ ad=8.49e+08 pd=278000 as=0 ps=0 
M2873 diff_82000_3097000# diff_2605000_4946000# diff_2698000_3826000# GND efet w=131500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2874 diff_94000_5193000# diff_2508000_3808000# diff_2508000_3808000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2875 diff_2269000_3389000# diff_742000_2973000# diff_82000_3097000# GND efet w=67000 l=9000
+ ad=-4.02967e+08 pd=590000 as=0 ps=0 
M2876 diff_905000_3225000# diff_93000_3550000# diff_82000_3097000# GND efet w=127500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2877 diff_82000_3097000# diff_2867000_3891000# diff_905000_3225000# GND efet w=134000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2878 diff_82000_3097000# diff_2911000_3917000# diff_2903000_3861000# GND efet w=82000 l=10000
+ ad=0 pd=0 as=1.591e+09 ps=328000 
M2879 diff_2910000_3803000# diff_2903000_3861000# diff_82000_3097000# GND efet w=68000 l=11000
+ ad=-1.49397e+09 pd=628000 as=0 ps=0 
M2880 diff_82000_3097000# diff_2964000_3935000# diff_2910000_3803000# GND efet w=65000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2881 diff_2964000_3935000# diff_71000_4514000# diff_3008000_3949000# GND efet w=15000 l=14000
+ ad=2.5e+08 pd=90000 as=7.83e+08 ps=188000 
M2882 diff_94000_5193000# diff_3034000_4153000# diff_3034000_4153000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2883 diff_2820000_3542000# diff_71000_4514000# diff_2937000_3466000# GND efet w=22000 l=13000
+ ad=-1.95497e+09 pd=518000 as=-2.00097e+09 ps=514000 
M2884 diff_3008000_3949000# diff_3008000_3949000# diff_94000_5193000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M2885 diff_82000_3097000# diff_2881000_3710000# diff_2910000_3803000# GND efet w=72500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M2886 diff_82000_3097000# diff_2269000_3389000# diff_2218000_3480000# GND efet w=177000 l=10000
+ ad=0 pd=0 as=1.927e+09 ps=488000 
M2887 diff_1715000_2865000# diff_64000_4219000# diff_82000_3097000# GND efet w=83000 l=11000
+ ad=-1.80697e+09 pd=476000 as=0 ps=0 
M2888 diff_2218000_3480000# diff_64000_4219000# diff_1732000_2882000# GND efet w=145500 l=10500
+ ad=0 pd=0 as=-1.26197e+09 ps=598000 
M2889 diff_1658000_2819000# diff_1658000_2819000# diff_94000_5193000# GND efet w=14000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M2890 diff_82000_3097000# diff_64000_4219000# diff_1501000_2924000# GND efet w=127500 l=9500
+ ad=0 pd=0 as=-7.89346e+07 ps=1.478e+06 
M2891 diff_1501000_2924000# diff_596000_3012000# diff_82000_3097000# GND efet w=112500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2892 diff_82000_3097000# diff_1603000_3122000# diff_1501000_2924000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2893 diff_1027000_3007000# diff_71000_4514000# diff_954000_2506000# GND efet w=30000 l=13000
+ ad=0 pd=0 as=1.034e+09 ps=212000 
M2894 diff_1047000_3118000# diff_71000_4514000# diff_1156000_2479000# GND efet w=29000 l=13000
+ ad=0 pd=0 as=1.208e+09 ps=230000 
M2895 diff_947000_2557000# diff_937000_2547000# diff_916000_2526000# GND efet w=140000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2896 diff_964000_2516000# diff_954000_2506000# diff_964000_2485000# GND efet w=345500 l=10500
+ ad=0 pd=0 as=-1.40093e+09 ps=1.056e+06 
M2897 diff_1125000_2750000# diff_964000_2485000# diff_964000_2485000# GND efet w=26000 l=10000
+ ad=5.46e+08 pd=94000 as=0 ps=0 
M2898 diff_1087000_2459000# diff_1087000_2459000# diff_1125000_2750000# GND efet w=26000 l=10000
+ ad=-9.14935e+08 pd=1.106e+06 as=0 ps=0 
M2899 diff_1084000_2522000# diff_1062000_2499000# diff_964000_2485000# GND efet w=336500 l=9500
+ ad=1.65065e+08 pd=646000 as=0 ps=0 
M2900 diff_82000_3097000# diff_122000_2373000# diff_133000_2383000# GND efet w=307500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2901 diff_1087000_2459000# diff_1062000_2499000# diff_1084000_2522000# GND efet w=294000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2902 diff_122000_2373000# diff_552000_1210000# diff_82000_3097000# GND efet w=416500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2903 diff_1167000_2490000# diff_1156000_2479000# diff_1087000_2459000# GND efet w=340500 l=9500
+ ad=1.45703e+09 pd=520000 as=0 ps=0 
M2904 diff_1258000_2793000# diff_67000_5287000# diff_1258000_2735000# GND efet w=15000 l=13000
+ ad=-8.68967e+08 pd=628000 as=9.79e+08 ps=180000 
M2905 diff_1458000_2942000# diff_1458000_2942000# diff_94000_5193000# GND efet w=15000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M2906 diff_1339000_3007000# diff_1339000_3007000# diff_94000_5193000# GND efet w=16000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M2907 diff_82000_3097000# diff_966000_2988000# diff_1501000_2924000# GND efet w=120000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2908 diff_1501000_2924000# diff_859000_2986000# diff_82000_3097000# GND efet w=125500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2909 diff_82000_3097000# diff_1585000_2911000# diff_1501000_2924000# GND efet w=126000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2910 diff_1501000_2924000# diff_1501000_2924000# diff_94000_5193000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M2911 diff_1458000_2942000# diff_67000_5287000# diff_1404000_2968000# GND efet w=14000 l=13000
+ ad=0 pd=0 as=6.46e+08 ps=138000 
M2912 diff_999000_2989000# diff_67000_5287000# diff_1585000_2911000# GND efet w=16000 l=13000
+ ad=0 pd=0 as=5.35e+08 ps=142000 
M2913 diff_82000_3097000# diff_93000_3550000# diff_2269000_3389000# GND efet w=63000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2914 diff_1816000_2933000# diff_93000_3550000# diff_82000_3097000# GND efet w=66500 l=10500
+ ad=1.493e+09 pd=312000 as=0 ps=0 
M2915 diff_94000_5193000# diff_1715000_2865000# diff_1715000_2865000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2916 diff_1816000_2933000# diff_1816000_2933000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2917 diff_94000_5193000# diff_1732000_2882000# diff_1732000_2882000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2918 diff_2269000_3389000# diff_2269000_3389000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2919 diff_2903000_3861000# diff_2903000_3861000# diff_94000_5193000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2920 diff_82000_3097000# diff_3023000_3903000# diff_3008000_3949000# GND efet w=44000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2921 diff_3004000_3815000# diff_67000_5287000# diff_3023000_3903000# GND efet w=13000 l=13000
+ ad=1.2e+09 pd=250000 as=3.86e+08 ps=136000 
M2922 diff_905000_3225000# diff_905000_3225000# diff_905000_3225000# GND efet w=2000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2923 diff_2910000_3803000# diff_67000_5287000# diff_2867000_3891000# GND efet w=15000 l=12000
+ ad=0 pd=0 as=7.39e+08 ps=184000 
M2924 diff_94000_5193000# diff_905000_3225000# diff_905000_3225000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M2925 diff_2910000_3803000# diff_2910000_3803000# diff_94000_5193000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2926 diff_82000_3097000# diff_3031000_3773000# diff_3004000_3815000# GND efet w=45000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2927 diff_3004000_3815000# diff_3004000_3815000# diff_94000_5193000# GND efet w=15000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M2928 diff_518000_3031000# diff_71000_4514000# diff_2659000_3492000# GND efet w=16000 l=15000
+ ad=0 pd=0 as=-2.09697e+09 ps=468000 
M2929 diff_2771000_3401000# diff_71000_4514000# diff_3031000_3773000# GND efet w=14000 l=14000
+ ad=-1.78997e+09 pd=546000 as=5.34e+08 ps=144000 
M2930 diff_82000_3097000# diff_2565000_3499000# diff_1603000_3122000# GND efet w=185000 l=10000
+ ad=0 pd=0 as=-1.04297e+09 ps=614000 
M2931 diff_82000_3097000# diff_2597000_3303000# diff_529000_4371000# GND efet w=293000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2932 diff_64000_4219000# diff_71000_4514000# diff_2881000_3710000# GND efet w=16000 l=12000
+ ad=0 pd=0 as=1.006e+09 ps=246000 
M2933 diff_529000_4371000# diff_529000_4371000# diff_94000_5193000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2934 diff_82000_3097000# diff_1839000_3082000# diff_1827000_2941000# GND efet w=186500 l=9500
+ ad=0 pd=0 as=-2.19673e+07 ps=874000 
M2935 diff_1750000_2973000# diff_1750000_2973000# diff_94000_5193000# GND efet w=14000 l=23000
+ ad=-1.56997e+09 pd=584000 as=0 ps=0 
M2936 diff_1809000_2941000# diff_64000_4219000# diff_1750000_2973000# GND efet w=177000 l=11000
+ ad=1.239e+09 pd=368000 as=0 ps=0 
M2937 diff_1827000_2941000# diff_1816000_2933000# diff_1809000_2941000# GND efet w=177000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2938 diff_82000_3097000# diff_742000_2973000# diff_1827000_2941000# GND efet w=27000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2939 diff_82000_3097000# diff_73000_3121000# diff_1839000_3082000# GND efet w=80500 l=10500
+ ad=0 pd=0 as=1.91e+09 ps=394000 
M2940 diff_1936000_3037000# diff_1809000_946000# diff_82000_3097000# GND efet w=117500 l=10500
+ ad=-6.01967e+08 pd=638000 as=0 ps=0 
M2941 diff_1961000_3116000# diff_67000_5287000# diff_2003000_3054000# GND efet w=14000 l=14000
+ ad=2.84e+08 pd=80000 as=-1.07897e+09 ps=572000 
M2942 diff_1999000_3197000# diff_71000_4514000# diff_1697000_2847000# GND efet w=15000 l=14000
+ ad=4.39e+08 pd=112000 as=-3.74967e+08 ps=828000 
M2943 diff_82000_3097000# diff_742000_2973000# diff_1827000_2941000# GND efet w=157500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2944 diff_1839000_3082000# diff_1839000_3082000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2945 diff_1555000_2818000# diff_71000_4514000# diff_1553000_2585000# GND efet w=22000 l=14000
+ ad=0 pd=0 as=9.37e+08 ps=164000 
M2946 diff_1189000_3106000# diff_71000_4514000# diff_1609000_2778000# GND efet w=23000 l=15000
+ ad=0 pd=0 as=9.06e+08 ps=160000 
M2947 diff_1658000_2819000# diff_71000_4514000# diff_1658000_2776000# GND efet w=23000 l=15000
+ ad=0 pd=0 as=9.98e+08 ps=162000 
M2948 diff_82000_3097000# diff_1961000_3116000# diff_1962000_2986000# GND efet w=71000 l=10000
+ ad=0 pd=0 as=2.126e+09 ps=434000 
M2949 diff_2003000_3054000# diff_1999000_3197000# diff_82000_3097000# GND efet w=65000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2950 diff_2109000_2944000# diff_71000_4514000# diff_2081000_3200000# GND efet w=15000 l=13000
+ ad=-1.08497e+09 pd=592000 as=6.5e+08 ps=150000 
M2951 diff_2652000_3483000# diff_2641000_3474000# diff_82000_3097000# GND efet w=136500 l=10500
+ ad=1.03e+09 pd=288000 as=0 ps=0 
M2952 diff_2634000_3303000# diff_2659000_3492000# diff_2652000_3483000# GND efet w=136000 l=10000
+ ad=-5.16967e+08 pd=662000 as=0 ps=0 
M2953 diff_82000_3097000# diff_93000_3550000# diff_2659000_3492000# GND efet w=67000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M2954 diff_3228000_4781000# diff_3228000_4781000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2955 diff_3047000_3538000# diff_67000_5287000# diff_2877000_4621000# GND efet w=15000 l=13000
+ ad=5.14e+08 pd=142000 as=0 ps=0 
M2956 diff_94000_5193000# diff_1603000_3122000# diff_1603000_3122000# GND efet w=15000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2957 diff_2634000_3303000# diff_2634000_3303000# diff_94000_5193000# GND efet w=15000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2958 diff_2634000_3303000# diff_67000_5287000# diff_2597000_3303000# GND efet w=24000 l=14000
+ ad=0 pd=0 as=4.93e+08 ps=106000 
M2959 diff_2065000_3012000# diff_2003000_3054000# diff_82000_3097000# GND efet w=117000 l=11000
+ ad=-2.10097e+09 pd=510000 as=0 ps=0 
M2960 diff_82000_3097000# diff_2081000_3200000# diff_2065000_3012000# GND efet w=117500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M2961 diff_2133000_3059000# diff_1096000_3118000# diff_82000_3097000# GND efet w=67000 l=10000
+ ad=-1.07197e+09 pd=562000 as=0 ps=0 
M2962 diff_2003000_3054000# diff_2003000_3054000# diff_94000_5193000# GND efet w=16000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M2963 diff_94000_5193000# diff_1962000_2986000# diff_1962000_2986000# GND efet w=13000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2964 diff_94000_5193000# diff_1936000_3037000# diff_1936000_3037000# GND efet w=16000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M2965 diff_2065000_3012000# diff_2065000_3012000# diff_94000_5193000# GND efet w=15000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M2966 diff_2133000_3059000# diff_2133000_3059000# diff_94000_5193000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2967 diff_82000_3097000# diff_2197000_2999000# diff_2292000_3173000# GND efet w=154500 l=9500
+ ad=0 pd=0 as=-7.63967e+08 ps=748000 
M2968 diff_82000_3097000# diff_2197000_2999000# diff_2183000_3047000# GND efet w=42000 l=11000
+ ad=0 pd=0 as=-1.89967e+08 ps=866000 
M2969 diff_2183000_3047000# diff_2133000_3059000# diff_82000_3097000# GND efet w=132000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2970 diff_82000_3097000# diff_2247000_3125000# diff_2183000_3047000# GND efet w=148000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2971 diff_2292000_3173000# diff_2247000_3125000# diff_82000_3097000# GND efet w=145000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2972 diff_2183000_3047000# diff_2172000_3037000# diff_2109000_2944000# GND efet w=155000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2973 diff_82000_3097000# diff_2197000_2999000# diff_2183000_3047000# GND efet w=105000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2974 diff_2355000_3006000# diff_2350000_3073000# diff_2292000_3173000# GND efet w=135000 l=10000
+ ad=-1.45597e+09 pd=428000 as=0 ps=0 
M2975 diff_2391000_3200000# diff_71000_4514000# diff_2355000_3006000# GND efet w=15000 l=14000
+ ad=2.81e+08 pd=104000 as=0 ps=0 
M2976 diff_2133000_3059000# diff_71000_4514000# diff_2419000_3101000# GND efet w=15000 l=13000
+ ad=0 pd=0 as=2.35e+08 ps=76000 
M2977 diff_2399000_2875000# diff_2391000_3200000# diff_82000_3097000# GND efet w=80000 l=11000
+ ad=1.427e+09 pd=316000 as=0 ps=0 
M2978 diff_82000_3097000# diff_2419000_3101000# diff_2399000_2875000# GND efet w=85000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2979 diff_82000_3097000# diff_2463000_2894000# diff_1258000_2793000# GND efet w=122000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2980 diff_1936000_3037000# diff_2182000_2692000# diff_2247000_3125000# GND efet w=15000 l=13000
+ ad=0 pd=0 as=1.8e+08 ps=54000 
M2981 diff_2109000_2944000# diff_2109000_2944000# diff_94000_5193000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2982 diff_1697000_2847000# diff_71000_4514000# diff_1711000_2777000# GND efet w=22000 l=15000
+ ad=0 pd=0 as=1.016e+09 ps=162000 
M2983 diff_1715000_2865000# diff_71000_4514000# diff_1775000_2769000# GND efet w=14000 l=13000
+ ad=0 pd=0 as=1.13e+09 ps=168000 
M2984 diff_1732000_2882000# diff_71000_4514000# diff_1815000_2508000# GND efet w=17000 l=14000
+ ad=0 pd=0 as=1.219e+09 ps=172000 
M2985 diff_1750000_2973000# diff_71000_4514000# diff_1873000_2768000# GND efet w=16000 l=13000
+ ad=0 pd=0 as=1.111e+09 ps=168000 
M2986 diff_1309000_2729000# diff_1277000_2573000# diff_1277000_2573000# GND efet w=15000 l=11000
+ ad=1.26e+09 pd=184000 as=2.10327e+07 ps=548000 
M2987 diff_1309000_2729000# diff_1317000_2486000# diff_1317000_2486000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=1.441e+09 ps=326000 
M2988 diff_1277000_2573000# diff_1258000_2735000# diff_1243000_2573000# GND efet w=118000 l=10000
+ ad=0 pd=0 as=-1.46297e+09 ps=284000 
M2989 diff_1280000_2491000# diff_1151000_1006000# diff_1277000_2573000# GND efet w=205500 l=10500
+ ad=2.136e+09 pd=474000 as=0 ps=0 
M2990 diff_133000_2006000# diff_122000_2206000# diff_82000_3097000# GND efet w=882500 l=10500
+ ad=2.04623e+09 pd=4.28e+06 as=0 ps=0 
M2991 diff_82000_3097000# diff_122000_2206000# diff_133000_2006000# GND efet w=307000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2992 diff_82000_3097000# diff_553000_2340000# diff_122000_2206000# GND efet w=416500 l=10500
+ ad=0 pd=0 as=1.51507e+09 ps=1.284e+06 
M2993 diff_1328000_2491000# diff_1317000_2486000# diff_1280000_2491000# GND efet w=200000 l=11000
+ ad=1.04707e+09 pd=998000 as=0 ps=0 
M2994 diff_1392000_2557000# diff_1392000_2557000# diff_1410000_2714000# GND efet w=14000 l=23000
+ ad=-1.00897e+09 pd=584000 as=5.81e+08 ps=124000 
M2995 diff_1513000_2747000# diff_1485000_2491000# diff_1485000_2491000# GND efet w=15000 l=11000
+ ad=6.82e+08 pd=136000 as=-9.31967e+08 ps=602000 
M2996 diff_1328000_2491000# diff_1333000_2957000# diff_1317000_2486000# GND efet w=79500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M2997 diff_1392000_2557000# diff_1333000_2957000# diff_1328000_2491000# GND efet w=74500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M2998 diff_1457000_2547000# diff_1447000_2541000# diff_1392000_2557000# GND efet w=83000 l=10000
+ ad=2.014e+09 pd=364000 as=0 ps=0 
M2999 diff_1328000_2491000# diff_1392000_2557000# diff_1384000_2467000# GND efet w=150500 l=11500
+ ad=0 pd=0 as=-1.63297e+09 ps=428000 
M3000 diff_1485000_2491000# diff_1333000_2957000# diff_1457000_2547000# GND efet w=162000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3001 diff_1590000_2747000# diff_1486000_840000# diff_1486000_840000# GND efet w=23000 l=9000
+ ad=5.18e+08 pd=92000 as=2.10403e+09 ps=1.006e+06 
M3002 diff_1546000_931000# diff_1546000_931000# diff_1590000_2747000# GND efet w=17000 l=10000
+ ad=5.90327e+07 pd=912000 as=0 ps=0 
M3003 diff_1507000_2551000# diff_1236000_1920000# diff_1485000_2491000# GND efet w=190000 l=11000
+ ad=-1.97797e+09 pd=388000 as=0 ps=0 
M3004 diff_82000_3097000# diff_581000_2216000# diff_122000_2206000# GND efet w=415500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3005 diff_82000_3097000# diff_122000_2206000# diff_133000_2006000# GND efet w=242000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3006 diff_857000_2350000# diff_847000_2341000# diff_82000_3097000# GND efet w=134000 l=10000
+ ad=1.689e+09 pd=330000 as=0 ps=0 
M3007 diff_94000_5193000# diff_857000_2350000# diff_857000_2350000# GND efet w=14000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3008 diff_816000_2341000# diff_801000_877000# diff_801000_877000# GND efet w=14000 l=105000
+ ad=-2.0159e+09 pd=2.218e+06 as=-1.14497e+09 ps=706000 
M3009 diff_94000_5193000# diff_913000_2209000# diff_913000_2209000# GND efet w=15000 l=9000
+ ad=0 pd=0 as=2.042e+09 ps=432000 
M3010 diff_969000_2376000# diff_890000_2283000# diff_931000_2160000# GND efet w=106500 l=10500
+ ad=-1.79797e+09 pd=506000 as=-8.98902e+08 ps=1.668e+06 
M3011 diff_931000_2160000# diff_816000_2341000# diff_913000_2209000# GND efet w=145000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3012 diff_94000_5193000# diff_969000_2376000# diff_969000_2376000# GND efet w=15000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3013 diff_1065000_2210000# diff_1065000_2210000# diff_94000_5193000# GND efet w=15000 l=23000
+ ad=-1.83797e+09 pd=452000 as=0 ps=0 
M3014 diff_890000_2283000# diff_876000_1127000# diff_857000_2350000# GND efet w=21000 l=13000
+ ad=4.2e+08 pd=82000 as=0 ps=0 
M3015 diff_913000_2209000# diff_900000_990000# diff_890000_2283000# GND efet w=21000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M3016 diff_450000_2165000# diff_122000_1996000# diff_133000_2006000# GND efet w=240500 l=10500
+ ad=-1.84093e+09 pd=652000 as=0 ps=0 
M3017 diff_122000_2206000# diff_122000_2206000# diff_450000_2165000# GND efet w=37000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3018 diff_581000_2216000# diff_679000_2183000# diff_718000_2179000# GND efet w=36000 l=13000
+ ad=5.16e+08 pd=106000 as=1.1e+09 ps=212000 
M3019 diff_450000_2165000# diff_122000_1996000# diff_122000_1996000# GND efet w=43000 l=11000
+ ad=0 pd=0 as=-1.9059e+09 ps=1.358e+06 
M3020 diff_133000_2006000# diff_122000_1996000# diff_105000_1847000# GND efet w=857000 l=11000
+ ad=0 pd=0 as=5.10131e+08 ps=2.114e+06 
M3021 diff_450000_2113000# diff_122000_1996000# diff_133000_2006000# GND efet w=240500 l=10500
+ ad=2.079e+09 pd=240000 as=0 ps=0 
M3022 diff_82000_3097000# diff_586000_2094000# diff_122000_1996000# GND efet w=181000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3023 diff_450000_2036000# diff_122000_1996000# diff_133000_2006000# GND efet w=344500 l=10500
+ ad=-1.81897e+09 pd=346000 as=0 ps=0 
M3024 diff_82000_3097000# diff_586000_2094000# diff_122000_1996000# GND efet w=271000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3025 diff_122000_1996000# diff_552000_1999000# diff_82000_3097000# GND efet w=415000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3026 diff_133000_1629000# diff_122000_1840000# diff_105000_1847000# GND efet w=861000 l=11000
+ ad=1.65923e+09 pd=4.28e+06 as=0 ps=0 
M3027 diff_82000_3097000# diff_552000_1210000# diff_122000_1840000# GND efet w=415500 l=10500
+ ad=0 pd=0 as=-1.6719e+09 ps=1.368e+06 
M3028 diff_94000_5193000# diff_122000_1840000# diff_133000_1629000# GND efet w=344500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3029 diff_82000_3097000# diff_122000_1619000# diff_122000_1840000# GND efet w=272000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3030 diff_94000_5193000# diff_122000_1840000# diff_133000_1629000# GND efet w=240500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3031 diff_82000_3097000# diff_122000_1619000# diff_122000_1840000# GND efet w=183000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3032 diff_94000_5193000# diff_122000_1840000# diff_133000_1629000# GND efet w=240500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3033 diff_122000_1840000# diff_122000_1840000# diff_94000_5193000# GND efet w=44000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3034 diff_801000_877000# diff_801000_877000# diff_816000_2039000# GND efet w=14000 l=105000
+ ad=0 pd=0 as=3.81e+08 ps=80000 
M3035 diff_857000_2021000# diff_847000_2015000# diff_82000_3097000# GND efet w=132000 l=10000
+ ad=1.672e+09 pd=332000 as=0 ps=0 
M3036 diff_1009000_2203000# diff_890000_2283000# diff_931000_2160000# GND efet w=38000 l=10000
+ ad=1.471e+09 pd=358000 as=0 ps=0 
M3037 diff_969000_2376000# diff_890000_2283000# diff_931000_2160000# GND efet w=49000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3038 diff_1009000_2203000# diff_890000_2283000# diff_931000_2160000# GND efet w=79500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3039 diff_1065000_2210000# diff_1036000_876000# diff_1009000_2203000# GND efet w=123000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3040 diff_1086000_2210000# diff_969000_2376000# diff_1065000_2210000# GND efet w=75500 l=10500
+ ad=1.342e+09 pd=332000 as=0 ps=0 
M3041 diff_82000_3097000# diff_1093000_1019000# diff_1086000_2210000# GND efet w=141000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3042 diff_1086000_2210000# diff_969000_2376000# diff_1065000_2210000# GND efet w=47000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3043 diff_1151000_1006000# diff_1065000_2210000# diff_82000_3097000# GND efet w=86000 l=10000
+ ad=9.95164e+08 pd=3.402e+06 as=0 ps=0 
M3044 diff_1151000_1006000# diff_1065000_2210000# diff_82000_3097000# GND efet w=45000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3045 diff_931000_2160000# diff_921000_2149000# diff_913000_2133000# GND efet w=143000 l=10000
+ ad=0 pd=0 as=2.041e+09 ps=430000 
M3046 diff_890000_2093000# diff_876000_1127000# diff_857000_2021000# GND efet w=21000 l=13000
+ ad=4.2e+08 pd=82000 as=0 ps=0 
M3047 diff_913000_2133000# diff_900000_990000# diff_890000_2093000# GND efet w=21000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M3048 diff_969000_2014000# diff_961000_2107000# diff_931000_2160000# GND efet w=49000 l=10000
+ ad=-1.71597e+09 pd=510000 as=0 ps=0 
M3049 diff_1009000_2186000# diff_1003000_2176000# diff_931000_2160000# GND efet w=82000 l=10000
+ ad=1.397e+09 pd=360000 as=0 ps=0 
M3050 diff_969000_2014000# diff_961000_2107000# diff_931000_2160000# GND efet w=104000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3051 diff_874000_2000000# diff_857000_2021000# diff_857000_2021000# GND efet w=14000 l=10000
+ ad=9.78e+08 pd=190000 as=0 ps=0 
M3052 diff_857000_1973000# diff_847000_1964000# diff_82000_3097000# GND efet w=134000 l=10000
+ ad=1.736e+09 pd=330000 as=0 ps=0 
M3053 diff_874000_2000000# diff_857000_1973000# diff_857000_1973000# GND efet w=15000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3054 diff_816000_1964000# diff_801000_877000# diff_801000_877000# GND efet w=14000 l=105000
+ ad=2.99e+08 pd=70000 as=0 ps=0 
M3055 diff_940000_2000000# diff_913000_2133000# diff_913000_2133000# GND efet w=15000 l=9000
+ ad=9.94e+08 pd=196000 as=0 ps=0 
M3056 diff_1009000_2186000# diff_1003000_2176000# diff_931000_2160000# GND efet w=39000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3057 diff_1065000_2063000# diff_1036000_876000# diff_1009000_2186000# GND efet w=123000 l=11000
+ ad=-1.78597e+09 pd=460000 as=0 ps=0 
M3058 diff_1086000_2100000# diff_1075000_2090000# diff_1065000_2063000# GND efet w=46000 l=11000
+ ad=1.378e+09 pd=326000 as=0 ps=0 
M3059 diff_82000_3097000# diff_1093000_1019000# diff_1086000_2100000# GND efet w=139000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3060 diff_1086000_2100000# diff_1075000_2090000# diff_1065000_2063000# GND efet w=74000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3061 diff_1151000_1006000# diff_1130000_2112000# diff_82000_3097000# GND efet w=45000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3062 diff_1013000_2000000# diff_969000_2014000# diff_969000_2014000# GND efet w=15000 l=10000
+ ad=1.006e+09 pd=192000 as=0 ps=0 
M3063 diff_940000_2000000# diff_913000_1832000# diff_913000_1832000# GND efet w=15000 l=9000
+ ad=0 pd=0 as=2.066e+09 ps=430000 
M3064 diff_969000_1999000# diff_961000_1837000# diff_931000_1783000# GND efet w=106500 l=10500
+ ad=-1.72397e+09 pd=506000 as=-1.0019e+09 ps=1.67e+06 
M3065 diff_931000_1783000# diff_921000_1827000# diff_913000_1832000# GND efet w=144000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3066 diff_1013000_2000000# diff_969000_1999000# diff_969000_1999000# GND efet w=14000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3067 diff_1065000_2063000# diff_1065000_2063000# diff_1049000_1986000# GND efet w=16000 l=23000
+ ad=0 pd=0 as=1.07e+09 ps=146000 
M3068 diff_1065000_1833000# diff_1065000_1833000# diff_1049000_1986000# GND efet w=15000 l=23000
+ ad=-1.83497e+09 pd=454000 as=0 ps=0 
M3069 diff_1151000_1006000# diff_1130000_2112000# diff_82000_3097000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3070 diff_890000_1906000# diff_876000_1127000# diff_857000_1973000# GND efet w=21000 l=12000
+ ad=4.2e+08 pd=82000 as=0 ps=0 
M3071 diff_913000_1832000# diff_900000_990000# diff_890000_1906000# GND efet w=21000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M3072 diff_133000_1629000# diff_122000_1619000# diff_82000_3097000# GND efet w=879000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3073 diff_82000_3097000# diff_122000_1619000# diff_133000_1629000# GND efet w=242000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3074 diff_94000_5193000# diff_122000_1619000# diff_122000_1619000# GND efet w=37000 l=10000
+ ad=0 pd=0 as=1.33607e+09 ps=1.28e+06 
M3075 diff_718000_1785000# diff_679000_1018000# diff_581000_1717000# GND efet w=36000 l=13000
+ ad=1.039e+09 pd=206000 as=5.88e+08 ps=112000 
M3076 diff_82000_3097000# diff_581000_1717000# diff_122000_1619000# GND efet w=414500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3077 diff_82000_3097000# diff_122000_1619000# diff_133000_1629000# GND efet w=307000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3078 diff_122000_1619000# diff_552000_1210000# diff_82000_3097000# GND efet w=417500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3079 diff_801000_877000# diff_801000_877000# diff_816000_1662000# GND efet w=14000 l=106000
+ ad=0 pd=0 as=3.65e+08 ps=78000 
M3080 diff_857000_1644000# diff_847000_1638000# diff_82000_3097000# GND efet w=132000 l=10000
+ ad=1.667e+09 pd=330000 as=0 ps=0 
M3081 diff_1009000_1826000# diff_1003000_1837000# diff_931000_1783000# GND efet w=39000 l=10000
+ ad=1.512e+09 pd=360000 as=0 ps=0 
M3082 diff_969000_1999000# diff_961000_1837000# diff_931000_1783000# GND efet w=50000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3083 diff_1009000_1826000# diff_1003000_1837000# diff_931000_1783000# GND efet w=79000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3084 diff_1065000_1833000# diff_1036000_876000# diff_1009000_1826000# GND efet w=124000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3085 diff_1086000_1833000# diff_1075000_1826000# diff_1065000_1833000# GND efet w=76500 l=10500
+ ad=1.327e+09 pd=332000 as=0 ps=0 
M3086 diff_82000_3097000# diff_1093000_1019000# diff_1086000_1833000# GND efet w=142500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3087 diff_1086000_1833000# diff_1075000_1826000# diff_1065000_1833000# GND efet w=47000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3088 diff_1151000_1006000# diff_1130000_1886000# diff_82000_3097000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3089 diff_1151000_1006000# diff_1130000_1886000# diff_82000_3097000# GND efet w=45000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3090 diff_931000_1783000# diff_921000_1772000# diff_913000_1756000# GND efet w=143000 l=10000
+ ad=0 pd=0 as=2.041e+09 ps=430000 
M3091 diff_133000_1252000# diff_122000_1452000# diff_82000_3097000# GND efet w=884500 l=10500
+ ad=1.52423e+09 pd=4.288e+06 as=0 ps=0 
M3092 diff_82000_3097000# diff_122000_1452000# diff_133000_1252000# GND efet w=307000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3093 diff_82000_3097000# diff_553000_1586000# diff_122000_1452000# GND efet w=416500 l=10500
+ ad=0 pd=0 as=1.51407e+09 ps=1.284e+06 
M3094 diff_889000_1716000# diff_876000_1127000# diff_857000_1644000# GND efet w=21000 l=12000
+ ad=4.2e+08 pd=82000 as=0 ps=0 
M3095 diff_913000_1756000# diff_900000_990000# diff_889000_1716000# GND efet w=21000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M3096 diff_969000_1637000# diff_961000_1731000# diff_931000_1783000# GND efet w=49000 l=10000
+ ad=-1.73197e+09 pd=512000 as=0 ps=0 
M3097 diff_1009000_1809000# diff_1003000_1799000# diff_931000_1783000# GND efet w=82000 l=10000
+ ad=1.396e+09 pd=360000 as=0 ps=0 
M3098 diff_969000_1637000# diff_961000_1731000# diff_931000_1783000# GND efet w=103500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3099 diff_874000_1624000# diff_857000_1644000# diff_857000_1644000# GND efet w=13000 l=10000
+ ad=9.67e+08 pd=190000 as=0 ps=0 
M3100 diff_82000_3097000# diff_581000_1462000# diff_122000_1452000# GND efet w=415500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3101 diff_82000_3097000# diff_122000_1452000# diff_133000_1252000# GND efet w=242500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M3102 diff_857000_1596000# diff_847000_1587000# diff_82000_3097000# GND efet w=134000 l=10000
+ ad=1.715e+09 pd=328000 as=0 ps=0 
M3103 diff_874000_1624000# diff_857000_1596000# diff_857000_1596000# GND efet w=15000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3104 diff_816000_1587000# diff_801000_877000# diff_801000_877000# GND efet w=14000 l=105000
+ ad=-2.0279e+09 pd=2.192e+06 as=0 ps=0 
M3105 diff_940000_1623000# diff_913000_1756000# diff_913000_1756000# GND efet w=15000 l=9000
+ ad=9.94e+08 pd=196000 as=0 ps=0 
M3106 diff_1009000_1809000# diff_1003000_1799000# diff_931000_1783000# GND efet w=39000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3107 diff_1065000_1686000# diff_1036000_876000# diff_1009000_1809000# GND efet w=123000 l=11000
+ ad=-1.81797e+09 pd=456000 as=0 ps=0 
M3108 diff_1086000_1724000# diff_1075000_1713000# diff_1065000_1686000# GND efet w=46000 l=11000
+ ad=1.361e+09 pd=328000 as=0 ps=0 
M3109 diff_82000_3097000# diff_1093000_1019000# diff_1086000_1724000# GND efet w=140000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3110 diff_1086000_1724000# diff_1075000_1713000# diff_1065000_1686000# GND efet w=74000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3111 diff_1151000_1006000# diff_1130000_1735000# diff_82000_3097000# GND efet w=45000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3112 diff_1013000_1623000# diff_969000_1637000# diff_969000_1637000# GND efet w=15000 l=10000
+ ad=1.006e+09 pd=192000 as=0 ps=0 
M3113 diff_940000_1623000# diff_913000_1455000# diff_913000_1455000# GND efet w=15000 l=9000
+ ad=0 pd=0 as=2.066e+09 ps=430000 
M3114 diff_969000_1622000# diff_890000_1529000# diff_931000_1406000# GND efet w=106500 l=10500
+ ad=-1.74497e+09 pd=504000 as=-9.86902e+08 ps=1.668e+06 
M3115 diff_931000_1406000# diff_816000_1587000# diff_913000_1455000# GND efet w=144000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3116 diff_1013000_1623000# diff_969000_1622000# diff_969000_1622000# GND efet w=14000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3117 diff_1065000_1686000# diff_1065000_1686000# diff_1049000_1609000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=1.068e+09 ps=146000 
M3118 diff_1064000_1456000# diff_1064000_1456000# diff_1049000_1609000# GND efet w=15000 l=23000
+ ad=-1.71097e+09 pd=456000 as=0 ps=0 
M3119 diff_1151000_1006000# diff_1130000_1735000# diff_82000_3097000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3120 diff_94000_5193000# diff_1188000_2358000# diff_1188000_2358000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=1.517e+09 ps=280000 
M3121 diff_1486000_840000# diff_1553000_2585000# diff_1541000_2447000# GND efet w=297500 l=10500
+ ad=0 pd=0 as=-4.39967e+08 ps=616000 
M3122 diff_1591000_2479000# diff_1581000_2469000# diff_1486000_840000# GND efet w=255000 l=10000
+ ad=3.41033e+08 pd=508000 as=0 ps=0 
M3123 diff_1546000_931000# diff_1581000_2469000# diff_1591000_2479000# GND efet w=233500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3124 diff_1643000_2549000# diff_1609000_2778000# diff_1546000_931000# GND efet w=257500 l=10500
+ ad=-4.39673e+07 pd=540000 as=0 ps=0 
M3125 diff_1642000_832000# diff_1658000_2776000# diff_1643000_2549000# GND efet w=248000 l=11000
+ ad=-1.01967e+08 pd=906000 as=0 ps=0 
M3126 diff_1694000_2749000# diff_1642000_832000# diff_1642000_832000# GND efet w=19000 l=10000
+ ad=4.18e+08 pd=82000 as=0 ps=0 
M3127 diff_1695000_985000# diff_1695000_985000# diff_1694000_2749000# GND efet w=19000 l=10000
+ ad=6.45033e+08 pd=918000 as=0 ps=0 
M3128 diff_1694000_2536000# diff_1684000_2526000# diff_1642000_832000# GND efet w=203000 l=10000
+ ad=-2.24967e+08 pd=438000 as=0 ps=0 
M3129 diff_1695000_985000# diff_1684000_2526000# diff_1694000_2536000# GND efet w=203000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3130 diff_1745000_2551000# diff_1711000_2777000# diff_1695000_985000# GND efet w=248500 l=9500
+ ad=4.42033e+08 pd=552000 as=0 ps=0 
M3131 diff_1779000_2705000# diff_1727000_2244000# diff_1727000_2244000# GND efet w=15000 l=17000
+ ad=6.32e+08 pd=112000 as=-1.74497e+09 ps=540000 
M3132 diff_1934000_2757000# diff_1930000_2738000# diff_1930000_2738000# GND efet w=14000 l=17000
+ ad=6.38e+08 pd=110000 as=1.355e+09 ps=270000 
M3133 diff_1977000_2723000# diff_1912000_2695000# diff_1986000_2692000# GND efet w=14000 l=12000
+ ad=5.69e+08 pd=106000 as=-1.22497e+09 ps=448000 
M3134 diff_1727000_2244000# diff_1756000_2491000# diff_1745000_2551000# GND efet w=104000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3135 diff_1797000_2536000# diff_1775000_2769000# diff_1727000_2244000# GND efet w=121500 l=9500
+ ad=1.878e+09 pd=262000 as=0 ps=0 
M3136 diff_1728000_2090000# diff_1815000_2508000# diff_1797000_2536000# GND efet w=110000 l=10000
+ ad=2.118e+09 pd=510000 as=0 ps=0 
M3137 diff_1836000_2676000# diff_1728000_2090000# diff_1728000_2090000# GND efet w=13000 l=16000
+ ad=-1.11597e+09 pd=270000 as=0 ps=0 
M3138 diff_1728000_1867000# diff_1728000_1867000# diff_1836000_2676000# GND efet w=13000 l=16000
+ ad=-1.82897e+09 pd=488000 as=0 ps=0 
M3139 diff_1930000_2738000# diff_1912000_2695000# diff_1915000_2537000# GND efet w=123500 l=9500
+ ad=0 pd=0 as=-6.18935e+08 ps=562000 
M3140 diff_1986000_2692000# diff_1967000_2491000# diff_1915000_2537000# GND efet w=172000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M3141 diff_2012000_2519000# diff_1930000_2738000# diff_1986000_2692000# GND efet w=178500 l=10500
+ ad=-1.53197e+09 pd=378000 as=0 ps=0 
M3142 diff_1846000_2538000# diff_1836000_2528000# diff_1728000_2090000# GND efet w=110000 l=10000
+ ad=-6.52967e+08 pd=282000 as=0 ps=0 
M3143 diff_1728000_1867000# diff_1836000_2528000# diff_1846000_2538000# GND efet w=109000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3144 diff_1915000_2537000# diff_1873000_2768000# diff_1728000_1867000# GND efet w=109500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3145 diff_2355000_3006000# diff_2355000_3006000# diff_94000_5193000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3146 diff_2399000_2875000# diff_2399000_2875000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3147 diff_1962000_2986000# diff_2052000_2804000# diff_2059000_2776000# GND efet w=23500 l=15500
+ ad=0 pd=0 as=1.009e+09 ps=162000 
M3148 diff_1258000_2793000# diff_1258000_2793000# diff_94000_5193000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M3149 diff_2562000_3212000# diff_71000_4514000# diff_2520000_3104000# GND efet w=16000 l=14000
+ ad=-1.01967e+08 pd=750000 as=2.84e+08 ps=100000 
M3150 diff_2463000_2894000# diff_2520000_3104000# diff_82000_3097000# GND efet w=82000 l=10000
+ ad=1.532e+09 pd=338000 as=0 ps=0 
M3151 diff_82000_3097000# diff_2399000_2875000# diff_2463000_2894000# GND efet w=81500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3152 diff_2562000_3212000# diff_2572000_3038000# diff_82000_3097000# GND efet w=72000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3153 diff_2463000_2894000# diff_2463000_2894000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3154 diff_82000_3097000# diff_2197000_2999000# diff_2562000_3212000# GND efet w=67000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3155 diff_3016000_3538000# diff_71000_4514000# diff_3013000_3474000# GND efet w=14000 l=13000
+ ad=4.68e+08 pd=144000 as=-7.15967e+08 ps=708000 
M3156 diff_82000_3097000# diff_2789000_3478000# diff_2771000_3401000# GND efet w=79500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3157 diff_82000_3097000# diff_93000_3550000# diff_2820000_3542000# GND efet w=68000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M3158 diff_82000_3097000# diff_2820000_3542000# diff_2809000_3351000# GND efet w=44000 l=11000
+ ad=0 pd=0 as=-1.21397e+09 ps=598000 
M3159 diff_3381000_4293000# diff_1252000_4406000# diff_3358000_4500000# GND efet w=201500 l=9500
+ ad=1.72e+09 pd=420000 as=0 ps=0 
M3160 diff_3400000_4293000# diff_3270000_4961000# diff_3381000_4293000# GND efet w=201500 l=10500
+ ad=1.477e+09 pd=420000 as=0 ps=0 
M3161 diff_82000_3097000# diff_3407000_4287000# diff_3400000_4293000# GND efet w=203500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3162 diff_3420000_4637000# diff_3407000_4287000# diff_82000_3097000# GND efet w=44000 l=11000
+ ad=2.069e+09 pd=474000 as=0 ps=0 
M3163 diff_3495000_4369000# diff_3359000_4961000# diff_82000_3097000# GND efet w=150500 l=10500
+ ad=1.524e+09 pd=318000 as=0 ps=0 
M3164 diff_3400000_3460000# diff_518000_3031000# diff_3495000_4369000# GND efet w=144000 l=10000
+ ad=-1.75597e+09 pd=606000 as=0 ps=0 
M3165 diff_3536000_4388000# diff_3388000_4961000# diff_3400000_3460000# GND efet w=150000 l=10000
+ ad=1.383e+09 pd=320000 as=0 ps=0 
M3166 diff_82000_3097000# diff_1000000_4393000# diff_3536000_4388000# GND efet w=152500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3167 diff_3420000_4637000# diff_3420000_4637000# diff_3420000_4637000# GND efet w=500 l=1500
+ ad=0 pd=0 as=0 ps=0 
M3168 diff_3420000_4637000# diff_3420000_4637000# diff_94000_5193000# GND efet w=15000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M3169 diff_3271000_3282000# diff_3359000_4961000# diff_82000_3097000# GND efet w=51500 l=9500
+ ad=8.93e+08 pd=224000 as=0 ps=0 
M3170 diff_2771000_3401000# diff_2771000_3401000# diff_94000_5193000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3171 diff_3271000_3282000# diff_3271000_3282000# diff_94000_5193000# GND efet w=14000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M3172 diff_529000_4371000# diff_71000_4514000# diff_3338000_4041000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=2.22e+08 ps=94000 
M3173 diff_3349000_3930000# diff_3338000_4041000# diff_3326000_3885000# GND efet w=146000 l=10000
+ ad=1.168e+09 pd=308000 as=-1.97297e+09 ps=472000 
M3174 diff_82000_3097000# diff_2605000_4946000# diff_3349000_3930000# GND efet w=146000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3175 diff_2789000_3478000# diff_67000_5287000# diff_2809000_3351000# GND efet w=16000 l=13000
+ ad=2.72e+08 pd=88000 as=0 ps=0 
M3176 diff_2809000_3351000# diff_2809000_3351000# diff_94000_5193000# GND efet w=15000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M3177 diff_2562000_3212000# diff_2133000_3059000# diff_82000_3097000# GND efet w=69500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3178 diff_82000_3097000# diff_2350000_3073000# diff_2562000_3212000# GND efet w=78500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3179 diff_2677000_3054000# diff_905000_3225000# diff_82000_3097000# GND efet w=74000 l=10000
+ ad=1.862e+09 pd=428000 as=0 ps=0 
M3180 diff_82000_3097000# diff_401000_4712000# diff_2677000_3054000# GND efet w=83000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3181 diff_1936000_3037000# diff_2182000_2692000# diff_2572000_3038000# GND efet w=15000 l=13000
+ ad=0 pd=0 as=3.25e+08 ps=100000 
M3182 diff_2562000_3212000# diff_2562000_3212000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3183 diff_2677000_3054000# diff_2677000_3054000# diff_94000_5193000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3184 diff_1658000_2819000# diff_2052000_2804000# diff_2112000_2777000# GND efet w=23000 l=15000
+ ad=0 pd=0 as=1.022e+09 ps=164000 
M3185 diff_2065000_3012000# diff_2182000_2692000# diff_2207000_2716000# GND efet w=20000 l=14000
+ ad=0 pd=0 as=1.065e+09 ps=254000 
M3186 diff_990000_3075000# diff_71000_4514000# diff_2528000_2776000# GND efet w=21500 l=15500
+ ad=0 pd=0 as=1.003e+09 ps=162000 
M3187 diff_1836000_1363000# diff_2059000_2776000# diff_2046000_2527000# GND efet w=248000 l=10000
+ ad=7.52033e+08 pd=1.046e+06 as=-1.36967e+08 ps=520000 
M3188 diff_2094000_2748000# diff_1836000_1363000# diff_1836000_1363000# GND efet w=20000 l=10000
+ ad=4.6e+08 pd=86000 as=0 ps=0 
M3189 diff_1857000_1018000# diff_1857000_1018000# diff_2094000_2748000# GND efet w=20000 l=9000
+ ad=6.45033e+08 pd=976000 as=0 ps=0 
M3190 diff_2095000_2536000# diff_2084000_2526000# diff_1836000_1363000# GND efet w=203500 l=10500
+ ad=-3.87967e+08 pd=438000 as=0 ps=0 
M3191 diff_1857000_1018000# diff_2084000_2526000# diff_2095000_2536000# GND efet w=204500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3192 diff_2147000_2552000# diff_2112000_2777000# diff_1857000_1018000# GND efet w=246500 l=10500
+ ad=-1.31967e+08 pd=524000 as=0 ps=0 
M3193 diff_2230000_2466000# diff_2230000_2466000# diff_2224000_2739000# GND efet w=20000 l=11000
+ ad=2.30327e+07 pd=722000 as=6.39e+08 ps=138000 
M3194 diff_2185000_2629000# diff_2185000_2629000# diff_2170000_2654000# GND efet w=21000 l=11000
+ ad=-9.46967e+08 pd=624000 as=1.13e+09 ps=218000 
M3195 diff_2219000_2489000# diff_2199000_2471000# diff_2185000_2629000# GND efet w=201500 l=10500
+ ad=-7.67967e+08 pd=468000 as=0 ps=0 
M3196 diff_2230000_2466000# diff_2207000_2716000# diff_2219000_2489000# GND efet w=224000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3197 diff_1251000_2260000# diff_1236000_1920000# diff_94000_5193000# GND efet w=14000 l=10000
+ ad=-2.69673e+07 pd=604000 as=0 ps=0 
M3198 diff_1195000_2101000# diff_1065000_2210000# diff_1175000_1642000# GND efet w=156500 l=10500
+ ad=4.33033e+08 pd=680000 as=-9.64902e+08 ps=2.104e+06 
M3199 diff_1188000_2358000# diff_1065000_2210000# diff_1195000_2101000# GND efet w=61000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3200 diff_1344000_2359000# diff_1344000_2359000# diff_94000_5193000# GND efet w=13000 l=22000
+ ad=-1.60897e+09 pd=534000 as=0 ps=0 
M3201 diff_1246000_2014000# diff_1188000_2358000# diff_1251000_2260000# GND efet w=53000 l=12000
+ ad=5.96033e+08 pd=802000 as=0 ps=0 
M3202 diff_94000_5193000# diff_1304000_2338000# diff_1304000_2338000# GND efet w=14000 l=26000
+ ad=0 pd=0 as=1.42e+09 ps=306000 
M3203 diff_1438000_2360000# diff_1354000_780000# diff_1344000_2359000# GND efet w=23000 l=13000
+ ad=2.29e+08 pd=66000 as=0 ps=0 
M3204 diff_1461000_2360000# diff_1439000_785000# diff_1438000_2360000# GND efet w=23500 l=13500
+ ad=4.01e+08 pd=120000 as=0 ps=0 
M3205 diff_1391000_2313000# diff_969000_2376000# diff_1344000_2359000# GND efet w=80500 l=9500
+ ad=1.208e+09 pd=292000 as=0 ps=0 
M3206 diff_1195000_2101000# diff_1184000_2091000# diff_1175000_1642000# GND efet w=157500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3207 diff_1246000_2014000# diff_1188000_2358000# diff_1251000_2260000# GND efet w=56000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M3208 diff_1188000_2022000# diff_1184000_2091000# diff_1195000_2101000# GND efet w=62000 l=10000
+ ad=1.409e+09 pd=270000 as=0 ps=0 
M3209 diff_1304000_2338000# diff_1251000_2260000# diff_1304000_2116000# GND efet w=65000 l=10000
+ ad=0 pd=0 as=2.37065e+08 ps=1.354e+06 
M3210 diff_1304000_2116000# diff_969000_2376000# diff_1304000_2338000# GND efet w=64500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3211 diff_1344000_2359000# diff_1304000_2338000# diff_1304000_2116000# GND efet w=52000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3212 diff_1391000_2313000# diff_969000_2376000# diff_1344000_2359000# GND efet w=26000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3213 diff_1304000_2116000# diff_1251000_2260000# diff_1391000_2313000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3214 diff_1188000_2022000# diff_1188000_2022000# diff_1194000_2002000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=1.038e+09 ps=174000 
M3215 diff_1246000_1991000# diff_1263000_2096000# diff_1246000_2014000# GND efet w=37000 l=12000
+ ad=7.14033e+08 pd=786000 as=0 ps=0 
M3216 diff_1304000_2037000# diff_1302000_2091000# diff_1304000_2116000# GND efet w=64000 l=10000
+ ad=1.402e+09 pd=308000 as=0 ps=0 
M3217 diff_1304000_2116000# diff_1334000_2128000# diff_1304000_2037000# GND efet w=64500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3218 diff_1246000_2014000# diff_1236000_1920000# diff_1194000_2002000# GND efet w=16000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3219 diff_1246000_1991000# diff_1263000_2096000# diff_1246000_2014000# GND efet w=73000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M3220 diff_1344000_2015000# diff_1304000_2037000# diff_1304000_2116000# GND efet w=52000 l=10000
+ ad=-1.64697e+09 pd=538000 as=0 ps=0 
M3221 diff_1391000_2051000# diff_1381000_2129000# diff_1344000_2015000# GND efet w=27000 l=10000
+ ad=1.202e+09 pd=288000 as=0 ps=0 
M3222 diff_1304000_2116000# diff_1402000_2164000# diff_1391000_2051000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3223 diff_1391000_2051000# diff_1381000_2129000# diff_1344000_2015000# GND efet w=77500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3224 diff_1304000_2037000# diff_1304000_2037000# diff_1312000_1986000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=1.504e+09 ps=170000 
M3225 diff_1194000_2002000# diff_1188000_1978000# diff_1188000_1978000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=1.527e+09 ps=272000 
M3226 diff_1246000_1991000# diff_1236000_1920000# diff_1194000_2002000# GND efet w=15000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3227 diff_1478000_2223000# diff_1461000_2360000# diff_82000_3097000# GND efet w=197500 l=9500
+ ad=-7.51967e+08 pd=688000 as=0 ps=0 
M3228 diff_1518000_2376000# diff_1478000_2223000# diff_1478000_2223000# GND efet w=15000 l=24000
+ ad=4.47e+08 pd=86000 as=0 ps=0 
M3229 diff_1575000_2219000# diff_1577000_2342000# diff_1577000_2378000# GND efet w=15000 l=35000
+ ad=9.63e+08 pd=182000 as=4.39e+08 ps=84000 
M3230 diff_1584000_2230000# diff_1577000_2342000# diff_1557000_2303000# GND efet w=14500 l=76500
+ ad=-4.81967e+08 pd=728000 as=5.29e+08 ps=188000 
M3231 diff_1655000_2366000# diff_1577000_2342000# diff_1584000_2230000# GND efet w=14000 l=24000
+ ad=4.74e+08 pd=88000 as=0 ps=0 
M3232 diff_1478000_2223000# diff_1486000_840000# diff_847000_2341000# GND efet w=110500 l=12500
+ ad=0 pd=0 as=1.64403e+09 ps=1.224e+06 
M3233 diff_1557000_2303000# diff_1546000_931000# diff_1478000_2223000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3234 diff_1478000_2075000# diff_1461000_2014000# diff_82000_3097000# GND efet w=205500 l=9500
+ ad=1.553e+09 pd=302000 as=0 ps=0 
M3235 diff_1513000_2024000# diff_1486000_840000# diff_1503000_2076000# GND efet w=111500 l=11500
+ ad=2.026e+09 pd=386000 as=1.125e+09 ps=242000 
M3236 diff_847000_2341000# diff_1642000_832000# diff_1584000_2230000# GND efet w=104500 l=12500
+ ad=0 pd=0 as=0 ps=0 
M3237 diff_1575000_2219000# diff_1557000_2303000# diff_82000_3097000# GND efet w=72500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3238 diff_1584000_2230000# diff_1575000_2219000# diff_82000_3097000# GND efet w=211000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3239 diff_816000_2341000# diff_1695000_985000# diff_1584000_2230000# GND efet w=106000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M3240 diff_1584000_2156000# diff_1575000_2145000# diff_82000_3097000# GND efet w=211000 l=10000
+ ad=-1.43697e+09 pd=490000 as=0 ps=0 
M3241 diff_1584000_2058000# diff_1557000_2075000# diff_82000_3097000# GND efet w=80500 l=9500
+ ad=9.77e+08 pd=180000 as=0 ps=0 
M3242 diff_1557000_2075000# diff_1546000_931000# diff_1513000_2024000# GND efet w=20000 l=11000
+ ad=5.65e+08 pd=174000 as=0 ps=0 
M3243 diff_1344000_2015000# diff_1344000_2015000# diff_1312000_1986000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3244 diff_1438000_2014000# diff_1354000_780000# diff_1344000_2015000# GND efet w=23000 l=14000
+ ad=2.3e+08 pd=66000 as=0 ps=0 
M3245 diff_1461000_2014000# diff_1439000_785000# diff_1438000_2014000# GND efet w=23000 l=13000
+ ad=4.12e+08 pd=110000 as=0 ps=0 
M3246 diff_1195000_1873000# diff_1184000_1863000# diff_1175000_1642000# GND efet w=154500 l=10500
+ ad=2.02303e+09 pd=798000 as=0 ps=0 
M3247 diff_1188000_1978000# diff_1184000_1863000# diff_1195000_1873000# GND efet w=60000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3248 diff_1344000_1982000# diff_1344000_1982000# diff_1312000_1986000# GND efet w=14000 l=22000
+ ad=-1.62897e+09 pd=532000 as=0 ps=0 
M3249 diff_1264000_1695000# diff_1263000_1901000# diff_1246000_1991000# GND efet w=55000 l=12000
+ ad=-6.59673e+07 pd=660000 as=0 ps=0 
M3250 diff_1312000_1986000# diff_1304000_1961000# diff_1304000_1961000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=1.435e+09 ps=308000 
M3251 diff_1438000_1983000# diff_1354000_780000# diff_1344000_1982000# GND efet w=23000 l=14000
+ ad=2.3e+08 pd=66000 as=0 ps=0 
M3252 diff_1461000_1983000# diff_1439000_785000# diff_1438000_1983000# GND efet w=23000 l=13000
+ ad=4.02e+08 pd=120000 as=0 ps=0 
M3253 diff_1391000_1936000# diff_1381000_1874000# diff_1344000_1982000# GND efet w=79500 l=9500
+ ad=1.197e+09 pd=290000 as=0 ps=0 
M3254 diff_1195000_1873000# diff_1188000_1668000# diff_1175000_1642000# GND efet w=127500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3255 diff_1264000_1695000# diff_1263000_1901000# diff_1246000_1991000# GND efet w=57000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M3256 diff_1201000_1632000# diff_1175000_1642000# diff_1195000_1873000# GND efet w=169500 l=11500
+ ad=4.89033e+08 pd=782000 as=0 ps=0 
M3257 diff_1195000_1873000# diff_1188000_1668000# diff_1175000_1642000# GND efet w=33000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3258 diff_1304000_1961000# diff_1302000_1910000# diff_1304000_1739000# GND efet w=65000 l=10000
+ ad=0 pd=0 as=2.37065e+08 ps=1.352e+06 
M3259 diff_1304000_1739000# diff_1334000_1840000# diff_1304000_1961000# GND efet w=65500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3260 diff_1344000_1982000# diff_1304000_1961000# diff_1304000_1739000# GND efet w=52000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3261 diff_1391000_1936000# diff_1381000_1874000# diff_1344000_1982000# GND efet w=26000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3262 diff_1304000_1739000# diff_1402000_1836000# diff_1391000_1936000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3263 diff_1304000_1660000# diff_1302000_1714000# diff_1304000_1739000# GND efet w=64000 l=10000
+ ad=1.4e+09 pd=306000 as=0 ps=0 
M3264 diff_1304000_1739000# diff_1334000_1751000# diff_1304000_1660000# GND efet w=64500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3265 diff_1344000_1638000# diff_1304000_1660000# diff_1304000_1739000# GND efet w=52000 l=10000
+ ad=-1.60497e+09 pd=538000 as=0 ps=0 
M3266 diff_1391000_1673000# diff_1381000_1752000# diff_1344000_1638000# GND efet w=27000 l=10000
+ ad=1.21e+09 pd=290000 as=0 ps=0 
M3267 diff_1304000_1739000# diff_1402000_1787000# diff_1391000_1673000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3268 diff_1264000_1695000# diff_1236000_1920000# diff_1258000_1634000# GND efet w=14000 l=11000
+ ad=0 pd=0 as=1.316e+09 ps=174000 
M3269 diff_1391000_1673000# diff_1381000_1752000# diff_1344000_1638000# GND efet w=78500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3270 diff_1304000_1660000# diff_1304000_1660000# diff_1312000_1609000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=1.506e+09 ps=170000 
M3271 diff_1258000_1634000# diff_1236000_1920000# diff_1201000_1632000# GND efet w=14000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3272 diff_890000_1529000# diff_876000_1127000# diff_857000_1596000# GND efet w=21000 l=13000
+ ad=4.2e+08 pd=82000 as=0 ps=0 
M3273 diff_913000_1455000# diff_900000_990000# diff_890000_1529000# GND efet w=21000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M3274 diff_450000_1411000# diff_122000_1242000# diff_133000_1252000# GND efet w=240500 l=10500
+ ad=-1.79793e+09 pd=652000 as=0 ps=0 
M3275 diff_122000_1452000# diff_122000_1452000# diff_450000_1411000# GND efet w=37000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3276 diff_581000_1462000# diff_679000_1428000# diff_718000_1425000# GND efet w=36000 l=13000
+ ad=5.16e+08 pd=106000 as=1.188e+09 ps=212000 
M3277 diff_450000_1411000# diff_122000_1242000# diff_122000_1242000# GND efet w=44000 l=11000
+ ad=0 pd=0 as=-1.9199e+09 ps=1.36e+06 
M3278 diff_133000_1252000# diff_122000_1242000# diff_104000_1093000# GND efet w=859000 l=11000
+ ad=0 pd=0 as=8.98131e+08 ps=2.116e+06 
M3279 diff_450000_1359000# diff_122000_1242000# diff_133000_1252000# GND efet w=240500 l=11500
+ ad=1.98e+09 pd=238000 as=0 ps=0 
M3280 diff_82000_3097000# diff_586000_1340000# diff_122000_1242000# GND efet w=180000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3281 diff_450000_1282000# diff_122000_1242000# diff_133000_1252000# GND efet w=344000 l=11000
+ ad=-1.88597e+09 pd=342000 as=0 ps=0 
M3282 diff_82000_3097000# diff_586000_1340000# diff_122000_1242000# GND efet w=271000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3283 diff_122000_1242000# diff_552000_1245000# diff_82000_3097000# GND efet w=415500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3284 diff_801000_877000# diff_801000_877000# diff_816000_1285000# GND efet w=14000 l=105000
+ ad=0 pd=0 as=3.65e+08 ps=78000 
M3285 diff_857000_1266000# diff_847000_1261000# diff_82000_3097000# GND efet w=133000 l=10000
+ ad=1.684e+09 pd=334000 as=0 ps=0 
M3286 diff_1009000_1449000# diff_890000_1529000# diff_931000_1406000# GND efet w=39000 l=10000
+ ad=1.512e+09 pd=360000 as=0 ps=0 
M3287 diff_969000_1622000# diff_890000_1529000# diff_931000_1406000# GND efet w=49000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3288 diff_1009000_1449000# diff_890000_1529000# diff_931000_1406000# GND efet w=79000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3289 diff_1064000_1456000# diff_1036000_876000# diff_1009000_1449000# GND efet w=124000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3290 diff_1086000_1456000# diff_969000_1622000# diff_1064000_1456000# GND efet w=76500 l=10500
+ ad=1.329e+09 pd=332000 as=0 ps=0 
M3291 diff_82000_3097000# diff_1093000_1019000# diff_1086000_1456000# GND efet w=142000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3292 diff_1086000_1456000# diff_969000_1622000# diff_1064000_1456000# GND efet w=47000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3293 diff_1151000_1006000# diff_1064000_1456000# diff_82000_3097000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3294 diff_94000_5193000# diff_1197000_1523000# diff_1197000_1523000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=1.181e+09 ps=232000 
M3295 diff_1478000_1847000# diff_1461000_1983000# diff_82000_3097000# GND efet w=197500 l=9500
+ ad=-7.01967e+08 pd=682000 as=0 ps=0 
M3296 diff_1513000_2024000# diff_1513000_2024000# diff_1519000_1998000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=5.1e+08 ps=94000 
M3297 diff_1519000_1998000# diff_1478000_1847000# diff_1478000_1847000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3298 diff_1669000_2093000# diff_1642000_832000# diff_1584000_2156000# GND efet w=101000 l=12000
+ ad=1.018e+09 pd=194000 as=0 ps=0 
M3299 diff_82000_3097000# diff_1727000_2244000# diff_816000_2341000# GND efet w=90000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M3300 diff_1707000_2129000# diff_1695000_985000# diff_1687000_2095000# GND efet w=106000 l=12000
+ ad=1.698e+09 pd=326000 as=9.6e+08 ps=228000 
M3301 diff_1584000_2058000# diff_1577000_1964000# diff_1577000_2001000# GND efet w=14000 l=35000
+ ad=0 pd=0 as=4.82e+08 ps=90000 
M3302 diff_1584000_2156000# diff_1577000_1964000# diff_1557000_2075000# GND efet w=14500 l=81500
+ ad=0 pd=0 as=0 ps=0 
M3303 diff_1584000_2156000# diff_1577000_1964000# diff_1655000_1988000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=8.9e+08 ps=132000 
M3304 diff_1577000_2001000# diff_1577000_1964000# diff_1575000_1842000# GND efet w=15000 l=35000
+ ad=0 pd=0 as=9.48e+08 ps=180000 
M3305 diff_1584000_1853000# diff_1577000_1964000# diff_1557000_1926000# GND efet w=14500 l=78500
+ ad=-4.30967e+08 pd=722000 as=5.37e+08 ps=186000 
M3306 diff_1655000_1988000# diff_1577000_1964000# diff_1584000_1853000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3307 diff_1478000_1847000# diff_1486000_840000# diff_1503000_1891000# GND efet w=110500 l=12500
+ ad=0 pd=0 as=1.53003e+09 ps=1.224e+06 
M3308 diff_1557000_1926000# diff_1546000_931000# diff_1478000_1847000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3309 diff_1478000_1698000# diff_1461000_1637000# diff_82000_3097000# GND efet w=206500 l=9500
+ ad=1.562e+09 pd=304000 as=0 ps=0 
M3310 diff_1513000_1647000# diff_1486000_840000# diff_1503000_1699000# GND efet w=111500 l=11500
+ ad=2.116e+09 pd=388000 as=1.015e+09 ps=240000 
M3311 diff_1740000_2095000# diff_1728000_2090000# diff_1707000_2129000# GND efet w=89000 l=12000
+ ad=1.587e+09 pd=262000 as=0 ps=0 
M3312 diff_1503000_1891000# diff_1642000_832000# diff_1584000_1853000# GND efet w=104000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M3313 diff_1575000_1842000# diff_1557000_1926000# diff_82000_3097000# GND efet w=73500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3314 diff_1584000_1853000# diff_1575000_1842000# diff_82000_3097000# GND efet w=211000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3315 diff_1707000_1881000# diff_1695000_985000# diff_1584000_1853000# GND efet w=105000 l=12000
+ ad=-2.0289e+09 pd=2.156e+06 as=0 ps=0 
M3316 diff_1584000_1779000# diff_1575000_1767000# diff_82000_3097000# GND efet w=211000 l=10000
+ ad=-1.37697e+09 pd=486000 as=0 ps=0 
M3317 diff_1584000_1682000# diff_1557000_1697000# diff_82000_3097000# GND efet w=80500 l=9500
+ ad=9.6e+08 pd=178000 as=0 ps=0 
M3318 diff_1557000_1697000# diff_1546000_931000# diff_1513000_1647000# GND efet w=21000 l=11000
+ ad=5.52e+08 pd=176000 as=0 ps=0 
M3319 diff_1344000_1638000# diff_1344000_1638000# diff_1312000_1609000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3320 diff_1438000_1637000# diff_1354000_780000# diff_1344000_1638000# GND efet w=23000 l=13000
+ ad=2.3e+08 pd=66000 as=0 ps=0 
M3321 diff_1461000_1637000# diff_1439000_785000# diff_1438000_1637000# GND efet w=23000 l=13000
+ ad=4.13e+08 pd=110000 as=0 ps=0 
M3322 diff_1344000_1605000# diff_1344000_1605000# diff_1312000_1609000# GND efet w=14000 l=22000
+ ad=-1.59897e+09 pd=534000 as=0 ps=0 
M3323 diff_1201000_1632000# diff_1197000_1523000# diff_1235000_1425000# GND efet w=122000 l=12000
+ ad=0 pd=0 as=-1.71967e+08 ps=646000 
M3324 diff_1151000_1006000# diff_1064000_1456000# diff_82000_3097000# GND efet w=45000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3325 diff_931000_1406000# diff_921000_1395000# diff_913000_1379000# GND efet w=143000 l=10000
+ ad=0 pd=0 as=2.062e+09 ps=434000 
M3326 diff_133000_875000# diff_122000_1086000# diff_104000_1093000# GND efet w=860500 l=10500
+ ad=1.51023e+09 pd=4.28e+06 as=0 ps=0 
M3327 diff_82000_3097000# diff_552000_1210000# diff_122000_1086000# GND efet w=415000 l=11000
+ ad=0 pd=0 as=-1.9419e+09 ps=1.362e+06 
M3328 diff_94000_5193000# diff_122000_1086000# diff_133000_875000# GND efet w=345000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3329 diff_890000_1339000# diff_876000_1127000# diff_857000_1266000# GND efet w=21000 l=13000
+ ad=4.2e+08 pd=82000 as=0 ps=0 
M3330 diff_913000_1379000# diff_900000_990000# diff_890000_1339000# GND efet w=21000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M3331 diff_969000_1260000# diff_961000_1354000# diff_931000_1406000# GND efet w=49000 l=10000
+ ad=-1.72997e+09 pd=514000 as=0 ps=0 
M3332 diff_1009000_1432000# diff_1003000_1422000# diff_931000_1406000# GND efet w=82000 l=10000
+ ad=1.396e+09 pd=360000 as=0 ps=0 
M3333 diff_969000_1260000# diff_961000_1354000# diff_931000_1406000# GND efet w=103500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3334 diff_874000_1246000# diff_857000_1266000# diff_857000_1266000# GND efet w=14000 l=10000
+ ad=9.68e+08 pd=190000 as=0 ps=0 
M3335 diff_82000_3097000# diff_122000_865000# diff_122000_1086000# GND efet w=271000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3336 diff_94000_5193000# diff_122000_1086000# diff_133000_875000# GND efet w=240500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3337 diff_82000_3097000# diff_122000_865000# diff_122000_1086000# GND efet w=182500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3338 diff_94000_5193000# diff_122000_1086000# diff_133000_875000# GND efet w=241000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3339 diff_122000_1086000# diff_122000_1086000# diff_94000_5193000# GND efet w=45000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3340 diff_857000_1219000# diff_847000_1210000# diff_82000_3097000# GND efet w=133000 l=10000
+ ad=1.683e+09 pd=324000 as=0 ps=0 
M3341 diff_874000_1246000# diff_857000_1219000# diff_857000_1219000# GND efet w=15000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3342 diff_816000_1210000# diff_801000_877000# diff_801000_877000# GND efet w=14000 l=105000
+ ad=1.31507e+09 pd=2.022e+06 as=0 ps=0 
M3343 diff_940000_1246000# diff_913000_1379000# diff_913000_1379000# GND efet w=16000 l=9000
+ ad=9.98e+08 pd=196000 as=0 ps=0 
M3344 diff_1009000_1432000# diff_1003000_1422000# diff_931000_1406000# GND efet w=39000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3345 diff_1064000_1309000# diff_1036000_876000# diff_1009000_1432000# GND efet w=123000 l=10000
+ ad=-1.66897e+09 pd=462000 as=0 ps=0 
M3346 diff_1086000_1347000# diff_1075000_1336000# diff_1064000_1309000# GND efet w=46000 l=11000
+ ad=1.35e+09 pd=326000 as=0 ps=0 
M3347 diff_82000_3097000# diff_1093000_1019000# diff_1086000_1347000# GND efet w=139500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3348 diff_1086000_1347000# diff_1075000_1336000# diff_1064000_1309000# GND efet w=74000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3349 diff_1151000_1006000# diff_1130000_1358000# diff_82000_3097000# GND efet w=45000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3350 diff_1197000_1523000# diff_1064000_1456000# diff_1175000_1427000# GND efet w=54000 l=10000
+ ad=0 pd=0 as=5.70327e+07 ps=496000 
M3351 diff_1235000_1425000# diff_1187000_1276000# diff_1235000_1244000# GND efet w=121500 l=11500
+ ad=0 pd=0 as=8.40327e+07 ps=756000 
M3352 diff_1013000_1246000# diff_969000_1260000# diff_969000_1260000# GND efet w=15000 l=10000
+ ad=9.96e+08 pd=192000 as=0 ps=0 
M3353 diff_940000_1246000# diff_913000_1078000# diff_913000_1078000# GND efet w=15000 l=9000
+ ad=0 pd=0 as=2.08e+09 ps=430000 
M3354 diff_774000_468000# diff_890000_1152000# diff_931000_1029000# GND efet w=106500 l=10500
+ ad=-1.72497e+09 pd=506000 as=-9.36902e+08 ps=1.67e+06 
M3355 diff_931000_1029000# diff_816000_1210000# diff_913000_1078000# GND efet w=144000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3356 diff_1013000_1246000# diff_774000_468000# diff_774000_468000# GND efet w=14000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3357 diff_1064000_1309000# diff_1064000_1309000# diff_1049000_1232000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=1.047e+09 ps=144000 
M3358 diff_1065000_1079000# diff_1065000_1079000# diff_1049000_1232000# GND efet w=15000 l=23000
+ ad=-1.83497e+09 pd=454000 as=0 ps=0 
M3359 diff_1151000_1006000# diff_1130000_1358000# diff_82000_3097000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3360 diff_890000_1152000# diff_876000_1127000# diff_857000_1219000# GND efet w=21000 l=14000
+ ad=4.2e+08 pd=82000 as=0 ps=0 
M3361 diff_913000_1078000# diff_900000_990000# diff_890000_1152000# GND efet w=21000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M3362 diff_133000_875000# diff_122000_865000# diff_82000_3097000# GND efet w=878500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3363 diff_82000_3097000# diff_122000_865000# diff_133000_875000# GND efet w=242500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3364 diff_94000_5193000# diff_122000_865000# diff_122000_865000# GND efet w=37000 l=11000
+ ad=0 pd=0 as=1.23407e+09 ps=1.28e+06 
M3365 diff_718000_1031000# diff_679000_1018000# diff_581000_963000# GND efet w=36000 l=14000
+ ad=-2.03897e+09 pd=440000 as=5.52e+08 ps=110000 
M3366 diff_82000_3097000# diff_581000_963000# diff_122000_865000# GND efet w=417000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3367 diff_82000_3097000# diff_122000_865000# diff_133000_875000# GND efet w=307500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3368 diff_122000_865000# diff_552000_1210000# diff_82000_3097000# GND efet w=417000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3369 diff_801000_877000# diff_801000_877000# diff_816000_908000# GND efet w=14000 l=106000
+ ad=0 pd=0 as=3.65e+08 ps=78000 
M3370 diff_857000_889000# diff_847000_884000# diff_82000_3097000# GND efet w=133000 l=10000
+ ad=1.702e+09 pd=332000 as=0 ps=0 
M3371 diff_1009000_1072000# diff_890000_1152000# diff_931000_1029000# GND efet w=40000 l=10000
+ ad=1.481e+09 pd=360000 as=0 ps=0 
M3372 diff_774000_468000# diff_890000_1152000# diff_931000_1029000# GND efet w=50000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3373 diff_1009000_1072000# diff_890000_1152000# diff_931000_1029000# GND efet w=79500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3374 diff_1065000_1079000# diff_1036000_876000# diff_1009000_1072000# GND efet w=124000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3375 diff_1086000_1079000# diff_774000_468000# diff_1065000_1079000# GND efet w=76500 l=10500
+ ad=1.328e+09 pd=332000 as=0 ps=0 
M3376 diff_82000_3097000# diff_1093000_1019000# diff_1086000_1079000# GND efet w=142500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3377 diff_1086000_1079000# diff_774000_468000# diff_1065000_1079000# GND efet w=47000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3378 diff_1151000_1006000# diff_1065000_1079000# diff_82000_3097000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3379 diff_1151000_1006000# diff_1065000_1079000# diff_82000_3097000# GND efet w=45000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3380 diff_931000_1029000# diff_921000_1018000# diff_913000_1002000# GND efet w=143000 l=10000
+ ad=0 pd=0 as=2.111e+09 ps=432000 
M3381 diff_890000_962000# diff_876000_1127000# diff_857000_889000# GND efet w=21000 l=13000
+ ad=4.2e+08 pd=82000 as=0 ps=0 
M3382 diff_913000_1002000# diff_900000_990000# diff_890000_962000# GND efet w=21000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M3383 diff_969000_883000# diff_961000_976000# diff_931000_1029000# GND efet w=49000 l=10000
+ ad=9.54033e+08 pd=954000 as=0 ps=0 
M3384 diff_1009000_1055000# diff_1003000_1045000# diff_931000_1029000# GND efet w=82000 l=10000
+ ad=1.396e+09 pd=360000 as=0 ps=0 
M3385 diff_969000_883000# diff_961000_976000# diff_931000_1029000# GND efet w=104000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3386 diff_873000_870000# diff_857000_889000# diff_857000_889000# GND efet w=14000 l=10000
+ ad=6.85e+08 pd=138000 as=0 ps=0 
M3387 diff_133000_497000# diff_122000_699000# diff_82000_3097000# GND efet w=881500 l=10500
+ ad=1.16823e+09 pd=4.228e+06 as=0 ps=0 
M3388 diff_82000_3097000# diff_122000_699000# diff_133000_497000# GND efet w=306500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3389 diff_82000_3097000# diff_553000_832000# diff_122000_699000# GND efet w=409000 l=11000
+ ad=0 pd=0 as=1.37007e+09 ps=1.274e+06 
M3390 diff_940000_870000# diff_913000_1002000# diff_913000_1002000# GND efet w=15000 l=9000
+ ad=6.71e+08 pd=136000 as=0 ps=0 
M3391 diff_1009000_1055000# diff_1003000_1045000# diff_931000_1029000# GND efet w=39000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3392 diff_1065000_932000# diff_1036000_876000# diff_1009000_1055000# GND efet w=123000 l=11000
+ ad=-1.83097e+09 pd=460000 as=0 ps=0 
M3393 diff_1086000_970000# diff_1075000_959000# diff_1065000_932000# GND efet w=46000 l=11000
+ ad=1.349e+09 pd=326000 as=0 ps=0 
M3394 diff_82000_3097000# diff_1093000_1019000# diff_1086000_970000# GND efet w=139000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3395 diff_1086000_970000# diff_1075000_959000# diff_1065000_932000# GND efet w=74000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3396 diff_1151000_1006000# diff_1130000_981000# diff_82000_3097000# GND efet w=45000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3397 diff_1187000_1276000# diff_1189000_1317000# diff_1175000_1427000# GND efet w=52500 l=9500
+ ad=1.931e+09 pd=404000 as=0 ps=0 
M3398 diff_1187000_1276000# diff_1187000_1276000# diff_1187000_1246000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=6.2e+08 ps=110000 
M3399 diff_1312000_1609000# diff_1304000_1584000# diff_1304000_1584000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=1.443e+09 ps=308000 
M3400 diff_1438000_1606000# diff_1354000_780000# diff_1344000_1605000# GND efet w=23000 l=13000
+ ad=2.29e+08 pd=66000 as=0 ps=0 
M3401 diff_1461000_1606000# diff_1439000_785000# diff_1438000_1606000# GND efet w=23500 l=13500
+ ad=4.12e+08 pd=118000 as=0 ps=0 
M3402 diff_1391000_1559000# diff_969000_1622000# diff_1344000_1605000# GND efet w=79500 l=9500
+ ad=1.197e+09 pd=290000 as=0 ps=0 
M3403 diff_1304000_1584000# diff_1201000_1632000# diff_1304000_1362000# GND efet w=65000 l=10000
+ ad=0 pd=0 as=2.26065e+08 ps=1.35e+06 
M3404 diff_1304000_1362000# diff_969000_1622000# diff_1304000_1584000# GND efet w=64500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3405 diff_1344000_1605000# diff_1304000_1584000# diff_1304000_1362000# GND efet w=51000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3406 diff_1391000_1559000# diff_969000_1622000# diff_1344000_1605000# GND efet w=26000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3407 diff_1304000_1362000# diff_1201000_1632000# diff_1391000_1559000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3408 diff_1304000_1283000# diff_1302000_1337000# diff_1304000_1362000# GND efet w=64000 l=10000
+ ad=1.4e+09 pd=306000 as=0 ps=0 
M3409 diff_1304000_1362000# diff_1334000_1374000# diff_1304000_1283000# GND efet w=64500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3410 diff_1344000_1261000# diff_1304000_1283000# diff_1304000_1362000# GND efet w=51000 l=10000
+ ad=-1.62797e+09 pd=538000 as=0 ps=0 
M3411 diff_1391000_1296000# diff_1381000_1375000# diff_1344000_1261000# GND efet w=27000 l=10000
+ ad=1.211e+09 pd=290000 as=0 ps=0 
M3412 diff_1304000_1362000# diff_1402000_1410000# diff_1391000_1296000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3413 diff_1391000_1296000# diff_1381000_1375000# diff_1344000_1261000# GND efet w=78500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3414 diff_1235000_1425000# diff_1236000_1920000# diff_1265000_1280000# GND efet w=15000 l=11000
+ ad=0 pd=0 as=1.11e+09 ps=162000 
M3415 diff_1304000_1283000# diff_1304000_1283000# diff_1312000_1232000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=1.504e+09 ps=170000 
M3416 diff_1187000_1246000# diff_1187000_1218000# diff_1187000_1218000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=1.446e+09 ps=276000 
M3417 diff_1265000_1280000# diff_1236000_1920000# diff_1235000_1244000# GND efet w=14000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3418 diff_1478000_1469000# diff_1461000_1606000# diff_82000_3097000# GND efet w=197500 l=9500
+ ad=-7.69967e+08 pd=684000 as=0 ps=0 
M3419 diff_1513000_1647000# diff_1513000_1647000# diff_1519000_1621000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=5.11e+08 ps=94000 
M3420 diff_1519000_1621000# diff_1478000_1469000# diff_1478000_1469000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3421 diff_1669000_1716000# diff_1642000_832000# diff_1584000_1779000# GND efet w=100500 l=11500
+ ad=1.018e+09 pd=194000 as=0 ps=0 
M3422 diff_1721000_1815000# diff_1728000_1867000# diff_1707000_1881000# GND efet w=89000 l=12000
+ ad=-1.83097e+09 pd=362000 as=0 ps=0 
M3423 diff_1707000_1752000# diff_1695000_985000# diff_1687000_1717000# GND efet w=107000 l=12000
+ ad=1.336e+09 pd=256000 as=9.75e+08 ps=230000 
M3424 diff_1584000_1682000# diff_1577000_1588000# diff_1577000_1624000# GND efet w=14000 l=36000
+ ad=0 pd=0 as=4.82e+08 ps=90000 
M3425 diff_1584000_1779000# diff_1577000_1588000# diff_1557000_1697000# GND efet w=14500 l=83500
+ ad=0 pd=0 as=0 ps=0 
M3426 diff_1584000_1779000# diff_1577000_1588000# diff_1655000_1612000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=8.76e+08 ps=130000 
M3427 diff_1577000_1624000# diff_1577000_1588000# diff_1575000_1465000# GND efet w=15000 l=34000
+ ad=0 pd=0 as=9.63e+08 ps=182000 
M3428 diff_1584000_1476000# diff_1577000_1588000# diff_1558000_1549000# GND efet w=14500 l=76500
+ ad=-4.02967e+08 pd=726000 as=5.28e+08 ps=184000 
M3429 diff_1655000_1612000# diff_1577000_1588000# diff_1584000_1476000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3430 diff_1478000_1469000# diff_1486000_840000# diff_847000_1587000# GND efet w=110000 l=12000
+ ad=0 pd=0 as=7.31033e+08 ps=1.04e+06 
M3431 diff_1558000_1549000# diff_1546000_931000# diff_1478000_1469000# GND efet w=20000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M3432 diff_1478000_1321000# diff_1461000_1260000# diff_82000_3097000# GND efet w=205500 l=9500
+ ad=1.552e+09 pd=302000 as=0 ps=0 
M3433 diff_1513000_1270000# diff_1486000_840000# diff_1503000_1322000# GND efet w=112500 l=11500
+ ad=2.038e+09 pd=388000 as=1.081e+09 ps=242000 
M3434 diff_847000_1587000# diff_1642000_832000# diff_1584000_1476000# GND efet w=104000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M3435 diff_1575000_1465000# diff_1558000_1549000# diff_82000_3097000# GND efet w=73500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3436 diff_1584000_1476000# diff_1575000_1465000# diff_82000_3097000# GND efet w=211000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3437 diff_816000_1587000# diff_1695000_985000# diff_1584000_1476000# GND efet w=105000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M3438 diff_1584000_1402000# diff_1575000_1390000# diff_82000_3097000# GND efet w=211000 l=10000
+ ad=-1.31797e+09 pd=486000 as=0 ps=0 
M3439 diff_1584000_1305000# diff_1558000_1320000# diff_82000_3097000# GND efet w=80500 l=9500
+ ad=9.6e+08 pd=178000 as=0 ps=0 
M3440 diff_1558000_1320000# diff_1546000_931000# diff_1513000_1270000# GND efet w=21000 l=12000
+ ad=5.32e+08 pd=174000 as=0 ps=0 
M3441 diff_1344000_1261000# diff_1344000_1261000# diff_1312000_1232000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3442 diff_1438000_1260000# diff_1354000_780000# diff_1344000_1261000# GND efet w=23000 l=14000
+ ad=2.3e+08 pd=66000 as=0 ps=0 
M3443 diff_1461000_1260000# diff_1439000_785000# diff_1438000_1260000# GND efet w=23000 l=13000
+ ad=4.12e+08 pd=110000 as=0 ps=0 
M3444 diff_1344000_1228000# diff_1344000_1228000# diff_1312000_1232000# GND efet w=13000 l=22000
+ ad=-1.61797e+09 pd=532000 as=0 ps=0 
M3445 diff_1187000_1218000# diff_1065000_1079000# diff_1183000_1061000# GND efet w=51000 l=10000
+ ad=0 pd=0 as=1.961e+09 ps=276000 
M3446 diff_1235000_1244000# diff_1187000_1218000# diff_1237000_974000# GND efet w=116000 l=11000
+ ad=0 pd=0 as=-1.66397e+09 ps=508000 
M3447 diff_1312000_1232000# diff_1304000_1207000# diff_1304000_1207000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=1.442e+09 ps=308000 
M3448 diff_1438000_1229000# diff_1354000_780000# diff_1344000_1228000# GND efet w=23000 l=14000
+ ad=2.3e+08 pd=66000 as=0 ps=0 
M3449 diff_1461000_1229000# diff_1439000_785000# diff_1438000_1229000# GND efet w=23000 l=13000
+ ad=4.11e+08 pd=118000 as=0 ps=0 
M3450 diff_1013000_869000# diff_969000_883000# diff_969000_883000# GND efet w=15000 l=10000
+ ad=7.44e+08 pd=138000 as=0 ps=0 
M3451 diff_82000_3097000# diff_581000_708000# diff_122000_699000# GND efet w=416000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3452 diff_82000_3097000# diff_122000_699000# diff_133000_497000# GND efet w=242500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3453 diff_450000_657000# diff_122000_487000# diff_133000_497000# GND efet w=241000 l=11000
+ ad=-2.08193e+09 pd=652000 as=0 ps=0 
M3454 diff_122000_699000# diff_122000_699000# diff_450000_657000# GND efet w=38000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3455 diff_753000_679000# diff_684000_665000# diff_581000_708000# GND efet w=37000 l=13000
+ ad=4.91e+08 pd=126000 as=4.9e+08 ps=116000 
M3456 diff_450000_657000# diff_122000_487000# diff_122000_487000# GND efet w=43000 l=11000
+ ad=0 pd=0 as=-1.7589e+09 ps=1.394e+06 
M3457 diff_450000_605000# diff_122000_487000# diff_133000_497000# GND efet w=240000 l=11000
+ ad=1.98e+09 pd=238000 as=0 ps=0 
M3458 diff_82000_3097000# diff_915000_743000# diff_876000_1127000# GND efet w=79000 l=12000
+ ad=0 pd=0 as=1.891e+09 ps=244000 
M3459 diff_900000_990000# diff_915000_743000# diff_82000_3097000# GND efet w=79000 l=12000
+ ad=1.639e+09 pd=250000 as=0 ps=0 
M3460 diff_1065000_932000# diff_1065000_932000# diff_1049000_876000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=5.85e+08 ps=100000 
M3461 diff_1151000_1006000# diff_1130000_981000# diff_82000_3097000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3462 diff_1178000_871000# diff_1151000_1006000# diff_1151000_1006000# GND efet w=14000 l=9000
+ ad=7.46e+08 pd=136000 as=0 ps=0 
M3463 diff_570000_477000# diff_588000_587000# diff_122000_487000# GND efet w=366500 l=10500
+ ad=-1.19019e+07 pd=1.432e+06 as=0 ps=0 
M3464 diff_122000_487000# diff_588000_587000# diff_570000_477000# GND efet w=40000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3465 diff_133000_497000# diff_122000_487000# diff_105000_354000# GND efet w=830500 l=10500
+ ad=0 pd=0 as=-1.39787e+09 ps=1.868e+06 
M3466 diff_450000_527000# diff_122000_487000# diff_133000_497000# GND efet w=345000 l=11000
+ ad=-1.87897e+09 pd=344000 as=0 ps=0 
M3467 diff_122000_487000# diff_561000_494000# diff_570000_477000# GND efet w=83000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3468 diff_82000_3097000# diff_826000_618000# diff_791000_355000# GND efet w=403500 l=9500
+ ad=0 pd=0 as=-1.12935e+08 ps=1.36e+06 
M3469 diff_82000_3097000# diff_905000_614000# diff_791000_355000# GND efet w=409500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3470 diff_570000_477000# diff_561000_494000# diff_122000_487000# GND efet w=383000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3471 diff_122000_487000# diff_122000_487000# diff_122000_487000# GND efet w=500 l=4500
+ ad=0 pd=0 as=0 ps=0 
M3472 diff_969000_883000# diff_989000_660000# diff_905000_614000# GND efet w=36000 l=14000
+ ad=0 pd=0 as=5.2e+08 ps=138000 
M3473 diff_1391000_1181000# diff_774000_468000# diff_1344000_1228000# GND efet w=79500 l=9500
+ ad=1.208e+09 pd=292000 as=0 ps=0 
M3474 diff_1304000_1207000# diff_1235000_1244000# diff_1304000_985000# GND efet w=65000 l=10000
+ ad=0 pd=0 as=2.19065e+08 ps=1.35e+06 
M3475 diff_1304000_985000# diff_774000_468000# diff_1304000_1207000# GND efet w=64500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3476 diff_1344000_1228000# diff_1304000_1207000# diff_1304000_985000# GND efet w=51000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3477 diff_1391000_1181000# diff_774000_468000# diff_1344000_1228000# GND efet w=27000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3478 diff_1304000_985000# diff_1235000_1244000# diff_1391000_1181000# GND efet w=107000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3479 diff_1267000_1004000# diff_1236000_1920000# diff_1237000_974000# GND efet w=15000 l=11000
+ ad=-1.63997e+09 pd=332000 as=0 ps=0 
M3480 diff_1304000_906000# diff_1302000_960000# diff_1304000_985000# GND efet w=64000 l=10000
+ ad=1.416e+09 pd=310000 as=0 ps=0 
M3481 diff_1304000_985000# diff_1334000_997000# diff_1304000_906000# GND efet w=64500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3482 diff_1344000_884000# diff_1304000_906000# diff_1304000_985000# GND efet w=51000 l=10000
+ ad=-1.68497e+09 pd=540000 as=0 ps=0 
M3483 diff_1391000_919000# diff_1381000_998000# diff_1344000_884000# GND efet w=26000 l=10000
+ ad=1.204e+09 pd=288000 as=0 ps=0 
M3484 diff_1304000_985000# diff_1402000_1033000# diff_1391000_919000# GND efet w=105000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3485 diff_1391000_919000# diff_1381000_998000# diff_1344000_884000# GND efet w=78500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3486 diff_1304000_906000# diff_1304000_906000# diff_1311000_876000# GND efet w=15000 l=25000
+ ad=0 pd=0 as=8.94e+08 ps=126000 
M3487 diff_1478000_1092000# diff_1461000_1229000# diff_82000_3097000# GND efet w=196500 l=9500
+ ad=-7.88967e+08 pd=682000 as=0 ps=0 
M3488 diff_1513000_1270000# diff_1513000_1270000# diff_1519000_1244000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=5.11e+08 ps=94000 
M3489 diff_1519000_1244000# diff_1478000_1092000# diff_1478000_1092000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3490 diff_1669000_1339000# diff_1642000_832000# diff_1584000_1402000# GND efet w=100500 l=11500
+ ad=1.018e+09 pd=194000 as=0 ps=0 
M3491 diff_1707000_1375000# diff_1695000_985000# diff_1687000_1340000# GND efet w=107000 l=12000
+ ad=1.351e+09 pd=258000 as=9.75e+08 ps=230000 
M3492 diff_1584000_1305000# diff_1577000_1211000# diff_1577000_1247000# GND efet w=14000 l=36000
+ ad=0 pd=0 as=4.82e+08 ps=90000 
M3493 diff_1584000_1402000# diff_1577000_1211000# diff_1558000_1320000# GND efet w=14500 l=82500
+ ad=0 pd=0 as=0 ps=0 
M3494 diff_1584000_1402000# diff_1577000_1211000# diff_1655000_1235000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=8.76e+08 ps=130000 
M3495 diff_1577000_1247000# diff_1577000_1211000# diff_1575000_1088000# GND efet w=15000 l=34000
+ ad=0 pd=0 as=9.64e+08 ps=182000 
M3496 diff_1584000_1099000# diff_1577000_1211000# diff_1557000_1172000# GND efet w=14500 l=77500
+ ad=-4.19967e+08 pd=724000 as=5.51e+08 ps=188000 
M3497 diff_1655000_1235000# diff_1577000_1211000# diff_1584000_1099000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3498 diff_1478000_1092000# diff_1486000_840000# diff_847000_1210000# GND efet w=110000 l=12000
+ ad=0 pd=0 as=6.87033e+08 ps=1.036e+06 
M3499 diff_1557000_1172000# diff_1546000_931000# diff_1478000_1092000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3500 diff_1478000_943000# diff_1461000_883000# diff_82000_3097000# GND efet w=204500 l=9500
+ ad=1.551e+09 pd=302000 as=0 ps=0 
M3501 diff_1513000_893000# diff_1486000_840000# diff_1503000_945000# GND efet w=112000 l=12000
+ ad=2.034e+09 pd=388000 as=1.092e+09 ps=242000 
M3502 diff_847000_1210000# diff_1642000_832000# diff_1584000_1099000# GND efet w=102500 l=12500
+ ad=0 pd=0 as=0 ps=0 
M3503 diff_1575000_1088000# diff_1557000_1172000# diff_82000_3097000# GND efet w=73500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3504 diff_1584000_1099000# diff_1575000_1088000# diff_82000_3097000# GND efet w=210000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3505 diff_816000_1210000# diff_1695000_985000# diff_1584000_1099000# GND efet w=105000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M3506 diff_1584000_1025000# diff_1575000_1013000# diff_82000_3097000# GND efet w=211000 l=10000
+ ad=-1.36997e+09 pd=490000 as=0 ps=0 
M3507 diff_1584000_927000# diff_1557000_943000# diff_82000_3097000# GND efet w=80500 l=9500
+ ad=9.74e+08 pd=180000 as=0 ps=0 
M3508 diff_1557000_943000# diff_1546000_931000# diff_1513000_893000# GND efet w=20000 l=11000
+ ad=5.61e+08 pd=172000 as=0 ps=0 
M3509 diff_1344000_884000# diff_1344000_884000# diff_1311000_876000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3510 diff_1438000_883000# diff_1354000_780000# diff_1344000_884000# GND efet w=22000 l=13000
+ ad=2.2e+08 pd=64000 as=0 ps=0 
M3511 diff_1461000_883000# diff_1439000_785000# diff_1438000_883000# GND efet w=22000 l=13000
+ ad=4.08e+08 pd=106000 as=0 ps=0 
M3512 diff_1513000_893000# diff_1513000_893000# diff_1518000_870000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=4.99e+08 ps=92000 
M3513 diff_1236000_1920000# diff_915000_743000# diff_82000_3097000# GND efet w=74000 l=12000
+ ad=1.624e+09 pd=208000 as=0 ps=0 
M3514 diff_1669000_962000# diff_1642000_832000# diff_1584000_1025000# GND efet w=101000 l=12000
+ ad=1.018e+09 pd=194000 as=0 ps=0 
M3515 diff_1707000_998000# diff_1695000_985000# diff_1687000_963000# GND efet w=108000 l=12000
+ ad=1.271e+09 pd=258000 as=1.042e+09 ps=232000 
M3516 diff_1584000_927000# diff_1577000_893000# diff_1577000_869000# GND efet w=14000 l=34000
+ ad=0 pd=0 as=4.82e+08 ps=90000 
M3517 diff_1584000_1025000# diff_1577000_893000# diff_1557000_943000# GND efet w=14500 l=81500
+ ad=0 pd=0 as=0 ps=0 
M3518 diff_1584000_1025000# diff_1577000_893000# diff_1654000_876000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=5.49e+08 ps=96000 
M3519 diff_1439000_785000# diff_1385000_840000# diff_1410000_785000# GND efet w=74000 l=11000
+ ad=-1.61897e+09 pd=430000 as=1.332e+09 ps=184000 
M3520 diff_1520000_785000# diff_1508000_759000# diff_1486000_840000# GND efet w=77000 l=12000
+ ad=1.528e+09 pd=194000 as=0 ps=0 
M3521 diff_1546000_931000# diff_1508000_759000# diff_1520000_785000# GND efet w=77000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3522 diff_1674000_771000# diff_1624000_777000# diff_1642000_832000# GND efet w=72000 l=12000
+ ad=1.512e+09 pd=186000 as=0 ps=0 
M3523 diff_1695000_985000# diff_1624000_777000# diff_1674000_771000# GND efet w=72000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M3524 diff_2248000_788000# diff_2248000_788000# diff_2337000_2732000# GND efet w=19000 l=11000
+ ad=1.12503e+09 pd=928000 as=1.759e+09 ps=268000 
M3525 diff_2337000_2732000# diff_2287000_2487000# diff_2287000_2487000# GND efet w=15000 l=25000
+ ad=0 pd=0 as=-2.08597e+09 ps=400000 
M3526 diff_2337000_2732000# diff_2326000_2476000# diff_2326000_2476000# GND efet w=14000 l=10000
+ ad=0 pd=0 as=1.56033e+08 ps=748000 
M3527 diff_2299000_2498000# diff_2287000_2487000# diff_2232000_2217000# GND efet w=137000 l=12000
+ ad=-4.10967e+08 pd=620000 as=-1.59967e+08 ps=698000 
M3528 diff_2287000_2487000# diff_2310000_2576000# diff_2299000_2498000# GND efet w=69500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3529 diff_2299000_2498000# diff_2316000_2469000# diff_2287000_2487000# GND efet w=70000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3530 diff_2326000_2476000# diff_2316000_2469000# diff_2299000_2498000# GND efet w=181500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3531 diff_2385000_2506000# diff_2374000_2501000# diff_2326000_2476000# GND efet w=174000 l=11000
+ ad=-1.22597e+09 pd=462000 as=0 ps=0 
M3532 diff_2248000_788000# diff_2283000_2432000# diff_2385000_2506000# GND efet w=201000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3533 diff_82000_3097000# diff_2961000_3295000# diff_2937000_3466000# GND efet w=64000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3534 diff_82000_3097000# diff_3016000_3538000# diff_2986000_3359000# GND efet w=44000 l=11000
+ ad=0 pd=0 as=-1.36597e+09 ps=588000 
M3535 diff_3013000_3474000# diff_3047000_3538000# diff_82000_3097000# GND efet w=81000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3536 diff_530000_4621000# diff_530000_4621000# diff_530000_4621000# GND efet w=3000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3537 diff_3326000_3885000# diff_67000_5287000# diff_3211000_3555000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=9.07e+08 ps=230000 
M3538 diff_94000_5193000# diff_530000_4621000# diff_530000_4621000# GND efet w=26000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3539 diff_3326000_3885000# diff_3326000_3885000# diff_94000_5193000# GND efet w=16000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3540 diff_3414000_3851000# diff_2605000_4946000# diff_1697000_2847000# GND efet w=205000 l=10000
+ ad=1.435e+09 pd=424000 as=0 ps=0 
M3541 diff_82000_3097000# diff_596000_3012000# diff_3414000_3851000# GND efet w=205000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3542 diff_1697000_2847000# diff_1697000_2847000# diff_94000_5193000# GND efet w=14000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M3543 diff_82000_3097000# diff_3211000_3555000# diff_530000_4621000# GND efet w=270500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3544 diff_2937000_3466000# diff_2937000_3466000# diff_94000_5193000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3545 diff_3400000_3460000# diff_3400000_3460000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3546 diff_3013000_3474000# diff_3013000_3474000# diff_94000_5193000# GND efet w=14000 l=18000
+ ad=0 pd=0 as=0 ps=0 
M3547 diff_2986000_3359000# diff_2986000_3359000# diff_94000_5193000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M3548 diff_82000_3097000# diff_3034000_4153000# diff_2987000_3090000# GND efet w=74000 l=10000
+ ad=0 pd=0 as=1.455e+09 ps=312000 
M3549 diff_3112000_3385000# diff_3105000_3437000# diff_82000_3097000# GND efet w=69000 l=11000
+ ad=1.323e+09 pd=296000 as=0 ps=0 
M3550 diff_82000_3097000# diff_783000_3632000# diff_3112000_3385000# GND efet w=81000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3551 diff_3755000_4643000# diff_790000_4021000# diff_3701000_4747000# GND efet w=85000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3552 diff_82000_3097000# diff_3624000_4961000# diff_3755000_4643000# GND efet w=91000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3553 diff_3665000_4489000# diff_3506000_4961000# diff_82000_3097000# GND efet w=150000 l=10000
+ ad=1.92033e+08 pd=824000 as=0 ps=0 
M3554 diff_3701000_4747000# diff_3701000_4747000# diff_94000_5193000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M3555 diff_94000_5193000# diff_3666000_4700000# diff_3666000_4700000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=-2.11597e+09 ps=488000 
M3556 diff_3665000_4489000# diff_790000_4021000# diff_3666000_4700000# GND efet w=153500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M3557 diff_3608000_4425000# diff_3418000_4961000# diff_82000_3097000# GND efet w=161000 l=10000
+ ad=-7.61967e+08 pd=716000 as=0 ps=0 
M3558 diff_82000_3097000# diff_3446000_4961000# diff_3608000_4425000# GND efet w=156500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3559 diff_82000_3097000# diff_3536000_4961000# diff_3665000_4489000# GND efet w=136500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3560 diff_82000_3097000# diff_3476000_4961000# diff_3657000_4141000# GND efet w=62500 l=10500
+ ad=0 pd=0 as=1.182e+09 ps=266000 
M3561 diff_3657000_4141000# diff_3657000_4141000# diff_94000_5193000# GND efet w=15000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M3562 diff_3667000_4148000# diff_3657000_4141000# diff_3608000_4425000# GND efet w=134000 l=10000
+ ad=1.072e+09 pd=284000 as=0 ps=0 
M3563 diff_3665000_4068000# diff_790000_4021000# diff_3667000_4148000# GND efet w=134000 l=10000
+ ad=-1.80497e+09 pd=486000 as=0 ps=0 
M3564 diff_94000_5193000# diff_3665000_4068000# diff_3665000_4068000# GND efet w=15000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M3565 diff_3534000_3824000# diff_67000_5287000# diff_3582000_4084000# GND efet w=15000 l=14000
+ ad=-3.37967e+08 pd=752000 as=2.5e+08 ps=100000 
M3566 diff_82000_3097000# diff_3447000_3516000# diff_3534000_3824000# GND efet w=67500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3567 diff_783000_3632000# diff_3582000_4084000# diff_82000_3097000# GND efet w=103000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3568 diff_3447000_3516000# diff_71000_4514000# diff_2569000_3911000# GND efet w=21000 l=13000
+ ad=-1.63097e+09 pd=504000 as=6.20327e+07 ps=808000 
M3569 diff_945000_3262000# diff_71000_4514000# diff_3676000_3846000# GND efet w=15000 l=12000
+ ad=0 pd=0 as=2.93e+08 ps=98000 
M3570 diff_82000_3097000# diff_3622000_3885000# diff_2569000_3911000# GND efet w=66000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3571 diff_3669000_3851000# diff_3531000_3484000# diff_3618000_3825000# GND efet w=146000 l=10000
+ ad=1.109e+09 pd=308000 as=2.111e+09 ps=472000 
M3572 diff_2987000_3090000# diff_2987000_3090000# diff_94000_5193000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3573 diff_3112000_3385000# diff_3112000_3385000# diff_94000_5193000# GND efet w=16000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M3574 diff_2734000_2819000# diff_2743000_3027000# diff_82000_3097000# GND efet w=87000 l=10000
+ ad=1.966e+09 pd=474000 as=0 ps=0 
M3575 diff_82000_3097000# diff_859000_2986000# diff_2734000_2819000# GND efet w=79000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3576 diff_2820000_3093000# diff_530000_4621000# diff_82000_3097000# GND efet w=134000 l=11000
+ ad=8.04e+08 pd=280000 as=0 ps=0 
M3577 diff_2807000_2819000# diff_511000_4351000# diff_2820000_3093000# GND efet w=134000 l=11000
+ ad=-1.55797e+09 pd=540000 as=0 ps=0 
M3578 diff_2743000_3027000# diff_67000_5287000# diff_999000_2989000# GND efet w=14000 l=13000
+ ad=2.76e+08 pd=90000 as=0 ps=0 
M3579 diff_2734000_2819000# diff_2734000_2819000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3580 diff_2807000_2819000# diff_2807000_2819000# diff_94000_5193000# GND efet w=15000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M3581 diff_2986000_3359000# diff_67000_5287000# diff_2961000_3295000# GND efet w=14000 l=13000
+ ad=0 pd=0 as=5.06e+08 ps=132000 
M3582 diff_2908000_3148000# diff_67000_5287000# diff_2873000_3144000# GND efet w=14000 l=14000
+ ad=1.721e+09 pd=348000 as=2.6e+08 ps=98000 
M3583 diff_82000_3097000# diff_2873000_3144000# diff_2601000_2819000# GND efet w=74000 l=10000
+ ad=0 pd=0 as=-1.86397e+09 ps=504000 
M3584 diff_2910000_2819000# diff_71000_4514000# diff_2921000_3077000# GND efet w=15000 l=13000
+ ad=-1.31297e+09 pd=614000 as=2.4e+08 ps=74000 
M3585 diff_82000_3097000# diff_2921000_3077000# diff_2908000_3148000# GND efet w=69500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3586 diff_2979000_3081000# diff_742000_2973000# diff_2910000_2819000# GND efet w=138000 l=10000
+ ad=1.314e+09 pd=342000 as=0 ps=0 
M3587 diff_82000_3097000# diff_2987000_3090000# diff_2979000_3081000# GND efet w=142500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3588 diff_3025000_3074000# diff_93000_3157000# diff_82000_3097000# GND efet w=136500 l=10500
+ ad=8.71e+08 pd=286000 as=0 ps=0 
M3589 diff_2908000_3148000# diff_2908000_3148000# diff_94000_5193000# GND efet w=15000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M3590 diff_2631000_2819000# diff_2987000_3090000# diff_3025000_3074000# GND efet w=135500 l=10500
+ ad=-4.34967e+08 pd=688000 as=0 ps=0 
M3591 diff_3073000_3192000# diff_71000_4514000# diff_2631000_2819000# GND efet w=15000 l=14000
+ ad=2.75e+08 pd=96000 as=0 ps=0 
M3592 diff_3121000_3079000# diff_67000_5287000# diff_3060000_3051000# GND efet w=14000 l=13000
+ ad=6.25e+08 pd=142000 as=-1.83997e+09 ps=414000 
M3593 diff_3060000_3051000# diff_3073000_3192000# diff_82000_3097000# GND efet w=65000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3594 diff_3534000_3824000# diff_3534000_3824000# diff_94000_5193000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3595 diff_82000_3097000# diff_3676000_3846000# diff_3669000_3851000# GND efet w=146000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3596 diff_3618000_3825000# diff_67000_5287000# diff_3622000_3885000# GND efet w=13000 l=13000
+ ad=0 pd=0 as=4.97e+08 ps=138000 
M3597 diff_4019000_4532000# diff_3839000_4961000# diff_82000_3097000# GND efet w=90500 l=10500
+ ad=-1.86497e+09 pd=474000 as=0 ps=0 
M3598 diff_82000_3097000# diff_3869000_4933000# diff_4019000_4532000# GND efet w=88000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M3599 diff_94000_5193000# diff_3980000_4516000# diff_3980000_4516000# GND efet w=15000 l=38000
+ ad=0 pd=0 as=-1.98393e+09 ps=1.27e+06 
M3600 diff_3980000_4516000# diff_1000000_4393000# diff_4019000_4532000# GND efet w=91500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3601 diff_3886000_4603000# diff_67000_5287000# diff_3908000_4368000# GND efet w=16000 l=13000
+ ad=2.6e+08 pd=84000 as=1.908e+09 ps=446000 
M3602 diff_783000_3632000# diff_783000_3632000# diff_94000_5193000# GND efet w=14000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M3603 diff_3618000_3825000# diff_3618000_3825000# diff_94000_5193000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3604 diff_94000_5193000# diff_2569000_3911000# diff_2569000_3911000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3605 diff_82000_3097000# diff_93000_3550000# diff_3447000_3516000# GND efet w=67500 l=12500
+ ad=0 pd=0 as=0 ps=0 
M3606 diff_3646000_3520000# diff_790000_4021000# diff_3443000_3166000# GND efet w=148000 l=11000
+ ad=1.036e+09 pd=310000 as=-1.46897e+09 ps=578000 
M3607 diff_82000_3097000# diff_3568000_3529000# diff_3531000_3484000# GND efet w=83500 l=10500
+ ad=0 pd=0 as=1.615e+09 ps=272000 
M3608 diff_3443000_3166000# diff_3443000_3166000# diff_94000_5193000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3609 diff_82000_3097000# diff_3653000_3514000# diff_3646000_3520000# GND efet w=148000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3610 diff_3487000_4661000# diff_71000_4514000# diff_3701000_3517000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.55e+08 ps=96000 
M3611 diff_82000_3097000# diff_3886000_4603000# diff_3980000_4516000# GND efet w=45500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3612 diff_82000_3097000# diff_3013000_3474000# diff_3980000_4516000# GND efet w=44000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3613 diff_4127000_4461000# diff_3956000_4961000# diff_82000_3097000# GND efet w=151500 l=11500
+ ad=-1.12797e+09 pd=650000 as=0 ps=0 
M3614 diff_4176000_4456000# diff_4016000_4961000# diff_82000_3097000# GND efet w=137000 l=11000
+ ad=-8.09967e+08 pd=744000 as=0 ps=0 
M3615 diff_82000_3097000# diff_4046000_4929000# diff_4176000_4456000# GND efet w=136000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3616 diff_4124000_2819000# diff_4074000_4961000# diff_82000_3097000# GND efet w=69000 l=12000
+ ad=6.42033e+08 pd=852000 as=0 ps=0 
M3617 diff_82000_3097000# diff_4322000_4961000# diff_4381000_4592000# GND efet w=61500 l=10500
+ ad=0 pd=0 as=1.854e+09 ps=352000 
M3618 diff_82000_3097000# diff_4292000_4961000# diff_4381000_4592000# GND efet w=44000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3619 diff_82000_3097000# diff_3986000_4961000# diff_4127000_4461000# GND efet w=142500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3620 diff_4176000_4456000# diff_3986000_4961000# diff_82000_3097000# GND efet w=150500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3621 diff_4067000_4316000# diff_3898000_4961000# diff_82000_3097000# GND efet w=88500 l=10500
+ ad=9.69e+08 pd=222000 as=0 ps=0 
M3622 diff_3980000_4516000# diff_529000_4371000# diff_4067000_4316000# GND efet w=87000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3623 diff_3940000_3885000# diff_790000_4021000# diff_2970000_4655000# GND efet w=132000 l=10000
+ ad=9.24e+08 pd=278000 as=-7.63967e+08 ps=638000 
M3624 diff_82000_3097000# diff_3780000_4961000# diff_3940000_3885000# GND efet w=132000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3625 diff_3908000_4368000# diff_3943000_3771000# diff_82000_3097000# GND efet w=47500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3626 diff_2970000_4655000# diff_2970000_4655000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3627 diff_3908000_4368000# diff_3908000_4368000# diff_94000_5193000# GND efet w=14000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M3628 diff_3943000_3771000# diff_71000_4514000# diff_2970000_4655000# GND efet w=15000 l=13000
+ ad=2.35e+08 pd=88000 as=0 ps=0 
M3629 diff_82000_3097000# diff_2859000_4569000# diff_2350000_3073000# GND efet w=207000 l=11000
+ ad=0 pd=0 as=-4.56967e+08 ps=644000 
M3630 diff_3792000_3499000# diff_3682000_4961000# diff_82000_3097000# GND efet w=145000 l=11000
+ ad=1.328e+09 pd=310000 as=0 ps=0 
M3631 diff_82000_3097000# diff_3121000_3079000# diff_2940000_2819000# GND efet w=66000 l=10000
+ ad=0 pd=0 as=1.522e+09 ps=380000 
M3632 diff_3049000_2819000# diff_3112000_3385000# diff_82000_3097000# GND efet w=81500 l=9500
+ ad=-2.04997e+09 pd=472000 as=0 ps=0 
M3633 diff_3232000_3141000# diff_529000_4371000# diff_3013000_2819000# GND efet w=133000 l=11000
+ ad=9.31e+08 pd=280000 as=1.24065e+08 ps=1.45e+06 
M3634 diff_82000_3097000# diff_511000_4351000# diff_3232000_3141000# GND efet w=133000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3635 diff_3283000_3143000# diff_3271000_3282000# diff_82000_3097000# GND efet w=131000 l=9000
+ ad=1.048e+09 pd=278000 as=0 ps=0 
M3636 diff_3013000_2819000# diff_518000_3031000# diff_3283000_3143000# GND efet w=131000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3637 diff_82000_3097000# diff_3173000_4961000# diff_3186000_3100000# GND efet w=146500 l=10500
+ ad=0 pd=0 as=1.688e+09 ps=428000 
M3638 diff_3186000_3100000# diff_905000_3225000# diff_3013000_2819000# GND efet w=142000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3639 diff_94000_5193000# diff_2601000_2819000# diff_2601000_2819000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3640 diff_3060000_3051000# diff_3060000_3051000# diff_94000_5193000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M3641 diff_2940000_2819000# diff_2940000_2819000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3642 diff_2631000_2819000# diff_2631000_2819000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3643 diff_94000_5193000# diff_2910000_2819000# diff_2910000_2819000# GND efet w=16000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3644 diff_3049000_2819000# diff_3049000_2819000# diff_94000_5193000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3645 diff_2631000_2819000# diff_71000_4514000# diff_2631000_2776000# GND efet w=22500 l=15500
+ ad=0 pd=0 as=9.95e+08 ps=162000 
M3646 diff_2601000_2819000# diff_71000_4514000# diff_2580000_2776000# GND efet w=21000 l=15000
+ ad=0 pd=0 as=1.004e+09 ps=162000 
M3647 diff_2677000_3054000# diff_71000_4514000# diff_2683000_2776000# GND efet w=21000 l=15000
+ ad=0 pd=0 as=9.92e+08 ps=162000 
M3648 diff_2734000_2819000# diff_71000_4514000# diff_2734000_2776000# GND efet w=21000 l=15000
+ ad=0 pd=0 as=9.92e+08 ps=162000 
M3649 diff_3013000_2819000# diff_168000_4544000# diff_82000_3097000# GND efet w=66000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3650 diff_3531000_3484000# diff_3531000_3484000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3651 diff_3550000_3278000# diff_93000_3550000# diff_82000_3097000# GND efet w=64000 l=9000
+ ad=-2.22967e+08 pd=818000 as=0 ps=0 
M3652 diff_82000_3097000# diff_3701000_3517000# diff_3550000_3278000# GND efet w=80500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3653 diff_3550000_3278000# diff_3550000_3278000# diff_94000_5193000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3654 diff_3550000_3278000# diff_67000_5287000# diff_3516000_3178000# GND efet w=15000 l=16000
+ ad=0 pd=0 as=3.09e+08 ps=104000 
M3655 diff_3013000_2819000# diff_3013000_2819000# diff_94000_5193000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3656 diff_3356000_3023000# diff_596000_3012000# diff_2837000_2819000# GND efet w=132000 l=10000
+ ad=1.03e+09 pd=278000 as=-1.21297e+09 ps=608000 
M3657 diff_82000_3097000# diff_3364000_3032000# diff_3356000_3023000# GND efet w=132500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M3658 diff_82000_3097000# diff_1603000_3122000# diff_3364000_3032000# GND efet w=79500 l=10500
+ ad=0 pd=0 as=-2.11497e+09 ps=374000 
M3659 diff_2837000_2819000# diff_2837000_2819000# diff_94000_5193000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M3660 diff_3364000_3032000# diff_3364000_3032000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3661 diff_2807000_2819000# diff_71000_4514000# diff_2787000_2776000# GND efet w=22000 l=15000
+ ad=0 pd=0 as=9.95e+08 ps=162000 
M3662 diff_2837000_2819000# diff_71000_4514000# diff_2837000_2776000# GND efet w=22000 l=15000
+ ad=0 pd=0 as=9.95e+08 ps=162000 
M3663 diff_2940000_2819000# diff_71000_4514000# diff_2940000_2776000# GND efet w=22500 l=15500
+ ad=0 pd=0 as=1.006e+09 ps=162000 
M3664 diff_2910000_2819000# diff_71000_4514000# diff_2890000_2776000# GND efet w=21000 l=15000
+ ad=0 pd=0 as=9.78e+08 ps=160000 
M3665 diff_3013000_2819000# diff_71000_4514000# diff_2993000_2776000# GND efet w=21000 l=15000
+ ad=0 pd=0 as=9.67e+08 ps=160000 
M3666 diff_3049000_2819000# diff_71000_4514000# diff_3046000_2782000# GND efet w=22000 l=15000
+ ad=0 pd=0 as=1.05e+09 ps=188000 
M3667 diff_2837000_2819000# diff_3106000_2804000# diff_3114000_2776000# GND efet w=21000 l=15000
+ ad=0 pd=0 as=1.003e+09 ps=162000 
M3668 diff_3187000_2819000# diff_3106000_2804000# diff_3167000_2776000# GND efet w=21000 l=15000
+ ad=5.60327e+07 pd=838000 as=9.67e+08 ps=160000 
M3669 diff_2464000_2760000# diff_2444000_2729000# diff_2444000_2729000# GND efet w=27000 l=10000
+ ad=4.85e+08 pd=94000 as=-1.72793e+09 ps=1.052e+06 
M3670 diff_2447000_2716000# diff_2447000_2716000# diff_2464000_2760000# GND efet w=20000 l=11000
+ ad=-1.00967e+08 pd=910000 as=0 ps=0 
M3671 diff_2444000_2729000# diff_2447000_2716000# diff_2441000_2691000# GND efet w=449000 l=11000
+ ad=0 pd=0 as=-2.11993e+09 ps=934000 
M3672 diff_2441000_2691000# diff_1439000_785000# diff_2248000_788000# GND efet w=216000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3673 diff_1851000_2289000# diff_1836000_1363000# diff_1833000_2289000# GND efet w=104000 l=12000
+ ad=1.055e+09 pd=226000 as=8.75e+08 ps=220000 
M3674 diff_1892000_2366000# diff_1891000_2340000# diff_1869000_2209000# GND efet w=14000 l=23000
+ ad=5.22e+08 pd=94000 as=-1.39397e+09 ps=500000 
M3675 diff_1931000_2307000# diff_1891000_2340000# diff_1869000_2209000# GND efet w=15000 l=81000
+ ad=5.9e+08 pd=138000 as=0 ps=0 
M3676 diff_2511000_2555000# diff_71000_4514000# diff_2447000_2716000# GND efet w=219500 l=10500
+ ad=-8.79967e+08 pd=522000 as=0 ps=0 
M3677 diff_1965000_2374000# diff_1891000_2340000# diff_1943000_2273000# GND efet w=15000 l=34000
+ ad=4.91e+08 pd=90000 as=1.183e+09 ps=208000 
M3678 diff_1869000_2209000# diff_1857000_1018000# diff_1850000_2209000# GND efet w=107500 l=12500
+ ad=0 pd=0 as=9.06e+08 ps=228000 
M3679 diff_1996000_2221000# diff_1996000_2221000# diff_2009000_2371000# GND efet w=14000 l=23000
+ ad=1.687e+09 pd=364000 as=4.7e+08 ps=88000 
M3680 diff_1889000_2181000# diff_1880000_2202000# diff_1869000_2209000# GND efet w=200500 l=9500
+ ad=-1.03093e+09 pd=788000 as=0 ps=0 
M3681 diff_1943000_2273000# diff_1931000_2307000# diff_1889000_2181000# GND efet w=63000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3682 diff_1996000_2221000# diff_1982000_1350000# diff_1981000_2297000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=3.96e+08 ps=80000 
M3683 diff_2103000_2359000# diff_1439000_785000# diff_2049000_2210000# GND efet w=24000 l=15000
+ ad=1.2e+08 pd=58000 as=3.7e+08 ps=108000 
M3684 diff_2123000_2359000# diff_2108000_871000# diff_2103000_2359000# GND efet w=24000 l=14500
+ ad=-1.37297e+09 pd=426000 as=0 ps=0 
M3685 diff_2015000_2221000# diff_2003000_996000# diff_1996000_2221000# GND efet w=122000 l=12000
+ ad=1.35e+09 pd=220000 as=0 ps=0 
M3686 diff_1869000_2161000# diff_1857000_1018000# diff_1850000_2129000# GND efet w=108000 l=12000
+ ad=-1.41497e+09 pd=494000 as=9.91e+08 ps=230000 
M3687 diff_1889000_2181000# diff_1880000_2170000# diff_1869000_2161000# GND efet w=199500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3688 diff_1851000_2073000# diff_1836000_1363000# diff_1833000_2037000# GND efet w=105000 l=12000
+ ad=1.07e+09 pd=228000 as=8.68e+08 ps=222000 
M3689 diff_1943000_2100000# diff_1931000_2081000# diff_1889000_2181000# GND efet w=64000 l=10000
+ ad=1.219e+09 pd=204000 as=0 ps=0 
M3690 diff_2052000_2279000# diff_2049000_2210000# diff_2035000_2184000# GND efet w=187500 l=10500
+ ad=1.26e+09 pd=306000 as=3.00033e+08 ps=858000 
M3691 diff_2015000_2139000# diff_2003000_996000# diff_1996000_2115000# GND efet w=118500 l=12500
+ ad=1.249e+09 pd=212000 as=1.787e+09 ps=362000 
M3692 diff_2052000_2101000# diff_2049000_2146000# diff_2035000_2184000# GND efet w=185500 l=10500
+ ad=1.262e+09 pd=306000 as=0 ps=0 
M3693 diff_1851000_1912000# diff_1836000_1363000# diff_1833000_1912000# GND efet w=104000 l=12000
+ ad=1.109e+09 pd=226000 as=8.14e+08 ps=220000 
M3694 diff_1996000_2115000# diff_1982000_1350000# diff_1981000_2078000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=3.78e+08 ps=78000 
M3695 diff_1869000_2161000# diff_1891000_1964000# diff_1892000_1989000# GND efet w=15500 l=24500
+ ad=0 pd=0 as=9.42e+08 ps=136000 
M3696 diff_1931000_2081000# diff_1891000_1964000# diff_1869000_2161000# GND efet w=14500 l=81500
+ ad=5.44e+08 pd=136000 as=0 ps=0 
M3697 diff_1943000_2100000# diff_1891000_1964000# diff_1965000_1997000# GND efet w=14000 l=34000
+ ad=0 pd=0 as=5.62e+08 ps=98000 
M3698 diff_1892000_1989000# diff_1891000_1964000# diff_1869000_1832000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=-1.32197e+09 ps=500000 
M3699 diff_1931000_1930000# diff_1891000_1964000# diff_1869000_1832000# GND efet w=15000 l=81000
+ ad=5.87e+08 pd=138000 as=0 ps=0 
M3700 diff_1965000_1997000# diff_1891000_1964000# diff_1943000_1896000# GND efet w=15000 l=34000
+ ad=0 pd=0 as=1.188e+09 ps=208000 
M3701 diff_1869000_1832000# diff_1857000_1018000# diff_1850000_1832000# GND efet w=108000 l=12000
+ ad=0 pd=0 as=9.54e+08 ps=230000 
M3702 diff_1996000_2115000# diff_1996000_2115000# diff_2009000_1994000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=8.13e+08 ps=122000 
M3703 diff_1996000_1844000# diff_1996000_1844000# diff_2009000_1994000# GND efet w=14500 l=24500
+ ad=1.703e+09 pd=364000 as=0 ps=0 
M3704 diff_1996000_1844000# diff_1982000_1350000# diff_1981000_1921000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=3.78e+08 ps=78000 
M3705 diff_2123000_2359000# diff_2129000_2349000# diff_2136000_2333000# GND efet w=68000 l=9000
+ ad=0 pd=0 as=1.716e+09 ps=374000 
M3706 diff_2197000_2356000# diff_2123000_2359000# diff_2123000_2359000# GND efet w=13000 l=23000
+ ad=1.324e+09 pd=160000 as=0 ps=0 
M3707 diff_2197000_2356000# diff_2183000_2247000# diff_2183000_2247000# GND efet w=14000 l=21000
+ ad=0 pd=0 as=1.63e+09 ps=340000 
M3708 diff_2533000_2491000# diff_2528000_2776000# diff_2511000_2555000# GND efet w=246000 l=10000
+ ad=4.10327e+07 pd=886000 as=0 ps=0 
M3709 diff_2562000_2748000# diff_2533000_2491000# diff_2533000_2491000# GND efet w=19000 l=10000
+ ad=4.18e+08 pd=82000 as=0 ps=0 
M3710 diff_2582000_2724000# diff_2582000_2724000# diff_2562000_2748000# GND efet w=19000 l=10000
+ ad=-4.39673e+07 pd=882000 as=0 ps=0 
M3711 diff_2562000_2537000# diff_2552000_2526000# diff_2533000_2491000# GND efet w=205500 l=10500
+ ad=-2.20967e+08 pd=442000 as=0 ps=0 
M3712 diff_2582000_2724000# diff_2552000_2526000# diff_2562000_2537000# GND efet w=206000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3713 diff_2615000_2552000# diff_2580000_2776000# diff_2582000_2724000# GND efet w=246000 l=10000
+ ad=2.70327e+07 pd=522000 as=0 ps=0 
M3714 diff_2637000_2491000# diff_2631000_2776000# diff_2615000_2552000# GND efet w=246500 l=10500
+ ad=-6.49673e+07 pd=882000 as=0 ps=0 
M3715 diff_2665000_2748000# diff_2637000_2491000# diff_2637000_2491000# GND efet w=19000 l=9000
+ ad=4.37e+08 pd=84000 as=0 ps=0 
M3716 diff_2640000_933000# diff_2640000_933000# diff_2665000_2748000# GND efet w=19000 l=10000
+ ad=-1.84967e+08 pd=882000 as=0 ps=0 
M3717 diff_2666000_2536000# diff_2655000_2527000# diff_2637000_2491000# GND efet w=205500 l=10500
+ ad=-3.90967e+08 pd=440000 as=0 ps=0 
M3718 diff_2640000_933000# diff_2655000_2527000# diff_2666000_2536000# GND efet w=205000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3719 diff_2718000_2552000# diff_2683000_2776000# diff_2640000_933000# GND efet w=246500 l=10500
+ ad=-3.29673e+07 pd=522000 as=0 ps=0 
M3720 diff_2712000_821000# diff_2734000_2776000# diff_2718000_2552000# GND efet w=246500 l=10500
+ ad=-1.28967e+08 pd=878000 as=0 ps=0 
M3721 diff_2769000_2748000# diff_2712000_821000# diff_2712000_821000# GND efet w=19000 l=10000
+ ad=4.18e+08 pd=82000 as=0 ps=0 
M3722 diff_2776000_764000# diff_2776000_764000# diff_2769000_2748000# GND efet w=19000 l=10000
+ ad=8.94033e+08 pd=978000 as=0 ps=0 
M3723 diff_2769000_2536000# diff_2759000_2526000# diff_2712000_821000# GND efet w=205000 l=10000
+ ad=-2.18967e+08 pd=442000 as=0 ps=0 
M3724 diff_2776000_764000# diff_2759000_2526000# diff_2769000_2536000# GND efet w=205500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3725 diff_2821000_2553000# diff_2787000_2776000# diff_2776000_764000# GND efet w=246000 l=11000
+ ad=-5.79673e+07 pd=522000 as=0 ps=0 
M3726 diff_2842000_1949000# diff_2837000_2776000# diff_2821000_2553000# GND efet w=246500 l=10500
+ ad=8.00327e+07 pd=884000 as=0 ps=0 
M3727 diff_2872000_2748000# diff_2842000_1949000# diff_2842000_1949000# GND efet w=19000 l=10000
+ ad=4.18e+08 pd=82000 as=0 ps=0 
M3728 diff_2892000_2724000# diff_2892000_2724000# diff_2872000_2748000# GND efet w=19000 l=10000
+ ad=2.31033e+08 pd=894000 as=0 ps=0 
M3729 diff_2872000_2536000# diff_2862000_2526000# diff_2842000_1949000# GND efet w=205000 l=10000
+ ad=-1.92967e+08 pd=442000 as=0 ps=0 
M3730 diff_2892000_2724000# diff_2862000_2526000# diff_2872000_2536000# GND efet w=205000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3731 diff_2924000_2553000# diff_2890000_2776000# diff_2892000_2724000# GND efet w=247000 l=10000
+ ad=1.53033e+08 pd=524000 as=0 ps=0 
M3732 diff_2938000_823000# diff_2940000_2776000# diff_2924000_2553000# GND efet w=247000 l=10000
+ ad=-1.54967e+08 pd=860000 as=0 ps=0 
M3733 diff_2975000_2748000# diff_2938000_823000# diff_2938000_823000# GND efet w=19000 l=10000
+ ad=4.37e+08 pd=84000 as=0 ps=0 
M3734 diff_2995000_2724000# diff_2995000_2724000# diff_2975000_2748000# GND efet w=19000 l=9000
+ ad=9.80327e+07 pd=892000 as=0 ps=0 
M3735 diff_2975000_2537000# diff_2965000_2526000# diff_2938000_823000# GND efet w=205500 l=10500
+ ad=-2.22967e+08 pd=442000 as=0 ps=0 
M3736 diff_2995000_2724000# diff_2965000_2526000# diff_2975000_2537000# GND efet w=205500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3737 diff_3027000_2553000# diff_2993000_2776000# diff_2995000_2724000# GND efet w=246500 l=10500
+ ad=-6.60967e+08 pd=522000 as=0 ps=0 
M3738 diff_3064000_2758000# diff_3042000_2722000# diff_3042000_2722000# GND efet w=15000 l=13000
+ ad=3.15e+08 pd=72000 as=-1.60967e+08 ps=690000 
M3739 diff_3119000_2491000# diff_3114000_2776000# diff_3098000_2440000# GND efet w=246000 l=10000
+ ad=-9.19673e+07 pd=892000 as=7.45033e+08 ps=698000 
M3740 diff_3149000_2748000# diff_3119000_2491000# diff_3119000_2491000# GND efet w=20000 l=10000
+ ad=4.4e+08 pd=84000 as=0 ps=0 
M3741 diff_3170000_2724000# diff_3170000_2724000# diff_3149000_2748000# GND efet w=20000 l=10000
+ ad=1.50033e+08 pd=864000 as=0 ps=0 
M3742 diff_3149000_2536000# diff_3139000_2526000# diff_3119000_2491000# GND efet w=204500 l=10500
+ ad=-2.33967e+08 pd=440000 as=0 ps=0 
M3743 diff_2292000_2348000# diff_2280000_2194000# diff_2280000_2194000# GND efet w=15000 l=23000
+ ad=1.919e+09 pd=236000 as=1.415e+09 ps=316000 
M3744 diff_2292000_2348000# diff_2248000_788000# diff_2291000_2206000# GND efet w=15000 l=11000
+ ad=0 pd=0 as=1.643e+09 ps=310000 
M3745 diff_2136000_2333000# diff_2126000_2298000# diff_2121000_2103000# GND efet w=127500 l=10500
+ ad=0 pd=0 as=9.84065e+08 ps=1.432e+06 
M3746 diff_2123000_2359000# diff_2129000_2349000# diff_2136000_2333000# GND efet w=74500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3747 diff_2121000_2103000# diff_2183000_2247000# diff_2123000_2359000# GND efet w=59000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3748 diff_2183000_2247000# diff_2206000_2293000# diff_2121000_2103000# GND efet w=66000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3749 diff_2121000_2103000# diff_2232000_2217000# diff_2183000_2247000# GND efet w=74000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3750 diff_2136000_2051000# diff_2126000_2081000# diff_2121000_2103000# GND efet w=131000 l=10000
+ ad=1.786e+09 pd=374000 as=0 ps=0 
M3751 diff_2123000_2013000# diff_2129000_2042000# diff_2136000_2051000# GND efet w=78000 l=10000
+ ad=-1.25097e+09 pd=458000 as=0 ps=0 
M3752 diff_2136000_2051000# diff_2129000_2042000# diff_2123000_2013000# GND efet w=64500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3753 diff_2121000_2103000# diff_2183000_2055000# diff_2123000_2013000# GND efet w=58000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3754 diff_2183000_2055000# diff_2129000_2042000# diff_2121000_2103000# GND efet w=66000 l=10000
+ ad=1.623e+09 pd=336000 as=0 ps=0 
M3755 diff_2121000_2103000# diff_2126000_2081000# diff_2183000_2055000# GND efet w=74000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3756 diff_2183000_2055000# diff_2183000_2055000# diff_2197000_1980000# GND efet w=14000 l=20000
+ ad=0 pd=0 as=-1.94797e+09 ps=226000 
M3757 diff_2103000_2013000# diff_1439000_785000# diff_2049000_2146000# GND efet w=23000 l=16000
+ ad=1.15e+08 pd=56000 as=3.62e+08 ps=98000 
M3758 diff_2123000_2013000# diff_2108000_871000# diff_2103000_2013000# GND efet w=23000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M3759 diff_2197000_1980000# diff_2123000_2013000# diff_2123000_2013000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3760 diff_2416000_2381000# diff_2409000_2357000# diff_2409000_2357000# GND efet w=14000 l=24000
+ ad=7.97e+08 pd=130000 as=2.107e+09 ps=434000 
M3761 diff_2475000_2369000# diff_2487000_2340000# diff_2487000_2340000# GND efet w=15000 l=24000
+ ad=8.84e+08 pd=144000 as=1.488e+09 ps=316000 
M3762 diff_2409000_2357000# diff_2392000_1580000# diff_2405000_2324000# GND efet w=152500 l=10500
+ ad=0 pd=0 as=1.295e+09 ps=306000 
M3763 diff_2291000_2206000# diff_2280000_2194000# diff_2126000_2081000# GND efet w=119500 l=11500
+ ad=0 pd=0 as=-1.48597e+09 ps=598000 
M3764 diff_2315000_2142000# diff_2319000_2260000# diff_2280000_2194000# GND efet w=57500 l=9500
+ ad=-7.54967e+08 pd=654000 as=0 ps=0 
M3765 diff_2303000_1745000# diff_2319000_2260000# diff_2315000_2142000# GND efet w=154000 l=11000
+ ad=4.30098e+08 pd=2.104e+06 as=0 ps=0 
M3766 diff_2405000_2324000# diff_2382000_2291000# diff_2385000_2111000# GND efet w=122000 l=11000
+ ad=0 pd=0 as=9.52033e+08 ps=508000 
M3767 diff_2292000_1877000# diff_2280000_2085000# diff_2126000_2081000# GND efet w=139000 l=11000
+ ad=-5.78967e+08 pd=650000 as=0 ps=0 
M3768 diff_2303000_1745000# diff_2319000_2129000# diff_2315000_2142000# GND efet w=156500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3769 diff_2315000_2142000# diff_2319000_2129000# diff_2280000_2085000# GND efet w=64000 l=10000
+ ad=0 pd=0 as=1.331e+09 ps=310000 
M3770 diff_2103000_1983000# diff_1439000_785000# diff_2049000_1833000# GND efet w=22000 l=16000
+ ad=1.1e+08 pd=54000 as=3.19e+08 ps=100000 
M3771 diff_2123000_1983000# diff_2108000_871000# diff_2103000_1983000# GND efet w=22000 l=15000
+ ad=-1.39797e+09 pd=426000 as=0 ps=0 
M3772 diff_2015000_1844000# diff_2003000_996000# diff_1996000_1844000# GND efet w=122000 l=12000
+ ad=1.351e+09 pd=220000 as=0 ps=0 
M3773 diff_1889000_1804000# diff_1880000_1825000# diff_1869000_1832000# GND efet w=200500 l=9500
+ ad=-1.01793e+09 pd=788000 as=0 ps=0 
M3774 diff_1943000_1896000# diff_1931000_1930000# diff_1889000_1804000# GND efet w=63000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3775 diff_1869000_1783000# diff_1857000_1018000# diff_1850000_1752000# GND efet w=108000 l=12000
+ ad=-1.43797e+09 pd=494000 as=1.007e+09 ps=230000 
M3776 diff_1889000_1804000# diff_1880000_1793000# diff_1869000_1783000# GND efet w=200500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3777 diff_1852000_1696000# diff_1836000_1363000# diff_1833000_1660000# GND efet w=103000 l=12000
+ ad=1.026e+09 pd=224000 as=9.08e+08 ps=220000 
M3778 diff_1943000_1723000# diff_1931000_1704000# diff_1889000_1804000# GND efet w=64000 l=10000
+ ad=1.218e+09 pd=204000 as=0 ps=0 
M3779 diff_2052000_1901000# diff_2049000_1833000# diff_2035000_1807000# GND efet w=186500 l=10500
+ ad=1.248e+09 pd=304000 as=2.75033e+08 ps=862000 
M3780 diff_2052000_1723000# diff_2049000_1769000# diff_2035000_1807000# GND efet w=187500 l=10500
+ ad=1.276e+09 pd=306000 as=0 ps=0 
M3781 diff_2015000_1762000# diff_2003000_996000# diff_1996000_1738000# GND efet w=119000 l=12000
+ ad=1.26e+09 pd=214000 as=1.764e+09 ps=362000 
M3782 diff_1851000_1534000# diff_1836000_1363000# diff_1833000_1534000# GND efet w=105000 l=12000
+ ad=1.128e+09 pd=228000 as=8.19e+08 ps=222000 
M3783 diff_1996000_1738000# diff_1982000_1350000# diff_1981000_1701000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=3.74e+08 ps=78000 
M3784 diff_1869000_1783000# diff_1891000_1587000# diff_1892000_1612000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=9.58e+08 ps=138000 
M3785 diff_1931000_1704000# diff_1891000_1587000# diff_1869000_1783000# GND efet w=14500 l=82500
+ ad=5.29e+08 pd=132000 as=0 ps=0 
M3786 diff_1943000_1723000# diff_1891000_1587000# diff_1965000_1620000# GND efet w=14000 l=34000
+ ad=0 pd=0 as=5.62e+08 ps=98000 
M3787 diff_1892000_1612000# diff_1891000_1587000# diff_1869000_1455000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=-1.32197e+09 ps=500000 
M3788 diff_1931000_1553000# diff_1891000_1587000# diff_1869000_1455000# GND efet w=15000 l=80000
+ ad=5.85e+08 pd=138000 as=0 ps=0 
M3789 diff_1965000_1620000# diff_1891000_1587000# diff_1943000_1520000# GND efet w=15000 l=34000
+ ad=0 pd=0 as=1.14e+09 ps=206000 
M3790 diff_1869000_1455000# diff_1857000_1018000# diff_1850000_1455000# GND efet w=107500 l=12500
+ ad=0 pd=0 as=8.89e+08 ps=228000 
M3791 diff_1996000_1738000# diff_1996000_1738000# diff_2009000_1617000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=8.13e+08 ps=122000 
M3792 diff_1996000_1467000# diff_1996000_1467000# diff_2009000_1617000# GND efet w=14500 l=23500
+ ad=1.719e+09 pd=366000 as=0 ps=0 
M3793 diff_1996000_1467000# diff_1982000_1350000# diff_1981000_1544000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=3.57e+08 ps=76000 
M3794 diff_2197000_1980000# diff_2123000_1983000# diff_2123000_1983000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3795 diff_2126000_2081000# diff_2248000_788000# diff_2272000_2002000# GND efet w=14000 l=11000
+ ad=0 pd=0 as=4.73e+08 ps=94000 
M3796 diff_2461000_2209000# diff_2392000_2433000# diff_2409000_2357000# GND efet w=153000 l=10000
+ ad=1.446e+09 pd=328000 as=0 ps=0 
M3797 diff_816000_2341000# diff_2591000_970000# diff_2549000_2332000# GND efet w=89500 l=10500
+ ad=0 pd=0 as=1.45003e+09 ps=534000 
M3798 diff_2480000_2122000# diff_2470000_2204000# diff_2461000_2209000# GND efet w=125500 l=9500
+ ad=-6.32967e+08 pd=588000 as=0 ps=0 
M3799 diff_2487000_2340000# diff_2470000_2204000# diff_2480000_2122000# GND efet w=60000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3800 diff_2549000_2332000# diff_2533000_2232000# diff_2533000_2232000# GND efet w=13000 l=17000
+ ad=0 pd=0 as=1.635e+09 ps=342000 
M3801 diff_94000_5193000# diff_94000_5193000# diff_2673000_2206000# GND efet w=13500 l=33500
+ ad=0 pd=0 as=9.95e+08 ps=188000 
M3802 diff_2684000_2216000# diff_94000_5193000# diff_2652000_2298000# GND efet w=14000 l=76000
+ ad=-3.50967e+08 pd=728000 as=5.3e+08 ps=198000 
M3803 diff_94000_5193000# diff_94000_5193000# diff_2684000_2216000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3804 diff_2652000_2298000# diff_2640000_933000# diff_816000_2341000# GND efet w=23000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M3805 diff_2652000_2298000# diff_2652000_2298000# diff_2652000_2298000# GND efet w=1500 l=3500
+ ad=0 pd=0 as=0 ps=0 
M3806 diff_2554000_2126000# diff_2544000_2207000# diff_2533000_2232000# GND efet w=86000 l=10000
+ ad=-1.75097e+09 pd=358000 as=0 ps=0 
M3807 diff_2533000_2232000# diff_2447000_2716000# diff_2470000_2204000# GND efet w=22000 l=15000
+ ad=0 pd=0 as=3.37e+08 ps=100000 
M3808 diff_2280000_2085000# diff_2280000_2085000# diff_2339000_1998000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=4.92e+08 ps=92000 
M3809 diff_2292000_1877000# diff_2248000_788000# diff_2272000_2002000# GND efet w=12000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3810 diff_2123000_1983000# diff_2129000_1971000# diff_2136000_1956000# GND efet w=67500 l=9500
+ ad=0 pd=0 as=1.703e+09 ps=372000 
M3811 diff_2197000_1980000# diff_2183000_1870000# diff_2183000_1870000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=1.641e+09 ps=338000 
M3812 diff_2136000_1956000# diff_2126000_1921000# diff_2121000_1727000# GND efet w=127500 l=10500
+ ad=0 pd=0 as=9.73065e+08 ps=1.43e+06 
M3813 diff_2123000_1983000# diff_2129000_1971000# diff_2136000_1956000# GND efet w=75000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3814 diff_2121000_1727000# diff_2183000_1870000# diff_2123000_1983000# GND efet w=58000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3815 diff_2183000_1870000# diff_2206000_1916000# diff_2121000_1727000# GND efet w=66000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3816 diff_2121000_1727000# diff_2232000_1840000# diff_2183000_1870000# GND efet w=74000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3817 diff_2136000_1674000# diff_2126000_1704000# diff_2121000_1727000# GND efet w=131000 l=10000
+ ad=1.79e+09 pd=374000 as=0 ps=0 
M3818 diff_2123000_1636000# diff_2129000_1665000# diff_2136000_1674000# GND efet w=77500 l=10500
+ ad=-1.26897e+09 pd=456000 as=0 ps=0 
M3819 diff_2136000_1674000# diff_2129000_1665000# diff_2123000_1636000# GND efet w=64500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3820 diff_2121000_1727000# diff_2183000_1678000# diff_2123000_1636000# GND efet w=59000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3821 diff_2183000_1678000# diff_2129000_1665000# diff_2121000_1727000# GND efet w=66000 l=10000
+ ad=1.636e+09 pd=334000 as=0 ps=0 
M3822 diff_2121000_1727000# diff_2126000_1704000# diff_2183000_1678000# GND efet w=73000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3823 diff_2280000_1865000# diff_2280000_1865000# diff_2339000_1998000# GND efet w=14500 l=22500
+ ad=1.53e+09 pd=322000 as=0 ps=0 
M3824 diff_2292000_1877000# diff_2280000_1865000# diff_2126000_1704000# GND efet w=119000 l=12000
+ ad=0 pd=0 as=-4.95967e+08 ps=606000 
M3825 diff_2406000_2068000# diff_2129000_2042000# diff_2385000_2111000# GND efet w=117500 l=10500
+ ad=1.282e+09 pd=296000 as=0 ps=0 
M3826 diff_2319000_2129000# diff_2392000_1580000# diff_2406000_2068000# GND efet w=148500 l=10500
+ ad=2.109e+09 pd=422000 as=0 ps=0 
M3827 diff_2461000_2102000# diff_2392000_2433000# diff_2319000_2129000# GND efet w=152000 l=10000
+ ad=1.442e+09 pd=326000 as=0 ps=0 
M3828 diff_2480000_2122000# diff_2470000_2111000# diff_2461000_2102000# GND efet w=125500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3829 diff_2549000_2332000# diff_2591000_970000# diff_2544000_2207000# GND efet w=87500 l=10500
+ ad=0 pd=0 as=-1.69593e+09 ps=1.348e+06 
M3830 diff_847000_2341000# diff_2591000_970000# diff_2549000_2332000# GND efet w=73000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3831 diff_2673000_2206000# diff_2652000_2298000# diff_2655000_2158000# GND efet w=65000 l=10000
+ ad=0 pd=0 as=1.25103e+09 ps=882000 
M3832 diff_2830000_2241000# diff_94000_5193000# diff_94000_5193000# GND efet w=13000 l=24000
+ ad=-1.33967e+08 pd=732000 as=0 ps=0 
M3833 diff_2914000_2317000# diff_94000_5193000# diff_2830000_2241000# GND efet w=14000 l=74000
+ ad=1.39e+09 pd=316000 as=0 ps=0 
M3834 diff_94000_5193000# diff_94000_5193000# diff_2875000_2204000# GND efet w=14000 l=32000
+ ad=0 pd=0 as=9.3e+08 ps=180000 
M3835 diff_3080000_2440000# diff_3064000_2691000# diff_3042000_2722000# GND efet w=246000 l=10000
+ ad=1.799e+09 pd=516000 as=0 ps=0 
M3836 diff_3098000_2440000# diff_3046000_2782000# diff_3080000_2440000# GND efet w=250500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3837 diff_3170000_2724000# diff_3139000_2526000# diff_3149000_2536000# GND efet w=204000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3838 diff_3201000_2552000# diff_3167000_2776000# diff_3170000_2724000# GND efet w=247500 l=10500
+ ad=1.31033e+08 pd=522000 as=0 ps=0 
M3839 diff_3302000_2723000# diff_3255000_1458000# diff_3255000_1458000# GND efet w=14000 l=16000
+ ad=1.011e+09 pd=144000 as=-7.70967e+08 ps=646000 
M3840 diff_3302000_2723000# diff_3282000_1425000# diff_3282000_1425000# GND efet w=15000 l=18000
+ ad=0 pd=0 as=-1.80897e+09 ps=520000 
M3841 diff_3282000_1425000# diff_3282000_1425000# diff_3282000_1425000# GND efet w=2000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3842 diff_3255000_1458000# diff_3253000_2508000# diff_3236000_2514000# GND efet w=104000 l=11000
+ ad=0 pd=0 as=1.768e+09 ps=242000 
M3843 diff_3488000_3125000# diff_2848000_2985000# diff_82000_3097000# GND efet w=131000 l=11000
+ ad=9.17e+08 pd=276000 as=0 ps=0 
M3844 diff_3432000_2819000# diff_530000_4621000# diff_3488000_3125000# GND efet w=131000 l=11000
+ ad=-1.24997e+09 pd=652000 as=0 ps=0 
M3845 diff_82000_3097000# diff_3516000_3178000# diff_3432000_2819000# GND efet w=77500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3846 diff_82000_3097000# diff_3516000_3069000# diff_3432000_2819000# GND efet w=66000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3847 diff_3187000_2819000# diff_3187000_2819000# diff_94000_5193000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3848 diff_3187000_2819000# diff_790000_4021000# diff_3792000_3499000# GND efet w=145500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3849 diff_82000_3097000# diff_2771000_3401000# diff_3187000_2819000# GND efet w=66000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3850 diff_4127000_4461000# diff_1000000_4393000# diff_4135000_4236000# GND efet w=141000 l=11000
+ ad=0 pd=0 as=2.068e+09 ps=418000 
M3851 diff_4124000_2819000# diff_790000_4021000# diff_4176000_4456000# GND efet w=132000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3852 diff_4248000_4332000# diff_4104000_4961000# diff_4124000_2819000# GND efet w=133000 l=11000
+ ad=9.31e+08 pd=280000 as=0 ps=0 
M3853 diff_82000_3097000# diff_945000_3262000# diff_4248000_4332000# GND efet w=133000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3854 diff_4381000_4592000# diff_4381000_4592000# diff_94000_5193000# GND efet w=14000 l=40000
+ ad=0 pd=0 as=0 ps=0 
M3855 diff_82000_3097000# diff_4380000_4961000# diff_4466000_4515000# GND efet w=44000 l=10000
+ ad=0 pd=0 as=8.46e+08 ps=212000 
M3856 diff_4317000_4211000# diff_4318000_4838000# diff_82000_3097000# GND efet w=79000 l=11000
+ ad=-3.91935e+08 pd=1.644e+06 as=0 ps=0 
M3857 diff_4124000_2819000# diff_4124000_2819000# diff_94000_5193000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3858 diff_4466000_4515000# diff_4466000_4515000# diff_94000_5193000# GND efet w=15000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M3859 diff_82000_3097000# diff_4558000_4961000# diff_4646000_4720000# GND efet w=42000 l=11000
+ ad=0 pd=0 as=-1.89697e+09 ps=434000 
M3860 diff_4646000_4720000# diff_4586000_4961000# diff_82000_3097000# GND efet w=46000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3861 diff_4646000_4720000# diff_4646000_4720000# diff_94000_5193000# GND efet w=14000 l=40000
+ ad=0 pd=0 as=0 ps=0 
M3862 diff_82000_3097000# diff_4616000_4961000# diff_4693000_4600000# GND efet w=46000 l=10000
+ ad=0 pd=0 as=1.802e+09 ps=412000 
M3863 diff_4693000_4600000# diff_4734000_4961000# diff_82000_3097000# GND efet w=51500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3864 diff_4317000_4211000# diff_4350000_4961000# diff_82000_3097000# GND efet w=67000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3865 diff_82000_3097000# diff_4381000_4592000# diff_4317000_4211000# GND efet w=63000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3866 diff_4469000_4299000# diff_4350000_4961000# diff_82000_3097000# GND efet w=44000 l=10000
+ ad=2.20327e+07 pd=846000 as=0 ps=0 
M3867 diff_82000_3097000# diff_4466000_4515000# diff_4469000_4299000# GND efet w=43000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3868 diff_4525000_4434000# diff_1000000_4393000# diff_82000_3097000# GND efet w=91000 l=10000
+ ad=6.71e+08 pd=196000 as=0 ps=0 
M3869 diff_94000_5193000# diff_4135000_4236000# diff_4135000_4236000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3870 diff_4170000_3958000# diff_71000_4514000# diff_4144000_3668000# GND efet w=15000 l=14000
+ ad=3.04e+08 pd=108000 as=-6.30967e+08 ps=704000 
M3871 diff_82000_3097000# diff_3928000_4961000# diff_4213000_3932000# GND efet w=45000 l=11000
+ ad=0 pd=0 as=-9.05967e+08 ps=586000 
M3872 diff_4144000_3668000# diff_3665000_4068000# diff_82000_3097000# GND efet w=42000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3873 diff_3187000_2819000# diff_71000_4514000# diff_3620000_3187000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=5.74e+08 ps=148000 
M3874 diff_3603000_3006000# diff_67000_5287000# diff_3578000_3163000# GND efet w=14000 l=14000
+ ad=1.867e+09 pd=344000 as=2.44e+08 ps=104000 
M3875 diff_3516000_3069000# diff_3443000_3166000# diff_82000_3097000# GND efet w=66000 l=10000
+ ad=1.419e+09 pd=282000 as=0 ps=0 
M3876 diff_82000_3097000# diff_3578000_3163000# diff_3505000_2819000# GND efet w=82000 l=10000
+ ad=0 pd=0 as=-1.19497e+09 ps=566000 
M3877 diff_3432000_2819000# diff_3432000_2819000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3878 diff_3516000_3069000# diff_3516000_3069000# diff_94000_5193000# GND efet w=15000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M3879 diff_82000_3097000# diff_3620000_3187000# diff_3603000_3006000# GND efet w=66000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3880 diff_3603000_3006000# diff_3603000_3006000# diff_94000_5193000# GND efet w=15000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M3881 diff_3818000_3048000# diff_3712000_4961000# diff_82000_3097000# GND efet w=82000 l=11000
+ ad=1.452e+09 pd=312000 as=0 ps=0 
M3882 diff_82000_3097000# diff_3665000_4068000# diff_3818000_3048000# GND efet w=80500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3883 diff_82000_3097000# diff_4170000_3958000# diff_4162000_3766000# GND efet w=55500 l=10500
+ ad=0 pd=0 as=2.12e+09 ps=458000 
M3884 diff_4219000_3817000# diff_4188000_3787000# diff_82000_3097000# GND efet w=87000 l=11000
+ ad=8.55e+08 pd=216000 as=0 ps=0 
M3885 diff_4213000_3932000# diff_4135000_4236000# diff_4219000_3817000# GND efet w=87000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3886 diff_4188000_3787000# diff_67000_5287000# diff_4162000_3766000# GND efet w=14000 l=14000
+ ad=2.45e+08 pd=86000 as=0 ps=0 
M3887 diff_4162000_3766000# diff_4162000_3766000# diff_94000_5193000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M3888 diff_4213000_3932000# diff_4213000_3932000# diff_94000_5193000# GND efet w=14000 l=40000
+ ad=0 pd=0 as=0 ps=0 
M3889 diff_94000_5193000# diff_4144000_3668000# diff_4144000_3668000# GND efet w=13000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M3890 diff_4045000_3494000# diff_790000_4021000# diff_3608000_2819000# GND efet w=136000 l=11000
+ ad=1.027e+09 pd=286000 as=-1.42397e+09 ps=638000 
M3891 diff_82000_3097000# diff_3810000_4961000# diff_4045000_3494000# GND efet w=136500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3892 diff_3638000_2819000# diff_1196000_3118000# diff_82000_3097000# GND efet w=67000 l=10000
+ ad=-5.40967e+08 pd=602000 as=0 ps=0 
M3893 diff_82000_3097000# diff_1603000_3122000# diff_3535000_2819000# GND efet w=79500 l=9500
+ ad=0 pd=0 as=1.7e+09 ps=392000 
M3894 diff_3638000_2819000# diff_1603000_3122000# diff_82000_3097000# GND efet w=80000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3895 diff_82000_3097000# diff_530000_4621000# diff_3638000_2819000# GND efet w=66000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3896 diff_3818000_3048000# diff_3818000_3048000# diff_94000_5193000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3897 diff_3550000_3278000# diff_67000_5287000# diff_3916000_3245000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=4.05e+08 ps=118000 
M3898 diff_3866000_3071000# diff_71000_4514000# diff_3608000_2819000# GND efet w=13000 l=13000
+ ad=5.19e+08 pd=148000 as=0 ps=0 
M3899 diff_82000_3097000# diff_2930000_4556000# diff_3711000_2819000# GND efet w=81500 l=10500
+ ad=0 pd=0 as=1.972e+09 ps=442000 
M3900 diff_3741000_2819000# diff_3818000_3048000# diff_82000_3097000# GND efet w=82000 l=11000
+ ad=-1.41097e+09 pd=556000 as=0 ps=0 
M3901 diff_94000_5193000# diff_3505000_2819000# diff_3505000_2819000# GND efet w=15000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3902 diff_3535000_2819000# diff_3535000_2819000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3903 diff_3638000_2819000# diff_3638000_2819000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3904 diff_3711000_2819000# diff_3711000_2819000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3905 diff_3741000_2819000# diff_3741000_2819000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3906 diff_3866000_2980000# diff_3866000_3071000# diff_82000_3097000# GND efet w=67000 l=10000
+ ad=1.948e+09 pd=386000 as=0 ps=0 
M3907 diff_3814000_2819000# diff_3916000_3245000# diff_82000_3097000# GND efet w=65000 l=10000
+ ad=-1.37397e+09 pd=590000 as=0 ps=0 
M3908 diff_4002000_3073000# diff_3701000_4747000# diff_82000_3097000# GND efet w=57000 l=11000
+ ad=1.175e+09 pd=278000 as=0 ps=0 
M3909 diff_82000_3097000# diff_3839000_4961000# diff_4002000_3073000# GND efet w=52000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3910 diff_4027000_3053000# diff_3980000_4516000# diff_82000_3097000# GND efet w=44000 l=10000
+ ad=-5.87967e+08 pd=764000 as=0 ps=0 
M3911 diff_82000_3097000# diff_4422000_4317000# diff_4317000_4211000# GND efet w=65000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3912 diff_82000_3097000# diff_4422000_4317000# diff_4469000_4299000# GND efet w=44000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3913 diff_4526000_4141000# diff_4410000_4961000# diff_4525000_4434000# GND efet w=91500 l=10500
+ ad=2.027e+09 pd=436000 as=0 ps=0 
M3914 diff_4693000_4600000# diff_4693000_4600000# diff_94000_5193000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M3915 diff_94000_5193000# diff_4526000_4141000# diff_4526000_4141000# GND efet w=14000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M3916 diff_4317000_4211000# diff_4317000_4211000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3917 diff_4469000_4299000# diff_4469000_4299000# diff_94000_5193000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M3918 diff_4375000_4011000# diff_3407000_4287000# diff_4317000_4211000# GND efet w=132000 l=11000
+ ad=7.92e+08 pd=276000 as=0 ps=0 
M3919 diff_82000_3097000# diff_4164000_4928000# diff_4375000_4011000# GND efet w=132000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3920 diff_82000_3097000# diff_4823000_4961000# diff_4787000_4475000# GND efet w=54500 l=10500
+ ad=0 pd=0 as=-1.90597e+09 ps=478000 
M3921 diff_82000_3097000# diff_4842000_4667000# diff_4787000_4475000# GND efet w=43000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3922 diff_5297000_4763000# diff_71000_4514000# diff_4901000_4753000# GND efet w=15000 l=14000
+ ad=3.54e+08 pd=76000 as=0 ps=0 
M3923 diff_6030000_4912000# diff_71000_4514000# diff_2350000_3073000# GND efet w=16000 l=14000
+ ad=2.52e+08 pd=102000 as=0 ps=0 
M3924 diff_5219000_4034000# diff_6030000_4912000# diff_82000_3097000# GND efet w=83500 l=10500
+ ad=1.525e+09 pd=288000 as=0 ps=0 
M3925 diff_94000_5193000# diff_5219000_4034000# diff_5219000_4034000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M3926 diff_6030000_4889000# diff_71000_4514000# diff_4317000_4211000# GND efet w=15000 l=14000
+ ad=3.39e+08 pd=110000 as=0 ps=0 
M3927 diff_82000_3097000# diff_6030000_4912000# diff_6077000_4886000# GND efet w=133000 l=10000
+ ad=0 pd=0 as=9.31e+08 ps=280000 
M3928 diff_6077000_4886000# diff_6030000_4889000# diff_5600000_3944000# GND efet w=133000 l=12000
+ ad=0 pd=0 as=-4.33935e+08 ps=1.142e+06 
M3929 diff_6030000_4850000# diff_71000_4514000# diff_4469000_4299000# GND efet w=16000 l=14000
+ ad=2.74e+08 pd=102000 as=0 ps=0 
M3930 diff_5600000_3944000# diff_6030000_4850000# diff_6077000_4837000# GND efet w=133000 l=10000
+ ad=0 pd=0 as=9.31e+08 ps=280000 
M3931 diff_82000_3097000# diff_5487000_4744000# diff_5412000_4657000# GND efet w=53500 l=9500
+ ad=0 pd=0 as=-1.32197e+09 ps=638000 
M3932 diff_4317000_4211000# diff_71000_4514000# diff_5487000_4744000# GND efet w=16000 l=14000
+ ad=0 pd=0 as=2.64e+08 ps=92000 
M3933 diff_4469000_4299000# diff_71000_4514000# diff_5488000_4717000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=6.99e+08 ps=150000 
M3934 diff_6077000_4837000# diff_5219000_4034000# diff_82000_3097000# GND efet w=133000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3935 diff_82000_3097000# diff_5488000_4717000# diff_5412000_4657000# GND efet w=54500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3936 diff_5642000_4716000# diff_67000_5287000# diff_5537000_2618000# GND efet w=15000 l=15000
+ ad=2.55e+08 pd=96000 as=1.33803e+09 ps=998000 
M3937 diff_82000_3097000# diff_5642000_4716000# diff_6077000_4788000# GND efet w=133000 l=11000
+ ad=0 pd=0 as=9.31e+08 ps=280000 
M3938 diff_6077000_4788000# diff_4926000_3399000# diff_5600000_3944000# GND efet w=133000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3939 diff_4921000_4668000# diff_71000_4514000# diff_3008000_4522000# GND efet w=14000 l=14000
+ ad=2.48e+08 pd=76000 as=0 ps=0 
M3940 diff_4926000_3399000# diff_4921000_4668000# diff_82000_3097000# GND efet w=165000 l=11000
+ ad=-1.92097e+09 pd=510000 as=0 ps=0 
M3941 diff_5600000_3944000# diff_4264000_3069000# diff_6077000_4739000# GND efet w=133000 l=10000
+ ad=0 pd=0 as=1.064e+09 ps=282000 
M3942 diff_5992000_4718000# diff_71000_4514000# diff_4919000_4771000# GND efet w=15000 l=15000
+ ad=4.3e+08 pd=108000 as=0 ps=0 
M3943 diff_6077000_4739000# diff_5992000_4718000# diff_82000_3097000# GND efet w=133000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3944 diff_5412000_4657000# diff_5412000_4657000# diff_94000_5193000# GND efet w=13500 l=38500
+ ad=0 pd=0 as=0 ps=0 
M3945 diff_4787000_4475000# diff_4787000_4475000# diff_94000_5193000# GND efet w=14000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M3946 diff_94000_5193000# diff_4926000_3399000# diff_4926000_3399000# GND efet w=15000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M3947 diff_82000_3097000# diff_4750000_4351000# diff_5126000_4638000# GND efet w=82000 l=11000
+ ad=0 pd=0 as=4.92e+08 ps=176000 
M3948 diff_5600000_3944000# diff_5336000_4601000# diff_82000_3097000# GND efet w=76500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3949 diff_5126000_4638000# diff_4693000_4600000# diff_5126000_4616000# GND efet w=82000 l=11000
+ ad=0 pd=0 as=2.04e+09 ps=352000 
M3950 diff_82000_3097000# diff_5475000_4642000# diff_5412000_4657000# GND efet w=49000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3951 diff_4919000_4771000# diff_71000_4514000# diff_5475000_4642000# GND efet w=16000 l=13000
+ ad=0 pd=0 as=2.42e+08 ps=78000 
M3952 diff_5412000_4657000# diff_5295000_4529000# diff_82000_3097000# GND efet w=45000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3953 diff_94000_5193000# diff_4805000_4500000# diff_4805000_4500000# GND efet w=15000 l=39000
+ ad=0 pd=0 as=-8.18967e+08 ps=668000 
M3954 diff_94000_5193000# diff_5126000_4616000# diff_5126000_4616000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M3955 diff_5336000_4601000# diff_5336000_4601000# diff_94000_5193000# GND efet w=13000 l=39000
+ ad=-1.78097e+09 pd=480000 as=0 ps=0 
M3956 diff_5412000_4657000# diff_4926000_3399000# diff_82000_3097000# GND efet w=47000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3957 diff_94000_5193000# diff_5600000_3944000# diff_5600000_3944000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3958 diff_5159000_4310000# diff_71000_4514000# diff_5126000_4616000# GND efet w=13000 l=13000
+ ad=4.11e+08 pd=92000 as=0 ps=0 
M3959 diff_5095000_4555000# diff_4693000_4600000# diff_82000_3097000# GND efet w=60000 l=11000
+ ad=1.769e+09 pd=322000 as=0 ps=0 
M3960 diff_5600000_3944000# diff_5412000_4657000# diff_6078000_4660000# GND efet w=132000 l=11000
+ ad=0 pd=0 as=9.24e+08 ps=278000 
M3961 diff_6078000_4660000# diff_6048000_4640000# diff_82000_3097000# GND efet w=132000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3962 diff_6048000_4640000# diff_71000_4514000# diff_3407000_4287000# GND efet w=13000 l=14000
+ ad=3.41e+08 pd=106000 as=-1.78397e+09 ps=514000 
M3963 diff_94000_5193000# diff_3407000_4287000# diff_3407000_4287000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M3964 diff_3407000_4287000# diff_5710000_4527000# diff_82000_3097000# GND efet w=118000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3965 diff_5095000_4555000# diff_5073000_4505000# diff_82000_3097000# GND efet w=44000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3966 diff_5230000_4553000# diff_71000_4514000# diff_5095000_4555000# GND efet w=14000 l=13000
+ ad=6.03e+08 pd=104000 as=0 ps=0 
M3967 diff_82000_3097000# diff_1000000_4393000# diff_5073000_4505000# GND efet w=66000 l=10000
+ ad=0 pd=0 as=1.442e+09 ps=264000 
M3968 diff_5336000_4568000# diff_5336000_4568000# diff_94000_5193000# GND efet w=12000 l=39000
+ ad=1.943e+09 pd=414000 as=0 ps=0 
M3969 diff_4750000_4351000# diff_4769000_4457000# diff_82000_3097000# GND efet w=72500 l=10500
+ ad=1.809e+09 pd=420000 as=0 ps=0 
M3970 diff_82000_3097000# diff_4422000_4317000# diff_4750000_4351000# GND efet w=81500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3971 diff_4805000_4500000# diff_4787000_4475000# diff_82000_3097000# GND efet w=46500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3972 diff_82000_3097000# diff_4422000_4317000# diff_4805000_4500000# GND efet w=45000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3973 diff_5095000_4555000# diff_5095000_4555000# diff_94000_5193000# GND efet w=14000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M3974 diff_82000_3097000# diff_5456000_4543000# diff_5336000_4601000# GND efet w=42000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3975 diff_5295000_4529000# diff_5295000_4529000# diff_94000_5193000# GND efet w=14000 l=38000
+ ad=1.346e+09 pd=216000 as=0 ps=0 
M3976 diff_94000_5193000# diff_4750000_4351000# diff_4750000_4351000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3977 diff_4375000_3895000# diff_4164000_4928000# diff_4357000_3757000# GND efet w=136500 l=10500
+ ad=9.52e+08 pd=286000 as=-1.71197e+09 ps=552000 
M3978 diff_82000_3097000# diff_790000_4021000# diff_4375000_3895000# GND efet w=136500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3979 diff_4420000_3821000# diff_790000_4021000# diff_82000_3097000# GND efet w=134500 l=10500
+ ad=9.41e+08 pd=282000 as=0 ps=0 
M3980 diff_4414000_3773000# diff_4427000_3812000# diff_4420000_3821000# GND efet w=134000 l=10000
+ ad=-9.20967e+08 pd=686000 as=0 ps=0 
M3981 diff_82000_3097000# diff_4192000_4961000# diff_4457000_3836000# GND efet w=142500 l=10500
+ ad=0 pd=0 as=-8.60967e+08 ps=748000 
M3982 diff_4457000_3836000# diff_4222000_4961000# diff_82000_3097000# GND efet w=148500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3983 diff_4461000_3007000# diff_4515000_3836000# diff_4457000_3836000# GND efet w=133000 l=10000
+ ad=-7.31967e+08 pd=704000 as=0 ps=0 
M3984 diff_82000_3097000# diff_1196000_3118000# diff_4515000_3836000# GND efet w=73000 l=10000
+ ad=0 pd=0 as=-6.33967e+08 ps=690000 
M3985 diff_94000_5193000# diff_4357000_3757000# diff_4357000_3757000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3986 diff_4414000_3773000# diff_4414000_3773000# diff_94000_5193000# GND efet w=15000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M3987 diff_94000_5193000# diff_4461000_3007000# diff_4461000_3007000# GND efet w=14500 l=24500
+ ad=0 pd=0 as=0 ps=0 
M3988 diff_4515000_3836000# diff_4515000_3836000# diff_94000_5193000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3989 diff_82000_3097000# diff_4213000_3932000# diff_4021000_2819000# GND efet w=74500 l=9500
+ ad=0 pd=0 as=1.74033e+08 ps=822000 
M3990 diff_82000_3097000# diff_3928000_4961000# diff_4027000_3053000# GND efet w=45000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3991 diff_4027000_3053000# diff_2967000_4961000# diff_82000_3097000# GND efet w=45000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3992 diff_3608000_2819000# diff_3608000_2819000# diff_94000_5193000# GND efet w=13000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3993 diff_4021000_2819000# diff_2937000_3466000# diff_82000_3097000# GND efet w=65000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3994 diff_4305000_3504000# diff_4134000_4961000# diff_4021000_2819000# GND efet w=133000 l=10000
+ ad=9.31e+08 pd=280000 as=0 ps=0 
M3995 diff_82000_3097000# diff_529000_4371000# diff_4305000_3504000# GND efet w=133000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3996 diff_4002000_3073000# diff_4002000_3073000# diff_94000_5193000# GND efet w=15000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M3997 diff_4027000_3053000# diff_4027000_3053000# diff_94000_5193000# GND efet w=15000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M3998 diff_4021000_2819000# diff_4021000_2819000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M3999 diff_3814000_2819000# diff_3905000_3048000# diff_82000_3097000# GND efet w=66000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4000 diff_82000_3097000# diff_1603000_3122000# diff_3814000_2819000# GND efet w=91000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4001 diff_3905000_3048000# diff_67000_5287000# diff_3866000_2980000# GND efet w=14000 l=13000
+ ad=2.94e+08 pd=82000 as=0 ps=0 
M4002 diff_3866000_2980000# diff_3866000_2980000# diff_94000_5193000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M4003 diff_3814000_2819000# diff_3814000_2819000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4004 diff_4296000_3177000# diff_4264000_3069000# diff_82000_3097000# GND efet w=71000 l=11000
+ ad=1.785e+09 pd=332000 as=0 ps=0 
M4005 diff_82000_3097000# diff_4002000_3073000# diff_3845000_2819000# GND efet w=69000 l=10000
+ ad=0 pd=0 as=-1.24497e+09 ps=600000 
M4006 diff_3948000_2819000# diff_4027000_3053000# diff_82000_3097000# GND efet w=81000 l=10000
+ ad=1.974e+09 pd=414000 as=0 ps=0 
M4007 diff_3948000_2819000# diff_3948000_2819000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4008 diff_3845000_2819000# diff_3845000_2819000# diff_94000_5193000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M4009 diff_3443000_3166000# diff_71000_4514000# diff_4094000_3084000# GND efet w=15000 l=13000
+ ad=0 pd=0 as=4.79e+08 ps=134000 
M4010 diff_4086000_3164000# diff_67000_5287000# diff_4067000_3123000# GND efet w=13000 l=14000
+ ad=5.85e+08 pd=126000 as=-1.80697e+09 ps=470000 
M4011 diff_82000_3097000# diff_4094000_3084000# diff_4067000_3123000# GND efet w=43000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4012 diff_4051000_2819000# diff_4086000_3164000# diff_82000_3097000# GND efet w=70000 l=10000
+ ad=-1.60497e+09 pd=562000 as=0 ps=0 
M4013 diff_4067000_3123000# diff_4067000_3123000# diff_94000_5193000# GND efet w=15000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M4014 diff_4155000_3009000# diff_2848000_2985000# diff_4051000_2819000# GND efet w=133000 l=10000
+ ad=1.264e+09 pd=320000 as=0 ps=0 
M4015 diff_82000_3097000# diff_529000_4371000# diff_4155000_3009000# GND efet w=152000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4016 diff_4051000_2819000# diff_4051000_2819000# diff_94000_5193000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4017 diff_4296000_3177000# diff_4296000_3177000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4018 diff_82000_3097000# diff_1936000_3037000# diff_4224000_2933000# GND efet w=81000 l=10000
+ ad=0 pd=0 as=-1.46097e+09 ps=480000 
M4019 diff_4307000_3184000# diff_4296000_3177000# diff_82000_3097000# GND efet w=116000 l=11000
+ ad=8.12e+08 pd=246000 as=0 ps=0 
M4020 diff_4261000_2986000# diff_3407000_4287000# diff_4307000_3184000# GND efet w=116500 l=10500
+ ad=5.33033e+08 pd=838000 as=0 ps=0 
M4021 diff_82000_3097000# diff_1096000_3118000# diff_4494000_3313000# GND efet w=84000 l=11000
+ ad=0 pd=0 as=-7.83967e+08 ps=676000 
M4022 diff_82000_3097000# diff_1000000_4393000# diff_4422000_4317000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=1.35e+09 ps=318000 
M4023 diff_94000_5193000# diff_5073000_4505000# diff_5073000_4505000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4024 diff_5023000_4456000# diff_71000_4514000# diff_4994000_4439000# GND efet w=14000 l=13000
+ ad=5.37e+08 pd=160000 as=1.302e+09 ps=290000 
M4025 diff_5336000_4568000# diff_71000_4514000# diff_5456000_4543000# GND efet w=14500 l=14500
+ ad=0 pd=0 as=2.52e+08 ps=90000 
M4026 diff_5600000_3944000# diff_67000_5287000# diff_5710000_4527000# GND efet w=16000 l=14000
+ ad=0 pd=0 as=2.96e+08 ps=108000 
M4027 diff_5336000_4568000# diff_5295000_4529000# diff_5390000_4497000# GND efet w=128000 l=11000
+ ad=0 pd=0 as=1.215e+09 ps=312000 
M4028 diff_5396000_4486000# diff_67000_5287000# diff_5537000_2618000# GND efet w=22000 l=15000
+ ad=5.55e+08 pd=152000 as=0 ps=0 
M4029 diff_82000_3097000# diff_5396000_4486000# diff_5390000_4497000# GND efet w=131500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4030 diff_5295000_4529000# diff_5023000_4456000# diff_82000_3097000# GND efet w=44000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4031 diff_6152000_4535000# diff_5097000_4893000# diff_82000_3097000# GND efet w=44000 l=10000
+ ad=1.977e+09 pd=394000 as=0 ps=0 
M4032 diff_6152000_4535000# diff_5979000_4396000# diff_82000_3097000# GND efet w=47000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4033 diff_94000_5193000# diff_6152000_4535000# diff_6152000_4535000# GND efet w=14000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M4034 diff_4181000_2527000# diff_5741000_4459000# diff_82000_3097000# GND efet w=82000 l=11000
+ ad=1.837e+09 pd=362000 as=0 ps=0 
M4035 diff_82000_3097000# diff_4926000_3399000# diff_5257000_4375000# GND efet w=45000 l=11000
+ ad=0 pd=0 as=-1.64297e+09 ps=462000 
M4036 diff_4994000_4439000# diff_4983000_4429000# diff_82000_3097000# GND efet w=61500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4037 diff_94000_5193000# diff_4994000_4439000# diff_4994000_4439000# GND efet w=14000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M4038 diff_5741000_4459000# diff_67000_5287000# diff_5388000_4407000# GND efet w=14000 l=13000
+ ad=3.01e+08 pd=96000 as=1.94107e+09 ps=1.874e+06 
M4039 diff_6222000_4301000# diff_5979000_4396000# diff_82000_3097000# GND efet w=43000 l=11000
+ ad=1.511e+09 pd=250000 as=0 ps=0 
M4040 diff_94000_5193000# diff_6222000_4301000# diff_6222000_4301000# GND efet w=14000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M4041 diff_82000_3097000# diff_4302000_2656000# diff_5948000_4451000# GND efet w=88000 l=11000
+ ad=0 pd=0 as=-1.99797e+09 ps=430000 
M4042 diff_82000_3097000# diff_4181000_2527000# diff_5948000_4451000# GND efet w=88000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4043 diff_5948000_4451000# diff_5825000_4380000# diff_5979000_4396000# GND efet w=90000 l=10000
+ ad=0 pd=0 as=1.772e+09 ps=338000 
M4044 diff_5055000_4360000# diff_67000_5287000# diff_4983000_4429000# GND efet w=16000 l=13000
+ ad=9.95e+08 pd=238000 as=2.78e+08 ps=78000 
M4045 diff_94000_5193000# diff_5055000_4360000# diff_5055000_4360000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M4046 diff_5388000_4407000# diff_5345000_4398000# diff_5388000_4390000# GND efet w=132000 l=9000
+ ad=0 pd=0 as=1.056e+09 ps=280000 
M4047 diff_5257000_4375000# diff_5257000_4375000# diff_94000_5193000# GND efet w=13000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M4048 diff_82000_3097000# diff_5560000_4417000# diff_5568000_4410000# GND efet w=131000 l=11000
+ ad=0 pd=0 as=9.17e+08 ps=276000 
M4049 diff_4181000_2527000# diff_71000_4514000# diff_5560000_4417000# GND efet w=15000 l=13000
+ ad=0 pd=0 as=2.28e+08 ps=88000 
M4050 diff_5568000_4410000# diff_5257000_4375000# diff_5388000_4407000# GND efet w=131000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4051 diff_82000_3097000# diff_5230000_4553000# diff_5257000_4375000# GND efet w=60000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4052 diff_5388000_4390000# diff_5230000_4553000# diff_82000_3097000# GND efet w=132000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4053 diff_94000_5193000# diff_5388000_4407000# diff_5388000_4407000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4054 diff_6186000_3964000# diff_6152000_4535000# diff_82000_3097000# GND efet w=50500 l=10500
+ ad=1.493e+09 pd=296000 as=0 ps=0 
M4055 diff_5979000_4396000# diff_5979000_4396000# diff_94000_5193000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M4056 diff_6186000_3964000# diff_6186000_3964000# diff_6186000_3964000# GND efet w=500 l=2500
+ ad=0 pd=0 as=0 ps=0 
M4057 diff_94000_5193000# diff_6186000_3964000# diff_6186000_3964000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M4058 diff_6186000_3964000# diff_5097000_4893000# diff_6145000_4382000# GND efet w=89000 l=10000
+ ad=0 pd=0 as=-1.92097e+09 ps=508000 
M4059 diff_4980000_4332000# diff_4980000_4332000# diff_4980000_4332000# GND efet w=500 l=3500
+ ad=2.25e+08 pd=78000 as=0 ps=0 
M4060 diff_5055000_4360000# diff_4980000_4332000# diff_82000_3097000# GND efet w=53000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4061 diff_4980000_4332000# diff_71000_4514000# diff_4414000_3773000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M4062 diff_5170000_4318000# diff_5159000_4310000# diff_82000_3097000# GND efet w=47000 l=11000
+ ad=8.52e+08 pd=180000 as=0 ps=0 
M4063 diff_94000_5193000# diff_5170000_4318000# diff_5170000_4318000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M4064 diff_5602000_4345000# diff_5297000_4763000# diff_82000_3097000# GND efet w=131000 l=10000
+ ad=1.048e+09 pd=278000 as=0 ps=0 
M4065 diff_5825000_4380000# diff_5825000_4380000# diff_94000_5193000# GND efet w=14000 l=38000
+ ad=9.11e+08 pd=244000 as=0 ps=0 
M4066 diff_6145000_4382000# diff_4240000_2639000# diff_82000_3097000# GND efet w=88000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4067 diff_6145000_4382000# diff_6222000_4301000# diff_82000_3097000# GND efet w=45000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4068 diff_6145000_4382000# diff_6222000_4301000# diff_82000_3097000# GND efet w=42000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4069 diff_82000_3097000# diff_5297000_4763000# diff_5257000_4375000# GND efet w=44000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4070 diff_5602000_4345000# diff_4264000_3069000# diff_5388000_4407000# GND efet w=131000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4071 diff_4422000_4317000# diff_4422000_4317000# diff_94000_5193000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M4072 diff_5056000_4274000# diff_71000_4514000# diff_4696000_3225000# GND efet w=15000 l=13000
+ ad=2.7e+08 pd=96000 as=4.97033e+08 ps=978000 
M4073 diff_94000_5193000# diff_5090000_4256000# diff_5090000_4256000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=1.681e+09 ps=332000 
M4074 diff_5257000_4375000# diff_5170000_4318000# diff_82000_3097000# GND efet w=44000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4075 diff_82000_3097000# diff_5056000_4274000# diff_5090000_4256000# GND efet w=66000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4076 diff_5388000_4407000# diff_4926000_3399000# diff_5602000_4299000# GND efet w=140500 l=11500
+ ad=0 pd=0 as=1.001e+09 ps=312000 
M4077 diff_5163000_4225000# diff_67000_5287000# diff_5090000_4256000# GND efet w=14000 l=13000
+ ad=5.44e+08 pd=136000 as=0 ps=0 
M4078 diff_5375000_4258000# diff_67000_5287000# diff_5375000_4231000# GND efet w=16000 l=14000
+ ad=5.02e+08 pd=116000 as=5.84e+08 ps=126000 
M4079 diff_5602000_4299000# diff_5375000_4258000# diff_82000_3097000# GND efet w=149000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4080 diff_5825000_4380000# diff_4181000_2527000# diff_6030000_4331000# GND efet w=88000 l=11000
+ ad=0 pd=0 as=7.04e+08 ps=192000 
M4081 diff_6030000_4331000# diff_4302000_2656000# diff_82000_3097000# GND efet w=88000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4082 diff_82000_3097000# diff_5067000_4961000# diff_5955000_4223000# GND efet w=45500 l=10500
+ ad=0 pd=0 as=7.71e+08 ps=166000 
M4083 diff_82000_3097000# diff_4240000_2639000# diff_6144000_4250000# GND efet w=44000 l=10000
+ ad=0 pd=0 as=-1.90397e+09 ps=438000 
M4084 diff_82000_3097000# diff_6222000_4301000# diff_6144000_4250000# GND efet w=43000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4085 diff_94000_5193000# diff_6144000_4250000# diff_6144000_4250000# GND efet w=15000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M4086 diff_5574000_4253000# diff_5170000_4318000# diff_82000_3097000# GND efet w=136000 l=10000
+ ad=1.023e+09 pd=288000 as=0 ps=0 
M4087 diff_5574000_4253000# diff_5566000_4242000# diff_5388000_4407000# GND efet w=137000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4088 diff_94000_5193000# diff_4181000_2527000# diff_4181000_2527000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4089 diff_5955000_4223000# diff_5955000_4223000# diff_94000_5193000# GND efet w=13000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M4090 diff_4716000_3890000# diff_790000_4021000# diff_4696000_3225000# GND efet w=145000 l=10000
+ ad=1.024e+09 pd=304000 as=0 ps=0 
M4091 diff_82000_3097000# diff_4498000_4961000# diff_4716000_3890000# GND efet w=145000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4092 diff_4526000_4141000# diff_71000_4514000# diff_5003000_4149000# GND efet w=14000 l=15000
+ ad=0 pd=0 as=2.15e+08 ps=76000 
M4093 diff_94000_5193000# diff_5027000_4157000# diff_5027000_4157000# GND efet w=14000 l=39000
+ ad=0 pd=0 as=1.357e+09 ps=272000 
M4094 diff_5027000_4157000# diff_5003000_4149000# diff_82000_3097000# GND efet w=44000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4095 diff_94000_5193000# diff_5113000_4072000# diff_94000_5193000# GND efet w=21500 l=19500
+ ad=0 pd=0 as=0 ps=0 
M4096 diff_5027000_4157000# diff_67000_5287000# diff_5018000_4115000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=4.75e+08 ps=120000 
M4097 diff_4779000_3876000# diff_4528000_4961000# diff_4761000_3820000# GND efet w=143000 l=10000
+ ad=1.112e+09 pd=300000 as=-1.71397e+09 ps=592000 
M4098 diff_82000_3097000# diff_4515000_3836000# diff_4779000_3876000# GND efet w=141500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4099 diff_82000_3097000# diff_5018000_4115000# diff_5028000_4063000# GND efet w=43000 l=11000
+ ad=0 pd=0 as=1.409e+09 ps=278000 
M4100 diff_94000_5193000# diff_5113000_4072000# diff_5113000_4072000# GND efet w=14000 l=39000
+ ad=0 pd=0 as=1.909e+09 ps=390000 
M4101 diff_5566000_4242000# diff_71000_4514000# diff_5673000_4155000# GND efet w=13000 l=14000
+ ad=1.91e+08 pd=66000 as=-1.49997e+09 ps=540000 
M4102 diff_94000_5193000# diff_5673000_4155000# diff_5673000_4155000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4103 diff_6157000_4261000# diff_6144000_4250000# diff_6157000_4244000# GND efet w=88000 l=11000
+ ad=-2.03497e+09 pd=386000 as=5.28e+08 ps=188000 
M4104 diff_94000_5193000# diff_6157000_4261000# diff_6157000_4261000# GND efet w=15000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M4105 diff_6157000_4244000# diff_5097000_4893000# diff_82000_3097000# GND efet w=88000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4106 diff_6157000_4261000# diff_6178000_4192000# diff_82000_3097000# GND efet w=44000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4107 diff_5673000_4155000# diff_5452000_4209000# diff_82000_3097000# GND efet w=69000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4108 diff_5673000_4155000# diff_5163000_4225000# diff_82000_3097000# GND efet w=69000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4109 diff_94000_5193000# diff_5028000_4063000# diff_5028000_4063000# GND efet w=14000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M4110 diff_5056000_4063000# diff_71000_4514000# diff_5028000_4063000# GND efet w=14000 l=13000
+ ad=2.45e+08 pd=96000 as=0 ps=0 
M4111 diff_5113000_4072000# diff_5056000_4063000# diff_82000_3097000# GND efet w=54000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4112 diff_6178000_4192000# diff_5097000_4893000# diff_82000_3097000# GND efet w=52500 l=10500
+ ad=1.765e+09 pd=364000 as=0 ps=0 
M4113 diff_82000_3097000# diff_6222000_4301000# diff_6178000_4192000# GND efet w=45000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4114 diff_82000_3097000# diff_5917000_4119000# diff_2119000_4000000# GND efet w=81500 l=10500
+ ad=0 pd=0 as=-2.36967e+08 ps=706000 
M4115 diff_5355000_4072000# diff_5330000_4061000# diff_5355000_4054000# GND efet w=145500 l=10500
+ ad=5.10065e+08 pd=1.71e+06 as=1.015e+09 ps=304000 
M4116 diff_5355000_4054000# diff_5219000_4034000# diff_5355000_4036000# GND efet w=145500 l=10500
+ ad=0 pd=0 as=9.68e+08 ps=304000 
M4117 diff_5355000_4036000# diff_5009000_3740000# diff_82000_3097000# GND efet w=144500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4118 diff_5611000_4009000# diff_5600000_3944000# diff_82000_3097000# GND efet w=120500 l=10500
+ ad=-1.02697e+09 pd=690000 as=0 ps=0 
M4119 diff_82000_3097000# diff_3407000_4287000# diff_5849000_3990000# GND efet w=44000 l=10000
+ ad=0 pd=0 as=-2.13197e+09 ps=444000 
M4120 diff_5849000_3990000# diff_5849000_3990000# diff_94000_5193000# GND efet w=14000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M4121 diff_5611000_4009000# diff_5370000_3653000# diff_82000_3097000# GND efet w=134000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4122 diff_4715000_3242000# diff_4646000_4720000# diff_82000_3097000# GND efet w=75000 l=10000
+ ad=-1.79897e+09 pd=596000 as=0 ps=0 
M4123 diff_82000_3097000# diff_4427000_3812000# diff_4715000_3242000# GND efet w=73500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4124 diff_4696000_3225000# diff_4696000_3225000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4125 diff_4761000_3820000# diff_4761000_3820000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4126 diff_4715000_3242000# diff_4715000_3242000# diff_94000_5193000# GND efet w=15000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4127 diff_82000_3097000# diff_1196000_3118000# diff_4715000_3242000# GND efet w=66000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4128 diff_82000_3097000# diff_3358000_4500000# diff_4813000_3334000# GND efet w=65000 l=11000
+ ad=0 pd=0 as=-1.51897e+09 ps=624000 
M4129 diff_82000_3097000# diff_1196000_3118000# diff_4813000_3334000# GND efet w=65000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4130 diff_4750000_4351000# diff_71000_4514000# diff_5060000_3958000# GND efet w=14000 l=13000
+ ad=0 pd=0 as=4.96e+08 ps=136000 
M4131 diff_82000_3097000# diff_5060000_3958000# diff_5273000_3954000# GND efet w=78500 l=10500
+ ad=0 pd=0 as=-1.20997e+09 ps=598000 
M4132 diff_5079000_3925000# diff_67000_5287000# diff_3550000_3278000# GND efet w=15000 l=14000
+ ad=5.36e+08 pd=156000 as=0 ps=0 
M4133 diff_5355000_4072000# diff_5330000_4061000# diff_5273000_3954000# GND efet w=163000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4134 diff_5068000_3913000# diff_71000_4514000# diff_4974000_3888000# GND efet w=14000 l=13000
+ ad=1.151e+09 pd=230000 as=3.94e+08 ps=116000 
M4135 diff_5068000_3913000# diff_5079000_3925000# diff_82000_3097000# GND efet w=47000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4136 diff_5273000_3954000# diff_5263000_3944000# diff_5262000_3934000# GND efet w=144500 l=9500
+ ad=0 pd=0 as=1.026e+09 ps=296000 
M4137 diff_5262000_3934000# diff_5113000_4072000# diff_82000_3097000# GND efet w=124000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4138 diff_82000_3097000# diff_4974000_3888000# diff_4972000_3873000# GND efet w=44000 l=12000
+ ad=0 pd=0 as=1.318e+09 ps=274000 
M4139 diff_94000_5193000# diff_5068000_3913000# diff_5068000_3913000# GND efet w=14000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M4140 diff_82000_3097000# diff_5113000_4072000# diff_5227000_3878000# GND efet w=43000 l=10000
+ ad=0 pd=0 as=5.10327e+07 ps=802000 
M4141 diff_4972000_3873000# diff_67000_5287000# diff_4972000_3833000# GND efet w=14000 l=13000
+ ad=0 pd=0 as=2.88e+08 ps=100000 
M4142 diff_94000_5193000# diff_4972000_3873000# diff_4972000_3873000# GND efet w=15000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M4143 diff_82000_3097000# diff_4926000_3399000# diff_5227000_3878000# GND efet w=51000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4144 diff_82000_3097000# diff_4972000_3833000# diff_4996000_3825000# GND efet w=46500 l=10500
+ ad=0 pd=0 as=1.228e+09 ps=254000 
M4145 diff_5345000_4398000# diff_5624000_3955000# diff_5611000_4009000# GND efet w=161000 l=10000
+ ad=-1.56397e+09 pd=444000 as=0 ps=0 
M4146 diff_94000_5193000# diff_5345000_4398000# diff_5345000_4398000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4147 diff_5849000_3990000# diff_3568000_3529000# diff_82000_3097000# GND efet w=44000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4148 diff_5849000_3990000# diff_4240000_2639000# diff_82000_3097000# GND efet w=43000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4149 diff_94000_5193000# diff_6178000_4192000# diff_6178000_4192000# GND efet w=13000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M4150 diff_5995000_3978000# diff_3568000_3529000# diff_82000_3097000# GND efet w=134000 l=10000
+ ad=1.31033e+08 pd=780000 as=0 ps=0 
M4151 diff_82000_3097000# diff_5849000_3990000# diff_5995000_3978000# GND efet w=133000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4152 diff_6197000_3984000# diff_6186000_3964000# diff_82000_3097000# GND efet w=89000 l=11000
+ ad=-1.61997e+09 pd=638000 as=0 ps=0 
M4153 diff_5917000_4119000# diff_5008000_4961000# diff_6197000_3984000# GND efet w=97500 l=10500
+ ad=-1.41597e+09 pd=566000 as=0 ps=0 
M4154 diff_94000_5193000# diff_5917000_4119000# diff_5917000_4119000# GND efet w=15000 l=35000
+ ad=0 pd=0 as=0 ps=0 
M4155 diff_5917000_4119000# diff_5955000_4223000# diff_82000_3097000# GND efet w=41000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4156 diff_82000_3097000# diff_5762000_4183000# diff_5917000_4119000# GND efet w=42000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4157 diff_6197000_3984000# diff_6157000_4261000# diff_5917000_4119000# GND efet w=115000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4158 diff_82000_3097000# diff_5695000_3193000# diff_6197000_3984000# GND efet w=95000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4159 diff_82000_3097000# diff_5695000_3193000# diff_6197000_3984000# GND efet w=34000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4160 diff_5995000_3978000# diff_5987000_3968000# diff_2119000_4000000# GND efet w=157000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4161 diff_5624000_3955000# diff_5600000_3944000# diff_5624000_3937000# GND efet w=132000 l=11000
+ ad=-1.99797e+09 pd=464000 as=9.24e+08 ps=278000 
M4162 diff_2119000_4000000# diff_2119000_4000000# diff_94000_5193000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4163 diff_5624000_3937000# diff_5370000_3653000# diff_82000_3097000# GND efet w=132000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4164 diff_94000_5193000# diff_5624000_3955000# diff_5624000_3955000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4165 diff_82000_3097000# diff_5982000_3916000# diff_2119000_4000000# GND efet w=65000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4166 diff_82000_3097000# diff_6075000_3941000# diff_2119000_4000000# GND efet w=66000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4167 diff_5762000_4183000# diff_5762000_4183000# diff_94000_5193000# GND efet w=15000 l=39000
+ ad=1.024e+09 pd=218000 as=0 ps=0 
M4168 diff_4996000_3825000# diff_71000_4514000# diff_4993000_3786000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=2.69e+08 ps=110000 
M4169 diff_94000_5193000# diff_4996000_3825000# diff_4996000_3825000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M4170 diff_4628000_3379000# diff_1697000_2847000# diff_82000_3097000# GND efet w=213000 l=11000
+ ad=1.52e+09 pd=438000 as=0 ps=0 
M4171 diff_4477000_4816000# diff_3228000_4781000# diff_4628000_3379000# GND efet w=211500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4172 diff_82000_3097000# diff_4510000_3501000# diff_4494000_3313000# GND efet w=72000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4173 diff_4510000_3501000# diff_4318000_4838000# diff_82000_3097000# GND efet w=80000 l=11000
+ ad=1.404e+09 pd=316000 as=0 ps=0 
M4174 diff_82000_3097000# diff_4422000_4317000# diff_4510000_3501000# GND efet w=66000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4175 diff_4510000_3501000# diff_4510000_3501000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4176 diff_4494000_3313000# diff_4494000_3313000# diff_94000_5193000# GND efet w=15000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M4177 diff_4477000_4816000# diff_4477000_4816000# diff_94000_5193000# GND efet w=14000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M4178 diff_82000_3097000# diff_4264000_3069000# diff_4277000_3057000# GND efet w=109500 l=10500
+ ad=0 pd=0 as=1.074e+09 ps=278000 
M4179 diff_4261000_2986000# diff_4224000_2933000# diff_4277000_3057000# GND efet w=102000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4180 diff_4362000_2477000# diff_4261000_2986000# diff_82000_3097000# GND efet w=180000 l=10000
+ ad=-1.77197e+09 pd=490000 as=0 ps=0 
M4181 diff_4261000_2986000# diff_4261000_2986000# diff_94000_5193000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4182 diff_94000_5193000# diff_4224000_2933000# diff_4224000_2933000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4183 diff_82000_3097000# diff_3568000_3529000# diff_4362000_2477000# GND efet w=171000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4184 diff_4436000_3014000# diff_4357000_3757000# diff_82000_3097000# GND efet w=198000 l=10000
+ ad=1.584e+09 pd=412000 as=0 ps=0 
M4185 diff_4454000_3014000# diff_4414000_3773000# diff_4436000_3014000# GND efet w=198000 l=10000
+ ad=1.386e+09 pd=410000 as=0 ps=0 
M4186 diff_4461000_2970000# diff_4461000_3007000# diff_4454000_3014000# GND efet w=198000 l=11000
+ ad=-2.22967e+08 pd=634000 as=0 ps=0 
M4187 diff_4592000_3171000# diff_4477000_4816000# diff_82000_3097000# GND efet w=66000 l=11000
+ ad=2.90327e+07 pd=688000 as=0 ps=0 
M4188 diff_82000_3097000# diff_4468000_4961000# diff_4592000_3171000# GND efet w=65000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4189 diff_4813000_3334000# diff_4813000_3334000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4190 diff_94000_5193000# diff_5009000_3740000# diff_5009000_3740000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=9.38e+08 ps=218000 
M4191 diff_5227000_3878000# diff_5227000_3878000# diff_94000_5193000# GND efet w=15000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M4192 diff_82000_3097000# diff_5060000_3958000# diff_5227000_3878000# GND efet w=61000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4193 diff_5009000_3740000# diff_4993000_3786000# diff_82000_3097000# GND efet w=54000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4194 diff_94000_5193000# diff_127000_4096000# diff_127000_4096000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4195 diff_127000_4096000# diff_5047000_3692000# diff_5038000_3681000# GND efet w=50500 l=10500
+ ad=0 pd=0 as=1.861e+09 ps=418000 
M4196 diff_5038000_3681000# diff_5047000_3692000# diff_127000_4096000# GND efet w=81500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4197 diff_5263000_3944000# diff_71000_4514000# diff_4240000_2639000# GND efet w=14000 l=13000
+ ad=2.24e+08 pd=72000 as=-1.82797e+09 ps=470000 
M4198 diff_5762000_4183000# diff_5038000_4961000# diff_82000_3097000# GND efet w=43000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4199 diff_5982000_3916000# diff_5762000_4183000# diff_82000_3097000# GND efet w=51500 l=9500
+ ad=1.952e+09 pd=360000 as=0 ps=0 
M4200 diff_94000_5193000# diff_5982000_3916000# diff_5982000_3916000# GND efet w=15000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M4201 diff_5500000_3808000# diff_4926000_3399000# diff_82000_3097000# GND efet w=104000 l=10000
+ ad=7.28e+08 pd=222000 as=0 ps=0 
M4202 diff_5500000_3808000# diff_5320000_3743000# diff_5355000_4072000# GND efet w=104500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4203 diff_94000_5193000# diff_5355000_4072000# diff_5355000_4072000# GND efet w=15000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M4204 diff_5355000_4072000# diff_5227000_3878000# diff_5500000_3769000# GND efet w=106000 l=11000
+ ad=0 pd=0 as=7.49e+08 ps=226000 
M4205 diff_5355000_4072000# diff_67000_5287000# diff_5677000_3739000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=3.3e+08 ps=74000 
M4206 diff_5227000_3878000# diff_5009000_3740000# diff_82000_3097000# GND efet w=51000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4207 diff_5982000_3916000# diff_5067000_4961000# diff_82000_3097000# GND efet w=58000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4208 diff_6160000_3829000# diff_6150000_3838000# diff_5982000_3916000# GND efet w=91000 l=11000
+ ad=1.966e+09 pd=432000 as=0 ps=0 
M4209 diff_6160000_3829000# diff_3568000_3529000# diff_82000_3097000# GND efet w=91000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4210 diff_6160000_3829000# diff_6154000_3763000# diff_82000_3097000# GND efet w=88000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4211 diff_5500000_3769000# diff_5490000_3759000# diff_82000_3097000# GND efet w=105500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4212 diff_3568000_3529000# diff_3568000_3529000# diff_94000_5193000# GND efet w=15000 l=25000
+ ad=9e+08 pd=140000 as=0 ps=0 
M4213 diff_82000_3097000# diff_5042000_3670000# diff_5038000_3681000# GND efet w=138000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4214 diff_5042000_3670000# diff_4926000_3399000# diff_82000_3097000# GND efet w=43000 l=11000
+ ad=9.27e+08 pd=192000 as=0 ps=0 
M4215 diff_94000_5193000# diff_5042000_3670000# diff_5042000_3670000# GND efet w=13000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M4216 diff_4240000_2639000# diff_71000_4514000# diff_5490000_3759000# GND efet w=14000 l=13000
+ ad=0 pd=0 as=2.65e+08 ps=92000 
M4217 diff_5320000_3743000# diff_67000_5287000# diff_4199000_2721000# GND efet w=14000 l=14000
+ ad=3.13e+08 pd=72000 as=1.458e+09 ps=324000 
M4218 diff_94000_5193000# diff_4240000_2639000# diff_4240000_2639000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4219 diff_4240000_2639000# diff_5677000_3739000# diff_82000_3097000# GND efet w=67000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4220 diff_82000_3097000# diff_5097000_4893000# diff_3568000_3529000# GND efet w=70500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4221 diff_5294000_3705000# diff_67000_5287000# diff_4305000_1753000# GND efet w=14000 l=13000
+ ad=3.52e+08 pd=106000 as=1.74033e+08 ps=806000 
M4222 diff_82000_3097000# diff_5294000_3705000# diff_5396000_3689000# GND efet w=99000 l=10000
+ ad=0 pd=0 as=7.14e+08 ps=212000 
M4223 diff_5396000_3689000# diff_4926000_3399000# diff_5396000_3663000# GND efet w=98500 l=10500
+ ad=0 pd=0 as=3.61033e+08 ps=838000 
M4224 diff_82000_3097000# diff_5008000_4961000# diff_6154000_3781000# GND efet w=88000 l=10000
+ ad=0 pd=0 as=6.16e+08 ps=190000 
M4225 diff_6154000_3781000# diff_4302000_2656000# diff_6154000_3763000# GND efet w=88000 l=10000
+ ad=0 pd=0 as=1.697e+09 ps=334000 
M4226 diff_6154000_3763000# diff_6145000_3753000# diff_82000_3097000# GND efet w=47000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4227 diff_94000_5193000# diff_6154000_3763000# diff_6154000_3763000# GND efet w=15000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M4228 diff_6145000_3753000# diff_4302000_2656000# diff_82000_3097000# GND efet w=46000 l=10000
+ ad=2.012e+09 pd=416000 as=0 ps=0 
M4229 diff_6145000_3753000# diff_5008000_4961000# diff_82000_3097000# GND efet w=42000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4230 diff_4870000_3350000# diff_4926000_3399000# diff_82000_3097000# GND efet w=49500 l=10500
+ ad=-1.75297e+09 pd=410000 as=0 ps=0 
M4231 diff_82000_3097000# diff_5021000_3614000# diff_4870000_3350000# GND efet w=45000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4232 diff_5021000_3614000# diff_71000_4514000# diff_4805000_4500000# GND efet w=14000 l=14000
+ ad=4.57e+08 pd=136000 as=0 ps=0 
M4233 diff_94000_5193000# diff_5227000_3586000# diff_5227000_3586000# GND efet w=15000 l=38000
+ ad=0 pd=0 as=-6.84967e+08 ps=766000 
M4234 diff_94000_5193000# diff_5396000_3663000# diff_5396000_3663000# GND efet w=17000 l=43000
+ ad=0 pd=0 as=0 ps=0 
M4235 diff_94000_5193000# diff_6145000_3753000# diff_6145000_3753000# GND efet w=13000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M4236 diff_5396000_3663000# diff_5370000_3653000# diff_5396000_3645000# GND efet w=99000 l=10000
+ ad=0 pd=0 as=6.91e+08 ps=210000 
M4237 diff_5396000_3663000# diff_5227000_3586000# diff_5512000_3640000# GND efet w=57000 l=10000
+ ad=0 pd=0 as=1.159e+09 ps=296000 
M4238 diff_5396000_3645000# diff_5060000_3958000# diff_82000_3097000# GND efet w=98500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4239 diff_5227000_3586000# diff_5060000_3958000# diff_82000_3097000# GND efet w=44000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4240 diff_5512000_3640000# diff_5503000_3629000# diff_82000_3097000# GND efet w=117500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4241 diff_5396000_3663000# diff_67000_5287000# diff_5659000_3639000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=3.72e+08 ps=114000 
M4242 diff_5396000_3663000# diff_5227000_3586000# diff_5512000_3640000# GND efet w=28000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4243 diff_4302000_2656000# diff_5659000_3639000# diff_82000_3097000# GND efet w=64000 l=10000
+ ad=2.033e+09 pd=414000 as=0 ps=0 
M4244 diff_82000_3097000# diff_4926000_3399000# diff_5227000_3586000# GND efet w=43000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4245 diff_6150000_3838000# diff_3568000_3529000# diff_6184000_3576000# GND efet w=146000 l=11000
+ ad=-1.96697e+09 pd=458000 as=-2.02097e+09 ps=472000 
M4246 diff_94000_5193000# diff_4870000_3350000# diff_4870000_3350000# GND efet w=14000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M4247 diff_4302000_2656000# diff_71000_4514000# diff_5503000_3629000# GND efet w=15000 l=13000
+ ad=0 pd=0 as=2.5e+08 ps=74000 
M4248 diff_94000_5193000# diff_4302000_2656000# diff_4302000_2656000# GND efet w=13000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4249 diff_6016000_3580000# diff_6016000_3580000# diff_94000_5193000# GND efet w=14000 l=37000
+ ad=1.722e+09 pd=342000 as=0 ps=0 
M4250 diff_82000_3097000# diff_5008000_4961000# diff_6184000_3601000# GND efet w=145500 l=10500
+ ad=0 pd=0 as=1.015e+09 ps=304000 
M4251 diff_82000_3097000# diff_4181000_2527000# diff_6016000_3580000# GND efet w=44000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4252 diff_6184000_3601000# diff_4181000_2527000# diff_6184000_3576000# GND efet w=145000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4253 diff_82000_3097000# diff_5008000_4961000# diff_6016000_3580000# GND efet w=43000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4254 diff_6184000_3576000# diff_6016000_3580000# diff_82000_3097000# GND efet w=73000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4255 diff_6150000_3838000# diff_6150000_3838000# diff_94000_5193000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M4256 diff_82000_3097000# diff_4926000_3399000# diff_5356000_3321000# GND efet w=45000 l=11000
+ ad=0 pd=0 as=-4.80967e+08 ps=678000 
M4257 diff_82000_3097000# diff_4926000_3399000# diff_5471000_3487000# GND efet w=96000 l=11000
+ ad=0 pd=0 as=5.76e+08 ps=204000 
M4258 diff_5471000_3487000# diff_5295000_3448000# diff_5047000_3692000# GND efet w=96000 l=11000
+ ad=0 pd=0 as=-1.47693e+09 ps=1.25e+06 
M4259 diff_6111000_3387000# diff_4240000_2639000# diff_6159000_3508000# GND efet w=89000 l=10000
+ ad=-6.77967e+08 pd=734000 as=5.34e+08 ps=190000 
M4260 diff_6159000_3508000# diff_5097000_4893000# diff_82000_3097000# GND efet w=89000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4261 diff_5295000_3448000# diff_67000_5287000# diff_816000_1587000# GND efet w=16000 l=13000
+ ad=2.56e+08 pd=106000 as=0 ps=0 
M4262 diff_5047000_3692000# diff_5431000_3450000# diff_5438000_3443000# GND efet w=99000 l=11000
+ ad=0 pd=0 as=6.93e+08 ps=212000 
M4263 diff_5047000_3692000# diff_67000_5287000# diff_5577000_3392000# GND efet w=15000 l=13000
+ ad=0 pd=0 as=3.86e+08 ps=84000 
M4264 diff_94000_5193000# diff_5047000_3692000# diff_5047000_3692000# GND efet w=14000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M4265 diff_82000_3097000# diff_3407000_4287000# diff_6159000_3458000# GND efet w=92500 l=10500
+ ad=0 pd=0 as=6.6e+08 ps=200000 
M4266 diff_4592000_3171000# diff_530000_4621000# diff_82000_3097000# GND efet w=69000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4267 diff_82000_3097000# diff_64000_4219000# diff_4592000_3171000# GND efet w=79500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4268 diff_4778000_3197000# diff_71000_4514000# diff_4696000_3225000# GND efet w=14000 l=13000
+ ad=5.95e+08 pd=154000 as=0 ps=0 
M4269 diff_3282000_2537000# diff_3272000_2527000# diff_3255000_1458000# GND efet w=125500 l=9500
+ ad=1.456e+09 pd=244000 as=0 ps=0 
M4270 diff_3282000_1425000# diff_3272000_2527000# diff_3282000_2537000# GND efet w=102000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4271 diff_3331000_2538000# diff_3320000_2526000# diff_3282000_1425000# GND efet w=128000 l=10000
+ ad=1.359e+09 pd=260000 as=0 ps=0 
M4272 diff_3432000_2819000# diff_71000_4514000# diff_3432000_2777000# GND efet w=22500 l=15500
+ ad=0 pd=0 as=9.94e+08 ps=158000 
M4273 diff_3400000_3460000# diff_71000_4514000# diff_3382000_2777000# GND efet w=21000 l=15000
+ ad=0 pd=0 as=9.57e+08 ps=156000 
M4274 diff_3505000_2819000# diff_71000_4514000# diff_3485000_2777000# GND efet w=21000 l=15000
+ ad=0 pd=0 as=9.57e+08 ps=156000 
M4275 diff_3535000_2819000# diff_71000_4514000# diff_3535000_2777000# GND efet w=22000 l=15000
+ ad=0 pd=0 as=9.84e+08 ps=158000 
M4276 diff_3608000_2819000# diff_71000_4514000# diff_3588000_2777000# GND efet w=21000 l=15000
+ ad=0 pd=0 as=9.67e+08 ps=156000 
M4277 diff_3638000_2819000# diff_71000_4514000# diff_3638000_2777000# GND efet w=21000 l=15000
+ ad=0 pd=0 as=9.82e+08 ps=158000 
M4278 diff_3711000_2819000# diff_71000_4514000# diff_3691000_2777000# GND efet w=21000 l=15000
+ ad=0 pd=0 as=9.57e+08 ps=156000 
M4279 diff_3741000_2819000# diff_71000_4514000# diff_3741000_2777000# GND efet w=21000 l=15000
+ ad=0 pd=0 as=9.82e+08 ps=158000 
M4280 diff_3845000_2819000# diff_71000_4514000# diff_3845000_2777000# GND efet w=21500 l=15500
+ ad=0 pd=0 as=9.57e+08 ps=156000 
M4281 diff_3814000_2819000# diff_71000_4514000# diff_3793000_2777000# GND efet w=21000 l=15000
+ ad=0 pd=0 as=9.91e+08 ps=158000 
M4282 diff_3666000_4700000# diff_71000_4514000# diff_3897000_2777000# GND efet w=22000 l=15000
+ ad=0 pd=0 as=9.94e+08 ps=158000 
M4283 diff_3948000_2819000# diff_71000_4514000# diff_3948000_2777000# GND efet w=21000 l=15000
+ ad=0 pd=0 as=9.81e+08 ps=158000 
M4284 diff_4021000_2819000# diff_71000_4514000# diff_4000000_2777000# GND efet w=21000 l=15000
+ ad=0 pd=0 as=9.82e+08 ps=158000 
M4285 diff_4051000_2819000# diff_71000_4514000# diff_4051000_2777000# GND efet w=21000 l=15000
+ ad=0 pd=0 as=9.82e+08 ps=158000 
M4286 diff_4124000_2819000# diff_71000_4514000# diff_4103000_2777000# GND efet w=21000 l=15000
+ ad=0 pd=0 as=9.81e+08 ps=158000 
M4287 diff_3353000_2408000# diff_3353000_2408000# diff_3367000_2749000# GND efet w=19000 l=10000
+ ad=9.90033e+08 pd=1.13e+06 as=3.61e+08 ps=76000 
M4288 diff_3353000_2408000# diff_3364000_2491000# diff_3367000_2515000# GND efet w=205000 l=10000
+ ad=0 pd=0 as=-6.32967e+08 ps=436000 
M4289 diff_3416000_2552000# diff_3382000_2777000# diff_3353000_2408000# GND efet w=246500 l=10500
+ ad=4.90327e+07 pd=522000 as=0 ps=0 
M4290 diff_3438000_2491000# diff_3432000_2777000# diff_3416000_2552000# GND efet w=246000 l=10000
+ ad=4.85033e+08 pd=900000 as=0 ps=0 
M4291 diff_3467000_2748000# diff_3438000_2491000# diff_3438000_2491000# GND efet w=20000 l=10000
+ ad=4.4e+08 pd=84000 as=0 ps=0 
M4292 diff_3488000_2724000# diff_3488000_2724000# diff_3467000_2748000# GND efet w=20000 l=10000
+ ad=3.98033e+08 pd=898000 as=0 ps=0 
M4293 diff_3467000_2537000# diff_3457000_2526000# diff_3438000_2491000# GND efet w=205500 l=10500
+ ad=-2.20967e+08 pd=442000 as=0 ps=0 
M4294 diff_2684000_2216000# diff_2673000_2206000# diff_2655000_2158000# GND efet w=220500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4295 diff_2544000_2207000# diff_2712000_821000# diff_2684000_2216000# GND efet w=105000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4296 diff_2533000_2142000# diff_2447000_2716000# diff_2470000_2111000# GND efet w=23000 l=14000
+ ad=1.647e+09 pd=340000 as=3.2e+08 ps=84000 
M4297 diff_2129000_2042000# diff_2470000_2111000# diff_2480000_2122000# GND efet w=60000 l=9000
+ ad=1.508e+09 pd=308000 as=0 ps=0 
M4298 diff_2554000_2126000# diff_2544000_2115000# diff_2533000_2142000# GND efet w=80500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4299 diff_2549000_1954000# diff_2591000_970000# diff_2544000_2115000# GND efet w=88500 l=10500
+ ad=-1.5939e+09 pd=918000 as=1.142e+09 ps=228000 
M4300 diff_2628000_2106000# diff_2591000_970000# diff_2549000_1954000# GND efet w=73000 l=11000
+ ad=1.007e+09 pd=184000 as=0 ps=0 
M4301 diff_816000_2341000# diff_2776000_764000# diff_2684000_2216000# GND efet w=109000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4302 diff_2830000_2241000# diff_2582000_2724000# diff_816000_2341000# GND efet w=88000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4303 diff_2914000_2317000# diff_2938000_823000# diff_816000_2341000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4304 diff_2914000_2317000# diff_2914000_2317000# diff_2914000_2317000# GND efet w=1500 l=12500
+ ad=0 pd=0 as=0 ps=0 
M4305 diff_2830000_2241000# diff_2842000_1949000# diff_847000_2341000# GND efet w=108500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M4306 diff_2684000_2154000# diff_2673000_2143000# diff_2655000_2158000# GND efet w=220500 l=10500
+ ad=-1.54897e+09 pd=488000 as=0 ps=0 
M4307 diff_2674000_2059000# diff_2652000_2076000# diff_2655000_2158000# GND efet w=68000 l=10000
+ ad=9.54e+08 pd=186000 as=0 ps=0 
M4308 diff_2759000_2135000# diff_2712000_821000# diff_2684000_2154000# GND efet w=105000 l=12000
+ ad=1.236e+09 pd=236000 as=0 ps=0 
M4309 diff_2533000_2142000# diff_2533000_2142000# diff_2549000_1954000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M4310 diff_2319000_2129000# diff_2319000_2129000# diff_2416000_2004000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=7.5e+08 ps=136000 
M4311 diff_2416000_2004000# diff_2409000_1980000# diff_2409000_1980000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=2.089e+09 ps=430000 
M4312 diff_2129000_2042000# diff_2129000_2042000# diff_2475000_1993000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=1.408e+09 ps=178000 
M4313 diff_2475000_1993000# diff_2487000_1963000# diff_2487000_1963000# GND efet w=15000 l=25000
+ ad=0 pd=0 as=1.519e+09 ps=314000 
M4314 diff_2409000_1980000# diff_2392000_1580000# diff_2405000_1947000# GND efet w=152500 l=10500
+ ad=0 pd=0 as=1.285e+09 ps=306000 
M4315 diff_2310000_1813000# diff_2319000_1882000# diff_2280000_1865000# GND efet w=58000 l=9000
+ ad=1.35903e+09 pd=724000 as=0 ps=0 
M4316 diff_2303000_1745000# diff_2319000_1882000# diff_2310000_1813000# GND efet w=154500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4317 diff_2405000_1947000# diff_2382000_1914000# diff_2385000_1734000# GND efet w=122000 l=11000
+ ad=0 pd=0 as=9.52033e+08 ps=508000 
M4318 diff_2310000_1813000# diff_2303000_1745000# diff_2271000_1558000# GND efet w=163500 l=9500
+ ad=0 pd=0 as=2.81033e+08 ps=788000 
M4319 diff_2303000_1745000# diff_2329000_1774000# diff_2310000_1813000# GND efet w=153000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4320 diff_2126000_1704000# diff_2248000_788000# diff_2271000_1624000# GND efet w=15000 l=10000
+ ad=0 pd=0 as=1.132e+09 ps=176000 
M4321 diff_2183000_1678000# diff_2183000_1678000# diff_2197000_1603000# GND efet w=14000 l=20000
+ ad=0 pd=0 as=-1.93097e+09 ps=226000 
M4322 diff_2103000_1636000# diff_1439000_785000# diff_2049000_1769000# GND efet w=23000 l=15000
+ ad=1.15e+08 pd=56000 as=3.94e+08 ps=98000 
M4323 diff_2123000_1636000# diff_2108000_871000# diff_2103000_1636000# GND efet w=23000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M4324 diff_2197000_1603000# diff_2123000_1636000# diff_2123000_1636000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4325 diff_2103000_1606000# diff_1439000_785000# diff_2049000_1456000# GND efet w=23000 l=15000
+ ad=1.15e+08 pd=56000 as=3.61e+08 ps=104000 
M4326 diff_2123000_1606000# diff_2108000_871000# diff_2103000_1606000# GND efet w=23000 l=15000
+ ad=-1.42397e+09 pd=426000 as=0 ps=0 
M4327 diff_2015000_1467000# diff_2003000_996000# diff_1996000_1467000# GND efet w=122000 l=12000
+ ad=1.35e+09 pd=220000 as=0 ps=0 
M4328 diff_1889000_1428000# diff_1880000_1449000# diff_1869000_1455000# GND efet w=200500 l=9500
+ ad=-9.97935e+08 pd=788000 as=0 ps=0 
M4329 diff_1943000_1520000# diff_1931000_1553000# diff_1889000_1428000# GND efet w=61000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4330 diff_1869000_1407000# diff_1857000_1018000# diff_1850000_1375000# GND efet w=107000 l=12000
+ ad=-1.32397e+09 pd=494000 as=9.57e+08 ps=228000 
M4331 diff_1889000_1428000# diff_1880000_1417000# diff_1869000_1407000# GND efet w=200500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4332 diff_1852000_1318000# diff_1836000_1363000# diff_1833000_1282000# GND efet w=104500 l=12500
+ ad=1.046e+09 pd=226000 as=8.78e+08 ps=222000 
M4333 diff_1943000_1345000# diff_1931000_1327000# diff_1889000_1428000# GND efet w=66000 l=10000
+ ad=1.268e+09 pd=206000 as=0 ps=0 
M4334 diff_2052000_1524000# diff_2049000_1456000# diff_2035000_1429000# GND efet w=185500 l=10500
+ ad=1.242e+09 pd=302000 as=2.64033e+08 ps=860000 
M4335 diff_2015000_1385000# diff_2003000_996000# diff_1996000_1361000# GND efet w=119000 l=12000
+ ad=1.26e+09 pd=214000 as=1.764e+09 ps=362000 
M4336 diff_2052000_1346000# diff_2049000_1392000# diff_2035000_1429000# GND efet w=187500 l=10500
+ ad=1.269e+09 pd=306000 as=0 ps=0 
M4337 diff_1851000_1157000# diff_1836000_1363000# diff_1833000_1157000# GND efet w=104500 l=11500
+ ad=1.13e+09 pd=228000 as=8.82e+08 ps=222000 
M4338 diff_1996000_1361000# diff_1982000_1350000# diff_1981000_1324000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=3.96e+08 ps=80000 
M4339 diff_1869000_1407000# diff_1891000_1210000# diff_1892000_1235000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=9.58e+08 ps=138000 
M4340 diff_1931000_1327000# diff_1891000_1210000# diff_1869000_1407000# GND efet w=14500 l=82500
+ ad=5.29e+08 pd=132000 as=0 ps=0 
M4341 diff_1943000_1345000# diff_1891000_1210000# diff_1965000_1244000# GND efet w=14000 l=33000
+ ad=0 pd=0 as=5.6e+08 ps=98000 
M4342 diff_1892000_1235000# diff_1891000_1210000# diff_1869000_1078000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=-1.36797e+09 ps=504000 
M4343 diff_1931000_1176000# diff_1891000_1210000# diff_1869000_1078000# GND efet w=15000 l=78000
+ ad=5.99e+08 pd=146000 as=0 ps=0 
M4344 diff_1965000_1244000# diff_1891000_1210000# diff_1943000_1143000# GND efet w=15000 l=34000
+ ad=0 pd=0 as=1.154e+09 ps=208000 
M4345 diff_1869000_1078000# diff_1857000_1018000# diff_1850000_1078000# GND efet w=106500 l=12500
+ ad=0 pd=0 as=8.82e+08 ps=226000 
M4346 diff_1996000_1361000# diff_1996000_1361000# diff_2009000_1240000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=8.14e+08 ps=122000 
M4347 diff_1996000_1090000# diff_1996000_1090000# diff_2009000_1240000# GND efet w=14500 l=23500
+ ad=1.705e+09 pd=362000 as=0 ps=0 
M4348 diff_1996000_1090000# diff_1982000_1350000# diff_1981000_1167000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=3.78e+08 ps=78000 
M4349 diff_2123000_1606000# diff_2129000_1594000# diff_2136000_1579000# GND efet w=67000 l=10000
+ ad=0 pd=0 as=1.703e+09 ps=372000 
M4350 diff_2197000_1603000# diff_2123000_1606000# diff_2123000_1606000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4351 diff_2197000_1603000# diff_2183000_1493000# diff_2183000_1493000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=1.607e+09 ps=336000 
M4352 diff_2136000_1579000# diff_2126000_1544000# diff_2121000_1350000# GND efet w=128500 l=10500
+ ad=0 pd=0 as=9.36065e+08 ps=1.434e+06 
M4353 diff_2123000_1606000# diff_2129000_1594000# diff_2136000_1579000# GND efet w=75500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4354 diff_2121000_1350000# diff_2183000_1493000# diff_2123000_1606000# GND efet w=59000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4355 diff_2183000_1493000# diff_2206000_1539000# diff_2121000_1350000# GND efet w=65000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4356 diff_2121000_1350000# diff_2232000_1463000# diff_2183000_1493000# GND efet w=73000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4357 diff_2136000_1297000# diff_2126000_1327000# diff_2121000_1350000# GND efet w=130000 l=10000
+ ad=1.786e+09 pd=374000 as=0 ps=0 
M4358 diff_2122000_1260000# diff_2129000_1288000# diff_2136000_1297000# GND efet w=78000 l=10000
+ ad=-1.28597e+09 pd=458000 as=0 ps=0 
M4359 diff_2136000_1297000# diff_2129000_1288000# diff_2122000_1260000# GND efet w=64500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4360 diff_2121000_1350000# diff_2183000_1301000# diff_2122000_1260000# GND efet w=59000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4361 diff_2183000_1301000# diff_2129000_1288000# diff_2121000_1350000# GND efet w=65000 l=10000
+ ad=1.625e+09 pd=332000 as=0 ps=0 
M4362 diff_2121000_1350000# diff_2126000_1327000# diff_2183000_1301000# GND efet w=73000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4363 diff_2183000_1301000# diff_2183000_1301000# diff_2197000_1226000# GND efet w=14000 l=20000
+ ad=0 pd=0 as=-1.93197e+09 ps=226000 
M4364 diff_2103000_1260000# diff_1439000_785000# diff_2049000_1392000# GND efet w=22000 l=15000
+ ad=1.1e+08 pd=54000 as=3.74e+08 ps=96000 
M4365 diff_2122000_1260000# diff_2108000_871000# diff_2103000_1260000# GND efet w=22000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M4366 diff_2197000_1226000# diff_2122000_1260000# diff_2122000_1260000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4367 diff_2461000_1832000# diff_2392000_2433000# diff_2409000_1980000# GND efet w=153000 l=10000
+ ad=1.457e+09 pd=328000 as=0 ps=0 
M4368 diff_2628000_2040000# diff_2591000_970000# diff_2549000_1954000# GND efet w=89500 l=10500
+ ad=-1.79397e+09 pd=484000 as=0 ps=0 
M4369 diff_2652000_2076000# diff_2640000_933000# diff_2628000_2040000# GND efet w=22000 l=12000
+ ad=5.25e+08 pd=190000 as=0 ps=0 
M4370 diff_2800000_2075000# diff_2776000_764000# diff_2781000_2075000# GND efet w=108000 l=12000
+ ad=1.48e+09 pd=314000 as=1.107e+09 ps=226000 
M4371 diff_2886000_2178000# diff_2875000_2204000# diff_2830000_2241000# GND efet w=217500 l=10500
+ ad=-1.27893e+09 pd=910000 as=0 ps=0 
M4372 diff_2875000_2204000# diff_2914000_2317000# diff_2886000_2178000# GND efet w=61500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4373 diff_1707000_1881000# diff_2591000_970000# diff_2549000_1954000# GND efet w=90500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4374 diff_2480000_1745000# diff_2470000_1827000# diff_2461000_1832000# GND efet w=126500 l=9500
+ ad=-6.12967e+08 pd=590000 as=0 ps=0 
M4375 diff_2487000_1963000# diff_2470000_1827000# diff_2480000_1745000# GND efet w=61000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4376 diff_2549000_1954000# diff_2532000_1854000# diff_2532000_1854000# GND efet w=13000 l=16000
+ ad=0 pd=0 as=1.705e+09 ps=346000 
M4377 diff_2674000_2059000# diff_94000_5193000# diff_94000_5193000# GND efet w=13500 l=33500
+ ad=0 pd=0 as=0 ps=0 
M4378 diff_2684000_2154000# diff_94000_5193000# diff_2652000_2076000# GND efet w=14500 l=82500
+ ad=0 pd=0 as=0 ps=0 
M4379 diff_2684000_2154000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4380 diff_94000_5193000# diff_94000_5193000# diff_2673000_1830000# GND efet w=13000 l=32000
+ ad=0 pd=0 as=9.88e+08 ps=188000 
M4381 diff_2684000_1840000# diff_94000_5193000# diff_2651000_1920000# GND efet w=14000 l=74000
+ ad=-4.07967e+08 pd=734000 as=5.58e+08 ps=204000 
M4382 diff_94000_5193000# diff_94000_5193000# diff_2684000_1840000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4383 diff_2651000_1920000# diff_2640000_933000# diff_1707000_1881000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4384 diff_2651000_1920000# diff_2651000_1920000# diff_2651000_1920000# GND efet w=2000 l=4000
+ ad=0 pd=0 as=0 ps=0 
M4385 diff_2830000_2069000# diff_2582000_2724000# diff_2800000_2075000# GND efet w=88000 l=12000
+ ad=1.097e+09 pd=214000 as=0 ps=0 
M4386 diff_2865000_2160000# diff_2842000_1949000# diff_2846000_2124000# GND efet w=108500 l=12500
+ ad=-1.37997e+09 pd=502000 as=9.77e+08 ps=230000 
M4387 diff_2886000_2178000# diff_2875000_2169000# diff_2865000_2160000# GND efet w=216500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4388 diff_2930000_2100000# diff_2913000_2059000# diff_2886000_2178000# GND efet w=70500 l=9500
+ ad=9.4e+08 pd=174000 as=0 ps=0 
M4389 diff_816000_2341000# diff_2637000_2491000# diff_3028000_2299000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=1.859e+09 ps=396000 
M4390 diff_94000_5193000# diff_94000_5193000# diff_3098000_2318000# GND efet w=14000 l=32000
+ ad=0 pd=0 as=1.063e+09 ps=192000 
M4391 diff_3118000_2218000# diff_94000_5193000# diff_3028000_2299000# GND efet w=14000 l=74000
+ ad=-4.30967e+08 pd=702000 as=0 ps=0 
M4392 diff_94000_5193000# diff_94000_5193000# diff_3118000_2218000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4393 diff_847000_2341000# diff_2995000_2724000# diff_2914000_2317000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4394 diff_3028000_2299000# diff_2995000_2724000# diff_2544000_2207000# GND efet w=21000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4395 diff_3028000_2040000# diff_2995000_2724000# diff_3005000_2149000# GND efet w=21000 l=12000
+ ad=1.609e+09 pd=310000 as=3.57e+08 ps=76000 
M4396 diff_3011000_2111000# diff_2995000_2724000# diff_2987000_2077000# GND efet w=22000 l=11000
+ ad=4.18e+08 pd=82000 as=1.167e+09 ps=228000 
M4397 diff_2865000_2160000# diff_94000_5193000# diff_94000_5193000# GND efet w=13000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M4398 diff_2913000_2059000# diff_94000_5193000# diff_2865000_2160000# GND efet w=14500 l=82500
+ ad=2.09e+08 pd=82000 as=0 ps=0 
M4399 diff_2930000_2100000# diff_94000_5193000# diff_94000_5193000# GND efet w=13000 l=33000
+ ad=0 pd=0 as=0 ps=0 
M4400 diff_2987000_2077000# diff_2938000_823000# diff_2962000_2041000# GND efet w=21000 l=13000
+ ad=0 pd=0 as=3.57e+08 ps=76000 
M4401 diff_2830000_1864000# diff_94000_5193000# diff_94000_5193000# GND efet w=13000 l=24000
+ ad=-1.47967e+08 pd=734000 as=0 ps=0 
M4402 diff_2914000_1941000# diff_94000_5193000# diff_2830000_1864000# GND efet w=14000 l=73000
+ ad=1.38e+09 pd=316000 as=0 ps=0 
M4403 diff_94000_5193000# diff_94000_5193000# diff_2875000_1828000# GND efet w=14000 l=31000
+ ad=0 pd=0 as=9.24e+08 ps=180000 
M4404 diff_2554000_1747000# diff_2544000_1829000# diff_2532000_1854000# GND efet w=85500 l=10500
+ ad=-1.75297e+09 pd=358000 as=0 ps=0 
M4405 diff_2532000_1854000# diff_2447000_2716000# diff_2470000_1827000# GND efet w=23000 l=13000
+ ad=0 pd=0 as=3.79e+08 ps=104000 
M4406 diff_2406000_1691000# diff_2129000_1665000# diff_2385000_1734000# GND efet w=117500 l=10500
+ ad=1.283e+09 pd=296000 as=0 ps=0 
M4407 diff_2329000_1774000# diff_2392000_1580000# diff_2406000_1691000# GND efet w=148500 l=10500
+ ad=2.118e+09 pd=420000 as=0 ps=0 
M4408 diff_2461000_1726000# diff_2392000_2433000# diff_2329000_1774000# GND efet w=152000 l=10000
+ ad=1.433e+09 pd=326000 as=0 ps=0 
M4409 diff_2480000_1745000# diff_2470000_1735000# diff_2461000_1726000# GND efet w=125500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4410 diff_2549000_1954000# diff_2591000_970000# diff_2544000_1829000# GND efet w=87500 l=10500
+ ad=0 pd=0 as=1.112e+09 ps=222000 
M4411 diff_1503000_1891000# diff_2591000_970000# diff_2549000_1954000# GND efet w=73000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4412 diff_2673000_1830000# diff_2651000_1920000# diff_2655000_1780000# GND efet w=63000 l=10000
+ ad=0 pd=0 as=1.27603e+09 ps=880000 
M4413 diff_2684000_1840000# diff_2673000_1830000# diff_2655000_1780000# GND efet w=219500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4414 diff_2759000_1832000# diff_2712000_821000# diff_2684000_1840000# GND efet w=105000 l=12000
+ ad=1.53103e+09 pd=1.126e+06 as=0 ps=0 
M4415 diff_2532000_1765000# diff_2447000_2716000# diff_2470000_1735000# GND efet w=23000 l=13000
+ ad=1.666e+09 pd=340000 as=3.19e+08 ps=84000 
M4416 diff_2271000_1558000# diff_2248000_788000# diff_2271000_1624000# GND efet w=14000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4417 diff_2126000_1327000# diff_2290000_1481000# diff_2271000_1558000# GND efet w=124000 l=12000
+ ad=4.13033e+08 pd=698000 as=0 ps=0 
M4418 diff_2329000_1617000# diff_2290000_1481000# diff_2290000_1481000# GND efet w=15000 l=22000
+ ad=4.45e+08 pd=88000 as=1.085e+09 ps=214000 
M4419 diff_2129000_1665000# diff_2470000_1735000# diff_2480000_1745000# GND efet w=60000 l=9000
+ ad=1.499e+09 pd=306000 as=0 ps=0 
M4420 diff_2554000_1747000# diff_2544000_1737000# diff_2532000_1765000# GND efet w=81000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4421 diff_2549000_1578000# diff_2591000_970000# diff_2544000_1737000# GND efet w=88500 l=10500
+ ad=-1.6429e+09 pd=914000 as=1.143e+09 ps=228000 
M4422 diff_2628000_1728000# diff_2591000_970000# diff_2549000_1578000# GND efet w=74000 l=11000
+ ad=1.016e+09 pd=186000 as=0 ps=0 
M4423 diff_1707000_1881000# diff_2776000_764000# diff_2684000_1840000# GND efet w=109500 l=12500
+ ad=0 pd=0 as=0 ps=0 
M4424 diff_2830000_1864000# diff_2582000_2724000# diff_1707000_1881000# GND efet w=88000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4425 diff_2914000_1941000# diff_2938000_823000# diff_1707000_1881000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4426 diff_2830000_1864000# diff_2842000_1949000# diff_2830000_1864000# GND efet w=4000 l=4000
+ ad=0 pd=0 as=0 ps=0 
M4427 diff_2914000_1941000# diff_2914000_1941000# diff_2914000_1941000# GND efet w=1000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4428 diff_2830000_1864000# diff_2842000_1949000# diff_1503000_1891000# GND efet w=109000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4429 diff_2684000_1778000# diff_2673000_1767000# diff_2655000_1780000# GND efet w=221500 l=10500
+ ad=-1.55597e+09 pd=492000 as=0 ps=0 
M4430 diff_2674000_1682000# diff_2652000_1699000# diff_2655000_1780000# GND efet w=71000 l=10000
+ ad=9.78e+08 pd=188000 as=0 ps=0 
M4431 diff_2759000_1758000# diff_2712000_821000# diff_2684000_1778000# GND efet w=105500 l=11500
+ ad=1.24e+09 pd=236000 as=0 ps=0 
M4432 diff_2532000_1765000# diff_2532000_1765000# diff_2549000_1578000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M4433 diff_2329000_1774000# diff_2329000_1774000# diff_2416000_1627000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=7.5e+08 ps=136000 
M4434 diff_2416000_1627000# diff_2409000_1603000# diff_2409000_1603000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=-2.10597e+09 ps=430000 
M4435 diff_2129000_1665000# diff_2129000_1665000# diff_2475000_1616000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=1.407e+09 ps=178000 
M4436 diff_2475000_1616000# diff_2487000_1586000# diff_2487000_1586000# GND efet w=15000 l=25000
+ ad=0 pd=0 as=1.494e+09 ps=314000 
M4437 diff_2409000_1603000# diff_2392000_1580000# diff_2406000_1570000# GND efet w=152000 l=10000
+ ad=0 pd=0 as=1.28e+09 ps=304000 
M4438 diff_82000_3097000# diff_2334000_1513000# diff_2290000_1481000# GND efet w=61000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4439 diff_2406000_1570000# diff_2382000_1537000# diff_82000_3097000# GND efet w=121000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4440 diff_2460000_1455000# diff_2392000_2433000# diff_2409000_1603000# GND efet w=153500 l=9500
+ ad=1.536e+09 pd=330000 as=0 ps=0 
M4441 diff_2628000_1664000# diff_2591000_970000# diff_2549000_1578000# GND efet w=89500 l=10500
+ ad=9.91e+08 pd=198000 as=0 ps=0 
M4442 diff_2652000_1699000# diff_2640000_933000# diff_2628000_1664000# GND efet w=22000 l=12000
+ ad=5.37e+08 pd=170000 as=0 ps=0 
M4443 diff_2800000_1698000# diff_2776000_764000# diff_2781000_1698000# GND efet w=108500 l=12500
+ ad=1.489e+09 pd=316000 as=1.044e+09 ps=226000 
M4444 diff_2886000_1802000# diff_2875000_1828000# diff_2830000_1864000# GND efet w=215500 l=10500
+ ad=-1.28193e+09 pd=908000 as=0 ps=0 
M4445 diff_2875000_1828000# diff_2914000_1941000# diff_2886000_1802000# GND efet w=61500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4446 diff_2628000_1544000# diff_2591000_970000# diff_2549000_1578000# GND efet w=89500 l=10500
+ ad=1.079e+09 pd=202000 as=0 ps=0 
M4447 diff_2480000_1368000# diff_2470000_1450000# diff_2460000_1455000# GND efet w=126500 l=9500
+ ad=-6.75967e+08 pd=590000 as=0 ps=0 
M4448 diff_2487000_1586000# diff_2470000_1450000# diff_2480000_1368000# GND efet w=61000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4449 diff_2549000_1578000# diff_2532000_1478000# diff_2532000_1478000# GND efet w=13000 l=17000
+ ad=0 pd=0 as=1.68e+09 ps=346000 
M4450 diff_2674000_1682000# diff_94000_5193000# diff_94000_5193000# GND efet w=13500 l=33500
+ ad=0 pd=0 as=0 ps=0 
M4451 diff_2684000_1778000# diff_94000_5193000# diff_2652000_1699000# GND efet w=14500 l=83500
+ ad=0 pd=0 as=0 ps=0 
M4452 diff_2684000_1778000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4453 diff_2673000_1453000# diff_94000_5193000# diff_94000_5193000# GND efet w=13500 l=33500
+ ad=9.84e+08 pd=188000 as=0 ps=0 
M4454 diff_2684000_1462000# diff_94000_5193000# diff_2652000_1544000# GND efet w=14000 l=76000
+ ad=-5.10967e+08 pd=732000 as=5.25e+08 ps=202000 
M4455 diff_94000_5193000# diff_94000_5193000# diff_2684000_1462000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4456 diff_2652000_1544000# diff_2640000_933000# diff_2628000_1544000# GND efet w=23000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4457 diff_2830000_1692000# diff_2582000_2724000# diff_2800000_1698000# GND efet w=88000 l=12000
+ ad=1.097e+09 pd=214000 as=0 ps=0 
M4458 diff_2865000_1783000# diff_2842000_1949000# diff_2846000_1747000# GND efet w=106500 l=11500
+ ad=-1.37197e+09 pd=500000 as=1.008e+09 ps=228000 
M4459 diff_2886000_1802000# diff_2875000_1792000# diff_2865000_1783000# GND efet w=214500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4460 diff_2930000_1723000# diff_2913000_1682000# diff_2886000_1802000# GND efet w=71500 l=9500
+ ad=9.61e+08 pd=176000 as=0 ps=0 
M4461 diff_2913000_1682000# diff_2913000_1682000# diff_2913000_1682000# GND efet w=500 l=11500
+ ad=2.14e+08 pd=86000 as=0 ps=0 
M4462 diff_3081000_2267000# diff_2533000_2491000# diff_2544000_2207000# GND efet w=108500 l=11500
+ ad=-1.50993e+09 pd=1.006e+06 as=0 ps=0 
M4463 diff_3098000_2318000# diff_3028000_2299000# diff_3081000_2267000# GND efet w=62500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4464 diff_3118000_2218000# diff_3098000_2318000# diff_3081000_2267000# GND efet w=215500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4465 diff_2544000_2207000# diff_3119000_2491000# diff_3118000_2218000# GND efet w=88000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4466 diff_816000_2341000# diff_2892000_2724000# diff_3118000_2218000# GND efet w=88000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M4467 diff_3081000_2267000# diff_2533000_2491000# diff_3062000_2095000# GND efet w=108500 l=12500
+ ad=0 pd=0 as=1.183e+09 ps=232000 
M4468 diff_3118000_2155000# diff_3108000_2143000# diff_3081000_2267000# GND efet w=214500 l=9500
+ ad=-1.54497e+09 pd=470000 as=0 ps=0 
M4469 diff_3098000_2060000# diff_3092000_2085000# diff_3081000_2267000# GND efet w=70500 l=10500
+ ad=9.88e+08 pd=188000 as=0 ps=0 
M4470 diff_3052000_2040000# diff_2637000_2491000# diff_3028000_2040000# GND efet w=22000 l=11000
+ ad=4.18e+08 pd=82000 as=0 ps=0 
M4471 diff_1707000_1881000# diff_2637000_2491000# diff_3028000_1922000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=1.856e+09 ps=396000 
M4472 diff_3197000_2095000# diff_3119000_2491000# diff_3118000_2155000# GND efet w=88000 l=12000
+ ad=1.222e+09 pd=214000 as=0 ps=0 
M4473 diff_2628000_2040000# diff_2892000_2724000# diff_3212000_2093000# GND efet w=88000 l=13000
+ ad=0 pd=0 as=9.15e+08 ps=210000 
M4474 diff_3098000_2060000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=34000
+ ad=0 pd=0 as=0 ps=0 
M4475 diff_3118000_2155000# diff_94000_5193000# diff_3092000_2085000# GND efet w=14000 l=85000
+ ad=0 pd=0 as=1.75e+08 ps=64000 
M4476 diff_94000_5193000# diff_94000_5193000# diff_3118000_2155000# GND efet w=13000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M4477 diff_94000_5193000# diff_94000_5193000# diff_3098000_1942000# GND efet w=14000 l=32000
+ ad=0 pd=0 as=1.062e+09 ps=192000 
M4478 diff_3118000_1842000# diff_94000_5193000# diff_3028000_1922000# GND efet w=14000 l=72000
+ ad=-4.07967e+08 pd=706000 as=0 ps=0 
M4479 diff_94000_5193000# diff_94000_5193000# diff_3118000_1842000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4480 diff_1503000_1891000# diff_2995000_2724000# diff_2914000_1941000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4481 diff_3028000_1922000# diff_2995000_2724000# diff_2759000_1832000# GND efet w=21000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4482 diff_3028000_1663000# diff_2995000_2724000# diff_3005000_1772000# GND efet w=21000 l=12000
+ ad=1.588e+09 pd=308000 as=3.57e+08 ps=76000 
M4483 diff_3011000_1734000# diff_2995000_2724000# diff_2987000_1700000# GND efet w=22000 l=12000
+ ad=4.18e+08 pd=82000 as=1.157e+09 ps=228000 
M4484 diff_2865000_1783000# diff_94000_5193000# diff_94000_5193000# GND efet w=13000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M4485 diff_2913000_1682000# diff_94000_5193000# diff_2865000_1783000# GND efet w=14500 l=82500
+ ad=0 pd=0 as=0 ps=0 
M4486 diff_2930000_1723000# diff_94000_5193000# diff_94000_5193000# GND efet w=13000 l=33000
+ ad=0 pd=0 as=0 ps=0 
M4487 diff_2987000_1700000# diff_2938000_823000# diff_2962000_1663000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=3.96e+08 ps=80000 
M4488 diff_94000_5193000# diff_94000_5193000# diff_2830000_1487000# GND efet w=13000 l=24000
+ ad=0 pd=0 as=-1.93967e+08 ps=728000 
M4489 diff_2914000_1564000# diff_94000_5193000# diff_2830000_1487000# GND efet w=14000 l=75000
+ ad=1.373e+09 pd=314000 as=0 ps=0 
M4490 diff_94000_5193000# diff_94000_5193000# diff_2875000_1450000# GND efet w=14000 l=32000
+ ad=0 pd=0 as=9.28e+08 ps=180000 
M4491 diff_2652000_1544000# diff_2652000_1544000# diff_2652000_1544000# GND efet w=1500 l=3500
+ ad=0 pd=0 as=0 ps=0 
M4492 diff_2554000_1371000# diff_2544000_1452000# diff_2532000_1478000# GND efet w=85000 l=10000
+ ad=-1.75197e+09 pd=358000 as=0 ps=0 
M4493 diff_2532000_1478000# diff_2447000_2716000# diff_2470000_1450000# GND efet w=22000 l=14000
+ ad=0 pd=0 as=3.37e+08 ps=100000 
M4494 diff_2271000_1166000# diff_2289000_1293000# diff_2126000_1327000# GND efet w=125000 l=12000
+ ad=-3.42967e+08 pd=728000 as=0 ps=0 
M4495 diff_2103000_1229000# diff_1439000_785000# diff_2049000_1080000# GND efet w=23000 l=15000
+ ad=1.15e+08 pd=56000 as=3.51e+08 ps=106000 
M4496 diff_2122000_1229000# diff_2108000_871000# diff_2103000_1229000# GND efet w=23000 l=14000
+ ad=-1.37397e+09 pd=428000 as=0 ps=0 
M4497 diff_2015000_1090000# diff_2003000_996000# diff_1996000_1090000# GND efet w=122000 l=12000
+ ad=1.369e+09 pd=220000 as=0 ps=0 
M4498 diff_1889000_1051000# diff_1880000_1072000# diff_1869000_1078000# GND efet w=199500 l=9500
+ ad=-1.04493e+09 pd=786000 as=0 ps=0 
M4499 diff_1943000_1143000# diff_1931000_1176000# diff_1889000_1051000# GND efet w=61000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4500 diff_1869000_1028000# diff_1857000_1018000# diff_1850000_998000# GND efet w=107000 l=12000
+ ad=-1.42497e+09 pd=490000 as=9.83e+08 ps=228000 
M4501 diff_1889000_1051000# diff_1880000_1040000# diff_1869000_1028000# GND efet w=199500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4502 diff_1851000_942000# diff_1836000_1363000# diff_1833000_905000# GND efet w=103500 l=11500
+ ad=1.061e+09 pd=226000 as=9.19e+08 ps=220000 
M4503 diff_1943000_969000# diff_1930000_948000# diff_1889000_1051000# GND efet w=65000 l=10000
+ ad=1.236e+09 pd=204000 as=0 ps=0 
M4504 diff_2052000_1147000# diff_2049000_1080000# diff_2035000_1052000# GND efet w=183500 l=10500
+ ad=1.239e+09 pd=302000 as=2.86033e+08 ps=856000 
M4505 diff_2015000_1008000# diff_2003000_996000# diff_1996000_984000# GND efet w=118500 l=11500
+ ad=1.26e+09 pd=214000 as=1.786e+09 ps=362000 
M4506 diff_2052000_969000# diff_2049000_1016000# diff_2035000_1052000# GND efet w=188500 l=10500
+ ad=1.279e+09 pd=308000 as=0 ps=0 
M4507 diff_1996000_984000# diff_1982000_1350000# diff_1981000_947000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=3.78e+08 ps=78000 
M4508 diff_1869000_1028000# diff_1891000_905000# diff_1891000_876000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=5.84e+08 ps=100000 
M4509 diff_1930000_948000# diff_1891000_905000# diff_1869000_1028000# GND efet w=13500 l=85500
+ ad=5.46e+08 pd=132000 as=0 ps=0 
M4510 diff_1943000_969000# diff_1891000_905000# diff_1965000_869000# GND efet w=14000 l=34000
+ ad=0 pd=0 as=5.25e+08 ps=94000 
M4511 diff_1996000_984000# diff_1996000_984000# diff_2009000_876000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=5.18e+08 ps=94000 
M4512 diff_2122000_1229000# diff_2129000_1218000# diff_2136000_1203000# GND efet w=67500 l=9500
+ ad=0 pd=0 as=1.665e+09 ps=372000 
M4513 diff_2197000_1226000# diff_2122000_1229000# diff_2122000_1229000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4514 diff_2126000_1327000# diff_2248000_788000# diff_2272000_1244000# GND efet w=14000 l=11000
+ ad=0 pd=0 as=4.91e+08 ps=96000 
M4515 diff_2272000_1244000# diff_2248000_788000# diff_2271000_1166000# GND efet w=14000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4516 diff_2197000_1226000# diff_2183000_1117000# diff_2183000_1117000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=1.608e+09 ps=336000 
M4517 diff_2136000_1203000# diff_2126000_1168000# diff_2122000_972000# GND efet w=128000 l=11000
+ ad=0 pd=0 as=9.38065e+08 ps=1.436e+06 
M4518 diff_2122000_1229000# diff_2129000_1218000# diff_2136000_1203000# GND efet w=75500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4519 diff_2122000_972000# diff_2183000_1117000# diff_2122000_1229000# GND efet w=59000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4520 diff_2183000_1117000# diff_2206000_1163000# diff_2122000_972000# GND efet w=66000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4521 diff_2122000_972000# diff_2232000_1087000# diff_2183000_1117000# GND efet w=74000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4522 diff_2136000_921000# diff_2126000_951000# diff_2122000_972000# GND efet w=131500 l=10500
+ ad=1.729e+09 pd=372000 as=0 ps=0 
M4523 diff_2122000_883000# diff_2129000_912000# diff_2136000_921000# GND efet w=77500 l=10500
+ ad=-1.26597e+09 pd=456000 as=0 ps=0 
M4524 diff_2136000_921000# diff_2129000_912000# diff_2122000_883000# GND efet w=64500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4525 diff_2122000_972000# diff_2183000_925000# diff_2122000_883000# GND efet w=59000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4526 diff_2183000_925000# diff_2206000_953000# diff_2122000_972000# GND efet w=66000 l=10000
+ ad=1.6e+09 pd=330000 as=0 ps=0 
M4527 diff_2122000_972000# diff_2232000_994000# diff_2183000_925000# GND efet w=74000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4528 diff_82000_3097000# diff_2334000_1371000# diff_2289000_1293000# GND efet w=66000 l=10000
+ ad=0 pd=0 as=1.228e+09 ps=222000 
M4529 diff_2405000_1314000# diff_2129000_1288000# diff_82000_3097000# GND efet w=118500 l=10500
+ ad=1.293e+09 pd=298000 as=0 ps=0 
M4530 diff_2334000_1371000# diff_2392000_1580000# diff_2405000_1314000# GND efet w=149000 l=10000
+ ad=-2.07797e+09 pd=420000 as=0 ps=0 
M4531 diff_2460000_1349000# diff_2392000_2433000# diff_2334000_1371000# GND efet w=153000 l=10000
+ ad=1.528e+09 pd=330000 as=0 ps=0 
M4532 diff_2480000_1368000# diff_2470000_1357000# diff_2460000_1349000# GND efet w=126500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4533 diff_2549000_1578000# diff_2591000_970000# diff_2544000_1452000# GND efet w=88500 l=10500
+ ad=0 pd=0 as=1.129e+09 ps=224000 
M4534 diff_2628000_1463000# diff_2591000_970000# diff_2549000_1578000# GND efet w=73000 l=11000
+ ad=9.55e+08 pd=184000 as=0 ps=0 
M4535 diff_2673000_1453000# diff_2652000_1544000# diff_2655000_1403000# GND efet w=62000 l=10000
+ ad=0 pd=0 as=1.29703e+09 ps=876000 
M4536 diff_2684000_1462000# diff_2673000_1453000# diff_2655000_1403000# GND efet w=219500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4537 diff_2759000_1455000# diff_2712000_821000# diff_2684000_1462000# GND efet w=104500 l=12500
+ ad=1.65703e+09 pd=1.144e+06 as=0 ps=0 
M4538 diff_2532000_1388000# diff_2447000_2716000# diff_2470000_1357000# GND efet w=23000 l=13000
+ ad=1.672e+09 pd=342000 as=3.2e+08 ps=84000 
M4539 diff_2289000_1293000# diff_2289000_1293000# diff_2328000_1245000# GND efet w=16000 l=24000
+ ad=0 pd=0 as=4.93e+08 ps=92000 
M4540 diff_2328000_1245000# diff_2289000_1090000# diff_2289000_1090000# GND efet w=15000 l=25000
+ ad=0 pd=0 as=1.384e+09 ps=242000 
M4541 diff_2292000_953000# diff_2289000_1090000# diff_2271000_1166000# GND efet w=123000 l=12000
+ ad=-9.30967e+08 pd=548000 as=0 ps=0 
M4542 diff_2129000_1288000# diff_2470000_1357000# diff_2480000_1368000# GND efet w=61000 l=10000
+ ad=1.426e+09 pd=306000 as=0 ps=0 
M4543 diff_2554000_1371000# diff_2544000_1361000# diff_2532000_1388000# GND efet w=81000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4544 diff_2549000_1201000# diff_2591000_970000# diff_2544000_1361000# GND efet w=87500 l=10500
+ ad=-1.6879e+09 pd=914000 as=1.141e+09 ps=226000 
M4545 diff_2628000_1352000# diff_2591000_970000# diff_2549000_1201000# GND efet w=73000 l=11000
+ ad=1.007e+09 pd=184000 as=0 ps=0 
M4546 diff_816000_1587000# diff_2776000_764000# diff_2684000_1462000# GND efet w=109500 l=12500
+ ad=0 pd=0 as=0 ps=0 
M4547 diff_2830000_1487000# diff_2582000_2724000# diff_816000_1587000# GND efet w=88000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4548 diff_2914000_1564000# diff_2938000_823000# diff_816000_1587000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4549 diff_2914000_1564000# diff_2914000_1564000# diff_2914000_1564000# GND efet w=1000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4550 diff_2830000_1487000# diff_2842000_1949000# diff_847000_1587000# GND efet w=107500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M4551 diff_2684000_1401000# diff_2673000_1390000# diff_2655000_1403000# GND efet w=220500 l=10500
+ ad=-1.66897e+09 pd=488000 as=0 ps=0 
M4552 diff_2674000_1305000# diff_2651000_1322000# diff_2655000_1403000# GND efet w=70000 l=10000
+ ad=9.62e+08 pd=186000 as=0 ps=0 
M4553 diff_2759000_1380000# diff_2712000_821000# diff_2684000_1401000# GND efet w=105500 l=12500
+ ad=1.246e+09 pd=236000 as=0 ps=0 
M4554 diff_2532000_1388000# diff_2532000_1388000# diff_2549000_1201000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M4555 diff_2334000_1371000# diff_2334000_1371000# diff_2415000_1250000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=7.62e+08 ps=140000 
M4556 diff_2415000_1250000# diff_2409000_1226000# diff_2409000_1226000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=2e+09 ps=430000 
M4557 diff_2129000_1288000# diff_2129000_1288000# diff_2475000_1238000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=1.422e+09 ps=180000 
M4558 diff_2475000_1238000# diff_2487000_1208000# diff_2487000_1208000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=1.495e+09 ps=314000 
M4559 diff_2409000_1226000# diff_2392000_1580000# diff_2405000_1193000# GND efet w=153500 l=11500
+ ad=0 pd=0 as=1.285e+09 ps=304000 
M4560 diff_2405000_1193000# diff_2382000_1160000# diff_2341000_1052000# GND efet w=122000 l=11000
+ ad=0 pd=0 as=5.35098e+08 ps=1.072e+06 
M4561 diff_2341000_1052000# diff_2334000_1126000# diff_2289000_1090000# GND efet w=62000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4562 diff_2461000_1078000# diff_2392000_2433000# diff_2409000_1226000# GND efet w=152500 l=10500
+ ad=1.445e+09 pd=328000 as=0 ps=0 
M4563 diff_2628000_1287000# diff_2591000_970000# diff_2549000_1201000# GND efet w=90500 l=10500
+ ad=1.012e+09 pd=200000 as=0 ps=0 
M4564 diff_2651000_1322000# diff_2640000_933000# diff_2628000_1287000# GND efet w=23000 l=11000
+ ad=5.69e+08 pd=194000 as=0 ps=0 
M4565 diff_2800000_1321000# diff_2776000_764000# diff_2781000_1321000# GND efet w=109500 l=12500
+ ad=1.479e+09 pd=316000 as=1.068e+09 ps=228000 
M4566 diff_2886000_1425000# diff_2875000_1450000# diff_2830000_1487000# GND efet w=216500 l=10500
+ ad=-1.27793e+09 pd=908000 as=0 ps=0 
M4567 diff_2875000_1450000# diff_2914000_1564000# diff_2886000_1425000# GND efet w=63500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4568 diff_2628000_1167000# diff_2591000_970000# diff_2549000_1201000# GND efet w=90500 l=10500
+ ad=1.078e+09 pd=204000 as=0 ps=0 
M4569 diff_2341000_1052000# diff_2470000_1073000# diff_2461000_1078000# GND efet w=125500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4570 diff_2487000_1208000# diff_2470000_1073000# diff_2341000_1052000# GND efet w=60000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4571 diff_2549000_1201000# diff_2532000_1101000# diff_2532000_1101000# GND efet w=13000 l=18000
+ ad=0 pd=0 as=1.685e+09 ps=342000 
M4572 diff_2674000_1305000# diff_94000_5193000# diff_94000_5193000# GND efet w=13500 l=33500
+ ad=0 pd=0 as=0 ps=0 
M4573 diff_2684000_1401000# diff_94000_5193000# diff_2651000_1322000# GND efet w=14500 l=83500
+ ad=0 pd=0 as=0 ps=0 
M4574 diff_2684000_1401000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M4575 diff_2673000_1076000# diff_94000_5193000# diff_94000_5193000# GND efet w=13000 l=33000
+ ad=9.87e+08 pd=188000 as=0 ps=0 
M4576 diff_2684000_1085000# diff_94000_5193000# diff_2652000_1167000# GND efet w=14000 l=76000
+ ad=-3.80967e+08 pd=732000 as=5.34e+08 ps=200000 
M4577 diff_94000_5193000# diff_94000_5193000# diff_2684000_1085000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4578 diff_2652000_1167000# diff_2640000_933000# diff_2628000_1167000# GND efet w=23000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4579 diff_2652000_1167000# diff_2652000_1167000# diff_2652000_1167000# GND efet w=1500 l=3500
+ ad=0 pd=0 as=0 ps=0 
M4580 diff_2554000_993000# diff_2544000_1075000# diff_2532000_1101000# GND efet w=84500 l=10500
+ ad=-1.75297e+09 pd=358000 as=0 ps=0 
M4581 diff_2532000_1101000# diff_2447000_2716000# diff_2470000_1073000# GND efet w=23000 l=14000
+ ad=0 pd=0 as=3.37e+08 ps=84000 
M4582 diff_2341000_1052000# diff_2408000_957000# diff_2384000_972000# GND efet w=66000 l=10000
+ ad=0 pd=0 as=1.752e+09 ps=360000 
M4583 diff_2549000_1201000# diff_2591000_970000# diff_2544000_1075000# GND efet w=87500 l=10500
+ ad=0 pd=0 as=1.107e+09 ps=222000 
M4584 diff_2628000_1087000# diff_2591000_970000# diff_2549000_1201000# GND efet w=73000 l=11000
+ ad=9.55e+08 pd=184000 as=0 ps=0 
M4585 diff_2673000_1076000# diff_2652000_1167000# diff_2655000_1026000# GND efet w=63000 l=10000
+ ad=0 pd=0 as=1.22803e+09 ps=880000 
M4586 diff_2830000_1315000# diff_2582000_2724000# diff_2800000_1321000# GND efet w=88000 l=12000
+ ad=1.097e+09 pd=214000 as=0 ps=0 
M4587 diff_2865000_1406000# diff_2842000_1949000# diff_2846000_1371000# GND efet w=107500 l=11500
+ ad=-1.40597e+09 pd=504000 as=1.062e+09 ps=230000 
M4588 diff_2886000_1425000# diff_2875000_1415000# diff_2865000_1406000# GND efet w=214500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4589 diff_2930000_1346000# diff_2913000_1305000# diff_2886000_1425000# GND efet w=69500 l=9500
+ ad=9.44e+08 pd=174000 as=0 ps=0 
M4590 diff_2913000_1305000# diff_2913000_1305000# diff_2913000_1305000# GND efet w=500 l=11500
+ ad=2.13e+08 pd=86000 as=0 ps=0 
M4591 diff_3081000_1718000# diff_2533000_2491000# diff_2759000_1832000# GND efet w=108000 l=12000
+ ad=-1.47493e+09 pd=1.008e+06 as=0 ps=0 
M4592 diff_3098000_1942000# diff_3028000_1922000# diff_3081000_1718000# GND efet w=62500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4593 diff_3118000_1842000# diff_3098000_1942000# diff_3081000_1718000# GND efet w=213500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4594 diff_2759000_1832000# diff_3119000_2491000# diff_3118000_1842000# GND efet w=88000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4595 diff_1707000_1881000# diff_2892000_2724000# diff_3118000_1842000# GND efet w=89000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M4596 diff_3081000_1718000# diff_2533000_2491000# diff_3062000_1718000# GND efet w=109000 l=12000
+ ad=0 pd=0 as=1.183e+09 ps=232000 
M4597 diff_3118000_1778000# diff_3108000_1767000# diff_3081000_1718000# GND efet w=214500 l=9500
+ ad=-1.46097e+09 pd=472000 as=0 ps=0 
M4598 diff_3098000_1682000# diff_3092000_1709000# diff_3081000_1718000# GND efet w=69500 l=10500
+ ad=1.014e+09 pd=190000 as=0 ps=0 
M4599 diff_3052000_1663000# diff_2637000_2491000# diff_3028000_1663000# GND efet w=22000 l=12000
+ ad=4.18e+08 pd=82000 as=0 ps=0 
M4600 diff_816000_1587000# diff_2637000_2491000# diff_3028000_1545000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=1.864e+09 ps=396000 
M4601 diff_3197000_1718000# diff_3119000_2491000# diff_3118000_1778000# GND efet w=88000 l=12000
+ ad=1.221e+09 pd=214000 as=0 ps=0 
M4602 diff_3238000_1681000# diff_2892000_2724000# diff_3212000_1716000# GND efet w=88000 l=13000
+ ad=1.49e+09 pd=286000 as=9.13e+08 ps=210000 
M4603 diff_3098000_1682000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=33000
+ ad=0 pd=0 as=0 ps=0 
M4604 diff_3118000_1778000# diff_94000_5193000# diff_3092000_1709000# GND efet w=14000 l=83000
+ ad=0 pd=0 as=1.97e+08 ps=66000 
M4605 diff_3118000_1778000# diff_94000_5193000# diff_94000_5193000# GND efet w=13000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4606 diff_94000_5193000# diff_94000_5193000# diff_3098000_1565000# GND efet w=14000 l=32000
+ ad=0 pd=0 as=1.062e+09 ps=192000 
M4607 diff_3118000_1465000# diff_94000_5193000# diff_3028000_1545000# GND efet w=14000 l=74000
+ ad=-4.47967e+08 pd=704000 as=0 ps=0 
M4608 diff_94000_5193000# diff_94000_5193000# diff_3118000_1465000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4609 diff_847000_1587000# diff_2995000_2724000# diff_2914000_1564000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4610 diff_3028000_1545000# diff_2995000_2724000# diff_2759000_1455000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4611 diff_3028000_1286000# diff_2995000_2724000# diff_3005000_1395000# GND efet w=21000 l=12000
+ ad=1.588e+09 pd=308000 as=3.57e+08 ps=76000 
M4612 diff_3011000_1357000# diff_2995000_2724000# diff_2987000_1323000# GND efet w=21000 l=12000
+ ad=3.99e+08 pd=80000 as=1.144e+09 ps=226000 
M4613 diff_2865000_1406000# diff_94000_5193000# diff_94000_5193000# GND efet w=13000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M4614 diff_2913000_1305000# diff_94000_5193000# diff_2865000_1406000# GND efet w=14500 l=82500
+ ad=0 pd=0 as=0 ps=0 
M4615 diff_2930000_1346000# diff_94000_5193000# diff_94000_5193000# GND efet w=13000 l=33000
+ ad=0 pd=0 as=0 ps=0 
M4616 diff_2987000_1323000# diff_2938000_823000# diff_2962000_1286000# GND efet w=21000 l=13000
+ ad=0 pd=0 as=3.57e+08 ps=76000 
M4617 diff_94000_5193000# diff_94000_5193000# diff_2830000_1110000# GND efet w=13000 l=24000
+ ad=0 pd=0 as=-1.93967e+08 ps=728000 
M4618 diff_2914000_1187000# diff_94000_5193000# diff_2830000_1110000# GND efet w=14000 l=76000
+ ad=1.358e+09 pd=310000 as=0 ps=0 
M4619 diff_94000_5193000# diff_94000_5193000# diff_2875000_1073000# GND efet w=14000 l=32000
+ ad=0 pd=0 as=9.28e+08 ps=180000 
M4620 diff_2684000_1085000# diff_2673000_1076000# diff_2655000_1026000# GND efet w=220500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4621 diff_2759000_1078000# diff_2712000_821000# diff_2684000_1085000# GND efet w=104000 l=12000
+ ad=-1.76693e+09 pd=1.358e+06 as=0 ps=0 
M4622 diff_2554000_993000# diff_2544000_983000# diff_2532000_968000# GND efet w=82000 l=10000
+ ad=0 pd=0 as=1.759e+09 ps=340000 
M4623 diff_2550000_879000# diff_2591000_970000# diff_2544000_983000# GND efet w=88500 l=10500
+ ad=1.43603e+09 pd=536000 as=1.156e+09 ps=228000 
M4624 diff_2292000_953000# diff_2248000_788000# diff_2197000_895000# GND efet w=14000 l=11000
+ ad=0 pd=0 as=-3.35967e+08 ps=360000 
M4625 diff_2183000_925000# diff_2183000_925000# diff_2197000_895000# GND efet w=14000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M4626 diff_2103000_883000# diff_1439000_785000# diff_2049000_1016000# GND efet w=22000 l=14000
+ ad=1.1e+08 pd=54000 as=4.2e+08 ps=100000 
M4627 diff_2122000_883000# diff_2108000_871000# diff_2103000_883000# GND efet w=22000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M4628 diff_2197000_895000# diff_2122000_883000# diff_2122000_883000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4629 diff_1888000_764000# diff_1876000_750000# diff_1836000_1363000# GND efet w=72000 l=12000
+ ad=1.512e+09 pd=186000 as=0 ps=0 
M4630 diff_1857000_1018000# diff_1876000_750000# diff_1888000_764000# GND efet w=72000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4631 diff_2027000_787000# diff_1978000_775000# diff_1982000_1350000# GND efet w=74000 l=12000
+ ad=1.463e+09 pd=190000 as=9.71e+08 ps=210000 
M4632 diff_2003000_996000# diff_1978000_775000# diff_2027000_787000# GND efet w=81500 l=11500
+ ad=1.584e+09 pd=290000 as=0 ps=0 
M4633 diff_2117000_758000# diff_2103000_843000# diff_1439000_785000# GND efet w=74000 l=12000
+ ad=1.406e+09 pd=186000 as=0 ps=0 
M4634 diff_2248000_788000# diff_2199000_774000# diff_2218000_809000# GND efet w=74000 l=12000
+ ad=0 pd=0 as=1.191e+09 ps=184000 
M4635 diff_2532000_968000# diff_2447000_2716000# diff_2500000_969000# GND efet w=24000 l=14000
+ ad=0 pd=0 as=4.3e+08 ps=84000 
M4636 diff_2628000_975000# diff_2591000_970000# diff_2550000_879000# GND efet w=74000 l=11000
+ ad=1.016e+09 pd=186000 as=0 ps=0 
M4637 diff_816000_1210000# diff_2776000_764000# diff_2684000_1085000# GND efet w=110500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M4638 diff_2830000_1110000# diff_2582000_2724000# diff_816000_1210000# GND efet w=88000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M4639 diff_2914000_1187000# diff_2938000_823000# diff_816000_1210000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4640 diff_2914000_1187000# diff_2914000_1187000# diff_2914000_1187000# GND efet w=1000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4641 diff_2830000_1110000# diff_2842000_1949000# diff_847000_1210000# GND efet w=108500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M4642 diff_2684000_1023000# diff_2673000_1012000# diff_2655000_1026000# GND efet w=220500 l=10500
+ ad=-1.52797e+09 pd=490000 as=0 ps=0 
M4643 diff_2408000_867000# diff_2384000_972000# diff_2384000_972000# GND efet w=16000 l=24000
+ ad=1.829e+09 pd=236000 as=0 ps=0 
M4644 diff_2365000_781000# diff_2342000_760000# diff_2338000_781000# GND efet w=104000 l=10000
+ ad=-1.97997e+09 pd=326000 as=1.768e+09 ps=242000 
M4645 diff_2408000_867000# diff_2365000_781000# diff_2365000_781000# GND efet w=16000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M4646 diff_2447000_2716000# diff_2476000_759000# diff_2468000_786000# GND efet w=74000 l=11000
+ ad=0 pd=0 as=1.479e+09 ps=188000 
M4647 diff_2674000_928000# diff_2651000_946000# diff_2655000_1026000# GND efet w=70000 l=10000
+ ad=9.75e+08 pd=186000 as=0 ps=0 
M4648 diff_2759000_1004000# diff_2712000_821000# diff_2684000_1023000# GND efet w=105500 l=11500
+ ad=1.24e+09 pd=236000 as=0 ps=0 
M4649 diff_2532000_968000# diff_2532000_968000# diff_2550000_879000# GND efet w=15000 l=18000
+ ad=0 pd=0 as=0 ps=0 
M4650 diff_2628000_910000# diff_2591000_970000# diff_2550000_879000# GND efet w=89500 l=10500
+ ad=1.002e+09 pd=198000 as=0 ps=0 
M4651 diff_2651000_946000# diff_2640000_933000# diff_2628000_910000# GND efet w=22000 l=11000
+ ad=5.42e+08 pd=188000 as=0 ps=0 
M4652 diff_2799000_944000# diff_2776000_764000# diff_2781000_945000# GND efet w=110000 l=11000
+ ad=1.449e+09 pd=318000 as=1.116e+09 ps=228000 
M4653 diff_2886000_1048000# diff_2875000_1073000# diff_2830000_1110000# GND efet w=215500 l=10500
+ ad=-1.28593e+09 pd=906000 as=0 ps=0 
M4654 diff_2875000_1073000# diff_2914000_1187000# diff_2886000_1048000# GND efet w=63500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4655 diff_2674000_928000# diff_2667000_894000# diff_2668000_869000# GND efet w=14000 l=34000
+ ad=0 pd=0 as=4.82e+08 ps=90000 
M4656 diff_2684000_1023000# diff_2667000_894000# diff_2651000_946000# GND efet w=14500 l=82500
+ ad=0 pd=0 as=0 ps=0 
M4657 diff_2684000_1023000# diff_2667000_894000# diff_2744000_876000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=5.46e+08 ps=96000 
M4658 diff_2830000_938000# diff_2582000_2724000# diff_2799000_944000# GND efet w=88000 l=13000
+ ad=1.097e+09 pd=214000 as=0 ps=0 
M4659 diff_2865000_1028000# diff_2842000_1949000# diff_2846000_994000# GND efet w=108000 l=12000
+ ad=-1.40297e+09 pd=504000 as=1.017e+09 ps=230000 
M4660 diff_2886000_1048000# diff_2875000_1038000# diff_2865000_1028000# GND efet w=214500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4661 diff_2930000_970000# diff_2914000_928000# diff_2886000_1048000# GND efet w=68500 l=9500
+ ad=9.43e+08 pd=174000 as=0 ps=0 
M4662 diff_82000_3097000# diff_791000_355000# diff_968000_455000# GND efet w=508500 l=10500
+ ad=0 pd=0 as=1.14507e+09 ps=1.51e+06 
M4663 diff_980000_464000# diff_791000_355000# diff_791000_355000# GND efet w=35000 l=11000
+ ad=-1.74967e+08 pd=550000 as=0 ps=0 
M4664 diff_968000_455000# diff_968000_455000# diff_980000_464000# GND efet w=44000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4665 diff_968000_455000# diff_1115000_636000# diff_82000_3097000# GND efet w=333000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4666 diff_968000_455000# diff_1115000_636000# diff_82000_3097000# GND efet w=65000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4667 diff_136000_354000# diff_125000_346000# diff_105000_354000# GND efet w=693500 l=10500
+ ad=7.29229e+08 pd=4.198e+06 as=0 ps=0 
M4668 diff_802000_365000# diff_791000_355000# diff_597000_373000# GND efet w=235000 l=11000
+ ad=8.61262e+08 pd=4.3e+06 as=1.54223e+09 ps=3.358e+06 
M4669 diff_597000_373000# diff_588000_420000# diff_125000_346000# GND efet w=277500 l=10500
+ ad=0 pd=0 as=1.63407e+09 ps=1.612e+06 
M4670 diff_876000_465000# diff_791000_355000# diff_802000_365000# GND efet w=197500 l=10500
+ ad=1.559e+09 pd=196000 as=0 ps=0 
M4671 diff_928000_464000# diff_791000_355000# diff_802000_365000# GND efet w=197500 l=9500
+ ad=1.638e+09 pd=198000 as=0 ps=0 
M4672 diff_980000_464000# diff_968000_455000# diff_802000_365000# GND efet w=353000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4673 diff_1228000_660000# diff_1218000_655000# diff_1203000_545000# GND efet w=442000 l=10000
+ ad=-1.11897e+09 pd=460000 as=-9.23902e+08 ps=2.038e+06 
M4674 diff_1286000_578000# diff_1276000_567000# diff_1203000_545000# GND efet w=488500 l=10500
+ ad=-1.56897e+09 pd=504000 as=0 ps=0 
M4675 diff_1360000_692000# diff_1203000_545000# diff_1203000_545000# GND efet w=54500 l=9500
+ ad=5e+08 pd=90000 as=0 ps=0 
M4676 diff_1405000_650000# diff_1398000_597000# diff_1384000_624000# GND efet w=233000 l=10000
+ ad=-1.79097e+09 pd=316000 as=-3.50967e+08 ps=648000 
M4677 diff_1452000_699000# diff_1384000_624000# diff_1384000_624000# GND efet w=18000 l=10000
+ ad=4.64e+08 pd=88000 as=0 ps=0 
M4678 diff_1547000_715000# diff_1537000_704000# diff_1429000_566000# GND efet w=300500 l=10500
+ ad=-9.77967e+08 pd=434000 as=1.88707e+09 ps=1.498e+06 
M4679 diff_1503000_592000# diff_1203000_545000# diff_1429000_566000# GND efet w=277000 l=11000
+ ad=-2.12197e+09 pd=280000 as=0 ps=0 
M4680 diff_1384000_624000# diff_1371000_619000# diff_1276000_567000# GND efet w=37000 l=13000
+ ad=0 pd=0 as=6.37e+08 ps=180000 
M4681 diff_1203000_545000# diff_1203000_545000# diff_1203000_545000# GND efet w=6000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M4682 diff_1429000_566000# diff_1203000_545000# diff_1429000_544000# GND efet w=48000 l=11000
+ ad=0 pd=0 as=2.025e+09 ps=306000 
M4683 diff_1082000_465000# diff_968000_455000# diff_802000_365000# GND efet w=173000 l=10000
+ ad=1.386e+09 pd=174000 as=0 ps=0 
M4684 diff_1134000_464000# diff_968000_455000# diff_802000_365000# GND efet w=174000 l=10000
+ ad=1.406e+09 pd=176000 as=0 ps=0 
M4685 diff_458000_404000# diff_125000_346000# diff_136000_354000# GND efet w=246500 l=10500
+ ad=2.059e+09 pd=246000 as=0 ps=0 
M4686 diff_597000_373000# diff_588000_420000# diff_125000_346000# GND efet w=122500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4687 diff_458000_352000# diff_125000_346000# diff_136000_354000# GND efet w=246000 l=10000
+ ad=2.06e+09 pd=246000 as=0 ps=0 
M4688 diff_597000_373000# diff_173000_152000# diff_125000_346000# GND efet w=501500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4689 diff_802000_365000# diff_791000_355000# diff_597000_373000# GND efet w=514500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4690 diff_457000_301000# diff_125000_346000# diff_136000_354000# GND efet w=490000 l=10000
+ ad=5.01033e+08 pd=552000 as=0 ps=0 
M4691 diff_125000_346000# diff_125000_346000# diff_457000_301000# GND efet w=44000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4692 diff_173000_152000# diff_173000_152000# diff_598000_271000# GND efet w=36000 l=11000
+ ad=1.67707e+09 pd=1.472e+06 as=5.32e+08 ps=106000 
M4693 diff_459000_154000# diff_173000_152000# diff_136000_354000# GND efet w=606000 l=10000
+ ad=7.70327e+07 pd=612000 as=0 ps=0 
M4694 diff_136000_354000# diff_173000_152000# diff_183000_100000# GND efet w=832000 l=11000
+ ad=0 pd=0 as=-1.2729e+09 ps=1.39e+06 
M4695 diff_597000_373000# diff_639000_113000# diff_173000_152000# GND efet w=379500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4696 diff_708000_309000# diff_679000_1018000# diff_691000_114000# GND efet w=36000 l=13000
+ ad=8.52e+08 pd=166000 as=5.29e+08 ps=138000 
M4697 diff_701000_124000# diff_691000_114000# diff_173000_152000# GND efet w=397500 l=9500
+ ad=-2.06967e+08 pd=410000 as=0 ps=0 
M4698 diff_802000_365000# diff_791000_355000# diff_597000_373000# GND efet w=278000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4699 diff_1049000_100000# diff_968000_455000# diff_802000_365000# GND efet w=122500 l=10500
+ ad=2.66196e+08 pd=2.65e+06 as=0 ps=0 
M4700 diff_1219000_196000# diff_1203000_545000# diff_1049000_100000# GND efet w=191000 l=10000
+ ad=2.12626e+09 pd=4.536e+06 as=0 ps=0 
M4701 diff_1292000_491000# diff_1203000_545000# diff_1219000_196000# GND efet w=205500 l=10500
+ ad=1.364e+09 pd=204000 as=0 ps=0 
M4702 diff_1219000_196000# diff_1203000_545000# diff_1049000_100000# GND efet w=652000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4703 diff_1345000_491000# diff_1203000_545000# diff_1219000_196000# GND efet w=205000 l=10000
+ ad=1.332e+09 pd=204000 as=0 ps=0 
M4704 diff_1398000_490000# diff_1203000_545000# diff_1219000_196000# GND efet w=208500 l=10500
+ ad=1.327e+09 pd=206000 as=0 ps=0 
M4705 diff_1429000_566000# diff_1429000_566000# diff_1490000_540000# GND efet w=37000 l=10000
+ ad=0 pd=0 as=6.66e+08 ps=110000 
M4706 diff_1429000_566000# diff_1537000_704000# diff_1547000_715000# GND efet w=56000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4707 diff_1429000_544000# diff_1429000_566000# diff_1219000_196000# GND efet w=193500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4708 diff_1641000_566000# diff_1631000_556000# diff_1619000_122000# GND efet w=57000 l=11000
+ ad=-8.44967e+08 pd=442000 as=1.75107e+09 ps=1.5e+06 
M4709 diff_1641000_566000# diff_1631000_556000# diff_1619000_122000# GND efet w=303000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4710 diff_1703000_589000# diff_1693000_584000# diff_1619000_122000# GND efet w=276000 l=10000
+ ad=-2.04597e+09 pd=280000 as=0 ps=0 
M4711 diff_2591000_970000# diff_2597000_842000# diff_2590000_764000# GND efet w=74000 l=13000
+ ad=9.78e+08 pd=208000 as=1.332e+09 ps=184000 
M4712 diff_2680000_788000# diff_2658000_766000# diff_2640000_933000# GND efet w=73000 l=11000
+ ad=1.605e+09 pd=190000 as=0 ps=0 
M4713 diff_3081000_1341000# diff_2533000_2491000# diff_2759000_1455000# GND efet w=109000 l=12000
+ ad=-1.64493e+09 pd=1.012e+06 as=0 ps=0 
M4714 diff_3098000_1565000# diff_3028000_1545000# diff_3081000_1341000# GND efet w=63500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4715 diff_3488000_2724000# diff_3457000_2526000# diff_3467000_2537000# GND efet w=205500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4716 diff_3519000_2552000# diff_3485000_2777000# diff_3488000_2724000# GND efet w=246500 l=10500
+ ad=1.78033e+08 pd=524000 as=0 ps=0 
M4717 diff_3473000_793000# diff_3535000_2777000# diff_3519000_2552000# GND efet w=246500 l=10500
+ ad=1.03903e+09 pd=982000 as=0 ps=0 
M4718 diff_3570000_2748000# diff_3473000_793000# diff_3473000_793000# GND efet w=20000 l=9000
+ ad=4.6e+08 pd=86000 as=0 ps=0 
M4719 diff_3566000_784000# diff_3566000_784000# diff_3570000_2748000# GND efet w=20000 l=9000
+ ad=1.47033e+08 pd=948000 as=0 ps=0 
M4720 diff_3571000_2536000# diff_3560000_2527000# diff_3473000_793000# GND efet w=205500 l=10500
+ ad=-2.20967e+08 pd=442000 as=0 ps=0 
M4721 diff_3566000_784000# diff_3560000_2527000# diff_3571000_2536000# GND efet w=205500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4722 diff_3622000_2553000# diff_3588000_2777000# diff_3566000_784000# GND efet w=247000 l=10000
+ ad=1.77033e+08 pd=524000 as=0 ps=0 
M4723 diff_3595000_2394000# diff_3638000_2777000# diff_3622000_2553000# GND efet w=246500 l=10500
+ ad=2.54033e+08 pd=862000 as=0 ps=0 
M4724 diff_3674000_2748000# diff_3595000_2394000# diff_3595000_2394000# GND efet w=20000 l=10000
+ ad=4.4e+08 pd=84000 as=0 ps=0 
M4725 diff_3694000_2724000# diff_3694000_2724000# diff_3674000_2748000# GND efet w=20000 l=10000
+ ad=6.84033e+08 pd=994000 as=0 ps=0 
M4726 diff_3674000_2536000# diff_3664000_2526000# diff_3595000_2394000# GND efet w=205000 l=10000
+ ad=-1.92967e+08 pd=442000 as=0 ps=0 
M4727 diff_3694000_2724000# diff_3664000_2526000# diff_3674000_2536000# GND efet w=205000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4728 diff_3726000_2552000# diff_3691000_2777000# diff_3694000_2724000# GND efet w=246500 l=10500
+ ad=-5.89673e+07 pd=522000 as=0 ps=0 
M4729 diff_3748000_2433000# diff_3741000_2777000# diff_3726000_2552000# GND efet w=247000 l=11000
+ ad=-1.26697e+09 pd=662000 as=0 ps=0 
M4730 diff_3777000_2748000# diff_3748000_2433000# diff_3748000_2433000# GND efet w=20000 l=10000
+ ad=4.4e+08 pd=84000 as=0 ps=0 
M4731 diff_3738000_825000# diff_3738000_825000# diff_3777000_2748000# GND efet w=20000 l=10000
+ ad=5.25033e+08 pd=926000 as=0 ps=0 
M4732 diff_3777000_2536000# diff_3766000_2527000# diff_3748000_2433000# GND efet w=206000 l=10000
+ ad=-2.19967e+08 pd=442000 as=0 ps=0 
M4733 diff_3118000_1465000# diff_3098000_1565000# diff_3081000_1341000# GND efet w=214500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4734 diff_2759000_1455000# diff_3119000_2491000# diff_3118000_1465000# GND efet w=87000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4735 diff_816000_1587000# diff_2892000_2724000# diff_3118000_1465000# GND efet w=89000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M4736 diff_82000_3097000# diff_3255000_1458000# diff_816000_1587000# GND efet w=93000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4737 diff_3738000_825000# diff_3766000_2527000# diff_3777000_2536000# GND efet w=205500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4738 diff_3829000_2552000# diff_3793000_2777000# diff_3738000_825000# GND efet w=246000 l=10000
+ ad=4.90327e+07 pd=522000 as=0 ps=0 
M4739 diff_3829000_786000# diff_3845000_2777000# diff_3829000_2552000# GND efet w=246500 l=10500
+ ad=4.49033e+08 pd=930000 as=0 ps=0 
M4740 diff_3880000_2748000# diff_3829000_786000# diff_3829000_786000# GND efet w=20000 l=10000
+ ad=4.4e+08 pd=84000 as=0 ps=0 
M4741 diff_3900000_2724000# diff_3900000_2724000# diff_3880000_2748000# GND efet w=20000 l=10000
+ ad=-1.06297e+09 pd=680000 as=0 ps=0 
M4742 diff_3880000_2536000# diff_3870000_2526000# diff_3829000_786000# GND efet w=206000 l=10000
+ ad=-1.76967e+08 pd=444000 as=0 ps=0 
M4743 diff_3900000_2724000# diff_3870000_2526000# diff_3880000_2536000# GND efet w=206000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4744 diff_3932000_2552000# diff_3897000_2777000# diff_3900000_2724000# GND efet w=246000 l=10000
+ ad=4.90327e+07 pd=522000 as=0 ps=0 
M4745 diff_3921000_785000# diff_3948000_2777000# diff_3932000_2552000# GND efet w=246500 l=10500
+ ad=4.03033e+08 pd=952000 as=0 ps=0 
M4746 diff_3983000_2748000# diff_3921000_785000# diff_3921000_785000# GND efet w=20000 l=10000
+ ad=4.4e+08 pd=84000 as=0 ps=0 
M4747 diff_4003000_2724000# diff_4003000_2724000# diff_3983000_2748000# GND efet w=20000 l=10000
+ ad=5.32033e+08 pd=890000 as=0 ps=0 
M4748 diff_3983000_2536000# diff_3973000_2526000# diff_3921000_785000# GND efet w=205000 l=10000
+ ad=-1.92967e+08 pd=442000 as=0 ps=0 
M4749 diff_94000_5193000# diff_94000_5193000# diff_94000_5193000# GND efet w=1000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M4750 diff_94000_5193000# diff_94000_5193000# diff_2544000_2207000# GND efet w=14000 l=106000
+ ad=0 pd=0 as=0 ps=0 
M4751 diff_94000_5193000# diff_94000_5193000# diff_3426000_2320000# GND efet w=14000 l=34000
+ ad=0 pd=0 as=1.014e+09 ps=184000 
M4752 diff_3437000_2232000# diff_94000_5193000# diff_3373000_2283000# GND efet w=14000 l=76000
+ ad=-3.73967e+08 pd=720000 as=1.726e+09 ps=372000 
M4753 diff_94000_5193000# diff_94000_5193000# diff_3437000_2232000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4754 diff_816000_2341000# diff_3170000_2724000# diff_3373000_2283000# GND efet w=21000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4755 diff_3437000_2232000# diff_3438000_2491000# diff_816000_2341000# GND efet w=108000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4756 diff_3578000_2264000# diff_3566000_784000# diff_3437000_2232000# GND efet w=111000 l=12000
+ ad=-9.54967e+08 pd=706000 as=0 ps=0 
M4757 diff_3373000_2283000# diff_3353000_2408000# diff_2544000_2207000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4758 diff_3373000_2059000# diff_3353000_2408000# diff_3334000_2135000# GND efet w=22000 l=12000
+ ad=1.468e+09 pd=290000 as=7.86e+08 ps=156000 
M4759 diff_3334000_2135000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=104000
+ ad=0 pd=0 as=0 ps=0 
M4760 diff_3426000_2320000# diff_3373000_2283000# diff_82000_3097000# GND efet w=68000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4761 diff_3437000_2232000# diff_3426000_2320000# diff_82000_3097000# GND efet w=206500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4762 diff_2544000_2207000# diff_3473000_793000# diff_3437000_2232000# GND efet w=88000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4763 diff_3437000_2161000# diff_3427000_2150000# diff_82000_3097000# GND efet w=207500 l=9500
+ ad=-1.51297e+09 pd=478000 as=0 ps=0 
M4764 diff_3427000_2063000# diff_3409000_2088000# diff_82000_3097000# GND efet w=74000 l=10000
+ ad=9.95e+08 pd=184000 as=0 ps=0 
M4765 diff_3521000_2100000# diff_3473000_793000# diff_3437000_2161000# GND efet w=88000 l=12000
+ ad=9.04e+08 pd=212000 as=0 ps=0 
M4766 diff_847000_2341000# diff_3595000_2394000# diff_3578000_2264000# GND efet w=121000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4767 diff_4003000_2724000# diff_3973000_2526000# diff_3983000_2536000# GND efet w=205000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4768 diff_4035000_2552000# diff_4000000_2777000# diff_4003000_2724000# GND efet w=246500 l=10500
+ ad=-3.69673e+07 pd=522000 as=0 ps=0 
M4769 diff_4056000_2491000# diff_4051000_2777000# diff_4035000_2552000# GND efet w=246500 l=10500
+ ad=-1.03197e+09 pd=678000 as=0 ps=0 
M4770 diff_4086000_2748000# diff_4056000_2491000# diff_4056000_2491000# GND efet w=20000 l=10000
+ ad=4.4e+08 pd=84000 as=0 ps=0 
M4771 diff_4107000_2724000# diff_4107000_2724000# diff_4086000_2748000# GND efet w=20000 l=10000
+ ad=-9.89673e+07 pd=894000 as=0 ps=0 
M4772 diff_4086000_2536000# diff_4076000_2526000# diff_4056000_2491000# GND efet w=205000 l=10000
+ ad=-1.92967e+08 pd=442000 as=0 ps=0 
M4773 diff_4107000_2724000# diff_4076000_2526000# diff_4086000_2536000# GND efet w=205000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4774 diff_4138000_2552000# diff_4103000_2777000# diff_4107000_2724000# GND efet w=247500 l=10500
+ ad=-2.83967e+08 pd=556000 as=0 ps=0 
M4775 diff_4223000_2738000# diff_4223000_2738000# diff_4213000_2744000# GND efet w=14000 l=16000
+ ad=6.43033e+08 pd=870000 as=5.35e+08 ps=120000 
M4776 diff_4276000_2780000# diff_4276000_2780000# diff_4266000_2739000# GND efet w=16000 l=15000
+ ad=-4.95967e+08 pd=824000 as=7.7e+08 ps=170000 
M4777 diff_94000_5193000# diff_4362000_2477000# diff_4362000_2477000# GND efet w=15000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4778 diff_4251000_2644000# diff_4240000_2639000# diff_4223000_2738000# GND efet w=130500 l=10500
+ ad=-5.99673e+07 pd=594000 as=0 ps=0 
M4779 diff_4161000_2693000# diff_4154000_2675000# diff_4154000_2675000# GND efet w=15000 l=18000
+ ad=8.77e+08 pd=134000 as=-7.57967e+08 ps=644000 
M4780 diff_4154000_2675000# diff_4154000_2620000# diff_4138000_2552000# GND efet w=102000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4781 diff_4192000_2538000# diff_4181000_2527000# diff_4154000_2675000# GND efet w=119500 l=10500
+ ad=1.549e+09 pd=258000 as=0 ps=0 
M4782 diff_816000_2341000# diff_3488000_2724000# diff_3633000_2300000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=1.069e+09 ps=238000 
M4783 diff_94000_5193000# diff_94000_5193000# diff_3685000_2316000# GND efet w=15000 l=34000
+ ad=0 pd=0 as=1.14e+09 ps=194000 
M4784 diff_3697000_2231000# diff_94000_5193000# diff_3633000_2300000# GND efet w=14000 l=74000
+ ad=-3.98967e+08 pd=718000 as=0 ps=0 
M4785 diff_94000_5193000# diff_94000_5193000# diff_3697000_2231000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4786 diff_3633000_2300000# diff_3353000_2408000# diff_847000_2341000# GND efet w=21000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4787 diff_3397000_2059000# diff_3170000_2724000# diff_3373000_2059000# GND efet w=21000 l=12000
+ ad=3.78e+08 pd=78000 as=0 ps=0 
M4788 diff_94000_5193000# diff_94000_5193000# diff_2759000_1832000# GND efet w=14000 l=106000
+ ad=0 pd=0 as=0 ps=0 
M4789 diff_3427000_2063000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=34000
+ ad=0 pd=0 as=0 ps=0 
M4790 diff_3437000_2161000# diff_94000_5193000# diff_3409000_2088000# GND efet w=14500 l=81500
+ ad=0 pd=0 as=2.75e+08 ps=100000 
M4791 diff_3437000_2161000# diff_94000_5193000# diff_94000_5193000# GND efet w=15000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M4792 diff_94000_5193000# diff_94000_5193000# diff_3426000_1943000# GND efet w=14000 l=34000
+ ad=0 pd=0 as=1.009e+09 ps=184000 
M4793 diff_3437000_1855000# diff_94000_5193000# diff_3373000_1906000# GND efet w=14000 l=74000
+ ad=-4.09967e+08 pd=718000 as=1.725e+09 ps=372000 
M4794 diff_94000_5193000# diff_94000_5193000# diff_3437000_1855000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4795 diff_1707000_1881000# diff_3170000_2724000# diff_3373000_1906000# GND efet w=21000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4796 diff_3557000_2087000# diff_3438000_2491000# diff_3538000_2051000# GND efet w=107500 l=11500
+ ad=1.102e+09 pd=234000 as=9.57e+08 ps=230000 
M4797 diff_3578000_2124000# diff_3566000_784000# diff_3557000_2087000# GND efet w=111000 l=12000
+ ad=1.496e+09 pd=290000 as=0 ps=0 
M4798 diff_3610000_2037000# diff_3595000_2394000# diff_3578000_2124000# GND efet w=122000 l=12000
+ ad=1.342e+09 pd=284000 as=0 ps=0 
M4799 diff_3633000_2077000# diff_3353000_2408000# diff_3610000_2037000# GND efet w=21000 l=13000
+ ad=7.97e+08 pd=154000 as=0 ps=0 
M4800 diff_816000_2341000# diff_3801000_831000# diff_3697000_2231000# GND efet w=104000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4801 diff_3847000_2257000# diff_3829000_786000# diff_816000_2341000# GND efet w=104000 l=12000
+ ad=-2.77967e+08 pd=716000 as=0 ps=0 
M4802 diff_3685000_2316000# diff_3633000_2300000# diff_82000_3097000# GND efet w=67500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4803 diff_3697000_2231000# diff_3685000_2316000# diff_82000_3097000# GND efet w=204000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4804 diff_3578000_2264000# diff_3738000_825000# diff_3697000_2231000# GND efet w=88000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4805 diff_94000_5193000# diff_94000_5193000# diff_3847000_2257000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4806 diff_3937000_2316000# diff_94000_5193000# diff_3847000_2257000# GND efet w=14000 l=74000
+ ad=8.49e+08 pd=270000 as=0 ps=0 
M4807 diff_94000_5193000# diff_94000_5193000# diff_3901000_2205000# GND efet w=15000 l=34000
+ ad=0 pd=0 as=1.094e+09 ps=190000 
M4808 diff_4307000_2532000# diff_4302000_2656000# diff_4276000_2780000# GND efet w=105000 l=11000
+ ad=-1.26797e+09 pd=550000 as=0 ps=0 
M4809 diff_4307000_2532000# diff_4292000_2626000# diff_4276000_2780000# GND efet w=125500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4810 diff_4251000_2644000# diff_4240000_2606000# diff_4223000_2738000# GND efet w=117000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4811 diff_3697000_2161000# diff_3687000_2150000# diff_82000_3097000# GND efet w=205000 l=10000
+ ad=-1.55197e+09 pd=476000 as=0 ps=0 
M4812 diff_3686000_2065000# diff_3670000_2092000# diff_82000_3097000# GND efet w=72500 l=10500
+ ad=1.078e+09 pd=192000 as=0 ps=0 
M4813 diff_3780000_2100000# diff_3738000_825000# diff_3697000_2161000# GND efet w=88000 l=12000
+ ad=9.72e+08 pd=212000 as=0 ps=0 
M4814 diff_3847000_2257000# diff_3694000_2724000# diff_3578000_2264000# GND efet w=88000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4815 diff_816000_2341000# diff_3921000_785000# diff_3937000_2316000# GND efet w=22000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M4816 diff_4038000_2326000# diff_4003000_2724000# diff_816000_2341000# GND efet w=22000 l=13000
+ ad=9.23e+08 pd=274000 as=0 ps=0 
M4817 diff_94000_5193000# diff_94000_5193000# diff_4056000_2221000# GND efet w=15000 l=34000
+ ad=0 pd=0 as=1.038e+09 ps=186000 
M4818 diff_4067000_2231000# diff_94000_5193000# diff_4038000_2326000# GND efet w=14500 l=74500
+ ad=-1.38197e+09 pd=484000 as=0 ps=0 
M4819 diff_94000_5193000# diff_94000_5193000# diff_4067000_2231000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4820 diff_82000_3097000# diff_3901000_2205000# diff_3847000_2257000# GND efet w=205000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4821 diff_3901000_2205000# diff_3937000_2316000# diff_82000_3097000# GND efet w=63500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4822 diff_3437000_1855000# diff_3438000_2491000# diff_1707000_1881000# GND efet w=107500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M4823 diff_3578000_1887000# diff_3566000_784000# diff_3437000_1855000# GND efet w=111000 l=12000
+ ad=-9.36967e+08 pd=708000 as=0 ps=0 
M4824 diff_3373000_1906000# diff_3353000_2408000# diff_2759000_1832000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4825 diff_3373000_1682000# diff_3353000_2408000# diff_3334000_1758000# GND efet w=22000 l=12000
+ ad=1.472e+09 pd=290000 as=7.87e+08 ps=156000 
M4826 diff_3334000_1758000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=104000
+ ad=0 pd=0 as=0 ps=0 
M4827 diff_3426000_1943000# diff_3373000_1906000# diff_82000_3097000# GND efet w=68000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4828 diff_3437000_1855000# diff_3426000_1943000# diff_82000_3097000# GND efet w=206500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4829 diff_2759000_1832000# diff_3473000_793000# diff_3437000_1855000# GND efet w=88000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4830 diff_3437000_1784000# diff_3427000_1773000# diff_82000_3097000# GND efet w=207500 l=9500
+ ad=-1.57897e+09 pd=478000 as=0 ps=0 
M4831 diff_3427000_1686000# diff_3409000_1711000# diff_82000_3097000# GND efet w=74000 l=10000
+ ad=1.009e+09 pd=186000 as=0 ps=0 
M4832 diff_3520000_1723000# diff_3473000_793000# diff_3437000_1784000# GND efet w=88000 l=12000
+ ad=1e+09 pd=214000 as=0 ps=0 
M4833 diff_1503000_1891000# diff_3595000_2394000# diff_3578000_1887000# GND efet w=122000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4834 diff_3659000_2040000# diff_3488000_2724000# diff_3633000_2077000# GND efet w=22000 l=12000
+ ad=4.07e+08 pd=86000 as=0 ps=0 
M4835 diff_3686000_2065000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=34000
+ ad=0 pd=0 as=0 ps=0 
M4836 diff_3697000_2161000# diff_94000_5193000# diff_3670000_2092000# GND efet w=14500 l=81500
+ ad=0 pd=0 as=2.8e+08 ps=94000 
M4837 diff_3697000_2161000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M4838 diff_1707000_1881000# diff_3488000_2724000# diff_3633000_1922000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=1.082e+09 ps=238000 
M4839 diff_94000_5193000# diff_94000_5193000# diff_3685000_1939000# GND efet w=15000 l=34000
+ ad=0 pd=0 as=1.147e+09 ps=194000 
M4840 diff_3697000_1854000# diff_94000_5193000# diff_3633000_1922000# GND efet w=14000 l=75000
+ ad=-3.41967e+08 pd=718000 as=0 ps=0 
M4841 diff_94000_5193000# diff_94000_5193000# diff_3697000_1854000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4842 diff_3633000_1922000# diff_3353000_2408000# diff_1503000_1891000# GND efet w=22000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M4843 diff_3397000_1682000# diff_3170000_2724000# diff_3373000_1682000# GND efet w=22000 l=12000
+ ad=3.96e+08 pd=80000 as=0 ps=0 
M4844 diff_3081000_1341000# diff_2533000_2491000# diff_3062000_1342000# GND efet w=109000 l=12000
+ ad=0 pd=0 as=1.223e+09 ps=232000 
M4845 diff_3118000_1401000# diff_3108000_1389000# diff_3081000_1341000# GND efet w=212500 l=9500
+ ad=-1.47497e+09 pd=474000 as=0 ps=0 
M4846 diff_3098000_1305000# diff_3092000_1332000# diff_3081000_1341000# GND efet w=69500 l=10500
+ ad=1.013e+09 pd=190000 as=0 ps=0 
M4847 diff_3051000_1286000# diff_2637000_2491000# diff_3028000_1286000# GND efet w=22000 l=11000
+ ad=4.4e+08 pd=84000 as=0 ps=0 
M4848 diff_816000_1210000# diff_2637000_2491000# diff_3028000_1167000# GND efet w=23000 l=11000
+ ad=0 pd=0 as=1.849e+09 ps=394000 
M4849 diff_3196000_1342000# diff_3119000_2491000# diff_3118000_1401000# GND efet w=87000 l=11000
+ ad=1.297e+09 pd=214000 as=0 ps=0 
M4850 diff_3238000_1305000# diff_3282000_1425000# diff_82000_3097000# GND efet w=91000 l=11000
+ ad=1.11103e+09 pd=880000 as=0 ps=0 
M4851 diff_94000_5193000# diff_94000_5193000# diff_2759000_1455000# GND efet w=14000 l=106000
+ ad=0 pd=0 as=0 ps=0 
M4852 diff_3427000_1686000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=34000
+ ad=0 pd=0 as=0 ps=0 
M4853 diff_3437000_1784000# diff_94000_5193000# diff_3409000_1711000# GND efet w=14500 l=80500
+ ad=0 pd=0 as=2.89e+08 ps=102000 
M4854 diff_3437000_1784000# diff_94000_5193000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4855 diff_94000_5193000# diff_94000_5193000# diff_3426000_1565000# GND efet w=14000 l=34000
+ ad=0 pd=0 as=9.93e+08 ps=182000 
M4856 diff_3437000_1477000# diff_94000_5193000# diff_3373000_1529000# GND efet w=14000 l=76000
+ ad=-4.76967e+08 pd=716000 as=1.732e+09 ps=372000 
M4857 diff_94000_5193000# diff_94000_5193000# diff_3437000_1477000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4858 diff_816000_1587000# diff_3170000_2724000# diff_3373000_1529000# GND efet w=21000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4859 diff_3557000_1710000# diff_3438000_2491000# diff_3538000_1674000# GND efet w=107000 l=12000
+ ad=1.044e+09 pd=232000 as=9.49e+08 ps=228000 
M4860 diff_3578000_1747000# diff_3566000_784000# diff_3557000_1710000# GND efet w=110000 l=12000
+ ad=1.494e+09 pd=290000 as=0 ps=0 
M4861 diff_3610000_1660000# diff_3595000_2394000# diff_3578000_1747000# GND efet w=122000 l=12000
+ ad=1.355e+09 pd=286000 as=0 ps=0 
M4862 diff_3633000_1700000# diff_3353000_2408000# diff_3610000_1660000# GND efet w=21000 l=12000
+ ad=8.12e+08 pd=156000 as=0 ps=0 
M4863 diff_3819000_2042000# diff_3801000_831000# diff_3795000_2097000# GND efet w=104000 l=12000
+ ad=1.292e+09 pd=242000 as=1.003e+09 ps=232000 
M4864 diff_3847000_2079000# diff_3829000_786000# diff_3819000_2042000# GND efet w=104500 l=11500
+ ad=1.208e+09 pd=236000 as=0 ps=0 
M4865 diff_3881000_2061000# diff_3694000_2724000# diff_3864000_2146000# GND efet w=87000 l=12000
+ ad=-1.51897e+09 pd=476000 as=8.76e+08 ps=208000 
M4866 diff_82000_3097000# diff_3901000_2171000# diff_3881000_2061000# GND efet w=206000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4867 diff_3949000_2094000# diff_3938000_2059000# diff_82000_3097000# GND efet w=65000 l=10000
+ ad=1.086e+09 pd=188000 as=0 ps=0 
M4868 diff_1707000_1881000# diff_3801000_831000# diff_3697000_1854000# GND efet w=104500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M4869 diff_3847000_1880000# diff_3829000_786000# diff_1707000_1881000# GND efet w=104500 l=11500
+ ad=-2.46967e+08 pd=716000 as=0 ps=0 
M4870 diff_3685000_1939000# diff_3633000_1922000# diff_82000_3097000# GND efet w=68500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4871 diff_3697000_1854000# diff_3685000_1939000# diff_82000_3097000# GND efet w=205000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4872 diff_3578000_1887000# diff_3738000_825000# diff_3697000_1854000# GND efet w=88000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4873 diff_4056000_2221000# diff_4038000_2326000# diff_82000_3097000# GND efet w=61500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4874 diff_4067000_2231000# diff_4056000_2221000# diff_82000_3097000# GND efet w=204500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4875 diff_816000_2341000# diff_4107000_2724000# diff_4067000_2231000# GND efet w=88000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4876 diff_4185000_2206000# diff_4162000_2432000# diff_4166000_2316000# GND efet w=87000 l=12000
+ ad=1.569e+09 pd=368000 as=9.16e+08 ps=208000 
M4877 diff_4067000_2161000# diff_4056000_2150000# diff_82000_3097000# GND efet w=206500 l=9500
+ ad=-1.39497e+09 pd=476000 as=0 ps=0 
M4878 diff_82000_3097000# diff_4037000_2050000# diff_4057000_2112000# GND efet w=62500 l=10500
+ ad=0 pd=0 as=9.89e+08 ps=180000 
M4879 diff_4150000_2101000# diff_4107000_2724000# diff_4067000_2161000# GND efet w=88000 l=12000
+ ad=1.04e+09 pd=212000 as=0 ps=0 
M4880 diff_4204000_2168000# diff_4192000_1025000# diff_4185000_2206000# GND efet w=108000 l=12000
+ ad=-1.23697e+09 pd=464000 as=0 ps=0 
M4881 diff_4204000_2168000# diff_4192000_1025000# diff_4184000_2136000# GND efet w=106000 l=12000
+ ad=0 pd=0 as=1.579e+09 ps=364000 
M4882 diff_4237000_2412000# diff_4154000_2675000# diff_4204000_2168000# GND efet w=91000 l=12000
+ ad=-2.66967e+08 pd=676000 as=0 ps=0 
M4883 diff_3881000_2061000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M4884 diff_3938000_2059000# diff_94000_5193000# diff_3881000_2061000# GND efet w=14500 l=80500
+ ad=8.93e+08 pd=248000 as=0 ps=0 
M4885 diff_3949000_2094000# diff_94000_5193000# diff_94000_5193000# GND efet w=15000 l=34000
+ ad=0 pd=0 as=0 ps=0 
M4886 diff_4005000_2050000# diff_3921000_785000# diff_3938000_2059000# GND efet w=22000 l=12000
+ ad=4.4e+08 pd=84000 as=0 ps=0 
M4887 diff_4037000_2050000# diff_4003000_2724000# diff_4005000_2050000# GND efet w=22000 l=12000
+ ad=9.33e+08 pd=232000 as=0 ps=0 
M4888 diff_3937000_1939000# diff_94000_5193000# diff_3847000_1880000# GND efet w=14000 l=76000
+ ad=8.69e+08 pd=272000 as=0 ps=0 
M4889 diff_94000_5193000# diff_94000_5193000# diff_3847000_1880000# GND efet w=13000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4890 diff_94000_5193000# diff_94000_5193000# diff_3901000_1828000# GND efet w=15000 l=34000
+ ad=0 pd=0 as=1.104e+09 ps=190000 
M4891 diff_4057000_2112000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=34000
+ ad=0 pd=0 as=0 ps=0 
M4892 diff_4067000_2161000# diff_94000_5193000# diff_4037000_2050000# GND efet w=14000 l=81000
+ ad=0 pd=0 as=0 ps=0 
M4893 diff_4067000_2161000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M4894 diff_1707000_1881000# diff_3921000_785000# diff_3937000_1939000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4895 diff_4037000_1949000# diff_4003000_2724000# diff_1707000_1881000# GND efet w=22000 l=12000
+ ad=9.18e+08 pd=250000 as=0 ps=0 
M4896 diff_94000_5193000# diff_94000_5193000# diff_4056000_1844000# GND efet w=15000 l=34000
+ ad=0 pd=0 as=1.046e+09 ps=186000 
M4897 diff_4067000_1854000# diff_94000_5193000# diff_4037000_1949000# GND efet w=14000 l=76000
+ ad=-1.34797e+09 pd=484000 as=0 ps=0 
M4898 diff_4184000_2136000# diff_4162000_2432000# diff_4165000_2061000# GND efet w=88000 l=12000
+ ad=0 pd=0 as=8.96e+08 ps=212000 
M4899 diff_94000_5193000# diff_94000_5193000# diff_4067000_1854000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4900 diff_3697000_1784000# diff_3687000_1773000# diff_82000_3097000# GND efet w=206000 l=10000
+ ad=-1.51997e+09 pd=480000 as=0 ps=0 
M4901 diff_3686000_1688000# diff_3670000_1715000# diff_82000_3097000# GND efet w=72500 l=10500
+ ad=1.091e+09 pd=194000 as=0 ps=0 
M4902 diff_3780000_1723000# diff_3738000_825000# diff_3697000_1784000# GND efet w=88000 l=12000
+ ad=9.72e+08 pd=212000 as=0 ps=0 
M4903 diff_3847000_1880000# diff_3694000_2724000# diff_3578000_1887000# GND efet w=88000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4904 diff_82000_3097000# diff_3901000_1828000# diff_3847000_1880000# GND efet w=206000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4905 diff_3901000_1828000# diff_3937000_1939000# diff_82000_3097000# GND efet w=64500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4906 diff_3437000_1477000# diff_3438000_2491000# diff_816000_1587000# GND efet w=108000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4907 diff_3578000_1510000# diff_3566000_784000# diff_3437000_1477000# GND efet w=111000 l=12000
+ ad=-9.16967e+08 pd=710000 as=0 ps=0 
M4908 diff_3238000_1305000# diff_2892000_2724000# diff_3212000_1340000# GND efet w=88000 l=13000
+ ad=0 pd=0 as=9.15e+08 ps=210000 
M4909 diff_3098000_1305000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=33000
+ ad=0 pd=0 as=0 ps=0 
M4910 diff_3118000_1401000# diff_94000_5193000# diff_3092000_1332000# GND efet w=14000 l=81000
+ ad=0 pd=0 as=1.97e+08 ps=66000 
M4911 diff_3118000_1401000# diff_94000_5193000# diff_94000_5193000# GND efet w=13000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4912 diff_94000_5193000# diff_94000_5193000# diff_3098000_1188000# GND efet w=14000 l=32000
+ ad=0 pd=0 as=1.065e+09 ps=192000 
M4913 diff_3118000_1088000# diff_94000_5193000# diff_3028000_1167000# GND efet w=14000 l=76000
+ ad=-3.90967e+08 pd=700000 as=0 ps=0 
M4914 diff_94000_5193000# diff_94000_5193000# diff_3118000_1088000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4915 diff_847000_1210000# diff_2995000_2724000# diff_2914000_1187000# GND efet w=21000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M4916 diff_3028000_1167000# diff_2995000_2724000# diff_2759000_1078000# GND efet w=21000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4917 diff_3028000_909000# diff_2995000_2724000# diff_3005000_1018000# GND efet w=21000 l=12000
+ ad=1.608e+09 pd=310000 as=3.57e+08 ps=76000 
M4918 diff_3011000_980000# diff_2995000_2724000# diff_2987000_946000# GND efet w=21000 l=11000
+ ad=3.99e+08 pd=80000 as=1.192e+09 ps=230000 
M4919 diff_2865000_1028000# diff_2860000_903000# diff_2860000_876000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=5.47e+08 ps=96000 
M4920 diff_2914000_928000# diff_2860000_903000# diff_2865000_1028000# GND efet w=14500 l=83500
+ ad=1.76e+08 pd=76000 as=0 ps=0 
M4921 diff_2930000_970000# diff_2860000_903000# diff_2937000_871000# GND efet w=14000 l=33000
+ ad=0 pd=0 as=4.77e+08 ps=90000 
M4922 diff_2987000_946000# diff_2938000_823000# diff_2962000_909000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=3.78e+08 ps=78000 
M4923 diff_3081000_1137000# diff_2533000_2491000# diff_2759000_1078000# GND efet w=108500 l=11500
+ ad=-1.49993e+09 pd=1.008e+06 as=0 ps=0 
M4924 diff_3098000_1188000# diff_3028000_1167000# diff_3081000_1137000# GND efet w=64500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4925 diff_3373000_1529000# diff_3353000_2408000# diff_2759000_1455000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4926 diff_3373000_1305000# diff_3353000_2408000# diff_3334000_1381000# GND efet w=22000 l=12000
+ ad=1.473e+09 pd=290000 as=7.7e+08 ps=156000 
M4927 diff_3334000_1381000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=104000
+ ad=0 pd=0 as=0 ps=0 
M4928 diff_3426000_1565000# diff_3373000_1529000# diff_82000_3097000# GND efet w=67000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4929 diff_3437000_1477000# diff_3426000_1565000# diff_82000_3097000# GND efet w=205500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4930 diff_2759000_1455000# diff_3473000_793000# diff_3437000_1477000# GND efet w=88000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4931 diff_3437000_1406000# diff_3427000_1395000# diff_82000_3097000# GND efet w=206500 l=9500
+ ad=-1.57797e+09 pd=476000 as=0 ps=0 
M4932 diff_3427000_1308000# diff_3409000_1334000# diff_82000_3097000# GND efet w=72000 l=10000
+ ad=9.86e+08 pd=184000 as=0 ps=0 
M4933 diff_3520000_1345000# diff_3473000_793000# diff_3437000_1406000# GND efet w=88000 l=12000
+ ad=9.94e+08 pd=214000 as=0 ps=0 
M4934 diff_847000_1587000# diff_3595000_2394000# diff_3578000_1510000# GND efet w=122000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4935 diff_3659000_1662000# diff_3488000_2724000# diff_3633000_1700000# GND efet w=22000 l=12000
+ ad=4.08e+08 pd=86000 as=0 ps=0 
M4936 diff_3686000_1688000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=34000
+ ad=0 pd=0 as=0 ps=0 
M4937 diff_3697000_1784000# diff_94000_5193000# diff_3670000_1715000# GND efet w=14500 l=80500
+ ad=0 pd=0 as=2.95e+08 ps=96000 
M4938 diff_3697000_1784000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4939 diff_816000_1587000# diff_3488000_2724000# diff_3633000_1545000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=1.073e+09 ps=238000 
M4940 diff_94000_5193000# diff_94000_5193000# diff_3685000_1561000# GND efet w=15000 l=34000
+ ad=0 pd=0 as=1.122e+09 ps=192000 
M4941 diff_3697000_1476000# diff_94000_5193000# diff_3633000_1545000# GND efet w=14000 l=76000
+ ad=-4.08967e+08 pd=712000 as=0 ps=0 
M4942 diff_94000_5193000# diff_94000_5193000# diff_3697000_1476000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4943 diff_3633000_1545000# diff_3353000_2408000# diff_847000_1587000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4944 diff_3397000_1305000# diff_3170000_2724000# diff_3373000_1305000# GND efet w=21000 l=12000
+ ad=3.78e+08 pd=78000 as=0 ps=0 
M4945 diff_3118000_1088000# diff_3098000_1188000# diff_3081000_1137000# GND efet w=214500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4946 diff_2759000_1078000# diff_3119000_2491000# diff_3118000_1088000# GND efet w=88000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4947 diff_816000_1210000# diff_2892000_2724000# diff_3118000_1088000# GND efet w=88000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4948 diff_3081000_1137000# diff_2533000_2491000# diff_3062000_965000# GND efet w=108500 l=12500
+ ad=0 pd=0 as=1.193e+09 ps=232000 
M4949 diff_3118000_1024000# diff_3108000_1012000# diff_3081000_1137000# GND efet w=215500 l=9500
+ ad=-1.53697e+09 pd=476000 as=0 ps=0 
M4950 diff_3098000_928000# diff_3092000_955000# diff_3081000_1137000# GND efet w=69500 l=10500
+ ad=1.052e+09 pd=190000 as=0 ps=0 
M4951 diff_3052000_908000# diff_2637000_2491000# diff_3028000_909000# GND efet w=23000 l=12000
+ ad=4.35e+08 pd=84000 as=0 ps=0 
M4952 diff_3196000_965000# diff_3119000_2491000# diff_3118000_1024000# GND efet w=88000 l=11000
+ ad=1.31e+09 pd=216000 as=0 ps=0 
M4953 diff_3238000_927000# diff_2892000_2724000# diff_3212000_963000# GND efet w=88000 l=12000
+ ad=1.49e+09 pd=286000 as=1.002e+09 ps=212000 
M4954 diff_3098000_928000# diff_3092000_894000# diff_3091000_870000# GND efet w=14000 l=34000
+ ad=0 pd=0 as=4.89e+08 ps=90000 
M4955 diff_3118000_1024000# diff_3092000_894000# diff_3092000_955000# GND efet w=14000 l=83000
+ ad=0 pd=0 as=2.18e+08 ps=72000 
M4956 diff_3118000_1024000# diff_3092000_894000# diff_3181000_876000# GND efet w=13000 l=25000
+ ad=0 pd=0 as=5.19e+08 ps=94000 
M4957 diff_2744000_764000# diff_2733000_743000# diff_2712000_821000# GND efet w=73000 l=11000
+ ad=1.46e+09 pd=186000 as=0 ps=0 
M4958 diff_2776000_764000# diff_2733000_743000# diff_2744000_764000# GND efet w=73000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4959 diff_2838000_765000# diff_2827000_743000# diff_2582000_2724000# GND efet w=72000 l=11000
+ ad=1.44e+09 pd=184000 as=0 ps=0 
M4960 diff_2842000_1949000# diff_2827000_743000# diff_2838000_765000# GND efet w=72000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4961 diff_2970000_767000# diff_2959000_743000# diff_2938000_823000# GND efet w=73000 l=11000
+ ad=1.533e+09 pd=188000 as=0 ps=0 
M4962 diff_2995000_2724000# diff_2959000_743000# diff_2970000_767000# GND efet w=73000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4963 diff_3065000_767000# diff_3054000_743000# diff_2637000_2491000# GND efet w=73000 l=11000
+ ad=1.46e+09 pd=186000 as=0 ps=0 
M4964 diff_2533000_2491000# diff_3054000_743000# diff_3065000_767000# GND efet w=73000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4965 diff_3183000_765000# diff_3171000_743000# diff_3119000_2491000# GND efet w=73000 l=12000
+ ad=1.46e+09 pd=186000 as=0 ps=0 
M4966 diff_2892000_2724000# diff_3171000_743000# diff_3183000_765000# GND efet w=73000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4967 diff_2759000_1078000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=105000
+ ad=0 pd=0 as=0 ps=0 
M4968 diff_3427000_1308000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=34000
+ ad=0 pd=0 as=0 ps=0 
M4969 diff_3437000_1406000# diff_94000_5193000# diff_3409000_1334000# GND efet w=14500 l=81500
+ ad=0 pd=0 as=2.75e+08 ps=100000 
M4970 diff_3437000_1406000# diff_94000_5193000# diff_94000_5193000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4971 diff_3426000_1188000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=35000
+ ad=9.91e+08 pd=182000 as=0 ps=0 
M4972 diff_3437000_1100000# diff_94000_5193000# diff_3373000_1152000# GND efet w=14000 l=76000
+ ad=-3.17967e+08 pd=720000 as=1.744e+09 ps=374000 
M4973 diff_94000_5193000# diff_94000_5193000# diff_3437000_1100000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4974 diff_816000_1210000# diff_3170000_2724000# diff_3373000_1152000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4975 diff_3557000_1333000# diff_3438000_2491000# diff_3538000_1297000# GND efet w=106500 l=11500
+ ad=1.094e+09 pd=232000 as=9.5e+08 ps=228000 
M4976 diff_3578000_1369000# diff_3566000_784000# diff_3557000_1333000# GND efet w=110000 l=12000
+ ad=1.505e+09 pd=290000 as=0 ps=0 
M4977 diff_3610000_1283000# diff_3595000_2394000# diff_3578000_1369000# GND efet w=122000 l=12000
+ ad=1.363e+09 pd=286000 as=0 ps=0 
M4978 diff_3633000_1323000# diff_3353000_2408000# diff_3610000_1283000# GND efet w=21000 l=12000
+ ad=8.13e+08 pd=156000 as=0 ps=0 
M4979 diff_3819000_1665000# diff_3801000_831000# diff_3795000_1720000# GND efet w=104500 l=11500
+ ad=1.279e+09 pd=242000 as=1.07e+09 ps=234000 
M4980 diff_3847000_1701000# diff_3829000_786000# diff_3819000_1665000# GND efet w=104500 l=11500
+ ad=1.205e+09 pd=236000 as=0 ps=0 
M4981 diff_3881000_1684000# diff_3694000_2724000# diff_3864000_1769000# GND efet w=88000 l=12000
+ ad=-1.49897e+09 pd=480000 as=8.84e+08 ps=210000 
M4982 diff_82000_3097000# diff_3901000_1794000# diff_3881000_1684000# GND efet w=206000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4983 diff_3949000_1717000# diff_3938000_1681000# diff_82000_3097000# GND efet w=65000 l=10000
+ ad=1.102e+09 pd=190000 as=0 ps=0 
M4984 diff_816000_1587000# diff_3801000_831000# diff_3697000_1476000# GND efet w=104000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4985 diff_3847000_1503000# diff_3829000_786000# diff_816000_1587000# GND efet w=104500 l=11500
+ ad=-2.62967e+08 pd=712000 as=0 ps=0 
M4986 diff_3685000_1561000# diff_3633000_1545000# diff_82000_3097000# GND efet w=67500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4987 diff_3697000_1476000# diff_3685000_1561000# diff_82000_3097000# GND efet w=205000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4988 diff_3578000_1510000# diff_3738000_825000# diff_3697000_1476000# GND efet w=88000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4989 diff_4056000_1844000# diff_4037000_1949000# diff_82000_3097000# GND efet w=62500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4990 diff_4067000_1854000# diff_4056000_1844000# diff_82000_3097000# GND efet w=205500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4991 diff_1707000_1881000# diff_4107000_2724000# diff_4067000_1854000# GND efet w=88000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4992 diff_4185000_1829000# diff_4162000_2432000# diff_4166000_1940000# GND efet w=88000 l=12000
+ ad=1.51e+09 pd=368000 as=9.23e+08 ps=210000 
M4993 diff_4461000_2970000# diff_4461000_2970000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M4994 diff_82000_3097000# diff_4494000_3313000# diff_4516000_3009000# GND efet w=74000 l=10000
+ ad=0 pd=0 as=1.178e+09 ps=274000 
M4995 diff_4592000_3171000# diff_4516000_3009000# diff_82000_3097000# GND efet w=66000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4996 diff_82000_3097000# diff_4592000_3171000# diff_4655000_3019000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=5.55033e+08 ps=938000 
M4997 diff_4655000_3019000# diff_859000_2986000# diff_82000_3097000# GND efet w=116000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4998 diff_82000_3097000# diff_905000_3225000# diff_4655000_3019000# GND efet w=115500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4999 diff_94000_5193000# diff_4592000_3171000# diff_4592000_3171000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M5000 diff_4516000_3009000# diff_4516000_3009000# diff_94000_5193000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M5001 diff_4655000_3019000# diff_4655000_3019000# diff_94000_5193000# GND efet w=15000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M5002 diff_4715000_3242000# diff_71000_4514000# diff_4842000_3180000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=5.78e+08 ps=148000 
M5003 diff_4813000_3334000# diff_71000_4514000# diff_4864000_3204000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=4.48e+08 ps=128000 
M5004 diff_82000_3097000# diff_4778000_3197000# diff_4776000_2950000# GND efet w=74500 l=10500
+ ad=0 pd=0 as=-9.12967e+08 ps=668000 
M5005 diff_4776000_2950000# diff_3568000_3529000# diff_82000_3097000# GND efet w=64000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5006 diff_82000_3097000# diff_4842000_3180000# diff_4842000_3066000# GND efet w=65000 l=10000
+ ad=0 pd=0 as=7.87033e+08 ps=882000 
M5007 diff_4842000_3066000# diff_4864000_3204000# diff_82000_3097000# GND efet w=65000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5008 diff_4805000_4500000# diff_71000_4514000# diff_4922000_2910000# GND efet w=13000 l=13000
+ ad=0 pd=0 as=3.65e+08 ps=118000 
M5009 diff_94000_5193000# diff_4776000_2950000# diff_4776000_2950000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M5010 diff_4904000_3016000# diff_67000_5287000# diff_3238000_1305000# GND efet w=14000 l=13000
+ ad=7.23e+08 pd=132000 as=0 ps=0 
M5011 diff_4967000_3078000# diff_4904000_3016000# diff_82000_3097000# GND efet w=133000 l=11000
+ ad=9.31e+08 pd=280000 as=0 ps=0 
M5012 diff_4984000_2921000# diff_4926000_3399000# diff_4967000_3078000# GND efet w=133000 l=10000
+ ad=8.06033e+08 pd=886000 as=0 ps=0 
M5013 diff_5438000_3443000# diff_5356000_3321000# diff_82000_3097000# GND efet w=99000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5014 diff_5919000_3448000# diff_5919000_3448000# diff_94000_5193000# GND efet w=14000 l=39000
+ ad=2.078e+09 pd=500000 as=0 ps=0 
M5015 diff_3253000_2508000# diff_71000_4514000# diff_5431000_3450000# GND efet w=15000 l=13000
+ ad=1.451e+09 pd=300000 as=3.38e+08 ps=86000 
M5016 diff_6005000_3448000# diff_5067000_4961000# diff_5919000_3448000# GND efet w=87000 l=11000
+ ad=6.09e+08 pd=188000 as=0 ps=0 
M5017 diff_94000_5193000# diff_6111000_3387000# diff_6111000_3387000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M5018 diff_6159000_3458000# diff_5919000_3448000# diff_6111000_3387000# GND efet w=92500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5019 diff_94000_5193000# diff_3253000_2508000# diff_3253000_2508000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M5020 diff_3253000_2508000# diff_5577000_3392000# diff_82000_3097000# GND efet w=74000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5021 diff_6005000_3448000# diff_5097000_4893000# diff_82000_3097000# GND efet w=87000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5022 diff_4882000_4961000# diff_71000_4514000# diff_5406000_3339000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=5.9e+08 ps=142000 
M5023 diff_5530000_3345000# diff_4264000_3069000# diff_82000_3097000# GND efet w=95000 l=10000
+ ad=7.93e+08 pd=224000 as=0 ps=0 
M5024 diff_5530000_3345000# diff_5406000_3339000# diff_5047000_3692000# GND efet w=105000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5025 diff_82000_3097000# diff_5406000_3339000# diff_5356000_3321000# GND efet w=50000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5026 diff_6075000_3941000# diff_5038000_4961000# diff_82000_3097000# GND efet w=44000 l=11000
+ ad=-1.49397e+09 pd=554000 as=0 ps=0 
M5027 diff_6121000_3398000# diff_6111000_3387000# diff_82000_3097000# GND efet w=105500 l=10500
+ ad=1.856e+09 pd=370000 as=0 ps=0 
M5028 diff_82000_3097000# diff_5695000_3193000# diff_6121000_3398000# GND efet w=92000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5029 diff_6075000_3941000# diff_6179000_3355000# diff_6121000_3398000# GND efet w=90000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5030 diff_94000_5193000# diff_6075000_3941000# diff_6075000_3941000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M5031 diff_82000_3097000# diff_5008000_4961000# diff_5695000_3193000# GND efet w=68000 l=11000
+ ad=0 pd=0 as=1.765e+09 ps=402000 
M5032 diff_82000_3097000# diff_5468000_3308000# diff_5356000_3321000# GND efet w=46000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5033 diff_5356000_3321000# diff_5356000_3321000# diff_94000_5193000# GND efet w=14000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M5034 diff_5047000_3692000# diff_5468000_3308000# diff_82000_3097000# GND efet w=44000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5035 diff_5468000_3308000# diff_71000_4514000# diff_64000_4219000# GND efet w=14000 l=14000
+ ad=2.57e+08 pd=74000 as=0 ps=0 
M5036 diff_5083000_3005000# diff_67000_5287000# diff_4984000_2921000# GND efet w=14000 l=14000
+ ad=6.18e+08 pd=144000 as=0 ps=0 
M5037 diff_94000_5193000# diff_4264000_3069000# diff_4264000_3069000# GND efet w=15000 l=25000
+ ad=0 pd=0 as=1.812e+09 ps=358000 
M5038 diff_4264000_3069000# diff_5575000_3240000# diff_82000_3097000# GND efet w=80500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5039 diff_5695000_3193000# diff_71000_4514000# diff_5575000_3240000# GND efet w=14500 l=13500
+ ad=0 pd=0 as=2.42e+08 ps=72000 
M5040 diff_94000_5193000# diff_4842000_3066000# diff_4842000_3066000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M5041 diff_82000_3097000# diff_4922000_2910000# diff_4911000_2899000# GND efet w=144000 l=9000
+ ad=0 pd=0 as=-1.73097e+09 ps=520000 
M5042 diff_4984000_2921000# diff_4974000_2909000# diff_4911000_2899000# GND efet w=144000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5043 diff_5011000_3005000# diff_4870000_3350000# diff_4984000_2921000# GND efet w=131000 l=10000
+ ad=9.17e+08 pd=276000 as=0 ps=0 
M5044 diff_82000_3097000# diff_5018000_2992000# diff_5011000_3005000# GND efet w=131000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5045 diff_3320000_2526000# diff_71000_4514000# diff_5018000_2992000# GND efet w=14000 l=12000
+ ad=2.062e+09 pd=392000 as=3.85e+08 ps=126000 
M5046 diff_82000_3097000# diff_5083000_3005000# diff_3320000_2526000# GND efet w=94500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5047 diff_5695000_3193000# diff_5695000_3193000# diff_94000_5193000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M5048 diff_94000_5193000# diff_6179000_3355000# diff_6179000_3355000# GND efet w=13500 l=37500
+ ad=0 pd=0 as=1.671e+09 ps=350000 
M5049 diff_6179000_3355000# diff_5695000_3193000# diff_6268000_3301000# GND efet w=133000 l=11000
+ ad=0 pd=0 as=9.31e+08 ps=280000 
M5050 diff_6268000_3301000# diff_5067000_4961000# diff_6268000_3283000# GND efet w=133000 l=10000
+ ad=0 pd=0 as=1.064e+09 ps=282000 
M5051 diff_6268000_3283000# diff_6251000_3156000# diff_82000_3097000# GND efet w=133000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5052 diff_94000_5193000# diff_4984000_2921000# diff_4984000_2921000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M5053 diff_94000_5193000# diff_3320000_2526000# diff_3320000_2526000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M5054 diff_5203000_3036000# diff_71000_4514000# diff_82000_3097000# GND efet w=274000 l=11000
+ ad=1.22003e+09 pd=856000 as=0 ps=0 
M5055 diff_82000_3097000# diff_5213000_3049000# diff_5203000_3036000# GND efet w=272000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5056 diff_82000_3097000# diff_5256000_3172000# diff_5213000_3049000# GND efet w=127500 l=10500
+ ad=0 pd=0 as=-2.12497e+09 ps=342000 
M5057 diff_5213000_3049000# diff_5213000_3049000# diff_94000_5193000# GND efet w=15000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5058 diff_4357000_3757000# diff_4382000_2804000# diff_4390000_2777000# GND efet w=21000 l=16000
+ ad=0 pd=0 as=9.67e+08 ps=156000 
M5059 diff_4461000_2970000# diff_4382000_2804000# diff_4493000_2777000# GND efet w=21500 l=15500
+ ad=0 pd=0 as=9.67e+08 ps=156000 
M5060 diff_4414000_3773000# diff_4382000_2804000# diff_4442000_2777000# GND efet w=22000 l=15000
+ ad=0 pd=0 as=9.94e+08 ps=158000 
M5061 diff_4461000_3007000# diff_4382000_2804000# diff_4545000_2777000# GND efet w=21000 l=15000
+ ad=0 pd=0 as=9.57e+08 ps=156000 
M5062 diff_4696000_3225000# diff_4734000_2812000# diff_4688000_2591000# GND efet w=14000 l=10000
+ ad=0 pd=0 as=1.057e+09 ps=156000 
M5063 diff_4623000_2773000# diff_4601000_2751000# diff_4601000_2751000# GND efet w=20000 l=10000
+ ad=4.78e+08 pd=100000 as=5.39033e+08 ps=980000 
M5064 diff_4373000_832000# diff_4390000_2777000# diff_4377000_2527000# GND efet w=247000 l=10000
+ ad=3.53033e+08 pd=958000 as=-5.04967e+08 ps=516000 
M5065 diff_4424000_2748000# diff_4373000_832000# diff_4373000_832000# GND efet w=20000 l=9000
+ ad=4.6e+08 pd=86000 as=0 ps=0 
M5066 diff_4416000_951000# diff_4416000_951000# diff_4424000_2748000# GND efet w=20000 l=9000
+ ad=1.40327e+07 pd=898000 as=0 ps=0 
M5067 diff_4425000_2536000# diff_4414000_2527000# diff_4373000_832000# GND efet w=205000 l=11000
+ ad=-3.89967e+08 pd=440000 as=0 ps=0 
M5068 diff_4416000_951000# diff_4414000_2527000# diff_4425000_2536000# GND efet w=205000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5069 diff_4477000_2552000# diff_4442000_2777000# diff_4416000_951000# GND efet w=246000 l=10000
+ ad=2.40327e+07 pd=522000 as=0 ps=0 
M5070 diff_4497000_2491000# diff_4493000_2777000# diff_4477000_2552000# GND efet w=247000 l=10000
+ ad=-9.09673e+07 pd=898000 as=0 ps=0 
M5071 diff_4528000_2748000# diff_4497000_2491000# diff_4497000_2491000# GND efet w=20000 l=10000
+ ad=4.4e+08 pd=84000 as=0 ps=0 
M5072 diff_4547000_2724000# diff_4547000_2724000# diff_4528000_2748000# GND efet w=20000 l=10000
+ ad=1.14033e+08 pd=898000 as=0 ps=0 
M5073 diff_4528000_2536000# diff_4517000_2527000# diff_4497000_2491000# GND efet w=206000 l=10000
+ ad=-2.19967e+08 pd=442000 as=0 ps=0 
M5074 diff_4547000_2724000# diff_4517000_2527000# diff_4528000_2536000# GND efet w=205500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5075 diff_4580000_2552000# diff_4545000_2777000# diff_4547000_2724000# GND efet w=246500 l=10500
+ ad=-3.19673e+07 pd=520000 as=0 ps=0 
M5076 diff_4642000_2735000# diff_4642000_2735000# diff_4623000_2773000# GND efet w=26000 l=10000
+ ad=1.60903e+09 pd=1.026e+06 as=0 ps=0 
M5077 diff_4715000_3242000# diff_4734000_2812000# diff_4784000_2782000# GND efet w=15000 l=11000
+ ad=0 pd=0 as=1.157e+09 ps=186000 
M5078 diff_4776000_2950000# diff_4825000_2753000# diff_4882000_2652000# GND efet w=15000 l=10000
+ ad=0 pd=0 as=1.006e+09 ps=170000 
M5079 diff_4628000_2513000# diff_4617000_2492000# diff_4601000_2751000# GND efet w=202500 l=10500
+ ad=-6.81967e+08 pd=436000 as=0 ps=0 
M5080 diff_4264000_1839000# diff_4223000_2738000# diff_4199000_2721000# GND efet w=89000 l=12000
+ ad=-9.30935e+08 pd=748000 as=0 ps=0 
M5081 diff_4067000_1784000# diff_4056000_1773000# diff_82000_3097000# GND efet w=205500 l=9500
+ ad=-1.38597e+09 pd=478000 as=0 ps=0 
M5082 diff_82000_3097000# diff_4038000_1673000# diff_4057000_1734000# GND efet w=62500 l=10500
+ ad=0 pd=0 as=1.005e+09 ps=182000 
M5083 diff_4149000_1723000# diff_4107000_2724000# diff_4067000_1784000# GND efet w=88000 l=11000
+ ad=1.136e+09 pd=214000 as=0 ps=0 
M5084 diff_4204000_1790000# diff_4192000_1025000# diff_4185000_1829000# GND efet w=107000 l=12000
+ ad=-1.25297e+09 pd=462000 as=0 ps=0 
M5085 diff_4235000_1746000# diff_4225000_1879000# diff_4204000_1790000# GND efet w=77000 l=10000
+ ad=-1.70497e+09 pd=406000 as=0 ps=0 
M5086 diff_4264000_1839000# diff_4251000_1918000# diff_4235000_1746000# GND efet w=74000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5087 diff_4204000_1790000# diff_4192000_1025000# diff_4184000_1760000# GND efet w=107500 l=12500
+ ad=0 pd=0 as=1.598e+09 ps=366000 
M5088 diff_3881000_1684000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M5089 diff_3938000_1681000# diff_94000_5193000# diff_3881000_1684000# GND efet w=14500 l=79500
+ ad=8.86e+08 pd=248000 as=0 ps=0 
M5090 diff_3949000_1717000# diff_94000_5193000# diff_94000_5193000# GND efet w=15000 l=33000
+ ad=0 pd=0 as=0 ps=0 
M5091 diff_4005000_1673000# diff_3921000_785000# diff_3938000_1681000# GND efet w=22000 l=13000
+ ad=4.4e+08 pd=84000 as=0 ps=0 
M5092 diff_4038000_1673000# diff_4003000_2724000# diff_4005000_1673000# GND efet w=22000 l=13000
+ ad=9.25e+08 pd=232000 as=0 ps=0 
M5093 diff_3937000_1562000# diff_94000_5193000# diff_3847000_1503000# GND efet w=14000 l=77000
+ ad=8.52e+08 pd=264000 as=0 ps=0 
M5094 diff_94000_5193000# diff_94000_5193000# diff_3847000_1503000# GND efet w=13000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M5095 diff_94000_5193000# diff_94000_5193000# diff_3901000_1450000# GND efet w=15000 l=34000
+ ad=0 pd=0 as=1.076e+09 ps=188000 
M5096 diff_4057000_1734000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=33000
+ ad=0 pd=0 as=0 ps=0 
M5097 diff_4067000_1784000# diff_94000_5193000# diff_4038000_1673000# GND efet w=14000 l=80000
+ ad=0 pd=0 as=0 ps=0 
M5098 diff_4067000_1784000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M5099 diff_4067000_1476000# diff_94000_5193000# diff_4038000_1572000# GND efet w=14000 l=77000
+ ad=-1.36697e+09 pd=480000 as=9.01e+08 ps=244000 
M5100 diff_816000_1587000# diff_3921000_785000# diff_3937000_1562000# GND efet w=22000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M5101 diff_4038000_1572000# diff_4003000_2724000# diff_816000_1587000# GND efet w=22000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M5102 diff_94000_5193000# diff_94000_5193000# diff_4056000_1466000# GND efet w=15000 l=34000
+ ad=0 pd=0 as=1.019e+09 ps=184000 
M5103 diff_4184000_1760000# diff_4162000_2432000# diff_4165000_1685000# GND efet w=89000 l=12000
+ ad=0 pd=0 as=9.05e+08 ps=214000 
M5104 diff_4225000_1648000# diff_4239000_1722000# diff_4235000_1746000# GND efet w=73000 l=10000
+ ad=-1.86397e+09 pd=406000 as=0 ps=0 
M5105 diff_94000_5193000# diff_94000_5193000# diff_4067000_1476000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M5106 diff_3697000_1406000# diff_3687000_1396000# diff_82000_3097000# GND efet w=206000 l=10000
+ ad=-1.51997e+09 pd=478000 as=0 ps=0 
M5107 diff_3686000_1310000# diff_3670000_1337000# diff_82000_3097000# GND efet w=72500 l=10500
+ ad=1.095e+09 pd=194000 as=0 ps=0 
M5108 diff_3780000_1346000# diff_3738000_825000# diff_3697000_1406000# GND efet w=88000 l=12000
+ ad=9.79e+08 pd=212000 as=0 ps=0 
M5109 diff_3847000_1503000# diff_3694000_2724000# diff_3578000_1510000# GND efet w=88000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5110 diff_82000_3097000# diff_3901000_1450000# diff_3847000_1503000# GND efet w=206000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5111 diff_3901000_1450000# diff_3937000_1562000# diff_82000_3097000# GND efet w=64000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5112 diff_3437000_1100000# diff_3438000_2491000# diff_816000_1210000# GND efet w=107500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M5113 diff_3578000_1133000# diff_3566000_784000# diff_3437000_1100000# GND efet w=111000 l=12000
+ ad=-9.25967e+08 pd=710000 as=0 ps=0 
M5114 diff_3373000_1152000# diff_3353000_2408000# diff_2759000_1078000# GND efet w=22000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5115 diff_3373000_928000# diff_3353000_2408000# diff_3334000_1004000# GND efet w=22000 l=11000
+ ad=1.488e+09 pd=292000 as=7.7e+08 ps=156000 
M5116 diff_3334000_1004000# diff_3323000_873000# diff_3323000_873000# GND efet w=14000 l=105000
+ ad=0 pd=0 as=5.94e+08 ps=124000 
M5117 diff_3426000_1188000# diff_3373000_1152000# diff_82000_3097000# GND efet w=66000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5118 diff_3437000_1100000# diff_3426000_1188000# diff_82000_3097000# GND efet w=206500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5119 diff_2759000_1078000# diff_3473000_793000# diff_3437000_1100000# GND efet w=88000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5120 diff_3437000_1029000# diff_3427000_1018000# diff_82000_3097000# GND efet w=207500 l=9500
+ ad=-1.47497e+09 pd=470000 as=0 ps=0 
M5121 diff_3427000_934000# diff_3409000_959000# diff_82000_3097000# GND efet w=74000 l=10000
+ ad=9.76e+08 pd=182000 as=0 ps=0 
M5122 diff_3520000_968000# diff_3473000_793000# diff_3437000_1029000# GND efet w=88000 l=11000
+ ad=1e+09 pd=214000 as=0 ps=0 
M5123 diff_847000_1210000# diff_3595000_2394000# diff_3578000_1133000# GND efet w=122000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5124 diff_3659000_1285000# diff_3488000_2724000# diff_3633000_1323000# GND efet w=23000 l=12000
+ ad=4.28e+08 pd=88000 as=0 ps=0 
M5125 diff_3686000_1310000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=34000
+ ad=0 pd=0 as=0 ps=0 
M5126 diff_3697000_1406000# diff_94000_5193000# diff_3670000_1337000# GND efet w=14500 l=80500
+ ad=0 pd=0 as=2.86e+08 ps=98000 
M5127 diff_3697000_1406000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M5128 diff_816000_1210000# diff_3488000_2724000# diff_3633000_1168000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=1.073e+09 ps=238000 
M5129 diff_94000_5193000# diff_94000_5193000# diff_3685000_1184000# GND efet w=15000 l=35000
+ ad=0 pd=0 as=1.12e+09 ps=192000 
M5130 diff_3697000_1099000# diff_94000_5193000# diff_3633000_1168000# GND efet w=14000 l=76000
+ ad=-3.16967e+08 pd=714000 as=0 ps=0 
M5131 diff_94000_5193000# diff_94000_5193000# diff_3697000_1099000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M5132 diff_3633000_1168000# diff_3353000_2408000# diff_847000_1210000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5133 diff_3397000_928000# diff_3170000_2724000# diff_3373000_928000# GND efet w=21000 l=12000
+ ad=3.78e+08 pd=78000 as=0 ps=0 
M5134 diff_3427000_934000# diff_3422000_893000# diff_3424000_872000# GND efet w=14000 l=35000
+ ad=0 pd=0 as=4.39e+08 ps=86000 
M5135 diff_3437000_1029000# diff_3422000_893000# diff_3409000_959000# GND efet w=14500 l=83500
+ ad=0 pd=0 as=2.68e+08 ps=104000 
M5136 diff_3499000_875000# diff_3422000_893000# diff_3437000_1029000# GND efet w=14000 l=24000
+ ad=5.55e+08 pd=98000 as=0 ps=0 
M5137 diff_3557000_956000# diff_3438000_2491000# diff_3538000_920000# GND efet w=106500 l=12500
+ ad=1.075e+09 pd=232000 as=9.12e+08 ps=226000 
M5138 diff_3578000_992000# diff_3566000_784000# diff_3557000_956000# GND efet w=109500 l=11500
+ ad=1.505e+09 pd=290000 as=0 ps=0 
M5139 diff_3610000_906000# diff_3595000_2394000# diff_3578000_992000# GND efet w=122000 l=12000
+ ad=1.341e+09 pd=284000 as=0 ps=0 
M5140 diff_3632000_946000# diff_3353000_2408000# diff_3610000_906000# GND efet w=21000 l=12000
+ ad=8.34e+08 pd=158000 as=0 ps=0 
M5141 diff_3819000_1288000# diff_3801000_831000# diff_3795000_1343000# GND efet w=104000 l=12000
+ ad=1.267e+09 pd=240000 as=1.008e+09 ps=232000 
M5142 diff_3847000_1324000# diff_3829000_786000# diff_3819000_1288000# GND efet w=104000 l=12000
+ ad=1.205e+09 pd=236000 as=0 ps=0 
M5143 diff_3881000_1306000# diff_3694000_2724000# diff_3864000_1391000# GND efet w=88000 l=12000
+ ad=-1.50997e+09 pd=478000 as=8.93e+08 ps=210000 
M5144 diff_82000_3097000# diff_3901000_1417000# diff_3881000_1306000# GND efet w=207000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5145 diff_3949000_1339000# diff_3938000_1304000# diff_82000_3097000# GND efet w=65500 l=9500
+ ad=1.112e+09 pd=190000 as=0 ps=0 
M5146 diff_816000_1210000# diff_3801000_831000# diff_3697000_1099000# GND efet w=103500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M5147 diff_3847000_1127000# diff_3829000_786000# diff_816000_1210000# GND efet w=103000 l=12000
+ ad=-1.94967e+08 pd=710000 as=0 ps=0 
M5148 diff_3685000_1184000# diff_3633000_1168000# diff_82000_3097000# GND efet w=66500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5149 diff_3697000_1099000# diff_3685000_1184000# diff_82000_3097000# GND efet w=204000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5150 diff_3578000_1133000# diff_3738000_825000# diff_3697000_1099000# GND efet w=88000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5151 diff_4056000_1466000# diff_4038000_1572000# diff_82000_3097000# GND efet w=62000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5152 diff_4067000_1476000# diff_4056000_1466000# diff_82000_3097000# GND efet w=205500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5153 diff_816000_1587000# diff_4107000_2724000# diff_4067000_1476000# GND efet w=88000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5154 diff_4185000_1452000# diff_4162000_2432000# diff_4166000_1562000# GND efet w=87000 l=12000
+ ad=1.501e+09 pd=366000 as=9.23e+08 ps=208000 
M5155 diff_4305000_1753000# diff_4276000_2780000# diff_4264000_1839000# GND efet w=86000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5156 diff_4264000_1839000# diff_3320000_2526000# diff_4274000_1612000# GND efet w=45000 l=11000
+ ad=0 pd=0 as=8.31e+08 ps=168000 
M5157 diff_4225000_1648000# diff_4225000_1648000# diff_4232000_1627000# GND efet w=13000 l=38000
+ ad=0 pd=0 as=3.79e+08 ps=80000 
M5158 diff_4274000_1612000# diff_4274000_1612000# diff_4274000_1612000# GND efet w=1000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M5159 diff_4274000_1612000# diff_4274000_1612000# diff_4287000_1631000# GND efet w=15000 l=38000
+ ad=0 pd=0 as=5.97e+08 ps=104000 
M5160 diff_4286000_1500000# diff_4286000_1500000# diff_4287000_1631000# GND efet w=14000 l=23000
+ ad=1.47e+09 pd=296000 as=0 ps=0 
M5161 diff_4067000_1406000# diff_4056000_1396000# diff_82000_3097000# GND efet w=206500 l=9500
+ ad=-1.39497e+09 pd=476000 as=0 ps=0 
M5162 diff_82000_3097000# diff_4037000_1296000# diff_4057000_1357000# GND efet w=63000 l=10000
+ ad=0 pd=0 as=1.012e+09 ps=182000 
M5163 diff_4149000_1346000# diff_4107000_2724000# diff_4067000_1406000# GND efet w=88000 l=11000
+ ad=1.128e+09 pd=214000 as=0 ps=0 
M5164 diff_4204000_1414000# diff_4192000_1025000# diff_4185000_1452000# GND efet w=108500 l=12500
+ ad=-6.14967e+08 pd=548000 as=0 ps=0 
M5165 diff_4204000_1414000# diff_4192000_1025000# diff_4184000_1383000# GND efet w=107000 l=12000
+ ad=0 pd=0 as=1.598e+09 ps=366000 
M5166 diff_4267000_1500000# diff_4225000_1648000# diff_4245000_1443000# GND efet w=103000 l=11000
+ ad=8.24e+08 pd=222000 as=-9.08935e+08 ps=976000 
M5167 diff_4286000_1500000# diff_4274000_1612000# diff_4267000_1500000# GND efet w=103000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5168 diff_4306000_1553000# diff_4267000_1478000# diff_4267000_1478000# GND efet w=14000 l=40000
+ ad=1.798e+09 pd=248000 as=9.94e+08 ps=202000 
M5169 diff_4380000_2279000# diff_4347000_2438000# diff_4354000_1418000# GND efet w=101500 l=10500
+ ad=1.089e+09 pd=216000 as=7.80164e+08 ps=3.294e+06 
M5170 diff_4379000_2146000# diff_4347000_2438000# diff_4354000_1418000# GND efet w=103000 l=11000
+ ad=1.06e+09 pd=218000 as=0 ps=0 
M5171 diff_4675000_2475000# diff_4601000_2751000# diff_4642000_2735000# GND efet w=451000 l=11000
+ ad=2.02003e+09 pd=858000 as=0 ps=0 
M5172 diff_4761000_2747000# diff_4741000_2690000# diff_4704000_2610000# GND efet w=16000 l=14000
+ ad=1.02e+09 pd=168000 as=2.041e+09 ps=398000 
M5173 diff_4739000_2640000# diff_4739000_2640000# diff_4718000_2635000# GND efet w=14000 l=10000
+ ad=-1.48997e+09 pd=616000 as=1.843e+09 ps=252000 
M5174 diff_4718000_2635000# diff_4704000_2610000# diff_4704000_2610000# GND efet w=15000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M5175 diff_4704000_2610000# diff_4688000_2591000# diff_4675000_2475000# GND efet w=68500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5176 diff_4777000_2518000# diff_4761000_2747000# diff_4739000_2640000# GND efet w=163500 l=10500
+ ad=6.61033e+08 pd=444000 as=0 ps=0 
M5177 diff_4837000_2673000# diff_4825000_2753000# diff_4804000_2758000# GND efet w=17000 l=13000
+ ad=1.08e+09 pd=176000 as=1.78e+09 ps=384000 
M5178 diff_4838000_2617000# diff_4838000_2617000# diff_4819000_2721000# GND efet w=14000 l=10000
+ ad=-1.59097e+09 pd=578000 as=2.002e+09 ps=322000 
M5179 diff_4905000_2664000# diff_4905000_2664000# diff_4896000_2688000# GND efet w=14000 l=10000
+ ad=-1.16397e+09 pd=646000 as=6.98e+08 ps=142000 
M5180 diff_4905000_2664000# diff_4882000_2652000# diff_4888000_2467000# GND efet w=169500 l=10500
+ ad=0 pd=0 as=-9.19967e+08 ps=402000 
M5181 diff_4819000_2721000# diff_4804000_2758000# diff_4804000_2758000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M5182 diff_4804000_2758000# diff_4784000_2782000# diff_4777000_2518000# GND efet w=78000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5183 diff_4434000_2245000# diff_4373000_832000# diff_4410000_2197000# GND efet w=22000 l=12000
+ ad=9.57e+08 pd=168000 as=1.054e+09 ps=184000 
M5184 diff_4460000_2077000# diff_4416000_951000# diff_4434000_2245000# GND efet w=22000 l=12000
+ ad=2.089e+09 pd=418000 as=0 ps=0 
M5185 diff_4481000_2228000# diff_4478000_2251000# diff_4478000_2251000# GND efet w=15000 l=105000
+ ad=4.02e+08 pd=82000 as=7.23e+08 ps=154000 
M5186 diff_4531000_2370000# diff_4517000_2326000# diff_4517000_2326000# GND efet w=14000 l=21000
+ ad=4.38e+08 pd=86000 as=1.859e+09 ps=338000 
M5187 diff_4517000_2326000# diff_4532000_2229000# diff_4519000_2127000# GND efet w=51000 l=10000
+ ad=0 pd=0 as=-1.47997e+09 ps=472000 
M5188 diff_4588000_2371000# diff_4574000_2327000# diff_4574000_2327000# GND efet w=14000 l=23000
+ ad=1.168e+09 pd=152000 as=1.672e+09 ps=304000 
M5189 diff_4588000_2371000# diff_4607000_2223000# diff_4607000_2223000# GND efet w=15000 l=22000
+ ad=0 pd=0 as=1.903e+09 ps=406000 
M5190 diff_4574000_2327000# diff_4497000_2491000# diff_4563000_2272000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=3.74e+08 ps=78000 
M5191 diff_4888000_2467000# diff_4837000_2673000# diff_4838000_2617000# GND efet w=162000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5192 diff_4996000_2788000# diff_4944000_2493000# diff_4944000_2493000# GND efet w=14000 l=23000
+ ad=5.29e+08 pd=94000 as=5.93033e+08 ps=732000 
M5193 diff_5171000_2829000# diff_71000_4514000# diff_4974000_2909000# GND efet w=15000 l=13000
+ ad=2.087e+09 pd=442000 as=9.28e+08 ps=214000 
M5194 diff_4761000_3820000# diff_71000_4514000# diff_4931000_2481000# GND efet w=17000 l=13000
+ ad=0 pd=0 as=1.189e+09 ps=166000 
M5195 diff_5013000_2754000# diff_4991000_2691000# diff_4958000_2607000# GND efet w=16000 l=13000
+ ad=1.098e+09 pd=178000 as=1.563e+09 ps=340000 
M5196 diff_4842000_3066000# diff_5085000_2690000# diff_5113000_2489000# GND efet w=22000 l=14000
+ ad=0 pd=0 as=5.5e+08 ps=126000 
M5197 diff_5203000_3036000# diff_5203000_3036000# diff_94000_5193000# GND efet w=23000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5198 diff_4494000_3313000# diff_5257000_2805000# diff_5264000_2777000# GND efet w=22000 l=14000
+ ad=0 pd=0 as=9.52e+08 ps=160000 
M5199 diff_4655000_3019000# diff_5257000_2805000# diff_5317000_2777000# GND efet w=22000 l=14000
+ ad=0 pd=0 as=9.64e+08 ps=140000 
M5200 diff_5052000_2756000# diff_4931000_826000# diff_4931000_826000# GND efet w=19000 l=11000
+ ad=3.04e+08 pd=70000 as=4.51033e+08 ps=932000 
M5201 diff_4993000_2633000# diff_4993000_2633000# diff_4971000_2631000# GND efet w=15000 l=10000
+ ad=2.084e+09 pd=492000 as=1.615e+09 ps=274000 
M5202 diff_5028000_2635000# diff_5013000_2754000# diff_4993000_2633000# GND efet w=178500 l=10500
+ ad=-1.10497e+09 pd=474000 as=0 ps=0 
M5203 diff_4931000_826000# diff_5034000_2443000# diff_5028000_2635000# GND efet w=235000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5204 diff_5074000_2676000# diff_5064000_2665000# diff_4931000_826000# GND efet w=214500 l=10500
+ ad=-7.58967e+08 pd=506000 as=0 ps=0 
M5205 diff_5186000_2411000# diff_5186000_2411000# diff_5190000_2733000# GND efet w=13000 l=17000
+ ad=-6.90967e+08 pd=662000 as=3.73e+08 ps=78000 
M5206 diff_4971000_2631000# diff_4958000_2607000# diff_4958000_2607000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M5207 diff_4958000_2607000# diff_4944000_2493000# diff_4968000_2493000# GND efet w=76000 l=10000
+ ad=0 pd=0 as=1.969e+09 ps=218000 
M5208 diff_4968000_2493000# diff_4931000_2481000# diff_4944000_2493000# GND efet w=65000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5209 diff_4701000_2373000# diff_4693000_2316000# diff_4693000_2316000# GND efet w=15000 l=27000
+ ad=1.446e+09 pd=178000 as=8.33e+08 ps=156000 
M5210 diff_4701000_2373000# diff_4726000_2237000# diff_4726000_2237000# GND efet w=15000 l=27000
+ ad=0 pd=0 as=1.638e+09 ps=296000 
M5211 diff_4481000_2154000# diff_4477000_1873000# diff_4477000_1873000# GND efet w=14000 l=105000
+ ad=3.34e+08 pd=74000 as=1.174e+09 ps=200000 
M5212 diff_4517000_2031000# diff_4532000_2086000# diff_4519000_2127000# GND efet w=51000 l=10000
+ ad=1.787e+09 pd=336000 as=0 ps=0 
M5213 diff_4617000_2117000# diff_4607000_2223000# diff_4574000_2327000# GND efet w=50000 l=10000
+ ad=-1.42397e+09 pd=390000 as=0 ps=0 
M5214 diff_4607000_2223000# diff_4624000_2286000# diff_4617000_2117000# GND efet w=69000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5215 diff_4672000_2273000# diff_4547000_2724000# diff_4607000_2223000# GND efet w=23000 l=12000
+ ad=4.6e+08 pd=86000 as=0 ps=0 
M5216 diff_4706000_2273000# diff_4601000_2751000# diff_4672000_2273000# GND efet w=23000 l=14000
+ ad=4.37e+08 pd=84000 as=0 ps=0 
M5217 diff_4574000_2030000# diff_4497000_2491000# diff_4563000_2106000# GND efet w=23000 l=12000
+ ad=1.684e+09 pd=304000 as=3.91e+08 ps=80000 
M5218 diff_4617000_2117000# diff_4607000_2076000# diff_4574000_2030000# GND efet w=52000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5219 diff_4607000_2076000# diff_4624000_2092000# diff_4617000_2117000# GND efet w=69000 l=10000
+ ad=1.892e+09 pd=404000 as=0 ps=0 
M5220 diff_4706000_2228000# diff_4601000_2751000# diff_4675000_2228000# GND efet w=22000 l=14000
+ ad=4.78e+08 pd=144000 as=3.74e+08 ps=78000 
M5221 diff_4753000_2186000# diff_4706000_2228000# diff_4726000_2237000# GND efet w=51000 l=10000
+ ad=1.61503e+09 pd=782000 as=0 ps=0 
M5222 diff_4787000_2229000# diff_4739000_2640000# diff_4753000_2186000# GND efet w=150500 l=10500
+ ad=1.658e+09 pd=366000 as=0 ps=0 
M5223 diff_4809000_2270000# diff_4798000_2261000# diff_4787000_2229000# GND efet w=128000 l=11000
+ ad=2.114e+09 pd=412000 as=0 ps=0 
M5224 diff_4831000_2306000# diff_4820000_2281000# diff_4809000_2270000# GND efet w=71000 l=11000
+ ad=-1.94497e+09 pd=394000 as=0 ps=0 
M5225 diff_4881000_2375000# diff_4870000_2312000# diff_4870000_2312000# GND efet w=14000 l=24000
+ ad=4.82e+08 pd=90000 as=-1.40597e+09 ps=460000 
M5226 diff_5200000_2422000# diff_3407000_4287000# diff_5186000_2411000# GND efet w=105000 l=11000
+ ad=-1.03193e+09 pd=918000 as=0 ps=0 
M5227 diff_5163000_2687000# diff_5123000_2494000# diff_5123000_2494000# GND efet w=15000 l=23000
+ ad=5.46e+08 pd=98000 as=-1.04897e+09 ps=570000 
M5228 diff_5163000_2687000# diff_4931000_826000# diff_5141000_2399000# GND efet w=15000 l=10000
+ ad=0 pd=0 as=1.43003e+09 ps=1.022e+06 
M5229 diff_5186000_2543000# diff_5174000_2532000# diff_5141000_2399000# GND efet w=165500 l=11500
+ ad=1.866e+09 pd=332000 as=0 ps=0 
M5230 diff_5123000_2494000# diff_5113000_2489000# diff_5074000_2676000# GND efet w=67000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5231 diff_5141000_2519000# diff_4931000_826000# diff_5123000_2494000# GND efet w=93500 l=9500
+ ad=1.02e+09 pd=190000 as=0 ps=0 
M5232 diff_4899000_2195000# diff_4904000_2299000# diff_4870000_2312000# GND efet w=53000 l=10000
+ ad=6.15033e+08 pd=810000 as=0 ps=0 
M5233 diff_4870000_2312000# diff_4838000_2617000# diff_4866000_2115000# GND efet w=63000 l=10000
+ ad=0 pd=0 as=-1.17297e+09 ps=460000 
M5234 diff_4831000_2306000# diff_4820000_2281000# diff_4809000_2270000# GND efet w=70500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5235 diff_4706000_2150000# diff_4601000_2751000# diff_4675000_2150000# GND efet w=22000 l=14000
+ ad=5.03e+08 pd=144000 as=3.74e+08 ps=78000 
M5236 diff_4809000_2270000# diff_4798000_2261000# diff_4787000_2229000# GND efet w=14000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5237 diff_4866000_2115000# diff_4838000_2617000# diff_4831000_2306000# GND efet w=53000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5238 diff_4809000_2023000# diff_4799000_2016000# diff_4787000_2161000# GND efet w=12000 l=10000
+ ad=2.098e+09 pd=412000 as=1.741e+09 ps=366000 
M5239 diff_4379000_1851000# diff_4347000_2438000# diff_4354000_1418000# GND efet w=104000 l=9000
+ ad=1.126e+09 pd=220000 as=0 ps=0 
M5240 diff_4459000_1939000# diff_4416000_951000# diff_4432000_2036000# GND efet w=21000 l=12000
+ ad=1.278e+09 pd=254000 as=1.937e+09 ps=364000 
M5241 diff_4432000_2036000# diff_4373000_832000# diff_4409000_1887000# GND efet w=21000 l=12000
+ ad=0 pd=0 as=-1.22097e+09 ps=540000 
M5242 diff_4517000_2031000# diff_4517000_2031000# diff_4531000_1993000# GND efet w=14000 l=21000
+ ad=0 pd=0 as=7.8e+08 ps=120000 
M5243 diff_4435000_1905000# diff_4373000_832000# diff_4409000_1887000# GND efet w=21000 l=12000
+ ad=8.28e+08 pd=172000 as=0 ps=0 
M5244 diff_4379000_1770000# diff_4347000_2438000# diff_4354000_1418000# GND efet w=102000 l=10000
+ ad=1.137e+09 pd=218000 as=0 ps=0 
M5245 diff_4460000_1689000# diff_4416000_951000# diff_4435000_1905000# GND efet w=23000 l=11000
+ ad=-1.97797e+09 pd=428000 as=0 ps=0 
M5246 diff_4477000_1873000# diff_4477000_1873000# diff_4480000_1851000# GND efet w=14000 l=106000
+ ad=0 pd=0 as=3.86e+08 ps=80000 
M5247 diff_4531000_1993000# diff_4517000_1949000# diff_4517000_1949000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=1.863e+09 ps=336000 
M5248 diff_4517000_1949000# diff_4532000_1851000# diff_4519000_1750000# GND efet w=51000 l=10000
+ ad=0 pd=0 as=-1.48797e+09 ps=470000 
M5249 diff_4672000_2104000# diff_4547000_2724000# diff_4607000_2076000# GND efet w=22000 l=12000
+ ad=4.4e+08 pd=84000 as=0 ps=0 
M5250 diff_4706000_2104000# diff_4601000_2751000# diff_4672000_2104000# GND efet w=22000 l=14000
+ ad=4.39e+08 pd=84000 as=0 ps=0 
M5251 diff_4753000_2186000# diff_4706000_2150000# diff_4726000_2137000# GND efet w=52000 l=10000
+ ad=0 pd=0 as=1.625e+09 ps=300000 
M5252 diff_4787000_2161000# diff_4739000_2640000# diff_4753000_2186000# GND efet w=149500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5253 diff_4574000_2030000# diff_4574000_2030000# diff_4588000_1994000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=1.566e+09 ps=180000 
M5254 diff_4607000_2076000# diff_4607000_2076000# diff_4588000_1994000# GND efet w=15000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5255 diff_4588000_1994000# diff_4574000_1950000# diff_4574000_1950000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=1.682e+09 ps=306000 
M5256 diff_4588000_1994000# diff_4607000_1846000# diff_4607000_1846000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=1.878e+09 ps=402000 
M5257 diff_4574000_1950000# diff_4497000_2491000# diff_4563000_1895000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=3.73e+08 ps=78000 
M5258 diff_4692000_2057000# diff_4692000_2057000# diff_4701000_1996000# GND efet w=15000 l=27000
+ ad=8.16e+08 pd=156000 as=1.917e+09 ps=202000 
M5259 diff_4726000_2137000# diff_4726000_2137000# diff_4701000_1996000# GND efet w=16000 l=26000
+ ad=0 pd=0 as=0 ps=0 
M5260 diff_4809000_2023000# diff_4799000_2016000# diff_4787000_2161000# GND efet w=127000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5261 diff_4831000_2023000# diff_4821000_2015000# diff_4809000_2023000# GND efet w=68500 l=10500
+ ad=-2.01397e+09 pd=388000 as=0 ps=0 
M5262 diff_4899000_2195000# diff_4893000_2206000# diff_4870000_2312000# GND efet w=60000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5263 diff_4951000_2235000# diff_4904000_2299000# diff_4899000_2195000# GND efet w=136000 l=10000
+ ad=1.224e+09 pd=290000 as=0 ps=0 
M5264 diff_4971000_2235000# diff_4905000_2664000# diff_4951000_2235000# GND efet w=136000 l=11000
+ ad=1.638e+09 pd=348000 as=0 ps=0 
M5265 diff_4991000_2210000# diff_4982000_2204000# diff_4971000_2235000# GND efet w=97000 l=9000
+ ad=-2.03097e+09 pd=394000 as=0 ps=0 
M5266 diff_5270000_2492000# diff_5264000_2777000# diff_5200000_2422000# GND efet w=247500 l=10500
+ ad=-1.06297e+09 pd=678000 as=0 ps=0 
M5267 diff_5299000_2749000# diff_5270000_2492000# diff_5270000_2492000# GND efet w=19000 l=10000
+ ad=4.97e+08 pd=94000 as=0 ps=0 
M5268 diff_5320000_2718000# diff_5320000_2718000# diff_5299000_2749000# GND efet w=24000 l=9000
+ ad=-4.06967e+08 pd=568000 as=0 ps=0 
M5269 diff_5300000_2536000# diff_5289000_2527000# diff_5270000_2492000# GND efet w=204500 l=10500
+ ad=1.52065e+08 pd=1.026e+06 as=0 ps=0 
M5270 diff_5200000_2422000# diff_5235000_2513000# diff_5186000_2411000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5271 diff_5320000_2718000# diff_5314000_2695000# diff_5300000_2536000# GND efet w=258000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5272 diff_5300000_2536000# diff_5317000_2777000# diff_5320000_2718000# GND efet w=127000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5273 diff_5387000_2603000# diff_5317000_2777000# diff_5300000_2536000# GND efet w=155000 l=9000
+ ad=2.13e+09 pd=360000 as=0 ps=0 
M5274 diff_5200000_2422000# diff_5186000_2411000# diff_5200000_2399000# GND efet w=91500 l=11500
+ ad=0 pd=0 as=1.82e+09 ps=294000 
M5275 diff_6212000_3182000# diff_3568000_3529000# diff_82000_3097000# GND efet w=94500 l=10500
+ ad=-1.68097e+09 pd=494000 as=0 ps=0 
M5276 diff_82000_3097000# diff_4240000_2639000# diff_6212000_3182000# GND efet w=94000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5277 diff_6251000_3156000# diff_5097000_4893000# diff_6212000_3182000# GND efet w=93500 l=10500
+ ad=-8.97967e+08 pd=604000 as=0 ps=0 
M5278 diff_82000_3097000# diff_5008000_4961000# diff_5987000_3968000# GND efet w=43000 l=11000
+ ad=0 pd=0 as=-2.02497e+09 ps=436000 
M5279 diff_6212000_3182000# diff_3407000_4287000# diff_6251000_3156000# GND efet w=88000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5280 diff_5987000_3968000# diff_5067000_4961000# diff_82000_3097000# GND efet w=43000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5281 diff_82000_3097000# diff_5038000_4961000# diff_5987000_3968000# GND efet w=43000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5282 diff_94000_5193000# diff_6251000_3156000# diff_6251000_3156000# GND efet w=15000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M5283 diff_5987000_3968000# diff_5987000_3968000# diff_94000_5193000# GND efet w=15000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M5284 diff_5625000_2883000# diff_5618000_2892000# diff_82000_3097000# GND efet w=158000 l=12000
+ ad=-2.08197e+09 pd=400000 as=0 ps=0 
M5285 diff_5625000_2883000# diff_71000_4514000# diff_5617000_2717000# GND efet w=21000 l=13000
+ ad=0 pd=0 as=1.155e+09 ps=238000 
M5286 diff_5768000_2822000# diff_5256000_3172000# diff_82000_3097000# GND efet w=486000 l=11000
+ ad=6.19065e+08 pd=1.632e+06 as=0 ps=0 
M5287 diff_94000_5193000# diff_5625000_2883000# diff_5625000_2883000# GND efet w=14000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M5288 diff_94000_5193000# diff_5768000_2822000# diff_5618000_2892000# GND efet w=733000 l=10000
+ ad=0 pd=0 as=4.53597e+07 ps=6.924e+06 
M5289 diff_94000_5193000# diff_5652000_2806000# diff_5617000_2717000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M5290 diff_5652000_2806000# diff_5631000_2728000# diff_82000_3097000# GND efet w=48500 l=9500
+ ad=1.126e+09 pd=208000 as=0 ps=0 
M5291 diff_94000_5193000# diff_5768000_2822000# diff_5618000_2892000# GND efet w=289000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5292 diff_82000_3097000# diff_82000_3097000# diff_5618000_2892000# GND efet w=82000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M5293 diff_5618000_2171000# diff_82000_3097000# diff_82000_3097000# GND efet w=82000 l=14000
+ ad=-6.69608e+08 pd=7.514e+06 as=0 ps=0 
M5294 diff_5768000_2822000# diff_5696000_2541000# diff_82000_3097000# GND efet w=480000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5295 diff_94000_5193000# diff_5768000_2822000# diff_5618000_2892000# GND efet w=287500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5296 diff_94000_5193000# diff_5652000_2806000# diff_5652000_2806000# GND efet w=13000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M5297 diff_5652000_2806000# diff_71000_4514000# diff_82000_3097000# GND efet w=29000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5298 diff_5631000_2728000# diff_5617000_2717000# diff_82000_3097000# GND efet w=224500 l=10500
+ ad=-5.83967e+08 pd=730000 as=0 ps=0 
M5299 diff_94000_5193000# diff_5631000_2728000# diff_5631000_2728000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M5300 diff_5618000_2892000# diff_5768000_2822000# diff_94000_5193000# GND efet w=289500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5301 diff_5768000_2822000# diff_5768000_2822000# diff_94000_5193000# GND efet w=46000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5302 diff_94000_5193000# diff_5696000_2541000# diff_5696000_2541000# GND efet w=35000 l=10000
+ ad=0 pd=0 as=1.47707e+09 ps=1.8e+06 
M5303 diff_82000_3097000# diff_5696000_2541000# diff_5618000_2892000# GND efet w=240500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M5304 diff_5696000_2541000# diff_5256000_3172000# diff_82000_3097000# GND efet w=478500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5305 diff_5631000_2728000# diff_5555000_2636000# diff_5537000_2618000# GND efet w=89000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M5306 diff_82000_3097000# diff_5650000_2540000# diff_5696000_2541000# GND efet w=515500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5307 diff_5028000_2372000# diff_5021000_2345000# diff_5021000_2345000# GND efet w=15000 l=27000
+ ad=5.07e+08 pd=92000 as=1.894e+09 ps=298000 
M5308 diff_5074000_2370000# diff_5068000_2348000# diff_5068000_2348000# GND efet w=15000 l=22000
+ ad=8.31e+08 pd=132000 as=1.693e+09 ps=364000 
M5309 diff_5124000_2368000# diff_4931000_826000# diff_5074000_2370000# GND efet w=14000 l=10000
+ ad=2.20327e+07 pd=874000 as=0 ps=0 
M5310 diff_5141000_2399000# diff_5151000_2372000# diff_5124000_2368000# GND efet w=131000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5311 diff_4899000_2195000# diff_4893000_2186000# diff_4869000_2081000# GND efet w=61000 l=10000
+ ad=0 pd=0 as=-1.29397e+09 ps=472000 
M5312 diff_4866000_2115000# diff_4838000_2617000# diff_4831000_2023000# GND efet w=51000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5313 diff_4991000_2210000# diff_4982000_2204000# diff_4971000_2235000# GND efet w=35000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5314 diff_5024000_2111000# diff_4993000_2633000# diff_4991000_2210000# GND efet w=57000 l=11000
+ ad=-1.59697e+09 pd=418000 as=0 ps=0 
M5315 diff_5021000_2345000# diff_5037000_2263000# diff_5024000_2111000# GND efet w=46000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5316 diff_5124000_2368000# diff_5132000_2347000# diff_5111000_2140000# GND efet w=92000 l=13000
+ ad=0 pd=0 as=-1.68193e+09 ps=808000 
M5317 diff_5068000_2348000# diff_5068000_2286000# diff_5070000_2118000# GND efet w=67500 l=10500
+ ad=0 pd=0 as=1.875e+09 ps=374000 
M5318 diff_5111000_2140000# diff_4931000_826000# diff_5068000_2348000# GND efet w=67000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5319 diff_5208000_2365000# diff_5201000_2341000# diff_5201000_2341000# GND efet w=15000 l=24000
+ ad=8.63e+08 pd=128000 as=1.628e+09 ps=348000 
M5320 diff_5242000_2359000# diff_5242000_2359000# diff_5208000_2365000# GND efet w=14000 l=23000
+ ad=-2.13697e+09 pd=494000 as=0 ps=0 
M5321 diff_5289000_2222000# diff_5278000_2280000# diff_5242000_2359000# GND efet w=79500 l=10500
+ ad=1.289e+09 pd=324000 as=0 ps=0 
M5322 diff_4831000_2023000# diff_4821000_2015000# diff_4809000_2023000# GND efet w=70000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5323 diff_4869000_2081000# diff_4838000_2617000# diff_4866000_2115000# GND efet w=59500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5324 diff_4701000_1996000# diff_4693000_1939000# diff_4693000_1939000# GND efet w=15000 l=27000
+ ad=0 pd=0 as=8.33e+08 ps=156000 
M5325 diff_4701000_1996000# diff_4726000_1860000# diff_4726000_1860000# GND efet w=15000 l=26000
+ ad=0 pd=0 as=1.627e+09 ps=296000 
M5326 diff_4267000_1478000# diff_4225000_1648000# diff_4245000_1443000# GND efet w=53500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5327 diff_3881000_1306000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M5328 diff_3938000_1304000# diff_94000_5193000# diff_3881000_1306000# GND efet w=14500 l=80500
+ ad=8.88e+08 pd=254000 as=0 ps=0 
M5329 diff_3949000_1339000# diff_94000_5193000# diff_94000_5193000# GND efet w=15000 l=33000
+ ad=0 pd=0 as=0 ps=0 
M5330 diff_4005000_1296000# diff_3921000_785000# diff_3938000_1304000# GND efet w=22000 l=12000
+ ad=4.4e+08 pd=84000 as=0 ps=0 
M5331 diff_4037000_1296000# diff_4003000_2724000# diff_4005000_1296000# GND efet w=22000 l=12000
+ ad=9.29e+08 pd=238000 as=0 ps=0 
M5332 diff_94000_5193000# diff_94000_5193000# diff_3847000_1127000# GND efet w=13000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M5333 diff_3937000_1185000# diff_94000_5193000# diff_3847000_1127000# GND efet w=14000 l=76000
+ ad=8.69e+08 pd=268000 as=0 ps=0 
M5334 diff_94000_5193000# diff_94000_5193000# diff_3901000_1073000# GND efet w=15000 l=35000
+ ad=0 pd=0 as=1.079e+09 ps=188000 
M5335 diff_4057000_1357000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=33000
+ ad=0 pd=0 as=0 ps=0 
M5336 diff_4067000_1406000# diff_94000_5193000# diff_4037000_1296000# GND efet w=14000 l=81000
+ ad=0 pd=0 as=0 ps=0 
M5337 diff_4067000_1406000# diff_94000_5193000# diff_94000_5193000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M5338 diff_3697000_1029000# diff_3687000_1019000# diff_82000_3097000# GND efet w=206000 l=10000
+ ad=-1.48897e+09 pd=470000 as=0 ps=0 
M5339 diff_3686000_934000# diff_3670000_960000# diff_82000_3097000# GND efet w=72500 l=10500
+ ad=1.042e+09 pd=192000 as=0 ps=0 
M5340 diff_3780000_968000# diff_3738000_825000# diff_3697000_1029000# GND efet w=89000 l=12000
+ ad=9.87e+08 pd=214000 as=0 ps=0 
M5341 diff_3847000_1127000# diff_3694000_2724000# diff_3578000_1133000# GND efet w=88000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5342 diff_816000_1210000# diff_3921000_785000# diff_3937000_1185000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5343 diff_4037000_1195000# diff_4003000_2724000# diff_816000_1210000# GND efet w=22000 l=12000
+ ad=9.17e+08 pd=246000 as=0 ps=0 
M5344 diff_94000_5193000# diff_94000_5193000# diff_4056000_1090000# GND efet w=15000 l=35000
+ ad=0 pd=0 as=1.022e+09 ps=184000 
M5345 diff_4067000_1099000# diff_94000_5193000# diff_4037000_1195000# GND efet w=14000 l=76000
+ ad=-1.29397e+09 pd=480000 as=0 ps=0 
M5346 diff_4184000_1383000# diff_4162000_2432000# diff_4165000_1308000# GND efet w=89000 l=12000
+ ad=0 pd=0 as=9.05e+08 ps=214000 
M5347 diff_94000_5193000# diff_94000_5193000# diff_4067000_1099000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M5348 diff_82000_3097000# diff_3901000_1073000# diff_3847000_1127000# GND efet w=205000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5349 diff_3901000_1073000# diff_3937000_1185000# diff_82000_3097000# GND efet w=64000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5350 diff_3353000_2408000# diff_3334000_772000# diff_3361000_767000# GND efet w=83000 l=12000
+ ad=0 pd=0 as=-1.79797e+09 ps=326000 
M5351 diff_3170000_2724000# diff_3411000_824000# diff_3361000_767000# GND efet w=86000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5352 diff_3659000_908000# diff_3488000_2724000# diff_3632000_946000# GND efet w=23000 l=12000
+ ad=4.28e+08 pd=88000 as=0 ps=0 
M5353 diff_3686000_934000# diff_3683000_893000# diff_3684000_872000# GND efet w=14000 l=35000
+ ad=0 pd=0 as=4.02e+08 ps=82000 
M5354 diff_3697000_1029000# diff_3683000_893000# diff_3670000_960000# GND efet w=14500 l=82500
+ ad=0 pd=0 as=2.81e+08 ps=104000 
M5355 diff_3473000_793000# diff_3411000_824000# diff_3473000_771000# GND efet w=80000 l=11000
+ ad=0 pd=0 as=1.81e+09 ps=258000 
M5356 diff_3438000_2491000# diff_3526000_822000# diff_3473000_771000# GND efet w=76000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5357 diff_3697000_1029000# diff_3683000_893000# diff_3758000_876000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=5.39e+08 ps=96000 
M5358 diff_3819000_912000# diff_3801000_831000# diff_3795000_966000# GND efet w=103500 l=11500
+ ad=1.246e+09 pd=238000 as=1.075e+09 ps=232000 
M5359 diff_3847000_947000# diff_3829000_786000# diff_3819000_912000# GND efet w=103000 l=12000
+ ad=1.206e+09 pd=234000 as=0 ps=0 
M5360 diff_3881000_929000# diff_3694000_2724000# diff_3864000_1014000# GND efet w=89000 l=12000
+ ad=-1.54897e+09 pd=472000 as=9.01e+08 ps=212000 
M5361 diff_82000_3097000# diff_3901000_1040000# diff_3881000_929000# GND efet w=207000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5362 diff_3949000_962000# diff_3938000_928000# diff_82000_3097000# GND efet w=65500 l=9500
+ ad=1.067e+09 pd=188000 as=0 ps=0 
M5363 diff_4056000_1090000# diff_4037000_1195000# diff_82000_3097000# GND efet w=62000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5364 diff_4067000_1099000# diff_4056000_1090000# diff_82000_3097000# GND efet w=204500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5365 diff_816000_1210000# diff_4107000_2724000# diff_4067000_1099000# GND efet w=88000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5366 diff_4185000_1075000# diff_4162000_2432000# diff_4166000_1185000# GND efet w=87000 l=12000
+ ad=1.513e+09 pd=366000 as=9.16e+08 ps=208000 
M5367 diff_4242000_1303000# diff_4226000_1550000# diff_4204000_1414000# GND efet w=110000 l=11000
+ ad=1.274e+09 pd=300000 as=0 ps=0 
M5368 diff_4262000_1287000# diff_4252000_1283000# diff_4242000_1303000# GND efet w=30000 l=11000
+ ad=1.62003e+09 pd=860000 as=0 ps=0 
M5369 diff_4262000_1287000# diff_4252000_1283000# diff_4242000_1303000# GND efet w=80000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5370 diff_4245000_1443000# diff_4275000_1328000# diff_4262000_1287000# GND efet w=74000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5371 diff_4373000_1474000# diff_4347000_2438000# diff_4354000_1418000# GND efet w=101000 l=10000
+ ad=1.089e+09 pd=200000 as=0 ps=0 
M5372 diff_4481000_1777000# diff_4477000_1497000# diff_4477000_1497000# GND efet w=14000 l=105000
+ ad=3.34e+08 pd=74000 as=1.164e+09 ps=200000 
M5373 diff_4517000_1654000# diff_4532000_1709000# diff_4519000_1750000# GND efet w=51000 l=10000
+ ad=1.797e+09 pd=336000 as=0 ps=0 
M5374 diff_4617000_1740000# diff_4607000_1846000# diff_4574000_1950000# GND efet w=50000 l=10000
+ ad=-1.44397e+09 pd=388000 as=0 ps=0 
M5375 diff_4607000_1846000# diff_4624000_1908000# diff_4617000_1740000# GND efet w=68000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5376 diff_4672000_1895000# diff_4547000_2724000# diff_4607000_1846000# GND efet w=23000 l=12000
+ ad=4.6e+08 pd=86000 as=0 ps=0 
M5377 diff_4706000_1895000# diff_4601000_2751000# diff_4672000_1895000# GND efet w=23000 l=14000
+ ad=4.37e+08 pd=84000 as=0 ps=0 
M5378 diff_4574000_1652000# diff_4497000_2491000# diff_4563000_1729000# GND efet w=23000 l=12000
+ ad=1.668e+09 pd=302000 as=3.91e+08 ps=80000 
M5379 diff_4617000_1740000# diff_4607000_1699000# diff_4574000_1652000# GND efet w=51000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5380 diff_4607000_1699000# diff_4624000_1715000# diff_4617000_1740000# GND efet w=69000 l=10000
+ ad=1.859e+09 pd=404000 as=0 ps=0 
M5381 diff_4706000_1850000# diff_4601000_2751000# diff_4675000_1850000# GND efet w=23000 l=14000
+ ad=5.03e+08 pd=146000 as=3.91e+08 ps=80000 
M5382 diff_4753000_1809000# diff_4706000_1850000# diff_4726000_1860000# GND efet w=51000 l=10000
+ ad=1.61903e+09 pd=782000 as=0 ps=0 
M5383 diff_4787000_1852000# diff_4739000_2640000# diff_4753000_1809000# GND efet w=150500 l=10500
+ ad=1.66e+09 pd=366000 as=0 ps=0 
M5384 diff_4809000_1892000# diff_4798000_1884000# diff_4787000_1852000# GND efet w=128000 l=11000
+ ad=2.115e+09 pd=412000 as=0 ps=0 
M5385 diff_4831000_1929000# diff_4820000_1904000# diff_4809000_1892000# GND efet w=71000 l=11000
+ ad=-1.94297e+09 pd=394000 as=0 ps=0 
M5386 diff_4899000_2195000# diff_4904000_2082000# diff_4869000_2081000# GND efet w=55000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5387 diff_4869000_2081000# diff_4869000_2081000# diff_4881000_1998000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=6.58e+08 ps=110000 
M5388 diff_4952000_2027000# diff_4904000_2082000# diff_4899000_2195000# GND efet w=137000 l=11000
+ ad=1.096e+09 pd=290000 as=0 ps=0 
M5389 diff_4971000_2027000# diff_4905000_2664000# diff_4952000_2027000# GND efet w=137000 l=11000
+ ad=1.649e+09 pd=350000 as=0 ps=0 
M5390 diff_4991000_2027000# diff_4982000_2020000# diff_4971000_2027000# GND efet w=34000 l=9000
+ ad=-2.09597e+09 pd=396000 as=0 ps=0 
M5391 diff_5334000_2356000# diff_5224000_815000# diff_5242000_2359000# GND efet w=22500 l=13500
+ ad=1.75e+08 pd=60000 as=0 ps=0 
M5392 diff_5355000_2355000# diff_5270000_856000# diff_5334000_2356000# GND efet w=22000 l=13000
+ ad=3.36e+08 pd=108000 as=0 ps=0 
M5393 diff_5124000_2368000# diff_5132000_2347000# diff_5111000_2140000# GND efet w=50000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5394 diff_5201000_2341000# diff_5141000_2399000# diff_5202000_2119000# GND efet w=79000 l=10000
+ ad=0 pd=0 as=1.915e+09 ps=362000 
M5395 diff_5124000_2017000# diff_5136000_2101000# diff_5111000_2140000# GND efet w=124000 l=11000
+ ad=8.60327e+07 pd=844000 as=0 ps=0 
M5396 diff_4991000_2027000# diff_4982000_2020000# diff_4971000_2027000# GND efet w=99000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5397 diff_5024000_2111000# diff_4993000_2633000# diff_4991000_2027000# GND efet w=55000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5398 diff_5021000_2029000# diff_5037000_2104000# diff_5024000_2111000# GND efet w=46000 l=8000
+ ad=1.819e+09 pd=296000 as=0 ps=0 
M5399 diff_5068000_2031000# diff_5068000_2093000# diff_5070000_2118000# GND efet w=66500 l=10500
+ ad=1.793e+09 pd=360000 as=0 ps=0 
M5400 diff_5111000_2140000# diff_4931000_826000# diff_5068000_2031000# GND efet w=67000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5401 diff_4881000_1998000# diff_4870000_1933000# diff_4870000_1933000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=-1.36897e+09 ps=464000 
M5402 diff_4899000_1818000# diff_4904000_1921000# diff_4870000_1933000# GND efet w=54000 l=10000
+ ad=6.30033e+08 pd=812000 as=0 ps=0 
M5403 diff_4870000_1933000# diff_4838000_2617000# diff_4866000_1738000# GND efet w=62000 l=9000
+ ad=0 pd=0 as=-1.15897e+09 ps=462000 
M5404 diff_4831000_1929000# diff_4820000_1904000# diff_4809000_1892000# GND efet w=70500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5405 diff_4706000_1772000# diff_4601000_2751000# diff_4675000_1772000# GND efet w=22000 l=14000
+ ad=5.01e+08 pd=146000 as=3.74e+08 ps=78000 
M5406 diff_4809000_1892000# diff_4798000_1884000# diff_4787000_1852000# GND efet w=14000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5407 diff_4866000_1738000# diff_4838000_2617000# diff_4831000_1929000# GND efet w=53000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5408 diff_4809000_1646000# diff_4799000_1639000# diff_4787000_1783000# GND efet w=12000 l=10000
+ ad=2.113e+09 pd=412000 as=1.748e+09 ps=366000 
M5409 diff_4460000_1561000# diff_4416000_951000# diff_4429000_1713000# GND efet w=22000 l=12000
+ ad=1.177e+09 pd=236000 as=1.46e+09 ps=280000 
M5410 diff_4429000_1713000# diff_4373000_832000# diff_4412000_1466000# GND efet w=21000 l=12000
+ ad=0 pd=0 as=-2.06297e+09 ps=456000 
M5411 diff_4517000_1654000# diff_4517000_1654000# diff_4531000_1616000# GND efet w=14000 l=21000
+ ad=0 pd=0 as=7.88e+08 ps=120000 
M5412 diff_4435000_1490000# diff_4373000_832000# diff_4412000_1466000# GND efet w=21000 l=12000
+ ad=7.36e+08 pd=154000 as=0 ps=0 
M5413 diff_4459000_1490000# diff_4416000_951000# diff_4435000_1490000# GND efet w=21000 l=12000
+ ad=-2.10197e+09 pd=438000 as=0 ps=0 
M5414 diff_4477000_1497000# diff_4477000_1497000# diff_4480000_1474000# GND efet w=14000 l=107000
+ ad=0 pd=0 as=3.9e+08 ps=80000 
M5415 diff_4531000_1616000# diff_4517000_1572000# diff_4517000_1572000# GND efet w=14000 l=21000
+ ad=0 pd=0 as=1.838e+09 ps=338000 
M5416 diff_4517000_1572000# diff_4532000_1475000# diff_4519000_1373000# GND efet w=51000 l=10000
+ ad=0 pd=0 as=-1.47397e+09 ps=472000 
M5417 diff_4672000_1727000# diff_4547000_2724000# diff_4607000_1699000# GND efet w=22000 l=12000
+ ad=4.4e+08 pd=84000 as=0 ps=0 
M5418 diff_4706000_1727000# diff_4601000_2751000# diff_4672000_1727000# GND efet w=22000 l=14000
+ ad=4.4e+08 pd=84000 as=0 ps=0 
M5419 diff_4753000_1809000# diff_4706000_1772000# diff_4726000_1760000# GND efet w=52000 l=10000
+ ad=0 pd=0 as=1.623e+09 ps=300000 
M5420 diff_4787000_1783000# diff_4739000_2640000# diff_4753000_1809000# GND efet w=149500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5421 diff_4574000_1652000# diff_4574000_1652000# diff_4588000_1617000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=1.522e+09 ps=174000 
M5422 diff_4607000_1699000# diff_4607000_1699000# diff_4588000_1617000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M5423 diff_4588000_1617000# diff_4574000_1573000# diff_4574000_1573000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=1.693e+09 ps=308000 
M5424 diff_4588000_1617000# diff_4607000_1470000# diff_4607000_1470000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=1.876e+09 ps=404000 
M5425 diff_4574000_1573000# diff_4497000_2491000# diff_4563000_1518000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=3.73e+08 ps=78000 
M5426 diff_4692000_1680000# diff_4692000_1680000# diff_4701000_1619000# GND efet w=15000 l=27000
+ ad=8.17e+08 pd=156000 as=1.919e+09 ps=196000 
M5427 diff_4726000_1760000# diff_4726000_1760000# diff_4701000_1619000# GND efet w=16000 l=27000
+ ad=0 pd=0 as=0 ps=0 
M5428 diff_4809000_1646000# diff_4799000_1639000# diff_4787000_1783000# GND efet w=128000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5429 diff_4831000_1646000# diff_4821000_1638000# diff_4809000_1646000# GND efet w=68500 l=10500
+ ad=-2.01297e+09 pd=388000 as=0 ps=0 
M5430 diff_4899000_1818000# diff_4893000_1829000# diff_4870000_1933000# GND efet w=60000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5431 diff_4951000_1858000# diff_4904000_1921000# diff_4899000_1818000# GND efet w=137000 l=10000
+ ad=1.233e+09 pd=292000 as=0 ps=0 
M5432 diff_4971000_1858000# diff_4905000_2664000# diff_4951000_1858000# GND efet w=137000 l=11000
+ ad=1.649e+09 pd=350000 as=0 ps=0 
M5433 diff_4991000_1833000# diff_4982000_1826000# diff_4971000_1858000# GND efet w=98000 l=9000
+ ad=-2.01097e+09 pd=396000 as=0 ps=0 
M5434 diff_5021000_2029000# diff_5021000_2029000# diff_5028000_1995000# GND efet w=15000 l=27000
+ ad=0 pd=0 as=6.82e+08 ps=110000 
M5435 diff_5068000_2031000# diff_5068000_2031000# diff_5074000_1993000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=1.488e+09 ps=180000 
M5436 diff_5124000_2368000# diff_5161000_2126000# diff_5124000_2017000# GND efet w=42000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5437 diff_5124000_2017000# diff_5136000_2101000# diff_5111000_2140000# GND efet w=23000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5438 diff_5124000_2368000# diff_5161000_2126000# diff_5124000_2017000# GND efet w=72000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5439 diff_5243000_2120000# diff_5233000_2294000# diff_5201000_2341000# GND efet w=72500 l=9500
+ ad=1.75203e+09 pd=966000 as=0 ps=0 
M5440 diff_5242000_2359000# diff_5201000_2341000# diff_5243000_2120000# GND efet w=65500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5441 diff_5289000_2222000# diff_5278000_2280000# diff_5242000_2359000# GND efet w=34000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5442 diff_5289000_2222000# diff_5281000_2212000# diff_5243000_2120000# GND efet w=117500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5443 diff_5200000_2037000# diff_5124000_2368000# diff_5202000_2119000# GND efet w=80000 l=10000
+ ad=1.544e+09 pd=340000 as=0 ps=0 
M5444 diff_5243000_2120000# diff_5233000_2092000# diff_5200000_2037000# GND efet w=72500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5445 diff_5243000_2120000# diff_5281000_2180000# diff_5289000_2044000# GND efet w=122000 l=11000
+ ad=0 pd=0 as=1.306e+09 ps=326000 
M5446 diff_5242000_2017000# diff_5200000_2037000# diff_5243000_2120000# GND efet w=65500 l=10500
+ ad=-1.97897e+09 pd=498000 as=0 ps=0 
M5447 diff_5289000_2044000# diff_5278000_2035000# diff_5242000_2017000# GND efet w=35000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5448 diff_5200000_2037000# diff_5200000_2037000# diff_5208000_1988000# GND efet w=15000 l=25000
+ ad=0 pd=0 as=1.544e+09 ps=184000 
M5449 diff_5124000_2017000# diff_4931000_826000# diff_5074000_1993000# GND efet w=15000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5450 diff_5289000_2044000# diff_5278000_2035000# diff_5242000_2017000# GND efet w=76000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5451 diff_5376000_2328000# diff_5376000_2328000# diff_5385000_2373000# GND efet w=15000 l=24000
+ ad=1.766e+09 pd=326000 as=7.18e+08 ps=114000 
M5452 diff_5376000_2328000# diff_5355000_2355000# diff_5358000_2058000# GND efet w=192000 l=10000
+ ad=0 pd=0 as=-9.34935e+08 ps=1.282e+06 
M5453 diff_5330000_4061000# diff_5376000_2328000# diff_5358000_2058000# GND efet w=157500 l=9500
+ ad=-1.02884e+09 pd=3.694e+06 as=0 ps=0 
M5454 diff_5465000_2330000# diff_5446000_801000# diff_5442000_2249000# GND efet w=88500 l=12500
+ ad=1.443e+09 pd=284000 as=9.09e+08 ps=210000 
M5455 diff_5376000_2057000# diff_5355000_2021000# diff_5358000_2058000# GND efet w=202000 l=11000
+ ad=1.795e+09 pd=304000 as=0 ps=0 
M5456 diff_5330000_4061000# diff_5376000_2057000# diff_5358000_2058000# GND efet w=156500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5457 diff_5242000_2017000# diff_5242000_2017000# diff_5208000_1988000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5458 diff_5335000_2021000# diff_5224000_815000# diff_5242000_2017000# GND efet w=21000 l=14000
+ ad=1.26e+08 pd=54000 as=0 ps=0 
M5459 diff_5355000_2021000# diff_5270000_856000# diff_5335000_2021000# GND efet w=21000 l=14000
+ ad=3.56e+08 pd=98000 as=0 ps=0 
M5460 diff_5376000_2057000# diff_5376000_2057000# diff_5385000_1996000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=1.292e+09 ps=152000 
M5461 diff_5465000_2048000# diff_5446000_801000# diff_5442000_2129000# GND efet w=88500 l=12500
+ ad=1.459e+09 pd=284000 as=9.09e+08 ps=210000 
M5462 diff_5537000_2618000# diff_5576000_2597000# diff_5650000_2540000# GND efet w=37000 l=14000
+ ad=0 pd=0 as=-1.39597e+09 ps=330000 
M5463 diff_82000_3097000# diff_5696000_2541000# diff_5618000_2892000# GND efet w=291000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5464 diff_82000_3097000# diff_5696000_2541000# diff_5618000_2892000# GND efet w=291500 l=12500
+ ad=0 pd=0 as=0 ps=0 
M5465 diff_5618000_2892000# diff_5696000_2541000# diff_82000_3097000# GND efet w=802500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M5466 diff_5695000_2525000# diff_5650000_2471000# diff_82000_3097000# GND efet w=518000 l=11000
+ ad=1.02207e+09 pd=1.816e+06 as=0 ps=0 
M5467 diff_82000_3097000# diff_5695000_2525000# diff_5618000_2171000# GND efet w=797500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M5468 diff_82000_3097000# diff_5751000_2392000# diff_5695000_2525000# GND efet w=476000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5469 diff_5650000_2471000# diff_5688000_2454000# diff_5562000_2269000# GND efet w=37000 l=13000
+ ad=-1.51497e+09 pd=300000 as=-1.77967e+08 ps=724000 
M5470 diff_5562000_2269000# diff_5633000_2428000# diff_5631000_2275000# GND efet w=89000 l=12000
+ ad=0 pd=0 as=-2.76967e+08 ps=748000 
M5471 diff_5631000_2275000# diff_5617000_2218000# diff_5619000_2361000# GND efet w=223000 l=10000
+ ad=0 pd=0 as=2.082e+09 ps=288000 
M5472 diff_82000_3097000# diff_5695000_2525000# diff_5618000_2171000# GND efet w=291500 l=12500
+ ad=0 pd=0 as=0 ps=0 
M5473 diff_82000_3097000# diff_5695000_2525000# diff_5618000_2171000# GND efet w=291000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5474 diff_5618000_2171000# diff_5695000_2525000# diff_82000_3097000# GND efet w=240500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M5475 diff_5695000_2525000# diff_5695000_2525000# diff_5695000_2525000# GND efet w=3000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5476 diff_5695000_2525000# diff_5695000_2525000# diff_94000_5193000# GND efet w=38000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5477 diff_5028000_1995000# diff_5021000_1967000# diff_5021000_1967000# GND efet w=15000 l=28000
+ ad=0 pd=0 as=1.88e+09 ps=296000 
M5478 diff_5074000_1993000# diff_5068000_1971000# diff_5068000_1971000# GND efet w=15000 l=22000
+ ad=0 pd=0 as=1.626e+09 ps=362000 
M5479 diff_5124000_1991000# diff_4931000_826000# diff_5074000_1993000# GND efet w=14000 l=10000
+ ad=4.20327e+07 pd=876000 as=0 ps=0 
M5480 diff_5124000_2017000# diff_5151000_1994000# diff_5124000_1991000# GND efet w=130500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M5481 diff_4899000_1818000# diff_4893000_1809000# diff_4869000_1704000# GND efet w=61000 l=10000
+ ad=0 pd=0 as=-1.24097e+09 ps=472000 
M5482 diff_4866000_1738000# diff_4838000_2617000# diff_4831000_1646000# GND efet w=52000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5483 diff_4991000_1833000# diff_4982000_1826000# diff_4971000_1858000# GND efet w=35000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5484 diff_5024000_1733000# diff_4993000_2633000# diff_4991000_1833000# GND efet w=57000 l=11000
+ ad=-1.58197e+09 pd=420000 as=0 ps=0 
M5485 diff_5021000_1967000# diff_5037000_1886000# diff_5024000_1733000# GND efet w=46000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5486 diff_5124000_1991000# diff_5132000_1970000# diff_5111000_1762000# GND efet w=91500 l=12500
+ ad=0 pd=0 as=-1.67293e+09 ps=808000 
M5487 diff_5068000_1971000# diff_5068000_1909000# diff_5070000_1741000# GND efet w=67500 l=10500
+ ad=0 pd=0 as=1.874e+09 ps=374000 
M5488 diff_5111000_1762000# diff_4931000_826000# diff_5068000_1971000# GND efet w=68000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5489 diff_5208000_1988000# diff_5201000_1963000# diff_5201000_1963000# GND efet w=15000 l=25000
+ ad=0 pd=0 as=1.612e+09 ps=346000 
M5490 diff_5242000_1982000# diff_5242000_1982000# diff_5208000_1988000# GND efet w=14000 l=23000
+ ad=-2.10097e+09 pd=496000 as=0 ps=0 
M5491 diff_5289000_1845000# diff_5278000_1902000# diff_5242000_1982000# GND efet w=78500 l=10500
+ ad=1.279e+09 pd=322000 as=0 ps=0 
M5492 diff_4831000_1646000# diff_4821000_1638000# diff_4809000_1646000# GND efet w=70000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5493 diff_4869000_1704000# diff_4838000_2617000# diff_4866000_1738000# GND efet w=60500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5494 diff_4701000_1619000# diff_4693000_1562000# diff_4693000_1562000# GND efet w=15000 l=26000
+ ad=0 pd=0 as=8.39e+08 ps=158000 
M5495 diff_4701000_1619000# diff_4726000_1482000# diff_4726000_1482000# GND efet w=15000 l=26000
+ ad=0 pd=0 as=1.673e+09 ps=300000 
M5496 diff_4379000_1393000# diff_4347000_2438000# diff_4354000_1418000# GND efet w=104500 l=10500
+ ad=1.155e+09 pd=222000 as=0 ps=0 
M5497 diff_4317000_998000# diff_4319000_1315000# diff_4245000_1443000# GND efet w=54500 l=10500
+ ad=6.71e+08 pd=144000 as=0 ps=0 
M5498 diff_4245000_1443000# diff_4276000_1307000# diff_4262000_1287000# GND efet w=85000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5499 diff_4228000_1258000# diff_4224000_1220000# diff_4224000_1220000# GND efet w=14000 l=37000
+ ad=3.34e+08 pd=74000 as=-1.50197e+09 ps=394000 
M5500 diff_4317000_998000# diff_4317000_998000# diff_4314000_1211000# GND efet w=14000 l=39000
+ ad=0 pd=0 as=1.298e+09 ps=174000 
M5501 diff_4314000_1211000# diff_4306000_1186000# diff_4306000_1186000# GND efet w=15000 l=25000
+ ad=0 pd=0 as=-1.72197e+09 ps=436000 
M5502 diff_4067000_1029000# diff_4056000_1019000# diff_82000_3097000# GND efet w=206500 l=9500
+ ad=-1.42197e+09 pd=472000 as=0 ps=0 
M5503 diff_82000_3097000# diff_4037000_919000# diff_4057000_979000# GND efet w=63000 l=10000
+ ad=0 pd=0 as=1.003e+09 ps=180000 
M5504 diff_4149000_968000# diff_4107000_2724000# diff_4067000_1029000# GND efet w=89000 l=11000
+ ad=1.145e+09 pd=216000 as=0 ps=0 
M5505 diff_4204000_1036000# diff_4192000_1025000# diff_4185000_1075000# GND efet w=107000 l=12000
+ ad=-1.11797e+09 pd=460000 as=0 ps=0 
M5506 diff_4262000_1287000# diff_4232000_995000# diff_4224000_1220000# GND efet w=111000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5507 diff_4204000_1036000# diff_4192000_1025000# diff_4184000_1005000# GND efet w=106500 l=11500
+ ad=0 pd=0 as=1.737e+09 ps=368000 
M5508 diff_3886000_876000# diff_3884000_904000# diff_3881000_929000# GND efet w=13000 l=24000
+ ad=5.38e+08 pd=96000 as=0 ps=0 
M5509 diff_3938000_928000# diff_3884000_904000# diff_3881000_929000# GND efet w=13500 l=82500
+ ad=8.5e+08 pd=254000 as=0 ps=0 
M5510 diff_3586000_784000# diff_3526000_822000# diff_3566000_784000# GND efet w=72000 l=11000
+ ad=-2.13997e+09 pd=310000 as=0 ps=0 
M5511 diff_3595000_2394000# diff_3604000_815000# diff_3586000_784000# GND efet w=95500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M5512 diff_3664000_845000# diff_3604000_815000# diff_3353000_2408000# GND efet w=72500 l=11500
+ ad=1.622e+09 pd=222000 as=0 ps=0 
M5513 diff_3488000_2724000# diff_3604000_815000# diff_3664000_845000# GND efet w=72000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5514 diff_3741000_766000# diff_3717000_755000# diff_3738000_825000# GND efet w=79000 l=12000
+ ad=1.865e+09 pd=248000 as=0 ps=0 
M5515 diff_3801000_831000# diff_3717000_755000# diff_3741000_766000# GND efet w=76000 l=12000
+ ad=1.633e+09 pd=258000 as=0 ps=0 
M5516 diff_3949000_962000# diff_3884000_904000# diff_3960000_872000# GND efet w=14000 l=35000
+ ad=0 pd=0 as=4.2e+08 ps=84000 
M5517 diff_4005000_919000# diff_3921000_785000# diff_3938000_928000# GND efet w=22000 l=12000
+ ad=4.4e+08 pd=84000 as=0 ps=0 
M5518 diff_4037000_919000# diff_4003000_2724000# diff_4005000_919000# GND efet w=22000 l=12000
+ ad=9.19e+08 pd=240000 as=0 ps=0 
M5519 diff_4057000_979000# diff_4052000_893000# diff_4052000_838000# GND efet w=14000 l=35000
+ ad=0 pd=0 as=9.66e+08 ps=152000 
M5520 diff_4067000_1029000# diff_4052000_893000# diff_4037000_919000# GND efet w=14000 l=83000
+ ad=0 pd=0 as=0 ps=0 
M5521 diff_3856000_786000# diff_3836000_763000# diff_3829000_786000# GND efet w=72000 l=12000
+ ad=1.311e+09 pd=194000 as=0 ps=0 
M5522 diff_3694000_2724000# diff_3836000_763000# diff_3856000_786000# GND efet w=98500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5523 diff_4067000_1029000# diff_4052000_893000# diff_4126000_876000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=5.39e+08 ps=96000 
M5524 diff_4184000_1005000# diff_4162000_2432000# diff_4165000_930000# GND efet w=88000 l=12000
+ ad=0 pd=0 as=8.08e+08 ps=210000 
M5525 diff_4308000_1009000# diff_4288000_1116000# diff_4280000_938000# GND efet w=103000 l=10000
+ ad=9.27e+08 pd=224000 as=-1.34693e+09 ps=702000 
M5526 diff_4306000_1186000# diff_4317000_998000# diff_4308000_1009000# GND efet w=103000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5527 diff_4481000_1400000# diff_4477000_1119000# diff_4477000_1119000# GND efet w=14000 l=106000
+ ad=3.34e+08 pd=74000 as=1.164e+09 ps=200000 
M5528 diff_4517000_1277000# diff_4532000_1332000# diff_4519000_1373000# GND efet w=51000 l=10000
+ ad=1.791e+09 pd=334000 as=0 ps=0 
M5529 diff_4617000_1363000# diff_4607000_1470000# diff_4574000_1573000# GND efet w=50000 l=10000
+ ad=-1.43197e+09 pd=388000 as=0 ps=0 
M5530 diff_4607000_1470000# diff_4624000_1532000# diff_4617000_1363000# GND efet w=68000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5531 diff_4672000_1518000# diff_4547000_2724000# diff_4607000_1470000# GND efet w=23000 l=12000
+ ad=4.6e+08 pd=86000 as=0 ps=0 
M5532 diff_4706000_1518000# diff_4601000_2751000# diff_4672000_1518000# GND efet w=23000 l=14000
+ ad=4.37e+08 pd=84000 as=0 ps=0 
M5533 diff_4574000_1276000# diff_4497000_2491000# diff_4563000_1352000# GND efet w=23000 l=12000
+ ad=1.673e+09 pd=302000 as=3.91e+08 ps=80000 
M5534 diff_4617000_1363000# diff_4607000_1322000# diff_4574000_1276000# GND efet w=52000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5535 diff_4607000_1322000# diff_4624000_1339000# diff_4617000_1363000# GND efet w=69000 l=10000
+ ad=1.852e+09 pd=402000 as=0 ps=0 
M5536 diff_4706000_1474000# diff_4601000_2751000# diff_4675000_1474000# GND efet w=22000 l=14000
+ ad=5.13e+08 pd=146000 as=3.74e+08 ps=78000 
M5537 diff_4753000_1432000# diff_4706000_1474000# diff_4726000_1482000# GND efet w=52000 l=10000
+ ad=1.63303e+09 pd=784000 as=0 ps=0 
M5538 diff_4787000_1475000# diff_4739000_2640000# diff_4753000_1432000# GND efet w=150500 l=10500
+ ad=1.658e+09 pd=366000 as=0 ps=0 
M5539 diff_4809000_1516000# diff_4798000_1507000# diff_4787000_1475000# GND efet w=128000 l=11000
+ ad=2.114e+09 pd=412000 as=0 ps=0 
M5540 diff_4831000_1552000# diff_4820000_1527000# diff_4809000_1516000# GND efet w=71000 l=11000
+ ad=-1.95697e+09 pd=394000 as=0 ps=0 
M5541 diff_4899000_1818000# diff_4904000_1705000# diff_4869000_1704000# GND efet w=55000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5542 diff_4869000_1704000# diff_4869000_1704000# diff_4881000_1621000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=6.49e+08 ps=108000 
M5543 diff_4952000_1650000# diff_4904000_1705000# diff_4899000_1818000# GND efet w=137000 l=11000
+ ad=1.096e+09 pd=290000 as=0 ps=0 
M5544 diff_4971000_1650000# diff_4905000_2664000# diff_4952000_1650000# GND efet w=137000 l=11000
+ ad=1.649e+09 pd=350000 as=0 ps=0 
M5545 diff_4991000_1650000# diff_4982000_1643000# diff_4971000_1650000# GND efet w=34000 l=9000
+ ad=-2.08597e+09 pd=396000 as=0 ps=0 
M5546 diff_5335000_1977000# diff_5224000_815000# diff_5242000_1982000# GND efet w=23000 l=14000
+ ad=1.38e+08 pd=58000 as=0 ps=0 
M5547 diff_5355000_1977000# diff_5270000_856000# diff_5335000_1977000# GND efet w=23000 l=14000
+ ad=3.45e+08 pd=112000 as=0 ps=0 
M5548 diff_5124000_1991000# diff_5132000_1970000# diff_5111000_1762000# GND efet w=50000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5549 diff_5201000_1963000# diff_5124000_2017000# diff_5202000_1742000# GND efet w=79000 l=10000
+ ad=0 pd=0 as=1.906e+09 ps=362000 
M5550 diff_5124000_1640000# diff_5136000_1724000# diff_5111000_1762000# GND efet w=125000 l=11000
+ ad=-1.69797e+09 pd=500000 as=0 ps=0 
M5551 diff_4991000_1650000# diff_4982000_1643000# diff_4971000_1650000# GND efet w=99000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5552 diff_5024000_1733000# diff_4993000_2633000# diff_4991000_1650000# GND efet w=56000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5553 diff_5021000_1652000# diff_5037000_1727000# diff_5024000_1733000# GND efet w=47000 l=8000
+ ad=1.8e+09 pd=296000 as=0 ps=0 
M5554 diff_5068000_1654000# diff_5068000_1716000# diff_5070000_1741000# GND efet w=66500 l=10500
+ ad=1.762e+09 pd=362000 as=0 ps=0 
M5555 diff_5111000_1762000# diff_4931000_826000# diff_5068000_1654000# GND efet w=67500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5556 diff_4881000_1621000# diff_4870000_1558000# diff_4870000_1558000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=-1.40597e+09 ps=458000 
M5557 diff_4899000_1441000# diff_4904000_1545000# diff_4870000_1558000# GND efet w=53000 l=10000
+ ad=6.35033e+08 pd=812000 as=0 ps=0 
M5558 diff_4870000_1558000# diff_4838000_2617000# diff_4866000_1360000# GND efet w=63500 l=10500
+ ad=0 pd=0 as=-1.16697e+09 ps=460000 
M5559 diff_4831000_1552000# diff_4820000_1527000# diff_4809000_1516000# GND efet w=70500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5560 diff_4706000_1395000# diff_4601000_2751000# diff_4675000_1395000# GND efet w=23000 l=14000
+ ad=5.16e+08 pd=146000 as=3.91e+08 ps=80000 
M5561 diff_4809000_1516000# diff_4798000_1507000# diff_4787000_1475000# GND efet w=14000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5562 diff_4866000_1360000# diff_4838000_2617000# diff_4831000_1552000# GND efet w=53000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5563 diff_4809000_1268000# diff_4799000_1262000# diff_4787000_1407000# GND efet w=12000 l=10000
+ ad=2.039e+09 pd=412000 as=1.611e+09 ps=368000 
M5564 diff_4517000_1277000# diff_4517000_1277000# diff_4531000_1239000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=7.81e+08 ps=120000 
M5565 diff_4432000_1347000# diff_4373000_832000# diff_4406000_1189000# GND efet w=22000 l=11000
+ ad=1.589e+09 pd=306000 as=1.435e+09 ps=266000 
M5566 diff_4458000_1182000# diff_4416000_951000# diff_4432000_1347000# GND efet w=22000 l=12000
+ ad=9.97e+08 pd=190000 as=0 ps=0 
M5567 diff_4378000_1100000# diff_4347000_2438000# diff_4354000_1418000# GND efet w=102500 l=10500
+ ad=1.175e+09 pd=222000 as=0 ps=0 
M5568 diff_4433000_1143000# diff_4373000_832000# diff_4406000_1189000# GND efet w=23000 l=11000
+ ad=8.9e+08 pd=166000 as=0 ps=0 
M5569 diff_4379000_974000# diff_4347000_2438000# diff_4354000_1418000# GND efet w=89000 l=11000
+ ad=1.115e+09 pd=204000 as=0 ps=0 
M5570 diff_3947000_785000# diff_3930000_764000# diff_3921000_785000# GND efet w=104500 l=11500
+ ad=1.758e+09 pd=258000 as=0 ps=0 
M5571 diff_1757000_612000# diff_1757000_612000# diff_1757000_699000# GND efet w=18000 l=10000
+ ad=-4.82967e+08 pd=644000 as=4.21e+08 ps=84000 
M5572 diff_1778000_637000# diff_1756000_738000# diff_1757000_612000# GND efet w=233000 l=10000
+ ad=-1.63797e+09 pd=316000 as=0 ps=0 
M5573 diff_1693000_584000# diff_1693000_584000# diff_1844000_692000# GND efet w=52500 l=9500
+ ad=-5.76902e+08 pd=2.026e+06 as=4.6e+08 ps=86000 
M5574 diff_1850000_578000# diff_1843000_567000# diff_1693000_584000# GND efet w=487500 l=10500
+ ad=-1.54697e+09 pd=504000 as=0 ps=0 
M5575 diff_1719000_540000# diff_1619000_122000# diff_1619000_122000# GND efet w=38000 l=10000
+ ad=7.21e+08 pd=114000 as=0 ps=0 
M5576 diff_1843000_567000# diff_1833000_667000# diff_1757000_612000# GND efet w=37000 l=13000
+ ad=8.06e+08 pd=184000 as=0 ps=0 
M5577 diff_1941000_635000# diff_1930000_625000# diff_1693000_584000# GND efet w=439000 l=10000
+ ad=-1.10497e+09 pd=452000 as=0 ps=0 
M5578 diff_1619000_122000# diff_1693000_584000# diff_1753000_545000# GND efet w=46000 l=11000
+ ad=0 pd=0 as=1.935e+09 ps=306000 
M5579 diff_2116000_578000# diff_2107000_567000# diff_2034000_544000# GND efet w=489500 l=10500
+ ad=-1.43997e+09 pd=504000 as=-6.92902e+08 ps=2.032e+06 
M5580 diff_2059000_661000# diff_2049000_625000# diff_2034000_544000# GND efet w=439000 l=10000
+ ad=-1.17297e+09 pd=456000 as=0 ps=0 
M5581 diff_2191000_692000# diff_2034000_544000# diff_2034000_544000# GND efet w=54500 l=9500
+ ad=5e+08 pd=90000 as=0 ps=0 
M5582 diff_2236000_651000# diff_2228000_597000# diff_2215000_624000# GND efet w=233500 l=10500
+ ad=-1.81997e+09 pd=316000 as=-4.24967e+08 ps=646000 
M5583 diff_2283000_699000# diff_2215000_624000# diff_2215000_624000# GND efet w=18000 l=10000
+ ad=4.61e+08 pd=88000 as=0 ps=0 
M5584 diff_2215000_624000# diff_2202000_619000# diff_2107000_567000# GND efet w=37000 l=13000
+ ad=0 pd=0 as=7.3e+08 ps=182000 
M5585 diff_2333000_592000# diff_2034000_544000# diff_2260000_566000# GND efet w=276000 l=10000
+ ad=-2.05297e+09 pd=280000 as=1.92807e+09 ps=1.504e+06 
M5586 diff_2377000_715000# diff_2367000_705000# diff_2260000_566000# GND efet w=301500 l=10500
+ ad=-8.87967e+08 pd=438000 as=0 ps=0 
M5587 diff_2260000_566000# diff_2034000_544000# diff_2260000_545000# GND efet w=47000 l=11000
+ ad=0 pd=0 as=2.01e+09 ps=304000 
M5588 diff_1506000_490000# diff_1429000_566000# diff_1219000_196000# GND efet w=185500 l=10500
+ ad=1.195e+09 pd=186000 as=0 ps=0 
M5589 diff_1465000_100000# diff_1429000_566000# diff_1219000_196000# GND efet w=184000 l=10000
+ ad=1.86716e+09 pd=2.898e+06 as=0 ps=0 
M5590 diff_1628000_457000# diff_1619000_122000# diff_1465000_100000# GND efet w=184000 l=10000
+ ad=-1.81571e+09 pd=4.532e+06 as=0 ps=0 
M5591 diff_1465000_100000# diff_1429000_566000# diff_1219000_196000# GND efet w=651500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5592 diff_1699000_492000# diff_1619000_122000# diff_1628000_457000# GND efet w=186000 l=10000
+ ad=1.229e+09 pd=188000 as=0 ps=0 
M5593 diff_1049000_100000# diff_968000_455000# diff_802000_365000# GND efet w=525000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5594 diff_802000_365000# diff_968000_455000# diff_1049000_100000# GND efet w=262000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5595 diff_1219000_196000# diff_1203000_545000# diff_1049000_100000# GND efet w=270500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5596 diff_1628000_457000# diff_1619000_122000# diff_1465000_100000# GND efet w=649500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5597 diff_1753000_545000# diff_1619000_122000# diff_1628000_457000# GND efet w=193500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5598 diff_1809000_491000# diff_1693000_584000# diff_1628000_457000# GND efet w=210000 l=10000
+ ad=1.369e+09 pd=208000 as=0 ps=0 
M5599 diff_1862000_492000# diff_1693000_584000# diff_1628000_457000# GND efet w=205500 l=10500
+ ad=1.36e+09 pd=204000 as=0 ps=0 
M5600 diff_1915000_492000# diff_1693000_584000# diff_1628000_457000# GND efet w=205500 l=10500
+ ad=1.36e+09 pd=204000 as=0 ps=0 
M5601 diff_1873000_101000# diff_1693000_584000# diff_1628000_457000# GND efet w=191500 l=10500
+ ad=-1.63877e+09 pd=2.932e+06 as=0 ps=0 
M5602 diff_2050000_195000# diff_2034000_544000# diff_1873000_101000# GND efet w=193000 l=10000
+ ad=-2.05171e+09 pd=4.538e+06 as=0 ps=0 
M5603 diff_1873000_101000# diff_1693000_584000# diff_1628000_457000# GND efet w=652000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5604 diff_2122000_492000# diff_2034000_544000# diff_2050000_195000# GND efet w=205500 l=10500
+ ad=1.328e+09 pd=204000 as=0 ps=0 
M5605 diff_2050000_195000# diff_2034000_544000# diff_1873000_101000# GND efet w=652000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5606 diff_1219000_196000# diff_1429000_566000# diff_1465000_100000# GND efet w=282000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5607 diff_1628000_457000# diff_1619000_122000# diff_1465000_100000# GND efet w=282000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5608 diff_2176000_491000# diff_2034000_544000# diff_2050000_195000# GND efet w=205500 l=10500
+ ad=1.36e+09 pd=204000 as=0 ps=0 
M5609 diff_2228000_491000# diff_2034000_544000# diff_2050000_195000# GND efet w=210000 l=10000
+ ad=1.337e+09 pd=208000 as=0 ps=0 
M5610 diff_2260000_566000# diff_2260000_566000# diff_2321000_541000# GND efet w=37000 l=10000
+ ad=0 pd=0 as=6.66e+08 ps=110000 
M5611 diff_2260000_566000# diff_2367000_705000# diff_2377000_715000# GND efet w=58000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5612 diff_2260000_545000# diff_2260000_566000# diff_2050000_195000# GND efet w=193500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5613 diff_2472000_566000# diff_2461000_557000# diff_2449000_122000# GND efet w=58000 l=10000
+ ad=-9.83967e+08 pd=440000 as=1.89807e+09 ps=1.5e+06 
M5614 diff_2472000_566000# diff_2461000_557000# diff_2449000_122000# GND efet w=301500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5615 diff_2534000_589000# diff_2523000_584000# diff_2449000_122000# GND efet w=276000 l=11000
+ ad=-2.13697e+09 pd=278000 as=0 ps=0 
M5616 diff_2588000_612000# diff_2588000_612000# diff_2587000_700000# GND efet w=18000 l=10000
+ ad=-6.16967e+08 pd=644000 as=4.24e+08 ps=84000 
M5617 diff_2608000_637000# diff_2598000_626000# diff_2588000_612000# GND efet w=233500 l=10500
+ ad=-1.66197e+09 pd=316000 as=0 ps=0 
M5618 diff_2523000_584000# diff_2523000_584000# diff_2675000_692000# GND efet w=52000 l=10000
+ ad=-6.84902e+08 pd=2.026e+06 as=4.4e+08 ps=84000 
M5619 diff_2681000_578000# diff_2673000_567000# diff_2523000_584000# GND efet w=485500 l=10500
+ ad=-1.58397e+09 pd=500000 as=0 ps=0 
M5620 diff_2549000_541000# diff_2449000_122000# diff_2449000_122000# GND efet w=36000 l=10000
+ ad=7.2e+08 pd=112000 as=0 ps=0 
M5621 diff_2673000_567000# diff_2664000_667000# diff_2588000_612000# GND efet w=37000 l=14000
+ ad=7.36e+08 pd=182000 as=0 ps=0 
M5622 diff_2771000_635000# diff_2760000_625000# diff_2523000_584000# GND efet w=441000 l=10000
+ ad=-9.89967e+08 pd=456000 as=0 ps=0 
M5623 diff_2449000_122000# diff_2523000_584000# diff_2583000_545000# GND efet w=47000 l=11000
+ ad=0 pd=0 as=1.991e+09 ps=306000 
M5624 diff_3279000_567000# diff_3269000_556000# diff_3257000_122000# GND efet w=58000 l=11000
+ ad=-8.66967e+08 pd=440000 as=1.67707e+09 ps=1.496e+06 
M5625 diff_3279000_567000# diff_3269000_556000# diff_3257000_122000# GND efet w=304000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5626 diff_3341000_590000# diff_3331000_584000# diff_3257000_122000# GND efet w=274000 l=10000
+ ad=-2.06597e+09 pd=278000 as=0 ps=0 
M5627 diff_2336000_490000# diff_2260000_566000# diff_2050000_195000# GND efet w=186500 l=10500
+ ad=1.231e+09 pd=188000 as=0 ps=0 
M5628 diff_2295000_101000# diff_2260000_566000# diff_2050000_195000# GND efet w=183000 l=10000
+ ad=1.65216e+09 pd=2.898e+06 as=0 ps=0 
M5629 diff_2459000_132000# diff_2449000_122000# diff_2295000_101000# GND efet w=185000 l=10000
+ ad=-1.61771e+09 pd=4.536e+06 as=0 ps=0 
M5630 diff_2295000_101000# diff_2260000_566000# diff_2050000_195000# GND efet w=648500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5631 diff_2530000_491000# diff_2449000_122000# diff_2459000_132000# GND efet w=186500 l=10500
+ ad=1.228e+09 pd=188000 as=0 ps=0 
M5632 diff_2459000_132000# diff_2449000_122000# diff_2295000_101000# GND efet w=650500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5633 diff_2583000_545000# diff_2449000_122000# diff_2459000_132000# GND efet w=193000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5634 diff_2639000_491000# diff_2523000_584000# diff_2459000_132000# GND efet w=210000 l=10000
+ ad=1.37e+09 pd=208000 as=0 ps=0 
M5635 diff_2693000_491000# diff_2523000_584000# diff_2459000_132000# GND efet w=205500 l=10500
+ ad=1.331e+09 pd=204000 as=0 ps=0 
M5636 diff_2746000_491000# diff_2523000_584000# diff_2459000_132000# GND efet w=205500 l=10500
+ ad=1.364e+09 pd=204000 as=0 ps=0 
M5637 diff_2705000_101000# diff_2523000_584000# diff_2459000_132000# GND efet w=191000 l=10000
+ ad=-1.05887e+09 pd=1.9e+06 as=0 ps=0 
M5638 diff_2705000_101000# diff_2523000_584000# diff_2459000_132000# GND efet w=648000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5639 diff_4003000_2724000# diff_3993000_764000# diff_3947000_785000# GND efet w=71000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5640 diff_4073000_749000# diff_4046000_762000# diff_4044000_822000# GND efet w=113000 l=10000
+ ad=-2.04097e+09 pd=314000 as=1.956e+09 ps=304000 
M5641 diff_4052000_838000# diff_4044000_822000# diff_4044000_822000# GND efet w=15000 l=17000
+ ad=0 pd=0 as=0 ps=0 
M5642 diff_4107000_2724000# diff_4120000_825000# diff_4073000_749000# GND efet w=76500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M5643 diff_4194000_784000# diff_4182000_762000# diff_4162000_2432000# GND efet w=76000 l=12000
+ ad=1.285e+09 pd=188000 as=9.34e+08 ps=204000 
M5644 diff_4192000_1025000# diff_4182000_762000# diff_4194000_784000# GND efet w=77000 l=12000
+ ad=1.009e+09 pd=208000 as=0 ps=0 
M5645 diff_4329000_909000# diff_4317000_839000# diff_4280000_938000# GND efet w=74000 l=12000
+ ad=1.406e+09 pd=186000 as=0 ps=0 
M5646 diff_4460000_935000# diff_4416000_951000# diff_4433000_1143000# GND efet w=23000 l=10000
+ ad=-2.14697e+09 pd=428000 as=0 ps=0 
M5647 diff_4477000_1119000# diff_4477000_1119000# diff_4480000_1097000# GND efet w=14000 l=106000
+ ad=0 pd=0 as=3.86e+08 ps=80000 
M5648 diff_4531000_1239000# diff_4517000_1195000# diff_4517000_1195000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=1.854e+09 ps=336000 
M5649 diff_4517000_1195000# diff_4532000_1098000# diff_4519000_996000# GND efet w=51000 l=10000
+ ad=0 pd=0 as=-1.48897e+09 ps=470000 
M5650 diff_4672000_1350000# diff_4547000_2724000# diff_4607000_1322000# GND efet w=22000 l=12000
+ ad=4.4e+08 pd=84000 as=0 ps=0 
M5651 diff_4706000_1350000# diff_4601000_2751000# diff_4672000_1350000# GND efet w=22000 l=14000
+ ad=4.4e+08 pd=84000 as=0 ps=0 
M5652 diff_4753000_1432000# diff_4706000_1395000# diff_4726000_1382000# GND efet w=52000 l=10000
+ ad=0 pd=0 as=1.622e+09 ps=300000 
M5653 diff_4787000_1407000# diff_4739000_2640000# diff_4753000_1432000# GND efet w=150000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5654 diff_4574000_1276000# diff_4574000_1276000# diff_4588000_1240000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=1.566e+09 ps=180000 
M5655 diff_4607000_1322000# diff_4607000_1322000# diff_4588000_1240000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M5656 diff_4588000_1240000# diff_4574000_1196000# diff_4574000_1196000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=1.676e+09 ps=300000 
M5657 diff_4588000_1240000# diff_4607000_1092000# diff_4607000_1092000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=1.865e+09 ps=400000 
M5658 diff_4574000_1196000# diff_4497000_2491000# diff_4563000_1140000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=3.74e+08 ps=78000 
M5659 diff_4692000_1303000# diff_4692000_1303000# diff_4701000_1242000# GND efet w=15000 l=27000
+ ad=7.8e+08 pd=154000 as=1.918e+09 ps=202000 
M5660 diff_4726000_1382000# diff_4726000_1382000# diff_4701000_1242000# GND efet w=16000 l=26000
+ ad=0 pd=0 as=0 ps=0 
M5661 diff_4809000_1268000# diff_4799000_1262000# diff_4787000_1407000# GND efet w=128000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5662 diff_4831000_1268000# diff_4820000_1262000# diff_4809000_1268000# GND efet w=68500 l=10500
+ ad=-1.99897e+09 pd=390000 as=0 ps=0 
M5663 diff_4899000_1441000# diff_4893000_1452000# diff_4870000_1558000# GND efet w=60000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5664 diff_4951000_1481000# diff_4904000_1545000# diff_4899000_1441000# GND efet w=136000 l=10000
+ ad=1.224e+09 pd=290000 as=0 ps=0 
M5665 diff_4971000_1481000# diff_4905000_2664000# diff_4951000_1481000# GND efet w=136000 l=11000
+ ad=1.639e+09 pd=348000 as=0 ps=0 
M5666 diff_4991000_1456000# diff_4982000_1450000# diff_4971000_1481000# GND efet w=97000 l=9000
+ ad=-2.03097e+09 pd=394000 as=0 ps=0 
M5667 diff_5021000_1652000# diff_5021000_1652000# diff_5028000_1618000# GND efet w=15000 l=27000
+ ad=0 pd=0 as=6.86e+08 ps=110000 
M5668 diff_5068000_1654000# diff_5068000_1654000# diff_5074000_1617000# GND efet w=14000 l=21000
+ ad=0 pd=0 as=1.495e+09 ps=178000 
M5669 diff_5124000_1991000# diff_5161000_1749000# diff_5124000_1640000# GND efet w=43000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5670 diff_5124000_1640000# diff_5136000_1724000# diff_5111000_1762000# GND efet w=23000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5671 diff_5124000_1991000# diff_5161000_1749000# diff_5124000_1640000# GND efet w=73000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5672 diff_5243000_1742000# diff_5233000_1916000# diff_5201000_1963000# GND efet w=72500 l=9500
+ ad=1.75003e+09 pd=966000 as=0 ps=0 
M5673 diff_5242000_1982000# diff_5201000_1963000# diff_5243000_1742000# GND efet w=65500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5674 diff_5289000_1845000# diff_5278000_1902000# diff_5242000_1982000# GND efet w=34000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5675 diff_5289000_1845000# diff_5281000_1835000# diff_5243000_1742000# GND efet w=117500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5676 diff_5200000_1659000# diff_5124000_1991000# diff_5202000_1742000# GND efet w=80000 l=10000
+ ad=1.554e+09 pd=342000 as=0 ps=0 
M5677 diff_5243000_1742000# diff_5233000_1714000# diff_5200000_1659000# GND efet w=73500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5678 diff_5243000_1742000# diff_5281000_1802000# diff_5289000_1667000# GND efet w=121500 l=11500
+ ad=0 pd=0 as=1.293e+09 ps=324000 
M5679 diff_5242000_1640000# diff_5200000_1659000# diff_5243000_1742000# GND efet w=65500 l=10500
+ ad=-2.00497e+09 pd=498000 as=0 ps=0 
M5680 diff_5289000_1667000# diff_5278000_1658000# diff_5242000_1640000# GND efet w=35000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5681 diff_5200000_1659000# diff_5200000_1659000# diff_5208000_1611000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=1.544e+09 ps=184000 
M5682 diff_5124000_1640000# diff_4931000_826000# diff_5074000_1617000# GND efet w=15000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5683 diff_5289000_1667000# diff_5278000_1658000# diff_5242000_1640000# GND efet w=76500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5684 diff_5385000_1996000# diff_5376000_1951000# diff_5376000_1951000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=1.777e+09 ps=328000 
M5685 diff_5376000_1951000# diff_5355000_1977000# diff_5358000_1681000# GND efet w=193000 l=10000
+ ad=0 pd=0 as=-9.05935e+08 ps=1.28e+06 
M5686 diff_5330000_4061000# diff_5376000_1951000# diff_5358000_1681000# GND efet w=157500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5687 diff_5520000_2087000# diff_5510000_2076000# diff_5171000_2829000# GND efet w=105500 l=10500
+ ad=1.608e+09 pd=202000 as=0 ps=0 
M5688 diff_5171000_2829000# diff_5171000_2829000# diff_5476000_1993000# GND efet w=14000 l=17000
+ ad=0 pd=0 as=-1.93697e+09 ps=238000 
M5689 diff_5465000_1953000# diff_5446000_801000# diff_5442000_1872000# GND efet w=90000 l=13000
+ ad=1.453e+09 pd=286000 as=9.02e+08 ps=212000 
M5690 diff_5476000_1993000# diff_5472000_1599000# diff_5472000_1599000# GND efet w=14000 l=16000
+ ad=0 pd=0 as=1.838e+09 ps=368000 
M5691 diff_5472000_1599000# diff_5472000_1599000# diff_5472000_1599000# GND efet w=1500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5692 diff_5376000_1680000# diff_5355000_1644000# diff_5358000_1681000# GND efet w=200500 l=10500
+ ad=1.801e+09 pd=306000 as=0 ps=0 
M5693 diff_5330000_4061000# diff_5376000_1680000# diff_5358000_1681000# GND efet w=156500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5694 diff_5472000_1599000# diff_5484000_1775000# diff_5476000_1801000# GND efet w=98000 l=10000
+ ad=0 pd=0 as=1.266e+09 ps=234000 
M5695 diff_94000_5193000# diff_5631000_2275000# diff_5631000_2275000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M5696 diff_5654000_2314000# diff_5645000_2303000# diff_5652000_2258000# GND efet w=30000 l=11000
+ ad=4.8e+08 pd=92000 as=1.182e+09 ps=212000 
M5697 diff_94000_5193000# diff_5768000_2160000# diff_5768000_2160000# GND efet w=46000 l=11000
+ ad=0 pd=0 as=6.80065e+08 ps=1.636e+06 
M5698 diff_82000_3097000# diff_5695000_2525000# diff_5768000_2160000# GND efet w=480000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5699 diff_5618000_2171000# diff_5768000_2160000# diff_94000_5193000# GND efet w=288000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5700 diff_5631000_2275000# diff_5631000_2275000# diff_5631000_2275000# GND efet w=2000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5701 diff_5956000_2270000# diff_5768000_2160000# diff_5618000_2171000# GND efet w=287500 l=10500
+ ad=2.047e+09 pd=282000 as=0 ps=0 
M5702 diff_5652000_2258000# diff_5631000_2275000# diff_5630000_2236000# GND efet w=45500 l=9500
+ ad=0 pd=0 as=9.68e+08 ps=176000 
M5703 diff_94000_5193000# diff_5652000_2258000# diff_5652000_2258000# GND efet w=14000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M5704 diff_5956000_2221000# diff_5768000_2160000# diff_5618000_2171000# GND efet w=287500 l=10500
+ ad=1.946e+09 pd=282000 as=0 ps=0 
M5705 diff_94000_5193000# diff_5652000_2258000# diff_5617000_2218000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=1.048e+09 ps=234000 
M5706 diff_82000_3097000# diff_5760000_2171000# diff_5768000_2160000# GND efet w=488000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5707 diff_5617000_2218000# diff_5647000_2195000# diff_5625000_2183000# GND efet w=21000 l=13000
+ ad=0 pd=0 as=2.06e+09 ps=394000 
M5708 diff_94000_5193000# diff_5625000_2183000# diff_5625000_2183000# GND efet w=15000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M5709 diff_5618000_2171000# diff_5768000_2160000# diff_5956000_2165000# GND efet w=777000 l=10000
+ ad=0 pd=0 as=5.44098e+08 ps=1.464e+06 
M5710 diff_5625000_2183000# diff_5618000_2171000# diff_5619000_2114000# GND efet w=156500 l=11500
+ ad=0 pd=0 as=-1.60967e+08 ps=394000 
M5711 diff_5625000_2090000# diff_5618000_2101000# diff_5619000_2114000# GND efet w=157000 l=11000
+ ad=-1.99997e+09 pd=400000 as=0 ps=0 
M5712 diff_5768000_2029000# diff_5256000_3172000# diff_82000_3097000# GND efet w=487000 l=11000
+ ad=8.04065e+08 pd=1.634e+06 as=0 ps=0 
M5713 diff_5625000_2090000# diff_71000_4514000# diff_5617000_1924000# GND efet w=21000 l=13000
+ ad=0 pd=0 as=1.135e+09 ps=238000 
M5714 diff_94000_5193000# diff_5625000_2090000# diff_5625000_2090000# GND efet w=14000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M5715 diff_94000_5193000# diff_5768000_2029000# diff_5618000_2101000# GND efet w=780000 l=10000
+ ad=0 pd=0 as=3.63327e+08 ps=6.556e+06 
M5716 diff_94000_5193000# diff_5652000_2013000# diff_5617000_1924000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M5717 diff_5652000_2013000# diff_5631000_1935000# diff_82000_3097000# GND efet w=49000 l=10000
+ ad=1.154e+09 pd=210000 as=0 ps=0 
M5718 diff_94000_5193000# diff_5768000_2029000# diff_5618000_2101000# GND efet w=288000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5719 diff_5768000_2029000# diff_5696000_1748000# diff_82000_3097000# GND efet w=480000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5720 diff_94000_5193000# diff_5768000_2029000# diff_5618000_2101000# GND efet w=287500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5721 diff_94000_5193000# diff_5652000_2013000# diff_5652000_2013000# GND efet w=14000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M5722 diff_5652000_2013000# diff_71000_4514000# diff_82000_3097000# GND efet w=30000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5723 diff_5631000_1935000# diff_5617000_1924000# diff_82000_3097000# GND efet w=224500 l=10500
+ ad=-5.28967e+08 pd=734000 as=0 ps=0 
M5724 diff_5242000_1640000# diff_5242000_1640000# diff_5208000_1611000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5725 diff_5334000_1644000# diff_5224000_815000# diff_5242000_1640000# GND efet w=21000 l=13000
+ ad=1.47e+08 pd=56000 as=0 ps=0 
M5726 diff_5355000_1644000# diff_5270000_856000# diff_5334000_1644000# GND efet w=21000 l=14000
+ ad=3.56e+08 pd=98000 as=0 ps=0 
M5727 diff_5376000_1680000# diff_5376000_1680000# diff_5385000_1619000# GND efet w=15000 l=22000
+ ad=0 pd=0 as=1.28e+09 ps=150000 
M5728 diff_5465000_1671000# diff_5446000_801000# diff_5442000_1752000# GND efet w=89500 l=11500
+ ad=1.477e+09 pd=288000 as=9.07e+08 ps=210000 
M5729 diff_5028000_1618000# diff_5021000_1591000# diff_5021000_1591000# GND efet w=15000 l=27000
+ ad=0 pd=0 as=1.892e+09 ps=298000 
M5730 diff_5074000_1617000# diff_5068000_1594000# diff_5068000_1594000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=1.687e+09 ps=364000 
M5731 diff_5124000_1613000# diff_4931000_826000# diff_5074000_1617000# GND efet w=15000 l=10000
+ ad=4.70327e+07 pd=876000 as=0 ps=0 
M5732 diff_5158000_1629000# diff_5151000_1618000# diff_5124000_1613000# GND efet w=131500 l=11500
+ ad=1.671e+09 pd=354000 as=0 ps=0 
M5733 diff_4899000_1441000# diff_4893000_1432000# diff_4869000_1327000# GND efet w=61000 l=10000
+ ad=0 pd=0 as=-1.26197e+09 ps=472000 
M5734 diff_4866000_1360000# diff_4838000_2617000# diff_4831000_1268000# GND efet w=52000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5735 diff_4991000_1456000# diff_4982000_1450000# diff_4971000_1481000# GND efet w=35000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5736 diff_5024000_1356000# diff_4993000_2633000# diff_4991000_1456000# GND efet w=57000 l=11000
+ ad=-1.58197e+09 pd=420000 as=0 ps=0 
M5737 diff_5021000_1591000# diff_5037000_1510000# diff_5024000_1356000# GND efet w=46000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5738 diff_5124000_1613000# diff_5132000_1593000# diff_5111000_1386000# GND efet w=92000 l=13000
+ ad=0 pd=0 as=-1.67393e+09 ps=810000 
M5739 diff_5068000_1594000# diff_5068000_1533000# diff_5070000_1364000# GND efet w=67500 l=10500
+ ad=0 pd=0 as=1.874e+09 ps=374000 
M5740 diff_5111000_1386000# diff_4931000_826000# diff_5068000_1594000# GND efet w=67000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5741 diff_5208000_1611000# diff_5201000_1587000# diff_5201000_1587000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=1.627e+09 ps=348000 
M5742 diff_5242000_1606000# diff_5242000_1606000# diff_5208000_1611000# GND efet w=14000 l=23000
+ ad=-2.13797e+09 pd=494000 as=0 ps=0 
M5743 diff_5289000_1468000# diff_5278000_1526000# diff_5242000_1606000# GND efet w=79500 l=10500
+ ad=1.288e+09 pd=324000 as=0 ps=0 
M5744 diff_4831000_1268000# diff_4820000_1262000# diff_4809000_1268000# GND efet w=71000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5745 diff_4869000_1327000# diff_4838000_2617000# diff_4866000_1360000# GND efet w=60000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5746 diff_4701000_1242000# diff_4693000_1184000# diff_4693000_1184000# GND efet w=15000 l=27000
+ ad=0 pd=0 as=8.57e+08 ps=156000 
M5747 diff_4701000_1242000# diff_4726000_1105000# diff_4726000_1105000# GND efet w=15000 l=26000
+ ad=0 pd=0 as=1.652e+09 ps=298000 
M5748 diff_4423000_963000# diff_4373000_832000# diff_4413000_1027000# GND efet w=22000 l=11000
+ ad=1.139e+09 pd=226000 as=6.58e+08 ps=146000 
M5749 diff_4423000_963000# diff_4416000_951000# diff_4423000_931000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=4.4e+08 ps=84000 
M5750 diff_4477000_914000# diff_4477000_914000# diff_4481000_1020000# GND efet w=15000 l=106000
+ ad=7.97e+08 pd=154000 as=3.42e+08 ps=74000 
M5751 diff_4517000_900000# diff_4532000_955000# diff_4519000_996000# GND efet w=51000 l=10000
+ ad=1.774e+09 pd=314000 as=0 ps=0 
M5752 diff_4617000_986000# diff_4607000_1092000# diff_4574000_1196000# GND efet w=50000 l=10000
+ ad=-1.43297e+09 pd=388000 as=0 ps=0 
M5753 diff_4607000_1092000# diff_4624000_1155000# diff_4617000_986000# GND efet w=68000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5754 diff_4672000_1141000# diff_4547000_2724000# diff_4607000_1092000# GND efet w=23000 l=12000
+ ad=4.6e+08 pd=86000 as=0 ps=0 
M5755 diff_4706000_1141000# diff_4601000_2751000# diff_4672000_1141000# GND efet w=23000 l=14000
+ ad=4.37e+08 pd=84000 as=0 ps=0 
M5756 diff_4574000_899000# diff_4497000_2491000# diff_4563000_975000# GND efet w=23000 l=12000
+ ad=1.653e+09 pd=300000 as=3.91e+08 ps=80000 
M5757 diff_4617000_986000# diff_4607000_945000# diff_4574000_899000# GND efet w=51000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5758 diff_4607000_945000# diff_4624000_962000# diff_4617000_986000# GND efet w=69000 l=10000
+ ad=1.862e+09 pd=402000 as=0 ps=0 
M5759 diff_4706000_1096000# diff_4601000_2751000# diff_4675000_1096000# GND efet w=23000 l=14000
+ ad=5.04e+08 pd=146000 as=3.91e+08 ps=80000 
M5760 diff_4753000_1054000# diff_4706000_1096000# diff_4726000_1105000# GND efet w=51000 l=10000
+ ad=1.20803e+09 pd=820000 as=0 ps=0 
M5761 diff_4786000_1098000# diff_4739000_2640000# diff_4753000_1054000# GND efet w=150500 l=10500
+ ad=1.538e+09 pd=366000 as=0 ps=0 
M5762 diff_4809000_1139000# diff_4798000_1130000# diff_4786000_1098000# GND efet w=128000 l=11000
+ ad=2.102e+09 pd=410000 as=0 ps=0 
M5763 diff_4831000_1174000# diff_4820000_1150000# diff_4809000_1139000# GND efet w=71000 l=11000
+ ad=-1.95197e+09 pd=392000 as=0 ps=0 
M5764 diff_4899000_1441000# diff_4904000_1328000# diff_4869000_1327000# GND efet w=56000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5765 diff_4869000_1327000# diff_4869000_1327000# diff_4881000_1243000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=6.44e+08 ps=108000 
M5766 diff_4952000_1272000# diff_4904000_1328000# diff_4899000_1441000# GND efet w=137000 l=11000
+ ad=1.096e+09 pd=290000 as=0 ps=0 
M5767 diff_4971000_1272000# diff_4905000_2664000# diff_4952000_1272000# GND efet w=137000 l=11000
+ ad=1.647e+09 pd=350000 as=0 ps=0 
M5768 diff_4991000_1272000# diff_4982000_1267000# diff_4971000_1272000# GND efet w=33000 l=9000
+ ad=-2.10097e+09 pd=396000 as=0 ps=0 
M5769 diff_5334000_1601000# diff_5224000_815000# diff_5242000_1606000# GND efet w=22000 l=13000
+ ad=1.54e+08 pd=58000 as=0 ps=0 
M5770 diff_5355000_1601000# diff_5270000_856000# diff_5334000_1601000# GND efet w=22000 l=14000
+ ad=3.27e+08 pd=110000 as=0 ps=0 
M5771 diff_5124000_1613000# diff_5132000_1593000# diff_5111000_1386000# GND efet w=49500 l=12500
+ ad=0 pd=0 as=0 ps=0 
M5772 diff_5201000_1587000# diff_5158000_1629000# diff_5202000_1366000# GND efet w=79000 l=10000
+ ad=0 pd=0 as=1.908e+09 ps=360000 
M5773 diff_5124000_1262000# diff_5136000_1347000# diff_5111000_1386000# GND efet w=124000 l=11000
+ ad=7.40327e+07 pd=846000 as=0 ps=0 
M5774 diff_4991000_1272000# diff_4982000_1267000# diff_4971000_1272000# GND efet w=99000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5775 diff_5024000_1356000# diff_4993000_2633000# diff_4991000_1272000# GND efet w=56000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5776 diff_5021000_1275000# diff_5037000_1351000# diff_5024000_1356000# GND efet w=47000 l=8000
+ ad=1.804e+09 pd=296000 as=0 ps=0 
M5777 diff_5068000_1277000# diff_5068000_1339000# diff_5070000_1364000# GND efet w=65500 l=10500
+ ad=1.788e+09 pd=358000 as=0 ps=0 
M5778 diff_5111000_1386000# diff_4931000_826000# diff_5068000_1277000# GND efet w=66000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5779 diff_5124000_1613000# diff_5161000_1372000# diff_5124000_1262000# GND efet w=43000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5780 diff_4881000_1243000# diff_4870000_1181000# diff_4870000_1181000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=-1.45097e+09 ps=460000 
M5781 diff_4899000_1064000# diff_4904000_1167000# diff_4870000_1181000# GND efet w=53000 l=10000
+ ad=2.10033e+08 pd=808000 as=0 ps=0 
M5782 diff_4870000_1181000# diff_4838000_2617000# diff_4866000_1100000# GND efet w=65000 l=10000
+ ad=0 pd=0 as=-1.32397e+09 ps=456000 
M5783 diff_4831000_1174000# diff_4820000_1150000# diff_4809000_1139000# GND efet w=70500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5784 diff_4809000_1139000# diff_4798000_1130000# diff_4786000_1098000# GND efet w=13000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5785 diff_4866000_1100000# diff_4838000_2617000# diff_4831000_1174000# GND efet w=53000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5786 diff_4706000_1018000# diff_4601000_2751000# diff_4675000_1018000# GND efet w=22000 l=14000
+ ad=5.01e+08 pd=122000 as=3.74e+08 ps=78000 
M5787 diff_4517000_900000# diff_4517000_900000# diff_4530000_879000# GND efet w=15000 l=22000
+ ad=0 pd=0 as=4.17e+08 ps=84000 
M5788 diff_4405000_795000# diff_4393000_785000# diff_4373000_832000# GND efet w=84000 l=11000
+ ad=1.536e+09 pd=204000 as=0 ps=0 
M5789 diff_4416000_951000# diff_4393000_785000# diff_4405000_795000# GND efet w=72000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5790 diff_4672000_973000# diff_4547000_2724000# diff_4607000_945000# GND efet w=22000 l=12000
+ ad=4.4e+08 pd=84000 as=0 ps=0 
M5791 diff_4706000_973000# diff_4601000_2751000# diff_4672000_973000# GND efet w=22000 l=14000
+ ad=4.4e+08 pd=84000 as=0 ps=0 
M5792 diff_4753000_1054000# diff_4706000_1018000# diff_4726000_1005000# GND efet w=52000 l=10000
+ ad=0 pd=0 as=1.607e+09 ps=298000 
M5793 diff_4787000_982000# diff_4767000_995000# diff_4753000_1054000# GND efet w=28000 l=11000
+ ad=1.709e+09 pd=392000 as=0 ps=0 
M5794 diff_4809000_920000# diff_4763000_779000# diff_4787000_982000# GND efet w=12000 l=11000
+ ad=2.03e+09 pd=428000 as=0 ps=0 
M5795 diff_4809000_920000# diff_4763000_779000# diff_4787000_982000# GND efet w=139000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5796 diff_4831000_883000# diff_4794000_778000# diff_4809000_920000# GND efet w=69500 l=10500
+ ad=-1.96197e+09 pd=402000 as=0 ps=0 
M5797 diff_4787000_982000# diff_4767000_995000# diff_4753000_1054000# GND efet w=110000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5798 diff_4574000_899000# diff_4574000_899000# diff_4588000_876000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=1.009e+09 ps=148000 
M5799 diff_4607000_945000# diff_4607000_945000# diff_4588000_876000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M5800 diff_4585000_783000# diff_4573000_760000# diff_4497000_2491000# GND efet w=77000 l=12000
+ ad=1.282e+09 pd=188000 as=0 ps=0 
M5801 diff_4547000_2724000# diff_4573000_760000# diff_4585000_783000# GND efet w=77000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5802 diff_4601000_2751000# diff_4643000_761000# diff_4638000_782000# GND efet w=76500 l=11500
+ ad=0 pd=0 as=1.034e+09 ps=182000 
M5803 diff_4692000_926000# diff_4692000_926000# diff_4692000_844000# GND efet w=14000 l=27000
+ ad=7.83e+08 pd=156000 as=1.817e+09 ps=258000 
M5804 diff_4726000_1005000# diff_4726000_1005000# diff_4692000_844000# GND efet w=16000 l=27000
+ ad=0 pd=0 as=0 ps=0 
M5805 diff_4831000_883000# diff_4794000_778000# diff_4809000_920000# GND efet w=78000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5806 diff_4899000_1064000# diff_4893000_1075000# diff_4870000_1181000# GND efet w=60000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5807 diff_4951000_1103000# diff_4904000_1167000# diff_4899000_1064000# GND efet w=137000 l=10000
+ ad=1.233e+09 pd=292000 as=0 ps=0 
M5808 diff_4971000_1103000# diff_4905000_2664000# diff_4951000_1103000# GND efet w=137000 l=11000
+ ad=1.649e+09 pd=350000 as=0 ps=0 
M5809 diff_4991000_1078000# diff_4982000_1073000# diff_4971000_1103000# GND efet w=98000 l=9000
+ ad=-1.96297e+09 pd=398000 as=0 ps=0 
M5810 diff_5021000_1275000# diff_5021000_1275000# diff_5028000_1241000# GND efet w=15000 l=27000
+ ad=0 pd=0 as=6.83e+08 ps=110000 
M5811 diff_5068000_1277000# diff_5068000_1277000# diff_5074000_1239000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=1.496e+09 ps=178000 
M5812 diff_5124000_1262000# diff_5136000_1347000# diff_5111000_1386000# GND efet w=24000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5813 diff_5124000_1613000# diff_5161000_1372000# diff_5124000_1262000# GND efet w=73000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5814 diff_5243000_1366000# diff_5233000_1540000# diff_5201000_1587000# GND efet w=72500 l=9500
+ ad=1.73103e+09 pd=966000 as=0 ps=0 
M5815 diff_5242000_1606000# diff_5201000_1587000# diff_5243000_1366000# GND efet w=65500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5816 diff_5289000_1468000# diff_5278000_1526000# diff_5242000_1606000# GND efet w=34000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5817 diff_5289000_1468000# diff_5281000_1458000# diff_5243000_1366000# GND efet w=117500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5818 diff_5200000_1283000# diff_5124000_1613000# diff_5202000_1366000# GND efet w=79000 l=10000
+ ad=1.55e+09 pd=340000 as=0 ps=0 
M5819 diff_5243000_1366000# diff_5233000_1338000# diff_5200000_1283000# GND efet w=72500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5820 diff_5289000_1290000# diff_5281000_1426000# diff_5243000_1366000# GND efet w=122500 l=11500
+ ad=1.308e+09 pd=326000 as=0 ps=0 
M5821 diff_5242000_1263000# diff_5200000_1283000# diff_5243000_1366000# GND efet w=66500 l=10500
+ ad=-2.02497e+09 pd=498000 as=0 ps=0 
M5822 diff_5289000_1290000# diff_5278000_1281000# diff_5242000_1263000# GND efet w=36000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5823 diff_5200000_1283000# diff_5200000_1283000# diff_5208000_1234000# GND efet w=15000 l=24000
+ ad=0 pd=0 as=1.559e+09 ps=186000 
M5824 diff_5124000_1262000# diff_4931000_826000# diff_5074000_1239000# GND efet w=15000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5825 diff_5289000_1290000# diff_5278000_1281000# diff_5242000_1263000# GND efet w=76000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5826 diff_5376000_1575000# diff_5376000_1575000# diff_5385000_1619000# GND efet w=15000 l=24000
+ ad=1.754e+09 pd=326000 as=0 ps=0 
M5827 diff_5376000_1575000# diff_5355000_1601000# diff_5358000_1304000# GND efet w=192000 l=10000
+ ad=0 pd=0 as=-9.54935e+08 ps=1.278e+06 
M5828 diff_5330000_4061000# diff_5376000_1575000# diff_5358000_1304000# GND efet w=157500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5829 diff_5465000_1576000# diff_5446000_801000# diff_5442000_1495000# GND efet w=89500 l=12500
+ ad=1.375e+09 pd=286000 as=9.11e+08 ps=210000 
M5830 diff_94000_5193000# diff_5631000_1935000# diff_5631000_1935000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M5831 diff_5618000_2101000# diff_5768000_2029000# diff_94000_5193000# GND efet w=289000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5832 diff_82000_3097000# diff_82000_3097000# diff_5618000_2101000# GND efet w=94500 l=14500
+ ad=0 pd=0 as=0 ps=0 
M5833 diff_5768000_2029000# diff_5768000_2029000# diff_94000_5193000# GND efet w=46000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5834 diff_94000_5193000# diff_5696000_1748000# diff_5696000_1748000# GND efet w=35000 l=10000
+ ad=0 pd=0 as=1.55307e+09 ps=1.802e+06 
M5835 diff_82000_3097000# diff_5696000_1748000# diff_5618000_2101000# GND efet w=241000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5836 diff_5696000_1748000# diff_5256000_3172000# diff_82000_3097000# GND efet w=477000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5837 diff_5631000_1935000# diff_5555000_2636000# diff_5569000_1916000# GND efet w=89000 l=13000
+ ad=0 pd=0 as=1.872e+09 ps=328000 
M5838 diff_82000_3097000# diff_5649000_1748000# diff_5696000_1748000# GND efet w=515000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5839 diff_5569000_1916000# diff_5576000_2597000# diff_5649000_1748000# GND efet w=37000 l=14000
+ ad=0 pd=0 as=-1.31297e+09 ps=330000 
M5840 diff_82000_3097000# diff_5696000_1748000# diff_5618000_2101000# GND efet w=291000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5841 diff_82000_3097000# diff_5696000_1748000# diff_5618000_2101000# GND efet w=292000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M5842 diff_5618000_2101000# diff_5696000_1748000# diff_82000_3097000# GND efet w=803500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M5843 diff_5695000_1732000# diff_5649000_1677000# diff_82000_3097000# GND efet w=516000 l=11000
+ ad=1.26207e+09 pd=1.82e+06 as=0 ps=0 
M5844 diff_82000_3097000# diff_5695000_1732000# diff_5618000_1380000# GND efet w=805000 l=12000
+ ad=0 pd=0 as=-7.76673e+08 ps=6.478e+06 
M5845 diff_82000_3097000# diff_5751000_1599000# diff_5695000_1732000# GND efet w=477500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5846 diff_5649000_1677000# diff_5688000_1661000# diff_5564000_1651000# GND efet w=37000 l=13000
+ ad=-1.34997e+09 pd=304000 as=1.589e+09 ps=308000 
M5847 diff_5631000_1484000# diff_5633000_1635000# diff_5564000_1651000# GND efet w=89500 l=13500
+ ad=-2.78967e+08 pd=738000 as=0 ps=0 
M5848 diff_5488000_1611000# diff_5488000_1611000# diff_5497000_1490000# GND efet w=15000 l=23000
+ ad=1.663e+09 pd=302000 as=1.892e+09 ps=354000 
M5849 diff_5497000_1490000# diff_5472000_1599000# diff_5482000_1425000# GND efet w=128000 l=12000
+ ad=0 pd=0 as=1.802e+09 ps=262000 
M5850 diff_5376000_1304000# diff_5355000_1268000# diff_5358000_1304000# GND efet w=200500 l=10500
+ ad=1.795e+09 pd=304000 as=0 ps=0 
M5851 diff_5330000_4061000# diff_5376000_1304000# diff_5358000_1304000# GND efet w=155500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5852 diff_5242000_1263000# diff_5242000_1263000# diff_5208000_1234000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5853 diff_5335000_1268000# diff_5224000_815000# diff_5242000_1263000# GND efet w=21000 l=14000
+ ad=1.26e+08 pd=54000 as=0 ps=0 
M5854 diff_5355000_1268000# diff_5270000_856000# diff_5335000_1268000# GND efet w=21000 l=14000
+ ad=3.5e+08 pd=100000 as=0 ps=0 
M5855 diff_5376000_1304000# diff_5376000_1304000# diff_5385000_1242000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=1.298e+09 ps=152000 
M5856 diff_5465000_1294000# diff_5446000_801000# diff_5442000_1375000# GND efet w=89500 l=12500
+ ad=1.391e+09 pd=286000 as=9.07e+08 ps=210000 
M5857 diff_5028000_1241000# diff_5021000_1214000# diff_5021000_1214000# GND efet w=15000 l=27000
+ ad=0 pd=0 as=1.922e+09 ps=298000 
M5858 diff_5074000_1239000# diff_5068000_1217000# diff_5068000_1217000# GND efet w=15000 l=22000
+ ad=0 pd=0 as=1.702e+09 ps=366000 
M5859 diff_5124000_1236000# diff_4931000_826000# diff_5074000_1239000# GND efet w=15000 l=10000
+ ad=3.63033e+08 pd=946000 as=0 ps=0 
M5860 diff_5124000_1262000# diff_5151000_1240000# diff_5124000_1236000# GND efet w=131500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M5861 diff_4899000_1064000# diff_4893000_1055000# diff_4869000_938000# GND efet w=62000 l=10000
+ ad=0 pd=0 as=-8.76967e+08 ps=606000 
M5862 diff_4991000_1078000# diff_4982000_1073000# diff_4971000_1103000# GND efet w=35000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5863 diff_5024000_982000# diff_4993000_2633000# diff_4991000_1078000# GND efet w=57000 l=10000
+ ad=-1.59297e+09 pd=422000 as=0 ps=0 
M5864 diff_5021000_1214000# diff_5037000_1132000# diff_5024000_982000# GND efet w=47000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5865 diff_5124000_1236000# diff_5132000_1216000# diff_5111000_1009000# GND efet w=92000 l=13000
+ ad=0 pd=0 as=-1.64493e+09 ps=810000 
M5866 diff_5068000_1217000# diff_5068000_1155000# diff_5070000_986000# GND efet w=67500 l=10500
+ ad=0 pd=0 as=1.884e+09 ps=374000 
M5867 diff_5111000_1009000# diff_4931000_826000# diff_5068000_1217000# GND efet w=68000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5868 diff_5208000_1234000# diff_5201000_1209000# diff_5201000_1209000# GND efet w=15000 l=25000
+ ad=0 pd=0 as=1.599e+09 ps=346000 
M5869 diff_5242000_1228000# diff_5242000_1228000# diff_5208000_1234000# GND efet w=15000 l=23000
+ ad=-2.07897e+09 pd=498000 as=0 ps=0 
M5870 diff_5289000_1091000# diff_5278000_1149000# diff_5242000_1228000# GND efet w=79500 l=10500
+ ad=1.29e+09 pd=324000 as=0 ps=0 
M5871 diff_4866000_1100000# diff_4838000_2617000# diff_4869000_938000# GND efet w=60000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5872 diff_4869000_938000# diff_4869000_938000# diff_4852000_874000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=1.24e+09 ps=152000 
M5873 diff_4899000_1064000# diff_4904000_951000# diff_4869000_938000# GND efet w=54500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5874 diff_4706000_839000# diff_4706000_839000# diff_4692000_844000# GND efet w=15000 l=38000
+ ad=1.424e+09 pd=258000 as=0 ps=0 
M5875 diff_4949000_896000# diff_4904000_951000# diff_4899000_1064000# GND efet w=135000 l=11000
+ ad=1.652e+09 pd=348000 as=0 ps=0 
M5876 diff_4970000_889000# diff_4905000_2664000# diff_4949000_896000# GND efet w=66000 l=11000
+ ad=1.749e+09 pd=408000 as=0 ps=0 
M5877 diff_4991000_889000# diff_4980000_886000# diff_4970000_889000# GND efet w=34000 l=9000
+ ad=-1.47967e+08 pd=702000 as=0 ps=0 
M5878 diff_5335000_1224000# diff_5224000_815000# diff_5242000_1228000# GND efet w=23000 l=14000
+ ad=1.38e+08 pd=58000 as=0 ps=0 
M5879 diff_5355000_1224000# diff_5270000_856000# diff_5335000_1224000# GND efet w=23000 l=14000
+ ad=3.46e+08 pd=110000 as=0 ps=0 
M5880 diff_5124000_1236000# diff_5132000_1216000# diff_5111000_1009000# GND efet w=49000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5881 diff_5201000_1209000# diff_5124000_1262000# diff_5202000_989000# GND efet w=79000 l=10000
+ ad=0 pd=0 as=1.897e+09 ps=360000 
M5882 diff_5124000_885000# diff_5136000_970000# diff_5111000_1009000# GND efet w=124000 l=11000
+ ad=-1.66897e+09 pd=542000 as=0 ps=0 
M5883 diff_4852000_874000# diff_4837000_813000# diff_4837000_813000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=1.056e+09 ps=210000 
M5884 diff_4970000_889000# diff_4905000_2664000# diff_4949000_896000# GND efet w=67000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5885 diff_4991000_889000# diff_4980000_886000# diff_4970000_889000# GND efet w=115500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5886 diff_5024000_982000# diff_4993000_2633000# diff_4991000_889000# GND efet w=52000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5887 diff_4991000_889000# diff_5037000_973000# diff_5024000_982000# GND efet w=47000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5888 diff_5068000_900000# diff_5068000_962000# diff_5070000_986000# GND efet w=66500 l=10500
+ ad=1.817e+09 pd=360000 as=0 ps=0 
M5889 diff_5111000_1009000# diff_4931000_826000# diff_5068000_900000# GND efet w=67000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5890 diff_5124000_1236000# diff_5161000_995000# diff_5124000_885000# GND efet w=43000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5891 diff_4991000_889000# diff_4991000_889000# diff_5029000_876000# GND efet w=14000 l=27000
+ ad=0 pd=0 as=4.36e+08 ps=86000 
M5892 diff_5068000_900000# diff_5068000_900000# diff_5074000_876000# GND efet w=14000 l=21000
+ ad=0 pd=0 as=9.06e+08 ps=136000 
M5893 diff_5124000_885000# diff_5136000_970000# diff_5111000_1009000# GND efet w=23000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5894 diff_5124000_1236000# diff_5161000_995000# diff_5124000_885000# GND efet w=73000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5895 diff_5243000_989000# diff_5233000_1162000# diff_5201000_1209000# GND efet w=73500 l=9500
+ ad=1.71403e+09 pd=966000 as=0 ps=0 
M5896 diff_5242000_1228000# diff_5201000_1209000# diff_5243000_989000# GND efet w=65500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5897 diff_5289000_1091000# diff_5278000_1149000# diff_5242000_1228000# GND efet w=35000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5898 diff_5289000_1091000# diff_5281000_1081000# diff_5243000_989000# GND efet w=117500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5899 diff_5200000_906000# diff_5124000_1236000# diff_5202000_989000# GND efet w=79000 l=10000
+ ad=1.557e+09 pd=340000 as=0 ps=0 
M5900 diff_5243000_989000# diff_5233000_961000# diff_5200000_906000# GND efet w=72500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5901 diff_5243000_989000# diff_5281000_1049000# diff_5289000_913000# GND efet w=121000 l=11000
+ ad=0 pd=0 as=1.298e+09 ps=326000 
M5902 diff_5242000_886000# diff_5200000_906000# diff_5243000_989000# GND efet w=66500 l=10500
+ ad=-2.02297e+09 pd=498000 as=0 ps=0 
M5903 diff_5289000_913000# diff_5278000_904000# diff_5242000_886000# GND efet w=36000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5904 diff_5124000_885000# diff_4931000_826000# diff_5074000_876000# GND efet w=15000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5905 diff_5200000_906000# diff_5200000_906000# diff_5208000_877000# GND efet w=15000 l=25000
+ ad=0 pd=0 as=8.75e+08 ps=132000 
M5906 diff_5289000_913000# diff_5278000_904000# diff_5242000_886000# GND efet w=76000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5907 diff_5385000_1242000# diff_5376000_1197000# diff_5376000_1197000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=1.791e+09 ps=328000 
M5908 diff_5376000_1197000# diff_5355000_1224000# diff_5358000_927000# GND efet w=195000 l=10000
+ ad=0 pd=0 as=-8.63935e+08 ps=1.278e+06 
M5909 diff_5330000_4061000# diff_5376000_1197000# diff_5358000_927000# GND efet w=157500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5910 diff_5465000_1199000# diff_5446000_801000# diff_5442000_1118000# GND efet w=89500 l=12500
+ ad=1.37e+09 pd=286000 as=9.12e+08 ps=210000 
M5911 diff_5376000_927000# diff_5355000_891000# diff_5358000_927000# GND efet w=199500 l=10500
+ ad=1.799e+09 pd=304000 as=0 ps=0 
M5912 diff_5330000_4061000# diff_5376000_927000# diff_5358000_927000# GND efet w=156500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5913 diff_5242000_886000# diff_5242000_886000# diff_5208000_877000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5914 diff_5334000_891000# diff_5224000_815000# diff_5242000_886000# GND efet w=21000 l=13000
+ ad=1.68e+08 pd=58000 as=0 ps=0 
M5915 diff_5355000_891000# diff_5270000_856000# diff_5334000_891000# GND efet w=21000 l=13000
+ ad=3.42e+08 pd=98000 as=0 ps=0 
M5916 diff_5376000_927000# diff_5376000_927000# diff_5384000_877000# GND efet w=15000 l=16000
+ ad=0 pd=0 as=1.483e+09 ps=176000 
M5917 diff_5465000_917000# diff_5446000_801000# diff_5442000_999000# GND efet w=90500 l=12500
+ ad=1.412e+09 pd=288000 as=9.15e+08 ps=212000 
M5918 diff_5631000_1484000# diff_5617000_1426000# diff_5619000_1567000# GND efet w=222500 l=10500
+ ad=0 pd=0 as=2.086e+09 ps=286000 
M5919 diff_82000_3097000# diff_5695000_1732000# diff_5618000_1380000# GND efet w=291500 l=12500
+ ad=0 pd=0 as=0 ps=0 
M5920 diff_82000_3097000# diff_5695000_1732000# diff_5618000_1380000# GND efet w=290500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M5921 diff_5618000_1380000# diff_5695000_1732000# diff_82000_3097000# GND efet w=240500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M5922 diff_5695000_1732000# diff_5695000_1732000# diff_5695000_1732000# GND efet w=3000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5923 diff_5695000_1732000# diff_5695000_1732000# diff_94000_5193000# GND efet w=38000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5924 diff_94000_5193000# diff_5631000_1484000# diff_5631000_1484000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M5925 diff_5654000_1521000# diff_5645000_1511000# diff_5652000_1465000# GND efet w=30000 l=11000
+ ad=5.39e+08 pd=96000 as=1.143e+09 ps=210000 
M5926 diff_94000_5193000# diff_5768000_1367000# diff_5768000_1367000# GND efet w=46000 l=10000
+ ad=0 pd=0 as=5.36065e+08 ps=1.636e+06 
M5927 diff_82000_3097000# diff_5695000_1732000# diff_5768000_1367000# GND efet w=480000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5928 diff_5618000_1380000# diff_5768000_1367000# diff_94000_5193000# GND efet w=287000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5929 diff_5956000_1477000# diff_5768000_1367000# diff_5618000_1380000# GND efet w=287500 l=10500
+ ad=2.07e+09 pd=284000 as=0 ps=0 
M5930 diff_5652000_1465000# diff_5631000_1484000# diff_5631000_1443000# GND efet w=45500 l=9500
+ ad=0 pd=0 as=9.64e+08 ps=174000 
M5931 diff_94000_5193000# diff_5652000_1465000# diff_5652000_1465000# GND efet w=13000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M5932 diff_5956000_1428000# diff_5768000_1367000# diff_5618000_1380000# GND efet w=288000 l=10000
+ ad=1.946e+09 pd=282000 as=0 ps=0 
M5933 diff_94000_5193000# diff_5652000_1465000# diff_5617000_1426000# GND efet w=16000 l=14000
+ ad=0 pd=0 as=1.133e+09 ps=236000 
M5934 diff_82000_3097000# diff_5760000_1378000# diff_5768000_1367000# GND efet w=487500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5935 diff_5617000_1426000# diff_5647000_1402000# diff_5625000_1391000# GND efet w=21000 l=12000
+ ad=0 pd=0 as=1.957e+09 ps=396000 
M5936 diff_94000_5193000# diff_5625000_1391000# diff_5625000_1391000# GND efet w=14000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M5937 diff_5618000_1380000# diff_5768000_1367000# diff_5956000_1373000# GND efet w=788000 l=10000
+ ad=0 pd=0 as=2.13807e+09 ps=1.454e+06 
M5938 diff_5625000_1391000# diff_5618000_1380000# diff_5619000_1321000# GND efet w=157000 l=11000
+ ad=0 pd=0 as=-1.22967e+08 ps=398000 
M5939 diff_6411000_1274000# diff_6411000_1274000# diff_5618000_1380000# GND efet w=99000 l=14000
+ ad=-2.07897e+09 pd=378000 as=0 ps=0 
M5940 diff_5625000_1298000# diff_5618000_1308000# diff_5619000_1321000# GND efet w=157500 l=11500
+ ad=-2.00797e+09 pd=400000 as=0 ps=0 
M5941 diff_5768000_1237000# diff_5256000_3172000# diff_82000_3097000# GND efet w=487000 l=11000
+ ad=6.31065e+08 pd=1.632e+06 as=0 ps=0 
M5942 diff_4772000_785000# diff_4763000_779000# diff_4706000_839000# GND efet w=44000 l=9000
+ ad=9.68e+08 pd=132000 as=0 ps=0 
M5943 diff_4775000_737000# diff_4794000_778000# diff_4772000_785000# GND efet w=44000 l=10000
+ ad=1.268e+09 pd=262000 as=0 ps=0 
M5944 diff_4890000_783000# diff_4869000_938000# diff_4837000_813000# GND efet w=45000 l=11000
+ ad=9e+08 pd=130000 as=0 ps=0 
M5945 diff_4962000_774000# diff_4950000_763000# diff_4931000_826000# GND efet w=73000 l=12000
+ ad=1.109e+09 pd=186000 as=0 ps=0 
M5946 diff_5008000_837000# diff_4977000_818000# diff_5008000_804000# GND efet w=139500 l=9500
+ ad=1.598e+09 pd=338000 as=1.336e+09 ps=260000 
M5947 diff_4775000_737000# diff_4775000_737000# diff_4751000_699000# GND efet w=14000 l=38000
+ ad=0 pd=0 as=1.152e+09 ps=176000 
M5948 diff_3395000_613000# diff_3395000_613000# diff_3395000_699000# GND efet w=18000 l=10000
+ ad=-5.05967e+08 pd=644000 as=4.21e+08 ps=84000 
M5949 diff_3416000_637000# diff_2759000_1455000# diff_3395000_613000# GND efet w=233000 l=10000
+ ad=-1.63897e+09 pd=316000 as=0 ps=0 
M5950 diff_3331000_584000# diff_3331000_584000# diff_3482000_692000# GND efet w=52500 l=9500
+ ad=-5.65902e+08 pd=2.026e+06 as=4.6e+08 ps=86000 
M5951 diff_3489000_578000# diff_3481000_567000# diff_3331000_584000# GND efet w=485500 l=10500
+ ad=-1.45997e+09 pd=500000 as=0 ps=0 
M5952 diff_3357000_541000# diff_3257000_122000# diff_3257000_122000# GND efet w=36000 l=10000
+ ad=6.84e+08 pd=110000 as=0 ps=0 
M5953 diff_3481000_567000# diff_3472000_667000# diff_3395000_613000# GND efet w=37000 l=13000
+ ad=7.98e+08 pd=186000 as=0 ps=0 
M5954 diff_3579000_635000# diff_3568000_625000# diff_3331000_584000# GND efet w=439000 l=10000
+ ad=-1.09397e+09 pd=452000 as=0 ps=0 
M5955 diff_3257000_122000# diff_3331000_584000# diff_3391000_545000# GND efet w=46000 l=11000
+ ad=0 pd=0 as=1.984e+09 ps=304000 
M5956 diff_3754000_578000# diff_3745000_567000# diff_3672000_544000# GND efet w=491500 l=10500
+ ad=-1.52597e+09 pd=508000 as=-6.76902e+08 ps=2.034e+06 
M5957 diff_3697000_661000# diff_3687000_625000# diff_3672000_544000# GND efet w=439000 l=10000
+ ad=-1.17297e+09 pd=456000 as=0 ps=0 
M5958 diff_3829000_692000# diff_3672000_544000# diff_3672000_544000# GND efet w=54500 l=9500
+ ad=5e+08 pd=90000 as=0 ps=0 
M5959 diff_3874000_651000# diff_3256000_1245000# diff_3853000_624000# GND efet w=233500 l=10500
+ ad=-1.79797e+09 pd=316000 as=-3.48967e+08 ps=648000 
M5960 diff_3921000_699000# diff_3853000_624000# diff_3853000_624000# GND efet w=18000 l=10000
+ ad=4.57e+08 pd=88000 as=0 ps=0 
M5961 diff_3853000_624000# diff_3840000_619000# diff_3745000_567000# GND efet w=37000 l=13000
+ ad=0 pd=0 as=7.08e+08 ps=180000 
M5962 diff_3971000_593000# diff_3672000_544000# diff_3898000_566000# GND efet w=275000 l=10000
+ ad=-2.05997e+09 pd=280000 as=1.95407e+09 ps=1.506e+06 
M5963 diff_4015000_715000# diff_4005000_705000# diff_3898000_566000# GND efet w=303500 l=10500
+ ad=-8.55967e+08 pd=436000 as=0 ps=0 
M5964 diff_3898000_566000# diff_3672000_544000# diff_3898000_545000# GND efet w=47000 l=11000
+ ad=0 pd=0 as=1.987e+09 ps=306000 
M5965 diff_3266000_457000# diff_3257000_122000# diff_2875000_456000# GND efet w=185000 l=10000
+ ad=-1.87371e+09 pd=4.538e+06 as=-1.22754e+09 ps=2.73e+06 
M5966 diff_3338000_491000# diff_3257000_122000# diff_3266000_457000# GND efet w=186000 l=10000
+ ad=1.229e+09 pd=188000 as=0 ps=0 
M5967 diff_1628000_457000# diff_1693000_584000# diff_1873000_101000# GND efet w=271000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5968 diff_2050000_195000# diff_2034000_544000# diff_1873000_101000# GND efet w=272000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5969 diff_2050000_195000# diff_2260000_566000# diff_2295000_101000# GND efet w=282000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5970 diff_2459000_132000# diff_2449000_122000# diff_2295000_101000# GND efet w=283000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5971 diff_2459000_132000# diff_2523000_584000# diff_2705000_101000# GND efet w=271000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5972 diff_3266000_457000# diff_3257000_122000# diff_2875000_456000# GND efet w=648500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5973 diff_3391000_545000# diff_3257000_122000# diff_3266000_457000# GND efet w=193000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5974 diff_3447000_491000# diff_3331000_584000# diff_3266000_457000# GND efet w=210000 l=10000
+ ad=1.337e+09 pd=208000 as=0 ps=0 
M5975 diff_3500000_492000# diff_3331000_584000# diff_3266000_457000# GND efet w=205500 l=10500
+ ad=1.36e+09 pd=204000 as=0 ps=0 
M5976 diff_3554000_491000# diff_3331000_584000# diff_3266000_457000# GND efet w=205500 l=10500
+ ad=1.328e+09 pd=204000 as=0 ps=0 
M5977 diff_3511000_102000# diff_3331000_584000# diff_3266000_457000# GND efet w=192000 l=10000
+ ad=-1.54777e+09 pd=2.938e+06 as=0 ps=0 
M5978 diff_3688000_195000# diff_3672000_544000# diff_3511000_102000# GND efet w=193000 l=10000
+ ad=-1.92171e+09 pd=4.536e+06 as=0 ps=0 
M5979 diff_3511000_102000# diff_3331000_584000# diff_3266000_457000# GND efet w=653000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5980 diff_3761000_491000# diff_3672000_544000# diff_3688000_195000# GND efet w=205500 l=10500
+ ad=1.36e+09 pd=204000 as=0 ps=0 
M5981 diff_3688000_195000# diff_3672000_544000# diff_3511000_102000# GND efet w=653000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5982 diff_3266000_457000# diff_3257000_122000# diff_2875000_456000# GND efet w=282000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5983 diff_3814000_491000# diff_3672000_544000# diff_3688000_195000# GND efet w=205500 l=10500
+ ad=1.36e+09 pd=204000 as=0 ps=0 
M5984 diff_3866000_491000# diff_3672000_544000# diff_3688000_195000# GND efet w=210000 l=10000
+ ad=1.369e+09 pd=208000 as=0 ps=0 
M5985 diff_3898000_566000# diff_3898000_566000# diff_3959000_541000# GND efet w=36000 l=10000
+ ad=0 pd=0 as=6.48e+08 ps=108000 
M5986 diff_3898000_566000# diff_4005000_705000# diff_4015000_715000# GND efet w=58000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5987 diff_3898000_545000# diff_3898000_566000# diff_3688000_195000# GND efet w=193000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5988 diff_4110000_566000# diff_4100000_556000# diff_4087000_122000# GND efet w=58000 l=10000
+ ad=-9.07967e+08 pd=440000 as=1.89807e+09 ps=1.498e+06 
M5989 diff_4110000_566000# diff_4100000_556000# diff_4087000_122000# GND efet w=302000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5990 diff_4172000_589000# diff_4161000_584000# diff_4087000_122000# GND efet w=274000 l=11000
+ ad=-2.14097e+09 pd=278000 as=0 ps=0 
M5991 diff_4226000_612000# diff_4226000_612000# diff_4225000_699000# GND efet w=18000 l=10000
+ ad=-5.89967e+08 pd=644000 as=4.42e+08 ps=86000 
M5992 diff_4246000_637000# diff_3907000_737000# diff_4226000_612000# GND efet w=234000 l=10000
+ ad=-1.66197e+09 pd=316000 as=0 ps=0 
M5993 diff_4161000_584000# diff_4161000_584000# diff_4312000_692000# GND efet w=53000 l=10000
+ ad=-7.29902e+08 pd=2.03e+06 as=4.6e+08 ps=86000 
M5994 diff_4319000_578000# diff_4311000_567000# diff_4161000_584000# GND efet w=485500 l=10500
+ ad=-1.58297e+09 pd=500000 as=0 ps=0 
M5995 diff_4187000_542000# diff_4087000_122000# diff_4087000_122000# GND efet w=36000 l=10000
+ ad=7.2e+08 pd=112000 as=0 ps=0 
M5996 diff_4311000_567000# diff_4302000_667000# diff_4226000_612000# GND efet w=37000 l=14000
+ ad=7.36e+08 pd=182000 as=0 ps=0 
M5997 diff_4409000_635000# diff_4398000_625000# diff_4161000_584000# GND efet w=441000 l=10000
+ ad=-9.89967e+08 pd=456000 as=0 ps=0 
M5998 diff_4087000_122000# diff_4161000_584000# diff_4221000_545000# GND efet w=46000 l=11000
+ ad=0 pd=0 as=1.955e+09 ps=306000 
M5999 diff_3974000_491000# diff_3898000_566000# diff_3688000_195000# GND efet w=186500 l=10500
+ ad=1.228e+09 pd=188000 as=0 ps=0 
M6000 diff_3932000_101000# diff_3898000_566000# diff_3688000_195000# GND efet w=183000 l=10000
+ ad=1.68716e+09 pd=2.896e+06 as=0 ps=0 
M6001 diff_4097000_195000# diff_4087000_122000# diff_3932000_101000# GND efet w=184000 l=10000
+ ad=-1.64071e+09 pd=4.524e+06 as=0 ps=0 
M6002 diff_3932000_101000# diff_3898000_566000# diff_3688000_195000# GND efet w=646500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M6003 diff_4168000_491000# diff_4087000_122000# diff_4097000_195000# GND efet w=183500 l=10500
+ ad=1.171e+09 pd=188000 as=0 ps=0 
M6004 diff_4585000_578000# diff_4575000_567000# diff_4502000_545000# GND efet w=489500 l=10500
+ ad=-1.56397e+09 pd=504000 as=-7.57902e+08 ps=2.034e+06 
M6005 diff_4527000_661000# diff_4517000_655000# diff_4502000_545000# GND efet w=441000 l=10000
+ ad=-1.02997e+09 pd=458000 as=0 ps=0 
M6006 diff_4660000_692000# diff_4502000_545000# diff_4502000_545000# GND efet w=54000 l=10000
+ ad=4.8e+08 pd=88000 as=0 ps=0 
M6007 diff_4704000_651000# diff_4302000_737000# diff_4684000_624000# GND efet w=232000 l=10000
+ ad=-1.78397e+09 pd=316000 as=-3.43967e+08 ps=646000 
M6008 diff_4751000_699000# diff_4684000_624000# diff_4684000_624000# GND efet w=18000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6009 diff_4802000_593000# diff_4502000_545000# diff_4728000_566000# GND efet w=275000 l=11000
+ ad=-2.14697e+09 pd=278000 as=2.04507e+09 ps=1.506e+06 
M6010 diff_4684000_624000# diff_4670000_619000# diff_4575000_567000# GND efet w=37000 l=14000
+ ad=0 pd=0 as=7.28e+08 ps=180000 
M6011 diff_4846000_715000# diff_4836000_704000# diff_4728000_566000# GND efet w=302000 l=10000
+ ad=-9.12967e+08 pd=434000 as=0 ps=0 
M6012 diff_4728000_566000# diff_4502000_545000# diff_4728000_545000# GND efet w=47000 l=11000
+ ad=0 pd=0 as=1.996e+09 ps=306000 
M6013 diff_4097000_195000# diff_4087000_122000# diff_3932000_101000# GND efet w=650500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M6014 diff_4221000_545000# diff_4087000_122000# diff_4097000_195000# GND efet w=190500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M6015 diff_4278000_490000# diff_4161000_584000# diff_4097000_195000# GND efet w=208500 l=10500
+ ad=1.327e+09 pd=206000 as=0 ps=0 
M6016 diff_4331000_491000# diff_4161000_584000# diff_4097000_195000# GND efet w=205000 l=10000
+ ad=1.332e+09 pd=204000 as=0 ps=0 
M6017 diff_4384000_491000# diff_4161000_584000# diff_4097000_195000# GND efet w=205500 l=10500
+ ad=1.364e+09 pd=204000 as=0 ps=0 
M6018 diff_4342000_102000# diff_4161000_584000# diff_4097000_195000# GND efet w=190000 l=10000
+ ad=-1.99077e+09 pd=2.926e+06 as=0 ps=0 
M6019 diff_4519000_195000# diff_4502000_545000# diff_4342000_102000# GND efet w=192000 l=10000
+ ad=-1.82371e+09 pd=4.542e+06 as=0 ps=0 
M6020 diff_4342000_102000# diff_4161000_584000# diff_4097000_195000# GND efet w=648000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M6021 diff_4591000_491000# diff_4502000_545000# diff_4519000_195000# GND efet w=207500 l=10500
+ ad=1.384e+09 pd=206000 as=0 ps=0 
M6022 diff_3266000_457000# diff_3331000_584000# diff_3511000_102000# GND efet w=272000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6023 diff_3688000_195000# diff_3672000_544000# diff_3511000_102000# GND efet w=272000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6024 diff_3688000_195000# diff_3898000_566000# diff_3932000_101000# GND efet w=281500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M6025 diff_4097000_195000# diff_4087000_122000# diff_3932000_101000# GND efet w=283000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6026 diff_4519000_195000# diff_4502000_545000# diff_4342000_102000# GND efet w=650000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M6027 diff_4644000_491000# diff_4502000_545000# diff_4519000_195000# GND efet w=207000 l=10000
+ ad=1.352e+09 pd=206000 as=0 ps=0 
M6028 diff_4697000_490000# diff_4502000_545000# diff_4519000_195000# GND efet w=212000 l=10000
+ ad=1.388e+09 pd=210000 as=0 ps=0 
M6029 diff_4728000_566000# diff_4728000_566000# diff_4790000_541000# GND efet w=37000 l=10000
+ ad=0 pd=0 as=6.29e+08 ps=108000 
M6030 diff_4728000_566000# diff_4836000_704000# diff_4846000_715000# GND efet w=58000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M6031 diff_5055000_793000# diff_4775000_737000# diff_5008000_837000# GND efet w=132500 l=10500
+ ad=1.978e+09 pd=368000 as=0 ps=0 
M6032 diff_5079000_824000# diff_5069000_814000# diff_5055000_793000# GND efet w=138500 l=10500
+ ad=1.369e+09 pd=256000 as=0 ps=0 
M6033 diff_5119000_786000# diff_5119000_786000# diff_5097000_842000# GND efet w=20000 l=9000
+ ad=-1.76967e+08 pd=690000 as=6.73e+08 ps=140000 
M6034 diff_5153000_743000# diff_5124000_885000# diff_5119000_786000# GND efet w=258500 l=10500
+ ad=1.914e+09 pd=254000 as=0 ps=0 
M6035 diff_5330000_4061000# diff_5330000_4061000# diff_5384000_877000# GND efet w=15000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M6036 diff_5270000_856000# diff_5243000_837000# diff_5270000_827000# GND efet w=73000 l=13000
+ ad=9.33e+08 pd=242000 as=2.033e+09 ps=206000 
M6037 diff_5625000_1298000# diff_71000_4514000# diff_5617000_1132000# GND efet w=21000 l=13000
+ ad=0 pd=0 as=1.154e+09 ps=238000 
M6038 diff_94000_5193000# diff_5625000_1298000# diff_5625000_1298000# GND efet w=15000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M6039 diff_94000_5193000# diff_5768000_1237000# diff_5618000_1308000# GND efet w=781000 l=10000
+ ad=0 pd=0 as=6.68327e+08 ps=6.646e+06 
M6040 diff_94000_5193000# diff_5652000_1221000# diff_5617000_1132000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M6041 diff_5652000_1221000# diff_5631000_1143000# diff_82000_3097000# GND efet w=49000 l=10000
+ ad=1.153e+09 pd=210000 as=0 ps=0 
M6042 diff_94000_5193000# diff_5768000_1237000# diff_5618000_1308000# GND efet w=288000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6043 diff_5768000_1237000# diff_5696000_956000# diff_82000_3097000# GND efet w=480000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6044 diff_94000_5193000# diff_5768000_1237000# diff_5618000_1308000# GND efet w=287500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M6045 diff_94000_5193000# diff_5652000_1221000# diff_5652000_1221000# GND efet w=14000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M6046 diff_5652000_1221000# diff_71000_4514000# diff_82000_3097000# GND efet w=30000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M6047 diff_5631000_1143000# diff_5617000_1132000# diff_82000_3097000# GND efet w=225500 l=10500
+ ad=-5.36967e+08 pd=734000 as=0 ps=0 
M6048 diff_94000_5193000# diff_5631000_1143000# diff_5631000_1143000# GND efet w=16000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M6049 diff_5618000_1308000# diff_5768000_1237000# diff_94000_5193000# GND efet w=289000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6050 diff_6411000_1274000# diff_6411000_1274000# diff_5618000_1308000# GND efet w=95500 l=14500
+ ad=0 pd=0 as=0 ps=0 
M6051 diff_5768000_1237000# diff_5768000_1237000# diff_94000_5193000# GND efet w=46000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6052 diff_94000_5193000# diff_5696000_956000# diff_5696000_956000# GND efet w=35000 l=10000
+ ad=0 pd=0 as=1.43807e+09 ps=1.798e+06 
M6053 diff_82000_3097000# diff_5696000_956000# diff_5618000_1308000# GND efet w=241000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M6054 diff_5696000_956000# diff_5256000_3172000# diff_82000_3097000# GND efet w=477000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6055 diff_5631000_1143000# diff_5555000_2636000# diff_5556000_1148000# GND efet w=89000 l=13000
+ ad=0 pd=0 as=-3.36967e+08 ps=632000 
M6056 diff_82000_3097000# diff_5650000_956000# diff_5696000_956000# GND efet w=515000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M6057 diff_5556000_1148000# diff_5576000_2597000# diff_5650000_956000# GND efet w=37000 l=14000
+ ad=0 pd=0 as=-1.43297e+09 ps=328000 
M6058 diff_82000_3097000# diff_5696000_956000# diff_5618000_1308000# GND efet w=291000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M6059 diff_82000_3097000# diff_5696000_956000# diff_5618000_1308000# GND efet w=292000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M6060 diff_5618000_1308000# diff_5696000_956000# diff_82000_3097000# GND efet w=802500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M6061 diff_5695000_940000# diff_5650000_887000# diff_82000_3097000# GND efet w=516000 l=11000
+ ad=1.06107e+09 pd=1.814e+06 as=0 ps=0 
M6062 diff_82000_3097000# diff_5695000_940000# diff_5599000_574000# GND efet w=806000 l=12000
+ ad=0 pd=0 as=-5.2664e+08 ps=7.096e+06 
M6063 diff_82000_3097000# diff_5751000_807000# diff_5695000_940000# GND efet w=477500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M6064 diff_5055000_793000# diff_5080000_704000# diff_5080000_704000# GND efet w=14000 l=13000
+ ad=0 pd=0 as=1.175e+09 ps=204000 
M6065 diff_5255000_745000# diff_5124000_1236000# diff_5069000_814000# GND efet w=57000 l=10000
+ ad=-1.75697e+09 pd=438000 as=9.55e+08 ps=214000 
M6066 diff_5069000_814000# diff_5069000_814000# diff_5213000_671000# GND efet w=12000 l=38000
+ ad=0 pd=0 as=1.234e+09 ps=186000 
M6067 diff_5388000_801000# diff_5323000_632000# diff_5370000_762000# GND efet w=174500 l=10500
+ ad=-5.88967e+08 pd=620000 as=1.785e+09 ps=364000 
M6068 diff_5650000_887000# diff_5483000_731000# diff_5550000_857000# GND efet w=37000 l=13000
+ ad=-1.56997e+09 pd=300000 as=-2.12797e+09 ps=416000 
M6069 diff_5417000_723000# diff_5342000_794000# diff_5388000_801000# GND efet w=166000 l=11000
+ ad=-2.10497e+09 pd=366000 as=0 ps=0 
M6070 diff_5323000_632000# diff_5124000_1236000# diff_5255000_745000# GND efet w=132500 l=10500
+ ad=-2.02497e+09 pd=402000 as=0 ps=0 
M6071 diff_5255000_745000# diff_5242000_710000# diff_5276000_709000# GND efet w=127500 l=10500
+ ad=0 pd=0 as=1.162e+09 ps=234000 
M6072 diff_4920000_663000# diff_4953000_638000# diff_4943000_579000# GND efet w=48000 l=13000
+ ad=-1.23097e+09 pd=436000 as=-2.08797e+09 ps=230000 
M6073 diff_5027000_596000# diff_5010000_575000# diff_4920000_663000# GND efet w=86000 l=13000
+ ad=-3.51967e+08 pd=574000 as=0 ps=0 
M6074 diff_5080000_704000# diff_5027000_596000# diff_5027000_596000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M6075 diff_5114000_586000# diff_5114000_586000# diff_5080000_704000# GND efet w=16000 l=38000
+ ad=-1.86697e+09 pd=480000 as=0 ps=0 
M6076 diff_4966000_476000# diff_5038000_606000# diff_5027000_596000# GND efet w=230000 l=10000
+ ad=1.64807e+09 pd=1.554e+06 as=0 ps=0 
M6077 diff_5114000_586000# diff_5027000_596000# diff_5114000_610000# GND efet w=36000 l=11000
+ ad=0 pd=0 as=6.24e+08 ps=112000 
M6078 diff_5114000_610000# diff_5105000_599000# diff_5114000_586000# GND efet w=28000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M6079 diff_5213000_671000# diff_5114000_586000# diff_5038000_606000# GND efet w=14000 l=13000
+ ad=0 pd=0 as=1.144e+09 ps=274000 
M6080 diff_5213000_671000# diff_5214000_614000# diff_5214000_614000# GND efet w=14000 l=13000
+ ad=0 pd=0 as=-2.10097e+09 ps=434000 
M6081 diff_5214000_614000# diff_5201000_599000# diff_5038000_606000# GND efet w=21000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M6082 diff_5446000_801000# diff_5430000_735000# diff_5417000_723000# GND efet w=75500 l=11500
+ ad=9.68e+08 pd=208000 as=0 ps=0 
M6083 diff_5550000_857000# diff_5500000_703000# diff_5631000_692000# GND efet w=89500 l=13500
+ ad=0 pd=0 as=-3.21967e+08 ps=740000 
M6084 diff_5631000_692000# diff_5617000_624000# diff_5618000_775000# GND efet w=221500 l=10500
+ ad=0 pd=0 as=2.13e+09 ps=286000 
M6085 diff_82000_3097000# diff_5695000_940000# diff_5599000_574000# GND efet w=291500 l=12500
+ ad=0 pd=0 as=0 ps=0 
M6086 diff_82000_3097000# diff_5695000_940000# diff_5599000_574000# GND efet w=290500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M6087 diff_5599000_574000# diff_5695000_940000# diff_82000_3097000# GND efet w=240500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M6088 diff_5695000_940000# diff_5695000_940000# diff_5695000_940000# GND efet w=3000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M6089 diff_5695000_940000# diff_5695000_940000# diff_94000_5193000# GND efet w=38000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M6090 diff_5339000_642000# diff_5339000_642000# diff_5323000_632000# GND efet w=15000 l=12000
+ ad=1.798e+09 pd=300000 as=0 ps=0 
M6091 diff_5339000_642000# diff_5388000_801000# diff_5388000_801000# GND efet w=17000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M6092 diff_94000_5193000# diff_5631000_692000# diff_5631000_692000# GND efet w=15000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M6093 diff_5654000_729000# diff_5645000_719000# diff_5652000_673000# GND efet w=30000 l=11000
+ ad=5.1e+08 pd=94000 as=1.151e+09 ps=210000 
M6094 diff_94000_5193000# diff_5768000_578000# diff_5768000_578000# GND efet w=46000 l=10000
+ ad=0 pd=0 as=1.14507e+09 ps=1.64e+06 
M6095 diff_82000_3097000# diff_5695000_940000# diff_5768000_578000# GND efet w=480000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M6096 diff_5599000_574000# diff_5768000_578000# diff_94000_5193000# GND efet w=287000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6097 diff_5956000_685000# diff_5768000_578000# diff_5599000_574000# GND efet w=287500 l=10500
+ ad=2.07e+09 pd=284000 as=0 ps=0 
M6098 diff_5652000_673000# diff_5631000_692000# diff_5631000_651000# GND efet w=44500 l=9500
+ ad=0 pd=0 as=1.024e+09 ps=174000 
M6099 diff_94000_5193000# diff_5652000_673000# diff_5652000_673000# GND efet w=14000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M6100 diff_5956000_636000# diff_5768000_578000# diff_5599000_574000# GND efet w=288000 l=10000
+ ad=1.946e+09 pd=282000 as=0 ps=0 
M6101 diff_94000_5193000# diff_5652000_673000# diff_5617000_624000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=1.245e+09 ps=246000 
M6102 diff_82000_3097000# diff_5760000_586000# diff_5768000_578000# GND efet w=487500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M6103 diff_5214000_614000# diff_4953000_397000# diff_5243000_579000# GND efet w=129000 l=13000
+ ad=0 pd=0 as=-1.2759e+09 ps=1.468e+06 
M6104 diff_4728000_545000# diff_4728000_566000# diff_4519000_195000# GND efet w=194500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M6105 diff_4805000_490000# diff_4728000_566000# diff_4519000_195000# GND efet w=186000 l=10000
+ ad=1.229e+09 pd=188000 as=0 ps=0 
M6106 diff_4763000_101000# diff_4728000_566000# diff_4519000_195000# GND efet w=183000 l=10000
+ ad=1.29629e+09 pd=3.654e+06 as=0 ps=0 
M6107 diff_4763000_101000# diff_4728000_566000# diff_4519000_195000# GND efet w=651500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M6108 diff_4966000_476000# diff_4943000_579000# diff_4941000_385000# GND efet w=560500 l=9500
+ ad=0 pd=0 as=-6.87902e+08 ps=1.754e+06 
M6109 diff_5617000_624000# diff_5507000_617000# diff_5609000_586000# GND efet w=21000 l=14000
+ ad=0 pd=0 as=-2.00197e+09 ps=396000 
M6110 diff_94000_5193000# diff_5609000_586000# diff_5609000_586000# GND efet w=14000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M6111 diff_5599000_574000# diff_5768000_578000# diff_5956000_580000# GND efet w=787000 l=10000
+ ad=0 pd=0 as=-1.7359e+09 ps=1.454e+06 
M6112 diff_4941000_385000# diff_5086000_471000# diff_4966000_476000# GND efet w=544000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6113 diff_5243000_579000# diff_4941000_385000# diff_5239000_451000# GND efet w=574500 l=10500
+ ad=0 pd=0 as=-1.1189e+09 ps=1.716e+06 
M6114 diff_5219000_459000# diff_4941000_385000# diff_4941000_385000# GND efet w=37000 l=11000
+ ad=8.54e+08 pd=182000 as=0 ps=0 
M6115 diff_5239000_451000# diff_5239000_451000# diff_5219000_459000# GND efet w=47000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6116 diff_5239000_451000# diff_5391000_471000# diff_5243000_579000# GND efet w=534500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M6117 diff_5609000_586000# diff_5599000_574000# diff_82000_3097000# GND efet w=149500 l=12500
+ ad=0 pd=0 as=0 ps=0 
M6118 diff_6411000_555000# diff_6411000_555000# diff_5599000_574000# GND efet w=99000 l=15000
+ ad=1.111e+09 pd=196000 as=0 ps=0 
M6119 diff_4953000_397000# diff_4941000_385000# diff_4763000_101000# GND efet w=243500 l=12500
+ ad=9.86294e+08 pd=5.36e+06 as=0 ps=0 
M6120 diff_4953000_397000# diff_4941000_385000# diff_4763000_101000# GND efet w=934500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M6121 diff_4953000_397000# diff_4941000_385000# diff_4763000_101000# GND efet w=418000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M6122 diff_4097000_195000# diff_4161000_584000# diff_4342000_102000# GND efet w=271000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6123 diff_4519000_195000# diff_4502000_545000# diff_4342000_102000# GND efet w=272000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6124 diff_4519000_195000# diff_4728000_566000# diff_4763000_101000# GND efet w=283000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6125 diff_5386000_199000# diff_5239000_451000# diff_5367000_123000# GND efet w=217000 l=10000
+ ad=-7.39869e+08 pd=2.16e+06 as=-1.73687e+09 ps=2.122e+06 
M6126 diff_5386000_199000# diff_5239000_451000# diff_5367000_123000# GND efet w=943000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6127 diff_5386000_199000# diff_5239000_451000# diff_5367000_123000# GND efet w=423500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M6128 diff_5607000_420000# diff_5595000_413000# diff_82000_3097000# GND efet w=145000 l=12000
+ ad=-1.58497e+09 pd=532000 as=0 ps=0 
M6129 diff_5768000_415000# diff_5256000_3172000# diff_82000_3097000# GND efet w=487000 l=11000
+ ad=7.12065e+08 pd=1.634e+06 as=0 ps=0 
M6130 diff_5607000_420000# diff_71000_4514000# diff_5617000_310000# GND efet w=22000 l=13000
+ ad=0 pd=0 as=1.188e+09 ps=240000 
M6131 diff_94000_5193000# diff_5607000_420000# diff_5607000_420000# GND efet w=15000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M6132 diff_94000_5193000# diff_5768000_415000# diff_5595000_413000# GND efet w=781000 l=10000
+ ad=0 pd=0 as=6.4636e+08 ps=7.01e+06 
M6133 diff_94000_5193000# diff_5652000_399000# diff_5617000_310000# GND efet w=15000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M6134 diff_5652000_399000# diff_5631000_321000# diff_82000_3097000# GND efet w=49000 l=10000
+ ad=1.132e+09 pd=210000 as=0 ps=0 
M6135 diff_5956000_434000# diff_5768000_415000# diff_5595000_413000# GND efet w=288000 l=10000
+ ad=1.946e+09 pd=282000 as=0 ps=0 
M6136 diff_5768000_415000# diff_5696000_134000# diff_82000_3097000# GND efet w=480000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6137 diff_5956000_384000# diff_5768000_415000# diff_5595000_413000# GND efet w=287500 l=10500
+ ad=2.07e+09 pd=284000 as=0 ps=0 
M6138 diff_94000_5193000# diff_5652000_399000# diff_5652000_399000# GND efet w=13000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M6139 diff_5652000_399000# diff_71000_4514000# diff_82000_3097000# GND efet w=30000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M6140 diff_5631000_321000# diff_5617000_310000# diff_82000_3097000# GND efet w=225500 l=10500
+ ad=-5.82967e+08 pd=734000 as=0 ps=0 
M6141 diff_94000_5193000# diff_5631000_321000# diff_5631000_321000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M6142 diff_5595000_413000# diff_5768000_415000# diff_94000_5193000# GND efet w=289000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6143 diff_6411000_452000# diff_6411000_452000# diff_5595000_413000# GND efet w=95000 l=15000
+ ad=1.018e+09 pd=180000 as=0 ps=0 
M6144 diff_5768000_415000# diff_5768000_415000# diff_94000_5193000# GND efet w=46000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6145 diff_94000_5193000# diff_5696000_134000# diff_5696000_134000# GND efet w=35000 l=10000
+ ad=0 pd=0 as=1.43307e+09 ps=1.798e+06 
M6146 diff_82000_3097000# diff_5696000_134000# diff_5595000_413000# GND efet w=241000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M6147 diff_5696000_134000# diff_5256000_3172000# diff_82000_3097000# GND efet w=477000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6148 diff_5631000_321000# diff_5555000_2636000# diff_5551000_265000# GND efet w=89000 l=13000
+ ad=0 pd=0 as=-1.78697e+09 ps=464000 
M6149 diff_82000_3097000# diff_5650000_134000# diff_5696000_134000# GND efet w=515000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M6150 diff_5551000_265000# diff_5576000_2597000# diff_5650000_134000# GND efet w=36000 l=14000
+ ad=0 pd=0 as=-1.44197e+09 ps=326000 
M6151 diff_82000_3097000# diff_5696000_134000# diff_5595000_413000# GND efet w=291000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M6152 diff_82000_3097000# diff_5696000_134000# diff_5595000_413000# GND efet w=292000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M6153 diff_5595000_413000# diff_5696000_134000# diff_82000_3097000# GND efet w=772500 l=11500
+ ad=0 pd=0 as=0 ps=0 
M6154 diff_5487000_89000# diff_5487000_89000# diff_4953000_397000# GND efet w=100500 l=13500
+ ad=1.433e+09 pd=200000 as=0 ps=0 
C0 metal_6090000_612000# gnd! 15.7fF ;**FLOATING
C1 metal_5920000_795000# gnd! 63.3fF ;**FLOATING
C2 metal_6090000_1404000# gnd! 15.7fF ;**FLOATING
C3 metal_6090000_2197000# gnd! 15.7fF ;**FLOATING
C4 metal_5920000_1587000# gnd! 63.3fF ;**FLOATING
C5 metal_5920000_2380000# gnd! 63.3fF ;**FLOATING
C6 metal_5418000_216000# gnd! 59.3fF ;**FLOATING
C7 metal_4964000_205000# gnd! 547.3fF ;**FLOATING
C8 metal_5253000_492000# gnd! 4.7fF ;**FLOATING
C9 metal_4565000_211000# gnd! 112.7fF ;**FLOATING
C10 metal_4144000_211000# gnd! 112.7fF ;**FLOATING
C11 metal_4024000_179000# gnd! 74.5fF ;**FLOATING
C12 metal_3735000_211000# gnd! 103.7fF ;**FLOATING
C13 metal_3314000_211000# gnd! 103.7fF ;**FLOATING
C14 metal_2506000_211000# gnd! 112.7fF ;**FLOATING
C15 metal_2097000_211000# gnd! 106.3fF ;**FLOATING
C16 metal_1676000_211000# gnd! 103.7fF ;**FLOATING
C17 metal_1266000_211000# gnd! 111.3fF ;**FLOATING
C18 metal_1142000_182000# gnd! 77.2fF ;**FLOATING
C19 metal_623000_199000# gnd! 137.8fF ;**FLOATING
C20 metal_808000_206000# gnd! 85.7fF ;**FLOATING
C21 metal_831000_251000# gnd! 209.7fF ;**FLOATING
C22 metal_752000_305000# gnd! 68.8fF ;**FLOATING
C23 metal_4754000_570000# gnd! 33.5fF ;**FLOATING
C24 metal_4157000_566000# gnd! 33.1fF ;**FLOATING
C25 metal_3923000_570000# gnd! 33.1fF ;**FLOATING
C26 metal_3326000_567000# gnd! 33.7fF ;**FLOATING
C27 metal_2519000_566000# gnd! 33.1fF ;**FLOATING
C28 metal_2285000_570000# gnd! 33.2fF ;**FLOATING
C29 metal_1688000_566000# gnd! 33.4fF ;**FLOATING
C30 metal_1454000_571000# gnd! 33.8fF ;**FLOATING
C31 metal_783000_608000# gnd! 163.7fF ;**FLOATING
C32 metal_5011000_580000# gnd! 88.3fF ;**FLOATING
C33 metal_784000_642000# gnd! 124.6fF ;**FLOATING
C34 metal_5277000_712000# gnd! 33.8fF ;**FLOATING
C35 metal_5546000_758000# gnd! 25.6fF ;**FLOATING
C36 metal_4957000_644000# gnd! 73.4fF ;**FLOATING
C37 metal_4337000_749000# gnd! 60.1fF ;**FLOATING
C38 metal_3249000_746000# gnd! 67.7fF ;**FLOATING
C39 metal_5550000_859000# gnd! 58.9fF ;**FLOATING
C40 metal_1842000_765000# gnd! 8.7fF ;**FLOATING
C41 metal_1777000_764000# gnd! 36.5fF ;**FLOATING
C42 metal_5009000_807000# gnd! 127.6fF ;**FLOATING
C43 metal_5185000_821000# gnd! 106.8fF ;**FLOATING
C44 metal_3267000_844000# gnd! 52.9fF ;**FLOATING
C45 metal_4076000_843000# gnd! 125.6fF ;**FLOATING
C46 metal_5393000_808000# gnd! 83.5fF ;**FLOATING
C47 metal_5207000_937000# gnd! 45.1fF ;**FLOATING
C48 metal_5097000_942000# gnd! 31.5fF ;**FLOATING
C49 metal_4692000_934000# gnd! 16.9fF ;**FLOATING
C50 metal_4708000_970000# gnd! 81.8fF ;**FLOATING
C51 metal_4460000_939000# gnd! 45.6fF ;**FLOATING
C52 metal_4332000_934000# gnd! 40.3fF ;**FLOATING
C53 metal_4432000_974000# gnd! 94.8fF ;**FLOATING
C54 metal_5004000_957000# gnd! 142.7fF ;**FLOATING
C55 metal_5525000_1024000# gnd! 73.8fF ;**FLOATING
C56 metal_5381000_963000# gnd! 87.3fF ;**FLOATING
C57 metal_4770000_999000# gnd! 75.8fF ;**FLOATING
C58 metal_4397000_993000# gnd! 38.0fF ;**FLOATING
C59 metal_4281000_977000# gnd! 39.8fF ;**FLOATING
C60 metal_4133000_935000# gnd! 79.4fF ;**FLOATING
C61 metal_4062000_967000# gnd! 34.7fF ;**FLOATING
C62 metal_3686000_939000# gnd! 29.6fF ;**FLOATING
C63 metal_3912000_954000# gnd! 23.6fF ;**FLOATING
C64 metal_3850000_968000# gnd! 42.3fF ;**FLOATING
C65 metal_3761000_935000# gnd! 41.3fF ;**FLOATING
C66 metal_3426000_935000# gnd! 29.6fF ;**FLOATING
C67 metal_3636000_951000# gnd! 22.2fF ;**FLOATING
C68 metal_3501000_935000# gnd! 36.6fF ;**FLOATING
C69 metal_3373000_963000# gnd! 23.9fF ;**FLOATING
C70 metal_3176000_935000# gnd! 32.4fF ;**FLOATING
C71 metal_3107000_935000# gnd! 34.3fF ;**FLOATING
C72 metal_3032000_952000# gnd! 37.8fF ;**FLOATING
C73 metal_2951000_964000# gnd! 28.2fF ;**FLOATING
C74 metal_2833000_934000# gnd! 30.1fF ;**FLOATING
C75 metal_2894000_965000# gnd! 36.5fF ;**FLOATING
C76 metal_2734000_934000# gnd! 36.4fF ;**FLOATING
C77 metal_2683000_961000# gnd! 32.8fF ;**FLOATING
C78 metal_2129000_936000# gnd! 73.9fF ;**FLOATING
C79 metal_1943000_933000# gnd! 28.4fF ;**FLOATING
C80 metal_2414000_963000# gnd! 46.6fF ;**FLOATING
C81 metal_2014000_938000# gnd! 42.9fF ;**FLOATING
C82 metal_1854000_945000# gnd! 27.6fF ;**FLOATING
C83 metal_1907000_960000# gnd! 30.9fF ;**FLOATING
C84 metal_4562000_1009000# gnd! 47.4fF ;**FLOATING
C85 metal_1481000_948000# gnd! 23.9fF ;**FLOATING
C86 metal_1661000_934000# gnd! 26.5fF ;**FLOATING
C87 metal_1590000_971000# gnd! 28.9fF ;**FLOATING
C88 metal_817000_912000# gnd! 493.7fF ;**FLOATING
C89 metal_1238000_978000# gnd! 99.8fF ;**FLOATING
C90 metal_1068000_940000# gnd! 55.6fF ;**FLOATING
C91 metal_893000_965000# gnd! 55.5fF ;**FLOATING
C92 metal_973000_1007000# gnd! 169.1fF ;**FLOATING
C93 metal_3581000_1011000# gnd! 313.2fF ;**FLOATING
C94 metal_4727000_1008000# gnd! 107.8fF ;**FLOATING
C95 metal_1833000_1002000# gnd! 121.5fF ;**FLOATING
C96 metal_4894000_1027000# gnd! 53.4fF ;**FLOATING
C97 metal_860000_1025000# gnd! 331.9fF ;**FLOATING
C98 metal_5382000_1122000# gnd! 57.4fF ;**FLOATING
C99 metal_4894000_1099000# gnd! 53.4fF ;**FLOATING
C100 metal_4727000_1099000# gnd! 111.3fF ;**FLOATING
C101 metal_4562000_1101000# gnd! 50.4fF ;**FLOATING
C102 metal_5097000_1176000# gnd! 47.3fF ;**FLOATING
C103 metal_5207000_1155000# gnd! 45.0fF ;**FLOATING
C104 metal_4994000_1167000# gnd! 156.2fF ;**FLOATING
C105 metal_4708000_1147000# gnd! 78.5fF ;**FLOATING
C106 metal_4692000_1189000# gnd! 13.8fF ;**FLOATING
C107 metal_4237000_1123000# gnd! 34.2fF ;**FLOATING
C108 metal_4438000_1149000# gnd! 93.9fF ;**FLOATING
C109 metal_4457000_1185000# gnd! 50.6fF ;**FLOATING
C110 metal_4328000_1126000# gnd! 57.0fF ;**FLOATING
C111 metal_2157000_1148000# gnd! 15.2fF ;**FLOATING
C112 metal_2014000_1151000# gnd! 41.7fF ;**FLOATING
C113 metal_1907000_1150000# gnd! 29.2fF ;**FLOATING
C114 metal_2359000_1182000# gnd! 36.8fF ;**FLOATING
C115 metal_2129000_1173000# gnd! 71.0fF ;**FLOATING
C116 metal_1943000_1178000# gnd! 28.4fF ;**FLOATING
C117 metal_1854000_1179000# gnd! 27.6fF ;**FLOATING
C118 metal_5381000_1340000# gnd! 56.8fF ;**FLOATING
C119 metal_5207000_1314000# gnd! 45.1fF ;**FLOATING
C120 metal_5097000_1319000# gnd! 31.5fF ;**FLOATING
C121 metal_4692000_1311000# gnd! 16.9fF ;**FLOATING
C122 metal_4708000_1347000# gnd! 80.5fF ;**FLOATING
C123 metal_4460000_1316000# gnd! 45.6fF ;**FLOATING
C124 metal_4133000_1312000# gnd! 70.0fF ;**FLOATING
C125 metal_4062000_1343000# gnd! 35.1fF ;**FLOATING
C126 metal_3686000_1316000# gnd! 29.6fF ;**FLOATING
C127 metal_3912000_1330000# gnd! 23.7fF ;**FLOATING
C128 metal_3850000_1345000# gnd! 42.3fF ;**FLOATING
C129 metal_3761000_1312000# gnd! 41.3fF ;**FLOATING
C130 metal_3426000_1311000# gnd! 31.1fF ;**FLOATING
C131 metal_3636000_1328000# gnd! 22.2fF ;**FLOATING
C132 metal_3501000_1312000# gnd! 37.0fF ;**FLOATING
C133 metal_3373000_1340000# gnd! 23.9fF ;**FLOATING
C134 metal_3107000_1312000# gnd! 32.5fF ;**FLOATING
C135 metal_3032000_1329000# gnd! 37.8fF ;**FLOATING
C136 metal_2951000_1341000# gnd! 28.2fF ;**FLOATING
C137 metal_2833000_1312000# gnd! 28.6fF ;**FLOATING
C138 metal_2894000_1342000# gnd! 35.1fF ;**FLOATING
C139 metal_2734000_1312000# gnd! 34.8fF ;**FLOATING
C140 metal_2683000_1338000# gnd! 34.3fF ;**FLOATING
C141 metal_1943000_1309000# gnd! 29.9fF ;**FLOATING
C142 metal_4432000_1351000# gnd! 94.8fF ;**FLOATING
C143 metal_4995000_1334000# gnd! 147.3fF ;**FLOATING
C144 metal_1854000_1322000# gnd! 28.1fF ;**FLOATING
C145 metal_2014000_1315000# gnd! 43.2fF ;**FLOATING
C146 metal_1907000_1336000# gnd! 30.9fF ;**FLOATING
C147 metal_4256000_1375000# gnd! 41.2fF ;**FLOATING
C148 metal_4562000_1386000# gnd! 47.4fF ;**FLOATING
C149 metal_1481000_1325000# gnd! 23.0fF ;**FLOATING
C150 metal_1661000_1311000# gnd! 26.5fF ;**FLOATING
C151 metal_1590000_1348000# gnd! 28.9fF ;**FLOATING
C152 metal_1263000_1314000# gnd! 79.3fF ;**FLOATING
C153 metal_1068000_1317000# gnd! 70.2fF ;**FLOATING
C154 metal_893000_1342000# gnd! 55.5fF ;**FLOATING
C155 metal_973000_1384000# gnd! 179.2fF ;**FLOATING
C156 metal_3581000_1388000# gnd! 314.1fF ;**FLOATING
C157 metal_4727000_1385000# gnd! 105.8fF ;**FLOATING
C158 metal_4894000_1404000# gnd! 53.4fF ;**FLOATING
C159 metal_860000_1401000# gnd! 335.1fF ;**FLOATING
C160 metal_5382000_1499000# gnd! 57.4fF ;**FLOATING
C161 metal_4894000_1476000# gnd! 53.4fF ;**FLOATING
C162 metal_4727000_1476000# gnd! 111.3fF ;**FLOATING
C163 metal_4562000_1478000# gnd! 50.4fF ;**FLOATING
C164 metal_5097000_1553000# gnd! 47.3fF ;**FLOATING
C165 metal_5207000_1532000# gnd! 167.0fF ;**FLOATING
C166 metal_4994000_1544000# gnd! 156.2fF ;**FLOATING
C167 metal_4708000_1524000# gnd! 78.5fF ;**FLOATING
C168 metal_4692000_1566000# gnd! 13.8fF ;**FLOATING
C169 metal_4440000_1530000# gnd! 93.5fF ;**FLOATING
C170 metal_4459000_1563000# gnd! 51.4fF ;**FLOATING
C171 metal_2157000_1525000# gnd! 12.3fF ;**FLOATING
C172 metal_2355000_1569000# gnd! 35.4fF ;**FLOATING
C173 metal_1907000_1527000# gnd! 30.9fF ;**FLOATING
C174 metal_2014000_1528000# gnd! 43.2fF ;**FLOATING
C175 metal_2129000_1549000# gnd! 60.8fF ;**FLOATING
C176 metal_1943000_1554000# gnd! 28.8fF ;**FLOATING
C177 metal_1854000_1556000# gnd! 27.6fF ;**FLOATING
C178 metal_5381000_1717000# gnd! 59.0fF ;**FLOATING
C179 metal_5207000_1690000# gnd! 48.2fF ;**FLOATING
C180 metal_5097000_1696000# gnd! 31.1fF ;**FLOATING
C181 metal_4692000_1688000# gnd! 9.5fF ;**FLOATING
C182 metal_4708000_1723000# gnd! 83.9fF ;**FLOATING
C183 metal_4460000_1693000# gnd! 49.9fF ;**FLOATING
C184 metal_4429000_1716000# gnd! 99.3fF ;**FLOATING
C185 metal_4133000_1689000# gnd! 62.8fF ;**FLOATING
C186 metal_4062000_1720000# gnd! 33.5fF ;**FLOATING
C187 metal_4995000_1710000# gnd! 147.4fF ;**FLOATING
C188 metal_4321000_1693000# gnd! 54.1fF ;**FLOATING
C189 metal_3686000_1693000# gnd! 29.6fF ;**FLOATING
C190 metal_3912000_1707000# gnd! 23.7fF ;**FLOATING
C191 metal_3426000_1688000# gnd! 31.1fF ;**FLOATING
C192 metal_3636000_1705000# gnd! 22.1fF ;**FLOATING
C193 metal_3501000_1688000# gnd! 38.3fF ;**FLOATING
C194 metal_3373000_1717000# gnd! 23.9fF ;**FLOATING
C195 metal_3107000_1689000# gnd! 32.8fF ;**FLOATING
C196 metal_3032000_1706000# gnd! 37.8fF ;**FLOATING
C197 metal_2951000_1718000# gnd! 28.2fF ;**FLOATING
C198 metal_2833000_1689000# gnd! 28.6fF ;**FLOATING
C199 metal_2894000_1719000# gnd! 35.1fF ;**FLOATING
C200 metal_3850000_1722000# gnd! 42.8fF ;**FLOATING
C201 metal_3761000_1688000# gnd! 41.8fF ;**FLOATING
C202 metal_2734000_1689000# gnd! 34.8fF ;**FLOATING
C203 metal_2683000_1715000# gnd! 32.8fF ;**FLOATING
C204 metal_1943000_1686000# gnd! 28.4fF ;**FLOATING
C205 metal_2014000_1691000# gnd! 41.8fF ;**FLOATING
C206 metal_1854000_1698000# gnd! 27.5fF ;**FLOATING
C207 metal_1907000_1713000# gnd! 29.2fF ;**FLOATING
C208 metal_4562000_1763000# gnd! 50.8fF ;**FLOATING
C209 metal_3581000_1764000# gnd! 179.7fF ;**FLOATING
C210 metal_1481000_1702000# gnd! 24.9fF ;**FLOATING
C211 metal_1661000_1688000# gnd! 26.5fF ;**FLOATING
C212 metal_1590000_1725000# gnd! 28.6fF ;**FLOATING
C213 metal_1265000_1702000# gnd! 79.8fF ;**FLOATING
C214 metal_1069000_1694000# gnd! 74.5fF ;**FLOATING
C215 metal_894000_1719000# gnd! 53.1fF ;**FLOATING
C216 metal_787000_1665000# gnd! 268.0fF ;**FLOATING
C217 metal_4727000_1762000# gnd! 113.0fF ;**FLOATING
C218 metal_1795000_1757000# gnd! 132.3fF ;**FLOATING
C219 metal_4894000_1781000# gnd! 53.4fF ;**FLOATING
C220 metal_860000_1778000# gnd! 350.5fF ;**FLOATING
C221 metal_5382000_1875000# gnd! 59.6fF ;**FLOATING
C222 metal_4894000_1853000# gnd! 53.4fF ;**FLOATING
C223 metal_4727000_1853000# gnd! 110.9fF ;**FLOATING
C224 metal_4562000_1855000# gnd! 47.4fF ;**FLOATING
C225 metal_5097000_1930000# gnd! 46.1fF ;**FLOATING
C226 metal_5523000_1856000# gnd! 54.3fF ;**FLOATING
C227 metal_5207000_1908000# gnd! 45.8fF ;**FLOATING
C228 metal_4994000_1921000# gnd! 159.2fF ;**FLOATING
C229 metal_4708000_1901000# gnd! 78.5fF ;**FLOATING
C230 metal_4692000_1943000# gnd! 2.5fF ;**FLOATING
C231 metal_4440000_1902000# gnd! 94.7fF ;**FLOATING
C232 metal_4459000_1939000# gnd! 48.2fF ;**FLOATING
C233 metal_2157000_1902000# gnd! 12.3fF ;**FLOATING
C234 metal_2014000_1905000# gnd! 41.7fF ;**FLOATING
C235 metal_1907000_1904000# gnd! 29.2fF ;**FLOATING
C236 metal_2339000_1941000# gnd! 41.6fF ;**FLOATING
C237 metal_2129000_1926000# gnd! 71.4fF ;**FLOATING
C238 metal_1943000_1932000# gnd! 27.2fF ;**FLOATING
C239 metal_1854000_1933000# gnd! 27.6fF ;**FLOATING
C240 metal_1219000_1902000# gnd! 32.9fF ;**FLOATING
C241 metal_786000_1790000# gnd! 277.3fF ;**FLOATING
C242 metal_894000_1912000# gnd! 53.1fF ;**FLOATING
C243 metal_1250000_1936000# gnd! 83.2fF ;**FLOATING
C244 metal_1069000_1938000# gnd! 69.5fF ;**FLOATING
C245 metal_5381000_2094000# gnd! 58.6fF ;**FLOATING
C246 metal_5207000_2068000# gnd! 45.0fF ;**FLOATING
C247 metal_5097000_2073000# gnd! 31.5fF ;**FLOATING
C248 metal_4692000_2065000# gnd! 16.5fF ;**FLOATING
C249 metal_4708000_2100000# gnd! 81.5fF ;**FLOATING
C250 metal_4460000_2077000# gnd! 50.9fF ;**FLOATING
C251 metal_4433000_2114000# gnd! 96.3fF ;**FLOATING
C252 metal_4133000_2066000# gnd! 62.4fF ;**FLOATING
C253 metal_4062000_2097000# gnd! 34.7fF ;**FLOATING
C254 metal_3686000_2070000# gnd! 29.6fF ;**FLOATING
C255 metal_3912000_2084000# gnd! 23.7fF ;**FLOATING
C256 metal_3426000_2065000# gnd! 31.1fF ;**FLOATING
C257 metal_3636000_2082000# gnd! 22.1fF ;**FLOATING
C258 metal_3501000_2065000# gnd! 38.3fF ;**FLOATING
C259 metal_3373000_2094000# gnd! 23.9fF ;**FLOATING
C260 metal_3107000_2066000# gnd! 32.8fF ;**FLOATING
C261 metal_3032000_2083000# gnd! 37.8fF ;**FLOATING
C262 metal_2951000_2095000# gnd! 28.2fF ;**FLOATING
C263 metal_2833000_2066000# gnd! 28.6fF ;**FLOATING
C264 metal_2894000_2096000# gnd! 35.1fF ;**FLOATING
C265 metal_3850000_2099000# gnd! 42.8fF ;**FLOATING
C266 metal_3761000_2065000# gnd! 41.8fF ;**FLOATING
C267 metal_2734000_2066000# gnd! 34.8fF ;**FLOATING
C268 metal_2683000_2092000# gnd! 32.8fF ;**FLOATING
C269 metal_1943000_2063000# gnd! 28.4fF ;**FLOATING
C270 metal_4995000_2087000# gnd! 147.6fF ;**FLOATING
C271 metal_2014000_2068000# gnd! 41.7fF ;**FLOATING
C272 metal_1854000_2075000# gnd! 28.2fF ;**FLOATING
C273 metal_1907000_2090000# gnd! 30.9fF ;**FLOATING
C274 metal_4562000_2140000# gnd! 50.4fF ;**FLOATING
C275 metal_3581000_2141000# gnd! 179.3fF ;**FLOATING
C276 metal_1661000_2065000# gnd! 26.0fF ;**FLOATING
C277 metal_1481000_2079000# gnd! 24.9fF ;**FLOATING
C278 metal_1590000_2102000# gnd! 28.6fF ;**FLOATING
C279 metal_1250000_2068000# gnd! 83.5fF ;**FLOATING
C280 metal_1219000_2103000# gnd! 40.2fF ;**FLOATING
C281 metal_1069000_2071000# gnd! 66.5fF ;**FLOATING
C282 metal_894000_2095000# gnd! 50.9fF ;**FLOATING
C283 metal_4727000_2139000# gnd! 109.6fF ;**FLOATING
C284 metal_4894000_2158000# gnd! 53.4fF ;**FLOATING
C285 metal_786000_2126000# gnd! 256.4fF ;**FLOATING
C286 metal_5382000_2252000# gnd! 59.6fF ;**FLOATING
C287 metal_4894000_2230000# gnd! 53.4fF ;**FLOATING
C288 metal_4727000_2230000# gnd! 110.8fF ;**FLOATING
C289 metal_4562000_2232000# gnd! 47.4fF ;**FLOATING
C290 metal_5097000_2307000# gnd! 46.1fF ;**FLOATING
C291 metal_5207000_2286000# gnd! 45.5fF ;**FLOATING
C292 metal_4994000_2298000# gnd! 157.0fF ;**FLOATING
C293 metal_4708000_2278000# gnd! 80.9fF ;**FLOATING
C294 metal_4692000_2320000# gnd! 14.1fF ;**FLOATING
C295 metal_4443000_2285000# gnd! 91.7fF ;**FLOATING
C296 metal_4513000_2316000# gnd! 27.7fF ;**FLOATING
C297 metal_2157000_2279000# gnd! 12.3fF ;**FLOATING
C298 metal_2014000_2282000# gnd! 42.8fF ;**FLOATING
C299 metal_1907000_2281000# gnd! 30.9fF ;**FLOATING
C300 metal_2129000_2303000# gnd! 66.1fF ;**FLOATING
C301 metal_2339000_2317000# gnd! 39.0fF ;**FLOATING
C302 metal_1943000_2308000# gnd! 28.8fF ;**FLOATING
C303 metal_1854000_2310000# gnd! 27.4fF ;**FLOATING
C304 metal_5382000_2450000# gnd! 31.3fF ;**FLOATING
C305 metal_4352000_2446000# gnd! 62.0fF ;**FLOATING
C306 metal_2329000_2464000# gnd! 48.7fF ;**FLOATING
C307 metal_2231000_2434000# gnd! 30.9fF ;**FLOATING
C308 metal_1121000_2414000# gnd! 93.4fF ;**FLOATING
C309 metal_1634000_2464000# gnd! 42.4fF ;**FLOATING
C310 metal_1060000_2414000# gnd! 62.1fF ;**FLOATING
C311 metal_4237000_2416000# gnd! 6.6fF ;**FLOATING
C312 metal_917000_2415000# gnd! 125.2fF ;**FLOATING
C313 metal_887000_2414000# gnd! 20.5fF ;**FLOATING
C314 metal_5127000_2637000# gnd! 25.4fF ;**FLOATING
C315 metal_5200000_2665000# gnd! 33.8fF ;**FLOATING
C316 metal_3053000_2614000# gnd! 120.6fF ;**FLOATING
C317 metal_1567000_2600000# gnd! 67.8fF ;**FLOATING
C318 metal_1280000_2610000# gnd! 238.8fF ;**FLOATING
C319 metal_1065000_2497000# gnd! 82.4fF ;**FLOATING
C320 metal_582000_319000# gnd! 82.6fF ;**FLOATING
C321 metal_564000_507000# gnd! 77.6fF ;**FLOATING
C322 metal_563000_690000# gnd! 163.4fF ;**FLOATING
C323 metal_555000_1277000# gnd! 117.0fF ;**FLOATING
C324 metal_563000_1444000# gnd! 148.1fF ;**FLOATING
C325 metal_187000_1256000# gnd! 118.9fF ;**FLOATING
C326 metal_555000_2031000# gnd! 117.0fF ;**FLOATING
C327 metal_563000_2198000# gnd! 147.2fF ;**FLOATING
C328 metal_1452000_2664000# gnd! 5.8fF ;**FLOATING
C329 metal_785000_2565000# gnd! 57.8fF ;**FLOATING
C330 metal_1237000_2700000# gnd! 97.1fF ;**FLOATING
C331 metal_187000_2011000# gnd! 117.2fF ;**FLOATING
C332 diff_5487000_89000# gnd! 266.0fF
C333 diff_5650000_134000# gnd! 631.3fF
C334 diff_5551000_265000# gnd! 357.8fF
C335 diff_5956000_384000# gnd! 235.4fF
C336 diff_5696000_134000# gnd! 2185.1fF
C337 diff_5956000_434000# gnd! 222.8fF
C338 diff_5631000_321000# gnd! 544.1fF
C339 diff_5652000_399000# gnd! 248.5fF
C340 diff_5617000_310000# gnd! 356.4fF
C341 diff_5768000_415000# gnd! 2146.0fF
C342 diff_5607000_420000# gnd! 360.9fF
C343 diff_6411000_452000# gnd! 227.0fF
C344 diff_5386000_199000# gnd! 1001.0fF
C345 diff_5367000_123000# gnd! 897.5fF
C346 diff_6411000_555000# gnd! 240.8fF
C347 diff_5391000_471000# gnd! 300.8fF
C348 diff_5219000_459000# gnd! 103.6fF
C349 diff_5239000_451000# gnd! 2277.4fF
C350 diff_5956000_580000# gnd! 830.8fF
C351 diff_5956000_636000# gnd! 222.8fF
C352 diff_5609000_586000# gnd! 301.9fF
C353 diff_5086000_471000# gnd! 311.6fF
C354 diff_4941000_385000# gnd! 2557.2fF
C355 diff_4763000_101000# gnd! 2213.0fF
C356 diff_4805000_490000# gnd! 141.7fF
C357 diff_5243000_579000# gnd! 878.2fF
C358 diff_5760000_586000# gnd! 285.6fF
C359 diff_5956000_685000# gnd! 235.4fF
C360 diff_5631000_651000# gnd! 119.8fF
C361 diff_5652000_673000# gnd! 246.8fF
C362 diff_5768000_578000# gnd! 2134.8fF
C363 diff_5645000_719000# gnd! 46.4fF
C364 diff_5654000_729000# gnd! 60.4fF
C365 diff_5507000_617000# gnd! 167.2fF
C366 diff_5618000_775000# gnd! 240.3fF
C367 diff_5631000_692000# gnd! 570.0fF
C368 diff_5617000_624000# gnd! 356.8fF
C369 diff_5500000_703000# gnd! 119.7fF
C370 diff_5417000_723000# gnd! 255.6fF
C371 diff_5339000_642000# gnd! 241.4fF
C372 diff_5201000_599000# gnd! 48.1fF
C373 diff_5214000_614000# gnd! 312.9fF
C374 diff_5105000_599000# gnd! 47.8fF
C375 diff_5114000_610000# gnd! 73.6fF
C376 diff_4966000_476000# gnd! 1179.2fF
C377 diff_5038000_606000# gnd! 323.1fF
C378 diff_5276000_709000# gnd! 139.6fF
C379 diff_5114000_586000# gnd! 396.6fF
C380 diff_4943000_579000# gnd! 551.5fF
C381 diff_4953000_638000# gnd! 61.8fF
C382 diff_5027000_596000# gnd! 547.5fF
C383 diff_5010000_575000# gnd! 82.3fF
C384 diff_5213000_671000# gnd! 142.0fF
C385 diff_5242000_710000# gnd! 114.3fF
C386 diff_5550000_857000# gnd! 258.2fF
C387 diff_5430000_735000# gnd! 66.5fF
C388 diff_5388000_801000# gnd! 463.4fF
C389 diff_5370000_762000# gnd! 214.8fF
C390 diff_5255000_745000# gnd! 297.6fF
C391 diff_5080000_704000# gnd! 181.3fF
C392 diff_5483000_731000# gnd! 197.3fF
C393 diff_5323000_632000# gnd! 424.8fF
C394 diff_5751000_807000# gnd! 277.4fF
C395 diff_5695000_940000# gnd! 2573.5fF
C396 diff_5650000_887000# gnd! 616.0fF
C397 diff_5650000_956000# gnd! 632.4fF
C398 diff_5696000_956000# gnd! 2224.5fF
C399 diff_5631000_1143000# gnd! 549.4fF
C400 diff_5556000_1019000# gnd! 146.1fF ;**FLOATING
C401 diff_5556000_1148000# gnd! 459.0fF
C402 diff_5652000_1221000# gnd! 250.6fF
C403 diff_5617000_1132000# gnd! 352.9fF
C404 diff_5270000_827000# gnd! 223.9fF
C405 diff_5342000_794000# gnd! 184.4fF
C406 diff_5243000_837000# gnd! 81.3fF
C407 diff_5153000_743000# gnd! 216.8fF
C408 diff_5119000_786000# gnd! 507.1fF
C409 diff_5097000_842000# gnd! 81.3fF
C410 diff_5079000_824000# gnd! 162.5fF
C411 diff_5055000_793000# gnd! 234.6fF
C412 diff_4920000_663000# gnd! 350.0fF
C413 diff_4790000_541000# gnd! 73.7fF
C414 diff_4697000_490000# gnd! 159.8fF
C415 diff_4644000_491000# gnd! 155.8fF
C416 diff_4591000_491000# gnd! 159.0fF
C417 diff_4342000_102000# gnd! 1382.0fF
C418 diff_4519000_195000# gnd! 3707.8fF
C419 diff_4728000_545000# gnd! 230.2fF
C420 diff_4384000_491000# gnd! 156.8fF
C421 diff_4331000_491000# gnd! 153.6fF
C422 diff_4278000_490000# gnd! 153.3fF
C423 diff_4802000_593000# gnd! 242.6fF
C424 diff_4846000_715000# gnd! 381.5fF
C425 diff_4836000_704000# gnd! 218.9fF
C426 diff_4728000_566000# gnd! 2131.5fF
C427 diff_4704000_651000# gnd! 282.7fF
C428 diff_4670000_619000# gnd! 56.6fF
C429 diff_4660000_692000# gnd! 56.8fF
C430 diff_4684000_624000# gnd! 484.7fF
C431 diff_4585000_578000# gnd! 323.5fF
C432 diff_4527000_661000# gnd! 372.3fF
C433 diff_4517000_655000# gnd! 253.6fF
C434 diff_4575000_567000# gnd! 375.6fF
C435 diff_4502000_545000# gnd! 2759.2fF
C436 diff_4168000_491000# gnd! 135.9fF
C437 diff_4097000_195000# gnd! 3724.3fF
C438 diff_3932000_101000# gnd! 887.8fF
C439 diff_3974000_491000# gnd! 141.6fF
C440 diff_4221000_545000# gnd! 226.1fF
C441 diff_4409000_635000# gnd! 376.1fF
C442 diff_4398000_625000# gnd! 252.4fF
C443 diff_4319000_578000# gnd! 321.2fF
C444 diff_4187000_542000# gnd! 83.2fF
C445 diff_4302000_667000# gnd! 56.6fF
C446 diff_4311000_567000# gnd! 371.4fF
C447 diff_4312000_692000# gnd! 54.6fF
C448 diff_4246000_637000# gnd! 294.9fF
C449 diff_4226000_612000# gnd! 459.9fF
C450 diff_4172000_589000# gnd! 243.2fF
C451 diff_4161000_584000# gnd! 2755.4fF
C452 diff_3959000_541000# gnd! 75.6fF
C453 diff_3866000_491000# gnd! 157.7fF
C454 diff_3814000_491000# gnd! 156.4fF
C455 diff_3761000_491000# gnd! 156.4fF
C456 diff_3511000_102000# gnd! 1427.5fF
C457 diff_3688000_195000# gnd! 3697.4fF
C458 diff_3898000_545000# gnd! 229.3fF
C459 diff_3554000_491000# gnd! 153.2fF
C460 diff_3500000_492000# gnd! 156.4fF
C461 diff_3447000_491000# gnd! 154.5fF
C462 diff_3338000_491000# gnd! 141.7fF
C463 diff_3266000_457000# gnd! 3702.4fF
C464 diff_3971000_593000# gnd! 251.5fF
C465 diff_4225000_699000# gnd! 52.8fF
C466 diff_4087000_122000# gnd! 2119.8fF
C467 diff_4110000_566000# gnd! 382.7fF
C468 diff_4100000_556000# gnd! 215.7fF
C469 diff_4015000_715000# gnd! 387.5fF
C470 diff_3874000_651000# gnd! 281.3fF
C471 diff_3840000_619000# gnd! 54.2fF
C472 diff_3829000_692000# gnd! 59.0fF
C473 diff_3921000_699000# gnd! 54.5fF
C474 diff_3853000_624000# gnd! 483.5fF
C475 diff_4005000_705000# gnd! 223.4fF
C476 diff_3898000_566000# gnd! 2120.5fF
C477 diff_3754000_578000# gnd! 327.7fF
C478 diff_3697000_661000# gnd! 357.8fF
C479 diff_3687000_625000# gnd! 255.4fF
C480 diff_3745000_567000# gnd! 369.2fF
C481 diff_3672000_544000# gnd! 2749.4fF
C482 diff_3391000_545000# gnd! 228.8fF
C483 diff_3579000_635000# gnd! 365.3fF
C484 diff_3568000_625000# gnd! 254.4fF
C485 diff_3357000_541000# gnd! 79.4fF
C486 diff_3472000_667000# gnd! 53.2fF
C487 diff_3489000_578000# gnd! 333.5fF
C488 diff_3482000_692000# gnd! 54.6fF
C489 diff_3481000_567000# gnd! 374.6fF
C490 diff_3416000_637000# gnd! 297.2fF
C491 diff_4751000_699000# gnd! 132.8fF
C492 diff_5008000_804000# gnd! 159.6fF
C493 diff_4977000_818000# gnd! 99.4fF
C494 diff_5008000_837000# gnd! 193.6fF
C495 diff_4962000_774000# gnd! 129.5fF
C496 diff_4890000_783000# gnd! 103.0fF
C497 diff_4772000_785000# gnd! 110.0fF
C498 diff_5069000_814000# gnd! 343.8fF
C499 diff_4775000_737000# gnd! 476.7fF
C500 diff_4950000_763000# gnd! 92.1fF
C501 diff_5384000_877000# gnd! 165.9fF
C502 diff_5524000_1020000# gnd! 151.9fF ;**FLOATING
C503 diff_5768000_1237000# gnd! 2137.3fF
C504 diff_5625000_1298000# gnd! 306.1fF
C505 diff_5618000_1308000# gnd! 3898.9fF
C506 diff_6411000_1274000# gnd! 465.2fF
C507 diff_5619000_1321000# gnd! 457.0fF
C508 diff_5956000_1373000# gnd! 788.7fF
C509 diff_5956000_1428000# gnd! 222.8fF
C510 diff_5625000_1391000# gnd! 269.4fF
C511 diff_5647000_1402000# gnd! 48.1fF
C512 diff_5760000_1378000# gnd! 285.6fF
C513 diff_5956000_1477000# gnd! 235.4fF
C514 diff_5631000_1443000# gnd! 113.8fF
C515 diff_5652000_1465000# gnd! 249.6fF
C516 diff_5768000_1367000# gnd! 2076.5fF
C517 diff_5645000_1511000# gnd! 46.4fF
C518 diff_5654000_1521000# gnd! 63.5fF
C519 diff_5618000_1380000# gnd! 4067.0fF
C520 diff_5619000_1567000# gnd! 236.0fF
C521 diff_5465000_917000# gnd! 170.0fF
C522 diff_5334000_891000# gnd! 22.6fF
C523 diff_5442000_999000# gnd! 112.7fF
C524 diff_5563000_1398000# gnd! 142.4fF ;**FLOATING
C525 diff_5355000_891000# gnd! 162.7fF
C526 diff_5376000_927000# gnd! 363.9fF
C527 diff_5442000_1118000# gnd! 112.2fF
C528 diff_5465000_1199000# gnd! 165.6fF
C529 diff_5358000_927000# gnd! 900.4fF
C530 diff_5376000_1197000# gnd! 372.1fF
C531 diff_5208000_877000# gnd! 100.7fF
C532 diff_5074000_876000# gnd! 104.2fF
C533 diff_5029000_876000# gnd! 52.2fF
C534 diff_5278000_904000# gnd! 87.8fF
C535 diff_5242000_886000# gnd! 315.3fF
C536 diff_5289000_913000# gnd! 162.4fF
C537 diff_5281000_1049000# gnd! 88.0fF
C538 diff_5200000_906000# gnd! 322.1fF
C539 diff_5233000_961000# gnd! 57.3fF
C540 diff_5124000_885000# gnd! 486.4fF
C541 diff_5068000_900000# gnd! 270.0fF
C542 diff_5037000_973000# gnd! 44.2fF
C543 diff_4837000_813000# gnd! 333.6fF
C544 diff_5161000_995000# gnd! 100.4fF
C545 diff_5136000_970000# gnd! 120.8fF
C546 diff_5068000_962000# gnd! 63.0fF
C547 diff_5202000_989000# gnd! 225.7fF
C548 diff_5243000_989000# gnd! 697.3fF
C549 diff_5281000_1081000# gnd! 88.0fF
C550 diff_5355000_1224000# gnd! 166.2fF
C551 diff_5335000_1224000# gnd! 19.6fF
C552 diff_4991000_889000# gnd! 543.5fF
C553 diff_4706000_839000# gnd! 236.9fF
C554 diff_4852000_874000# gnd! 139.2fF
C555 diff_4949000_896000# gnd! 200.0fF
C556 diff_4904000_951000# gnd! 146.1fF
C557 diff_4970000_889000# gnd! 215.7fF
C558 diff_4980000_886000# gnd! 107.3fF
C559 diff_5233000_1162000# gnd! 57.3fF
C560 diff_5289000_1091000# gnd! 159.6fF
C561 diff_5278000_1149000# gnd! 89.2fF
C562 diff_5201000_1209000# gnd! 322.8fF
C563 diff_5242000_1228000# gnd! 311.1fF
C564 diff_5070000_986000# gnd! 225.8fF
C565 diff_5111000_1009000# gnd! 775.5fF
C566 diff_5132000_1216000# gnd! 128.3fF
C567 diff_5068000_1155000# gnd! 63.5fF
C568 diff_5024000_982000# gnd! 312.3fF
C569 diff_4869000_938000# gnd! 524.4fF
C570 diff_4893000_1055000# gnd! 59.3fF
C571 diff_5037000_1132000# gnd! 43.8fF
C572 diff_5151000_1240000# gnd! 108.0fF
C573 diff_5124000_1236000# gnd! 900.9fF
C574 diff_5068000_1217000# gnd! 261.0fF
C575 diff_5021000_1214000# gnd! 282.1fF
C576 diff_5385000_1242000# gnd! 145.0fF
C577 diff_5465000_1294000# gnd! 167.7fF
C578 diff_5335000_1268000# gnd! 18.0fF
C579 diff_5442000_1375000# gnd! 111.7fF
C580 diff_5355000_1268000# gnd! 164.8fF
C581 diff_5376000_1304000# gnd! 370.1fF
C582 diff_5482000_1425000# gnd! 206.4fF
C583 diff_5497000_1490000# gnd! 224.6fF
C584 diff_5631000_1484000# gnd! 571.7fF
C585 diff_5617000_1426000# gnd! 350.6fF
C586 diff_5633000_1635000# gnd! 111.2fF
C587 diff_5688000_1661000# gnd! 55.2fF
C588 diff_5564000_1651000# gnd! 247.1fF
C589 diff_5751000_1599000# gnd! 277.4fF
C590 diff_5695000_1732000# gnd! 2594.2fF
C591 diff_5649000_1677000# gnd! 640.7fF
C592 diff_5649000_1748000# gnd! 644.6fF
C593 diff_5442000_1495000# gnd! 112.1fF
C594 diff_5465000_1576000# gnd! 166.1fF
C595 diff_5488000_1611000# gnd! 248.2fF
C596 diff_5358000_1304000# gnd! 891.2fF
C597 diff_5376000_1575000# gnd! 372.0fF
C598 diff_5208000_1234000# gnd! 174.5fF
C599 diff_5074000_1239000# gnd! 167.4fF
C600 diff_5028000_1241000# gnd! 79.3fF
C601 diff_5278000_1281000# gnd! 87.7fF
C602 diff_5242000_1263000# gnd! 315.1fF
C603 diff_5289000_1290000# gnd! 163.4fF
C604 diff_5281000_1426000# gnd! 87.8fF
C605 diff_5200000_1283000# gnd! 318.9fF
C606 diff_5233000_1338000# gnd! 56.6fF
C607 diff_4991000_1078000# gnd! 273.0fF
C608 diff_4971000_1103000# gnd! 199.9fF
C609 diff_4951000_1103000# gnd! 152.5fF
C610 diff_4692000_844000# gnd! 207.5fF
C611 diff_4692000_926000# gnd! 153.8fF
C612 diff_4638000_782000# gnd! 121.6fF
C613 diff_4643000_761000# gnd! 74.0fF
C614 diff_4585000_783000# gnd! 147.0fF
C615 diff_4302000_737000# gnd! 164.5fF
C616 diff_4573000_760000# gnd! 147.7fF
C617 diff_4588000_876000# gnd! 115.7fF
C618 diff_4831000_883000# gnd! 273.5fF
C619 diff_4809000_920000# gnd! 245.8fF
C620 diff_4706000_973000# gnd! 52.4fF
C621 diff_4672000_973000# gnd! 52.4fF
C622 diff_4405000_795000# gnd! 174.0fF
C623 diff_4530000_879000# gnd! 50.1fF
C624 diff_4726000_1005000# gnd! 262.3fF
C625 diff_4787000_982000# gnd! 210.1fF
C626 diff_4794000_778000# gnd! 182.2fF
C627 diff_4767000_995000# gnd! 112.2fF
C628 diff_4675000_1018000# gnd! 45.2fF
C629 diff_4706000_1018000# gnd! 123.8fF
C630 diff_4763000_779000# gnd! 185.9fF
C631 diff_4893000_1075000# gnd! 59.3fF
C632 diff_4866000_1100000# gnd! 342.7fF
C633 diff_4899000_1064000# gnd! 531.3fF
C634 diff_4982000_1073000# gnd! 91.7fF
C635 diff_4870000_1181000# gnd! 383.4fF
C636 diff_4904000_1167000# gnd! 142.0fF
C637 diff_5124000_1262000# gnd! 596.1fF
C638 diff_5068000_1277000# gnd! 266.6fF
C639 diff_5021000_1275000# gnd! 268.1fF
C640 diff_5037000_1351000# gnd! 43.8fF
C641 diff_5161000_1372000# gnd! 99.8fF
C642 diff_5136000_1347000# gnd! 121.5fF
C643 diff_5068000_1339000# gnd! 63.0fF
C644 diff_5202000_1366000# gnd! 226.8fF
C645 diff_5243000_1366000# gnd! 698.3fF
C646 diff_5281000_1458000# gnd! 87.9fF
C647 diff_5355000_1601000# gnd! 166.2fF
C648 diff_5334000_1601000# gnd! 21.1fF
C649 diff_5233000_1540000# gnd! 57.5fF
C650 diff_4991000_1272000# gnd! 259.0fF
C651 diff_4952000_1272000# gnd! 138.6fF
C652 diff_4881000_1243000# gnd! 75.2fF
C653 diff_4831000_1174000# gnd! 273.5fF
C654 diff_4809000_1139000# gnd! 251.2fF
C655 diff_4786000_1098000# gnd! 190.4fF
C656 diff_4675000_1096000# gnd! 47.1fF
C657 diff_4563000_975000# gnd! 47.1fF
C658 diff_4574000_899000# gnd! 254.8fF
C659 diff_4624000_962000# gnd! 61.1fF
C660 diff_4607000_945000# gnd! 345.2fF
C661 diff_4706000_1096000# gnd! 124.1fF
C662 diff_4706000_1141000# gnd! 52.1fF
C663 diff_4672000_1141000# gnd! 54.6fF
C664 diff_4617000_986000# gnd! 325.0fF
C665 diff_4517000_900000# gnd! 266.4fF
C666 diff_4532000_955000# gnd! 55.6fF
C667 diff_4477000_914000# gnd! 282.8fF
C668 diff_4393000_785000# gnd! 129.6fF
C669 diff_4423000_931000# gnd! 52.4fF
C670 diff_4481000_1020000# gnd! 41.3fF
C671 diff_4423000_963000# gnd! 136.5fF
C672 diff_4413000_1027000# gnd! 80.4fF
C673 diff_4480000_1097000# gnd! 46.6fF
C674 diff_4753000_1054000# gnd! 632.3fF
C675 diff_4726000_1105000# gnd! 261.5fF
C676 diff_4693000_1184000# gnd! 159.2fF
C677 diff_4820000_1150000# gnd! 112.3fF
C678 diff_4798000_1130000# gnd! 113.3fF
C679 diff_4971000_1272000# gnd! 199.7fF
C680 diff_4982000_1267000# gnd! 91.7fF
C681 diff_5289000_1468000# gnd! 159.5fF
C682 diff_5278000_1526000# gnd! 89.2fF
C683 diff_5201000_1587000# gnd! 322.7fF
C684 diff_5242000_1606000# gnd! 303.1fF
C685 diff_5070000_1364000# gnd! 224.8fF
C686 diff_5111000_1386000# gnd! 772.5fF
C687 diff_5132000_1593000# gnd! 129.5fF
C688 diff_5068000_1533000# gnd! 64.4fF
C689 diff_5024000_1356000# gnd! 313.3fF
C690 diff_4904000_1328000# gnd! 149.8fF
C691 diff_4869000_1327000# gnd! 410.1fF
C692 diff_4893000_1432000# gnd! 59.3fF
C693 diff_5037000_1510000# gnd! 44.1fF
C694 diff_5151000_1618000# gnd! 107.3fF
C695 diff_5124000_1613000# gnd! 595.5fF
C696 diff_5068000_1594000# gnd! 260.5fF
C697 diff_5021000_1591000# gnd! 279.8fF
C698 diff_5158000_1629000# gnd! 275.4fF
C699 diff_5385000_1619000# gnd! 142.9fF
C700 diff_5465000_1671000# gnd! 176.5fF
C701 diff_5334000_1644000# gnd! 20.3fF
C702 diff_5442000_1752000# gnd! 111.7fF
C703 diff_5509000_1567000# gnd! 203.3fF ;**FLOATING
C704 diff_5696000_1748000# gnd! 2666.6fF
C705 diff_5631000_1935000# gnd! 550.9fF
C706 diff_5569000_1916000# gnd! 374.1fF
C707 diff_5652000_2013000# gnd! 250.7fF
C708 diff_5617000_1924000# gnd! 350.9fF
C709 diff_5768000_2029000# gnd! 2154.8fF
C710 diff_5625000_2090000# gnd! 305.9fF
C711 diff_5618000_2101000# gnd! 4308.1fF
C712 diff_5956000_2165000# gnd! 630.3fF
C713 diff_5619000_2114000# gnd! 452.8fF
C714 diff_5956000_2221000# gnd! 222.8fF
C715 diff_5625000_2183000# gnd! 278.9fF
C716 diff_5647000_2195000# gnd! 49.8fF
C717 diff_5760000_2171000# gnd! 288.9fF
C718 diff_5956000_2270000# gnd! 232.9fF
C719 diff_5630000_2236000# gnd! 114.4fF
C720 diff_5652000_2258000# gnd! 253.7fF
C721 diff_5768000_2160000# gnd! 2094.8fF
C722 diff_5645000_2303000# gnd! 46.4fF
C723 diff_5654000_2314000# gnd! 57.2fF
C724 diff_5476000_1801000# gnd! 150.0fF
C725 diff_5355000_1644000# gnd! 163.3fF
C726 diff_5376000_1680000# gnd! 370.9fF
C727 diff_5484000_1775000# gnd! 80.2fF
C728 diff_5472000_1599000# gnd! 544.8fF
C729 diff_5442000_1872000# gnd! 111.4fF
C730 diff_5465000_1953000# gnd! 173.9fF
C731 diff_5476000_1993000# gnd! 259.6fF
C732 diff_5520000_2087000# gnd! 181.0fF
C733 diff_5358000_1681000# gnd! 896.3fF
C734 diff_5376000_1951000# gnd! 371.1fF
C735 diff_5208000_1611000# gnd! 172.8fF
C736 diff_5074000_1617000# gnd! 167.3fF
C737 diff_5028000_1618000# gnd! 79.6fF
C738 diff_5278000_1658000# gnd! 89.0fF
C739 diff_5242000_1640000# gnd! 316.0fF
C740 diff_5289000_1667000# gnd! 161.7fF
C741 diff_5281000_1802000# gnd! 88.0fF
C742 diff_5200000_1659000# gnd! 321.1fF
C743 diff_5233000_1714000# gnd! 57.5fF
C744 diff_4991000_1456000# gnd! 265.8fF
C745 diff_4971000_1481000# gnd! 198.7fF
C746 diff_4951000_1481000# gnd! 151.4fF
C747 diff_4831000_1268000# gnd! 268.6fF
C748 diff_4701000_1242000# gnd! 212.0fF
C749 diff_4692000_1303000# gnd! 152.7fF
C750 diff_4624000_1155000# gnd! 61.1fF
C751 diff_4563000_1140000# gnd! 45.2fF
C752 diff_4607000_1092000# gnd! 347.0fF
C753 diff_4574000_1196000# gnd! 258.6fF
C754 diff_4588000_1240000# gnd! 174.6fF
C755 diff_4706000_1350000# gnd! 52.4fF
C756 diff_4672000_1350000# gnd! 52.4fF
C757 diff_4519000_996000# gnd! 327.6fF
C758 diff_4532000_1098000# gnd! 55.6fF
C759 diff_4517000_1195000# gnd! 274.4fF
C760 diff_4460000_935000# gnd! 257.6fF
C761 diff_4379000_974000# gnd! 131.9fF
C762 diff_4329000_909000# gnd! 159.2fF
C763 diff_4073000_749000# gnd! 256.8fF
C764 diff_4194000_784000# gnd! 147.3fF
C765 diff_4182000_762000# gnd! 147.0fF
C766 diff_4264000_908000# gnd! 363.6fF ;**FLOATING
C767 diff_4120000_825000# gnd! 88.8fF
C768 diff_4046000_762000# gnd! 90.8fF
C769 diff_4044000_822000# gnd! 269.2fF
C770 diff_3395000_613000# gnd! 468.3fF
C771 diff_3395000_699000# gnd! 50.5fF
C772 diff_3341000_590000# gnd! 250.7fF
C773 diff_2875000_456000# gnd! 1009.2fF
C774 diff_2705000_101000# gnd! 1372.6fF
C775 diff_2746000_491000# gnd! 156.8fF
C776 diff_2693000_491000# gnd! 153.5fF
C777 diff_2639000_491000# gnd! 157.8fF
C778 diff_2530000_491000# gnd! 141.6fF
C779 diff_2295000_101000# gnd! 884.5fF
C780 diff_2336000_490000# gnd! 141.9fF
C781 diff_2459000_132000# gnd! 3727.8fF
C782 diff_2583000_545000# gnd! 229.7fF
C783 diff_3331000_584000# gnd! 2761.4fF
C784 diff_3257000_122000# gnd! 2088.6fF
C785 diff_2771000_635000# gnd! 376.1fF
C786 diff_2760000_625000# gnd! 252.5fF
C787 diff_2681000_578000# gnd! 321.1fF
C788 diff_2549000_541000# gnd! 83.2fF
C789 diff_2664000_667000# gnd! 56.6fF
C790 diff_2675000_692000# gnd! 52.4fF
C791 diff_2673000_567000# gnd! 377.2fF
C792 diff_2608000_637000# gnd! 294.9fF
C793 diff_3279000_567000# gnd! 386.8fF
C794 diff_3269000_556000# gnd! 219.9fF
C795 diff_2588000_612000# gnd! 457.2fF
C796 diff_2534000_589000# gnd! 243.6fF
C797 diff_2523000_584000# gnd! 2762.1fF
C798 diff_2321000_541000# gnd! 77.6fF
C799 diff_2228000_491000# gnd! 154.5fF
C800 diff_2176000_491000# gnd! 156.4fF
C801 diff_2122000_492000# gnd! 153.2fF
C802 diff_1873000_101000# gnd! 1417.8fF
C803 diff_2050000_195000# gnd! 3684.6fF
C804 diff_2260000_545000# gnd! 231.4fF
C805 diff_1915000_492000# gnd! 156.4fF
C806 diff_1862000_492000# gnd! 156.4fF
C807 diff_1809000_491000# gnd! 157.7fF
C808 diff_1699000_492000# gnd! 141.7fF
C809 diff_1465000_100000# gnd! 906.0fF
C810 diff_1506000_490000# gnd! 138.1fF
C811 diff_1628000_457000# gnd! 3707.6fF
C812 diff_2333000_592000# gnd! 252.2fF
C813 diff_2587000_700000# gnd! 50.8fF
C814 diff_2449000_122000# gnd! 2116.0fF
C815 diff_2472000_566000# gnd! 375.1fF
C816 diff_2461000_557000# gnd! 220.2fF
C817 diff_2377000_715000# gnd! 384.5fF
C818 diff_2367000_705000# gnd! 223.5fF
C819 diff_2260000_566000# gnd! 2118.8fF
C820 diff_2236000_651000# gnd! 279.1fF
C821 diff_2202000_619000# gnd! 53.2fF
C822 diff_2191000_692000# gnd! 59.0fF
C823 diff_2283000_699000# gnd! 54.9fF
C824 diff_2215000_624000# gnd! 476.6fF
C825 diff_2116000_578000# gnd! 335.9fF
C826 diff_2059000_661000# gnd! 357.8fF
C827 diff_2049000_625000# gnd! 255.4fF
C828 diff_2107000_567000# gnd! 367.0fF
C829 diff_2034000_544000# gnd! 2752.6fF
C830 diff_1753000_545000# gnd! 224.1fF
C831 diff_1941000_635000# gnd! 364.2fF
C832 diff_1930000_625000# gnd! 254.3fF
C833 diff_1850000_578000# gnd! 325.2fF
C834 diff_1719000_540000# gnd! 83.5fF
C835 diff_1833000_667000# gnd! 54.2fF
C836 diff_1843000_567000# gnd! 379.8fF
C837 diff_1844000_692000# gnd! 54.6fF
C838 diff_1778000_637000# gnd! 297.3fF
C839 diff_3947000_785000# gnd! 201.6fF
C840 diff_3930000_764000# gnd! 91.0fF
C841 diff_4317000_839000# gnd! 105.5fF
C842 diff_4433000_1143000# gnd! 105.6fF
C843 diff_4378000_1100000# gnd! 139.7fF
C844 diff_4458000_1182000# gnd! 118.7fF
C845 diff_4406000_1189000# gnd! 165.1fF
C846 diff_4531000_1239000# gnd! 90.1fF
C847 diff_4726000_1382000# gnd! 262.5fF
C848 diff_4809000_1268000# gnd! 245.1fF
C849 diff_4787000_1407000# gnd! 197.9fF
C850 diff_4820000_1262000# gnd! 112.3fF
C851 diff_4799000_1262000# gnd! 104.0fF
C852 diff_4893000_1452000# gnd! 60.4fF
C853 diff_4675000_1395000# gnd! 47.1fF
C854 diff_4706000_1395000# gnd! 122.5fF
C855 diff_4866000_1360000# gnd! 358.8fF
C856 diff_4899000_1441000# gnd! 573.0fF
C857 diff_4982000_1450000# gnd! 91.6fF
C858 diff_4870000_1558000# gnd! 389.8fF
C859 diff_4904000_1545000# gnd! 142.8fF
C860 diff_5124000_1640000# gnd! 309.6fF
C861 diff_5068000_1654000# gnd! 264.7fF
C862 diff_5021000_1652000# gnd! 267.6fF
C863 diff_5037000_1727000# gnd! 44.2fF
C864 diff_5136000_1724000# gnd! 120.2fF
C865 diff_5161000_1749000# gnd! 100.0fF
C866 diff_5068000_1716000# gnd! 62.1fF
C867 diff_5202000_1742000# gnd! 226.8fF
C868 diff_5243000_1742000# gnd! 701.0fF
C869 diff_5281000_1835000# gnd! 87.2fF
C870 diff_5355000_1977000# gnd! 167.2fF
C871 diff_5335000_1977000# gnd! 19.5fF
C872 diff_5289000_1845000# gnd! 158.3fF
C873 diff_5233000_1916000# gnd! 56.6fF
C874 diff_4991000_1650000# gnd! 260.5fF
C875 diff_4952000_1650000# gnd! 138.6fF
C876 diff_4881000_1621000# gnd! 75.7fF
C877 diff_4831000_1552000# gnd! 273.2fF
C878 diff_4809000_1516000# gnd! 252.6fF
C879 diff_4787000_1475000# gnd! 202.4fF
C880 diff_4675000_1474000# gnd! 45.2fF
C881 diff_4563000_1352000# gnd! 47.1fF
C882 diff_4574000_1276000# gnd! 257.0fF
C883 diff_4624000_1339000# gnd! 61.6fF
C884 diff_4607000_1322000# gnd! 344.2fF
C885 diff_4706000_1474000# gnd! 122.2fF
C886 diff_4706000_1518000# gnd! 52.1fF
C887 diff_4672000_1518000# gnd! 54.6fF
C888 diff_4617000_1363000# gnd! 325.1fF
C889 diff_4517000_1277000# gnd! 266.8fF
C890 diff_4532000_1332000# gnd! 55.6fF
C891 diff_4477000_1119000# gnd! 523.5fF
C892 diff_4481000_1400000# gnd! 40.8fF
C893 diff_4432000_1347000# gnd! 189.5fF
C894 diff_4308000_1009000# gnd! 115.1fF
C895 diff_4165000_930000# gnd! 101.8fF
C896 diff_4126000_876000# gnd! 63.5fF
C897 diff_3993000_764000# gnd! 67.5fF
C898 diff_3907000_737000# gnd! 183.8fF
C899 diff_3856000_786000# gnd! 150.5fF
C900 diff_3836000_763000# gnd! 133.4fF
C901 diff_4052000_838000# gnd! 111.8fF
C902 diff_4052000_893000# gnd! 207.7fF
C903 diff_3960000_872000# gnd! 50.4fF
C904 diff_4005000_919000# gnd! 52.4fF
C905 diff_3741000_766000# gnd! 211.3fF
C906 diff_3717000_755000# gnd! 173.6fF
C907 diff_3664000_845000# gnd! 184.4fF
C908 diff_3604000_815000# gnd! 206.2fF
C909 diff_3586000_784000# gnd! 246.5fF
C910 diff_3886000_876000# gnd! 63.4fF
C911 diff_3884000_904000# gnd! 204.1fF
C912 diff_4184000_1005000# gnd! 210.5fF
C913 diff_4280000_938000# gnd! 794.5fF
C914 diff_4288000_1116000# gnd! 84.0fF
C915 diff_4204000_1036000# gnd! 363.7fF
C916 diff_4149000_968000# gnd! 136.1fF
C917 diff_4057000_979000# gnd! 118.3fF
C918 diff_4037000_919000# gnd! 195.4fF
C919 diff_4067000_1029000# gnd! 334.5fF
C920 diff_4056000_1019000# gnd! 132.3fF
C921 diff_4306000_1186000# gnd! 357.1fF
C922 diff_4232000_995000# gnd! 129.6fF
C923 diff_4314000_1211000# gnd! 147.2fF
C924 diff_4224000_1220000# gnd! 396.9fF
C925 diff_4228000_1258000# gnd! 40.8fF
C926 diff_4276000_1307000# gnd! 108.3fF
C927 diff_4317000_998000# gnd! 389.4fF
C928 diff_4379000_1393000# gnd! 137.6fF
C929 diff_4480000_1474000# gnd! 46.9fF
C930 diff_4726000_1482000# gnd! 263.9fF
C931 diff_4693000_1562000# gnd! 157.2fF
C932 diff_4753000_1432000# gnd! 671.2fF
C933 diff_4820000_1527000# gnd! 111.4fF
C934 diff_4798000_1507000# gnd! 113.3fF
C935 diff_4971000_1650000# gnd! 199.9fF
C936 diff_4982000_1643000# gnd! 91.6fF
C937 diff_5278000_1902000# gnd! 88.8fF
C938 diff_5201000_1963000# gnd! 324.1fF
C939 diff_5242000_1982000# gnd! 308.0fF
C940 diff_5070000_1741000# gnd! 224.8fF
C941 diff_5111000_1762000# gnd! 772.5fF
C942 diff_5132000_1970000# gnd! 127.2fF
C943 diff_5068000_1909000# gnd! 63.5fF
C944 diff_5024000_1733000# gnd! 313.3fF
C945 diff_4904000_1705000# gnd! 149.6fF
C946 diff_4869000_1704000# gnd! 410.1fF
C947 diff_4893000_1809000# gnd! 59.3fF
C948 diff_5037000_1886000# gnd! 43.8fF
C949 diff_5151000_1994000# gnd! 108.0fF
C950 diff_5124000_1991000# gnd! 596.8fF
C951 diff_5068000_1971000# gnd! 252.9fF
C952 diff_5021000_1967000# gnd! 279.6fF
C953 diff_5385000_1996000# gnd! 144.4fF
C954 diff_5510000_2076000# gnd! 129.6fF
C955 diff_5619000_2361000# gnd! 237.0fF
C956 diff_5631000_2275000# gnd! 578.0fF
C957 diff_5617000_2218000# gnd! 342.1fF
C958 diff_5633000_2428000# gnd! 104.8fF
C959 diff_5562000_2269000# gnd! 484.0fF
C960 diff_5688000_2454000# gnd! 54.2fF
C961 diff_5751000_2392000# gnd! 275.5fF
C962 diff_5695000_2525000# gnd! 2552.8fF
C963 diff_5650000_2471000# gnd! 622.1fF
C964 diff_5465000_2048000# gnd! 174.3fF
C965 diff_5335000_2021000# gnd! 18.0fF
C966 diff_5442000_2129000# gnd! 111.9fF
C967 diff_5355000_2021000# gnd! 164.5fF
C968 diff_5376000_2057000# gnd! 370.5fF
C969 diff_5442000_2249000# gnd! 111.9fF
C970 diff_5465000_2330000# gnd! 172.7fF
C971 diff_5358000_2058000# gnd! 893.7fF
C972 diff_5376000_2328000# gnd! 371.9fF
C973 diff_5208000_1988000# gnd! 172.8fF
C974 diff_5074000_1993000# gnd! 166.8fF
C975 diff_5028000_1995000# gnd! 79.2fF
C976 diff_5278000_2035000# gnd! 87.8fF
C977 diff_5242000_2017000# gnd! 320.3fF
C978 diff_5289000_2044000# gnd! 163.2fF
C979 diff_5281000_2180000# gnd! 86.1fF
C980 diff_5200000_2037000# gnd! 320.8fF
C981 diff_5233000_2092000# gnd! 57.3fF
C982 diff_4991000_1833000# gnd! 268.0fF
C983 diff_4971000_1858000# gnd! 199.9fF
C984 diff_4951000_1858000# gnd! 152.5fF
C985 diff_4831000_1646000# gnd! 267.0fF
C986 diff_4701000_1619000# gnd! 211.5fF
C987 diff_4692000_1680000# gnd! 156.6fF
C988 diff_4624000_1532000# gnd! 61.6fF
C989 diff_4563000_1518000# gnd! 45.1fF
C990 diff_4607000_1470000# gnd! 351.0fF
C991 diff_4574000_1573000# gnd! 259.9fF
C992 diff_4588000_1617000# gnd! 169.6fF
C993 diff_4706000_1727000# gnd! 52.4fF
C994 diff_4672000_1727000# gnd! 52.4fF
C995 diff_4519000_1373000# gnd! 329.3fF
C996 diff_4532000_1475000# gnd! 55.6fF
C997 diff_4517000_1572000# gnd! 271.5fF
C998 diff_4459000_1490000# gnd! 263.1fF
C999 diff_4435000_1490000# gnd! 87.6fF
C1000 diff_4531000_1616000# gnd! 90.8fF
C1001 diff_4412000_1466000# gnd! 268.8fF
C1002 diff_4460000_1561000# gnd! 141.3fF
C1003 diff_4726000_1760000# gnd! 264.1fF
C1004 diff_4809000_1646000# gnd! 252.5fF
C1005 diff_4787000_1783000# gnd! 211.4fF
C1006 diff_4799000_1639000# gnd! 102.8fF
C1007 diff_4821000_1638000# gnd! 107.0fF
C1008 diff_4893000_1829000# gnd! 59.3fF
C1009 diff_4675000_1772000# gnd! 45.2fF
C1010 diff_4706000_1772000# gnd! 123.8fF
C1011 diff_4866000_1738000# gnd! 359.8fF
C1012 diff_4899000_1818000# gnd! 573.7fF
C1013 diff_4870000_1933000# gnd! 393.4fF
C1014 diff_4982000_1826000# gnd! 92.1fF
C1015 diff_4904000_1921000# gnd! 141.5fF
C1016 diff_5124000_2017000# gnd! 597.1fF
C1017 diff_5068000_2031000# gnd! 268.6fF
C1018 diff_5021000_2029000# gnd! 269.6fF
C1019 diff_5037000_2104000# gnd! 44.2fF
C1020 diff_5161000_2126000# gnd! 100.4fF
C1021 diff_5136000_2101000# gnd! 120.8fF
C1022 diff_5068000_2093000# gnd! 62.5fF
C1023 diff_5202000_2119000# gnd! 227.6fF
C1024 diff_5243000_2120000# gnd! 701.2fF
C1025 diff_5281000_2212000# gnd! 88.0fF
C1026 diff_5385000_2373000# gnd! 83.1fF
C1027 diff_5355000_2355000# gnd! 165.7fF
C1028 diff_5334000_2356000# gnd! 23.5fF
C1029 diff_5233000_2294000# gnd! 57.2fF
C1030 diff_4991000_2027000# gnd! 259.5fF
C1031 diff_4952000_2027000# gnd! 138.6fF
C1032 diff_4881000_1998000# gnd! 76.8fF
C1033 diff_4831000_1929000# gnd! 274.6fF
C1034 diff_4809000_1892000# gnd! 252.7fF
C1035 diff_4787000_1852000# gnd! 202.6fF
C1036 diff_4675000_1850000# gnd! 47.1fF
C1037 diff_4563000_1729000# gnd! 47.1fF
C1038 diff_4574000_1652000# gnd! 256.1fF
C1039 diff_4624000_1715000# gnd! 62.6fF
C1040 diff_4607000_1699000# gnd! 346.8fF
C1041 diff_4706000_1850000# gnd! 124.0fF
C1042 diff_4706000_1895000# gnd! 52.1fF
C1043 diff_4672000_1895000# gnd! 54.6fF
C1044 diff_4617000_1740000# gnd! 323.9fF
C1045 diff_4517000_1654000# gnd! 267.4fF
C1046 diff_4532000_1709000# gnd! 56.1fF
C1047 diff_4477000_1497000# gnd! 523.3fF
C1048 diff_4481000_1777000# gnd! 40.8fF
C1049 diff_4429000_1713000# gnd! 174.0fF
C1050 diff_4373000_1474000# gnd! 128.9fF
C1051 diff_4262000_1287000# gnd! 677.5fF
C1052 diff_4185000_1075000# gnd! 181.3fF
C1053 diff_4166000_1185000# gnd! 112.4fF
C1054 diff_4067000_1099000# gnd! 419.3fF
C1055 diff_3949000_962000# gnd! 125.5fF
C1056 diff_3938000_928000# gnd! 185.3fF
C1057 diff_3881000_929000# gnd! 321.7fF
C1058 diff_3847000_947000# gnd! 143.8fF
C1059 diff_3819000_912000# gnd! 148.4fF
C1060 diff_3758000_876000# gnd! 63.5fF
C1061 diff_3473000_771000# gnd! 206.8fF
C1062 diff_3526000_822000# gnd! 135.5fF
C1063 diff_3684000_872000# gnd! 48.4fF
C1064 diff_3683000_893000# gnd! 201.1fF
C1065 diff_3659000_908000# gnd! 51.6fF
C1066 diff_3361000_767000# gnd! 282.3fF
C1067 diff_3411000_824000# gnd! 131.8fF
C1068 diff_3334000_772000# gnd! 81.0fF
C1069 diff_3795000_966000# gnd! 130.7fF
C1070 diff_3864000_1014000# gnd! 111.3fF
C1071 diff_3901000_1040000# gnd! 132.6fF
C1072 diff_4056000_1090000# gnd! 287.6fF
C1073 diff_4165000_1308000# gnd! 111.9fF
C1074 diff_4037000_1195000# gnd! 198.2fF
C1075 diff_3901000_1073000# gnd! 282.9fF
C1076 diff_3780000_968000# gnd! 120.1fF
C1077 diff_3686000_934000# gnd! 123.4fF
C1078 diff_3670000_960000# gnd! 123.9fF
C1079 diff_3697000_1029000# gnd! 327.6fF
C1080 diff_3687000_1019000# gnd! 131.1fF
C1081 diff_3937000_1185000# gnd! 193.6fF
C1082 diff_4005000_1296000# gnd! 52.4fF
C1083 diff_4242000_1303000# gnd! 157.4fF
C1084 diff_4275000_1328000# gnd! 68.7fF
C1085 diff_4252000_1283000# gnd! 90.6fF
C1086 diff_4480000_1851000# gnd! 46.6fF
C1087 diff_4726000_1860000# gnd! 259.7fF
C1088 diff_4693000_1939000# gnd! 157.4fF
C1089 diff_4753000_1809000# gnd! 669.6fF
C1090 diff_4798000_1884000# gnd! 112.2fF
C1091 diff_4820000_1904000# gnd! 111.9fF
C1092 diff_4971000_2027000# gnd! 199.9fF
C1093 diff_4982000_2020000# gnd! 91.7fF
C1094 diff_5289000_2222000# gnd! 159.6fF
C1095 diff_5278000_2280000# gnd! 89.2fF
C1096 diff_5201000_2341000# gnd! 325.1fF
C1097 diff_5242000_2359000# gnd! 304.1fF
C1098 diff_5208000_2365000# gnd! 99.1fF
C1099 diff_5070000_2118000# gnd! 224.9fF
C1100 diff_5111000_2140000# gnd! 771.6fF
C1101 diff_5132000_2347000# gnd! 128.3fF
C1102 diff_5068000_2286000# gnd! 63.4fF
C1103 diff_5024000_2111000# gnd! 311.6fF
C1104 diff_4904000_2082000# gnd! 148.7fF
C1105 diff_4869000_2081000# gnd! 404.8fF
C1106 diff_4893000_2186000# gnd! 59.3fF
C1107 diff_5037000_2263000# gnd! 43.8fF
C1108 diff_5124000_2368000# gnd! 592.5fF
C1109 diff_5068000_2348000# gnd! 259.9fF
C1110 diff_5021000_2345000# gnd! 280.0fF
C1111 diff_5151000_2372000# gnd! 108.0fF
C1112 diff_5446000_801000# gnd! 1158.0fF
C1113 diff_5576000_2597000# gnd! 676.1fF
C1114 diff_5650000_2540000# gnd! 634.6fF
C1115 diff_5555000_2636000# gnd! 486.3fF
C1116 diff_5696000_2541000# gnd! 2232.7fF
C1117 diff_5631000_2728000# gnd! 542.9fF
C1118 diff_5652000_2806000# gnd! 247.2fF
C1119 diff_5617000_2717000# gnd! 355.4fF
C1120 diff_5625000_2883000# gnd! 299.4fF
C1121 diff_5768000_2822000# gnd! 2119.7fF
C1122 diff_6212000_3182000# gnd! 310.8fF
C1123 diff_5270000_856000# gnd! 200.1fF
C1124 diff_5200000_2399000# gnd! 211.4fF
C1125 diff_5224000_815000# gnd! 410.1fF
C1126 diff_5387000_2603000# gnd! 248.5fF
C1127 diff_5235000_2513000# gnd! 83.0fF
C1128 diff_5314000_2695000# gnd! 165.6fF
C1129 diff_5300000_2536000# gnd! 547.3fF
C1130 diff_5289000_2527000# gnd! 145.8fF
C1131 diff_5299000_2749000# gnd! 59.1fF
C1132 diff_5074000_2370000# gnd! 96.3fF
C1133 diff_5028000_2372000# gnd! 59.9fF
C1134 diff_4991000_2210000# gnd! 265.8fF
C1135 diff_4971000_2235000# gnd! 198.6fF
C1136 diff_4951000_2235000# gnd! 151.4fF
C1137 diff_4831000_2023000# gnd! 266.9fF
C1138 diff_4701000_1996000# gnd! 211.9fF
C1139 diff_4692000_2057000# gnd! 156.4fF
C1140 diff_4624000_1908000# gnd! 62.4fF
C1141 diff_4563000_1895000# gnd! 45.1fF
C1142 diff_4607000_1846000# gnd! 349.4fF
C1143 diff_4574000_1950000# gnd! 259.0fF
C1144 diff_4588000_1994000# gnd! 174.6fF
C1145 diff_4706000_2104000# gnd! 52.3fF
C1146 diff_4672000_2104000# gnd! 52.4fF
C1147 diff_4519000_1750000# gnd! 327.7fF
C1148 diff_4532000_1851000# gnd! 56.1fF
C1149 diff_4517000_1949000# gnd! 273.8fF
C1150 diff_4460000_1689000# gnd! 274.5fF
C1151 diff_4379000_1770000# gnd! 135.5fF
C1152 diff_4435000_1905000# gnd! 100.0fF
C1153 diff_4531000_1993000# gnd! 90.0fF
C1154 diff_4409000_1887000# gnd! 361.4fF
C1155 diff_4459000_1939000# gnd! 153.2fF
C1156 diff_4379000_1851000# gnd! 134.6fF
C1157 diff_4726000_2137000# gnd! 262.8fF
C1158 diff_4809000_2023000# gnd! 251.0fF
C1159 diff_4787000_2161000# gnd! 210.7fF
C1160 diff_4821000_2015000# gnd! 107.2fF
C1161 diff_4799000_2016000# gnd! 104.0fF
C1162 diff_4893000_2206000# gnd! 59.3fF
C1163 diff_4675000_2150000# gnd! 45.2fF
C1164 diff_4706000_2150000# gnd! 121.0fF
C1165 diff_4866000_2115000# gnd! 358.2fF
C1166 diff_4899000_2195000# gnd! 572.0fF
C1167 diff_4982000_2204000# gnd! 91.7fF
C1168 diff_5186000_2543000# gnd! 219.8fF
C1169 diff_5141000_2519000# gnd! 121.0fF
C1170 diff_5174000_2532000# gnd! 126.8fF
C1171 diff_5156000_2419000# gnd! 183.3fF ;**FLOATING
C1172 diff_5141000_2399000# gnd! 747.6fF
C1173 diff_5163000_2687000# gnd! 64.4fF
C1174 diff_5123000_2494000# gnd! 424.2fF
C1175 diff_4870000_2312000# gnd! 389.8fF
C1176 diff_4904000_2299000# gnd! 143.4fF
C1177 diff_4881000_2375000# gnd! 57.2fF
C1178 diff_4831000_2306000# gnd! 274.4fF
C1179 diff_4809000_2270000# gnd! 252.6fF
C1180 diff_4787000_2229000# gnd! 202.4fF
C1181 diff_4675000_2228000# gnd! 45.2fF
C1182 diff_4563000_2106000# gnd! 47.1fF
C1183 diff_4574000_2030000# gnd! 257.8fF
C1184 diff_4624000_2092000# gnd! 62.6fF
C1185 diff_4607000_2076000# gnd! 348.3fF
C1186 diff_4706000_2228000# gnd! 121.3fF
C1187 diff_4706000_2273000# gnd! 52.1fF
C1188 diff_4672000_2273000# gnd! 54.6fF
C1189 diff_4617000_2117000# gnd! 326.1fF
C1190 diff_4517000_2031000# gnd! 266.4fF
C1191 diff_4532000_2086000# gnd! 55.7fF
C1192 diff_4477000_1873000# gnd! 522.7fF
C1193 diff_4481000_2154000# gnd! 40.8fF
C1194 diff_4432000_2036000# gnd! 230.1fF
C1195 diff_4481000_2228000# gnd! 48.4fF
C1196 diff_4726000_2237000# gnd! 261.0fF
C1197 diff_4693000_2316000# gnd! 157.4fF
C1198 diff_4753000_2186000# gnd! 669.2fF
C1199 diff_4820000_2281000# gnd! 112.3fF
C1200 diff_4798000_2261000# gnd! 113.3fF
C1201 diff_4701000_2373000# gnd! 162.4fF
C1202 diff_4968000_2493000# gnd! 218.7fF
C1203 diff_5074000_2676000# gnd! 404.2fF
C1204 diff_5190000_2733000# gnd! 45.1fF
C1205 diff_5186000_2411000# gnd! 583.5fF
C1206 diff_5200000_2422000# gnd! 847.6fF
C1207 diff_5320000_2718000# gnd! 472.4fF
C1208 diff_5270000_2492000# gnd! 534.4fF
C1209 diff_5113000_2489000# gnd! 214.6fF
C1210 diff_5064000_2665000# gnd! 144.8fF
C1211 diff_5028000_2635000# gnd! 366.4fF
C1212 diff_5034000_2443000# gnd! 170.3fF
C1213 diff_4993000_2633000# gnd! 1144.4fF
C1214 diff_4931000_826000# gnd! 1775.0fF
C1215 diff_4971000_2631000# gnd! 188.9fF
C1216 diff_5317000_2777000# gnd! 301.9fF
C1217 diff_5264000_2777000# gnd! 262.0fF
C1218 diff_5257000_2805000# gnd! 88.8fF
C1219 diff_5085000_2690000# gnd! 99.7fF
C1220 diff_5052000_2756000# gnd! 37.4fF
C1221 diff_5013000_2754000# gnd! 257.0fF
C1222 diff_4958000_2607000# gnd! 339.4fF
C1223 diff_4991000_2691000# gnd! 61.5fF
C1224 diff_5171000_2829000# gnd! 312.6fF
C1225 diff_4996000_2788000# gnd! 62.3fF
C1226 diff_4944000_2493000# gnd! 669.9fF
C1227 diff_4624000_2286000# gnd! 61.2fF
C1228 diff_4563000_2272000# gnd! 45.2fF
C1229 diff_4607000_2223000# gnd! 352.0fF
C1230 diff_4574000_2327000# gnd! 258.5fF
C1231 diff_4588000_2371000# gnd! 132.0fF
C1232 diff_4519000_2127000# gnd! 328.7fF
C1233 diff_4532000_2229000# gnd! 55.1fF
C1234 diff_4517000_2326000# gnd! 273.6fF
C1235 diff_4460000_2077000# gnd! 250.7fF
C1236 diff_4410000_2197000# gnd! 123.8fF
C1237 diff_4531000_2370000# gnd! 52.4fF
C1238 diff_4478000_2251000# gnd! 270.8fF
C1239 diff_4905000_2664000# gnd! 1299.2fF
C1240 diff_4896000_2688000# gnd! 84.0fF
C1241 diff_4838000_2617000# gnd! 1402.5fF
C1242 diff_4819000_2721000# gnd! 232.4fF
C1243 diff_4882000_2652000# gnd! 303.1fF
C1244 diff_4804000_2758000# gnd! 367.3fF
C1245 diff_4837000_2673000# gnd! 322.4fF
C1246 diff_4777000_2518000# gnd! 540.0fF
C1247 diff_4739000_2640000# gnd! 1108.9fF
C1248 diff_4718000_2635000# gnd! 209.5fF
C1249 diff_4761000_2747000# gnd! 266.0fF
C1250 diff_4704000_2610000# gnd! 392.9fF
C1251 diff_4741000_2690000# gnd! 62.8fF
C1252 diff_4675000_2475000# gnd! 717.3fF
C1253 diff_4434000_2245000# gnd! 112.5fF
C1254 diff_4379000_2146000# gnd! 127.7fF
C1255 diff_4380000_2279000# gnd! 130.5fF
C1256 diff_4354000_1418000# gnd! 1266.4fF
C1257 diff_4267000_1478000# gnd! 282.4fF
C1258 diff_4306000_1553000# gnd! 204.6fF
C1259 diff_4267000_1500000# gnd! 104.6fF
C1260 diff_4245000_1443000# gnd! 865.7fF
C1261 diff_4184000_1383000# gnd! 189.9fF
C1262 diff_4204000_1414000# gnd! 422.8fF
C1263 diff_4149000_1346000# gnd! 134.2fF
C1264 diff_4057000_1357000# gnd! 119.4fF
C1265 diff_4037000_1296000# gnd! 195.4fF
C1266 diff_4067000_1406000# gnd! 337.6fF
C1267 diff_4056000_1396000# gnd! 132.4fF
C1268 diff_4226000_1550000# gnd! 162.6fF
C1269 diff_4287000_1631000# gnd! 70.0fF
C1270 diff_4286000_1500000# gnd! 291.2fF
C1271 diff_4232000_1627000# gnd! 45.9fF
C1272 diff_4274000_1612000# gnd! 268.9fF
C1273 diff_4319000_1315000# gnd! 206.6fF
C1274 diff_4347000_2438000# gnd! 889.8fF
C1275 diff_4185000_1452000# gnd! 180.2fF
C1276 diff_4166000_1562000# gnd! 113.1fF
C1277 diff_4067000_1476000# gnd! 403.0fF
C1278 diff_3949000_1339000# gnd! 130.2fF
C1279 diff_3847000_1127000# gnd! 523.3fF
C1280 diff_3938000_1304000# gnd! 188.5fF
C1281 diff_3881000_1306000# gnd! 326.3fF
C1282 diff_3847000_1324000# gnd! 144.1fF
C1283 diff_3819000_1288000# gnd! 150.7fF
C1284 diff_3697000_1099000# gnd! 510.5fF
C1285 diff_3632000_946000# gnd! 99.2fF
C1286 diff_3610000_906000# gnd! 162.5fF
C1287 diff_3557000_956000# gnd! 130.7fF
C1288 diff_3538000_920000# gnd! 113.8fF
C1289 diff_3499000_875000# gnd! 65.3fF
C1290 diff_3424000_872000# gnd! 52.5fF
C1291 diff_3422000_893000# gnd! 202.7fF
C1292 diff_3397000_928000# gnd! 45.6fF
C1293 diff_3578000_992000# gnd! 179.5fF
C1294 diff_3685000_1184000# gnd! 290.4fF
C1295 diff_3633000_1168000# gnd! 241.8fF
C1296 diff_3659000_1285000# gnd! 51.6fF
C1297 diff_3520000_968000# gnd! 121.4fF
C1298 diff_3427000_934000# gnd! 115.8fF
C1299 diff_3409000_959000# gnd! 116.3fF
C1300 diff_3437000_1029000# gnd! 328.5fF
C1301 diff_3427000_1018000# gnd! 133.7fF
C1302 diff_3323000_873000# gnd! 232.9fF
C1303 diff_3373000_928000# gnd! 178.0fF
C1304 diff_3334000_1004000# gnd! 92.6fF
C1305 diff_3578000_1133000# gnd! 586.8fF
C1306 diff_3795000_1343000# gnd! 124.0fF
C1307 diff_3864000_1391000# gnd! 110.3fF
C1308 diff_3901000_1417000# gnd! 132.5fF
C1309 diff_3780000_1346000# gnd! 119.1fF
C1310 diff_3686000_1310000# gnd! 128.9fF
C1311 diff_3670000_1337000# gnd! 122.2fF
C1312 diff_3697000_1406000# gnd! 325.3fF
C1313 diff_3687000_1396000# gnd! 131.1fF
C1314 diff_4056000_1466000# gnd! 289.1fF
C1315 diff_4225000_1648000# gnd! 478.4fF
C1316 diff_4239000_1722000# gnd! 64.0fF
C1317 diff_4165000_1685000# gnd! 111.9fF
C1318 diff_4038000_1572000# gnd! 195.0fF
C1319 diff_3901000_1450000# gnd! 284.4fF
C1320 diff_3937000_1562000# gnd! 190.3fF
C1321 diff_4005000_1673000# gnd! 52.4fF
C1322 diff_4184000_1760000# gnd! 189.9fF
C1323 diff_4251000_1918000# gnd! 69.8fF
C1324 diff_4235000_1746000# gnd! 299.6fF
C1325 diff_4204000_1790000# gnd! 350.4fF
C1326 diff_4149000_1723000# gnd! 135.0fF
C1327 diff_4057000_1734000# gnd! 118.7fF
C1328 diff_4038000_1673000# gnd! 194.4fF
C1329 diff_4067000_1784000# gnd! 338.7fF
C1330 diff_4056000_1773000# gnd! 134.1fF
C1331 diff_4264000_1839000# gnd! 840.7fF
C1332 diff_4617000_2492000# gnd! 138.3fF
C1333 diff_4825000_2753000# gnd! 157.9fF
C1334 diff_4784000_2782000# gnd! 320.1fF
C1335 diff_4580000_2552000# gnd! 48.8fF
C1336 diff_4528000_2536000# gnd! 22.2fF
C1337 diff_4517000_2527000# gnd! 265.0fF
C1338 diff_4528000_2748000# gnd! 52.4fF
C1339 diff_4477000_2552000# gnd! 54.6fF
C1340 diff_4425000_2536000# gnd! 5.0fF
C1341 diff_4414000_2527000# gnd! 276.4fF
C1342 diff_4424000_2748000# gnd! 54.6fF
C1343 diff_4642000_2735000# gnd! 294.8fF
C1344 diff_4623000_2773000# gnd! 57.8fF
C1345 diff_4547000_2724000# gnd! 1504.6fF
C1346 diff_4497000_2491000# gnd! 1588.6fF
C1347 diff_4416000_951000# gnd! 1479.7fF
C1348 diff_4373000_832000# gnd! 1605.0fF
C1349 diff_4601000_2751000# gnd! 1791.8fF
C1350 diff_4545000_2777000# gnd! 267.6fF
C1351 diff_4493000_2777000# gnd! 256.0fF
C1352 diff_4442000_2777000# gnd! 265.4fF
C1353 diff_4390000_2777000# gnd! 262.6fF
C1354 diff_4688000_2591000# gnd! 309.4fF
C1355 diff_4931000_2481000# gnd! 202.5fF
C1356 diff_4734000_2812000# gnd! 50.9fF
C1357 diff_4382000_2804000# gnd! 181.8fF
C1358 diff_5203000_3036000# gnd! 774.3fF
C1359 diff_5213000_3049000# gnd! 451.6fF
C1360 diff_6251000_3156000# gnd! 687.5fF
C1361 diff_6268000_3283000# gnd! 134.6fF
C1362 diff_6268000_3301000# gnd! 121.1fF
C1363 diff_5011000_3005000# gnd! 119.3fF
C1364 diff_4911000_2899000# gnd! 308.4fF
C1365 diff_4974000_2909000# gnd! 287.7fF
C1366 diff_5018000_2992000# gnd! 160.5fF
C1367 diff_5575000_3240000# gnd! 115.5fF
C1368 diff_5083000_3005000# gnd! 191.1fF
C1369 diff_5468000_3308000# gnd! 121.8fF
C1370 diff_6179000_3355000# gnd! 410.6fF
C1371 diff_6121000_3398000# gnd! 222.6fF
C1372 diff_5530000_3345000# gnd! 101.7fF
C1373 diff_5406000_3339000# gnd! 196.4fF
C1374 diff_6005000_3448000# gnd! 79.7fF
C1375 diff_6159000_3458000# gnd! 86.0fF
C1376 diff_4967000_3078000# gnd! 121.1fF
C1377 diff_4984000_2921000# gnd! 798.5fF
C1378 diff_4904000_3016000# gnd! 233.1fF
C1379 diff_4922000_2910000# gnd! 257.6fF
C1380 diff_4842000_3066000# gnd! 856.8fF
C1381 diff_4864000_3204000# gnd! 111.6fF
C1382 diff_4842000_3180000# gnd! 128.1fF
C1383 diff_4776000_2950000# gnd! 555.3fF
C1384 diff_4185000_1829000# gnd! 181.1fF
C1385 diff_4166000_1940000# gnd! 113.3fF
C1386 diff_4067000_1854000# gnd! 405.2fF
C1387 diff_3949000_1717000# gnd! 129.2fF
C1388 diff_3847000_1503000# gnd! 517.2fF
C1389 diff_3938000_1681000# gnd! 187.7fF
C1390 diff_3881000_1684000# gnd! 327.5fF
C1391 diff_3847000_1701000# gnd! 144.1fF
C1392 diff_3819000_1665000# gnd! 152.1fF
C1393 diff_3697000_1476000# gnd! 501.6fF
C1394 diff_3633000_1323000# gnd! 96.9fF
C1395 diff_3610000_1283000# gnd! 164.9fF
C1396 diff_3557000_1333000# gnd! 132.6fF
C1397 diff_3538000_1297000# gnd! 117.8fF
C1398 diff_3437000_1100000# gnd! 506.3fF
C1399 diff_3426000_1188000# gnd! 280.5fF
C1400 diff_3373000_1152000# gnd! 318.5fF
C1401 diff_3183000_765000# gnd! 164.6fF
C1402 diff_2598000_626000# gnd! 162.8fF
C1403 diff_3171000_743000# gnd! 146.8fF
C1404 diff_3065000_767000# gnd! 164.6fF
C1405 diff_2970000_767000# gnd! 172.1fF
C1406 diff_2838000_765000# gnd! 162.4fF
C1407 diff_2744000_764000# gnd! 164.6fF
C1408 diff_3054000_743000# gnd! 142.6fF
C1409 diff_3181000_876000# gnd! 61.3fF
C1410 diff_3091000_870000# gnd! 57.9fF
C1411 diff_3092000_894000# gnd! 239.4fF
C1412 diff_3244000_742000# gnd! 193.2fF ;**FLOATING
C1413 diff_3238000_927000# gnd! 177.6fF
C1414 diff_3212000_963000# gnd! 121.4fF
C1415 diff_3196000_965000# gnd! 152.6fF
C1416 diff_2959000_743000# gnd! 138.6fF
C1417 diff_3052000_908000# gnd! 51.9fF
C1418 diff_3098000_928000# gnd! 124.2fF
C1419 diff_3092000_955000# gnd! 115.0fF
C1420 diff_3118000_1024000# gnd! 323.4fF
C1421 diff_3108000_1012000# gnd! 140.6fF
C1422 diff_3062000_965000# gnd! 142.5fF
C1423 diff_3397000_1305000# gnd! 45.6fF
C1424 diff_3578000_1369000# gnd! 179.5fF
C1425 diff_3685000_1561000# gnd! 293.8fF
C1426 diff_3633000_1545000# gnd! 241.6fF
C1427 diff_3659000_1662000# gnd! 49.4fF
C1428 diff_3520000_1345000# gnd! 120.8fF
C1429 diff_3427000_1308000# gnd! 117.0fF
C1430 diff_3409000_1334000# gnd! 117.0fF
C1431 diff_3437000_1406000# gnd! 319.3fF
C1432 diff_3427000_1395000# gnd! 133.7fF
C1433 diff_3373000_1305000# gnd! 176.3fF
C1434 diff_3334000_1381000# gnd! 92.6fF
C1435 diff_3118000_1088000# gnd! 493.8fF
C1436 diff_3081000_1137000# gnd! 809.8fF
C1437 diff_3098000_1188000# gnd! 297.4fF
C1438 diff_2827000_743000# gnd! 137.4fF
C1439 diff_2937000_871000# gnd! 56.7fF
C1440 diff_2962000_909000# gnd! 45.6fF
C1441 diff_2860000_876000# gnd! 64.3fF
C1442 diff_2860000_903000# gnd! 217.2fF
C1443 diff_3011000_980000# gnd! 47.9fF
C1444 diff_2987000_946000# gnd! 142.2fF
C1445 diff_3028000_909000# gnd! 191.8fF
C1446 diff_3005000_1018000# gnd! 43.3fF
C1447 diff_3256000_1245000# gnd! 648.9fF
C1448 diff_3212000_1340000# gnd! 144.9fF
C1449 diff_3578000_1510000# gnd! 586.1fF
C1450 diff_3795000_1720000# gnd! 130.4fF
C1451 diff_3864000_1769000# gnd! 109.4fF
C1452 diff_3901000_1794000# gnd! 134.3fF
C1453 diff_3780000_1723000# gnd! 118.4fF
C1454 diff_3686000_1688000# gnd! 128.5fF
C1455 diff_3670000_1715000# gnd! 122.1fF
C1456 diff_3697000_1784000# gnd! 325.5fF
C1457 diff_3687000_1773000# gnd! 132.8fF
C1458 diff_4056000_1844000# gnd! 290.7fF
C1459 diff_4225000_1879000# gnd! 154.9fF
C1460 diff_4165000_2061000# gnd! 110.8fF
C1461 diff_4037000_1949000# gnd! 197.6fF
C1462 diff_3901000_1828000# gnd! 286.9fF
C1463 diff_3937000_1939000# gnd! 193.0fF
C1464 diff_4005000_2050000# gnd! 52.4fF
C1465 diff_4184000_2136000# gnd! 187.7fF
C1466 diff_4204000_2168000# gnd! 352.2fF
C1467 diff_4150000_2101000# gnd! 125.2fF
C1468 diff_4057000_2112000# gnd! 116.9fF
C1469 diff_4037000_2050000# gnd! 195.2fF
C1470 diff_4067000_2161000# gnd! 337.6fF
C1471 diff_4056000_2150000# gnd! 134.1fF
C1472 diff_4237000_2412000# gnd! 40.9fF
C1473 diff_4185000_2206000# gnd! 193.7fF
C1474 diff_4166000_2316000# gnd! 112.4fF
C1475 diff_4067000_2231000# gnd! 387.9fF
C1476 diff_3949000_2094000# gnd! 127.4fF
C1477 diff_3847000_1880000# gnd! 519.2fF
C1478 diff_3938000_2059000# gnd! 188.3fF
C1479 diff_3881000_2061000# gnd! 325.2fF
C1480 diff_3847000_2079000# gnd! 144.4fF
C1481 diff_3819000_2042000# gnd! 153.4fF
C1482 diff_3697000_1854000# gnd! 508.9fF
C1483 diff_3633000_1700000# gnd! 96.8fF
C1484 diff_3610000_1660000# gnd! 164.1fF
C1485 diff_3557000_1710000# gnd! 127.6fF
C1486 diff_3538000_1674000# gnd! 117.7fF
C1487 diff_3437000_1477000# gnd! 491.7fF
C1488 diff_3426000_1565000# gnd! 282.3fF
C1489 diff_3373000_1529000# gnd! 320.0fF
C1490 diff_3196000_1342000# gnd! 151.1fF
C1491 diff_3028000_1167000# gnd! 345.3fF
C1492 diff_3051000_1286000# gnd! 52.4fF
C1493 diff_3098000_1305000# gnd! 120.3fF
C1494 diff_3092000_1332000# gnd! 109.2fF
C1495 diff_3118000_1401000# gnd! 329.4fF
C1496 diff_3108000_1389000# gnd! 138.8fF
C1497 diff_3062000_1342000# gnd! 145.5fF
C1498 diff_3397000_1682000# gnd! 47.6fF
C1499 diff_3578000_1747000# gnd! 178.4fF
C1500 diff_3685000_1939000# gnd! 294.7fF
C1501 diff_3633000_1922000# gnd! 241.9fF
C1502 diff_3659000_2040000# gnd! 49.3fF
C1503 diff_3520000_1723000# gnd! 121.4fF
C1504 diff_3427000_1686000# gnd! 119.5fF
C1505 diff_3409000_1711000# gnd! 119.7fF
C1506 diff_3437000_1784000# gnd! 319.4fF
C1507 diff_3427000_1773000# gnd! 131.9fF
C1508 diff_3373000_1682000# gnd! 176.2fF
C1509 diff_3334000_1758000# gnd! 94.3fF
C1510 diff_3578000_1887000# gnd! 719.0fF
C1511 diff_3795000_2097000# gnd! 123.5fF
C1512 diff_3864000_2146000# gnd! 108.4fF
C1513 diff_3901000_2171000# gnd! 134.2fF
C1514 diff_4056000_2221000# gnd! 290.5fF
C1515 diff_4192000_1025000# gnd! 947.9fF
C1516 diff_4038000_2326000# gnd! 198.1fF
C1517 diff_3901000_2205000# gnd! 288.1fF
C1518 diff_3780000_2100000# gnd! 118.4fF
C1519 diff_3686000_2065000# gnd! 127.0fF
C1520 diff_3670000_2092000# gnd! 119.5fF
C1521 diff_3697000_2161000# gnd! 321.9fF
C1522 diff_3687000_2150000# gnd! 132.8fF
C1523 diff_3937000_2316000# gnd! 190.8fF
C1524 diff_4162000_2432000# gnd! 1170.0fF
C1525 diff_4292000_2626000# gnd! 98.8fF
C1526 diff_4240000_2606000# gnd! 88.3fF
C1527 diff_4307000_2532000# gnd! 357.7fF
C1528 diff_3847000_2257000# gnd! 516.0fF
C1529 diff_3697000_2231000# gnd! 503.2fF
C1530 diff_3633000_2077000# gnd! 95.1fF
C1531 diff_3610000_2037000# gnd! 162.6fF
C1532 diff_3557000_2087000# gnd! 133.6fF
C1533 diff_3538000_2051000# gnd! 118.7fF
C1534 diff_3437000_1855000# gnd! 497.4fF
C1535 diff_3426000_1943000# gnd! 284.0fF
C1536 diff_3373000_1906000# gnd! 319.7fF
C1537 diff_3397000_2059000# gnd! 45.6fF
C1538 diff_3578000_2124000# gnd! 178.6fF
C1539 diff_3685000_2316000# gnd! 296.3fF
C1540 diff_3633000_2300000# gnd! 241.6fF
C1541 diff_3801000_831000# gnd! 1133.8fF
C1542 diff_4192000_2538000# gnd! 180.7fF
C1543 diff_4154000_2620000# gnd! 73.5fF
C1544 diff_4154000_2675000# gnd! 679.0fF
C1545 diff_4251000_2644000# gnd! 482.9fF
C1546 diff_4266000_2739000# gnd! 94.0fF
C1547 diff_4276000_2780000# gnd! 699.1fF
C1548 diff_4223000_2738000# gnd! 695.5fF
C1549 diff_4213000_2744000# gnd! 65.4fF
C1550 diff_4161000_2693000# gnd! 101.1fF
C1551 diff_4138000_2552000# gnd! 456.7fF
C1552 diff_4086000_2536000# gnd! 24.9fF
C1553 diff_4076000_2526000# gnd! 254.8fF
C1554 diff_4086000_2748000# gnd! 52.4fF
C1555 diff_4035000_2552000# gnd! 48.5fF
C1556 diff_3983000_2536000# gnd! 24.9fF
C1557 diff_3521000_2100000# gnd! 111.6fF
C1558 diff_3427000_2063000# gnd! 117.9fF
C1559 diff_3409000_2088000# gnd! 118.2fF
C1560 diff_3437000_2161000# gnd! 326.0fF
C1561 diff_3427000_2150000# gnd! 131.9fF
C1562 diff_3373000_2059000# gnd! 175.8fF
C1563 diff_3334000_2135000# gnd! 94.1fF
C1564 diff_3578000_2264000# gnd! 739.2fF
C1565 diff_3437000_2232000# gnd! 502.4fF
C1566 diff_3373000_2283000# gnd! 319.4fF
C1567 diff_3426000_2320000# gnd! 284.5fF
C1568 diff_3973000_2526000# gnd! 254.8fF
C1569 diff_3983000_2748000# gnd! 52.4fF
C1570 diff_3932000_2552000# gnd! 57.1fF
C1571 diff_3880000_2536000# gnd! 25.1fF
C1572 diff_3870000_2526000# gnd! 254.8fF
C1573 diff_3880000_2748000# gnd! 52.4fF
C1574 diff_3829000_2552000# gnd! 57.1fF
C1575 diff_3777000_2536000# gnd! 22.2fF
C1576 diff_3766000_2527000# gnd! 265.0fF
C1577 diff_3777000_2748000# gnd! 52.4fF
C1578 diff_3726000_2552000# gnd! 46.3fF
C1579 diff_3674000_2536000# gnd! 24.9fF
C1580 diff_3664000_2526000# gnd! 254.8fF
C1581 diff_3674000_2748000# gnd! 52.4fF
C1582 diff_3622000_2553000# gnd! 70.1fF
C1583 diff_3571000_2536000# gnd! 22.1fF
C1584 diff_3560000_2527000# gnd! 266.6fF
C1585 diff_3570000_2748000# gnd! 54.6fF
C1586 diff_3519000_2552000# gnd! 70.2fF
C1587 diff_3467000_2537000# gnd! 22.1fF
C1588 diff_3118000_1465000# gnd! 487.8fF
C1589 diff_3081000_1341000# gnd! 795.7fF
C1590 diff_3098000_1565000# gnd! 299.2fF
C1591 diff_2733000_743000# gnd! 137.4fF
C1592 diff_2680000_788000# gnd! 179.5fF
C1593 diff_2590000_764000# gnd! 151.6fF
C1594 diff_2228000_597000# gnd! 169.6fF
C1595 diff_1757000_612000# gnd! 470.6fF
C1596 diff_1757000_699000# gnd! 50.5fF
C1597 diff_1703000_589000# gnd! 252.9fF
C1598 diff_1693000_584000# gnd! 2765.2fF
C1599 diff_1490000_540000# gnd! 77.6fF
C1600 diff_1398000_490000# gnd! 153.3fF
C1601 diff_1345000_491000# gnd! 153.6fF
C1602 diff_1292000_491000# gnd! 156.8fF
C1603 diff_701000_124000# gnd! 20.3fF
C1604 diff_691000_114000# gnd! 280.8fF
C1605 diff_708000_309000# gnd! 101.8fF
C1606 diff_459000_154000# gnd! 68.9fF
C1607 diff_183000_100000# gnd! 870.7fF
C1608 diff_598000_271000# gnd! 63.8fF
C1609 diff_639000_113000# gnd! 232.0fF
C1610 diff_457000_301000# gnd! 534.8fF
C1611 diff_458000_352000# gnd! 230.6fF
C1612 diff_173000_152000# gnd! 2310.2fF
C1613 diff_458000_404000# gnd! 230.5fF
C1614 diff_1134000_464000# gnd! 158.2fF
C1615 diff_1082000_465000# gnd! 156.0fF
C1616 diff_1049000_100000# gnd! 2439.1fF
C1617 diff_1219000_196000# gnd! 3672.6fF
C1618 diff_1429000_544000# gnd! 233.1fF
C1619 diff_1503000_592000# gnd! 245.3fF
C1620 diff_1619000_122000# gnd! 2100.9fF
C1621 diff_1641000_566000# gnd! 389.2fF
C1622 diff_1631000_556000# gnd! 219.8fF
C1623 diff_1547000_715000# gnd! 375.0fF
C1624 diff_1429000_566000# gnd! 2120.2fF
C1625 diff_1405000_650000# gnd! 282.0fF
C1626 diff_1371000_619000# gnd! 54.2fF
C1627 diff_1360000_692000# gnd! 59.0fF
C1628 diff_1452000_699000# gnd! 55.2fF
C1629 diff_1384000_624000# gnd! 484.2fF
C1630 diff_1537000_704000# gnd! 218.9fF
C1631 diff_1286000_578000# gnd! 323.0fF
C1632 diff_1276000_567000# gnd! 362.0fF
C1633 diff_1228000_660000# gnd! 363.6fF
C1634 diff_1218000_655000# gnd! 256.6fF
C1635 diff_1203000_545000# gnd! 2739.2fF
C1636 diff_928000_464000# gnd! 183.6fF
C1637 diff_876000_465000# gnd! 175.5fF
C1638 diff_588000_420000# gnd! 240.6fF
C1639 diff_802000_365000# gnd! 3522.6fF
C1640 diff_597000_373000# gnd! 2206.8fF
C1641 diff_136000_354000# gnd! 2210.7fF
C1642 diff_125000_346000# gnd! 2221.8fF
C1643 diff_968000_455000# gnd! 2178.2fF
C1644 diff_980000_464000# gnd! 467.0fF
C1645 diff_1115000_636000# gnd! 229.5fF
C1646 diff_2930000_970000# gnd! 111.7fF
C1647 diff_2914000_928000# gnd! 104.0fF
C1648 diff_2875000_1038000# gnd! 143.2fF
C1649 diff_2865000_1028000# gnd! 339.6fF
C1650 diff_2846000_994000# gnd! 124.7fF
C1651 diff_2830000_938000# gnd! 131.1fF
C1652 diff_2658000_766000# gnd! 66.0fF
C1653 diff_2744000_876000# gnd! 63.5fF
C1654 diff_2668000_869000# gnd! 57.2fF
C1655 diff_2667000_894000# gnd! 218.3fF
C1656 diff_2597000_842000# gnd! 78.5fF
C1657 diff_2799000_944000# gnd! 176.7fF
C1658 diff_2781000_945000# gnd! 134.4fF
C1659 diff_2628000_910000# gnd! 120.0fF
C1660 diff_2759000_1004000# gnd! 147.6fF
C1661 diff_2674000_928000# gnd! 116.0fF
C1662 diff_2651000_946000# gnd! 154.7fF
C1663 diff_2468000_786000# gnd! 166.6fF
C1664 diff_2476000_759000# gnd! 74.5fF
C1665 diff_2338000_781000# gnd! 200.9fF
C1666 diff_2365000_781000# gnd! 298.3fF
C1667 diff_2342000_760000# gnd! 80.0fF
C1668 diff_2408000_867000# gnd! 206.5fF
C1669 diff_2684000_1023000# gnd! 325.7fF
C1670 diff_2673000_1012000# gnd! 147.7fF
C1671 diff_2886000_1048000# gnd! 821.0fF
C1672 diff_2875000_1073000# gnd! 290.5fF
C1673 diff_2914000_1187000# gnd! 274.5fF
C1674 diff_2759000_1078000# gnd! 1380.0fF
C1675 diff_2628000_975000# gnd! 120.2fF
C1676 diff_2218000_809000# gnd! 137.1fF
C1677 diff_2117000_758000# gnd! 159.2fF
C1678 diff_2199000_774000# gnd! 106.2fF
C1679 diff_2103000_843000# gnd! 71.3fF
C1680 diff_2027000_787000# gnd! 165.3fF
C1681 diff_1888000_764000# gnd! 169.8fF
C1682 diff_1876000_750000# gnd! 199.9fF
C1683 diff_1978000_775000# gnd! 161.1fF
C1684 diff_2103000_883000# gnd! 16.4fF
C1685 diff_2197000_895000# gnd! 431.9fF
C1686 diff_2500000_969000# gnd! 51.4fF
C1687 diff_2550000_879000# gnd! 626.7fF
C1688 diff_2532000_968000# gnd! 254.8fF
C1689 diff_2830000_1110000# gnd! 511.5fF
C1690 diff_2962000_1286000# gnd! 43.3fF
C1691 diff_3011000_1357000# gnd! 47.9fF
C1692 diff_2987000_1323000# gnd! 137.0fF
C1693 diff_3028000_1286000# gnd! 189.6fF
C1694 diff_3005000_1395000# gnd! 43.3fF
C1695 diff_3238000_1681000# gnd! 696.0fF
C1696 diff_3212000_1716000# gnd! 144.7fF
C1697 diff_3197000_1718000# gnd! 143.5fF
C1698 diff_3028000_1545000# gnd! 347.8fF
C1699 diff_3052000_1663000# gnd! 50.0fF
C1700 diff_3098000_1682000# gnd! 120.4fF
C1701 diff_3092000_1709000# gnd! 110.0fF
C1702 diff_3118000_1778000# gnd! 330.6fF
C1703 diff_3108000_1767000# gnd! 138.3fF
C1704 diff_3062000_1718000# gnd! 141.5fF
C1705 diff_3118000_1842000# gnd! 491.7fF
C1706 diff_3081000_1718000# gnd! 812.3fF
C1707 diff_3098000_1942000# gnd! 297.0fF
C1708 diff_2930000_1346000# gnd! 111.8fF
C1709 diff_2913000_1305000# gnd! 111.5fF
C1710 diff_2875000_1415000# gnd! 143.3fF
C1711 diff_2865000_1406000# gnd! 339.3fF
C1712 diff_2846000_1371000# gnd! 129.2fF
C1713 diff_2830000_1315000# gnd! 131.1fF
C1714 diff_2655000_1026000# gnd! 640.3fF
C1715 diff_2628000_1087000# gnd! 113.9fF
C1716 diff_2544000_983000# gnd! 197.8fF
C1717 diff_2554000_993000# gnd! 290.0fF
C1718 diff_2384000_972000# gnd! 277.7fF
C1719 diff_2408000_957000# gnd! 60.5fF
C1720 diff_2544000_1075000# gnd! 193.4fF
C1721 diff_2684000_1085000# gnd! 501.0fF
C1722 diff_2652000_1167000# gnd! 157.8fF
C1723 diff_2673000_1076000# gnd! 298.1fF
C1724 diff_2532000_1101000# gnd! 244.8fF
C1725 diff_2628000_1167000# gnd! 128.2fF
C1726 diff_2800000_1321000# gnd! 179.5fF
C1727 diff_2781000_1321000# gnd! 129.6fF
C1728 diff_2628000_1287000# gnd! 121.2fF
C1729 diff_2470000_1073000# gnd! 171.1fF
C1730 diff_2461000_1078000# gnd! 177.3fF
C1731 diff_2341000_1052000# gnd! 1019.7fF
C1732 diff_2382000_1160000# gnd! 99.6fF
C1733 diff_2405000_1193000# gnd! 158.9fF
C1734 diff_2334000_1126000# gnd! 64.4fF
C1735 diff_2292000_953000# gnd! 391.2fF
C1736 diff_2487000_1208000# gnd! 223.7fF
C1737 diff_2475000_1238000# gnd! 160.2fF
C1738 diff_2409000_1226000# gnd! 285.5fF
C1739 diff_2415000_1250000# gnd! 90.1fF
C1740 diff_2759000_1380000# gnd! 148.2fF
C1741 diff_2674000_1305000# gnd! 114.7fF
C1742 diff_2651000_1322000# gnd! 157.9fF
C1743 diff_2684000_1401000# gnd! 311.4fF
C1744 diff_2673000_1390000# gnd! 150.5fF
C1745 diff_2886000_1425000# gnd! 822.0fF
C1746 diff_2875000_1450000# gnd! 290.5fF
C1747 diff_2914000_1564000# gnd! 277.4fF
C1748 diff_2759000_1455000# gnd! 1200.2fF
C1749 diff_2628000_1352000# gnd! 119.1fF
C1750 diff_2549000_1201000# gnd! 352.1fF
C1751 diff_2289000_1090000# gnd! 308.4fF
C1752 diff_2328000_1245000# gnd! 58.4fF
C1753 diff_2532000_1388000# gnd! 242.1fF
C1754 diff_2655000_1403000# gnd! 646.8fF
C1755 diff_2628000_1463000# gnd! 113.9fF
C1756 diff_2544000_1361000# gnd! 196.1fF
C1757 diff_2554000_1371000# gnd! 290.1fF
C1758 diff_2460000_1349000# gnd! 185.8fF
C1759 diff_2405000_1314000# gnd! 159.1fF
C1760 diff_2334000_1371000# gnd! 402.9fF
C1761 diff_2183000_925000# gnd! 286.5fF
C1762 diff_2122000_883000# gnd! 405.8fF
C1763 diff_2129000_912000# gnd! 96.5fF
C1764 diff_2232000_994000# gnd! 58.4fF
C1765 diff_2206000_953000# gnd! 55.0fF
C1766 diff_2136000_921000# gnd! 210.1fF
C1767 diff_2126000_951000# gnd! 87.1fF
C1768 diff_2232000_1087000# gnd! 57.9fF
C1769 diff_2122000_972000# gnd! 666.9fF
C1770 diff_2206000_1163000# gnd! 55.2fF
C1771 diff_2126000_1168000# gnd! 92.4fF
C1772 diff_2183000_1117000# gnd! 289.1fF
C1773 diff_2136000_1203000# gnd! 203.7fF
C1774 diff_2272000_1244000# gnd! 58.7fF
C1775 diff_2129000_1218000# gnd! 97.0fF
C1776 diff_2009000_876000# gnd! 61.2fF
C1777 diff_1965000_869000# gnd! 61.9fF
C1778 diff_1891000_876000# gnd! 68.3fF
C1779 diff_1891000_905000# gnd! 210.8fF
C1780 diff_1981000_947000# gnd! 45.6fF
C1781 diff_2052000_969000# gnd! 158.7fF
C1782 diff_2049000_1016000# gnd! 169.4fF
C1783 diff_2015000_1008000# gnd! 147.4fF
C1784 diff_1996000_984000# gnd! 266.2fF
C1785 diff_2035000_1052000# gnd! 543.7fF
C1786 diff_2052000_1147000# gnd! 154.1fF
C1787 diff_2015000_1090000# gnd! 158.9fF
C1788 diff_1943000_969000# gnd! 144.0fF
C1789 diff_1930000_948000# gnd! 116.0fF
C1790 diff_1851000_942000# gnd! 128.7fF
C1791 diff_1833000_905000# gnd! 113.9fF
C1792 diff_1869000_1028000# gnd! 336.0fF
C1793 diff_1850000_998000# gnd! 121.1fF
C1794 diff_1880000_1040000# gnd! 129.9fF
C1795 diff_1889000_1051000# gnd! 833.1fF
C1796 diff_2103000_1229000# gnd! 17.1fF
C1797 diff_2049000_1080000# gnd! 166.9fF
C1798 diff_2122000_1229000# gnd! 390.5fF
C1799 diff_2271000_1166000# gnd! 468.0fF
C1800 diff_2289000_1293000# gnd! 332.7fF
C1801 diff_2470000_1357000# gnd! 171.3fF
C1802 diff_2544000_1452000# gnd! 193.9fF
C1803 diff_2830000_1487000# gnd! 511.5fF
C1804 diff_2962000_1663000# gnd! 47.6fF
C1805 diff_3011000_1734000# gnd! 50.0fF
C1806 diff_2987000_1700000# gnd! 138.5fF
C1807 diff_3028000_1663000# gnd! 189.6fF
C1808 diff_3005000_1772000# gnd! 43.3fF
C1809 diff_3212000_2093000# gnd! 144.9fF
C1810 diff_3197000_2095000# gnd! 143.6fF
C1811 diff_3028000_1922000# gnd! 347.9fF
C1812 diff_3052000_2040000# gnd! 50.0fF
C1813 diff_3098000_2060000# gnd! 117.5fF
C1814 diff_3092000_2085000# gnd! 109.3fF
C1815 diff_3118000_2155000# gnd! 321.0fF
C1816 diff_3108000_2143000# gnd! 140.5fF
C1817 diff_3062000_2095000# gnd! 141.5fF
C1818 diff_3118000_2218000# gnd! 490.0fF
C1819 diff_3081000_2267000# gnd! 808.6fF
C1820 diff_3098000_2318000# gnd! 295.4fF
C1821 diff_2930000_1723000# gnd! 113.7fF
C1822 diff_2913000_1682000# gnd! 111.1fF
C1823 diff_2865000_1783000# gnd! 342.3fF
C1824 diff_2846000_1747000# gnd! 123.6fF
C1825 diff_2830000_1692000# gnd! 131.1fF
C1826 diff_2684000_1462000# gnd! 487.2fF
C1827 diff_2652000_1544000# gnd! 156.2fF
C1828 diff_2673000_1453000# gnd! 297.7fF
C1829 diff_2532000_1478000# gnd! 242.1fF
C1830 diff_2628000_1544000# gnd! 128.1fF
C1831 diff_2480000_1368000# gnd! 420.9fF
C1832 diff_2875000_1792000# gnd! 143.8fF
C1833 diff_2800000_1698000# gnd! 180.5fF
C1834 diff_2781000_1698000# gnd! 127.0fF
C1835 diff_2628000_1664000# gnd! 118.9fF
C1836 diff_2470000_1450000# gnd! 164.6fF
C1837 diff_2460000_1455000# gnd! 186.6fF
C1838 diff_2382000_1537000# gnd! 99.6fF
C1839 diff_2406000_1570000# gnd! 158.4fF
C1840 diff_2334000_1513000# gnd! 63.5fF
C1841 diff_2487000_1586000# gnd! 224.8fF
C1842 diff_2475000_1616000# gnd! 158.5fF
C1843 diff_2409000_1603000# gnd! 304.4fF
C1844 diff_2416000_1627000# gnd! 88.6fF
C1845 diff_2759000_1758000# gnd! 147.6fF
C1846 diff_2674000_1682000# gnd! 116.5fF
C1847 diff_2652000_1699000# gnd! 154.2fF
C1848 diff_2684000_1778000# gnd! 323.1fF
C1849 diff_2673000_1767000# gnd! 147.7fF
C1850 diff_2886000_1802000# gnd! 820.7fF
C1851 diff_2875000_1828000# gnd! 289.6fF
C1852 diff_2914000_1941000# gnd! 279.1fF
C1853 diff_2759000_1832000# gnd! 982.2fF
C1854 diff_2628000_1728000# gnd! 120.2fF
C1855 diff_2549000_1578000# gnd! 356.4fF
C1856 diff_2290000_1481000# gnd! 273.4fF
C1857 diff_2329000_1617000# gnd! 53.3fF
C1858 diff_2532000_1765000# gnd! 237.8fF
C1859 diff_2655000_1780000# gnd! 645.1fF
C1860 diff_2544000_1737000# gnd! 196.5fF
C1861 diff_2554000_1747000# gnd! 290.0fF
C1862 diff_2461000_1726000# gnd! 175.9fF
C1863 diff_2406000_1691000# gnd! 157.9fF
C1864 diff_2470000_1735000# gnd! 168.4fF
C1865 diff_2544000_1829000# gnd! 193.9fF
C1866 diff_2830000_1864000# gnd! 516.6fF
C1867 diff_2962000_2041000# gnd! 43.3fF
C1868 diff_3011000_2111000# gnd! 50.0fF
C1869 diff_2987000_2077000# gnd! 139.5fF
C1870 diff_3028000_2040000# gnd! 191.9fF
C1871 diff_3005000_2149000# gnd! 43.3fF
C1872 diff_3028000_2299000# gnd! 346.9fF
C1873 diff_2930000_2100000# gnd! 111.4fF
C1874 diff_2913000_2059000# gnd! 110.2fF
C1875 diff_2875000_2169000# gnd! 139.1fF
C1876 diff_2865000_2160000# gnd! 341.7fF
C1877 diff_2846000_2124000# gnd! 120.7fF
C1878 diff_2830000_2069000# gnd! 131.1fF
C1879 diff_2684000_1840000# gnd! 497.8fF
C1880 diff_2651000_1920000# gnd! 161.4fF
C1881 diff_2673000_1830000# gnd! 300.8fF
C1882 diff_2532000_1854000# gnd! 242.0fF
C1883 diff_2480000_1745000# gnd! 427.2fF
C1884 diff_2800000_2075000# gnd! 179.4fF
C1885 diff_2781000_2075000# gnd! 133.3fF
C1886 diff_2628000_2040000# gnd! 1033.3fF
C1887 diff_2470000_1827000# gnd! 169.2fF
C1888 diff_2461000_1832000# gnd! 178.5fF
C1889 diff_2271000_1624000# gnd! 130.2fF
C1890 diff_2103000_1260000# gnd! 16.4fF
C1891 diff_2197000_1226000# gnd! 258.9fF
C1892 diff_2183000_1301000# gnd! 285.9fF
C1893 diff_2122000_1260000# gnd! 402.6fF
C1894 diff_2129000_1288000# gnd! 475.4fF
C1895 diff_2136000_1297000# gnd! 216.0fF
C1896 diff_2126000_1327000# gnd! 745.5fF
C1897 diff_2232000_1463000# gnd! 57.7fF
C1898 diff_2206000_1539000# gnd! 55.2fF
C1899 diff_2121000_1350000# gnd! 666.5fF
C1900 diff_2126000_1544000# gnd! 89.3fF
C1901 diff_2183000_1493000# gnd! 287.1fF
C1902 diff_2136000_1579000# gnd! 207.5fF
C1903 diff_2129000_1594000# gnd! 98.0fF
C1904 diff_1981000_1167000# gnd! 45.6fF
C1905 diff_1996000_1090000# gnd! 256.0fF
C1906 diff_2009000_1240000# gnd! 93.4fF
C1907 diff_1943000_1143000# gnd! 136.2fF
C1908 diff_1880000_1072000# gnd! 132.8fF
C1909 diff_1850000_1078000# gnd! 110.8fF
C1910 diff_1931000_1176000# gnd! 125.2fF
C1911 diff_1869000_1078000# gnd! 343.1fF
C1912 diff_1965000_1244000# gnd! 65.8fF
C1913 diff_1892000_1235000# gnd! 109.5fF
C1914 diff_1891000_1210000# gnd! 357.1fF
C1915 diff_1981000_1324000# gnd! 47.6fF
C1916 diff_1851000_1157000# gnd! 135.8fF
C1917 diff_1833000_1157000# gnd! 110.4fF
C1918 diff_2052000_1346000# gnd! 157.5fF
C1919 diff_2049000_1392000# gnd! 165.8fF
C1920 diff_2015000_1385000# gnd! 147.4fF
C1921 diff_1996000_1361000# gnd! 265.6fF
C1922 diff_2035000_1429000# gnd! 541.9fF
C1923 diff_2052000_1524000# gnd! 154.4fF
C1924 diff_2015000_1467000# gnd! 157.0fF
C1925 diff_1943000_1345000# gnd! 147.4fF
C1926 diff_1931000_1327000# gnd! 114.5fF
C1927 diff_1852000_1318000# gnd! 127.2fF
C1928 diff_1833000_1282000# gnd! 110.0fF
C1929 diff_1869000_1407000# gnd! 346.5fF
C1930 diff_1850000_1375000# gnd! 118.5fF
C1931 diff_1880000_1417000# gnd! 128.2fF
C1932 diff_1889000_1428000# gnd! 838.0fF
C1933 diff_2103000_1606000# gnd! 17.1fF
C1934 diff_2049000_1456000# gnd! 167.9fF
C1935 diff_2123000_1606000# gnd! 388.6fF
C1936 diff_2103000_1636000# gnd! 17.1fF
C1937 diff_2197000_1603000# gnd! 259.0fF
C1938 diff_2329000_1774000# gnd! 440.9fF
C1939 diff_2271000_1558000# gnd! 536.4fF
C1940 diff_2382000_1914000# gnd! 99.6fF
C1941 diff_2310000_1813000# gnd! 637.8fF
C1942 diff_2405000_1947000# gnd! 159.1fF
C1943 diff_2487000_1963000# gnd! 227.3fF
C1944 diff_2475000_1993000# gnd! 158.6fF
C1945 diff_2409000_1980000# gnd! 294.4fF
C1946 diff_2416000_2004000# gnd! 88.6fF
C1947 diff_2759000_2135000# gnd! 147.2fF
C1948 diff_2674000_2059000# gnd! 113.9fF
C1949 diff_2652000_2076000# gnd! 154.1fF
C1950 diff_2684000_2154000# gnd! 323.4fF
C1951 diff_2673000_2143000# gnd! 146.3fF
C1952 diff_2886000_2178000# gnd! 821.1fF
C1953 diff_2875000_2204000# gnd! 292.1fF
C1954 diff_2914000_2317000# gnd! 278.0fF
C1955 diff_2628000_2106000# gnd! 468.4fF
C1956 diff_2549000_1954000# gnd! 361.9fF
C1957 diff_2533000_2142000# gnd! 237.2fF
C1958 diff_2830000_2241000# gnd! 517.9fF
C1959 diff_3457000_2526000# gnd! 266.6fF
C1960 diff_3467000_2748000# gnd! 52.4fF
C1961 diff_3416000_2552000# gnd! 57.1fF
C1962 diff_3364000_2491000# gnd! 148.7fF
C1963 diff_3367000_2749000# gnd! 43.7fF
C1964 diff_4107000_2724000# gnd! 1549.3fF
C1965 diff_4056000_2491000# gnd! 462.3fF
C1966 diff_4003000_2724000# gnd! 708.3fF
C1967 diff_3921000_785000# gnd! 732.3fF
C1968 diff_3900000_2724000# gnd! 463.7fF
C1969 diff_3829000_786000# gnd! 1607.1fF
C1970 diff_3738000_825000# gnd! 1717.8fF
C1971 diff_3748000_2433000# gnd! 464.0fF
C1972 diff_3694000_2724000# gnd! 1820.5fF
C1973 diff_3595000_2394000# gnd! 1622.3fF
C1974 diff_3566000_784000# gnd! 1629.0fF
C1975 diff_3473000_793000# gnd! 1667.5fF
C1976 diff_3488000_2724000# gnd! 807.1fF
C1977 diff_3438000_2491000# gnd! 1711.4fF
C1978 diff_3353000_2408000# gnd! 2631.2fF
C1979 diff_4103000_2777000# gnd! 270.3fF
C1980 diff_4051000_2777000# gnd! 270.3fF
C1981 diff_4000000_2777000# gnd! 270.4fF
C1982 diff_3948000_2777000# gnd! 270.1fF
C1983 diff_3897000_2777000# gnd! 265.4fF
C1984 diff_3845000_2777000# gnd! 267.4fF
C1985 diff_3793000_2777000# gnd! 265.1fF
C1986 diff_3741000_2777000# gnd! 271.6fF
C1987 diff_3691000_2777000# gnd! 267.7fF
C1988 diff_3638000_2777000# gnd! 270.2fF
C1989 diff_3588000_2777000# gnd! 256.1fF
C1990 diff_3535000_2777000# gnd! 263.6fF
C1991 diff_3485000_2777000# gnd! 267.4fF
C1992 diff_3432000_2777000# gnd! 265.4fF
C1993 diff_3382000_2777000# gnd! 267.4fF
C1994 diff_3331000_2538000# gnd! 161.9fF
C1995 diff_3282000_2537000# gnd! 170.0fF
C1996 diff_4516000_3009000# gnd! 247.9fF
C1997 diff_4655000_3019000# gnd! 994.7fF
C1998 diff_4778000_3197000# gnd! 189.1fF
C1999 diff_5438000_3443000# gnd! 90.5fF
C2000 diff_5919000_3448000# gnd! 409.5fF
C2001 diff_5431000_3450000# gnd! 173.1fF
C2002 diff_5577000_3392000# gnd! 157.8fF
C2003 diff_6159000_3508000# gnd! 72.4fF
C2004 diff_5295000_3448000# gnd! 212.5fF
C2005 diff_5471000_3487000# gnd! 78.0fF
C2006 diff_5356000_3321000# gnd! 686.2fF
C2007 diff_6111000_3387000# gnd! 589.4fF
C2008 diff_6184000_3576000# gnd! 274.6fF
C2009 diff_6184000_3601000# gnd! 131.9fF
C2010 diff_6016000_3580000# gnd! 350.3fF
C2011 diff_5659000_3639000# gnd! 107.2fF
C2012 diff_5503000_3629000# gnd! 130.6fF
C2013 diff_5512000_3640000# gnd! 145.5fF
C2014 diff_5396000_3645000# gnd! 90.1fF
C2015 diff_4870000_3350000# gnd! 1017.8fF
C2016 diff_5021000_3614000# gnd! 117.8fF
C2017 diff_5227000_3586000# gnd! 849.2fF
C2018 diff_5396000_3663000# gnd! 624.2fF
C2019 diff_6145000_3753000# gnd! 383.4fF
C2020 diff_6154000_3781000# gnd! 80.6fF
C2021 diff_5396000_3689000# gnd! 92.6fF
C2022 diff_5294000_3705000# gnd! 151.2fF
C2023 diff_5490000_3759000# gnd! 118.3fF
C2024 diff_6154000_3763000# gnd! 398.4fF
C2025 diff_6160000_3829000# gnd! 239.8fF
C2026 diff_6150000_3838000# gnd! 422.7fF
C2027 diff_5500000_3769000# gnd! 97.5fF
C2028 diff_5042000_3670000# gnd! 299.1fF
C2029 diff_5677000_3739000# gnd! 131.0fF
C2030 diff_5500000_3808000# gnd! 95.0fF
C2031 diff_5038000_3681000# gnd! 227.9fF
C2032 diff_5047000_3692000# gnd! 1277.5fF
C2033 diff_4592000_3171000# gnd! 715.0fF
C2034 diff_4461000_2970000# gnd! 181.5fF
C2035 diff_4454000_3014000# gnd! 179.6fF
C2036 diff_4436000_3014000# gnd! 199.6fF
C2037 diff_4362000_2477000# gnd! 1025.6fF
C2038 diff_4305000_1753000# gnd! 740.9fF
C2039 diff_4199000_2721000# gnd! 437.9fF
C2040 diff_4277000_3057000# gnd! 135.2fF
C2041 diff_4628000_3379000# gnd! 195.8fF
C2042 diff_4993000_3786000# gnd! 97.2fF
C2043 diff_6075000_3941000# gnd! 515.7fF
C2044 diff_5982000_3916000# gnd! 525.1fF
C2045 diff_5624000_3937000# gnd! 120.2fF
C2046 diff_5987000_3968000# gnd! 585.9fF
C2047 diff_5695000_3193000# gnd! 944.3fF
C2048 diff_6197000_3984000# gnd! 331.3fF
C2049 diff_5995000_3978000# gnd! 518.8fF
C2050 diff_5320000_3743000# gnd! 286.1fF
C2051 diff_4996000_3825000# gnd! 218.9fF
C2052 diff_4972000_3833000# gnd! 83.0fF
C2053 diff_5227000_3878000# gnd! 832.1fF
C2054 diff_4972000_3873000# gnd! 237.7fF
C2055 diff_5262000_3934000# gnd! 132.2fF
C2056 diff_5263000_3944000# gnd! 302.2fF
C2057 diff_5068000_3913000# gnd! 211.4fF
C2058 diff_4974000_3888000# gnd! 102.5fF
C2059 diff_5273000_3954000# gnd! 368.3fF
C2060 diff_5079000_3925000# gnd! 124.0fF
C2061 diff_4813000_3334000# gnd! 495.9fF
C2062 diff_4715000_3242000# gnd! 568.1fF
C2063 diff_5060000_3958000# gnd! 698.7fF
C2064 diff_5849000_3990000# gnd! 574.2fF
C2065 diff_5624000_3955000# gnd! 450.1fF
C2066 diff_5611000_4009000# gnd! 395.7fF
C2067 diff_5009000_3740000# gnd! 644.9fF
C2068 diff_5355000_4036000# gnd! 127.2fF
C2069 diff_5355000_4054000# gnd! 131.9fF
C2070 diff_5355000_4072000# gnd! 1242.8fF
C2071 diff_5330000_4061000# gnd! 2945.5fF
C2072 diff_5370000_3653000# gnd! 1814.2fF
C2073 diff_5056000_4063000# gnd! 93.0fF
C2074 diff_5917000_4119000# gnd! 815.2fF
C2075 diff_5762000_4183000# gnd! 831.7fF
C2076 diff_6178000_4192000# gnd! 371.5fF
C2077 diff_6157000_4244000# gnd! 71.6fF
C2078 diff_5673000_4155000# gnd! 390.5fF
C2079 diff_5028000_4063000# gnd! 253.9fF
C2080 diff_4779000_3876000# gnd! 141.2fF
C2081 diff_4761000_3820000# gnd! 870.2fF
C2082 diff_5018000_4115000# gnd! 115.1fF
C2083 diff_5113000_4072000# gnd! 561.4fF
C2084 diff_5003000_4149000# gnd! 77.8fF
C2085 diff_5027000_4157000# gnd! 238.2fF
C2086 diff_4716000_3890000# gnd! 132.8fF
C2087 diff_5452000_4209000# gnd! 578.4fF
C2088 diff_6157000_4261000# gnd! 401.3fF
C2089 diff_5163000_4225000# gnd! 408.2fF
C2090 diff_5375000_4231000# gnd! 169.0fF
C2091 diff_5566000_4242000# gnd! 123.9fF
C2092 diff_5574000_4253000# gnd! 131.1fF
C2093 diff_6144000_4250000# gnd! 453.2fF
C2094 diff_5955000_4223000# gnd! 517.0fF
C2095 diff_6030000_4331000# gnd! 89.6fF
C2096 diff_5602000_4299000# gnd! 131.3fF
C2097 diff_5056000_4274000# gnd! 96.4fF
C2098 diff_4696000_3225000# gnd! 1085.7fF
C2099 diff_5090000_4256000# gnd! 253.9fF
C2100 diff_5375000_4258000# gnd! 321.4fF
C2101 diff_5602000_4345000# gnd! 132.6fF
C2102 diff_4240000_2639000# gnd! 1904.8fF
C2103 diff_4980000_4332000# gnd! 111.2fF
C2104 diff_6145000_4382000# gnd! 288.2fF
C2105 diff_6186000_3964000# gnd! 284.2fF
C2106 diff_5170000_4318000# gnd! 517.8fF
C2107 diff_5568000_4410000# gnd! 119.3fF
C2108 diff_5388000_4390000# gnd! 133.6fF
C2109 diff_5345000_4398000# gnd! 730.8fF
C2110 diff_5560000_4417000# gnd! 128.3fF
C2111 diff_5055000_4360000# gnd! 200.8fF
C2112 diff_5825000_4380000# gnd! 458.6fF
C2113 diff_5948000_4451000# gnd! 272.7fF
C2114 diff_6222000_4301000# gnd! 548.7fF
C2115 diff_4302000_2656000# gnd! 1578.5fF
C2116 diff_5257000_4375000# gnd! 710.2fF
C2117 diff_4983000_4429000# gnd! 93.0fF
C2118 diff_5388000_4407000# gnd! 1451.5fF
C2119 diff_4181000_2527000# gnd! 1445.4fF
C2120 diff_5741000_4459000# gnd! 105.8fF
C2121 diff_5979000_4396000# gnd! 469.9fF
C2122 diff_6152000_4535000# gnd! 491.8fF
C2123 diff_5390000_4497000# gnd! 152.7fF
C2124 diff_5396000_4486000# gnd! 164.5fF
C2125 diff_4994000_4439000# gnd! 226.9fF
C2126 diff_5023000_4456000# gnd! 277.9fF
C2127 diff_4510000_3501000# gnd! 286.6fF
C2128 diff_4494000_3313000# gnd! 825.3fF
C2129 diff_4261000_2986000# gnd! 734.6fF
C2130 diff_4307000_3184000# gnd! 105.8fF
C2131 diff_4224000_2933000# gnd! 509.6fF
C2132 diff_4051000_2819000# gnd! 465.1fF
C2133 diff_4155000_3009000# gnd! 158.4fF
C2134 diff_4296000_3177000# gnd! 413.0fF
C2135 diff_4086000_3164000# gnd! 173.4fF
C2136 diff_4067000_3123000# gnd! 359.9fF
C2137 diff_4094000_3084000# gnd! 149.4fF
C2138 diff_3948000_2819000# gnd! 438.9fF
C2139 diff_3845000_2819000# gnd! 529.3fF
C2140 diff_3905000_3048000# gnd! 102.8fF
C2141 diff_4305000_3504000# gnd! 121.1fF
C2142 diff_4021000_2819000# gnd! 818.5fF
C2143 diff_4461000_3007000# gnd! 735.8fF
C2144 diff_4414000_3773000# gnd! 1202.0fF
C2145 diff_4420000_3821000# gnd! 122.3fF
C2146 diff_4375000_3895000# gnd! 123.8fF
C2147 diff_4357000_3757000# gnd! 703.3fF
C2148 diff_4457000_3836000# gnd! 418.2fF
C2149 diff_4515000_3836000# gnd! 657.3fF
C2150 diff_5456000_4543000# gnd! 84.0fF
C2151 diff_5230000_4553000# gnd! 317.4fF
C2152 diff_5073000_4505000# gnd! 284.9fF
C2153 diff_5095000_4555000# gnd! 276.6fF
C2154 diff_5710000_4527000# gnd! 369.9fF
C2155 diff_6078000_4660000# gnd! 120.2fF
C2156 diff_6048000_4640000# gnd! 132.2fF
C2157 diff_5336000_4568000# gnd! 306.2fF
C2158 diff_5159000_4310000# gnd! 217.5fF
C2159 diff_5475000_4642000# gnd! 81.6fF
C2160 diff_5126000_4616000# gnd! 323.1fF
C2161 diff_4805000_4500000# gnd! 889.8fF
C2162 diff_5126000_4638000# gnd! 66.8fF
C2163 diff_5295000_4529000# gnd! 473.8fF
C2164 diff_5336000_4601000# gnd! 619.0fF
C2165 diff_5992000_4718000# gnd! 161.9fF
C2166 diff_6077000_4739000# gnd! 134.6fF
C2167 diff_4921000_4668000# gnd! 193.5fF
C2168 diff_6077000_4788000# gnd! 121.1fF
C2169 diff_5537000_2618000# gnd! 745.2fF
C2170 diff_5642000_4716000# gnd! 401.2fF
C2171 diff_4926000_3399000# gnd! 2945.3fF
C2172 diff_5488000_4717000# gnd! 179.8fF
C2173 diff_6077000_4837000# gnd! 121.1fF
C2174 diff_5487000_4744000# gnd! 143.9fF
C2175 diff_6030000_4850000# gnd! 137.9fF
C2176 diff_5412000_4657000# gnd! 1069.5fF
C2177 diff_5600000_3944000# gnd! 1502.1fF
C2178 diff_6077000_4886000# gnd! 121.1fF
C2179 diff_6030000_4889000# gnd! 164.3fF
C2180 diff_6030000_4912000# gnd! 206.4fF
C2181 diff_5297000_4763000# gnd! 354.2fF
C2182 diff_5219000_4034000# gnd! 1088.4fF
C2183 diff_5097000_4893000# gnd! 1405.8fF
C2184 diff_5067000_4961000# gnd! 1011.0fF
C2185 diff_5038000_4961000# gnd! 1051.7fF
C2186 diff_5008000_4961000# gnd! 1892.6fF
C2187 diff_4750000_4351000# gnd! 598.5fF
C2188 diff_4787000_4475000# gnd! 481.6fF
C2189 diff_4375000_4011000# gnd! 106.8fF
C2190 diff_4264000_3069000# gnd! 1915.2fF
C2191 diff_4526000_4141000# gnd! 367.9fF
C2192 diff_4027000_3053000# gnd! 774.0fF
C2193 diff_4002000_3073000# gnd! 498.8fF
C2194 diff_3814000_2819000# gnd! 578.5fF
C2195 diff_3916000_3245000# gnd! 105.8fF
C2196 diff_3866000_2980000# gnd! 300.8fF
C2197 diff_3741000_2819000# gnd! 488.1fF
C2198 diff_3711000_2819000# gnd! 414.3fF
C2199 diff_3866000_3071000# gnd! 144.9fF
C2200 diff_3535000_2819000# gnd! 420.3fF
C2201 diff_3638000_2819000# gnd! 625.7fF
C2202 diff_4045000_3494000# gnd! 131.3fF
C2203 diff_3608000_2819000# gnd! 739.0fF
C2204 diff_4219000_3817000# gnd! 107.1fF
C2205 diff_4188000_3787000# gnd! 110.2fF
C2206 diff_4162000_3766000# gnd! 322.1fF
C2207 diff_3818000_3048000# gnd! 538.4fF
C2208 diff_3505000_2819000# gnd! 531.0fF
C2209 diff_3603000_3006000# gnd! 311.4fF
C2210 diff_3578000_3163000# gnd! 98.3fF
C2211 diff_3620000_3187000# gnd! 163.7fF
C2212 diff_4213000_3932000# gnd! 597.0fF
C2213 diff_4170000_3958000# gnd! 107.6fF
C2214 diff_4144000_3668000# gnd! 500.1fF
C2215 diff_4422000_4317000# gnd! 980.2fF
C2216 diff_4525000_4434000# gnd! 86.7fF
C2217 diff_4469000_4299000# gnd! 1146.9fF
C2218 diff_4693000_4600000# gnd! 839.7fF
C2219 diff_4646000_4720000# gnd! 886.9fF
C2220 diff_4317000_4211000# gnd! 2050.0fF
C2221 diff_4248000_4332000# gnd! 121.1fF
C2222 diff_4135000_4236000# gnd! 535.5fF
C2223 diff_3792000_3499000# gnd! 163.8fF
C2224 diff_3516000_3069000# gnd! 319.7fF
C2225 diff_3516000_3178000# gnd! 100.6fF
C2226 diff_3432000_2819000# gnd! 575.1fF
C2227 diff_3488000_3125000# gnd! 119.3fF
C2228 diff_3272000_2527000# gnd! 154.4fF
C2229 diff_3236000_2514000# gnd! 201.0fF
C2230 diff_3282000_1425000# gnd! 531.3fF
C2231 diff_3302000_2723000# gnd! 115.4fF
C2232 diff_3255000_1458000# gnd! 571.3fF
C2233 diff_3320000_2526000# gnd! 640.1fF
C2234 diff_3201000_2552000# gnd! 65.3fF
C2235 diff_3149000_2536000# gnd! 20.6fF
C2236 diff_3080000_2440000# gnd! 231.5fF
C2237 diff_2655000_2158000# gnd! 642.8fF
C2238 diff_2544000_2115000# gnd! 331.7fF
C2239 diff_2554000_2126000# gnd! 290.2fF
C2240 diff_2461000_2102000# gnd! 176.8fF
C2241 diff_2406000_2068000# gnd! 157.8fF
C2242 diff_2319000_1882000# gnd! 143.3fF
C2243 diff_2280000_1865000# gnd! 337.4fF
C2244 diff_2183000_1678000# gnd! 287.3fF
C2245 diff_2123000_1636000# gnd! 404.1fF
C2246 diff_2129000_1665000# gnd! 483.4fF
C2247 diff_2136000_1674000# gnd! 216.4fF
C2248 diff_2126000_1704000# gnd! 653.4fF
C2249 diff_2232000_1840000# gnd! 57.8fF
C2250 diff_2206000_1916000# gnd! 55.2fF
C2251 diff_2121000_1727000# gnd! 669.8fF
C2252 diff_2126000_1921000# gnd! 89.3fF
C2253 diff_2183000_1870000# gnd! 290.6fF
C2254 diff_2136000_1956000# gnd! 207.5fF
C2255 diff_2129000_1971000# gnd! 95.3fF
C2256 diff_2339000_1998000# gnd! 58.3fF
C2257 diff_2470000_2111000# gnd! 168.4fF
C2258 diff_2544000_2207000# gnd! 1282.3fF
C2259 diff_2684000_2216000# gnd! 502.9fF
C2260 diff_2652000_2298000# gnd! 157.4fF
C2261 diff_2673000_2206000# gnd! 297.4fF
C2262 diff_2533000_2232000# gnd! 236.6fF
C2263 diff_2480000_2122000# gnd! 425.0fF
C2264 diff_2549000_2332000# gnd! 198.2fF
C2265 diff_2470000_2204000# gnd! 165.1fF
C2266 diff_2461000_2209000# gnd! 177.4fF
C2267 diff_2272000_2002000# gnd! 56.7fF
C2268 diff_1981000_1544000# gnd! 43.3fF
C2269 diff_1996000_1467000# gnd! 258.9fF
C2270 diff_2009000_1617000# gnd! 93.3fF
C2271 diff_1943000_1520000# gnd! 134.6fF
C2272 diff_1880000_1449000# gnd! 128.2fF
C2273 diff_1850000_1455000# gnd! 111.7fF
C2274 diff_1931000_1553000# gnd! 121.0fF
C2275 diff_1869000_1455000# gnd! 347.3fF
C2276 diff_1965000_1620000# gnd! 66.0fF
C2277 diff_1892000_1612000# gnd! 109.5fF
C2278 diff_1891000_1587000# gnd! 361.6fF
C2279 diff_1981000_1701000# gnd! 45.2fF
C2280 diff_1851000_1534000# gnd! 135.6fF
C2281 diff_1833000_1534000# gnd! 104.1fF
C2282 diff_2052000_1723000# gnd! 158.2fF
C2283 diff_2015000_1762000# gnd! 147.4fF
C2284 diff_1996000_1738000# gnd! 265.6fF
C2285 diff_2049000_1769000# gnd! 167.9fF
C2286 diff_2035000_1807000# gnd! 543.2fF
C2287 diff_2015000_1844000# gnd! 157.1fF
C2288 diff_1943000_1723000# gnd! 142.2fF
C2289 diff_1931000_1704000# gnd! 114.0fF
C2290 diff_1852000_1696000# gnd! 125.0fF
C2291 diff_1833000_1660000# gnd! 112.8fF
C2292 diff_1869000_1783000# gnd! 335.1fF
C2293 diff_1850000_1752000# gnd! 123.7fF
C2294 diff_1880000_1793000# gnd! 132.8fF
C2295 diff_1889000_1804000# gnd! 836.0fF
C2296 diff_2052000_1901000# gnd! 155.2fF
C2297 diff_2103000_1983000# gnd! 16.4fF
C2298 diff_2049000_1833000# gnd! 163.3fF
C2299 diff_2123000_1983000# gnd! 386.2fF
C2300 diff_2319000_2129000# gnd! 476.3fF
C2301 diff_2292000_1877000# gnd! 436.6fF
C2302 diff_2280000_2085000# gnd! 331.1fF
C2303 diff_2382000_2291000# gnd! 99.6fF
C2304 diff_2315000_2142000# gnd! 419.4fF
C2305 diff_2405000_2324000# gnd! 160.1fF
C2306 diff_2487000_2340000# gnd! 223.2fF
C2307 diff_2475000_2369000# gnd! 102.8fF
C2308 diff_2591000_970000# gnd! 1662.9fF
C2309 diff_2409000_2357000# gnd! 297.3fF
C2310 diff_2416000_2381000# gnd! 92.7fF
C2311 diff_2319000_2260000# gnd! 147.9fF
C2312 diff_2103000_2013000# gnd! 17.1fF
C2313 diff_2197000_1980000# gnd! 257.3fF
C2314 diff_2183000_2055000# gnd! 286.1fF
C2315 diff_2123000_2013000# gnd! 406.1fF
C2316 diff_2129000_2042000# gnd! 483.9fF
C2317 diff_2136000_2051000# gnd! 216.0fF
C2318 diff_2126000_2081000# gnd! 546.3fF
C2319 diff_2291000_2206000# gnd! 195.3fF
C2320 diff_2206000_2293000# gnd! 55.2fF
C2321 diff_2121000_2103000# gnd! 671.0fF
C2322 diff_2280000_2194000# gnd! 338.8fF
C2323 diff_2292000_2348000# gnd! 215.5fF
C2324 diff_2392000_1580000# gnd! 885.0fF
C2325 diff_3139000_2526000# gnd! 256.5fF
C2326 diff_3149000_2748000# gnd! 52.4fF
C2327 diff_3098000_2440000# gnd! 573.8fF
C2328 diff_3170000_2724000# gnd! 1662.5fF
C2329 diff_3119000_2491000# gnd! 1642.2fF
C2330 diff_3042000_2722000# gnd! 532.1fF
C2331 diff_3064000_2758000# gnd! 38.7fF
C2332 diff_3027000_2553000# gnd! 415.6fF
C2333 diff_2975000_2537000# gnd! 21.9fF
C2334 diff_2965000_2526000# gnd! 266.8fF
C2335 diff_2975000_2748000# gnd! 52.1fF
C2336 diff_2924000_2553000# gnd! 67.7fF
C2337 diff_2872000_2536000# gnd! 24.9fF
C2338 diff_2862000_2526000# gnd! 254.8fF
C2339 diff_2872000_2748000# gnd! 50.0fF
C2340 diff_2821000_2553000# gnd! 46.4fF
C2341 diff_2769000_2536000# gnd! 22.3fF
C2342 diff_2759000_2526000# gnd! 256.5fF
C2343 diff_2769000_2748000# gnd! 50.0fF
C2344 diff_2718000_2552000# gnd! 48.9fF
C2345 diff_2666000_2536000# gnd! 4.9fF
C2346 diff_2655000_2527000# gnd! 275.2fF
C2347 diff_2665000_2748000# gnd! 52.1fF
C2348 diff_2615000_2552000# gnd! 54.9fF
C2349 diff_2562000_2537000# gnd! 22.1fF
C2350 diff_2552000_2526000# gnd! 265.1fF
C2351 diff_2562000_2748000# gnd! 50.0fF
C2352 diff_2392000_2433000# gnd! 768.2fF
C2353 diff_2126000_2298000# gnd! 89.3fF
C2354 diff_2183000_2247000# gnd! 288.6fF
C2355 diff_2136000_2333000# gnd! 209.0fF
C2356 diff_2129000_2349000# gnd! 95.5fF
C2357 diff_1981000_1921000# gnd! 45.6fF
C2358 diff_1996000_1844000# gnd! 258.4fF
C2359 diff_2009000_1994000# gnd! 93.3fF
C2360 diff_1943000_1896000# gnd! 139.6fF
C2361 diff_1880000_1825000# gnd! 129.9fF
C2362 diff_1850000_1832000# gnd! 118.4fF
C2363 diff_1931000_1930000# gnd! 121.7fF
C2364 diff_1869000_1832000# gnd! 347.3fF
C2365 diff_1965000_1997000# gnd! 66.0fF
C2366 diff_1892000_1989000# gnd! 107.7fF
C2367 diff_1891000_1964000# gnd! 362.7fF
C2368 diff_1981000_2078000# gnd! 45.6fF
C2369 diff_1851000_1912000# gnd! 133.5fF
C2370 diff_1833000_1912000# gnd! 103.4fF
C2371 diff_2052000_2101000# gnd! 156.8fF
C2372 diff_2049000_2146000# gnd! 164.3fF
C2373 diff_2015000_2139000# gnd! 146.1fF
C2374 diff_1996000_2115000# gnd! 265.6fF
C2375 diff_2035000_2184000# gnd! 545.3fF
C2376 diff_2052000_2279000# gnd! 156.6fF
C2377 diff_2015000_2221000# gnd! 157.0fF
C2378 diff_1943000_2100000# gnd! 142.3fF
C2379 diff_1931000_2081000# gnd! 116.7fF
C2380 diff_1851000_2073000# gnd! 129.8fF
C2381 diff_1833000_2037000# gnd! 109.0fF
C2382 diff_1869000_2161000# gnd! 337.4fF
C2383 diff_1850000_2129000# gnd! 122.1fF
C2384 diff_1880000_2170000# gnd! 130.3fF
C2385 diff_2197000_2356000# gnd! 148.4fF
C2386 diff_2103000_2359000# gnd! 17.8fF
C2387 diff_2049000_2210000# gnd! 169.2fF
C2388 diff_2123000_2359000# gnd! 389.8fF
C2389 diff_2303000_1745000# gnd! 1643.7fF
C2390 diff_1981000_2297000# gnd! 47.6fF
C2391 diff_1889000_2181000# gnd! 834.7fF
C2392 diff_1996000_2221000# gnd! 255.2fF
C2393 diff_2009000_2371000# gnd! 55.7fF
C2394 diff_1943000_2273000# gnd! 139.1fF
C2395 diff_1880000_2202000# gnd! 132.8fF
C2396 diff_1850000_2209000# gnd! 113.4fF
C2397 diff_1931000_2307000# gnd! 121.8fF
C2398 diff_1869000_2209000# gnd! 340.1fF
C2399 diff_2511000_2555000# gnd! 393.7fF
C2400 diff_2995000_2724000# gnd! 1623.8fF
C2401 diff_2938000_823000# gnd! 682.3fF
C2402 diff_2892000_2724000# gnd! 1721.2fF
C2403 diff_2842000_1949000# gnd! 1646.3fF
C2404 diff_2776000_764000# gnd! 1706.5fF
C2405 diff_2712000_821000# gnd! 1657.0fF
C2406 diff_2640000_933000# gnd! 1563.0fF
C2407 diff_2637000_2491000# gnd! 782.7fF
C2408 diff_2582000_2724000# gnd! 1698.6fF
C2409 diff_2533000_2491000# gnd! 1699.8fF
C2410 diff_3167000_2776000# gnd! 269.8fF
C2411 diff_3114000_2776000# gnd! 267.6fF
C2412 diff_3046000_2782000# gnd! 330.9fF
C2413 diff_2993000_2776000# gnd! 263.1fF
C2414 diff_2940000_2776000# gnd! 261.5fF
C2415 diff_2890000_2776000# gnd! 258.5fF
C2416 diff_2837000_2776000# gnd! 273.0fF
C2417 diff_2787000_2776000# gnd! 267.0fF
C2418 diff_2734000_2776000# gnd! 272.4fF
C2419 diff_2683000_2776000# gnd! 272.6fF
C2420 diff_2631000_2776000# gnd! 266.0fF
C2421 diff_2580000_2776000# gnd! 267.6fF
C2422 diff_2528000_2776000# gnd! 267.6fF
C2423 diff_2108000_871000# gnd! 181.0fF
C2424 diff_1965000_2374000# gnd! 58.1fF
C2425 diff_1891000_2340000# gnd! 209.7fF
C2426 diff_1892000_2366000# gnd! 61.6fF
C2427 diff_1851000_2289000# gnd! 128.1fF
C2428 diff_1833000_2289000# gnd! 109.5fF
C2429 diff_2441000_2691000# gnd! 740.4fF
C2430 diff_2464000_2760000# gnd! 57.9fF
C2431 diff_2447000_2716000# gnd! 1838.2fF
C2432 diff_2444000_2729000# gnd! 825.8fF
C2433 diff_3106000_2804000# gnd! 91.7fF
C2434 diff_3253000_2508000# gnd! 811.6fF
C2435 diff_3238000_1305000# gnd! 1605.6fF
C2436 diff_3356000_3023000# gnd! 130.8fF
C2437 diff_3364000_3032000# gnd! 403.1fF
C2438 diff_3550000_3278000# gnd! 941.3fF
C2439 diff_2837000_2819000# gnd! 696.6fF
C2440 diff_3186000_3100000# gnd! 211.6fF
C2441 diff_3283000_3143000# gnd! 132.6fF
C2442 diff_3232000_3141000# gnd! 121.1fF
C2443 diff_3013000_2819000# gnd! 1425.4fF
C2444 diff_3049000_2819000# gnd! 457.1fF
C2445 diff_2940000_2819000# gnd! 448.6fF
C2446 diff_3187000_2819000# gnd! 1107.7fF
C2447 diff_3943000_3771000# gnd! 148.9fF
C2448 diff_3940000_3885000# gnd! 120.2fF
C2449 diff_4067000_4316000# gnd! 119.1fF
C2450 diff_4466000_4515000# gnd! 245.9fF
C2451 diff_4919000_4771000# gnd! 712.4fF
C2452 diff_4901000_4753000# gnd! 196.0fF
C2453 diff_4882000_4961000# gnd! 724.3fF
C2454 diff_4842000_4667000# gnd! 246.8fF
C2455 diff_4823000_4961000# gnd! 165.6fF
C2456 diff_4769000_4457000# gnd! 149.7fF
C2457 diff_4427000_3812000# gnd! 599.9fF
C2458 diff_4734000_4961000# gnd! 206.2fF
C2459 diff_4381000_4592000# gnd! 411.9fF
C2460 diff_4124000_2819000# gnd! 1097.9fF
C2461 diff_4176000_4456000# gnd! 422.9fF
C2462 diff_4127000_4461000# gnd! 381.7fF
C2463 diff_3908000_4368000# gnd! 371.2fF
C2464 diff_3701000_3517000# gnd! 107.0fF
C2465 diff_3646000_3520000# gnd! 134.6fF
C2466 diff_3443000_3166000# gnd! 883.8fF
C2467 diff_3568000_3529000# gnd! 1820.4fF
C2468 diff_3980000_4516000# gnd! 1102.0fF
C2469 diff_4019000_4532000# gnd! 290.0fF
C2470 diff_3669000_3851000# gnd! 141.7fF
C2471 diff_3121000_3079000# gnd! 140.9fF
C2472 diff_3060000_3051000# gnd! 364.7fF
C2473 diff_3073000_3192000# gnd! 97.3fF
C2474 diff_3025000_3074000# gnd! 115.7fF
C2475 diff_2979000_3081000# gnd! 165.6fF
C2476 diff_2910000_2819000# gnd! 509.0fF
C2477 diff_2908000_3148000# gnd! 289.0fF
C2478 diff_2873000_3144000# gnd! 94.8fF
C2479 diff_2921000_3077000# gnd! 95.1fF
C2480 diff_2807000_2819000# gnd! 495.4fF
C2481 diff_2820000_3093000# gnd! 108.4fF
C2482 diff_2734000_2819000# gnd! 425.0fF
C2483 diff_2743000_3027000# gnd! 113.2fF
C2484 diff_3618000_3825000# gnd! 313.4fF
C2485 diff_3531000_3484000# gnd! 569.6fF
C2486 diff_3676000_3846000# gnd! 130.1fF
C2487 diff_3622000_3885000# gnd! 113.9fF
C2488 diff_3447000_3516000# gnd! 702.7fF
C2489 diff_3582000_4084000# gnd! 108.2fF
C2490 diff_3665000_4068000# gnd! 832.5fF
C2491 diff_3667000_4148000# gnd! 135.6fF
C2492 diff_3534000_3824000# gnd! 525.6fF
C2493 diff_3657000_4141000# gnd! 316.3fF
C2494 diff_3608000_4425000# gnd! 424.9fF
C2495 diff_3886000_4603000# gnd! 277.4fF
C2496 diff_3665000_4489000# gnd! 585.4fF
C2497 diff_3112000_3385000# gnd! 172.1fF
C2498 diff_2987000_3090000# gnd! 534.8fF
C2499 diff_3414000_3851000# gnd! 185.9fF
C2500 diff_2986000_3359000# gnd! 472.5fF
C2501 diff_2316000_2469000# gnd! 173.6fF
C2502 diff_2232000_2217000# gnd! 552.4fF
C2503 diff_2299000_2498000# gnd! 450.4fF
C2504 diff_2385000_2506000# gnd! 353.1fF
C2505 diff_2374000_2501000# gnd! 114.0fF
C2506 diff_2283000_2432000# gnd! 233.2fF
C2507 diff_2310000_2576000# gnd! 58.2fF
C2508 diff_2287000_2487000# gnd! 465.1fF
C2509 diff_2326000_2476000# gnd! 548.5fF
C2510 diff_2337000_2732000# gnd! 202.7fF
C2511 diff_2248000_788000# gnd! 904.3fF
C2512 diff_1790000_797000# gnd! 188.0fF ;**FLOATING
C2513 diff_1773000_759000# gnd! 4.1fF ;**FLOATING
C2514 diff_1674000_771000# gnd! 169.8fF
C2515 diff_1398000_597000# gnd! 159.3fF
C2516 diff_1624000_777000# gnd! 191.6fF
C2517 diff_1520000_785000# gnd! 172.2fF
C2518 diff_1410000_785000# gnd! 151.6fF
C2519 diff_1654000_876000# gnd! 64.5fF
C2520 diff_1577000_869000# gnd! 57.2fF
C2521 diff_1577000_893000# gnd! 195.8fF
C2522 diff_1687000_963000# gnd! 127.4fF
C2523 diff_1707000_998000# gnd! 152.9fF
C2524 diff_1669000_962000# gnd! 121.2fF
C2525 diff_1508000_759000# gnd! 153.4fF
C2526 diff_1518000_870000# gnd! 59.1fF
C2527 diff_1385000_840000# gnd! 115.8fF
C2528 diff_1438000_883000# gnd! 28.4fF
C2529 diff_1584000_927000# gnd! 115.4fF
C2530 diff_1557000_943000# gnd! 154.2fF
C2531 diff_1584000_1025000# gnd! 341.5fF
C2532 diff_1575000_1013000# gnd! 141.3fF
C2533 diff_1584000_1099000# gnd! 486.4fF
C2534 diff_1513000_893000# gnd! 283.6fF
C2535 diff_1503000_945000# gnd! 133.4fF
C2536 diff_1478000_943000# gnd! 185.3fF
C2537 diff_1461000_883000# gnd! 172.9fF
C2538 diff_1557000_1172000# gnd! 161.2fF
C2539 diff_1575000_1088000# gnd! 285.3fF
C2540 diff_1655000_1235000# gnd! 100.6fF
C2541 diff_1577000_1247000# gnd! 57.2fF
C2542 diff_1577000_1211000# gnd! 366.4fF
C2543 diff_1687000_1340000# gnd! 120.5fF
C2544 diff_1707000_1375000# gnd! 160.9fF
C2545 diff_1669000_1339000# gnd! 121.2fF
C2546 diff_1519000_1244000# gnd! 60.5fF
C2547 diff_1478000_1092000# gnd! 485.1fF
C2548 diff_1311000_876000# gnd! 102.0fF
C2549 diff_1391000_919000# gnd! 149.2fF
C2550 diff_1344000_884000# gnd! 356.6fF
C2551 diff_1304000_906000# gnd! 291.8fF
C2552 diff_1402000_1033000# gnd! 72.1fF
C2553 diff_1381000_998000# gnd! 74.2fF
C2554 diff_1334000_997000# gnd! 53.0fF
C2555 diff_1302000_960000# gnd! 58.3fF
C2556 diff_1304000_985000# gnd! 586.2fF
C2557 diff_1391000_1181000# gnd! 150.0fF
C2558 diff_989000_660000# gnd! 54.5fF
C2559 diff_791000_355000# gnd! 2203.2fF
C2560 diff_905000_614000# gnd! 307.0fF
C2561 diff_826000_618000# gnd! 232.2fF
C2562 diff_561000_494000# gnd! 263.3fF
C2563 diff_450000_527000# gnd! 276.0fF
C2564 diff_570000_477000# gnd! 1001.0fF
C2565 diff_105000_354000# gnd! 906.0fF
C2566 diff_588000_587000# gnd! 275.8fF
C2567 diff_450000_605000# gnd! 221.8fF
C2568 diff_1178000_871000# gnd! 88.2fF
C2569 diff_1049000_876000# gnd! 68.5fF
C2570 diff_915000_743000# gnd! 1392.6fF
C2571 diff_450000_657000# gnd! 285.9fF
C2572 diff_122000_487000# gnd! 1924.9fF
C2573 diff_684000_665000# gnd! 215.1fF
C2574 diff_581000_708000# gnd! 314.2fF
C2575 diff_1013000_869000# gnd! 88.2fF
C2576 diff_1461000_1229000# gnd! 177.7fF
C2577 diff_1438000_1229000# gnd! 29.6fF
C2578 diff_1304000_1207000# gnd! 291.7fF
C2579 diff_1237000_974000# gnd! 312.3fF
C2580 diff_1183000_1061000# gnd! 223.7fF
C2581 diff_1344000_1228000# gnd! 360.1fF
C2582 diff_1438000_1260000# gnd! 29.6fF
C2583 diff_1584000_1305000# gnd! 113.7fF
C2584 diff_1558000_1320000# gnd! 153.2fF
C2585 diff_1584000_1402000# gnd! 346.3fF
C2586 diff_1575000_1390000# gnd! 139.3fF
C2587 diff_1584000_1476000# gnd! 488.3fF
C2588 diff_1513000_1270000# gnd! 284.0fF
C2589 diff_1503000_1322000# gnd! 132.3fF
C2590 diff_1478000_1321000# gnd! 185.4fF
C2591 diff_1461000_1260000# gnd! 176.2fF
C2592 diff_1558000_1549000# gnd! 157.4fF
C2593 diff_1575000_1465000# gnd! 282.2fF
C2594 diff_1655000_1612000# gnd! 100.6fF
C2595 diff_1577000_1624000# gnd! 57.2fF
C2596 diff_1577000_1588000# gnd! 366.4fF
C2597 diff_1687000_1717000# gnd! 120.5fF
C2598 diff_1707000_1752000# gnd! 159.2fF
C2599 diff_1756000_738000# gnd! 484.1fF
C2600 diff_1721000_1815000# gnd! 282.6fF
C2601 diff_1669000_1716000# gnd! 121.2fF
C2602 diff_1519000_1621000# gnd! 60.5fF
C2603 diff_1478000_1469000# gnd! 485.3fF
C2604 diff_1312000_1232000# gnd! 167.4fF
C2605 diff_1187000_1218000# gnd! 319.0fF
C2606 diff_1265000_1280000# gnd! 127.2fF
C2607 diff_1391000_1296000# gnd! 150.1fF
C2608 diff_1344000_1261000# gnd! 360.4fF
C2609 diff_1304000_1283000# gnd! 291.3fF
C2610 diff_1402000_1410000# gnd! 72.0fF
C2611 diff_1381000_1375000# gnd! 74.2fF
C2612 diff_1302000_1337000# gnd! 58.4fF
C2613 diff_1334000_1374000# gnd! 52.9fF
C2614 diff_1304000_1362000# gnd! 586.9fF
C2615 diff_1391000_1559000# gnd! 148.7fF
C2616 diff_1461000_1606000# gnd! 178.2fF
C2617 diff_1438000_1606000# gnd! 29.4fF
C2618 diff_1304000_1584000# gnd! 293.1fF
C2619 diff_1187000_1246000# gnd! 73.0fF
C2620 diff_1235000_1244000# gnd! 723.4fF
C2621 diff_753000_679000# gnd! 456.2fF
C2622 diff_1130000_981000# gnd! 101.0fF
C2623 diff_1086000_970000# gnd! 167.5fF
C2624 diff_1065000_932000# gnd! 333.2fF
C2625 diff_940000_870000# gnd! 80.7fF
C2626 diff_553000_832000# gnd! 252.2fF
C2627 diff_133000_497000# gnd! 2687.1fF
C2628 diff_122000_699000# gnd! 1588.3fF
C2629 diff_873000_870000# gnd! 82.3fF
C2630 diff_1003000_1045000# gnd! 92.1fF
C2631 diff_1075000_959000# gnd! 96.1fF
C2632 diff_1009000_1055000# gnd! 175.6fF
C2633 diff_969000_883000# gnd! 646.5fF
C2634 diff_890000_962000# gnd! 50.2fF
C2635 diff_816000_908000# gnd! 44.3fF
C2636 diff_961000_976000# gnd! 112.8fF
C2637 diff_913000_1002000# gnd! 280.2fF
C2638 diff_1086000_1079000# gnd! 166.0fF
C2639 diff_921000_1018000# gnd! 101.2fF
C2640 diff_1009000_1072000# gnd! 184.1fF
C2641 diff_857000_889000# gnd! 233.4fF
C2642 diff_847000_884000# gnd! 95.7fF
C2643 diff_581000_963000# gnd! 319.8fF
C2644 diff_1065000_1079000# gnd! 553.4fF
C2645 diff_1049000_1232000# gnd! 119.1fF
C2646 diff_931000_1029000# gnd! 1361.8fF
C2647 diff_890000_1152000# gnd! 313.6fF
C2648 diff_774000_468000# gnd! 1210.2fF
C2649 diff_913000_1078000# gnd! 276.0fF
C2650 diff_1013000_1246000# gnd! 118.8fF
C2651 diff_1189000_1317000# gnd! 54.1fF
C2652 diff_1187000_1276000# gnd! 359.9fF
C2653 diff_1235000_1425000# gnd! 476.9fF
C2654 diff_1130000_1358000# gnd! 101.0fF
C2655 diff_1086000_1347000# gnd! 167.6fF
C2656 diff_1064000_1309000# gnd! 349.6fF
C2657 diff_940000_1246000# gnd! 119.4fF
C2658 diff_857000_1219000# gnd! 228.3fF
C2659 diff_816000_1210000# gnd! 2055.3fF
C2660 diff_847000_1210000# gnd! 1161.5fF
C2661 diff_122000_865000# gnd! 2429.2fF
C2662 diff_874000_1246000# gnd! 115.8fF
C2663 diff_1003000_1422000# gnd! 92.5fF
C2664 diff_1075000_1336000# gnd! 95.6fF
C2665 diff_1009000_1432000# gnd! 175.6fF
C2666 diff_969000_1260000# gnd! 334.8fF
C2667 diff_890000_1339000# gnd! 50.2fF
C2668 diff_816000_1285000# gnd! 44.3fF
C2669 diff_718000_1031000# gnd! 228.0fF
C2670 diff_133000_875000# gnd! 3575.6fF
C2671 diff_122000_1086000# gnd! 2434.0fF
C2672 diff_961000_1354000# gnd! 113.5fF
C2673 diff_913000_1379000# gnd! 276.0fF
C2674 diff_1175000_1427000# gnd! 484.8fF
C2675 diff_1344000_1605000# gnd! 362.9fF
C2676 diff_1438000_1637000# gnd! 29.6fF
C2677 diff_1584000_1682000# gnd! 113.7fF
C2678 diff_1557000_1697000# gnd! 155.2fF
C2679 diff_1584000_1779000# gnd! 340.4fF
C2680 diff_1575000_1767000# gnd! 141.3fF
C2681 diff_1707000_1881000# gnd! 1967.5fF
C2682 diff_1727000_741000# gnd! 20.5fF ;**FLOATING
C2683 diff_1584000_1853000# gnd! 485.2fF
C2684 diff_1513000_1647000# gnd! 291.8fF
C2685 diff_1503000_1699000# gnd! 125.5fF
C2686 diff_1478000_1698000# gnd! 186.6fF
C2687 diff_1461000_1637000# gnd! 175.5fF
C2688 diff_1557000_1926000# gnd! 159.7fF
C2689 diff_1503000_1891000# gnd! 1294.5fF
C2690 diff_1575000_1842000# gnd! 280.1fF
C2691 diff_1655000_1988000# gnd! 102.2fF
C2692 diff_1577000_2001000# gnd! 57.2fF
C2693 diff_1577000_1964000# gnd! 365.3fF
C2694 diff_1687000_2095000# gnd! 118.8fF
C2695 diff_1707000_2129000# gnd! 202.4fF
C2696 diff_1982000_1350000# gnd! 1183.4fF
C2697 diff_1740000_2095000# gnd! 184.9fF
C2698 diff_1669000_2093000# gnd! 121.2fF
C2699 diff_1519000_1998000# gnd! 60.4fF
C2700 diff_1478000_1847000# gnd! 493.7fF
C2701 diff_1312000_1609000# gnd! 167.6fF
C2702 diff_1197000_1523000# gnd! 280.1fF
C2703 diff_1086000_1456000# gnd! 166.1fF
C2704 diff_921000_1395000# gnd! 100.3fF
C2705 diff_1009000_1449000# gnd! 187.2fF
C2706 diff_857000_1266000# gnd! 231.3fF
C2707 diff_847000_1261000# gnd! 95.3fF
C2708 diff_552000_1245000# gnd! 259.1fF
C2709 diff_450000_1282000# gnd! 275.1fF
C2710 diff_450000_1359000# gnd! 221.8fF
C2711 diff_104000_1093000# gnd! 730.9fF
C2712 diff_586000_1340000# gnd! 259.8fF
C2713 diff_718000_1425000# gnd! 140.0fF
C2714 diff_679000_1428000# gnd! 65.1fF
C2715 diff_450000_1411000# gnd! 744.4fF
C2716 diff_122000_1242000# gnd! 2334.2fF
C2717 diff_1258000_1634000# gnd! 149.0fF
C2718 diff_1391000_1673000# gnd! 150.0fF
C2719 diff_1344000_1638000# gnd! 362.1fF
C2720 diff_1304000_1660000# gnd! 291.3fF
C2721 diff_1402000_1787000# gnd! 72.0fF
C2722 diff_1381000_1752000# gnd! 74.2fF
C2723 diff_1302000_1714000# gnd! 58.4fF
C2724 diff_1334000_1751000# gnd! 52.9fF
C2725 diff_1304000_1739000# gnd! 588.4fF
C2726 diff_1201000_1632000# gnd! 765.2fF
C2727 diff_1188000_1668000# gnd! 112.2fF
C2728 diff_1402000_1836000# gnd! 72.8fF
C2729 diff_1391000_1936000# gnd! 148.7fF
C2730 diff_1334000_1840000# gnd! 53.0fF
C2731 diff_1302000_1910000# gnd! 58.8fF
C2732 diff_1381000_1874000# gnd! 74.8fF
C2733 diff_1461000_1983000# gnd! 179.4fF
C2734 diff_1438000_1983000# gnd! 29.5fF
C2735 diff_1304000_1961000# gnd! 292.2fF
C2736 diff_1264000_1695000# gnd! 488.9fF
C2737 diff_1195000_1873000# gnd! 711.6fF
C2738 diff_1184000_1863000# gnd! 151.3fF
C2739 diff_1263000_1901000# gnd! 105.2fF
C2740 diff_1344000_1982000# gnd! 359.5fF
C2741 diff_1438000_2014000# gnd! 29.6fF
C2742 diff_1584000_2058000# gnd! 115.6fF
C2743 diff_1557000_2075000# gnd! 155.1fF
C2744 diff_1584000_2156000# gnd! 334.8fF
C2745 diff_1575000_2145000# gnd! 139.3fF
C2746 diff_1584000_2230000# gnd! 479.9fF
C2747 diff_1513000_2024000# gnd! 282.4fF
C2748 diff_1503000_2076000# gnd! 136.7fF
C2749 diff_1478000_2075000# gnd! 185.5fF
C2750 diff_1461000_2014000# gnd! 176.1fF
C2751 diff_1557000_2303000# gnd! 158.6fF
C2752 diff_1575000_2219000# gnd! 284.4fF
C2753 diff_1655000_2366000# gnd! 56.2fF
C2754 diff_1577000_2342000# gnd! 196.8fF
C2755 diff_1577000_2378000# gnd! 51.8fF
C2756 diff_1518000_2376000# gnd! 53.3fF
C2757 diff_1478000_2223000# gnd! 490.4fF
C2758 diff_1312000_1986000# gnd! 167.4fF
C2759 diff_1188000_1978000# gnd! 228.8fF
C2760 diff_1391000_2051000# gnd! 149.0fF
C2761 diff_1194000_2002000# gnd! 121.2fF
C2762 diff_1344000_2015000# gnd! 359.6fF
C2763 diff_1304000_2037000# gnd! 290.2fF
C2764 diff_1246000_1991000# gnd! 579.5fF
C2765 diff_1188000_2022000# gnd! 219.8fF
C2766 diff_1263000_2096000# gnd! 108.2fF
C2767 diff_1402000_2164000# gnd! 72.1fF
C2768 diff_1381000_2129000# gnd! 74.2fF
C2769 diff_1334000_2128000# gnd! 53.0fF
C2770 diff_1302000_2091000# gnd! 58.3fF
C2771 diff_1304000_2116000# gnd! 588.6fF
C2772 diff_1184000_2091000# gnd! 150.0fF
C2773 diff_1391000_2313000# gnd! 150.0fF
C2774 diff_1461000_2360000# gnd! 178.7fF
C2775 diff_1438000_2360000# gnd! 29.4fF
C2776 diff_1304000_2338000# gnd! 291.9fF
C2777 diff_1246000_2014000# gnd! 569.3fF
C2778 diff_1344000_2359000# gnd! 361.7fF
C2779 diff_1195000_2101000# gnd! 540.8fF
C2780 diff_2003000_996000# gnd! 1511.5fF
C2781 diff_2185000_2629000# gnd! 428.2fF
C2782 diff_2219000_2489000# gnd! 399.5fF
C2783 diff_2199000_2471000# gnd! 124.5fF
C2784 diff_2230000_2466000# gnd! 535.4fF
C2785 diff_2224000_2739000# gnd! 77.7fF
C2786 diff_2207000_2716000# gnd! 279.6fF
C2787 diff_2170000_2654000# gnd! 134.8fF
C2788 diff_2147000_2552000# gnd! 468.7fF
C2789 diff_2095000_2536000# gnd! 5.0fF
C2790 diff_2084000_2526000# gnd! 274.3fF
C2791 diff_2094000_2748000# gnd! 54.6fF
C2792 diff_2046000_2527000# gnd! 38.3fF
C2793 diff_1857000_1018000# gnd! 1818.5fF
C2794 diff_1836000_1363000# gnd! 1737.0fF
C2795 diff_2112000_2777000# gnd! 275.9fF
C2796 diff_2059000_2776000# gnd! 261.7fF
C2797 diff_2601000_2819000# gnd! 419.7fF
C2798 diff_2631000_2819000# gnd! 636.3fF
C2799 diff_2677000_3054000# gnd! 400.3fF
C2800 diff_2961000_3295000# gnd! 199.0fF
C2801 diff_3211000_3555000# gnd! 331.4fF
C2802 diff_3349000_3930000# gnd! 147.6fF
C2803 diff_3326000_3885000# gnd! 331.2fF
C2804 diff_3338000_4041000# gnd! 126.6fF
C2805 diff_3271000_3282000# gnd! 686.1fF
C2806 diff_3536000_4388000# gnd! 170.3fF
C2807 diff_3400000_3460000# gnd! 969.6fF
C2808 diff_3495000_4369000# gnd! 184.2fF
C2809 diff_3400000_4293000# gnd! 189.7fF
C2810 diff_3381000_4293000# gnd! 214.0fF
C2811 diff_3407000_4287000# gnd! 3808.6fF
C2812 diff_2789000_3478000# gnd! 121.3fF
C2813 diff_2809000_3351000# gnd! 468.3fF
C2814 diff_3016000_3538000# gnd! 232.9fF
C2815 diff_2572000_3038000# gnd! 124.4fF
C2816 diff_2562000_3212000# gnd! 548.0fF
C2817 diff_2520000_3104000# gnd! 106.8fF
C2818 diff_2052000_2804000# gnd! 91.5fF
C2819 diff_1967000_2491000# gnd! 120.3fF
C2820 diff_1915000_2537000# gnd! 423.8fF
C2821 diff_1836000_2528000# gnd! 159.9fF
C2822 diff_1797000_2536000# gnd! 213.9fF
C2823 diff_1728000_1867000# gnd! 538.4fF
C2824 diff_1728000_2090000# gnd! 358.5fF
C2825 diff_1756000_2491000# gnd! 85.8fF
C2826 diff_1986000_2692000# gnd! 351.8fF
C2827 diff_1912000_2695000# gnd! 144.1fF
C2828 diff_1977000_2723000# gnd! 67.5fF
C2829 diff_1930000_2738000# gnd! 372.1fF
C2830 diff_1934000_2757000# gnd! 74.8fF
C2831 diff_1727000_2244000# gnd! 545.0fF
C2832 diff_1779000_2705000# gnd! 74.4fF
C2833 diff_1873000_2768000# gnd! 274.4fF
C2834 diff_1745000_2551000# gnd! 528.9fF
C2835 diff_1694000_2536000# gnd! 21.3fF
C2836 diff_1684000_2526000# gnd! 254.8fF
C2837 diff_1694000_2749000# gnd! 50.0fF
C2838 diff_1591000_2479000# gnd! 84.9fF
C2839 diff_1581000_2469000# gnd! 71.2fF
C2840 diff_1541000_2447000# gnd! 447.1fF
C2841 diff_1354000_780000# gnd! 156.3fF
C2842 diff_1251000_2260000# gnd! 704.3fF
C2843 diff_1188000_2358000# gnd! 358.9fF
C2844 diff_1064000_1456000# gnd! 565.3fF
C2845 diff_1049000_1609000# gnd! 121.4fF
C2846 diff_931000_1406000# gnd! 1356.6fF
C2847 diff_890000_1529000# gnd! 311.6fF
C2848 diff_969000_1622000# gnd! 865.2fF
C2849 diff_913000_1455000# gnd! 274.6fF
C2850 diff_1013000_1623000# gnd! 119.8fF
C2851 diff_1130000_1735000# gnd! 101.0fF
C2852 diff_1086000_1724000# gnd! 168.9fF
C2853 diff_1065000_1686000# gnd! 333.3fF
C2854 diff_940000_1623000# gnd! 119.0fF
C2855 diff_857000_1596000# gnd! 231.6fF
C2856 diff_816000_1587000# gnd! 2609.5fF
C2857 diff_581000_1462000# gnd! 309.2fF
C2858 diff_847000_1587000# gnd! 1289.9fF
C2859 diff_874000_1624000# gnd! 115.7fF
C2860 diff_1003000_1799000# gnd! 92.5fF
C2861 diff_1075000_1713000# gnd! 95.6fF
C2862 diff_1009000_1809000# gnd! 175.6fF
C2863 diff_969000_1637000# gnd! 333.6fF
C2864 diff_889000_1716000# gnd! 50.2fF
C2865 diff_816000_1662000# gnd! 44.3fF
C2866 diff_785000_1585000# gnd! 148.0fF ;**FLOATING
C2867 diff_553000_1586000# gnd! 251.9fF
C2868 diff_133000_1252000# gnd! 2728.7fF
C2869 diff_122000_1452000# gnd! 1619.2fF
C2870 diff_961000_1731000# gnd! 113.5fF
C2871 diff_913000_1756000# gnd! 272.4fF
C2872 diff_1086000_1833000# gnd! 165.9fF
C2873 diff_1075000_1826000# gnd! 97.2fF
C2874 diff_921000_1772000# gnd! 101.2fF
C2875 diff_1009000_1826000# gnd! 187.2fF
C2876 diff_857000_1644000# gnd! 228.8fF
C2877 diff_847000_1638000# gnd! 95.3fF
C2878 diff_581000_1717000# gnd! 319.9fF
C2879 diff_718000_1785000# gnd! 124.5fF
C2880 diff_890000_1906000# gnd! 50.2fF
C2881 diff_1130000_1886000# gnd! 101.0fF
C2882 diff_1003000_1837000# gnd! 92.5fF
C2883 diff_1065000_1833000# gnd! 329.8fF
C2884 diff_1049000_1986000# gnd! 121.6fF
C2885 diff_921000_1827000# gnd! 101.3fF
C2886 diff_931000_1783000# gnd! 1355.3fF
C2887 diff_961000_1837000# gnd! 113.5fF
C2888 diff_969000_1999000# gnd! 331.4fF
C2889 diff_913000_1832000# gnd! 274.6fF
C2890 diff_1013000_2000000# gnd! 119.8fF
C2891 diff_1130000_2112000# gnd! 101.0fF
C2892 diff_1086000_2100000# gnd! 170.4fF
C2893 diff_1065000_2063000# gnd! 337.7fF
C2894 diff_940000_2000000# gnd! 119.0fF
C2895 diff_857000_1973000# gnd! 233.9fF
C2896 diff_816000_1964000# gnd! 36.9fF
C2897 diff_847000_1964000# gnd! 95.4fF
C2898 diff_874000_2000000# gnd! 116.8fF
C2899 diff_1003000_2176000# gnd! 92.1fF
C2900 diff_1075000_2090000# gnd! 95.2fF
C2901 diff_1009000_2186000# gnd! 175.7fF
C2902 diff_969000_2014000# gnd! 334.2fF
C2903 diff_890000_2093000# gnd! 50.2fF
C2904 diff_816000_2039000# gnd! 46.1fF
C2905 diff_961000_2107000# gnd! 112.7fF
C2906 diff_913000_2133000# gnd! 272.4fF
C2907 diff_1086000_2210000# gnd! 167.4fF
C2908 diff_921000_2149000# gnd! 101.2fF
C2909 diff_1009000_2203000# gnd! 182.9fF
C2910 diff_857000_2021000# gnd! 230.4fF
C2911 diff_847000_2015000# gnd! 95.7fF
C2912 diff_122000_1619000# gnd! 2432.2fF
C2913 diff_133000_1629000# gnd! 3585.8fF
C2914 diff_122000_1840000# gnd! 2457.8fF
C2915 diff_552000_1999000# gnd! 266.9fF
C2916 diff_450000_2036000# gnd! 282.2fF
C2917 diff_450000_2113000# gnd! 231.9fF
C2918 diff_586000_2094000# gnd! 259.1fF
C2919 diff_105000_1847000# gnd! 691.9fF
C2920 diff_718000_2179000# gnd! 131.2fF
C2921 diff_679000_2183000# gnd! 64.9fF
C2922 diff_450000_2165000# gnd! 740.0fF
C2923 diff_122000_1996000# gnd! 2319.5fF
C2924 diff_1175000_1642000# gnd! 1529.1fF
C2925 diff_1065000_2210000# gnd! 651.0fF
C2926 diff_931000_2160000# gnd! 1365.4fF
C2927 diff_890000_2283000# gnd! 310.8fF
C2928 diff_913000_2209000# gnd! 272.4fF
C2929 diff_969000_2376000# gnd! 807.7fF
C2930 diff_1093000_1019000# gnd! 977.1fF
C2931 diff_1036000_876000# gnd! 926.2fF
C2932 diff_900000_990000# gnd! 1171.7fF
C2933 diff_857000_2350000# gnd! 229.5fF
C2934 diff_816000_2341000# gnd! 2031.5fF
C2935 diff_581000_2216000# gnd! 309.2fF
C2936 diff_847000_2341000# gnd! 1400.8fF
C2937 diff_876000_1127000# gnd! 1219.7fF
C2938 diff_1507000_2551000# gnd! 270.5fF
C2939 diff_1643000_2549000# gnd! 49.6fF
C2940 diff_1695000_985000# gnd! 1679.4fF
C2941 diff_1642000_832000# gnd! 1648.7fF
C2942 diff_1815000_2508000# gnd! 288.4fF
C2943 diff_1775000_2769000# gnd! 295.1fF
C2944 diff_1546000_931000# gnd! 714.1fF
C2945 diff_1590000_2747000# gnd! 61.0fF
C2946 diff_1486000_840000# gnd! 1843.0fF
C2947 diff_1711000_2777000# gnd! 255.9fF
C2948 diff_1658000_2776000# gnd! 273.9fF
C2949 diff_1236000_1920000# gnd! 1204.7fF
C2950 diff_1384000_2467000# gnd! 309.0fF
C2951 diff_1457000_2547000# gnd! 237.8fF
C2952 diff_1447000_2541000# gnd! 88.0fF
C2953 diff_1485000_2491000# gnd! 425.4fF
C2954 diff_1513000_2747000# gnd! 81.8fF
C2955 diff_1392000_2557000# gnd! 548.7fF
C2956 diff_1410000_2714000# gnd! 70.5fF
C2957 diff_1328000_2491000# gnd! 1063.5fF
C2958 diff_801000_877000# gnd! 2371.9fF
C2959 diff_785000_2340000# gnd! 139.9fF ;**FLOATING
C2960 diff_553000_2340000# gnd! 251.9fF
C2961 diff_133000_2006000# gnd! 2780.1fF
C2962 diff_122000_2206000# gnd! 1611.5fF
C2963 diff_1280000_2491000# gnd! 261.0fF
C2964 diff_1151000_1006000# gnd! 2834.8fF
C2965 diff_1317000_2486000# gnd! 141.5fF
C2966 diff_1309000_2729000# gnd! 144.4fF
C2967 diff_1277000_2573000# gnd! 83.7fF
C2968 diff_1609000_2778000# gnd! 271.4fF
C2969 diff_1553000_2585000# gnd! 300.6fF
C2970 diff_2182000_2692000# gnd! 573.0fF
C2971 diff_2399000_2875000# gnd! 357.3fF
C2972 diff_2463000_2894000# gnd! 488.4fF
C2973 diff_2419000_3101000# gnd! 115.2fF
C2974 diff_2391000_3200000# gnd! 121.4fF
C2975 diff_2355000_3006000# gnd! 387.3fF
C2976 diff_2183000_3047000# gnd! 497.1fF
C2977 diff_2247000_3125000# gnd! 239.9fF
C2978 diff_2292000_3173000# gnd! 427.9fF
C2979 diff_2065000_3012000# gnd! 488.1fF
C2980 diff_2133000_3059000# gnd! 726.4fF
C2981 diff_3047000_3538000# gnd! 301.6fF
C2982 diff_2634000_3303000# gnd! 485.9fF
C2983 diff_2652000_3483000# gnd! 131.8fF
C2984 diff_2109000_2944000# gnd! 608.0fF
C2985 diff_2081000_3200000# gnd! 159.6fF
C2986 diff_1962000_2986000# gnd! 431.1fF
C2987 diff_1999000_3197000# gnd! 117.5fF
C2988 diff_2003000_3054000# gnd! 566.5fF
C2989 diff_1936000_3037000# gnd! 541.7fF
C2990 diff_1809000_946000# gnd! 336.4fF
C2991 diff_1809000_2941000# gnd! 160.7fF
C2992 diff_1750000_2973000# gnd! 482.4fF
C2993 diff_1839000_3082000# gnd! 387.9fF
C2994 diff_1827000_2941000# gnd! 514.7fF
C2995 diff_1961000_3116000# gnd! 224.7fF
C2996 diff_2350000_3073000# gnd! 2307.9fF
C2997 diff_2597000_3303000# gnd! 262.6fF
C2998 diff_2659000_3492000# gnd! 505.1fF
C2999 diff_2771000_3401000# gnd! 1047.7fF
C3000 diff_3004000_3815000# gnd! 212.3fF
C3001 diff_3031000_3773000# gnd! 142.8fF
C3002 diff_1697000_2847000# gnd! 1339.0fF
C3003 diff_1816000_2933000# gnd! 645.8fF
C3004 diff_1732000_2882000# gnd! 997.2fF
C3005 diff_1439000_785000# gnd! 1476.9fF
C3006 diff_1585000_2911000# gnd! 168.1fF
C3007 diff_1258000_2735000# gnd! 217.7fF
C3008 diff_1258000_2793000# gnd! 611.0fF
C3009 diff_1167000_2490000# gnd! 197.7fF
C3010 diff_1084000_2522000# gnd! 510.6fF
C3011 diff_1062000_2499000# gnd! 131.3fF
C3012 diff_1125000_2750000# gnd! 64.0fF
C3013 diff_1087000_2459000# gnd! 52.4fF
C3014 diff_964000_2485000# gnd! 857.9fF
C3015 diff_1156000_2479000# gnd! 131.1fF
C3016 diff_954000_2506000# gnd! 323.6fF
C3017 diff_1715000_2865000# gnd! 893.4fF
C3018 diff_2218000_3480000# gnd! 241.5fF
C3019 diff_2881000_3710000# gnd! 256.9fF
C3020 diff_3023000_3903000# gnd! 108.8fF
C3021 diff_3008000_3949000# gnd! 162.1fF
C3022 diff_2820000_3542000# gnd! 688.5fF
C3023 diff_2910000_3803000# gnd! 414.1fF
C3024 diff_2903000_3861000# gnd! 293.6fF
C3025 diff_2867000_3891000# gnd! 182.6fF
C3026 diff_2964000_3935000# gnd! 130.4fF
C3027 diff_2698000_3826000# gnd! 112.7fF
C3028 diff_2269000_3389000# gnd! 683.7fF
C3029 diff_964000_2516000# gnd! 135.1fF
C3030 diff_947000_2557000# gnd! 239.8fF
C3031 diff_916000_2526000# gnd! 357.1fF
C3032 diff_886000_2526000# gnd! 227.9fF
C3033 diff_581000_2471000# gnd! 320.4fF
C3034 diff_679000_1018000# gnd! 729.9fF
C3035 diff_718000_2539000# gnd! 190.8fF
C3036 diff_855000_2599000# gnd! 162.2fF
C3037 diff_122000_2373000# gnd! 2427.6fF
C3038 diff_133000_2383000# gnd! 3639.9fF
C3039 diff_122000_2594000# gnd! 2482.9fF
C3040 diff_552000_1210000# gnd! 3053.4fF
C3041 diff_937000_2547000# gnd! 487.0fF
C3042 diff_1404000_2968000# gnd! 178.9fF
C3043 diff_1458000_2942000# gnd! 427.2fF
C3044 diff_1481000_3102000# gnd! 129.5fF
C3045 diff_1410000_3065000# gnd! 123.3fF
C3046 diff_1333000_2957000# gnd! 792.6fF
C3047 diff_1339000_3007000# gnd! 630.6fF
C3048 diff_1603000_3122000# gnd! 1447.8fF
C3049 diff_1329000_3050000# gnd! 391.5fF
C3050 diff_1250000_3050000# gnd! 125.0fF
C3051 diff_2339000_3696000# gnd! 215.8fF
C3052 diff_2911000_3917000# gnd! 182.8fF
C3053 diff_2937000_3466000# gnd! 946.9fF
C3054 diff_2852000_4057000# gnd! 80.6fF
C3055 diff_2798000_4039000# gnd! 505.6fF
C3056 diff_3666000_4700000# gnd! 1320.3fF
C3057 diff_3755000_4643000# gnd! 277.5fF
C3058 diff_3701000_4747000# gnd! 1015.7fF
C3059 diff_3540000_4682000# gnd! 90.6fF
C3060 diff_3273000_4384000# gnd! 161.3fF
C3061 diff_3431000_4646000# gnd! 141.7fF
C3062 diff_3420000_4637000# gnd! 440.0fF
C3063 diff_3487000_4661000# gnd! 739.5fF
C3064 diff_3358000_4500000# gnd! 1744.7fF
C3065 diff_3183000_4335000# gnd! 440.7fF
C3066 diff_3034000_4153000# gnd! 705.6fF
C3067 diff_3013000_3474000# gnd! 1099.0fF
C3068 diff_3011000_4153000# gnd! 404.8fF
C3069 diff_2558000_3888000# gnd! 885.0fF
C3070 diff_2896000_4349000# gnd! 109.3fF
C3071 diff_2912000_4303000# gnd! 366.7fF
C3072 diff_3063000_4309000# gnd! 409.0fF
C3073 diff_2876000_4436000# gnd! 112.7fF
C3074 diff_3008000_4522000# gnd! 705.1fF
C3075 diff_2970000_4655000# gnd! 986.0fF
C3076 diff_2930000_4556000# gnd! 1051.9fF
C3077 diff_2916000_4681000# gnd! 71.6fF
C3078 diff_2877000_4621000# gnd! 544.1fF
C3079 diff_2905000_4657000# gnd! 429.4fF
C3080 diff_2859000_4569000# gnd! 643.6fF
C3081 diff_2508000_3808000# gnd! 439.9fF
C3082 diff_2489000_3878000# gnd! 137.4fF
C3083 diff_2470000_3861000# gnd! 114.0fF
C3084 diff_2688000_4367000# gnd! 121.8fF
C3085 diff_2641000_3474000# gnd! 978.5fF
C3086 diff_2648000_4396000# gnd! 134.6fF
C3087 diff_2183000_3680000# gnd! 561.8fF
C3088 diff_2173000_3676000# gnd! 479.8fF
C3089 diff_2027000_3554000# gnd! 417.7fF
C3090 diff_1555000_2818000# gnd! 752.0fF
C3091 diff_1501000_2924000# gnd! 1801.7fF
C3092 diff_1275000_3248000# gnd! 87.8fF
C3093 diff_1189000_3106000# gnd! 744.7fF
C3094 diff_1280000_3070000# gnd! 658.9fF
C3095 diff_1147000_3108000# gnd! 137.0fF
C3096 diff_1027000_3007000# gnd! 503.2fF
C3097 diff_1047000_3118000# gnd! 1283.5fF
C3098 diff_966000_2988000# gnd! 726.9fF
C3099 diff_963000_3081000# gnd! 134.6fF
C3100 diff_916000_3185000# gnd! 119.1fF
C3101 diff_913000_3047000# gnd! 366.2fF
C3102 diff_1978000_3618000# gnd! 214.5fF
C3103 diff_1658000_2819000# gnd! 1124.7fF
C3104 diff_1835000_3560000# gnd! 120.2fF
C3105 diff_874000_3124000# gnd! 126.8fF
C3106 diff_945000_3224000# gnd! 137.7fF
C3107 diff_2072000_3805000# gnd! 305.8fF
C3108 diff_2049000_3806000# gnd! 444.9fF
C3109 diff_2323000_3767000# gnd! 381.6fF
C3110 diff_2336000_4017000# gnd! 105.4fF
C3111 diff_2255000_3931000# gnd! 94.0fF
C3112 diff_2569000_4387000# gnd! 121.1fF
C3113 diff_2155000_3996000# gnd! 537.5fF
C3114 diff_2221000_4171000# gnd! 460.1fF
C3115 diff_2130000_4010000# gnd! 966.1fF
C3116 diff_2112000_3993000# gnd! 201.4fF
C3117 diff_2094000_3974000# gnd! 207.2fF
C3118 diff_2119000_4000000# gnd! 1484.6fF
C3119 diff_1945000_3755000# gnd! 132.8fF
C3120 diff_1464000_3203000# gnd! 721.5fF
C3121 diff_1994000_3920000# gnd! 179.6fF
C3122 diff_1977000_3920000# gnd! 179.6fF
C3123 diff_2197000_2999000# gnd! 1495.1fF
C3124 diff_2565000_3499000# gnd! 1211.1fF
C3125 diff_2404000_4386000# gnd! 338.6fF
C3126 diff_2569000_3911000# gnd! 1045.2fF
C3127 diff_2172000_3037000# gnd! 1430.5fF
C3128 diff_1952000_3749000# gnd! 410.8fF
C3129 diff_1903000_3916000# gnd! 134.6fF
C3130 diff_2193000_4239000# gnd! 214.6fF
C3131 diff_2186000_4494000# gnd! 1008.5fF
C3132 diff_2062000_4303000# gnd! 775.4fF
C3133 diff_2059000_4466000# gnd! 116.2fF
C3134 diff_1474000_3479000# gnd! 107.3fF
C3135 diff_1621000_3413000# gnd! 246.4fF
C3136 diff_1538000_3466000# gnd! 224.0fF
C3137 diff_1560000_3638000# gnd! 291.6fF
C3138 diff_1458000_3631000# gnd! 109.1fF
C3139 diff_1647000_3413000# gnd! 801.2fF
C3140 diff_1712000_3884000# gnd! 313.6fF
C3141 diff_1740000_3999000# gnd! 100.2fF
C3142 diff_1588000_4011000# gnd! 128.9fF
C3143 diff_2004000_4583000# gnd! 245.6fF
C3144 diff_2134000_4720000# gnd! 771.8fF
C3145 diff_1965000_4583000# gnd! 194.9fF
C3146 diff_1275000_3286000# gnd! 2215.2fF
C3147 diff_816000_3049000# gnd! 328.3fF
C3148 diff_742000_2973000# gnd! 1372.7fF
C3149 diff_1096000_3118000# gnd! 1869.3fF
C3150 diff_822000_3288000# gnd! 252.8fF
C3151 diff_1271000_3499000# gnd! 84.7fF
C3152 diff_1339000_3494000# gnd! 163.7fF
C3153 diff_1509000_3891000# gnd! 88.7fF
C3154 diff_1515000_3899000# gnd! 787.2fF
C3155 diff_1692000_4258000# gnd! 251.2fF
C3156 diff_1482000_3489000# gnd! 1165.0fF
C3157 diff_1437000_3777000# gnd! 370.6fF
C3158 diff_1420000_3777000# gnd! 146.5fF
C3159 diff_1405000_3518000# gnd! 406.1fF
C3160 diff_1476000_3931000# gnd! 385.3fF
C3161 diff_639000_3021000# gnd! 106.7fF
C3162 diff_668000_2929000# gnd! 727.8fF
C3163 diff_686000_3100000# gnd! 930.7fF
C3164 diff_1741000_4512000# gnd! 209.6fF
C3165 diff_1550000_4376000# gnd! 96.3fF
C3166 diff_1594000_4501000# gnd! 412.7fF
C3167 diff_1522000_4350000# gnd! 124.8fF
C3168 diff_558000_2987000# gnd! 442.6fF
C3169 diff_533000_2988000# gnd! 165.1fF
C3170 diff_82000_3132000# gnd! 181.4fF
C3171 diff_82000_3149000# gnd! 249.7fF
C3172 diff_103000_3168000# gnd! 439.6fF
C3173 diff_110000_3253000# gnd! 101.1fF
C3174 diff_89000_3264000# gnd! 316.1fF
C3175 diff_1236000_3460000# gnd! 698.1fF
C3176 diff_905000_3225000# gnd! 2150.9fF
C3177 diff_1691000_4496000# gnd! 166.3fF
C3178 diff_1540000_4609000# gnd! 499.4fF
C3179 diff_1673000_4605000# gnd! 745.4fF
C3180 diff_859000_2986000# gnd! 1861.4fF
C3181 diff_127000_3342000# gnd! 269.2fF
C3182 diff_205000_3371000# gnd! 98.5fF
C3183 diff_110000_3357000# gnd! 522.7fF
C3184 diff_905000_3510000# gnd! 199.8fF
C3185 diff_945000_3262000# gnd! 1571.2fF
C3186 diff_1143000_3813000# gnd! 135.6fF
C3187 diff_1151000_3808000# gnd! 153.3fF
C3188 diff_1133000_3806000# gnd! 143.4fF
C3189 diff_1049000_3791000# gnd! 134.6fF
C3190 diff_783000_3632000# gnd! 1368.1fF
C3191 diff_730000_3543000# gnd! 166.8fF
C3192 diff_1078000_3957000# gnd! 105.3fF
C3193 diff_1030000_3948000# gnd! 141.8fF
C3194 diff_986000_3873000# gnd! 225.4fF
C3195 diff_1054000_3958000# gnd! 127.7fF
C3196 diff_857000_3300000# gnd! 1100.7fF
C3197 diff_786000_3668000# gnd! 92.7fF
C3198 diff_110000_3413000# gnd! 129.1fF
C3199 diff_103000_3449000# gnd! 492.1fF
C3200 diff_103000_3495000# gnd! 118.8fF
C3201 diff_87000_3356000# gnd! 285.0fF
C3202 diff_123000_3548000# gnd! 124.0fF
C3203 diff_928000_3955000# gnd! 103.2fF
C3204 diff_996000_3890000# gnd! 122.2fF
C3205 diff_1179000_3098000# gnd! 648.1fF
C3206 diff_1447000_4597000# gnd! 418.9fF
C3207 diff_999000_2989000# gnd! 2014.5fF
C3208 diff_1263000_4412000# gnd! 107.6fF
C3209 diff_1196000_4347000# gnd! 139.7fF
C3210 diff_1150000_4300000# gnd! 186.1fF
C3211 diff_1199000_4479000# gnd! 127.8fF
C3212 diff_1234000_4460000# gnd! 740.4fF
C3213 diff_3228000_4781000# gnd! 1569.6fF
C3214 diff_990000_3075000# gnd! 1606.4fF
C3215 diff_806000_3039000# gnd! 1022.9fF
C3216 diff_93000_3157000# gnd! 2323.4fF
C3217 diff_4616000_4961000# gnd! 245.3fF
C3218 diff_4586000_4961000# gnd! 219.2fF
C3219 diff_4558000_4961000# gnd! 222.6fF
C3220 diff_4528000_4961000# gnd! 834.9fF
C3221 diff_4498000_4961000# gnd! 784.9fF
C3222 diff_4468000_4961000# gnd! 711.5fF
C3223 diff_4318000_4838000# gnd! 1155.5fF
C3224 diff_4410000_4961000# gnd! 391.5fF
C3225 diff_4380000_4961000# gnd! 306.4fF
C3226 diff_4350000_4961000# gnd! 521.9fF
C3227 diff_4322000_4961000# gnd! 250.2fF
C3228 diff_4292000_4961000# gnd! 288.4fF
C3229 diff_4222000_4961000# gnd! 578.9fF
C3230 diff_4192000_4961000# gnd! 784.1fF
C3231 diff_4164000_4928000# gnd! 795.0fF
C3232 diff_4134000_4961000# gnd! 712.4fF
C3233 diff_4104000_4961000# gnd! 472.1fF
C3234 diff_4074000_4961000# gnd! 358.8fF
C3235 diff_4046000_4929000# gnd! 350.2fF
C3236 diff_4016000_4961000# gnd! 346.1fF
C3237 diff_3986000_4961000# gnd! 333.9fF
C3238 diff_3956000_4961000# gnd! 218.8fF
C3239 diff_3928000_4961000# gnd! 679.0fF
C3240 diff_3898000_4961000# gnd! 514.2fF
C3241 diff_3869000_4933000# gnd! 274.8fF
C3242 diff_3839000_4961000# gnd! 776.2fF
C3243 diff_3810000_4961000# gnd! 802.2fF
C3244 diff_3780000_4961000# gnd! 518.6fF
C3245 diff_3712000_4961000# gnd! 593.5fF
C3246 diff_3682000_4961000# gnd! 844.7fF
C3247 diff_3653000_3514000# gnd! 749.4fF
C3248 diff_3624000_4961000# gnd! 247.6fF
C3249 diff_3594000_4961000# gnd! 215.9fF
C3250 diff_3564000_4961000# gnd! 214.1fF
C3251 diff_3536000_4961000# gnd! 435.4fF
C3252 diff_3506000_4961000# gnd! 382.6fF
C3253 diff_3476000_4961000# gnd! 448.9fF
C3254 diff_3446000_4961000# gnd! 444.4fF
C3255 diff_3418000_4961000# gnd! 454.9fF
C3256 diff_3388000_4961000# gnd! 399.0fF
C3257 diff_3359000_4961000# gnd! 446.9fF
C3258 diff_3329000_4961000# gnd! 318.4fF
C3259 diff_3300000_4961000# gnd! 212.2fF
C3260 diff_3270000_4961000# gnd! 436.9fF
C3261 diff_3203000_4961000# gnd! 245.1fF
C3262 diff_3173000_4961000# gnd! 968.0fF
C3263 diff_3105000_3437000# gnd! 583.6fF
C3264 diff_3115000_4961000# gnd! 276.4fF
C3265 diff_3085000_4961000# gnd! 419.9fF
C3266 diff_3055000_4961000# gnd! 210.6fF
C3267 diff_3027000_4946000# gnd! 439.6fF
C3268 diff_2997000_4961000# gnd! 416.4fF
C3269 diff_2967000_4961000# gnd! 466.0fF
C3270 diff_2848000_2985000# gnd! 933.2fF
C3271 diff_2909000_4961000# gnd! 353.2fF
C3272 diff_2879000_4961000# gnd! 276.6fF
C3273 diff_2850000_4961000# gnd! 348.9fF
C3274 diff_2820000_4961000# gnd! 221.1fF
C3275 diff_2791000_4961000# gnd! 226.8fF
C3276 diff_2761000_4961000# gnd! 242.7fF
C3277 diff_2693000_4961000# gnd! 291.4fF
C3278 diff_2663000_4961000# gnd! 485.4fF
C3279 diff_2635000_4961000# gnd! 255.2fF
C3280 diff_2605000_4946000# gnd! 680.0fF
C3281 diff_2576000_4948000# gnd! 364.6fF
C3282 diff_2546000_4961000# gnd! 428.8fF
C3283 diff_2517000_4961000# gnd! 302.7fF
C3284 diff_2487000_4961000# gnd! 285.4fF
C3285 diff_2428000_4961000# gnd! 204.4fF
C3286 diff_2398000_4961000# gnd! 396.8fF
C3287 diff_2370000_4961000# gnd! 311.8fF
C3288 diff_2340000_4961000# gnd! 168.2fF
C3289 diff_2311000_4961000# gnd! 204.1fF
C3290 diff_2281000_4961000# gnd! 215.5fF
C3291 diff_2252000_4961000# gnd! 198.4fF
C3292 diff_2222000_4961000# gnd! 201.4fF
C3293 diff_2154000_4961000# gnd! 228.9fF
C3294 diff_2124000_4961000# gnd! 439.9fF
C3295 diff_2096000_4961000# gnd! 434.8fF
C3296 diff_2066000_4961000# gnd! 422.4fF
C3297 diff_2036000_4961000# gnd! 351.8fF
C3298 diff_2006000_4961000# gnd! 346.4fF
C3299 diff_1978000_4961000# gnd! 688.6fF
C3300 diff_1948000_4961000# gnd! 263.9fF
C3301 diff_1830000_4961000# gnd! 304.4fF
C3302 diff_1800000_4961000# gnd! 424.5fF
C3303 diff_1771000_4961000# gnd! 320.7fF
C3304 diff_1741000_4961000# gnd! 329.9fF
C3305 diff_1712000_4961000# gnd! 308.7fF
C3306 diff_1682000_4961000# gnd! 398.3fF
C3307 diff_1654000_4961000# gnd! 531.9fF
C3308 diff_1624000_4961000# gnd! 746.1fF
C3309 diff_872000_3937000# gnd! 689.1fF
C3310 diff_810000_3855000# gnd! 147.7fF
C3311 diff_791000_3824000# gnd! 525.8fF
C3312 diff_100000_3536000# gnd! 497.2fF
C3313 diff_751000_3796000# gnd! 123.8fF
C3314 diff_731000_3737000# gnd! 439.4fF
C3315 diff_696000_3857000# gnd! 120.2fF
C3316 diff_634000_3799000# gnd! 781.0fF
C3317 diff_651000_3858000# gnd! 131.4fF
C3318 diff_181000_3690000# gnd! 105.3fF
C3319 diff_686000_3825000# gnd! 165.1fF
C3320 diff_607000_3764000# gnd! 357.7fF
C3321 diff_186000_3711000# gnd! 204.8fF
C3322 diff_117000_3657000# gnd! 149.4fF
C3323 diff_91000_3713000# gnd! 1510.6fF
C3324 diff_569000_3596000# gnd! 1029.2fF
C3325 diff_659000_3852000# gnd! 418.1fF
C3326 diff_1125000_4458000# gnd! 132.9fF
C3327 diff_1162000_4604000# gnd! 940.4fF
C3328 diff_1052000_4266000# gnd! 565.8fF
C3329 diff_992000_4387000# gnd! 148.3fF
C3330 diff_974000_4363000# gnd! 349.6fF
C3331 diff_1000000_4393000# gnd! 2152.0fF
C3332 diff_1176000_4477000# gnd! 379.1fF
C3333 diff_1196000_3118000# gnd! 2301.1fF
C3334 diff_1252000_4406000# gnd! 1169.8fF
C3335 diff_1159000_4672000# gnd! 133.6fF
C3336 diff_1075000_4556000# gnd! 709.5fF
C3337 diff_1025000_4535000# gnd! 494.8fF
C3338 diff_690000_4134000# gnd! 669.5fF
C3339 diff_658000_4116000# gnd! 602.8fF
C3340 diff_636000_4099000# gnd! 487.6fF
C3341 diff_726000_4203000# gnd! 554.5fF
C3342 diff_93000_3752000# gnd! 589.5fF
C3343 diff_140000_3843000# gnd! 289.4fF
C3344 diff_131000_3834000# gnd! 146.8fF
C3345 diff_233000_3859000# gnd! 374.2fF
C3346 diff_129000_3948000# gnd! 375.1fF
C3347 diff_105000_3784000# gnd! 479.6fF
C3348 diff_281000_4043000# gnd! 442.2fF
C3349 diff_127000_4096000# gnd! 1018.0fF
C3350 diff_223000_4164000# gnd! 112.9fF
C3351 diff_679000_4313000# gnd! 810.2fF
C3352 diff_772000_4077000# gnd! 869.8fF
C3353 diff_518000_3031000# gnd! 3261.8fF
C3354 diff_935000_4585000# gnd! 546.5fF
C3355 diff_854000_4511000# gnd! 198.0fF
C3356 diff_837000_4492000# gnd! 198.6fF
C3357 diff_794000_4432000# gnd! 122.3fF
C3358 diff_756000_4474000# gnd! 994.3fF
C3359 diff_790000_4021000# gnd! 4994.9fF
C3360 diff_653000_4323000# gnd! 129.2fF
C3361 diff_596000_3012000# gnd! 2839.7fF
C3362 diff_1015000_4729000# gnd! 525.0fF
C3363 diff_1556000_4961000# gnd! 524.4fF
C3364 diff_1527000_4961000# gnd! 241.5fF
C3365 diff_1498000_4961000# gnd! 237.3fF
C3366 diff_1468000_4961000# gnd! 462.6fF
C3367 diff_1439000_4961000# gnd! 273.6fF
C3368 diff_1409000_4961000# gnd! 279.9fF
C3369 diff_1380000_4961000# gnd! 453.1fF
C3370 diff_1350000_4961000# gnd! 813.0fF
C3371 diff_1321000_4961000# gnd! 295.3fF
C3372 diff_1291000_4961000# gnd! 272.4fF
C3373 diff_1262000_4961000# gnd! 252.2fF
C3374 diff_1232000_4961000# gnd! 265.8fF
C3375 diff_1203000_4961000# gnd! 398.7fF
C3376 diff_1144000_4573000# gnd! 423.6fF
C3377 diff_1145000_4961000# gnd! 195.2fF
C3378 diff_1037000_4589000# gnd! 444.6fF
C3379 diff_860000_4691000# gnd! 388.6fF
C3380 diff_740000_4507000# gnd! 733.4fF
C3381 diff_582000_4389000# gnd! 104.2fF
C3382 diff_577000_4446000# gnd! 375.1fF
C3383 diff_685000_4520000# gnd! 1131.6fF
C3384 diff_724000_4489000# gnd! 797.0fF
C3385 diff_100000_4085000# gnd! 791.0fF
C3386 diff_353000_4246000# gnd! 178.2fF
C3387 diff_315000_4257000# gnd! 277.7fF
C3388 diff_97000_4259000# gnd! 237.3fF
C3389 diff_77000_4234000# gnd! 745.5fF
C3390 diff_105000_4267000# gnd! 174.9fF
C3391 diff_529000_4371000# gnd! 3206.4fF
C3392 diff_511000_4351000# gnd! 1706.5fF
C3393 diff_521000_4361000# gnd! 349.9fF
C3394 diff_479000_4479000# gnd! 522.7fF
C3395 diff_87000_4248000# gnd! 407.4fF
C3396 diff_108000_4358000# gnd! 248.8fF
C3397 diff_80000_4320000# gnd! 256.2fF
C3398 diff_82000_4447000# gnd! 337.1fF
C3399 diff_64000_4219000# gnd! 3515.6fF
C3400 diff_166000_4460000# gnd! 663.1fF
C3401 diff_781000_4736000# gnd! 372.1fF
C3402 diff_641000_4582000# gnd! 557.3fF
C3403 diff_530000_4621000# gnd! 4563.4fF
C3404 diff_558000_4357000# gnd! 1098.4fF
C3405 diff_73000_3121000# gnd! 1006.8fF
C3406 diff_336000_4527000# gnd! 1289.6fF
C3407 diff_154000_4529000# gnd! 257.1fF
C3408 diff_168000_4544000# gnd! 2283.6fF
C3409 diff_215000_4573000# gnd! 105.1fF
C3410 diff_105000_4535000# gnd! 119.0fF
C3411 diff_80000_4528000# gnd! 152.4fF
C3412 diff_229000_4600000# gnd! 1245.1fF
C3413 diff_120000_4668000# gnd! 274.4fF
C3414 diff_624000_4564000# gnd! 640.8fF
C3415 diff_230000_4714000# gnd! 213.5fF
C3416 diff_204000_4723000# gnd! 100.3fF
C3417 diff_84000_4682000# gnd! 646.4fF
C3418 diff_200000_4773000# gnd! 163.4fF
C3419 diff_410000_4782000# gnd! 312.2fF
C3420 diff_77000_4694000# gnd! 943.0fF
C3421 diff_983000_4376000# gnd! 463.1fF
C3422 diff_1017000_4961000# gnd! 181.0fF
C3423 diff_987000_4961000# gnd! 189.4fF
C3424 diff_885000_3952000# gnd! 468.4fF
C3425 diff_887000_4705000# gnd! 204.7fF
C3426 diff_860000_4715000# gnd! 190.6fF
C3427 diff_830000_4715000# gnd! 192.2fF
C3428 diff_763000_4720000# gnd! 375.2fF
C3429 diff_667000_4503000# gnd! 570.0fF
C3430 diff_699000_4693000# gnd! 239.8fF
C3431 diff_666000_3268000# gnd! 2017.8fF
C3432 diff_4953000_397000# gnd! 2461.2fF
C3433 diff_5595000_413000# gnd! 5337.0fF
C3434 diff_6227000_5160000# gnd! 443.3fF
C3435 diff_777000_5045000# gnd! 2722.2fF
C3436 diff_445000_4909000# gnd! 1025.1fF
C3437 diff_377000_4962000# gnd! 4925.9fF
C3438 diff_5699000_5119000# gnd! 233.2fF
C3439 diff_5501000_5119000# gnd! 191.7fF
C3440 diff_5971000_5105000# gnd! 356.9fF
C3441 diff_6073000_5170000# gnd! 114.8fF
C3442 diff_5500000_5151000# gnd! 102.8fF
C3443 diff_774000_5075000# gnd! 2963.3fF
C3444 diff_6227000_5190000# gnd! 378.8fF
C3445 diff_6073000_5194000# gnd! 119.0fF
C3446 diff_5971000_5180000# gnd! 327.5fF
C3447 diff_774000_5102000# gnd! 1836.6fF
C3448 diff_5699000_5194000# gnd! 236.4fF
C3449 diff_5501000_5194000# gnd! 195.0fF
C3450 diff_5500000_5226000# gnd! 101.4fF
C3451 diff_774000_5133000# gnd! 2330.7fF
C3452 diff_6171000_5281000# gnd! 454.1fF
C3453 diff_6011000_5271000# gnd! 132.8fF
C3454 diff_5971000_5255000# gnd! 271.1fF
C3455 diff_5599000_574000# gnd! 4163.1fF
C3456 diff_774000_5159000# gnd! 2064.2fF
C3457 diff_5699000_5269000# gnd! 237.5fF
C3458 diff_5501000_5269000# gnd! 193.0fF
C3459 diff_5500000_5301000# gnd! 100.0fF
C3460 diff_464000_5068000# gnd! 526.7fF
C3461 diff_76000_4826000# gnd! 302.6fF
C3462 diff_486000_5097000# gnd! 515.2fF
C3463 diff_513000_5203000# gnd! 261.2fF
C3464 diff_774000_5191000# gnd! 2325.7fF
C3465 diff_5970000_2952000# gnd! 519.2fF
C3466 diff_5971000_5330000# gnd! 302.6fF
C3467 diff_6171000_5341000# gnd! 366.8fF
C3468 diff_6011000_5359000# gnd! 123.9fF
C3469 diff_5699000_5344000# gnd! 236.7fF
C3470 diff_774000_5217000# gnd! 1873.1fF
C3471 diff_5501000_5345000# gnd! 202.8fF
C3472 diff_5500000_5376000# gnd! 98.7fF
C3473 diff_774000_5248000# gnd! 3008.3fF
C3474 diff_94000_5159000# gnd! 3501.6fF
C3475 diff_84000_5212000# gnd! 9.0fF
C3476 diff_99000_3991000# gnd! 2683.2fF
C3477 diff_464000_5279000# gnd! 381.6fF
C3478 diff_501000_5321000# gnd! 154.3fF
C3479 diff_63000_4638000# gnd! 662.9fF
C3480 diff_6016000_5421000# gnd! 118.9fF
C3481 diff_6171000_5415000# gnd! 368.8fF
C3482 diff_5999000_2952000# gnd! 580.1fF
C3483 diff_5971000_5405000# gnd! 281.4fF
C3484 diff_5699000_5420000# gnd! 237.3fF
C3485 diff_774000_5274000# gnd! 1895.1fF
C3486 diff_498000_5333000# gnd! 190.8fF
C3487 diff_492000_5342000# gnd! 176.8fF
C3488 diff_5501000_5420000# gnd! 193.6fF
C3489 diff_5500000_5452000# gnd! 125.7fF
C3490 diff_774000_5305000# gnd! 3065.2fF
C3491 diff_472000_5334000# gnd! 142.2fF
C3492 diff_74000_5300000# gnd! 316.6fF
C3493 diff_6039000_2950000# gnd! 458.8fF
C3494 diff_6195000_5480000# gnd! 327.8fF
C3495 diff_5971000_5481000# gnd! 295.8fF
C3496 diff_6016000_5509000# gnd! 141.9fF
C3497 diff_5699000_5495000# gnd! 228.4fF
C3498 diff_774000_5332000# gnd! 1904.9fF
C3499 diff_5501000_5495000# gnd! 206.8fF
C3500 diff_5500000_5527000# gnd! 113.9fF
C3501 diff_774000_5363000# gnd! 3251.4fF
C3502 diff_6015000_5534000# gnd! 145.9fF
C3503 diff_6195000_5552000# gnd! 328.9fF
C3504 diff_5618000_2171000# gnd! 3750.2fF
C3505 diff_5971000_5556000# gnd! 261.4fF
C3506 diff_5618000_2892000# gnd! 4730.0fF
C3507 diff_5699000_5570000# gnd! 226.4fF
C3508 diff_774000_5389000# gnd! 2338.6fF
C3509 diff_5501000_5570000# gnd! 187.0fF
C3510 diff_6021000_5609000# gnd! 119.3fF
C3511 diff_5500000_5602000# gnd! 103.9fF
C3512 diff_774000_5420000# gnd! 2205.8fF
C3513 diff_6175000_5603000# gnd! 383.9fF
C3514 diff_5971000_5631000# gnd! 343.2fF
C3515 diff_6061000_5631000# gnd! 1160.9fF
C3516 diff_5699000_5645000# gnd! 228.1fF
C3517 diff_401000_4712000# gnd! 2180.0fF
C3518 diff_5081000_5586000# gnd! 838.8fF
C3519 diff_774000_5447000# gnd! 1283.7fF
C3520 diff_5023000_5586000# gnd! 853.0fF
C3521 diff_5501000_5645000# gnd! 187.0fF
C3522 diff_5251000_5061000# gnd! 2560.9fF
C3523 diff_5061000_5620000# gnd! 969.1fF
C3524 diff_5003000_5620000# gnd! 958.1fF
C3525 diff_4925000_5586000# gnd! 870.0fF
C3526 diff_4866000_5586000# gnd! 875.1fF
C3527 diff_4807000_5586000# gnd! 869.5fF
C3528 diff_4905000_5620000# gnd! 968.2fF
C3529 diff_4749000_5586000# gnd! 862.6fF
C3530 diff_4601000_5586000# gnd! 861.7fF
C3531 diff_4542000_5586000# gnd! 853.4fF
C3532 diff_4483000_5586000# gnd! 872.0fF
C3533 diff_4424000_5586000# gnd! 870.6fF
C3534 diff_4365000_5586000# gnd! 850.8fF
C3535 diff_4846000_5620000# gnd! 990.5fF
C3536 diff_4787000_5620000# gnd! 963.4fF
C3537 diff_4729000_5620000# gnd! 976.8fF
C3538 diff_5500000_5677000# gnd! 103.9fF
C3539 diff_774000_5478000# gnd! 2693.0fF
C3540 diff_5953000_5146000# gnd! 751.8fF
C3541 diff_6104000_5744000# gnd! 169.6fF
C3542 diff_5488000_5788000# gnd! 34.7fF
C3543 diff_5774000_5846000# gnd! 2390.3fF
C3544 diff_5927000_6129000# gnd! 2891.0fF
C3545 diff_5508000_5788000# gnd! 693.4fF
C3546 diff_5403000_5746000# gnd! 654.4fF
C3547 diff_5258000_5769000# gnd! 1077.3fF
C3548 diff_4581000_5620000# gnd! 963.3fF
C3549 diff_4522000_5620000# gnd! 995.9fF
C3550 diff_4463000_5620000# gnd! 953.5fF
C3551 diff_4306000_5586000# gnd! 861.4fF
C3552 diff_4404000_5620000# gnd! 976.6fF
C3553 diff_4345000_5620000# gnd! 951.3fF
C3554 diff_4287000_5620000# gnd! 985.1fF
C3555 diff_4207000_5586000# gnd! 880.3fF
C3556 diff_4148000_5586000# gnd! 881.9fF
C3557 diff_4089000_5586000# gnd! 845.8fF
C3558 diff_4187000_5620000# gnd! 944.3fF
C3559 diff_4030000_5586000# gnd! 867.4fF
C3560 diff_3971000_5586000# gnd! 864.4fF
C3561 diff_3912000_5586000# gnd! 862.6fF
C3562 diff_3853000_5586000# gnd! 863.7fF
C3563 diff_3795000_5586000# gnd! 877.7fF
C3564 diff_4128000_5620000# gnd! 989.3fF
C3565 diff_4069000_5620000# gnd! 980.7fF
C3566 diff_4010000_5620000# gnd! 982.8fF
C3567 diff_3951000_5620000# gnd! 972.6fF
C3568 diff_3892000_5620000# gnd! 983.8fF
C3569 diff_3833000_5620000# gnd! 1001.5fF
C3570 diff_3775000_5620000# gnd! 962.9fF
C3571 diff_3697000_5586000# gnd! 852.4fF
C3572 diff_3638000_5586000# gnd! 887.6fF
C3573 diff_3579000_5586000# gnd! 882.5fF
C3574 diff_3520000_5586000# gnd! 856.8fF
C3575 diff_3677000_5620000# gnd! 989.1fF
C3576 diff_3618000_5620000# gnd! 974.5fF
C3577 diff_3461000_5586000# gnd! 874.5fF
C3578 diff_3402000_5586000# gnd! 853.4fF
C3579 diff_3343000_5586000# gnd! 868.7fF
C3580 diff_3285000_5586000# gnd! 859.9fF
C3581 diff_3559000_5620000# gnd! 989.5fF
C3582 diff_3500000_5620000# gnd! 964.4fF
C3583 diff_3441000_5620000# gnd! 958.3fF
C3584 diff_3382000_5620000# gnd! 988.4fF
C3585 diff_3323000_5620000# gnd! 980.8fF
C3586 diff_3265000_5620000# gnd! 978.9fF
C3587 diff_3188000_5586000# gnd! 871.2fF
C3588 diff_3129000_5586000# gnd! 892.6fF
C3589 diff_3070000_5586000# gnd! 870.1fF
C3590 diff_3168000_5620000# gnd! 955.1fF
C3591 diff_3011000_5586000# gnd! 883.1fF
C3592 diff_2952000_5586000# gnd! 870.1fF
C3593 diff_2893000_5586000# gnd! 883.7fF
C3594 diff_2834000_5586000# gnd! 877.5fF
C3595 diff_2776000_5586000# gnd! 860.5fF
C3596 diff_3109000_5620000# gnd! 968.6fF
C3597 diff_3050000_5620000# gnd! 974.9fF
C3598 diff_2991000_5620000# gnd! 963.9fF
C3599 diff_2932000_5620000# gnd! 965.2fF
C3600 diff_2873000_5620000# gnd! 984.7fF
C3601 diff_2814000_5620000# gnd! 992.4fF
C3602 diff_2756000_5620000# gnd! 959.3fF
C3603 diff_2678000_5586000# gnd! 871.9fF
C3604 diff_2619000_5586000# gnd! 881.1fF
C3605 diff_2560000_5586000# gnd! 869.2fF
C3606 diff_2502000_5586000# gnd! 886.3fF
C3607 diff_2413000_5586000# gnd! 857.6fF
C3608 diff_2354000_5586000# gnd! 885.7fF
C3609 diff_2295000_5586000# gnd! 849.6fF
C3610 diff_2237000_5586000# gnd! 872.2fF
C3611 diff_2658000_5620000# gnd! 969.2fF
C3612 diff_2599000_5620000# gnd! 967.8fF
C3613 diff_2540000_5620000# gnd! 965.9fF
C3614 diff_2482000_5620000# gnd! 974.8fF
C3615 diff_4477000_4816000# gnd! 1927.3fF
C3616 diff_5172000_5734000# gnd! 967.2fF
C3617 diff_5429000_5897000# gnd! 372.6fF
C3618 diff_5452000_5801000# gnd! 384.3fF
C3619 diff_5771000_6154000# gnd! 290.4fF
C3620 diff_5760000_6139000# gnd! 2454.8fF
C3621 diff_5256000_3172000# gnd! 5999.0fF
C3622 diff_5405000_5991000# gnd! 729.7fF
C3623 diff_4426000_5700000# gnd! 428.8fF
C3624 diff_4355000_5716000# gnd! 685.3fF
C3625 diff_3961000_5823000# gnd! 314.9fF
C3626 diff_4197000_5802000# gnd! 324.4fF
C3627 diff_3902000_5736000# gnd! 469.1fF
C3628 diff_3871000_5818000# gnd! 766.9fF
C3629 diff_3883000_5843000# gnd! 509.7fF
C3630 diff_3756000_5781000# gnd! 322.6fF
C3631 diff_3676000_5838000# gnd! 605.7fF
C3632 diff_3694000_5840000# gnd! 484.2fF
C3633 diff_2393000_5620000# gnd! 959.5fF
C3634 diff_2334000_5620000# gnd! 983.6fF
C3635 diff_2275000_5620000# gnd! 1017.5fF
C3636 diff_2217000_5620000# gnd! 969.8fF
C3637 diff_2138000_5586000# gnd! 873.7fF
C3638 diff_2080000_5586000# gnd! 857.0fF
C3639 diff_2021000_5586000# gnd! 862.8fF
C3640 diff_1963000_5586000# gnd! 862.6fF
C3641 diff_1814000_5586000# gnd! 856.8fF
C3642 diff_1756000_5586000# gnd! 881.5fF
C3643 diff_1697000_5586000# gnd! 887.0fF
C3644 diff_1638000_5586000# gnd! 850.8fF
C3645 diff_2118000_5620000# gnd! 1002.6fF
C3646 diff_2060000_5620000# gnd! 961.8fF
C3647 diff_2001000_5620000# gnd! 954.8fF
C3648 diff_1943000_5620000# gnd! 954.8fF
C3649 diff_3504000_5808000# gnd! 645.2fF
C3650 diff_3100000_5786000# gnd! 315.1fF
C3651 diff_2984000_5745000# gnd! 190.7fF
C3652 diff_3582000_5809000# gnd! 557.4fF
C3653 diff_5066000_5899000# gnd! 905.4fF
C3654 diff_4397000_6170000# gnd! 848.7fF
C3655 diff_2747000_5771000# gnd! 239.6fF
C3656 diff_1580000_4324000# gnd! 1757.2fF
C3657 diff_2522000_5769000# gnd! 337.1fF
C3658 diff_2612000_5826000# gnd! 125.2fF
C3659 diff_2622000_5835000# gnd! 465.2fF
C3660 diff_2834000_5760000# gnd! 165.0fF
C3661 diff_2840000_5927000# gnd! 693.0fF
C3662 diff_2878000_5744000# gnd! 865.9fF
C3663 diff_2974000_5982000# gnd! 73.3fF ;**FLOATING
C3664 diff_2932000_6014000# gnd! 55.5fF ;**FLOATING
C3665 diff_2886000_5983000# gnd! 92.5fF ;**FLOATING
C3666 diff_2876000_6027000# gnd! 345.5fF ;**FLOATING
C3667 diff_2158000_5725000# gnd! 23.6fF
C3668 diff_2093000_5822000# gnd! 58.5fF
C3669 diff_2072000_5822000# gnd! 15.6fF
C3670 diff_1794000_5620000# gnd! 986.9fF
C3671 diff_1736000_5620000# gnd! 948.5fF
C3672 diff_1677000_5620000# gnd! 975.6fF
C3673 diff_1618000_5620000# gnd! 976.8fF
C3674 diff_1541000_5586000# gnd! 853.6fF
C3675 diff_1483000_5586000# gnd! 853.9fF
C3676 diff_1423000_5586000# gnd! 886.2fF
C3677 diff_1365000_5586000# gnd! 887.5fF
C3678 diff_1305000_5586000# gnd! 864.7fF
C3679 diff_1247000_5586000# gnd! 862.9fF
C3680 diff_1187000_5586000# gnd! 857.4fF
C3681 diff_1129000_5586000# gnd! 860.3fF
C3682 diff_1521000_5620000# gnd! 996.2fF
C3683 diff_1463000_5620000# gnd! 968.4fF
C3684 diff_1403000_5620000# gnd! 956.5fF
C3685 diff_1345000_5620000# gnd! 944.2fF
C3686 diff_1285000_5620000# gnd! 965.3fF
C3687 diff_1227000_5620000# gnd! 946.7fF
C3688 diff_1168000_5620000# gnd! 995.2fF
C3689 diff_1109000_5620000# gnd! 977.5fF
C3690 diff_1031000_5586000# gnd! 895.1fF
C3691 diff_972000_5586000# gnd! 867.7fF
C3692 diff_913000_5586000# gnd! 860.6fF
C3693 diff_854000_5586000# gnd! 845.8fF
C3694 diff_796000_5586000# gnd! 871.5fF
C3695 diff_760000_5560000# gnd! 879.4fF
C3696 diff_1011000_5620000# gnd! 962.5fF
C3697 diff_952000_5620000# gnd! 982.5fF
C3698 diff_893000_5620000# gnd! 977.1fF
C3699 diff_834000_5620000# gnd! 974.9fF
C3700 diff_134000_5506000# gnd! 2039.8fF
C3701 diff_90000_5336000# gnd! 2289.2fF
C3702 diff_505000_5536000# gnd! 2879.8fF
C3703 diff_475000_5142000# gnd! 4732.6fF
C3704 diff_572000_4609000# gnd! 905.4fF
C3705 diff_300000_4193000# gnd! 1468.8fF
C3706 diff_2048000_5822000# gnd! 264.6fF
C3707 diff_2195000_5725000# gnd! 646.2fF
C3708 diff_87000_5399000# gnd! 1520.4fF
C3709 diff_968000_5799000# gnd! 305.9fF
C3710 diff_234000_3316000# gnd! 1039.8fF
C3711 diff_895000_5770000# gnd! 375.3fF
C3712 diff_835000_5745000# gnd! 316.4fF
C3713 diff_508000_5592000# gnd! 132.8fF
C3714 diff_773000_5784000# gnd! 190.6fF
C3715 diff_71000_4514000# gnd! 16730.0fF
C3716 diff_67000_5287000# gnd! 13880.6fF
C3717 diff_93000_3550000# gnd! 5693.3fF
C3718 diff_513000_5775000# gnd! 682.7fF
C3719 diff_1585000_5875000# gnd! 258.4fF
C3720 diff_1647000_5846000# gnd! 559.0fF
C3721 diff_196000_5469000# gnd! 3245.2fF
C3722 diff_94000_5193000# gnd! 138847.0fF
C3723 diff_1585000_6056000# gnd! 1380.4fF
C3724 diff_1119000_5759000# gnd! 1956.3fF
C3725 diff_1277000_5967000# gnd! 1973.1fF
C3726 diff_1129000_5768000# gnd! 4689.3fF
C3727 diff_743000_5833000# gnd! 593.7fF
C3728 diff_1747000_6169000# gnd! 1322.5fF
C3729 diff_4055000_6170000# gnd! 645.2fF
C3730 diff_82000_3097000# gnd! 298862.0fF
C3731 diff_420000_6061000# gnd! 59.0fF ;**FLOATING
C3732 diff_378000_6061000# gnd! 64.0fF ;**FLOATING
C3733 diff_337000_6061000# gnd! 64.0fF ;**FLOATING
C3734 diff_296000_6061000# gnd! 69.6fF ;**FLOATING
C3735 diff_258000_6061000# gnd! 48.0fF ;**FLOATING
C3736 diff_220000_6060000# gnd! 45.6fF ;**FLOATING
C3737 diff_160000_6061000# gnd! 84.5fF ;**FLOATING
C3738 diff_616000_6169000# gnd! 1075.8fF
