* SPICE3 file created from 4004.ext - technology: 4004-nmos-buried-stacked

.option scale=0.001u

M1000 GND N0770 N0385 GND efet w=89900 l=11600
+ ad=-5.44009e+08 pd=4.4776e+06 as=0 ps=0 
M1001 GND GND test GND efet w=119625 l=15225
+ ad=0 pd=0 as=-1.74253e+09 ps=530700 
M1002 reset GND GND GND efet w=118175 l=15225
+ ad=1.54113e+09 pd=301600 as=0 ps=0 
M1003 GND N0754 N0761 GND efet w=26100 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1004 GND PC0_11 N0785 GND efet w=30450 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1005 N0785 N0406 N0770 GND efet w=26100 l=13050
+ ad=0 pd=0 as=1.61262e+09 ps=324800 
M1006 GND N0301 N0754 GND efet w=21750 l=11600
+ ad=0 pd=0 as=7.88438e+08 ps=147900 
M1007 N0761 N0301 N0753 GND efet w=78300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1008 N0754 Vdd Vdd GND efet w=7250 l=69600
+ ad=0 pd=0 as=2.78377e+08 ps=6.03548e+07 
M1009 N0754 N0289 GND GND efet w=23925 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1010 Vdd Vdd N0761 GND efet w=8700 l=30450
+ ad=0 pd=0 as=0 ps=0 
M1011 N0753 N0289 GND GND efet w=136300 l=20300
+ ad=0 pd=0 as=0 ps=0 
M1012 D3 RADB1 N0386 GND efet w=44225 l=13775
+ ad=-1.40613e+09 pd=522000 as=0 ps=0 
M1013 N0385 RADB2 D3 GND efet w=49300 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1014 N0770 WADB2 N0761 GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1015 GND N0289 N0311 GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1016 Vdd N0325 N0301 GND efet w=9425 l=13775
+ ad=0 pd=0 as=-9.51992e+08 ps=582900 
M1017 N0289 M12_M22_CLK1__M11_M12_ D3 GND efet w=21025 l=12325
+ ad=-4.55802e+08 pd=722100 as=0 ps=0 
M1018 N0387 RADB0 D3 GND efet w=44950 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1019 N0290 M12_M22_CLK1__M11_M12_ D2 GND efet w=20300 l=11600
+ ad=4.714e+08 pd=884500 as=1.07438e+09 ps=208800 
M1020 N0311 N0290 N0312 GND efet w=14500 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1021 N0301 N0290 N0302 GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1022 GND N0290 N0755 GND efet w=123250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1023 GND N0740 sync GND efet w=1224525 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1024 N0740 S00531 N0740 GND efet w=70325 l=13050
+ ad=1.77373e+09 pd=2.6738e+06 as=0 ps=0 
M1025 Vdd Vdd S00531 GND efet w=5800 l=13050
+ ad=0 pd=0 as=1.83759e+09 ps=275500 
M1026 Vdd S00531 N0740 GND efet w=10150 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1027 N0738 S00536 N0738 GND efet w=69600 l=13050
+ ad=1.28341e+09 pd=1.8473e+06 as=0 ps=0 
M1028 Vdd S00536 N0738 GND efet w=11600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1029 Vdd Vdd S00536 GND efet w=6525 l=13775
+ ad=0 pd=0 as=1.82918e+09 ps=272600 
M1030 sync N0738 Vdd GND efet w=679325 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1031 N0388 RADB0 D2 GND efet w=42050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1032 Vdd N0325 N0298 GND efet w=13050 l=14500
+ ad=0 pd=0 as=-1.66053e+09 ps=501700 
M1033 N0762 N0298 N0755 GND efet w=68150 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1034 GND N0290 N0756 GND efet w=23200 l=10150
+ ad=0 pd=0 as=6.70697e+08 ps=139200 
M1035 N0756 Vdd Vdd GND efet w=7250 l=68150
+ ad=0 pd=0 as=0 ps=0 
M1036 Vdd Vdd N0762 GND efet w=7250 l=27550
+ ad=0 pd=0 as=0 ps=0 
M1037 N0756 N0298 GND GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1038 N0762 N0756 GND GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1039 GND N0758 N0763 GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1040 GND N0293 N0758 GND efet w=23925 l=11600
+ ad=0 pd=0 as=6.66492e+08 ps=136300 
M1041 N0763 N0293 N0757 GND efet w=70325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1042 N0758 Vdd Vdd GND efet w=7975 l=67425
+ ad=0 pd=0 as=0 ps=0 
M1043 N0758 N0291 GND GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1044 Vdd Vdd N0763 GND efet w=7975 l=29725
+ ad=0 pd=0 as=0 ps=0 
M1045 N0757 N0291 GND GND efet w=125425 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1046 N0298 N0291 N0299 GND efet w=23200 l=18850
+ ad=0 pd=0 as=0 ps=0 
M1047 N0312 N0291 N0313 GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1048 N0302 N0291 N0303 GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1049 Vdd N0325 N0293 GND efet w=9425 l=13775
+ ad=0 pd=0 as=-1.69838e+09 ps=501700 
M1050 N0291 M12_M22_CLK1__M11_M12_ D1 GND efet w=20300 l=11600
+ ad=1.45747e+09 pd=1.0614e+06 as=1.02812e+09 ps=205900 
M1051 N0761 WADB1 N0774 GND efet w=14500 l=13775
+ ad=0 pd=0 as=1.19212e+09 ps=237800 
M1052 N0778 WADB0 N0761 GND efet w=14500 l=11600
+ ad=1.17109e+09 pd=234900 as=0 ps=0 
M1053 N0779 WADB0 N0762 GND efet w=17400 l=10150
+ ad=1.18581e+09 pd=240700 as=0 ps=0 
M1054 N0762 WADB1 N0775 GND efet w=15950 l=13050
+ ad=0 pd=0 as=1.12694e+09 ps=220400 
M1055 D2 RADB1 N0389 GND efet w=44225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1056 N0390 RADB2 D2 GND efet w=47125 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1057 D1 RADB1 N0392 GND efet w=44225 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1058 N0391 RADB2 D1 GND efet w=53650 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1059 N0393 RADB0 D1 GND efet w=43500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1060 N0313 N0292 N0305 GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1061 N0303 N0292 N0294 GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1062 N0299 N0292 N0294 GND efet w=17400 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1063 N0293 N0292 N0294 GND efet w=8700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1064 N0292 M12_M22_CLK1__M11_M12_ D0 GND efet w=23200 l=12325
+ ad=9.21335e+08 pd=954100 as=1.82077e+09 ps=319000 
M1065 GND N0292 N0759 GND efet w=125425 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1066 N0305 N0325 Vdd GND efet w=7975 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1067 N0394 RADB0 D0 GND efet w=43500 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1068 Vdd N0325 N0752 GND efet w=10875 l=14500
+ ad=0 pd=0 as=1.89015e+09 ps=374100 
M1069 N0764 N0752 N0759 GND efet w=69600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1070 GND N0292 N0760 GND efet w=29000 l=11600
+ ad=0 pd=0 as=6.18135e+08 ps=145000 
M1071 N0760 Vdd Vdd GND efet w=7975 l=67425
+ ad=0 pd=0 as=0 ps=0 
M1072 Vdd Vdd N0764 GND efet w=7250 l=27550
+ ad=0 pd=0 as=0 ps=0 
M1073 GND N0307 N0294 GND efet w=31900 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1074 N0760 N0752 GND GND efet w=21750 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1075 N0752 N0307 GND GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1076 N0764 N0760 GND GND efet w=27550 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1077 GND N0738 N0740 GND efet w=101500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1078 N0305 N0307 N0306 GND efet w=14500 l=11600
+ ad=0 pd=0 as=1.50749e+09 ps=292900 
M1079 GND N0295 N0738 GND efet w=112375 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1080 GND PC2_11 N0821 GND efet w=26100 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1081 N0806 PC1_11 GND GND efet w=19575 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1082 N0770 N0424 N0806 GND efet w=26825 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1083 N0821 N0434 N0770 GND efet w=26100 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1084 N0770 N0444 N0834 GND efet w=28275 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1085 N0834 PC3_11 GND GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1086 N0386 N0774 GND GND efet w=72500 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1087 N0385 N0381 PC0_11 GND efet w=6525 l=12325
+ ad=0 pd=0 as=5.61367e+08 ps=130500 
M1088 PC1_11 N0410 N0385 GND efet w=7975 l=10875
+ ad=5.02498e+08 pd=118900 as=0 ps=0 
M1089 N0386 N0381 PC0_7 GND efet w=6525 l=12325
+ ad=0 pd=0 as=5.57162e+08 ps=121800 
M1090 PC1_7 N0410 N0386 GND efet w=5800 l=10150
+ ad=5.40343e+08 pd=118900 as=0 ps=0 
M1091 N0786 N0406 N0774 GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1092 GND PC0_7 N0786 GND efet w=25375 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1093 N0385 N0426 PC2_11 GND efet w=6525 l=12325
+ ad=0 pd=0 as=5.8029e+08 ps=124700 
M1094 PC3_11 N0439 N0385 GND efet w=5800 l=11600
+ ad=4.91985e+08 pd=124700 as=0 ps=0 
M1095 N0386 N0426 PC2_7 GND efet w=6525 l=12325
+ ad=0 pd=0 as=5.02498e+08 ps=121800 
M1096 GND N0778 N0387 GND efet w=72500 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1097 N0787 N0406 N0778 GND efet w=24650 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1098 GND PC0_3 N0787 GND efet w=24650 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1099 N0807 PC1_7 GND GND efet w=22475 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1100 N0774 N0424 N0807 GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1101 N0822 N0434 N0774 GND efet w=26825 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1102 GND PC2_7 N0822 GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1103 N0388 N0779 GND GND efet w=71050 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1104 N0387 N0381 PC0_3 GND efet w=7975 l=12325
+ ad=0 pd=0 as=5.40343e+08 ps=118900 
M1105 N0808 PC1_3 GND GND efet w=23925 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1106 PC3_7 N0439 N0386 GND efet w=5800 l=13050
+ ad=5.50855e+08 pd=121800 as=0 ps=0 
M1107 Vdd __INH__X11_X31_CLK1 N0770 GND efet w=8700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1108 D0 M12_M22_CLK1__M11_M12_ N0497 GND efet w=14500 l=13050
+ ad=0 pd=0 as=1.71354e+09 ps=324800 
M1109 N0862 WRAB1 N0866 GND efet w=17400 l=13050
+ ad=0 pd=0 as=1.1795e+09 ps=229100 
M1110 GND N0866 N0531 GND efet w=63800 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1111 Vdd Vdd N0385 GND efet w=6525 l=31175
+ ad=0 pd=0 as=0 ps=0 
M1112 GND N0497 N0862 GND efet w=109475 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1113 Vdd Vdd N0386 GND efet w=7250 l=30450
+ ad=0 pd=0 as=0 ps=0 
M1114 GND PC2_3 N0823 GND efet w=25375 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1115 N0778 N0424 N0808 GND efet w=25375 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1116 N0823 N0434 N0778 GND efet w=26825 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1117 N0835 PC3_7 GND GND efet w=23925 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1118 N0774 N0444 N0835 GND efet w=26825 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1119 Vdd __INH__X11_X31_CLK1 N0774 GND efet w=9425 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1120 D0 RRAB1 N0531 GND efet w=46400 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1121 N0532 RRAB0 D0 GND efet w=45675 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1122 N0862 Vdd Vdd GND efet w=7975 l=22475
+ ad=0 pd=0 as=0 ps=0 
M1123 N0836 PC3_3 GND GND efet w=23925 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1124 N0778 N0444 N0836 GND efet w=28275 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1125 PC1_3 N0410 N0387 GND efet w=6525 l=10150
+ ad=5.2983e+08 pd=116000 as=0 ps=0 
M1126 N0388 N0381 PC0_2 GND efet w=5800 l=10150
+ ad=0 pd=0 as=5.50855e+08 ps=121800 
M1127 PC1_2 N0410 N0388 GND efet w=5800 l=10150
+ ad=5.36138e+08 pd=121800 as=0 ps=0 
M1128 N0788 N0406 N0779 GND efet w=28275 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1129 GND PC0_2 N0788 GND efet w=24650 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1130 N0387 N0426 PC2_3 GND efet w=6525 l=12325
+ ad=0 pd=0 as=4.83575e+08 ps=116000 
M1131 Vdd __INH__X11_X31_CLK1 N0778 GND efet w=9425 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1132 N0863 Vdd Vdd GND efet w=7975 l=21025
+ ad=0 pd=0 as=0 ps=0 
M1133 PC3_3 N0439 N0387 GND efet w=5800 l=11600
+ ad=5.34035e+08 pd=118900 as=0 ps=0 
M1134 N0388 N0426 PC2_2 GND efet w=6525 l=10150
+ ad=0 pd=0 as=4.89882e+08 ps=118900 
M1135 PC3_2 N0439 N0388 GND efet w=5800 l=11600
+ ad=5.40343e+08 pd=118900 as=0 ps=0 
M1136 GND N0775 N0389 GND efet w=63800 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1137 GND N0771 N0390 GND efet w=68875 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1138 N0771 WADB2 N0762 GND efet w=13050 l=11600
+ ad=1.35401e+09 pd=255200 as=0 ps=0 
M1139 N0789 N0406 N0775 GND efet w=24650 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1140 GND PC0_6 N0789 GND efet w=24650 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1141 N0809 PC1_2 GND GND efet w=23925 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1142 N0779 N0424 N0809 GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1143 N0824 N0434 N0779 GND efet w=26825 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1144 GND PC2_2 N0824 GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1145 GND N0498 N0863 GND efet w=114550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1146 Vdd Vdd N0387 GND efet w=7250 l=31900
+ ad=0 pd=0 as=0 ps=0 
M1147 Vdd Vdd N0388 GND efet w=7975 l=29725
+ ad=0 pd=0 as=0 ps=0 
M1148 N0837 PC3_2 GND GND efet w=23925 l=18125
+ ad=0 pd=0 as=0 ps=0 
M1149 N0810 PC1_6 GND GND efet w=22475 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1150 GND PC2_6 N0825 GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1151 N0775 N0424 N0810 GND efet w=26825 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1152 N0825 N0434 N0775 GND efet w=25375 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1153 N0779 N0444 N0837 GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1154 Vdd __INH__X11_X31_CLK1 N0779 GND efet w=8700 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1155 D1 RRAB1 N0534 GND efet w=44950 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1156 N0533 RRAB0 D1 GND efet w=46400 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1157 N0880 WRAB0 N0862 GND efet w=13775 l=13050
+ ad=1.11853e+09 pd=211700 as=0 ps=0 
M1158 N0532 N0880 GND GND efet w=59450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1159 N0903 N0543 N0866 GND efet w=24650 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1160 GND R1_0 N0903 GND efet w=26100 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1161 N0920 R3_0 GND GND efet w=24650 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1162 N0866 N0565 N0920 GND efet w=24650 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1163 N0929 N0581 N0866 GND efet w=26100 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1164 GND R5_0 N0929 GND efet w=23925 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1165 N0947 R7_0 GND GND efet w=25375 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1166 N0866 N0591 N0947 GND efet w=24650 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1167 N0956 N0616 N0866 GND efet w=26100 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1168 GND R9_0 N0956 GND efet w=26825 l=19575
+ ad=0 pd=0 as=0 ps=0 
M1169 N0966 R11_0 GND GND efet w=25375 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1170 N0531 N0529 R1_0 GND efet w=5800 l=11600
+ ad=0 pd=0 as=6.09725e+08 ps=124700 
M1171 R3_0 N0544 N0531 GND efet w=5800 l=11600
+ ad=6.16033e+08 pd=124700 as=0 ps=0 
M1172 N0531 N0569 R5_0 GND efet w=6525 l=12325
+ ad=0 pd=0 as=5.59265e+08 ps=121800 
M1173 N0532 N0529 R0_0 GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.52958e+08 ps=130500 
M1174 R2_0 N0544 N0532 GND efet w=5800 l=11600
+ ad=5.69777e+08 pd=136300 as=0 ps=0 
M1175 N0904 N0543 N0880 GND efet w=27550 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1176 GND R0_0 N0904 GND efet w=24650 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1177 R7_0 N0583 N0531 GND efet w=5800 l=11600
+ ad=6.16033e+08 pd=127600 as=0 ps=0 
M1178 GND R0_1 N0905 GND efet w=23925 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1179 N0498 M12_M22_CLK1__M11_M12_ D1 GND efet w=13050 l=11600
+ ad=1.63785e+09 pd=330600 as=0 ps=0 
M1180 N0838 PC3_6 GND GND efet w=24650 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1181 N0775 N0444 N0838 GND efet w=25375 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1182 N0389 N0381 PC0_6 GND efet w=7975 l=12325
+ ad=0 pd=0 as=5.2983e+08 ps=121800 
M1183 PC1_6 N0410 N0389 GND efet w=5800 l=12325
+ ad=5.36138e+08 pd=118900 as=0 ps=0 
M1184 N0390 N0381 PC0_10 GND efet w=5800 l=10150
+ ad=0 pd=0 as=5.34035e+08 ps=118900 
M1185 PC1_10 N0410 N0390 GND efet w=5800 l=10150
+ ad=5.36138e+08 pd=116000 as=0 ps=0 
M1186 N0790 N0406 N0771 GND efet w=27550 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1187 GND PC0_10 N0790 GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1188 N0389 N0426 PC2_6 GND efet w=6525 l=10875
+ ad=0 pd=0 as=4.89882e+08 ps=118900 
M1189 PC3_6 N0439 N0389 GND efet w=5800 l=10150
+ ad=5.36138e+08 pd=121800 as=0 ps=0 
M1190 N0390 N0426 PC2_10 GND efet w=5800 l=10150
+ ad=0 pd=0 as=4.8778e+08 ps=118900 
M1191 PC3_10 N0439 N0390 GND efet w=5800 l=10150
+ ad=5.40343e+08 pd=118900 as=0 ps=0 
M1192 GND N0772 N0391 GND efet w=73225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1193 N0772 WADB2 N0763 GND efet w=14500 l=10875
+ ad=1.35191e+09 pd=261000 as=0 ps=0 
M1194 N0763 WADB1 N0776 GND efet w=14500 l=13050
+ ad=0 pd=0 as=1.16058e+09 ps=232000 
M1195 N0791 N0406 N0772 GND efet w=26825 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1196 GND PC0_9 N0791 GND efet w=24650 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1197 N0811 PC1_10 GND GND efet w=23200 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1198 N0771 N0424 N0811 GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1199 N0826 N0434 N0771 GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1200 GND PC2_10 N0826 GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1201 Vdd __INH__X11_X31_CLK1 N0775 GND efet w=8700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1202 N0499 M12_M22_CLK1__M11_M12_ D2 GND efet w=14500 l=13050
+ ad=1.67359e+09 pd=316100 as=0 ps=0 
M1203 N0780 WADB0 N0763 GND efet w=14500 l=13050
+ ad=1.1732e+09 pd=229100 as=0 ps=0 
M1204 N0781 WADB0 N0764 GND efet w=15225 l=12325
+ ad=1.18371e+09 pd=229100 as=0 ps=0 
M1205 N0392 N0776 GND GND efet w=65975 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1206 N0391 N0381 PC0_9 GND efet w=6525 l=13050
+ ad=0 pd=0 as=5.25625e+08 ps=116000 
M1207 N0812 PC1_9 GND GND efet w=23200 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1208 GND PC2_9 N0827 GND efet w=26100 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1209 N0772 N0424 N0812 GND efet w=25375 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1210 N0827 N0434 N0772 GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1211 N0839 PC3_10 GND GND efet w=24650 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1212 N0771 N0444 N0839 GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1213 Vdd Vdd N0389 GND efet w=6525 l=29725
+ ad=0 pd=0 as=0 ps=0 
M1214 D2 RRAB1 N0535 GND efet w=44225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1215 GND N0499 N0864 GND efet w=109475 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1216 Vdd Vdd N0390 GND efet w=7975 l=28275
+ ad=0 pd=0 as=0 ps=0 
M1217 Vdd __INH__X11_X31_CLK1 N0771 GND efet w=10150 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1218 N0881 WRAB0 N0863 GND efet w=13050 l=13050
+ ad=1.08489e+09 pd=208800 as=0 ps=0 
M1219 N0863 WRAB1 N0867 GND efet w=13050 l=11600
+ ad=0 pd=0 as=1.10592e+09 ps=214600 
M1220 N0864 WRAB1 N0868 GND efet w=13050 l=11600
+ ad=0 pd=0 as=1.11643e+09 ps=211700 
M1221 N0840 PC3_9 GND GND efet w=25375 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1222 PC1_9 N0410 N0391 GND efet w=5800 l=11600
+ ad=4.91985e+08 pd=118900 as=0 ps=0 
M1223 PC1_5 N0410 N0392 GND efet w=5800 l=13050
+ ad=4.94087e+08 pd=121800 as=0 ps=0 
M1224 N0392 N0381 PC0_5 GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.23522e+08 ps=116000 
M1225 N0792 N0406 N0776 GND efet w=28275 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1226 GND PC0_5 N0792 GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1227 N0391 N0426 PC2_9 GND efet w=5800 l=10150
+ ad=0 pd=0 as=5.2142e+08 ps=130500 
M1228 N0772 N0444 N0840 GND efet w=25375 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1229 PC3_9 N0439 N0391 GND efet w=5800 l=10150
+ ad=5.50855e+08 pd=121800 as=0 ps=0 
M1230 N0392 N0426 PC2_5 GND efet w=5800 l=10150
+ ad=0 pd=0 as=5.19318e+08 ps=130500 
M1231 N0813 PC1_5 GND GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1232 GND PC0_1 N0793 GND efet w=25375 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1233 GND N0780 N0393 GND efet w=69600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1234 N0793 N0406 N0780 GND efet w=25375 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1235 N0776 N0424 N0813 GND efet w=26825 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1236 N0828 N0434 N0776 GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1237 GND PC2_5 N0828 GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1238 PC3_5 N0439 N0392 GND efet w=5800 l=11600
+ ad=5.57162e+08 pd=121800 as=0 ps=0 
M1239 N0841 PC3_5 GND GND efet w=23925 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1240 N0776 N0444 N0841 GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1241 N0394 N0781 GND GND efet w=68150 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1242 N0393 N0381 PC0_1 GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.31933e+08 ps=118900 
M1243 N0814 PC1_1 GND GND efet w=24650 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1244 GND PC2_1 N0829 GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1245 N0780 N0424 N0814 GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1246 N0829 N0434 N0780 GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1247 N0864 Vdd Vdd GND efet w=7250 l=20300
+ ad=0 pd=0 as=0 ps=0 
M1248 Vdd __INH__X11_X31_CLK1 N0772 GND efet w=9425 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1249 Vdd Vdd N0391 GND efet w=7975 l=28275
+ ad=0 pd=0 as=0 ps=0 
M1250 N0865 Vdd Vdd GND efet w=7975 l=20300
+ ad=0 pd=0 as=0 ps=0 
M1251 GND N0500 N0865 GND efet w=114550 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1252 N0536 RRAB0 D2 GND efet w=44950 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1253 GND N0881 N0533 GND efet w=59450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1254 N0534 N0867 GND GND efet w=60175 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1255 N0905 N0543 N0881 GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1256 N0921 R2_0 GND GND efet w=29000 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1257 N0880 N0565 N0921 GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1258 N0930 N0581 N0880 GND efet w=26100 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1259 N0532 N0569 R4_0 GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.50855e+08 ps=121800 
M1260 GND R4_0 N0930 GND efet w=21750 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1261 N0922 R2_1 GND GND efet w=26825 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1262 N0533 N0529 R0_1 GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.48753e+08 ps=130500 
M1263 R6_0 N0583 N0532 GND efet w=5800 l=11600
+ ad=5.73983e+08 pd=124700 as=0 ps=0 
M1264 N0948 R6_0 GND GND efet w=24650 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1265 N0866 N0632 N0966 GND efet w=30450 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1266 N0975 N0645 N0866 GND efet w=27550 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1267 GND R13_0 N0975 GND efet w=26825 l=18850
+ ad=0 pd=0 as=0 ps=0 
M1268 N0984 R15_0 GND GND efet w=27550 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1269 N0866 N0657 N0984 GND efet w=29000 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1270 N0880 N0591 N0948 GND efet w=26825 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1271 N0531 N0598 R9_0 GND efet w=5800 l=13050
+ ad=0 pd=0 as=6.1393e+08 ps=136300 
M1272 R11_0 N0619 N0531 GND efet w=7975 l=12325
+ ad=6.16033e+08 pd=124700 as=0 ps=0 
M1273 N0532 N0598 R8_0 GND efet w=7250 l=13050
+ ad=0 pd=0 as=5.50855e+08 ps=121800 
M1274 GND R8_0 N0957 GND efet w=21750 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1275 R10_0 N0619 N0532 GND efet w=6525 l=12325
+ ad=5.86598e+08 pd=127600 as=0 ps=0 
M1276 N0957 N0616 N0880 GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1277 GND R4_1 N0931 GND efet w=23200 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1278 N0881 N0565 N0922 GND efet w=28275 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1279 N0931 N0581 N0881 GND efet w=25375 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1280 N0531 N0634 R13_0 GND efet w=5800 l=13050
+ ad=0 pd=0 as=6.24442e+08 ps=124700 
M1281 R15_0 N0647 N0531 GND efet w=5800 l=14500
+ ad=6.26545e+08 pd=127600 as=0 ps=0 
M1282 N0532 N0634 R12_0 GND efet w=7250 l=13775
+ ad=0 pd=0 as=5.48753e+08 ps=118900 
M1283 N0949 R6_1 GND GND efet w=25375 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1284 N0881 N0591 N0949 GND efet w=27550 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1285 R2_1 N0544 N0533 GND efet w=5800 l=11600
+ ad=5.19318e+08 pd=130500 as=0 ps=0 
M1286 N0534 N0529 R1_1 GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.52958e+08 ps=121800 
M1287 R3_1 N0544 N0534 GND efet w=5800 l=11600
+ ad=5.36138e+08 pd=130500 as=0 ps=0 
M1288 N0906 N0543 N0867 GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1289 GND R1_1 N0906 GND efet w=23200 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1290 N0533 N0569 R4_1 GND efet w=6525 l=10875
+ ad=0 pd=0 as=5.3824e+08 ps=118900 
M1291 N0958 N0616 N0881 GND efet w=25375 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1292 GND R8_1 N0958 GND efet w=22475 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1293 N0967 R10_0 GND GND efet w=26825 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1294 N0880 N0632 N0967 GND efet w=25375 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1295 N0976 N0645 N0880 GND efet w=25375 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1296 GND R12_0 N0976 GND efet w=20300 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1297 R14_0 N0647 N0532 GND efet w=7975 l=15225
+ ad=6.26545e+08 pd=124700 as=0 ps=0 
M1298 N0968 R10_1 GND GND efet w=26100 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1299 N0881 N0632 N0968 GND efet w=26100 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1300 N0985 R14_0 GND GND efet w=26100 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1301 N0880 N0657 N0985 GND efet w=26100 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1302 R6_1 N0583 N0533 GND efet w=5800 l=11600
+ ad=5.34035e+08 pd=121800 as=0 ps=0 
M1303 N0534 N0569 R5_1 GND efet w=5800 l=10875
+ ad=0 pd=0 as=5.3824e+08 ps=118900 
M1304 R7_1 N0583 N0534 GND efet w=5800 l=11600
+ ad=5.4665e+08 pd=118900 as=0 ps=0 
M1305 N0923 R3_1 GND GND efet w=24650 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1306 GND R1_2 N0907 GND efet w=23925 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1307 GND N0868 N0535 GND efet w=58725 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1308 N0907 N0543 N0868 GND efet w=25375 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1309 N0867 N0565 N0923 GND efet w=29000 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1310 N0932 N0581 N0867 GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1311 GND R5_1 N0932 GND efet w=23200 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1312 N0533 N0598 R8_1 GND efet w=5800 l=13050
+ ad=0 pd=0 as=5.36138e+08 ps=118900 
M1313 N0977 N0645 N0881 GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1314 GND R12_1 N0977 GND efet w=21025 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1315 Vdd SC_A22_M22_CLK2 N0866 GND efet w=11600 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1316 Vdd Vdd N0531 GND efet w=8700 l=33350
+ ad=0 pd=0 as=0 ps=0 
M1317 Vdd Vdd N0532 GND efet w=8700 l=33350
+ ad=0 pd=0 as=0 ps=0 
M1318 Vdd SC_A22_M22_CLK2 N0880 GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1319 N0986 R14_1 GND GND efet w=26100 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1320 R10_1 N0619 N0533 GND efet w=5800 l=11600
+ ad=5.5506e+08 pd=124700 as=0 ps=0 
M1321 N0534 N0598 R9_1 GND efet w=5800 l=14500
+ ad=0 pd=0 as=5.40343e+08 ps=118900 
M1322 N0536 N0882 GND GND efet w=62350 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1323 N0882 WRAB0 N0864 GND efet w=13050 l=11600
+ ad=1.13325e+09 pd=220400 as=0 ps=0 
M1324 N0924 R3_2 GND GND efet w=23200 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1325 N0868 N0565 N0924 GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1326 N0933 N0581 N0868 GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1327 GND R5_2 N0933 GND efet w=23200 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1328 N0950 R7_1 GND GND efet w=23925 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1329 N0867 N0591 N0950 GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1330 N0959 N0616 N0867 GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1331 GND R9_1 N0959 GND efet w=23200 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1332 R11_1 N0619 N0534 GND efet w=7250 l=13050
+ ad=5.40343e+08 pd=121800 as=0 ps=0 
M1333 N0533 N0634 R12_1 GND efet w=5800 l=13050
+ ad=0 pd=0 as=5.44548e+08 ps=118900 
M1334 N0881 N0657 N0986 GND efet w=26100 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1335 R14_1 N0647 N0533 GND efet w=6525 l=13775
+ ad=5.9711e+08 pd=121800 as=0 ps=0 
M1336 N0534 N0634 R13_1 GND efet w=7250 l=13050
+ ad=0 pd=0 as=5.3824e+08 ps=118900 
M1337 N0969 R11_1 GND GND efet w=23200 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1338 N0867 N0632 N0969 GND efet w=25375 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1339 N0978 N0645 N0867 GND efet w=24650 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1340 GND R13_1 N0978 GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1341 N0951 R7_2 GND GND efet w=23200 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1342 N0535 N0529 R1_2 GND efet w=5800 l=12325
+ ad=0 pd=0 as=5.5506e+08 ps=121800 
M1343 R3_2 N0544 N0535 GND efet w=6525 l=12325
+ ad=5.4665e+08 pd=121800 as=0 ps=0 
M1344 N0536 N0529 R0_2 GND efet w=7975 l=10875
+ ad=0 pd=0 as=5.50855e+08 ps=121800 
M1345 R2_2 N0544 N0536 GND efet w=5800 l=11600
+ ad=5.4665e+08 pd=121800 as=0 ps=0 
M1346 N0908 N0543 N0882 GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1347 GND R0_2 N0908 GND efet w=23200 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1348 N0868 N0591 N0951 GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1349 N0960 N0616 N0868 GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1350 GND R9_2 N0960 GND efet w=23925 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1351 R15_1 N0647 N0534 GND efet w=7975 l=15225
+ ad=5.90802e+08 pd=124700 as=0 ps=0 
M1352 N0987 R15_1 GND GND efet w=27550 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1353 N0970 R11_2 GND GND efet w=23200 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1354 N0535 N0569 R5_2 GND efet w=5800 l=13050
+ ad=0 pd=0 as=5.40343e+08 ps=118900 
M1355 R7_2 N0583 N0535 GND efet w=7250 l=10875
+ ad=5.3824e+08 pd=118900 as=0 ps=0 
M1356 N0536 N0569 R4_2 GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.48753e+08 ps=124700 
M1357 GND R0_3 N0909 GND efet w=23925 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1358 Vdd Vdd N0392 GND efet w=7250 l=29000
+ ad=0 pd=0 as=0 ps=0 
M1359 Vdd __INH__X11_X31_CLK1 N0776 GND efet w=10875 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1360 N0500 M12_M22_CLK1__M11_M12_ D3 GND efet w=13050 l=11600
+ ad=1.66097e+09 pd=327700 as=0 ps=0 
M1361 D3 RRAB1 N0538 GND efet w=46400 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1362 N0537 RRAB0 D3 GND efet w=44950 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1363 N0842 PC3_1 GND GND efet w=23925 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1364 PC1_1 N0410 N0393 GND efet w=5800 l=11600
+ ad=5.2983e+08 pd=127600 as=0 ps=0 
M1365 N0780 N0444 N0842 GND efet w=25375 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1366 N0393 N0426 PC2_1 GND efet w=5800 l=10150
+ ad=0 pd=0 as=4.98293e+08 ps=124700 
M1367 PC3_1 N0439 N0393 GND efet w=5800 l=10150
+ ad=5.4665e+08 pd=121800 as=0 ps=0 
M1368 N0394 N0381 PC0_0 GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.34035e+08 ps=124700 
M1369 N0794 N0406 N0781 GND efet w=27550 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1370 GND PC0_0 N0794 GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1371 PC1_0 N0410 N0394 GND efet w=5800 l=11600
+ ad=5.27727e+08 pd=130500 as=0 ps=0 
M1372 N0815 PC1_0 GND GND efet w=23925 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1373 N0394 N0426 PC2_0 GND efet w=5800 l=10150
+ ad=0 pd=0 as=5.2142e+08 ps=133400 
M1374 GND N0777 N0395 GND efet w=68150 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1375 GND PC0_4 N0795 GND efet w=24650 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1376 N0764 WADB1 N0777 GND efet w=14500 l=11600
+ ad=0 pd=0 as=1.16058e+09 ps=232000 
M1377 D0 RADB1 N0395 GND efet w=43500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1378 N0396 RADB2 D0 GND efet w=48575 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1379 Vdd N0325 N0306 GND efet w=7250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1380 N0314 N0306 GND GND efet w=29000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1381 N0795 N0406 N0777 GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1382 N0781 N0424 N0815 GND efet w=25375 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1383 N0830 N0434 N0781 GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1384 GND PC2_0 N0830 GND efet w=23925 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1385 PC3_0 N0439 N0394 GND efet w=5800 l=10875
+ ad=5.48753e+08 pd=121800 as=0 ps=0 
M1386 N0843 PC3_0 GND GND efet w=22475 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1387 N0816 PC1_4 GND GND efet w=21750 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1388 N0777 N0424 N0816 GND efet w=25375 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1389 GND N0773 N0396 GND efet w=68875 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1390 N0773 WADB2 N0764 GND efet w=13050 l=11600
+ ad=1.37083e+09 pd=261000 as=0 ps=0 
M1391 N0395 N0381 PC0_4 GND efet w=6525 l=13775
+ ad=0 pd=0 as=5.27727e+08 ps=118900 
M1392 N0831 N0434 N0777 GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1393 GND PC2_4 N0831 GND efet w=23200 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1394 N0781 N0444 N0843 GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1395 Vdd __INH__X11_X31_CLK1 N0780 GND efet w=8700 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1396 N0883 WRAB0 N0865 GND efet w=13050 l=11600
+ ad=1.12273e+09 pd=214600 as=0 ps=0 
M1397 N0865 WRAB1 N0869 GND efet w=15225 l=10150
+ ad=0 pd=0 as=1.11432e+09 ps=214600 
M1398 GND N0883 N0537 GND efet w=59450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1399 N0909 N0543 N0883 GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1400 N0925 R2_2 GND GND efet w=23925 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1401 N0882 N0565 N0925 GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1402 N0934 N0581 N0882 GND efet w=24650 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1403 GND R4_2 N0934 GND efet w=25375 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1404 N0926 R2_3 GND GND efet w=23200 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1405 R6_2 N0583 N0536 GND efet w=5800 l=11600
+ ad=5.42445e+08 pd=118900 as=0 ps=0 
M1406 N0868 N0632 N0970 GND efet w=25375 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1407 N0979 N0645 N0868 GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1408 GND R13_2 N0979 GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1409 N0535 N0598 R9_2 GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.40343e+08 ps=121800 
M1410 R11_2 N0619 N0535 GND efet w=6525 l=13050
+ ad=5.4665e+08 pd=121800 as=0 ps=0 
M1411 N0867 N0657 N0987 GND efet w=25375 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1412 Vdd SC_A22_M22_CLK2 N0881 GND efet w=11600 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1413 Vdd Vdd N0533 GND efet w=7250 l=37700
+ ad=0 pd=0 as=0 ps=0 
M1414 Vdd Vdd N0534 GND efet w=7975 l=35525
+ ad=0 pd=0 as=0 ps=0 
M1415 Vdd SC_A22_M22_CLK2 N0867 GND efet w=12325 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1416 N0988 R15_2 GND GND efet w=27550 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1417 N0868 N0657 N0988 GND efet w=26100 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1418 N0536 N0598 R8_2 GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.5506e+08 ps=130500 
M1419 N0538 N0869 GND GND efet w=59450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1420 N0883 N0565 N0926 GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1421 N0935 N0581 N0883 GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1422 GND R4_3 N0935 GND efet w=26825 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1423 N0952 R6_2 GND GND efet w=23925 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1424 N0882 N0591 N0952 GND efet w=28275 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1425 N0961 N0616 N0882 GND efet w=29725 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1426 GND R8_2 N0961 GND efet w=25375 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1427 R10_2 N0619 N0536 GND efet w=5800 l=11600
+ ad=5.44548e+08 pd=121800 as=0 ps=0 
M1428 N0535 N0634 R13_2 GND efet w=5800 l=12325
+ ad=0 pd=0 as=5.36138e+08 ps=118900 
M1429 R15_2 N0647 N0535 GND efet w=6525 l=13775
+ ad=5.90802e+08 pd=124700 as=0 ps=0 
M1430 N0536 N0634 R12_2 GND efet w=6525 l=13775
+ ad=0 pd=0 as=5.69777e+08 ps=124700 
M1431 R14_2 N0647 N0536 GND efet w=6525 l=15225
+ ad=5.76085e+08 pd=127600 as=0 ps=0 
M1432 N0971 R10_2 GND GND efet w=24650 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1433 N0882 N0632 N0971 GND efet w=26825 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1434 N0980 N0645 N0882 GND efet w=29000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1435 N0953 R6_3 GND GND efet w=23200 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1436 N0537 N0529 R0_3 GND efet w=6525 l=13775
+ ad=0 pd=0 as=5.5506e+08 ps=121800 
M1437 R2_3 N0544 N0537 GND efet w=4350 l=12325
+ ad=5.50855e+08 pd=121800 as=0 ps=0 
M1438 N0538 N0529 R1_3 GND efet w=7250 l=11600
+ ad=0 pd=0 as=5.4665e+08 ps=121800 
M1439 R3_3 N0544 N0538 GND efet w=5800 l=11600
+ ad=5.40343e+08 pd=121800 as=0 ps=0 
M1440 N0910 N0543 N0869 GND efet w=24650 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1441 GND R1_3 N0910 GND efet w=23200 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1442 N0537 N0569 R4_3 GND efet w=7250 l=11600
+ ad=0 pd=0 as=5.69777e+08 ps=133400 
M1443 N0883 N0591 N0953 GND efet w=26825 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1444 N0962 N0616 N0883 GND efet w=26825 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1445 GND R8_3 N0962 GND efet w=26100 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1446 GND R12_2 N0980 GND efet w=21025 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1447 N0972 R10_3 GND GND efet w=24650 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1448 R6_3 N0583 N0537 GND efet w=6525 l=13775
+ ad=5.44548e+08 pd=121800 as=0 ps=0 
M1449 N0538 N0569 R5_3 GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.2142e+08 ps=130500 
M1450 Vdd Vdd N0393 GND efet w=5800 l=30450
+ ad=0 pd=0 as=0 ps=0 
M1451 GND N0461 N0469 GND efet w=13050 l=13050
+ ad=0 pd=0 as=1.66308e+09 ps=324800 
M1452 N0469 Vdd Vdd GND efet w=8700 l=65250
+ ad=0 pd=0 as=0 ps=0 
M1453 N0461 N0469 GND GND efet w=11600 l=11600
+ ad=1.4255e+09 pd=295800 as=0 ps=0 
M1454 N0927 R3_3 GND GND efet w=23925 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1455 N0869 N0565 N0927 GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1456 N0936 N0581 N0869 GND efet w=27550 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1457 GND R5_3 N0936 GND efet w=27550 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1458 R7_3 N0583 N0538 GND efet w=5800 l=11600
+ ad=5.36138e+08 pd=118900 as=0 ps=0 
M1459 N0883 N0632 N0972 GND efet w=26100 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1460 N0981 N0645 N0883 GND efet w=31175 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1461 GND R12_3 N0981 GND efet w=22475 l=17400
+ ad=0 pd=0 as=0 ps=0 
M1462 N0989 R14_2 GND GND efet w=29725 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1463 N0882 N0657 N0989 GND efet w=27550 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1464 Vdd SC_A22_M22_CLK2 N0868 GND efet w=14500 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1465 Vdd Vdd N0535 GND efet w=8700 l=34075
+ ad=0 pd=0 as=0 ps=0 
M1466 Vdd Vdd N0536 GND efet w=7975 l=32625
+ ad=0 pd=0 as=0 ps=0 
M1467 Vdd SC_A22_M22_CLK2 N0882 GND efet w=11600 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1468 N0990 R14_3 GND GND efet w=29000 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1469 N0883 N0657 N0990 GND efet w=29000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1470 N0537 N0598 R8_3 GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.76085e+08 ps=124700 
M1471 R10_3 N0619 N0537 GND efet w=5800 l=13775
+ ad=5.52958e+08 pd=127600 as=0 ps=0 
M1472 N0538 N0598 R9_3 GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.5506e+08 ps=130500 
M1473 N0954 R7_3 GND GND efet w=23925 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1474 N0869 N0591 N0954 GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1475 N0963 N0616 N0869 GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1476 GND R9_3 N0963 GND efet w=25375 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1477 R11_3 N0619 N0538 GND efet w=5800 l=11600
+ ad=5.67675e+08 pd=130500 as=0 ps=0 
M1478 N0973 R11_3 GND GND efet w=26825 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1479 N0537 N0634 R12_3 GND efet w=5800 l=11600
+ ad=0 pd=0 as=6.01315e+08 ps=124700 
M1480 Vdd SC_A22_M22_CLK2 N0883 GND efet w=11600 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1481 R14_3 N0647 N0537 GND efet w=5800 l=13050
+ ad=5.90802e+08 pd=139200 as=0 ps=0 
M1482 N0538 N0634 R13_3 GND efet w=5800 l=13050
+ ad=0 pd=0 as=5.78188e+08 ps=133400 
M1483 R15_3 N0647 N0538 GND efet w=7250 l=14500
+ ad=6.03417e+08 pd=127600 as=0 ps=0 
M1484 N0869 N0632 N0973 GND efet w=26100 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1485 N0982 N0645 N0869 GND efet w=26100 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1486 GND R13_3 N0982 GND efet w=27550 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1487 Vdd Vdd N0537 GND efet w=8700 l=34075
+ ad=0 pd=0 as=0 ps=0 
M1488 GND GND clk2 GND efet w=118175 l=13775
+ ad=0 pd=0 as=-8.51217e+08 ps=1.24294e+07 
M1489 GND GND clk1 GND efet w=113100 l=13050
+ ad=0 pd=0 as=1.86634e+09 ps=6.6033e+06 
M1490 Vdd Vdd N0538 GND efet w=8700 l=34075
+ ad=0 pd=0 as=0 ps=0 
M1491 N0991 R15_3 GND GND efet w=26100 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1492 N0869 N0657 N0991 GND efet w=26825 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1493 Vdd SC_A22_M22_CLK2 N0869 GND efet w=11600 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1494 Vdd Vdd N0394 GND efet w=5800 l=29000
+ ad=0 pd=0 as=0 ps=0 
M1495 Vdd Vdd N0461 GND efet w=5800 l=65250
+ ad=0 pd=0 as=0 ps=0 
M1496 ADDR_RFSH_1 Vdd Vdd GND efet w=8700 l=66700
+ ad=0 pd=0 as=0 ps=0 
M1497 GND N0461 ADDR_RFSH_1 GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1498 N0453 N0469 GND GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1499 GND N0902 N0543 GND efet w=14500 l=11600
+ ad=0 pd=0 as=1.27456e+09 ps=1.0034e+06 
M1500 GND N0902 N0529 GND efet w=11600 l=11600
+ ad=0 pd=0 as=1.15051e+09 ps=1.0179e+06 
M1501 GND N0919 N0544 GND efet w=11600 l=11600
+ ad=0 pd=0 as=1.1442e+09 ps=997600 
M1502 GND N0919 N0565 GND efet w=14500 l=11600
+ ad=0 pd=0 as=1.15682e+09 ps=1.0295e+06 
M1503 Vdd Vdd N0453 GND efet w=9425 l=65975
+ ad=0 pd=0 as=0 ps=0 
M1504 Vdd __INH__X11_X31_CLK1 N0781 GND efet w=9425 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1505 N0902 Vdd Vdd GND efet w=6525 l=61625
+ ad=1.15638e+09 pd=229100 as=0 ps=0 
M1506 N0543 N0530 __POC__CLK2_SC_A32_X12_ GND efet w=16675 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1507 N0529 N0530 CLK2_SC_A12_M12_ GND efet w=13775 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1508 N0544 N0545 CLK2_SC_A12_M12_ GND efet w=12325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1509 N0565 N0545 __POC__CLK2_SC_A32_X12_ GND efet w=16675 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1510 N0844 PC3_4 GND GND efet w=22475 l=18125
+ ad=0 pd=0 as=0 ps=0 
M1511 ADDR_RFSH_1 N0455 N0489 GND efet w=8700 l=10150
+ ad=0 pd=0 as=8.30487e+08 ps=185600 
M1512 N0453 N0455 N0454 GND efet w=8700 l=13050
+ ad=0 pd=0 as=1.08489e+09 ps=229100 
M1513 PC1_4 N0410 N0395 GND efet w=6525 l=12325
+ ad=5.48753e+08 pd=121800 as=0 ps=0 
M1514 N0396 N0381 PC0_8 GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.2142e+08 ps=116000 
M1515 N0796 N0406 N0773 GND efet w=27550 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1516 Vdd Vdd N0314 GND efet w=7250 l=65250
+ ad=0 pd=0 as=0 ps=0 
M1517 GND A32 N0712 GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1518 N0314 clk2 N0315 GND efet w=13050 l=14500
+ ad=0 pd=0 as=6.3916e+08 ps=136300 
M1519 cm_rom N0717 Vdd GND efet w=417600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1520 GND N0737 cm_rom GND efet w=607550 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1521 N0712 A22 GND GND efet w=26825 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1522 N0325 Vdd clk1 GND efet w=34800 l=11600
+ ad=9.0872e+08 pd=983100 as=0 ps=0 
M1523 Vdd Vdd WADB1 GND efet w=5800 l=27550
+ ad=0 pd=0 as=-8.52735e+08 ps=1.421e+06 
M1524 GND A12 N0711 GND efet w=13050 l=12325
+ ad=0 pd=0 as=9.62945e+08 ps=217500 
M1525 N0316 N0315 GND GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1526 WADB0 Vdd Vdd GND efet w=7250 l=27550
+ ad=-9.43142e+08 pd=1.4268e+06 as=0 ps=0 
M1527 GND N0300 WADB0 GND efet w=29000 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1528 Vdd Vdd N0316 GND efet w=6525 l=51475
+ ad=0 pd=0 as=0 ps=0 
M1529 N0711 Vdd Vdd GND efet w=6525 l=67425
+ ad=0 pd=0 as=0 ps=0 
M1530 N0317 clk1 N0316 GND efet w=8700 l=11600
+ ad=5.40343e+08 pd=118900 as=0 ps=0 
M1531 GND N0326 WADB0 GND efet w=36250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1532 GND PC0_8 N0796 GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1533 PC1_8 N0410 N0396 GND efet w=5800 l=11600
+ ad=5.3824e+08 pd=133400 as=0 ps=0 
M1534 N0777 N0444 N0844 GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1535 N0395 N0426 PC2_4 GND efet w=6525 l=10875
+ ad=0 pd=0 as=5.42445e+08 ps=124700 
M1536 PC3_4 N0439 N0395 GND efet w=5800 l=10150
+ ad=5.52958e+08 pd=121800 as=0 ps=0 
M1537 N0396 N0426 PC2_8 GND efet w=5800 l=10150
+ ad=0 pd=0 as=5.3824e+08 ps=127600 
M1538 PC3_8 N0439 N0396 GND efet w=5800 l=10150
+ ad=5.57162e+08 pd=121800 as=0 ps=0 
M1539 N0817 PC1_8 GND GND efet w=26100 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1540 N0773 N0424 N0817 GND efet w=27550 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1541 N0832 N0434 N0773 GND efet w=25375 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1542 WADB2 Vdd Vdd GND efet w=7975 l=31175
+ ad=-5.3736e+08 pd=1.4471e+06 as=0 ps=0 
M1543 GND PC2_8 N0832 GND efet w=25375 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1544 N0845 PC3_8 GND GND efet w=23925 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1545 N0773 N0444 N0845 GND efet w=26825 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1546 Vdd __INH__X11_X31_CLK1 N0777 GND efet w=8700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1547 N0488 N0463 N0469 GND efet w=21750 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1548 Vdd Vdd N0395 GND efet w=6525 l=32625
+ ad=0 pd=0 as=0 ps=0 
M1549 GND N0489 N0488 GND efet w=34075 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1550 N0462 N0454 GND GND efet w=34800 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1551 N0461 N0463 N0462 GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1552 Vdd Vdd N0396 GND efet w=6525 l=31175
+ ad=0 pd=0 as=0 ps=0 
M1553 GND N0928 N0581 GND efet w=14500 l=10150
+ ad=0 pd=0 as=1.18415e+09 ps=1.0092e+06 
M1554 GND N0928 N0569 GND efet w=11600 l=10150
+ ad=0 pd=0 as=1.16102e+09 ps=1.0382e+06 
M1555 GND N0938 N0583 GND efet w=13050 l=10150
+ ad=0 pd=0 as=1.12738e+09 ps=1.015e+06 
M1556 GND N0938 N0591 GND efet w=15950 l=10150
+ ad=0 pd=0 as=1.35445e+09 ps=1.0266e+06 
M1557 GND N0955 N0616 GND efet w=13775 l=10875
+ ad=0 pd=0 as=1.28297e+09 ps=1.0266e+06 
M1558 N0581 N0570 __POC__CLK2_SC_A32_X12_ GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1559 N0569 N0570 CLK2_SC_A12_M12_ GND efet w=12325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1560 N0583 N0584 CLK2_SC_A12_M12_ GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1561 N0591 N0584 __POC__CLK2_SC_A32_X12_ GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1562 GND N0530 N0902 GND efet w=11600 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1563 N0919 N0545 GND GND efet w=10150 l=11600
+ ad=1.58739e+09 pd=324800 as=0 ps=0 
M1564 GND N0570 N0928 GND efet w=10875 l=12325
+ ad=0 pd=0 as=1.54113e+09 ps=330600 
M1565 N0938 N0584 GND GND efet w=10150 l=13050
+ ad=1.6e+09 pd=330600 as=0 ps=0 
M1566 GND N0955 N0598 GND efet w=13050 l=10875
+ ad=0 pd=0 as=1.38389e+09 ps=1.0063e+06 
M1567 GND N0965 N0619 GND efet w=11600 l=11600
+ ad=0 pd=0 as=1.24302e+09 ps=1.0179e+06 
M1568 GND N0965 N0632 GND efet w=13050 l=12325
+ ad=0 pd=0 as=1.42594e+09 ps=1.0121e+06 
M1569 N0616 N0599 __POC__CLK2_SC_A32_X12_ GND efet w=14500 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1570 CLK2_SC_A12_M12_ N0599 N0598 GND efet w=12325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1571 N0619 N0620 CLK2_SC_A12_M12_ GND efet w=12325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1572 N0632 N0620 __POC__CLK2_SC_A32_X12_ GND efet w=13050 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1573 GND N0599 N0955 GND efet w=12325 l=12325
+ ad=0 pd=0 as=1.6021e+09 ps=342200 
M1574 RRAB1 S00557 RRAB1 GND efet w=77575 l=6525
+ ad=6.79548e+08 pd=881600 as=0 ps=0 
M1575 RRAB1 S00557 Vdd GND efet w=10150 l=23200
+ ad=0 pd=0 as=0 ps=0 
M1576 S00557 Vdd Vdd GND efet w=6525 l=13775
+ ad=-1.77617e+09 pd=304500 as=0 ps=0 
M1577 Vdd __INH__X11_X31_CLK1 N0773 GND efet w=10150 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1578 N0463 Vdd Vdd GND efet w=6525 l=71775
+ ad=-1.82032e+09 pd=466900 as=0 ps=0 
M1579 GND N0455 N0463 GND efet w=11600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1580 N0455 N0463 GND GND efet w=13050 l=11600
+ ad=-1.13095e+08 pd=797500 as=0 ps=0 
M1581 N0919 Vdd Vdd GND efet w=6525 l=45675
+ ad=0 pd=0 as=0 ps=0 
M1582 Vdd Vdd N0928 GND efet w=7975 l=51475
+ ad=0 pd=0 as=0 ps=0 
M1583 N0965 N0620 GND GND efet w=11600 l=13050
+ ad=1.67359e+09 pd=319000 as=0 ps=0 
M1584 GND N0974 N0645 GND efet w=14500 l=11600
+ ad=0 pd=0 as=1.44906e+09 ps=1.0353e+06 
M1585 GND N0974 N0634 GND efet w=11600 l=11600
+ ad=0 pd=0 as=1.47429e+09 ps=1.0208e+06 
M1586 GND N0983 N0647 GND efet w=11600 l=11600
+ ad=0 pd=0 as=1.61096e+09 ps=1.0092e+06 
M1587 GND N0983 N0657 GND efet w=14500 l=11600
+ ad=0 pd=0 as=1.71818e+09 ps=1.0324e+06 
M1588 N0645 N0635 __POC__CLK2_SC_A32_X12_ GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1589 N0634 N0635 CLK2_SC_A12_M12_ GND efet w=12325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1590 N0647 N0648 CLK2_SC_A12_M12_ GND efet w=12325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1591 N0657 N0648 __POC__CLK2_SC_A32_X12_ GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1592 N0938 Vdd Vdd GND efet w=5800 l=47850
+ ad=0 pd=0 as=0 ps=0 
M1593 Vdd Vdd N0955 GND efet w=6525 l=52925
+ ad=0 pd=0 as=0 ps=0 
M1594 GND N0635 N0974 GND efet w=10150 l=13050
+ ad=0 pd=0 as=1.67359e+09 ps=316100 
M1595 N0983 N0648 GND GND efet w=10150 l=13050
+ ad=1.69251e+09 pd=327700 as=0 ps=0 
M1596 Vdd Vdd N0613 GND efet w=13050 l=45675
+ ad=0 pd=0 as=4.14633e+08 ps=936700 
M1597 N0965 Vdd Vdd GND efet w=6525 l=48575
+ ad=0 pd=0 as=0 ps=0 
M1598 Vdd Vdd N0974 GND efet w=5800 l=47850
+ ad=0 pd=0 as=0 ps=0 
M1599 N0983 Vdd Vdd GND efet w=5800 l=47850
+ ad=0 pd=0 as=0 ps=0 
M1600 N0539 N0540 GND GND efet w=27550 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1601 Vdd Vdd N0540 GND efet w=7250 l=29000
+ ad=0 pd=0 as=2.13193e+09 ps=426300 
M1602 Vdd Vdd N0455 GND efet w=6525 l=68875
+ ad=0 pd=0 as=0 ps=0 
M1603 ADDR_RFSH_0 Vdd Vdd GND efet w=9425 l=73950
+ ad=0 pd=0 as=0 ps=0 
M1604 GND N0455 ADDR_RFSH_0 GND efet w=13775 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1605 N0503 N0463 GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1606 Vdd Vdd N0503 GND efet w=8700 l=66700
+ ad=0 pd=0 as=0 ps=0 
M1607 S00564 Vdd Vdd GND efet w=6525 l=13775
+ ad=-1.83925e+09 pd=313200 as=0 ps=0 
M1608 RRAB0 S00564 RRAB0 GND efet w=57275 l=15225
+ ad=7.46828e+08 pd=887400 as=0 ps=0 
M1609 RRAB0 S00564 Vdd GND efet w=7250 l=21750
+ ad=0 pd=0 as=0 ps=0 
M1610 WADB1 N0318 GND GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1611 GND N0304 WADB2 GND efet w=29000 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1612 GND N0300 WADB1 GND efet w=27550 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1613 WADB2 N0300 GND GND efet w=29725 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1614 GND N0783 N0406 GND efet w=15950 l=10150
+ ad=0 pd=0 as=-6.59305e+08 ps=1.4761e+06 
M1615 GND N0783 N0381 GND efet w=11600 l=10150
+ ad=0 pd=0 as=-7.60225e+08 ps=1.5283e+06 
M1616 GND N0804 N0410 GND efet w=11600 l=11600
+ ad=0 pd=0 as=-6.3828e+08 ps=1.4877e+06 
M1617 GND N0804 N0424 GND efet w=15950 l=10150
+ ad=0 pd=0 as=-8.92682e+08 ps=1.4732e+06 
M1618 N0406 N0382 __POC_CLK2_X12_X32__INH GND efet w=15950 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1619 N0381 N0382 ___SC__JIN_FIN__CLK1_M11_X21_INH_ GND efet w=10150 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1620 N0410 N0411 ___SC__JIN_FIN__CLK1_M11_X21_INH_ GND efet w=12325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1621 N0424 N0411 __POC_CLK2_X12_X32__INH GND efet w=15950 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1622 N0737 Vdd Vdd GND efet w=9425 l=13775
+ ad=-1.48769e+09 pd=1.4355e+06 as=0 ps=0 
M1623 N0711 N0732 N0712 GND efet w=23200 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1624 GND N0820 N0434 GND efet w=15950 l=10150
+ ad=0 pd=0 as=-8.63247e+08 ps=1.4616e+06 
M1625 N0426 N0820 GND GND efet w=11600 l=11600
+ ad=-8.08582e+08 pd=1.5051e+06 as=0 ps=0 
M1626 GND N0833 N0439 GND efet w=11600 l=11600
+ ad=0 pd=0 as=-9.59962e+08 ps=1.4848e+06 
M1627 N0444 N0833 GND GND efet w=15950 l=13050
+ ad=-6.48792e+08 pd=1.4616e+06 as=0 ps=0 
M1628 ADDR_RFSH_0 clk1 N0519 GND efet w=7250 l=11600
+ ad=0 pd=0 as=7.37977e+08 ps=156600 
M1629 N0545 N0540 GND GND efet w=14500 l=10150
+ ad=1.79553e+09 pd=377000 as=0 ps=0 
M1630 N0570 N0540 GND GND efet w=14500 l=11600
+ ad=2.06886e+09 pd=414700 as=0 ps=0 
M1631 N0584 N0540 GND GND efet w=13775 l=14500
+ ad=1.91117e+09 pd=377000 as=0 ps=0 
M1632 N0599 N0613 GND GND efet w=13775 l=13775
+ ad=1.74507e+09 pd=388600 as=0 ps=0 
M1633 GND N0613 N0540 GND efet w=32625 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1634 N0620 N0613 GND GND efet w=15225 l=12325
+ ad=1.94902e+09 pd=403100 as=0 ps=0 
M1635 N0635 N0613 GND GND efet w=13775 l=13775
+ ad=1.96584e+09 pd=388600 as=0 ps=0 
M1636 N0648 N0613 GND GND efet w=16675 l=13050
+ ad=1.83548e+09 pd=359600 as=0 ps=0 
M1637 N0613 N0646 GND GND efet w=52925 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1638 N0539 N0541 GND GND efet w=27550 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1639 N0545 N0541 GND GND efet w=14500 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1640 GND N0541 N0599 GND efet w=13775 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1641 GND N0541 N0620 GND efet w=13775 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1642 N0570 N0577 GND GND efet w=13775 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1643 GND N0542 N0539 GND efet w=29000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1644 N0584 N0577 GND GND efet w=13775 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1645 N0503 clk1 N0504 GND efet w=7250 l=13050
+ ad=0 pd=0 as=9.5033e+08 ps=200100 
M1646 N0635 N0577 GND GND efet w=13050 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1647 N0648 N0577 GND GND efet w=15950 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1648 Vdd Vdd N0541 GND efet w=9425 l=38425
+ ad=0 pd=0 as=-2.0028e+09 ps=1.3311e+06 
M1649 N0570 N0542 GND GND efet w=14500 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1650 N0434 N0427 __POC_CLK2_X12_X32__INH GND efet w=15950 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1651 N0426 N0427 ___SC__JIN_FIN__CLK1_M11_X21_INH_ GND efet w=10875 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1652 N0439 N0440 ___SC__JIN_FIN__CLK1_M11_X21_INH_ GND efet w=11600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1653 N0444 N0440 __POC_CLK2_X12_X32__INH GND efet w=18125 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1654 GND N0519 N0518 GND efet w=40600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1655 GND N0382 N0783 GND efet w=12325 l=12325
+ ad=0 pd=0 as=1.6799e+09 ps=353800 
M1656 N0804 N0411 GND GND efet w=11600 l=11600
+ ad=1.66938e+09 pd=350900 as=0 ps=0 
M1657 N0518 __INH__X32_CLK2 N0463 GND efet w=21750 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1658 N0508 N0504 GND GND efet w=38425 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1659 GND N0542 N0599 GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1660 GND N0542 N0635 GND efet w=13050 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1661 N0541 N0577 GND GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1662 N0577 N0617 GND GND efet w=52200 l=13050
+ ad=1.06431e+09 pd=1.0005e+06 as=0 ps=0 
M1663 N0455 __INH__X32_CLK2 N0508 GND efet w=19575 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1664 N0539 __FIN_X12_ N0530 GND efet w=41325 l=12325
+ ad=0 pd=0 as=1.65887e+09 ps=345100 
M1665 N0561 Vdd Vdd GND efet w=8700 l=40600
+ ad=1.93895e+09 pd=1.1948e+06 as=0 ps=0 
M1666 GND __FIN_X12_ N0561 GND efet w=29000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1667 Vdd Vdd N0833 GND efet w=5800 l=60900
+ ad=0 pd=0 as=1.38975e+09 ps=281300 
M1668 GND N0427 N0820 GND efet w=11600 l=10875
+ ad=0 pd=0 as=1.59159e+09 ps=336400 
M1669 N0833 N0440 GND GND efet w=11600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1670 N0732 N0317 GND GND efet w=19575 l=12325
+ ad=1.65467e+09 pd=356700 as=0 ps=0 
M1671 Vdd Vdd N0732 GND efet w=8700 l=65250
+ ad=0 pd=0 as=0 ps=0 
M1672 GND N0711 N0307 GND efet w=13775 l=11600
+ ad=0 pd=0 as=-1.89812e+09 ps=452400 
M1673 GND N0416 RADB0 GND efet w=43500 l=13050
+ ad=0 pd=0 as=-1.41831e+09 ps=1.2963e+06 
M1674 RADB2 Vdd Vdd GND efet w=7975 l=23200
+ ad=-2.5983e+08 pd=1.5921e+06 as=0 ps=0 
M1675 N0300 clk2 GND GND efet w=26100 l=13050
+ ad=-1.82663e+09 pd=495900 as=0 ps=0 
M1676 N0307 Vdd Vdd GND efet w=10150 l=50750
+ ad=0 pd=0 as=0 ps=0 
M1677 GND clk1 N0307 GND efet w=15950 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1678 Vdd Vdd N0300 GND efet w=6525 l=29725
+ ad=0 pd=0 as=0 ps=0 
M1679 GND N0717 N0737 GND efet w=94250 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1680 M12_M22_CLK1__M11_M12_ N0710 Vdd GND efet w=23925 l=15225
+ ad=-1.84722e+09 pd=1.2586e+06 as=0 ps=0 
M1681 GND N0708 M12_M22_CLK1__M11_M12_ GND efet w=20300 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1682 N0710 S00609 N0710 GND efet w=57275 l=14500
+ ad=6.8121e+08 pd=145000 as=0 ps=0 
M1683 S00609 Vdd Vdd GND efet w=7250 l=11600
+ ad=-2.01165e+09 pd=290000 as=0 ps=0 
M1684 GND N0708 N0710 GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1685 N0402 Vdd Vdd GND efet w=7975 l=60900
+ ad=0 pd=0 as=0 ps=0 
M1686 GND X32 N0402 GND efet w=15950 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1687 RADB1 Vdd Vdd GND efet w=7975 l=26825
+ ad=-2.32497e+08 pd=1.4993e+06 as=0 ps=0 
M1688 RADB0 Vdd Vdd GND efet w=8700 l=21750
+ ad=0 pd=0 as=0 ps=0 
M1689 RADB1 clk2 GND GND efet w=50750 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1690 GND N0384 RADB1 GND efet w=42775 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1691 RADB2 clk2 GND GND efet w=53650 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1692 GND N0374 RADB2 GND efet w=50025 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1693 Vdd Vdd N0783 GND efet w=5800 l=62350
+ ad=0 pd=0 as=0 ps=0 
M1694 Vdd Vdd N0804 GND efet w=6525 l=50025
+ ad=0 pd=0 as=0 ps=0 
M1695 N0820 Vdd Vdd GND efet w=5800 l=52200
+ ad=0 pd=0 as=0 ps=0 
M1696 N0400 N0409 GND GND efet w=23925 l=10875
+ ad=-2.32937e+08 pd=870000 as=0 ps=0 
M1697 GND N0560 N0545 GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1698 N0584 N0560 GND GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1699 N0620 N0560 GND GND efet w=14500 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1700 N0648 N0560 GND GND efet w=14500 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1701 N0545 N0561 GND GND efet w=14500 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1702 N0570 N0561 GND GND efet w=15225 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1703 N0584 N0561 GND GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1704 N0599 N0561 GND GND efet w=16675 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1705 N0620 N0561 GND GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1706 N0635 N0561 GND GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1707 N0648 N0561 GND GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1708 N0545 S00579 N0545 GND efet w=58725 l=29725
+ ad=0 pd=0 as=0 ps=0 
M1709 Vdd Vdd N0400 GND efet w=8700 l=65250
+ ad=0 pd=0 as=0 ps=0 
M1710 N0530 S00578 N0530 GND efet w=15950 l=50750
+ ad=0 pd=0 as=0 ps=0 
M1711 N0427 N0400 GND GND efet w=11600 l=13050
+ ad=1.49488e+09 pd=307400 as=0 ps=0 
M1712 N0475 Vdd Vdd GND efet w=7250 l=65250
+ ad=1.5958e+09 pd=319000 as=0 ps=0 
M1713 GND N0464 N0475 GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1714 ADDR_PTR_1 Vdd Vdd GND efet w=8700 l=68150
+ ad=0 pd=0 as=0 ps=0 
M1715 GND N0464 ADDR_PTR_1 GND efet w=15225 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1716 N0464 N0475 GND GND efet w=13050 l=11600
+ ad=1.48437e+09 pd=301600 as=0 ps=0 
M1717 Vdd Vdd N0464 GND efet w=6525 l=67425
+ ad=0 pd=0 as=0 ps=0 
M1718 N0457 N0475 GND GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1719 Vdd Vdd N0457 GND efet w=8700 l=66700
+ ad=0 pd=0 as=0 ps=0 
M1720 N0440 N0409 GND GND efet w=19575 l=12325
+ ad=1.5979e+09 pd=316100 as=0 ps=0 
M1721 ADDR_PTR_1 N0459 N0492 GND efet w=8700 l=11600
+ ad=0 pd=0 as=7.4008e+08 ps=153700 
M1722 N0457 N0459 N0458 GND efet w=9425 l=12325
+ ad=0 pd=0 as=9.48228e+08 ps=194300 
M1723 N0402 clk2 N0416 GND efet w=7250 l=13050
+ ad=0 pd=0 as=8.01052e+08 ps=162400 
M1724 N0384 clk2 N0379 GND efet w=7250 l=11600
+ ad=7.94745e+08 pd=162400 as=0 ps=0 
M1725 N0374 clk2 N0365 GND efet w=7975 l=13775
+ ad=8.19975e+08 pd=176900 as=0 ps=0 
M1726 N0710 S00609 Vdd GND efet w=7975 l=37700
+ ad=0 pd=0 as=0 ps=0 
M1727 N0379 A12 GND GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1728 GND A22 N0365 GND efet w=15950 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1729 Vdd Vdd N0365 GND efet w=9425 l=55825
+ ad=0 pd=0 as=0 ps=0 
M1730 Vdd Vdd N0708 GND efet w=8700 l=34800
+ ad=0 pd=0 as=1.1816e+09 ps=255200 
M1731 N0708 clk1 N0709 GND efet w=48575 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1732 N0709 N0278 GND GND efet w=44225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1733 Vdd Vdd N0279 GND efet w=6525 l=41325
+ ad=0 pd=0 as=0 ps=0 
M1734 GND M12 N0708 GND efet w=22475 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1735 N0708 M22 GND GND efet w=23200 l=8700
+ ad=0 pd=0 as=0 ps=0 
M1736 Vdd Vdd N0379 GND efet w=6525 l=52925
+ ad=0 pd=0 as=0 ps=0 
M1737 N0278 clk2 N0279 GND efet w=14500 l=11600
+ ad=7.9895e+08 pd=162400 as=0 ps=0 
M1738 GND M12 N0279 GND efet w=21025 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1739 RADB0 clk2 GND GND efet w=43500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1740 N0382 N0400 GND GND efet w=13050 l=10150
+ ad=-2.09996e+09 pd=452400 as=0 ps=0 
M1741 N0411 N0409 GND GND efet w=20300 l=10150
+ ad=1.81025e+09 pd=368300 as=0 ps=0 
M1742 N0382 N0401 GND GND efet w=12325 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1743 N0411 N0401 GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1744 GND N0420 N0427 GND efet w=20300 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1745 N0440 N0420 GND GND efet w=20300 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1746 N0382 S00598 N0382 GND efet w=30450 l=35525
+ ad=0 pd=0 as=0 ps=0 
M1747 GND A32 N0279 GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1748 Vdd Vdd N0304 GND efet w=7250 l=69600
+ ad=0 pd=0 as=1.77872e+09 ps=356700 
M1749 N0382 S00598 Vdd GND efet w=7250 l=56550
+ ad=0 pd=0 as=0 ps=0 
M1750 N0411 S00599 N0411 GND efet w=60900 l=30450
+ ad=0 pd=0 as=0 ps=0 
M1751 N0427 S00600 N0427 GND efet w=29725 l=60175
+ ad=0 pd=0 as=0 ps=0 
M1752 GND N0492 N0491 GND efet w=39150 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1753 N0440 S00601 N0440 GND efet w=62350 l=31900
+ ad=0 pd=0 as=0 ps=0 
M1754 N0411 S00599 Vdd GND efet w=7250 l=55100
+ ad=0 pd=0 as=0 ps=0 
M1755 N0427 S00600 Vdd GND efet w=7250 l=56550
+ ad=0 pd=0 as=0 ps=0 
M1756 N0401 N0420 GND GND efet w=24650 l=11600
+ ad=-1.36829e+09 pd=661200 as=0 ps=0 
M1757 Vdd Vdd N0401 GND efet w=8700 l=66700
+ ad=0 pd=0 as=0 ps=0 
M1758 N0491 N0466 N0475 GND efet w=21750 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1759 N0465 N0458 GND GND efet w=39150 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1760 N0464 N0466 N0465 GND efet w=19575 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1761 N0530 S00578 Vdd GND efet w=10150 l=55825
+ ad=0 pd=0 as=0 ps=0 
M1762 N0570 S00580 N0570 GND efet w=28275 l=31175
+ ad=0 pd=0 as=0 ps=0 
M1763 N0545 S00579 Vdd GND efet w=7975 l=60175
+ ad=0 pd=0 as=0 ps=0 
M1764 N0570 S00580 Vdd GND efet w=7250 l=56550
+ ad=0 pd=0 as=0 ps=0 
M1765 N0584 S00581 N0584 GND efet w=29725 l=55100
+ ad=0 pd=0 as=0 ps=0 
M1766 N0599 S00582 N0599 GND efet w=29725 l=52925
+ ad=0 pd=0 as=0 ps=0 
M1767 N0620 S00583 N0620 GND efet w=29725 l=52925
+ ad=0 pd=0 as=0 ps=0 
M1768 N0635 S00584 N0635 GND efet w=30450 l=31175
+ ad=0 pd=0 as=0 ps=0 
M1769 N0584 S00581 Vdd GND efet w=7250 l=56550
+ ad=0 pd=0 as=0 ps=0 
M1770 N0599 S00582 Vdd GND efet w=8700 l=59450
+ ad=0 pd=0 as=0 ps=0 
M1771 N0620 S00583 Vdd GND efet w=9425 l=54375
+ ad=0 pd=0 as=0 ps=0 
M1772 N0635 S00584 Vdd GND efet w=9425 l=55825
+ ad=0 pd=0 as=0 ps=0 
M1773 Vdd Vdd N0577 GND efet w=8700 l=37700
+ ad=0 pd=0 as=0 ps=0 
M1774 Vdd Vdd N0542 GND efet w=11600 l=42775
+ ad=0 pd=0 as=-1.8367e+09 ps=1.2644e+06 
M1775 N0648 S00585 N0648 GND efet w=30450 l=31175
+ ad=0 pd=0 as=0 ps=0 
M1776 N0542 N0560 GND GND efet w=26100 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1777 N0560 N0582 GND GND efet w=48575 l=10875
+ ad=1.40912e+09 pd=1.1484e+06 as=0 ps=0 
M1778 Vdd Vdd N0560 GND efet w=10150 l=44225
+ ad=0 pd=0 as=0 ps=0 
M1779 N0648 S00585 Vdd GND efet w=7250 l=53650
+ ad=0 pd=0 as=0 ps=0 
M1780 D1 SC_M22_CLK2 N0582 GND efet w=8700 l=13050
+ ad=0 pd=0 as=1.35191e+09 ps=252300 
M1781 D2 SC_M22_CLK2 N0617 GND efet w=7250 l=13050
+ ad=0 pd=0 as=1.15427e+09 ps=214600 
M1782 S00578 Vdd Vdd GND efet w=8700 l=11600
+ ad=-1.1286e+09 pd=319000 as=0 ps=0 
M1783 S00579 Vdd Vdd GND efet w=8700 l=12325
+ ad=-1.16434e+09 pd=301600 as=0 ps=0 
M1784 S00580 Vdd Vdd GND efet w=10150 l=10150
+ ad=-1.19588e+09 pd=304500 as=0 ps=0 
M1785 S00581 Vdd Vdd GND efet w=10150 l=10150
+ ad=-1.17906e+09 pd=298700 as=0 ps=0 
M1786 S00582 Vdd Vdd GND efet w=8700 l=10150
+ ad=-1.13281e+09 pd=307400 as=0 ps=0 
M1787 S00583 Vdd Vdd GND efet w=9425 l=10875
+ ad=-1.10758e+09 pd=316100 as=0 ps=0 
M1788 S00584 Vdd Vdd GND efet w=10875 l=14500
+ ad=-1.16224e+09 pd=307400 as=0 ps=0 
M1789 S00585 Vdd Vdd GND efet w=10150 l=11600
+ ad=-1.19168e+09 pd=295800 as=0 ps=0 
M1790 Vdd Vdd N0571 GND efet w=5800 l=68875
+ ad=0 pd=0 as=-1.69862e+08 ps=817800 
M1791 Vdd Vdd N0574 GND efet w=6525 l=65975
+ ad=0 pd=0 as=2.0205e+09 ps=429200 
M1792 Vdd Vdd N0573 GND efet w=5800 l=66700
+ ad=0 pd=0 as=0 ps=0 
M1793 Vdd Vdd N0600 GND efet w=5800 l=63800
+ ad=0 pd=0 as=-1.173e+08 ps=797500 
M1794 N0582 SC_A22 REG_RFSH_0 GND efet w=8700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1795 Vdd Vdd REG_RFSH_0 GND efet w=5800 l=33350
+ ad=0 pd=0 as=0 ps=0 
M1796 Vdd Vdd N0610 GND efet w=5800 l=72500
+ ad=0 pd=0 as=1.94481e+09 ps=435000 
M1797 Vdd Vdd N0609 GND efet w=5800 l=63800
+ ad=0 pd=0 as=0 ps=0 
M1798 Vdd Vdd REG_RFSH_1 GND efet w=6525 l=41325
+ ad=0 pd=0 as=0 ps=0 
M1799 N0617 SC_A22 REG_RFSH_1 GND efet w=10875 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1800 N0440 S00601 Vdd GND efet w=7250 l=53650
+ ad=0 pd=0 as=0 ps=0 
M1801 N0409 X12 ADDR_RFSH_1 GND efet w=8700 l=11600
+ ad=-9.89837e+08 pd=664100 as=0 ps=0 
M1802 ADDR_PTR_1 X32 N0409 GND efet w=8700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1803 N0420 X12 ADDR_RFSH_0 GND efet w=8700 l=11600
+ ad=-6.74462e+08 pd=765600 as=0 ps=0 
M1804 ADDR_PTR_0 X32 N0420 GND efet w=7975 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1805 N0449 S00613 N0449 GND efet w=73950 l=29000
+ ad=1.77241e+09 pd=350900 as=0 ps=0 
M1806 Vdd Vdd N0450 GND efet w=7250 l=59450
+ ad=0 pd=0 as=8.87255e+08 ps=179800 
M1807 S00598 Vdd Vdd GND efet w=10150 l=11600
+ ad=-1.1307e+09 pd=290000 as=0 ps=0 
M1808 S00599 Vdd Vdd GND efet w=11600 l=10150
+ ad=-1.23793e+09 pd=298700 as=0 ps=0 
M1809 S00600 Vdd Vdd GND efet w=10875 l=10150
+ ad=-1.28629e+09 pd=301600 as=0 ps=0 
M1810 S00601 Vdd Vdd GND efet w=11600 l=11600
+ ad=-1.26526e+09 pd=304500 as=0 ps=0 
M1811 __POC_CLK2_X12_X32__INH N0449 Vdd GND efet w=41325 l=21025
+ ad=0 pd=0 as=0 ps=0 
M1812 Vdd Vdd S00613 GND efet w=7975 l=12325
+ ad=0 pd=0 as=-1.76776e+09 ps=350900 
M1813 GND JUN_JMS N0309 GND efet w=34075 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1814 Vdd S00613 N0449 GND efet w=5800 l=43500
+ ad=0 pd=0 as=0 ps=0 
M1815 GND N0450 __POC_CLK2_X12_X32__INH GND efet w=29725 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1816 Vdd Vdd N0318 GND efet w=6525 l=68875
+ ad=0 pd=0 as=1.70136e+09 ps=1.189e+06 
M1817 N0308 X22 N0304 GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1818 N0309 N0310 N0308 GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1819 N0323 M12 GND GND efet w=32625 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1820 N0304 A32 GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1821 N0323 JUN_JMS N0324 GND efet w=36975 l=20300
+ ad=0 pd=0 as=0 ps=0 
M1822 N0320 SC GND GND efet w=30450 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1823 N0319 JIN_FIN N0320 GND efet w=29000 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1824 N0318 X22 N0319 GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1825 N0324 N0310 N0318 GND efet w=29000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1826 N0321 JCN_ISZ N0323 GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1827 N0318 N0322 N0321 GND efet w=31175 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1828 N0450 N0449 GND GND efet w=13050 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1829 Vdd Vdd N0437 GND efet w=8700 l=51475
+ ad=0 pd=0 as=4.5414e+08 ps=110200 
M1830 GND N0437 ___SC__JIN_FIN__CLK1_M11_X21_INH_ GND efet w=20300 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1831 Vdd S00612 N0436 GND efet w=7250 l=40600
+ ad=0 pd=0 as=-2.10837e+09 ps=449500 
M1832 Vdd Vdd S00612 GND efet w=5800 l=10150
+ ad=0 pd=0 as=-2.0495e+09 ps=249400 
M1833 S00628 Vdd Vdd GND efet w=5800 l=11600
+ ad=2.01209e+09 pd=310300 as=0 ps=0 
M1834 Vdd S00628 __INH__X11_X31_CLK1 GND efet w=7975 l=18125
+ ad=0 pd=0 as=1.83358e+08 ps=954100 
M1835 N0436 S00612 N0436 GND efet w=48575 l=23200
+ ad=0 pd=0 as=0 ps=0 
M1836 Vdd N0436 ___SC__JIN_FIN__CLK1_M11_X21_INH_ GND efet w=21025 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1837 GND N0436 N0437 GND efet w=13775 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1838 __INH__X11_X31_CLK1 S00628 __INH__X11_X31_CLK1 GND efet w=81925 l=22475
+ ad=0 pd=0 as=0 ps=0 
M1839 __INH__X11_X31_CLK1 N0517 GND GND efet w=35525 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1840 GND INH __INH__X11_X31_CLK1 GND efet w=36250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1841 GND N0522 __INH__X11_X31_CLK1 GND efet w=34800 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1842 Vdd Vdd N0451 GND efet w=5800 l=50750
+ ad=0 pd=0 as=4.91985e+08 ps=110200 
M1843 N0449 INH GND GND efet w=13775 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1844 N0436 N0443 GND GND efet w=13775 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1845 N0436 N0435 N0441 GND efet w=29725 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1846 N0449 POC GND GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1847 GND N0447 N0449 GND efet w=14500 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1848 N0449 N0451 GND GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1849 N0441 JIN_FIN GND GND efet w=29725 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1850 GND N0438 N0436 GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1851 GND A22 N0318 GND efet w=18125 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1852 N0451 clk2 GND GND efet w=14500 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1853 GND _CN N0322 GND efet w=34075 l=13775
+ ad=0 pd=0 as=-1.03189e+09 ps=669900 
M1854 N0322 SC GND GND efet w=26825 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1855 N0333 SC N0326 GND efet w=32625 l=10150
+ ad=0 pd=0 as=8.2418e+08 ps=171100 
M1856 N0326 A12 GND GND efet w=12325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1857 N0334 JIN_FIN N0333 GND efet w=31900 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1858 GND X32 N0334 GND efet w=30450 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1859 Vdd Vdd N0326 GND efet w=7975 l=64525
+ ad=0 pd=0 as=0 ps=0 
M1860 N0341 N0310 N0339 GND efet w=36250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1861 N0326 JUN_JMS N0341 GND efet w=38425 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1862 N0338 JCN_ISZ N0326 GND efet w=33350 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1863 N0339 N0322 N0338 GND efet w=33350 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1864 GND M22 N0339 GND efet w=34800 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1865 GND SC N0310 GND efet w=27550 l=10875
+ ad=0 pd=0 as=-1.13095e+08 ps=878700 
M1866 N0310 Vdd Vdd GND efet w=5800 l=27550
+ ad=0 pd=0 as=0 ps=0 
M1867 N0322 Vdd Vdd GND efet w=6525 l=28275
+ ad=0 pd=0 as=0 ps=0 
M1868 N0344 S00654 Vdd GND efet w=6525 l=28275
+ ad=7.94745e+08 pd=182700 as=0 ps=0 
M1869 Vdd N0344 SC GND efet w=37700 l=11600
+ ad=0 pd=0 as=-1.23509e+08 ps=4.8256e+06 
M1870 Vdd Vdd S00654 GND efet w=6525 l=13050
+ ad=0 pd=0 as=2.06886e+09 ps=284200 
M1871 GND X12 N0447 GND efet w=15225 l=12325
+ ad=0 pd=0 as=5.95007e+08 ps=133400 
M1872 GND X32 N0447 GND efet w=12325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1873 Vdd Vdd N0443 GND efet w=6525 l=51475
+ ad=0 pd=0 as=9.86073e+08 ps=217500 
M1874 N0447 Vdd Vdd GND efet w=5800 l=66700
+ ad=0 pd=0 as=0 ps=0 
M1875 N0443 clk1 GND GND efet w=14500 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1876 Vdd Vdd _INH GND efet w=5800 l=27550
+ ad=0 pd=0 as=-1.0403e+09 ps=655400 
M1877 Vdd Vdd INH GND efet w=5800 l=29000
+ ad=0 pd=0 as=-2.68923e+07 ps=913500 
M1878 N0511 Vdd Vdd GND efet w=7975 l=54375
+ ad=0 pd=0 as=0 ps=0 
M1879 N0517 clk2 N0511 GND efet w=9425 l=15225
+ ad=1.27201e+09 pd=272600 as=0 ps=0 
M1880 N0466 Vdd Vdd GND efet w=6525 l=73225
+ ad=-1.92965e+09 pd=452400 as=0 ps=0 
M1881 GND N0459 N0466 GND efet w=11600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1882 GND N0459 ADDR_PTR_0 GND efet w=18850 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1883 ADDR_PTR_0 Vdd Vdd GND efet w=7975 l=68875
+ ad=0 pd=0 as=0 ps=0 
M1884 N0459 N0466 GND GND efet w=13050 l=11600
+ ad=-2.83397e+08 pd=829400 as=0 ps=0 
M1885 Vdd Vdd N0459 GND efet w=6525 l=65250
+ ad=0 pd=0 as=0 ps=0 
M1886 N0505 N0466 GND GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1887 Vdd Vdd N0505 GND efet w=9425 l=76125
+ ad=0 pd=0 as=0 ps=0 
M1888 N0521 clk1 ADDR_PTR_0 GND efet w=8700 l=10875
+ ad=7.37977e+08 pd=153700 as=0 ps=0 
M1889 N0505 clk1 N0506 GND efet w=7250 l=10150
+ ad=0 pd=0 as=9.1669e+08 ps=194300 
M1890 REG_RFSH_0 clk1 N0566 GND efet w=7975 l=15225
+ ad=0 pd=0 as=1.08069e+09 ps=214600 
M1891 N0571 SC_A12_CLK2 N0572 GND efet w=24650 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1892 N0572 N0566 GND GND efet w=34075 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1893 GND N0574 REG_RFSH_0 GND efet w=21750 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1894 GND N0574 N0571 GND efet w=12325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1895 N0586 clk1 N0573 GND efet w=7975 l=13775
+ ad=1.1816e+09 pd=243600 as=0 ps=0 
M1896 N0573 N0571 GND GND efet w=12325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1897 N0574 N0571 GND GND efet w=12325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1898 REG_RFSH_1 N0571 N0593 GND efet w=10150 l=12325
+ ad=0 pd=0 as=1.13114e+09 ps=220400 
M1899 GND N0521 N0520 GND efet w=39150 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1900 Vdd Vdd N0494 GND efet w=7250 l=65250
+ ad=0 pd=0 as=1.22155e+09 ps=266800 
M1901 __INH__X32_CLK2 Vdd Vdd GND efet w=6525 l=28275
+ ad=1.55585e+09 pd=307400 as=0 ps=0 
M1902 N0520 CLK2_JMS_DC_M22_BBL_M22_X12_X22__ N0466 GND efet w=19575 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1903 N0509 N0506 GND GND efet w=39150 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1904 N0459 CLK2_JMS_DC_M22_BBL_M22_X12_X22__ N0509 GND efet w=20300 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1905 GND N0592 RRAB1 GND efet w=40600 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1906 GND N0494 __INH__X32_CLK2 GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1907 Vdd Vdd N0522 GND efet w=5800 l=36250
+ ad=0 pd=0 as=1.45493e+09 ps=313200 
M1908 CLK2_JMS_DC_M22_BBL_M22_X12_X22__ N0467 GND GND efet w=26825 l=13050
+ ad=1.03233e+09 pd=232000 as=0 ps=0 
M1909 GND DC RRAB1 GND efet w=31175 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1910 N0574 SC_A12_CLK2 N0585 GND efet w=21025 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1911 N0625 N0571 N0609 GND efet w=8700 l=13050
+ ad=1.24678e+09 pd=255200 as=0 ps=0 
M1912 GND N0600 N0609 GND efet w=13050 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1913 N0600 N0574 N0601 GND efet w=21750 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1914 GND N0610 REG_RFSH_1 GND efet w=21750 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1915 N0600 N0610 GND GND efet w=11600 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1916 N0585 N0586 GND GND efet w=35525 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1917 N0601 N0593 GND GND efet w=33350 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1918 RRAB1 clk2 GND GND efet w=29000 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1919 Vdd Vdd CLK2_JMS_DC_M22_BBL_M22_X12_X22__ GND efet w=9425 l=30450
+ ad=0 pd=0 as=0 ps=0 
M1920 GND clk2 N0496 GND efet w=29725 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1921 N0496 X32 N0495 GND efet w=31175 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1922 GND INH _INH GND efet w=26100 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1923 GND N0524 INH GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1924 GND M22 N0511 GND efet w=18850 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1925 N0522 clk1 GND GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1926 N0495 _INH N0494 GND efet w=29000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1927 N0429 X12 GND GND efet w=21750 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1928 N0438 clk2 N0428 GND efet w=7975 l=12325
+ ad=1.38555e+09 pd=298700 as=0 ps=0 
M1929 N0428 _INH N0429 GND efet w=21750 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1930 N0435 SC GND GND efet w=14500 l=10875
+ ad=-1.93596e+09 pd=478500 as=0 ps=0 
M1931 Vdd Vdd N0528 GND efet w=5800 l=52200
+ ad=0 pd=0 as=1.0912e+09 ps=229100 
M1932 N0428 Vdd Vdd GND efet w=5800 l=65250
+ ad=0 pd=0 as=0 ps=0 
M1933 N0428 A32 GND GND efet w=14500 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1934 N0435 Vdd Vdd GND efet w=7250 l=47850
+ ad=0 pd=0 as=0 ps=0 
M1935 GND X22 N0511 GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1936 GND DC N0526 GND efet w=29725 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1937 GND _CN N0528 GND efet w=16675 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1938 GND SC N0525 GND efet w=21750 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1939 N0525 JIN_FIN N0524 GND efet w=25375 l=10875
+ ad=0 pd=0 as=-1.2989e+09 ps=585800 
M1940 N0526 N0528 N0527 GND efet w=29725 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1941 Vdd Vdd N0467 GND efet w=5800 l=63800
+ ad=0 pd=0 as=1.39606e+09 ps=301600 
M1942 N0485 JMS GND GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1943 N0484 M22 N0485 GND efet w=31900 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1944 N0467 DC N0484 GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1945 Vdd Vdd N0460 GND efet w=5800 l=33350
+ ad=0 pd=0 as=7.84233e+08 ps=171100 
M1946 Vdd Vdd N0588 GND efet w=5800 l=70325
+ ad=0 pd=0 as=0 ps=0 
M1947 N0592 clk2 N0588 GND efet w=13050 l=13050
+ ad=1.89856e+09 pd=391500 as=0 ps=0 
M1948 GND clk2 N0460 GND efet w=21750 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1949 N0610 N0600 GND GND efet w=12325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1950 N0610 N0574 N0624 GND efet w=21750 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1951 N0624 N0625 GND GND efet w=36250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1952 D3 SC_M22_CLK2 N0646 GND efet w=10150 l=13050
+ ad=0 pd=0 as=9.4192e+08 ps=194300 
M1953 Vdd Vdd N0637 GND efet w=5800 l=65250
+ ad=0 pd=0 as=1.33298e+09 ps=278400 
M1954 Vdd Vdd N0642 GND efet w=6525 l=67425
+ ad=0 pd=0 as=8.22078e+08 ps=174000 
M1955 Vdd Vdd N0641 GND efet w=7250 l=69600
+ ad=0 pd=0 as=0 ps=0 
M1956 N0646 SC_A22 REG_RFSH_2 GND efet w=7250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1957 Vdd Vdd REG_RFSH_2 GND efet w=5075 l=34075
+ ad=0 pd=0 as=0 ps=0 
M1958 REG_RFSH_2 N0600 N0633 GND efet w=7975 l=12325
+ ad=0 pd=0 as=1.06807e+09 ps=229100 
M1959 N0637 N0610 N0638 GND efet w=21025 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1960 GND N0642 REG_RFSH_2 GND efet w=21750 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1961 N0637 N0642 GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1962 N0638 N0633 GND GND efet w=36250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1963 N0653 N0600 N0641 GND efet w=10875 l=15225
+ ad=1.25729e+09 pd=240700 as=0 ps=0 
M1964 N0641 N0637 GND GND efet w=11600 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1965 N0642 N0637 GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1966 Vdd Vdd __FIN_X12_ GND efet w=5800 l=51475
+ ad=0 pd=0 as=1.80394e+09 ps=365400 
M1967 GND N0578 WRAB1 GND efet w=24650 l=11600
+ ad=0 pd=0 as=9.5918e+08 ps=997600 
M1968 GND N0649 SC_A12_CLK2 GND efet w=21025 l=12325
+ ad=0 pd=0 as=1.53482e+09 ps=333500 
M1969 SC_A22_M22_CLK2 S00624 SC_A22_M22_CLK2 GND efet w=55825 l=27550
+ ad=-8.78405e+08 pd=698900 as=0 ps=0 
M1970 RRAB0 DC GND GND efet w=39150 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1971 Vdd Vdd N0608 GND efet w=5800 l=71050
+ ad=0 pd=0 as=0 ps=0 
M1972 GND N0615 RRAB0 GND efet w=36975 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1973 GND N0460 CLK2_JMS_DC_M22_BBL_M22_X12_X22__ GND efet w=29725 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1974 N0608 clk2 N0615 GND efet w=16675 l=10875
+ ad=0 pd=0 as=1.66518e+09 ps=330600 
M1975 N0589 X22 GND GND efet w=22475 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1976 N0594 N0580 N0588 GND efet w=32625 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1977 N0588 FIN_FIM_SRC_JIN N0589 GND efet w=21750 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1978 N0595 X12 N0594 GND efet w=29725 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1979 N0468 BBL GND GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1980 N0527 JCN_ISZ N0524 GND efet w=29000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1981 N0524 JUN_JMS N0526 GND efet w=21750 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1982 N0468 M22 N0467 GND efet w=25375 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1983 N0467 X22 N0468 GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1984 N0467 X12 N0468 GND efet w=21750 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1985 GND INC_ISZ_ADD_SUB_XCH_LD N0595 GND efet w=30450 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1986 GND clk2 RRAB0 GND efet w=34800 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1987 N0608 X12 N0602 GND efet w=31175 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1988 __FIN_X12_ X12 N0639 GND efet w=42775 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1989 Vdd Vdd DC GND efet w=8700 l=24650
+ ad=0 pd=0 as=-1.58607e+09 ps=2.1344e+06 
M1990 WRAB1 Vdd Vdd GND efet w=5800 l=33350
+ ad=0 pd=0 as=0 ps=0 
M1991 N0547 Vdd Vdd GND efet w=5800 l=69600
+ ad=-1.93596e+09 pd=432100 as=0 ps=0 
M1992 Vdd Vdd WRAB0 GND efet w=7250 l=29000
+ ad=0 pd=0 as=2.7797e+08 ps=817800 
M1993 SC_A12_CLK2 Vdd Vdd GND efet w=5800 l=36250
+ ad=0 pd=0 as=0 ps=0 
M1994 SC_A22_M22_CLK2 S00624 Vdd GND efet w=10150 l=27550
+ ad=0 pd=0 as=0 ps=0 
M1995 SC_A22_M22_CLK2 N0655 GND GND efet w=37700 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1996 N0642 N0610 N0652 GND efet w=24650 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1997 N0652 N0653 GND GND efet w=33350 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1998 GND N0622 N0621 GND efet w=12325 l=12325
+ ad=0 pd=0 as=5.25625e+08 ps=118900 
M1999 N0621 S00620 N0621 GND efet w=52925 l=29000
+ ad=0 pd=0 as=0 ps=0 
M2000 Vdd S00620 N0621 GND efet w=6525 l=54375
+ ad=0 pd=0 as=0 ps=0 
M2001 GND N0622 CLK2_SC_A12_M12_ GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2002 GND N0626 N0627 GND efet w=11600 l=11600
+ ad=0 pd=0 as=5.27727e+08 ps=133400 
M2003 N0626 S00627 N0626 GND efet w=52925 l=18125
+ ad=-1.97801e+09 pd=490100 as=0 ps=0 
M2004 CLK2_SC_A12_M12_ N0621 Vdd GND efet w=18850 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2005 __POC__CLK2_SC_A32_X12_ N0627 GND GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2006 S00624 Vdd Vdd GND efet w=6525 l=10875
+ ad=-1.71099e+09 pd=287100 as=0 ps=0 
M2007 WRAB0 N0547 GND GND efet w=33350 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2008 N0602 _OPA_0 N0614 GND efet w=52925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2009 N0640 _OPA_0 N0639 GND efet w=80475 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2010 GND N0636 N0640 GND efet w=42775 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2011 GND INC_ISZ_ADD_SUB_XCH_LD N0614 GND efet w=29725 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2012 GND SC N0612 GND efet w=29725 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2013 DC SC GND GND efet w=60175 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2014 GND FIN_FIM_SRC_JIN N0602 GND efet w=21750 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2015 N0580 _OPA_0 GND GND efet w=55100 l=11600
+ ad=-8.80507e+08 pd=672800 as=0 ps=0 
M2016 GND DC N0597 GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2017 N0597 FIN_FIM_SRC_JIN N0596 GND efet w=31175 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2018 N0649 Vdd Vdd GND efet w=5800 l=71050
+ ad=-2.0516e+09 pd=432100 as=0 ps=0 
M2019 Vdd Vdd N0655 GND efet w=5800 l=71050
+ ad=0 pd=0 as=8.13668e+08 ps=153700 
M2020 S00620 Vdd Vdd GND efet w=7250 l=11600
+ ad=-1.57643e+09 pd=348000 as=0 ps=0 
M2021 N0655 clk2 N0656 GND efet w=30450 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2022 N0649 clk2 N0650 GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2023 N0626 S00627 Vdd GND efet w=5800 l=52200
+ ad=0 pd=0 as=0 ps=0 
M2024 N0612 X32 N0611 GND efet w=36975 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2025 N0564 N0590 GND GND efet w=29725 l=14500
+ ad=1.87122e+09 pd=365400 as=0 ps=0 
M2026 N0524 Vdd Vdd GND efet w=5800 l=60900
+ ad=0 pd=0 as=0 ps=0 
M2027 GND _OPR_3 IO GND efet w=31900 l=12325
+ ad=0 pd=0 as=9.54535e+08 ps=214600 
M2028 OPE _OPR_3 GND GND efet w=32625 l=10875
+ ad=1.08279e+09 pd=220400 as=0 ps=0 
M2029 GND DC INC_ISZ GND efet w=24650 l=11600
+ ad=0 pd=0 as=3.3684e+08 ps=910600 
M2030 N0580 Vdd Vdd GND efet w=5800 l=27550
+ ad=0 pd=0 as=0 ps=0 
M2031 GND N0603 N0568 GND efet w=28275 l=14500
+ ad=0 pd=0 as=1.57898e+09 ps=281300 
M2032 N0596 _OPA_0 N0590 GND efet w=54375 l=12325
+ ad=0 pd=0 as=7.25362e+08 ps=145000 
M2033 N0568 Vdd Vdd GND efet w=5800 l=27550
+ ad=0 pd=0 as=0 ps=0 
M2034 N0563 N0564 N0562 GND efet w=34075 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2035 GND M12 N0563 GND efet w=34075 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2036 N0576 M22 GND GND efet w=31175 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2037 N0575 N0564 N0576 GND efet w=30450 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2038 N0562 clk2 N0547 GND efet w=34075 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2039 N0567 _OPA_0 N0562 GND efet w=53650 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2040 N0603 INC_ISZ_XCH N0611 GND efet w=31175 l=12325
+ ad=7.84233e+08 pd=174000 as=0 ps=0 
M2041 Vdd Vdd N0603 GND efet w=6525 l=64525
+ ad=0 pd=0 as=0 ps=0 
M2042 N0564 Vdd Vdd GND efet w=5800 l=27550
+ ad=0 pd=0 as=0 ps=0 
M2043 N0579 N0568 GND GND efet w=31175 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2044 GND N0568 N0567 GND efet w=30450 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2045 N0575 N0580 N0579 GND efet w=30450 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2046 N0654 SC N0656 GND efet w=32625 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2047 N0651 A12 N0650 GND efet w=32625 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2048 GND SC N0651 GND efet w=30450 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2049 GND M22 N0654 GND efet w=31175 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2050 Vdd Vdd N0622 GND efet w=7250 l=68150
+ ad=0 pd=0 as=9.60842e+08 ps=185600 
M2051 S00627 Vdd Vdd GND efet w=6525 l=10875
+ ad=-1.51756e+09 pd=330600 as=0 ps=0 
M2052 Vdd Vdd N0627 GND efet w=5800 l=52200
+ ad=0 pd=0 as=0 ps=0 
M2053 N0622 clk2 N0623 GND efet w=36975 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2054 GND M12 N0618 GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2055 N0682 X12 N0683 GND efet w=84825 l=16675
+ ad=0 pd=0 as=0 ps=0 
M2056 N0618 A12 GND GND efet w=36250 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2057 GND A22 N0654 GND efet w=29725 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2058 N0578 clk2 N0575 GND efet w=31900 l=13050
+ ad=-2.41347e+08 pd=754000 as=0 ps=0 
M2059 Vdd Vdd N0578 GND efet w=7975 l=67425
+ ad=0 pd=0 as=0 ps=0 
M2060 N0590 Vdd Vdd GND efet w=5800 l=65250
+ ad=0 pd=0 as=0 ps=0 
M2061 N0618 SC N0623 GND efet w=34075 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2062 GND POC N0683 GND efet w=86275 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2063 Vdd Vdd SC_A22 GND efet w=5800 l=34800
+ ad=0 pd=0 as=1.73666e+09 ps=371200 
M2064 __POC__CLK2_SC_A32_X12_ N0626 Vdd GND efet w=21750 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2065 Vdd Vdd N0679 GND efet w=9425 l=65975
+ ad=0 pd=0 as=9.14588e+08 ps=179800 
M2066 Vdd Vdd SC_M22_CLK2 GND efet w=7975 l=25375
+ ad=0 pd=0 as=1.62822e+09 ps=1.7603e+06 
M2067 SC_M22_CLK2 N0679 GND GND efet w=37700 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2068 N0626 N0630 GND GND efet w=13775 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2069 GND POC N0626 GND efet w=16675 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2070 N0679 M22 N0680 GND efet w=32625 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2071 GND N0643 SC_A22 GND efet w=25375 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2072 N0703 clk2 N0682 GND efet w=14500 l=13050
+ ad=-1.85186e+09 pd=443700 as=0 ps=0 
M2073 N0681 clk2 N0680 GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2074 N0681 SC GND GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2075 N0629 X12 GND GND efet w=31175 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2076 XCH _OPR_3 GND GND efet w=30450 l=15225
+ ad=-1.08655e+09 pd=643800 as=0 ps=0 
M2077 GND _OPR_3 BBL GND efet w=30450 l=13050
+ ad=0 pd=0 as=2.07306e+09 ps=423400 
M2078 N0628 _OPR_3 GND GND efet w=53650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2079 INC_ISZ_XCH _OPR_3 N0587 GND efet w=47850 l=11600
+ ad=7.4849e+08 pd=156600 as=0 ps=0 
M2080 LD _OPR_3 GND GND efet w=31175 l=11600
+ ad=5.17215e+08 pd=124700 as=0 ps=0 
M2081 SUB _OPR_3 GND GND efet w=30450 l=10875
+ ad=1.94481e+09 pd=374100 as=0 ps=0 
M2082 ADD _OPR_3 GND GND efet w=31175 l=13050
+ ad=1.3456e+09 pd=272600 as=0 ps=0 
M2083 JCN_ISZ OPR_3 GND GND efet w=50025 l=11600
+ ad=1.29138e+09 pd=1.1339e+06 as=0 ps=0 
M2084 GND OPR_3 JCN GND efet w=25375 l=13050
+ ad=0 pd=0 as=1.1774e+09 ps=249400 
M2085 FIN_FIM OPR_3 GND GND efet w=23925 l=13775
+ ad=1.80815e+09 pd=368300 as=0 ps=0 
M2086 N0361 Vdd Vdd GND efet w=6525 l=35525
+ ad=0 pd=0 as=0 ps=0 
M2087 N0344 S00654 N0344 GND efet w=69600 l=5075
+ ad=0 pd=0 as=0 ps=0 
M2088 GND N0343 SC GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2089 N0344 N0343 GND GND efet w=29000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2090 GND OPR_3 ISZ GND efet w=24650 l=11600
+ ad=0 pd=0 as=1.64416e+09 ps=336400 
M2091 GND OPR_3 FIM_SRC GND efet w=23925 l=12325
+ ad=0 pd=0 as=1.90697e+09 ps=388600 
M2092 GND OPR_3 JIN_FIN GND efet w=44950 l=11600
+ ad=0 pd=0 as=-1.9986e+09 ps=1.3079e+06 
M2093 JUN_JMS OPR_3 GND GND efet w=44225 l=11600
+ ad=1.73711e+09 pd=1.2441e+06 as=0 ps=0 
M2094 GND OPR_3 INC_ISZ GND efet w=23200 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2095 ISZ _OPR_2 GND GND efet w=31175 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2096 IO _OPR_2 GND GND efet w=29725 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2097 OPE _OPR_2 GND GND efet w=31175 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2098 JUN_JMS _OPR_2 GND GND efet w=55825 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2099 GND OPR_3 JMS GND efet w=24650 l=11600
+ ad=0 pd=0 as=-1.22321e+09 ps=635100 
M2100 GND OPR_3 N0636 GND efet w=23200 l=11600
+ ad=0 pd=0 as=-1.0889e+08 ps=835200 
M2101 LDM_BBL _OPR_3 GND GND efet w=31900 l=13050
+ ad=-9.18352e+08 pd=603200 as=0 ps=0 
M2102 GND A32 N0629 GND efet w=29725 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2103 N0629 SC N0631 GND efet w=34075 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2104 GND IOR N0683 GND efet w=81925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2105 GND A32 N0682 GND efet w=51475 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2106 N0682 M12 GND GND efet w=36975 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2107 GND N0703 L GND efet w=52925 l=13775
+ ad=0 pd=0 as=-7.01795e+08 ps=710500 
M2108 L N0703 GND GND efet w=60900 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2109 N0631 clk2 N0630 GND efet w=30450 l=8700
+ ad=0 pd=0 as=8.17873e+08 ps=185600 
M2110 GND M12 N0662 GND efet w=29725 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2111 N0662 SC N0661 GND efet w=29725 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2112 N0644 A22 N0643 GND efet w=23925 l=9425
+ ad=0 pd=0 as=1.42129e+09 ps=290000 
M2113 GND SC N0644 GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2114 N0661 clk2 N0660 GND efet w=30450 l=10150
+ ad=0 pd=0 as=8.36795e+08 ps=188500 
M2115 N0682 Vdd Vdd GND efet w=9425 l=35525
+ ad=0 pd=0 as=0 ps=0 
M2116 Vdd Vdd N0630 GND efet w=6525 l=64525
+ ad=0 pd=0 as=0 ps=0 
M2117 INC_ISZ_ADD_SUB_XCH_LD OPR_3 N0628 GND efet w=47850 l=13050
+ ad=-1.02137e+09 pd=652500 as=0 ps=0 
M2118 N0587 OPR_3 GND GND efet w=39875 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2119 GND _OPR_2 N0523 GND efet w=92075 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2120 INC_ISZ _OPR_2 GND GND efet w=30450 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2121 BBL _OPR_2 GND GND efet w=30450 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2122 N0373 JCN_ISZ N0372 GND efet w=36250 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2123 N0372 FIN_FIM N0373 GND efet w=33350 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2124 JMS _OPR_2 GND GND efet w=31900 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2125 GND OPR_3 FIN_FIM_SRC_JIN GND efet w=24650 l=11600
+ ad=0 pd=0 as=1.62401e+09 ps=1.972e+06 
M2126 GND OPR_3 JUN2_JMS2 GND efet w=24650 l=11600
+ ad=0 pd=0 as=-1.64582e+09 ps=469800 
M2127 N0628 _OPR_2 INC_ISZ_ADD_SUB_XCH_LD GND efet w=56550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2128 N0587 _OPR_2 GND GND efet w=46400 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2129 LDM_BBL _OPR_2 GND GND efet w=32625 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2130 N0523 OPR_2 JCN_ISZ GND efet w=98600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2131 GND OPR_2 FIN_FIM GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2132 GND OPR_2 JCN GND efet w=23925 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2133 FIM_SRC OPR_2 GND GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2134 JUN2_JMS2 _OPR_2 GND GND efet w=32625 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2135 GND OPR_2 JIN_FIN GND efet w=44950 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2136 FIN_FIM _OPR_1 GND GND efet w=31175 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2137 ISZ _OPR_1 GND GND efet w=31900 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2138 GND OPR_2 XCH GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2139 GND OPR_2 N0636 GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2140 N0628 OPR_2 GND GND efet w=46400 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2141 OPR_2 N0995 Vdd GND efet w=47850 l=20300
+ ad=1.01683e+09 pd=2.5404e+06 as=0 ps=0 
M2142 Vdd N0994 _OPR_2 GND efet w=33350 l=15950
+ ad=0 pd=0 as=1.43943e+09 ps=2.8014e+06 
M2143 N0587 OPR_2 INC_ISZ_XCH GND efet w=40600 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2144 GND OPR_2 FIN_FIM_SRC_JIN GND efet w=25375 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2145 FIM_SRC _OPR_1 GND GND efet w=29725 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2146 IO _OPR_1 GND GND efet w=29725 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2147 OPE _OPR_1 GND GND efet w=30450 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2148 JIN_FIN _OPR_1 GND GND efet w=53650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2149 INC_ISZ _OPR_1 GND GND efet w=29725 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2150 N0523 _OPR_1 GND GND efet w=89175 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2151 XCH _OPR_1 GND GND efet w=30450 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2152 GND OPR_2 LD GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2153 GND OPR_2 SUB GND efet w=23200 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2154 GND OPR_2 ADD GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2155 N0628 _OPR_1 INC_ISZ_ADD_SUB_XCH_LD GND efet w=57275 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2156 GND _OPR_1 N0587 GND efet w=45675 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2157 N0361 clk1 N0343 GND efet w=14500 l=13050
+ ad=0 pd=0 as=-2.12729e+09 ps=437900 
M2158 N0372 X32 GND GND efet w=37700 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2159 N0352 Vdd Vdd GND efet w=7975 l=64525
+ ad=1.20894e+09 pd=266800 as=0 ps=0 
M2160 GND N0362 N0361 GND efet w=22475 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2161 N0373 JUN_JMS N0372 GND efet w=31900 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2162 N0368 SC N0373 GND efet w=34800 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2163 GND OPR_1 JCN GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2164 GND OPR_1 JUN_JMS GND efet w=46400 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2165 N0636 _OPR_1 GND GND efet w=23200 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2166 N0523 OPR_1 JCN_ISZ GND efet w=96425 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2167 GND OPR_1 BBL GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2168 GND OPR_1 JMS GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2169 INC_ISZ_XCH _OPR_1 N0587 GND efet w=46400 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2170 FIN_FIM_SRC_JIN _OPR_1 GND GND efet w=30450 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2171 LD _OPR_1 GND GND efet w=31900 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2172 GND N0995 _OPR_2 GND efet w=32625 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2173 OPR_2 N0994 GND GND efet w=29725 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2174 L Vdd Vdd GND efet w=10150 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2175 OPR_3 N0993 Vdd GND efet w=39150 l=14500
+ ad=1.31118e+09 pd=2.5404e+06 as=0 ps=0 
M2176 Vdd N0992 _OPR_3 GND efet w=20300 l=14500
+ ad=0 pd=0 as=3.70631e+07 ps=2.5636e+06 
M2177 Vdd Vdd N0643 GND efet w=7250 l=60900
+ ad=0 pd=0 as=0 ps=0 
M2178 N0660 Vdd Vdd GND efet w=6525 l=63075
+ ad=0 pd=0 as=0 ps=0 
M2179 GND N0660 SC_M12_CLK2 GND efet w=36975 l=9425
+ ad=0 pd=0 as=-2.11047e+09 ps=423400 
M2180 SC_M12_CLK2 Vdd Vdd GND efet w=6525 l=26100
+ ad=0 pd=0 as=0 ps=0 
M2181 D0 SC_M12_CLK2 N1011 GND efet w=11600 l=12325
+ ad=0 pd=0 as=-3.23345e+08 ps=870000 
M2182 D2 SC_M12_CLK2 N1009 GND efet w=10875 l=11600
+ ad=0 pd=0 as=-8.95225e+08 ps=701800 
M2183 OPR_3 N0992 GND GND efet w=29725 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2184 GND N0993 _OPR_3 GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2185 N0998 Vdd Vdd GND efet w=8700 l=30450
+ ad=-8.3215e+08 pd=701800 as=0 ps=0 
M2186 N0994 Vdd Vdd GND efet w=10150 l=32625
+ ad=-1.95488e+09 pd=458200 as=0 ps=0 
M2187 GND N1011 N0998 GND efet w=58725 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2188 GND N1008 N0992 GND efet w=62350 l=11600
+ ad=0 pd=0 as=2.13824e+09 ps=429200 
M2189 D1 SC_M12_CLK2 N1010 GND efet w=10875 l=12325
+ ad=0 pd=0 as=-1.72781e+09 ps=524900 
M2190 N0996 Vdd Vdd GND efet w=12325 l=29000
+ ad=8.56158e+08 pd=1.0643e+06 as=0 ps=0 
M2191 GND N1009 N0994 GND efet w=61625 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2192 N0992 Vdd Vdd GND efet w=8700 l=33350
+ ad=0 pd=0 as=0 ps=0 
M2193 GND OPR_1 SUB GND efet w=23925 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2194 GND OPR_1 ADD GND efet w=23925 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2195 LDM_BBL OPR_1 GND GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2196 ISZ _OPR_0 GND GND efet w=31900 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2197 JCN _OPR_0 GND GND efet w=31175 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2198 OPE _OPR_0 GND GND efet w=30450 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2199 JIN_FIN _OPR_0 GND GND efet w=52200 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2200 GND X32 N0352 GND efet w=12325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2201 N0367 N0352 GND GND efet w=21750 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2202 N0368 N0343 N0367 GND efet w=21750 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2203 N0362 clk2 N0368 GND efet w=8700 l=11600
+ ad=5.3824e+08 pd=121800 as=0 ps=0 
M2204 Vdd Vdd N0368 GND efet w=6525 l=67425
+ ad=0 pd=0 as=0 ps=0 
M2205 XCH _OPR_0 GND GND efet w=29725 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2206 GND _OPR_0 JCN_ISZ GND efet w=53650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2207 JMS _OPR_0 GND GND efet w=31175 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2208 GND OPR_1 JUN2_JMS2 GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2209 INC_ISZ_XCH _OPR_0 N0587 GND efet w=52200 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2210 N0636 _OPR_0 GND GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2211 SUB _OPR_0 GND GND efet w=31175 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2212 Vdd N0998 _OPR_0 GND efet w=39875 l=21750
+ ad=0 pd=0 as=4.51256e+08 ps=2.7289e+06 
M2213 GND OPA_0 FIN_FIM GND efet w=21750 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2214 GND OPR_0 FIM_SRC GND efet w=25375 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2215 GND OPR_0 IO GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2216 Vdd Vdd N0769 GND efet w=6525 l=39875
+ ad=0 pd=0 as=6.16033e+08 ps=145000 
M2217 POC Vdd Vdd GND efet w=7975 l=22475
+ ad=-9.88858e+08 pd=6.3336e+06 as=0 ps=0 
M2218 _CN Vdd Vdd GND efet w=10150 l=28275
+ ad=-4.66315e+08 pd=626400 as=0 ps=0 
M2219 N0769 A12 GND GND efet w=18125 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2220 FIN_FIM Vdd Vdd GND efet w=5800 l=59450
+ ad=0 pd=0 as=0 ps=0 
M2221 GND OPR_0 BBL GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2222 OPR_0 N0999 Vdd GND efet w=20300 l=17400
+ ad=-8.96447e+08 pd=2.3171e+06 as=0 ps=0 
M2223 GND OPR_0 LD GND efet w=24650 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2224 GND OPR_0 ADD GND efet w=23200 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2225 ISZ Vdd Vdd GND efet w=7250 l=63800
+ ad=0 pd=0 as=0 ps=0 
M2226 JCN Vdd Vdd GND efet w=5800 l=62350
+ ad=0 pd=0 as=0 ps=0 
M2227 FIM_SRC Vdd Vdd GND efet w=5800 l=63075
+ ad=0 pd=0 as=0 ps=0 
M2228 IO Vdd Vdd GND efet w=9425 l=73225
+ ad=0 pd=0 as=0 ps=0 
M2229 N0493 Vdd Vdd GND efet w=7250 l=72500
+ ad=5.6347e+08 pd=121800 as=0 ps=0 
M2230 Vdd Vdd OPE GND efet w=7250 l=56550
+ ad=0 pd=0 as=0 ps=0 
M2231 JIN_FIN Vdd Vdd GND efet w=7250 l=36975
+ ad=0 pd=0 as=0 ps=0 
M2232 Vdd Vdd N0510 GND efet w=7250 l=50750
+ ad=0 pd=0 as=8.53615e+08 ps=182700 
M2233 JUN_JMS Vdd Vdd GND efet w=8700 l=39150
+ ad=0 pd=0 as=0 ps=0 
M2234 JCN_ISZ Vdd Vdd GND efet w=8700 l=34800
+ ad=0 pd=0 as=0 ps=0 
M2235 INC_ISZ Vdd Vdd GND efet w=7250 l=55100
+ ad=0 pd=0 as=0 ps=0 
M2236 Vdd Vdd DCL GND efet w=5800 l=63800
+ ad=0 pd=0 as=7.0644e+08 ps=153700 
M2237 GND OPA_0 N0516 GND efet w=38425 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2238 N0516 FIM_SRC _SRC GND efet w=23200 l=13050
+ ad=0 pd=0 as=1.46754e+09 ps=298700 
M2239 GND SC N0417 GND efet w=33350 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2240 GND reset N0327 GND efet w=35525 l=12325
+ ad=0 pd=0 as=1.55165e+09 ps=313200 
M2241 GND N0397 _CN GND efet w=57275 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2242 GND N0327 N0769 GND efet w=19575 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2243 POC N0327 GND GND efet w=55825 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2244 N0412 N0397 GND GND efet w=21750 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2245 N0399 X32 GND GND efet w=13775 l=12325
+ ad=5.02498e+08 pd=127600 as=0 ps=0 
M2246 N0417 X32 N0418 GND efet w=34075 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2247 GND IO N0493 GND efet w=13775 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2248 N0510 OPE GND GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2249 Vdd N0510 _OPE GND efet w=29000 l=11600
+ ad=0 pd=0 as=1.77004e+07 ps=1.6646e+06 
M2250 GND IO _I_O GND efet w=34800 l=11600
+ ad=0 pd=0 as=1.38477e+09 ps=2.9058e+06 
M2251 _I_O N0493 Vdd GND efet w=13775 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2252 GND ISZ N0456 GND efet w=13050 l=11600
+ ad=0 pd=0 as=8.53615e+08 ps=171100 
M2253 GND JCN N0476 GND efet w=13775 l=12325
+ ad=0 pd=0 as=5.65572e+08 ps=124700 
M2254 _OPE OPE GND GND efet w=29725 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2255 Vdd Vdd O_IB GND efet w=7250 l=53650
+ ad=0 pd=0 as=-1.76776e+09 ps=481400 
M2256 Vdd Vdd KBP GND efet w=5800 l=65975
+ ad=0 pd=0 as=2.11301e+09 ps=475600 
M2257 Vdd Vdd TCS GND efet w=8700 l=43500
+ ad=0 pd=0 as=-4.15415e+08 ps=1.5341e+06 
M2258 Vdd Vdd DAA GND efet w=8700 l=43500
+ ad=0 pd=0 as=-8.74246e+07 ps=1.5863e+06 
M2259 XCH Vdd Vdd GND efet w=5800 l=57275
+ ad=0 pd=0 as=0 ps=0 
M2260 BBL Vdd Vdd GND efet w=6525 l=57275
+ ad=0 pd=0 as=0 ps=0 
M2261 JMS Vdd Vdd GND efet w=7250 l=55100
+ ad=0 pd=0 as=0 ps=0 
M2262 N0636 Vdd Vdd GND efet w=6525 l=60900
+ ad=0 pd=0 as=0 ps=0 
M2263 INC_ISZ_ADD_SUB_XCH_LD Vdd Vdd GND efet w=10150 l=65250
+ ad=0 pd=0 as=0 ps=0 
M2264 Vdd Vdd IOW GND efet w=5800 l=56550
+ ad=0 pd=0 as=-1.14542e+09 ps=617700 
M2265 Vdd Vdd RAR GND efet w=7250 l=55100
+ ad=0 pd=0 as=-1.54279e+09 ps=519100 
M2266 RAL Vdd Vdd GND efet w=6525 l=55100
+ ad=-1.09917e+09 pd=580000 as=0 ps=0 
M2267 CMA Vdd Vdd GND efet w=6525 l=55825
+ ad=-1.25685e+09 pd=591600 as=0 ps=0 
M2268 Vdd Vdd TCC GND efet w=7250 l=56550
+ ad=0 pd=0 as=1.34981e+09 ps=269700 
M2269 STC Vdd Vdd GND efet w=5800 l=61625
+ ad=1.53062e+09 pd=298700 as=0 ps=0 
M2270 INC_ISZ_XCH Vdd Vdd GND efet w=5800 l=65250
+ ad=0 pd=0 as=0 ps=0 
M2271 LD Vdd Vdd GND efet w=6525 l=67425
+ ad=0 pd=0 as=0 ps=0 
M2272 FIN_FIM_SRC_JIN Vdd Vdd GND efet w=7250 l=50750
+ ad=0 pd=0 as=0 ps=0 
M2273 IOW _I_O GND GND efet w=38425 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2274 Vdd Vdd CMC GND efet w=7250 l=53650
+ ad=0 pd=0 as=-2.10626e+09 ps=423400 
M2275 Vdd Vdd DAC GND efet w=6525 l=52925
+ ad=0 pd=0 as=8.7464e+08 ps=203000 
M2276 Vdd Vdd IAC GND efet w=5800 l=56550
+ ad=0 pd=0 as=1.54954e+09 ps=304500 
M2277 Vdd Vdd CLC GND efet w=7250 l=63075
+ ad=0 pd=0 as=7.94745e+08 ps=165300 
M2278 SUB Vdd Vdd GND efet w=7250 l=60900
+ ad=0 pd=0 as=0 ps=0 
M2279 ADD Vdd Vdd GND efet w=7250 l=59450
+ ad=0 pd=0 as=0 ps=0 
M2280 LDM_BBL Vdd Vdd GND efet w=7975 l=58725
+ ad=0 pd=0 as=0 ps=0 
M2281 JUN2_JMS2 Vdd Vdd GND efet w=7250 l=63800
+ ad=0 pd=0 as=0 ps=0 
M2282 Vdd Vdd CLB GND efet w=7975 l=65250
+ ad=0 pd=0 as=8.95665e+08 ps=197200 
M2283 Vdd Vdd SBM GND efet w=7250 l=56550
+ ad=0 pd=0 as=1.67149e+09 ps=350900 
M2284 ADM Vdd Vdd GND efet w=5800 l=56550
+ ad=1.36663e+09 pd=269700 as=0 ps=0 
M2285 OPR_0 N0998 GND GND efet w=21025 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2286 GND N0999 _OPR_0 GND efet w=29725 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2287 _OPR_1 N0996 Vdd GND efet w=38425 l=15950
+ ad=1.61394e+09 pd=2.8768e+06 as=0 ps=0 
M2288 Vdd N0997 OPR_1 GND efet w=24650 l=13050
+ ad=0 pd=0 as=-2.82517e+08 ps=2.4244e+06 
M2289 N0999 N0998 GND GND efet w=27550 l=11600
+ ad=-1.39308e+09 pd=1.4239e+06 as=0 ps=0 
M2290 GND N1010 N0996 GND efet w=58000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2291 N0995 N0994 GND GND efet w=29000 l=11600
+ ad=1.26825e+09 pd=1.0324e+06 as=0 ps=0 
M2292 N0997 N0996 GND GND efet w=29000 l=10150
+ ad=-2.01375e+09 pd=466900 as=0 ps=0 
M2293 D3 SC_M12_CLK2 N1008 GND efet w=10150 l=12325
+ ad=0 pd=0 as=1.31196e+09 ps=263900 
M2294 N0993 N0992 GND GND efet w=26825 l=10875
+ ad=-9.73017e+08 pd=600300 as=0 ps=0 
M2295 N0999 Vdd Vdd GND efet w=13050 l=42050
+ ad=0 pd=0 as=0 ps=0 
M2296 _OPR_1 N0997 GND GND efet w=34075 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2297 GND N0996 OPR_1 GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2298 N0995 Vdd Vdd GND efet w=14500 l=43500
+ ad=0 pd=0 as=0 ps=0 
M2299 N0997 Vdd Vdd GND efet w=9425 l=36975
+ ad=0 pd=0 as=0 ps=0 
M2300 N0993 Vdd Vdd GND efet w=15950 l=38425
+ ad=0 pd=0 as=0 ps=0 
M2301 D3 OPA_IB OPA_3 GND efet w=58725 l=13775
+ ad=0 pd=0 as=2.44481e+07 ps=2.2939e+06 
M2302 Vdd Vdd IOR GND efet w=10875 l=41325
+ ad=0 pd=0 as=1.44065e+09 ps=1.0962e+06 
M2303 SBM _I_O GND GND efet w=31900 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2304 ADM _I_O GND GND efet w=31900 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2305 Vdd Vdd N0477 GND efet w=5800 l=49300
+ ad=0 pd=0 as=1.95743e+09 ps=359600 
M2306 GND __X31__CLK2_ N0480 GND efet w=13775 l=12325
+ ad=0 pd=0 as=5.92905e+08 ps=139200 
M2307 N0480 Vdd Vdd GND efet w=7250 l=67425
+ ad=0 pd=0 as=0 ps=0 
M2308 N0482 N0480 N0477 GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2309 N0479 Vdd Vdd GND efet w=7250 l=77575
+ ad=6.09725e+08 pd=136300 as=0 ps=0 
M2310 N0482 N0479 GND GND efet w=26825 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2311 N0479 IOR GND GND efet w=12325 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2312 N0412 N0399 N0413 GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2313 N0418 N0419 N0413 GND efet w=30450 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2314 GND N0769 N0327 GND efet w=33350 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2315 N0297 clk2 GND GND efet w=26100 l=11600
+ ad=6.60185e+08 pd=145000 as=0 ps=0 
M2316 N0297 S00678 N0297 GND efet w=74675 l=5075
+ ad=0 pd=0 as=0 ps=0 
M2317 X22 clk2 N0280 GND efet w=13775 l=12325
+ ad=-1.35269e+09 pd=2.2359e+06 as=1.18791e+09 ps=237800 
M2318 Vdd S00678 N0297 GND efet w=7975 l=32625
+ ad=0 pd=0 as=0 ps=0 
M2319 Vdd Vdd S00678 GND efet w=5800 l=13050
+ ad=0 pd=0 as=2.11722e+09 ps=298700 
M2320 N0295 N0297 N0296 GND efet w=27550 l=11600
+ ad=2.02681e+09 pd=388600 as=0 ps=0 
M2321 N0296 N0280 GND GND efet w=62350 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2322 Vdd Vdd N0296 GND efet w=7975 l=21025
+ ad=0 pd=0 as=0 ps=0 
M2323 N0739 clk1 N0296 GND efet w=11600 l=11600
+ ad=1.97215e+09 pd=408900 as=0 ps=0 
M2324 N0404 clk1 N0397 GND efet w=14500 l=11600
+ ad=0 pd=0 as=1.50329e+09 ps=295800 
M2325 GND N0405 N0404 GND efet w=26825 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2326 N0413 clk2 N0405 GND efet w=8700 l=11600
+ ad=0 pd=0 as=6.37057e+08 ps=139200 
M2327 Vdd Vdd N0399 GND efet w=7250 l=84100
+ ad=0 pd=0 as=0 ps=0 
M2328 GND test N0432 GND efet w=36250 l=10150
+ ad=0 pd=0 as=-1.81612e+09 ps=519100 
M2329 Vdd Vdd N0432 GND efet w=7250 l=55100
+ ad=0 pd=0 as=0 ps=0 
M2330 N0327 Vdd Vdd GND efet w=5800 l=26100
+ ad=0 pd=0 as=0 ps=0 
M2331 Vdd Vdd N0404 GND efet w=7250 l=36250
+ ad=0 pd=0 as=0 ps=0 
M2332 Vdd Vdd N0784 GND efet w=5800 l=50750
+ ad=0 pd=0 as=5.15113e+08 ps=113100 
M2333 N0741 N0739 GND GND efet w=31900 l=10875
+ ad=1.30565e+09 pd=261000 as=0 ps=0 
M2334 Vdd Vdd N0329 GND efet w=8700 l=20300
+ ad=0 pd=0 as=-1.79299e+09 ps=545200 
M2335 N0413 Vdd Vdd GND efet w=6525 l=63075
+ ad=0 pd=0 as=0 ps=0 
M2336 N0456 Vdd Vdd GND efet w=10875 l=65975
+ ad=0 pd=0 as=0 ps=0 
M2337 GND N0476 N0478 GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2338 GND _OPE DCL GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2339 O_IB _OPE GND GND efet w=23200 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2340 GND _OPE KBP GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2341 GND _OPE TCS GND efet w=38425 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2342 DAA _OPE GND GND efet w=34075 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2343 RAR _OPE GND GND efet w=23925 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2344 GND _OPE RAL GND efet w=23925 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2345 GND _OPE CMA GND efet w=25375 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2346 N0478 N0487 N0481 GND efet w=44225 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2347 N0478 _OPA_3 N0481 GND efet w=63800 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2348 N0478 N0456 N0419 GND efet w=41325 l=13775
+ ad=0 pd=0 as=6.68595e+08 ps=150800 
M2349 GND _I_O N0329 GND efet w=59450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2350 N0476 Vdd Vdd GND efet w=5800 l=58000
+ ad=0 pd=0 as=0 ps=0 
M2351 N0478 ADD_0 N0419 GND efet w=47125 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2352 N0419 Vdd Vdd GND efet w=5800 l=50025
+ ad=0 pd=0 as=0 ps=0 
M2353 Vdd Vdd _SRC GND efet w=5800 l=68875
+ ad=0 pd=0 as=0 ps=0 
M2354 DCL _OPA_3 GND GND efet w=30450 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2355 KBP _OPA_3 GND GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2356 TCS _OPA_3 GND GND efet w=40600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2357 DAA _OPA_3 GND GND efet w=40600 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2358 GND N0486 N0481 GND efet w=50750 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2359 GND OPA_3 N0481 GND efet w=75400 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2360 GND _OPE TCC GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2361 STC _OPE GND GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2362 GND _OPE CMC GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2363 GND _OPE DAC GND efet w=23200 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2364 GND _OPE IAC GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2365 GND _I_O IOR GND efet w=39875 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2366 N0477 A12 N0483 GND efet w=31900 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2367 D2 OPA_IB OPA_2 GND efet w=61625 l=16675
+ ad=0 pd=0 as=3.28581e+07 ps=2.2707e+06 
M2368 GND IOR N0483 GND efet w=31175 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2369 GND _OPE CLC GND efet w=23200 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2370 CLB _OPE GND GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2371 STC _OPA_3 GND GND efet w=31175 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2372 DAC _OPA_3 GND GND efet w=30450 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2373 SBM _OPA_3 GND GND efet w=32625 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2374 ADM _OPA_3 GND GND efet w=30450 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2375 IOR _OPA_3 GND GND efet w=44950 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2376 GND N1001 _OPA_3 GND efet w=29725 l=11600
+ ad=0 pd=0 as=8.50731e+08 ps=2.5868e+06 
M2377 OPA_3 N1000 GND GND efet w=57275 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2378 GND OPA_3 O_IB GND efet w=23200 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2379 GND OPA_3 IOW GND efet w=31900 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2380 GND OPA_3 RAR GND efet w=24650 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2381 GND OPA_3 RAL GND efet w=23925 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2382 GND OPA_3 CMA GND efet w=23200 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2383 GND OPA_3 TCC GND efet w=23200 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2384 GND OPA_3 CMC GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2385 GND OPA_3 IAC GND efet w=23925 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2386 GND N0486 N0487 GND efet w=13050 l=11600
+ ad=0 pd=0 as=1.59369e+09 ps=330600 
M2387 DCL _OPA_2 GND GND efet w=30450 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2388 GND OPA_2 N0501 GND efet w=44950 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2389 N0501 ACC_0 N0486 GND efet w=29000 l=10875
+ ad=0 pd=0 as=1.19422e+09 ps=261000 
M2390 N0487 Vdd Vdd GND efet w=5800 l=50750
+ ad=0 pd=0 as=0 ps=0 
M2391 Vdd Vdd N0398 GND efet w=6525 l=26100
+ ad=0 pd=0 as=7.6531e+08 ps=171100 
M2392 KBP _OPA_2 GND GND efet w=30450 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2393 RAR _OPA_2 GND GND efet w=31900 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2394 RAL _OPA_2 GND GND efet w=31175 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2395 GND OPA_3 CLC GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2396 GND OPA_3 CLB GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2397 CMA _OPA_2 GND GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2398 TCC _OPA_2 GND GND efet w=31175 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2399 N0486 Vdd Vdd GND efet w=5800 l=47850
+ ad=0 pd=0 as=0 ps=0 
M2400 GND OPA_2 TCS GND efet w=34075 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2401 GND OPA_2 DAA GND efet w=34800 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2402 GND N1003 _OPA_2 GND efet w=36975 l=15225
+ ad=0 pd=0 as=-2.32057e+08 ps=2.3635e+06 
M2403 OPA_2 N1002 GND GND efet w=54375 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2404 Vdd N1000 _OPA_3 GND efet w=22475 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2405 OPA_3 N1001 Vdd GND efet w=25375 l=9425
+ ad=0 pd=0 as=0 ps=0 
M2406 GND OPA_2 STC GND efet w=23200 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2407 GND OPA_2 CMC GND efet w=24650 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2408 GND OPA_2 DAC GND efet w=23925 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2409 GND OPA_2 IAC GND efet w=27550 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2410 GND OPA_2 CLC GND efet w=27550 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2411 CLB OPA_2 GND GND efet w=23200 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2412 DAA _OPA_1 GND GND efet w=43500 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2413 GND clk2 N0398 GND efet w=47850 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2414 Vdd Vdd N0799 GND efet w=6525 l=67425
+ ad=0 pd=0 as=6.09725e+08 ps=133400 
M2415 N0741 S00690 N0741 GND efet w=72500 l=5800
+ ad=0 pd=0 as=0 ps=0 
M2416 Vdd S00690 N0741 GND efet w=6525 l=26825
+ ad=0 pd=0 as=0 ps=0 
M2417 Vdd Vdd S00690 GND efet w=5800 l=13050
+ ad=0 pd=0 as=-2.08524e+09 ps=263900 
M2418 X32 N0739 GND GND efet w=31900 l=11600
+ ad=1.50339e+09 pd=4.5907e+06 as=0 ps=0 
M2419 GND N0782 N0784 GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2420 Vdd N0741 X32 GND efet w=36250 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2421 N0414 clk2 A22 GND efet w=8700 l=11600
+ ad=5.2983e+08 pd=118900 as=-2.22471e+07 ps=1.7168e+06 
M2422 N0799 _SRC GND GND efet w=13050 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2423 N0407 N0414 GND GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2424 N0407 N0398 N0408 GND efet w=8700 l=13050
+ ad=0 pd=0 as=4.66755e+08 ps=127600 
M2425 Vdd Vdd S00685 GND efet w=6525 l=11600
+ ad=0 pd=0 as=-1.90863e+09 ps=287100 
M2426 Vdd S00685 N0415 GND efet w=5800 l=16675
+ ad=0 pd=0 as=-1.23749e+09 ps=1.3804e+06 
M2427 N0415 S00685 N0415 GND efet w=69600 l=26825
+ ad=0 pd=0 as=0 ps=0 
M2428 N0507 CY_1 N0486 GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2429 RAR _OPA_1 GND GND efet w=31175 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2430 TCC _OPA_1 GND GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2431 GND OPA_1 N0507 GND efet w=45675 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2432 STC _OPA_1 GND GND efet w=31900 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2433 CMC _OPA_1 GND GND efet w=31175 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2434 IAC _OPA_1 GND GND efet w=31900 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2435 GND OPA_2 SBM GND efet w=28275 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2436 GND OPA_2 ADM GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2437 ADM _OPA_1 GND GND efet w=29725 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2438 _COM N0782 Vdd GND efet w=20300 l=11600
+ ad=-1.58817e+09 pd=2.2823e+06 as=0 ps=0 
M2439 GND N0784 _COM GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2440 N0800 N0801 N0782 GND efet w=30450 l=10150
+ ad=0 pd=0 as=1.48437e+09 ps=330600 
M2441 GND N0329 N0800 GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2442 N0798 N0805 GND GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2443 N0782 N0799 N0798 GND efet w=29725 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2444 GND N0797 N0782 GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2445 GND clk2 N0375 GND efet w=16675 l=12325
+ ad=0 pd=0 as=1.19422e+09 ps=246500 
M2446 N0797 N0408 GND GND efet w=20300 l=12325
+ ad=5.90802e+08 pd=130500 as=0 ps=0 
M2447 Vdd Vdd N0797 GND efet w=7975 l=55100
+ ad=0 pd=0 as=0 ps=0 
M2448 Vdd N0742 X22 GND efet w=39150 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2449 X22 N0719 GND GND efet w=36975 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2450 GND X22 N0288 GND efet w=25375 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2451 N0742 N0719 GND GND efet w=30450 l=11600
+ ad=1.38344e+09 pd=272600 as=0 ps=0 
M2452 N0742 S00710 N0742 GND efet w=70325 l=5800
+ ad=0 pd=0 as=0 ps=0 
M2453 Vdd Vdd S00710 GND efet w=6525 l=13775
+ ad=0 pd=0 as=2.14245e+09 ps=263900 
M2454 Vdd S00710 N0742 GND efet w=7250 l=27550
+ ad=0 pd=0 as=0 ps=0 
M2455 N0718 N0281 GND GND efet w=26825 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2456 N0281 clk2 X12 GND efet w=13050 l=13775
+ ad=5.69777e+08 pd=127600 as=2.34698e+08 ps=2.6187e+06 
M2457 N0719 clk1 N0718 GND efet w=14500 l=11600
+ ad=1.89015e+09 pd=429200 as=0 ps=0 
M2458 Vdd Vdd N0718 GND efet w=8700 l=37700
+ ad=0 pd=0 as=0 ps=0 
M2459 N0383 X22 GND GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2460 N0782 S00699 N0782 GND efet w=15950 l=58000
+ ad=0 pd=0 as=0 ps=0 
M2461 N0288 X12 GND GND efet w=21750 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2462 Vdd N0743 X12 GND efet w=35525 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2463 X12 N0721 GND GND efet w=36975 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2464 N0743 S00725 N0743 GND efet w=75400 l=5800
+ ad=1.79974e+09 pd=353800 as=0 ps=0 
M2465 N0743 N0721 GND GND efet w=26100 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2466 Vdd Vdd S00725 GND efet w=5800 l=11600
+ ad=0 pd=0 as=-2.10416e+09 ps=263900 
M2467 Vdd S00725 N0743 GND efet w=7975 l=26825
+ ad=0 pd=0 as=0 ps=0 
M2468 Vdd S00699 N0782 GND efet w=5800 l=39875
+ ad=0 pd=0 as=0 ps=0 
M2469 N0380 clk2 N0383 GND efet w=8700 l=11600
+ ad=7.50593e+08 pd=171100 as=0 ps=0 
M2470 Vdd Vdd N0407 GND efet w=5800 l=49300
+ ad=0 pd=0 as=0 ps=0 
M2471 GND OPA_1 DCL GND efet w=24650 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2472 GND OPA_1 KBP GND efet w=29000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2473 GND OPA_1 TCS GND efet w=33350 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2474 GND OPA_1 RAL GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2475 GND OPA_1 CMA GND efet w=24650 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2476 GND OPA_1 DAC GND efet w=23200 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2477 GND OPA_1 CLC GND efet w=23200 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2478 GND OPA_1 CLB GND efet w=24650 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2479 GND OPA_1 SBM GND efet w=23925 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2480 N0512 N0432 N0486 GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2481 GND OPA_0 N0512 GND efet w=49300 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2482 DCL _OPA_0 GND GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2483 TCS _OPA_0 GND GND efet w=42050 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2484 DAA _OPA_0 GND GND efet w=41325 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2485 RAL _OPA_0 GND GND efet w=31175 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2486 TCC _OPA_0 GND GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2487 CMC _OPA_0 GND GND efet w=31900 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2488 CLC _OPA_0 GND GND efet w=31175 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2489 ADM _OPA_0 GND GND efet w=29725 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2490 GND OPA_0 KBP GND efet w=24650 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2491 GND OPA_0 RAR GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2492 GND OPA_0 DAC GND efet w=26100 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2493 Vdd N1002 _OPA_2 GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2494 OPA_1 N1004 GND GND efet w=68875 l=12325
+ ad=2.13673e+08 pd=2.2475e+06 as=0 ps=0 
M2495 GND OPA_0 CMA GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2496 GND OPA_0 STC GND efet w=23200 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2497 GND OPA_0 IAC GND efet w=23200 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2498 GND OPA_0 CLB GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2499 GND OPA_0 SBM GND efet w=24650 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2500 GND _OPE N0415 GND efet w=44225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2501 GND N0353 N0351 GND efet w=22475 l=10875
+ ad=0 pd=0 as=1.04749e+09 ps=1.1078e+06 
M2502 N0351 __X21__CLK2_ GND GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2503 GND DCL N0353 GND efet w=14500 l=10150
+ ad=0 pd=0 as=4.83575e+08 ps=118900 
M2504 WRITE_ACC_1_ KBP GND GND efet w=14500 l=10150
+ ad=1.48857e+09 pd=310300 as=0 ps=0 
M2505 N0415 __X21__CLK2_ GND GND efet w=44225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2506 Vdd Vdd N0383 GND efet w=5800 l=47850
+ ad=0 pd=0 as=0 ps=0 
M2507 N0375 N0380 GND GND efet w=21750 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2508 Vdd Vdd __X31__CLK2_ GND efet w=5800 l=15950
+ ad=0 pd=0 as=-1.60753e+09 ps=1.4239e+06 
M2509 N0353 Vdd Vdd GND efet w=6525 l=64525
+ ad=0 pd=0 as=0 ps=0 
M2510 GND TCS WRITE_ACC_1_ GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2511 WRITE_ACC_1_ DAA GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2512 S00699 Vdd Vdd GND efet w=5800 l=11600
+ ad=-1.97381e+09 pd=310300 as=0 ps=0 
M2513 Vdd Vdd __X21__CLK2_ GND efet w=6525 l=18850
+ ad=0 pd=0 as=-1.71525e+08 ps=1.6182e+06 
M2514 __X31__CLK2_ N0375 GND GND efet w=65250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2515 N0375 Vdd Vdd GND efet w=5800 l=36250
+ ad=0 pd=0 as=0 ps=0 
M2516 N0369 Vdd Vdd GND efet w=5800 l=56550
+ ad=0 pd=0 as=0 ps=0 
M2517 N0337 Vdd Vdd GND efet w=5800 l=29000
+ ad=1.59369e+09 pd=330600 as=0 ps=0 
M2518 Vdd Vdd N0328 GND efet w=6525 l=64525
+ ad=0 pd=0 as=6.74903e+08 ps=142100 
M2519 N0720 N0282 GND GND efet w=26825 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2520 N0282 clk2 M22 GND efet w=15950 l=11600
+ ad=5.7188e+08 pd=127600 as=5.79508e+08 ps=2.6651e+06 
M2521 N0721 clk1 N0720 GND efet w=14500 l=11600
+ ad=1.95743e+09 pd=400200 as=0 ps=0 
M2522 Vdd Vdd N0720 GND efet w=7250 l=30450
+ ad=0 pd=0 as=0 ps=0 
M2523 N0337 N0360 GND GND efet w=34800 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2524 GND clk2 N0337 GND efet w=28275 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2525 __X21__CLK2_ N0337 GND GND efet w=53650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2526 GND N0329 N0328 GND efet w=13775 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2527 N0328 POC GND GND efet w=11600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2528 N0330 X22 N0331 GND efet w=29000 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2529 GND clk2 N0330 GND efet w=29725 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2530 N0369 X12 GND GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2531 N0360 clk2 N0369 GND efet w=9425 l=12325
+ ad=9.12485e+08 pd=208800 as=0 ps=0 
M2532 N0335 clk1 GND GND efet w=31175 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2533 N0336 N0337 N0335 GND efet w=31175 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2534 N0332 N0328 N0336 GND efet w=29725 l=12325
+ ad=1.08279e+09 pd=258100 as=0 ps=0 
M2535 N0331 N0329 N0332 GND efet w=30450 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2536 GND clk2 N0423 GND efet w=21750 l=13050
+ ad=0 pd=0 as=-1.83294e+09 ps=516200 
M2537 N0332 POC N0331 GND efet w=29000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2538 N0351 Vdd Vdd GND efet w=7250 l=43500
+ ad=0 pd=0 as=0 ps=0 
M2539 GND INC_ISZ N0442 GND efet w=15950 l=10150
+ ad=0 pd=0 as=-1.47762e+09 ps=559700 
M2540 N0442 Vdd Vdd GND efet w=6525 l=58725
+ ad=0 pd=0 as=0 ps=0 
M2541 GND TCS WRITE_CARRY_2_ GND efet w=11600 l=11600
+ ad=0 pd=0 as=-2.07707e+08 ps=826500 
M2542 GND TCS ADD_GROUP_4_ GND efet w=12325 l=12325
+ ad=0 pd=0 as=-1.76566e+09 ps=484300 
M2543 READ_ACC_3_ DAA GND GND efet w=13050 l=11600
+ ad=-9.09942e+08 pd=678600 as=0 ps=0 
M2544 GND N0446 N0448 GND efet w=76125 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2545 N0342 N0332 Vdd GND efet w=21025 l=11600
+ ad=-1.70845e+09 pd=1.4036e+06 as=0 ps=0 
M2546 Vdd Vdd N0423 GND efet w=6525 l=31175
+ ad=0 pd=0 as=0 ps=0 
M2547 GND M22 N0288 GND efet w=22475 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2548 Vdd N0744 M22 GND efet w=40600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2549 M22 N0723 GND GND efet w=34800 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2550 N0744 S00740 N0744 GND efet w=70325 l=5800
+ ad=1.29935e+09 pd=281300 as=0 ps=0 
M2551 N0744 N0723 GND GND efet w=27550 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2552 Vdd Vdd S00740 GND efet w=5800 l=11600
+ ad=0 pd=0 as=-2.11467e+09 ps=258100 
M2553 Vdd S00740 N0744 GND efet w=4350 l=31175
+ ad=0 pd=0 as=0 ps=0 
M2554 Vdd Vdd N0430 GND efet w=5800 l=49300
+ ad=0 pd=0 as=0 ps=0 
M2555 N0340 Vdd Vdd GND efet w=7250 l=72500
+ ad=6.49673e+08 pd=139200 as=0 ps=0 
M2556 N0430 N0423 N0431 GND efet w=10150 l=10875
+ ad=0 pd=0 as=1.41709e+09 ps=301600 
M2557 N0722 N0283 GND GND efet w=26825 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2558 N0283 clk2 M12 GND efet w=13775 l=15225
+ ad=5.44548e+08 pd=124700 as=6.40602e+06 ps=4.4138e+06 
M2559 N0723 clk1 N0722 GND efet w=14500 l=11600
+ ad=1.98686e+09 pd=394400 as=0 ps=0 
M2560 M12 clk2 N0433 GND efet w=8700 l=12325
+ ad=0 pd=0 as=7.37977e+08 ps=174000 
M2561 N0342 N0340 GND GND efet w=20300 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2562 GND N0332 N0340 GND efet w=11600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2563 Vdd S00731 N0332 GND efet w=6525 l=52925
+ ad=0 pd=0 as=0 ps=0 
M2564 S00731 Vdd Vdd GND efet w=6525 l=12325
+ ad=-1.20429e+09 pd=420500 as=0 ps=0 
M2565 N0332 S00731 N0332 GND efet w=70325 l=5075
+ ad=0 pd=0 as=0 ps=0 
M2566 Vdd Vdd N0805 GND efet w=11600 l=54375
+ ad=0 pd=0 as=1.08699e+09 ps=240700 
M2567 N0853 Vdd Vdd GND efet w=7975 l=67425
+ ad=1.14797e+09 pd=266800 as=0 ps=0 
M2568 X12 clk2 N0425 GND efet w=7975 l=13050
+ ad=0 pd=0 as=4.0368e+08 ps=104400 
M2569 N0421 Vdd Vdd GND efet w=5800 l=56550
+ ad=0 pd=0 as=0 ps=0 
M2570 N0421 N0423 N0422 GND efet w=10875 l=10875
+ ad=0 pd=0 as=5.3824e+08 ps=139200 
M2571 GND N0422 N0805 GND efet w=31175 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2572 N0853 X12 GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2573 GND N0433 N0430 GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2574 GND N0425 N0421 GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2575 N0801 Vdd Vdd GND efet w=6525 l=51475
+ ad=4.73503e+08 pd=948300 as=0 ps=0 
M2576 Vdd Vdd N0722 GND efet w=7975 l=38425
+ ad=0 pd=0 as=0 ps=0 
M2577 GND N0431 N0801 GND efet w=23925 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2578 N0288 M12 GND GND efet w=21750 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2579 Vdd N0745 M12 GND efet w=39150 l=21750
+ ad=0 pd=0 as=0 ps=0 
M2580 GND N0803 N0403 GND efet w=24650 l=10150
+ ad=0 pd=0 as=2.0228e+08 ps=843900 
M2581 M12 N0725 GND GND efet w=38425 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2582 N0717 S00757 N0717 GND efet w=65975 l=7250
+ ad=-1.65379e+09 pd=1.392e+06 as=0 ps=0 
M2583 GND POC N0717 GND efet w=70325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2584 N0717 S00757 Vdd GND efet w=10150 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2585 N0745 S00761 N0745 GND efet w=78300 l=8700
+ ad=1.90697e+09 pd=365400 as=0 ps=0 
M2586 N0403 N0802 GND GND efet w=21750 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2587 GND __X21__CLK2_ N0448 GND efet w=73950 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2588 GND XCH WRITE_ACC_1_ GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2589 WRITE_ACC_1_ POC GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2590 INC_GROUP_5_ INC_ISZ GND GND efet w=11600 l=12325
+ ad=-1.34516e+09 pd=539400 as=0 ps=0 
M2591 WRITE_CARRY_2_ POC GND GND efet w=15950 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2592 GND CMA WRITE_ACC_1_ GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2593 WRITE_ACC_1_ TCC GND GND efet w=13775 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2594 GND DAC WRITE_ACC_1_ GND efet w=11600 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2595 WRITE_ACC_1_ IAC GND GND efet w=11600 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2596 GND N1005 _OPA_1 GND efet w=34075 l=15225
+ ad=0 pd=0 as=-2.11379e+09 ps=1.972e+06 
M2597 WRITE_ACC_1_ CLB GND GND efet w=12325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2598 Vdd N1004 _OPA_1 GND efet w=30450 l=26100
+ ad=0 pd=0 as=0 ps=0 
M2599 OPA_1 N1005 Vdd GND efet w=26825 l=16675
+ ad=0 pd=0 as=0 ps=0 
M2600 GND LD WRITE_ACC_1_ GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2601 WRITE_ACC_1_ SUB GND GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2602 GND ADD WRITE_ACC_1_ GND efet w=13775 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2603 WRITE_ACC_1_ LDM_BBL GND GND efet w=13775 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2604 WRITE_CARRY_2_ SUB GND GND efet w=16675 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2605 WRITE_CARRY_2_ TCC GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2606 GND STC WRITE_CARRY_2_ GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2607 WRITE_CARRY_2_ CMC GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2608 GND DAC WRITE_CARRY_2_ GND efet w=13775 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2609 WRITE_CARRY_2_ IAC GND GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2610 GND CLC WRITE_CARRY_2_ GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2611 WRITE_CARRY_2_ CLB GND GND efet w=13775 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2612 GND SBM WRITE_CARRY_2_ GND efet w=13050 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2613 WRITE_CARRY_2_ ADM GND GND efet w=13775 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2614 GND RAR READ_ACC_3_ GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2615 READ_ACC_3_ RAL GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2616 N0448 N0445 ACB_IB GND efet w=74675 l=10875
+ ad=0 pd=0 as=1.52686e+09 ps=1.1397e+06 
M2617 ACB_IB __X31__CLK2_ N0448 GND efet w=76125 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2618 GND N0442 ADD_IB GND efet w=39150 l=12325
+ ad=0 pd=0 as=5.99653e+08 ps=965700 
M2619 GND XCH N0445 GND efet w=21750 l=11600
+ ad=0 pd=0 as=1.11853e+09 ps=237800 
M2620 GND N0446 CY_IB GND efet w=14500 l=11600
+ ad=0 pd=0 as=-8.59482e+08 ps=684400 
M2621 GND IOW N0446 GND efet w=21750 l=11600
+ ad=0 pd=0 as=-1.10968e+09 ps=638000 
M2622 ADD_GROUP_4_ TCC GND GND efet w=13050 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2623 READ_ACC_3_ IAC GND GND efet w=12325 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2624 GND DAC READ_ACC_3_ GND efet w=12325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2625 GND SBM READ_ACC_3_ GND efet w=11600 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2626 SUB_GROUP_6_ S00709 SUB_GROUP_6_ GND efet w=65250 l=14500
+ ad=6.12708e+08 pd=1.7893e+06 as=0 ps=0 
M2627 GND STC INC_GROUP_5_ GND efet w=11600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2628 N0502 RAL GND GND efet w=15225 l=10875
+ ad=4.43627e+08 pd=110200 as=0 ps=0 
M2629 CY_IB __X31__CLK2_ GND GND efet w=15950 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2630 SUB_GROUP_6_ CMC GND GND efet w=23925 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2631 SUB_GROUP_6_ S00709 Vdd GND efet w=5800 l=40600
+ ad=0 pd=0 as=0 ps=0 
M2632 INC_GROUP_5_ IAC GND GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2633 INC_GROUP_5_ Vdd Vdd GND efet w=7250 l=66700
+ ad=0 pd=0 as=0 ps=0 
M2634 READ_ACC_3_ Vdd Vdd GND efet w=7250 l=69600
+ ad=0 pd=0 as=0 ps=0 
M2635 GND RAR N0490 GND efet w=15225 l=15225
+ ad=0 pd=0 as=4.39422e+08 ps=104400 
M2636 GND __X31__CLK2_ ADSL GND efet w=17400 l=10875
+ ad=0 pd=0 as=1.54157e+09 ps=1.1774e+06 
M2637 GND __X31__CLK2_ ADD_IB GND efet w=38425 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2638 ADD_IB S00729 ADD_IB GND efet w=84100 l=28275
+ ad=0 pd=0 as=0 ps=0 
M2639 ADD_IB S00729 Vdd GND efet w=8700 l=24650
+ ad=0 pd=0 as=0 ps=0 
M2640 ACB_IB S00724 ACB_IB GND efet w=74675 l=50025
+ ad=0 pd=0 as=0 ps=0 
M2641 N0445 Vdd Vdd GND efet w=8700 l=41325
+ ad=0 pd=0 as=0 ps=0 
M2642 GND N0502 ADSL GND efet w=13050 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2643 CY_IB Vdd Vdd GND efet w=7975 l=70325
+ ad=0 pd=0 as=0 ps=0 
M2644 N0446 Vdd Vdd GND efet w=8700 l=43500
+ ad=0 pd=0 as=0 ps=0 
M2645 GND __X31__CLK2_ ADSR GND efet w=14500 l=11600
+ ad=0 pd=0 as=7.7416e+08 ps=1.0063e+06 
M2646 ADSR N0490 GND GND efet w=15950 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2647 GND CMA N0515 GND efet w=11600 l=11600
+ ad=0 pd=0 as=5.08805e+08 ps=116000 
M2648 Vdd Vdd S00709 GND efet w=6525 l=13775
+ ad=0 pd=0 as=-1.92335e+09 ps=263900 
M2649 ACB_IB S00724 Vdd GND efet w=10875 l=29725
+ ad=0 pd=0 as=0 ps=0 
M2650 Vdd Vdd ADSL GND efet w=8700 l=65250
+ ad=0 pd=0 as=0 ps=0 
M2651 N0502 Vdd Vdd GND efet w=5800 l=60900
+ ad=0 pd=0 as=0 ps=0 
M2652 Vdd Vdd N0490 GND efet w=7975 l=84825
+ ad=0 pd=0 as=0 ps=0 
M2653 ADSR Vdd Vdd GND efet w=7250 l=65250
+ ad=0 pd=0 as=0 ps=0 
M2654 ACC_ADAC N0515 GND GND efet w=13775 l=11600
+ ad=-1.23793e+09 pd=600300 as=0 ps=0 
M2655 GND N0342 ACC_ADAC GND efet w=13050 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2656 WRITE_CARRY_2_ Vdd Vdd GND efet w=6525 l=63800
+ ad=0 pd=0 as=0 ps=0 
M2657 N0515 Vdd Vdd GND efet w=7250 l=84100
+ ad=0 pd=0 as=0 ps=0 
M2658 GND N0853 N0854 GND efet w=19575 l=13775
+ ad=0 pd=0 as=-1.25055e+09 ps=591600 
M2659 READ_ACC_3_ ADM GND GND efet w=13050 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2660 ADD_GROUP_4_ ADM GND GND efet w=12325 l=16675
+ ad=0 pd=0 as=0 ps=0 
M2661 GND SBM SUB_GROUP_6_ GND efet w=21750 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2662 ADD_GROUP_4_ Vdd Vdd GND efet w=6525 l=60175
+ ad=0 pd=0 as=0 ps=0 
M2663 GND ADD WRITE_CARRY_2_ GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2664 READ_ACC_3_ SUB GND GND efet w=13050 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2665 GND IOR WRITE_ACC_1_ GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2666 GND ADD READ_ACC_3_ GND efet w=13775 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2667 GND ADD ADD_GROUP_4_ GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2668 SUB_GROUP_6_ SUB GND GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2669 Vdd Vdd N1001 GND efet w=13050 l=37700
+ ad=0 pd=0 as=8.51953e+08 ps=1.0034e+06 
M2670 OPA_2 N1003 Vdd GND efet w=32625 l=25375
+ ad=0 pd=0 as=0 ps=0 
M2671 N1001 N1000 GND GND efet w=27550 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2672 Vdd Vdd N1005 GND efet w=13050 l=33350
+ ad=0 pd=0 as=7.80468e+08 ps=922200 
M2673 D1 OPA_IB OPA_1 GND efet w=58725 l=18125
+ ad=0 pd=0 as=0 ps=0 
M2674 GND clk2 N0702 GND efet w=54375 l=12325
+ ad=0 pd=0 as=1.54157e+09 ps=1.1629e+06 
M2675 N0702 S00676 N0702 GND efet w=65250 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2676 S00676 Vdd Vdd GND efet w=8700 l=15950
+ ad=2.08358e+09 pd=249400 as=0 ps=0 
M2677 Vdd Vdd N0671 GND efet w=13050 l=33350
+ ad=0 pd=0 as=0 ps=0 
M2678 D0 OPA_IB OPA_0 GND efet w=65250 l=13050
+ ad=0 pd=0 as=1.64783e+07 ps=3.3031e+06 
M2679 GND N1007 _OPA_0 GND efet w=37700 l=14500
+ ad=0 pd=0 as=8.81046e+08 ps=4.2572e+06 
M2680 OPA_0 N1006 GND GND efet w=70325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2681 N0702 S00676 Vdd GND efet w=13050 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2682 N0671 N0702 N0688 GND efet w=27550 l=13775
+ ad=0 pd=0 as=3.1161e+08 ps=817800 
M2683 N0671 D3 GND GND efet w=53650 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2684 Vdd N1006 _OPA_0 GND efet w=52925 l=25375
+ ad=0 pd=0 as=0 ps=0 
M2685 OPA_0 N1007 Vdd GND efet w=29000 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2686 Vdd Vdd N1003 GND efet w=12325 l=35525
+ ad=0 pd=0 as=1.17994e+09 ps=962800 
M2687 N1005 N1004 GND GND efet w=26825 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2688 GND N1012 N1000 GND efet w=56550 l=13050
+ ad=0 pd=0 as=1.11873e+08 ps=838100 
M2689 GND N1014 N1004 GND efet w=55825 l=12325
+ ad=0 pd=0 as=-1.00245e+09 ps=585800 
M2690 GND JUN2_JMS2 N0658 GND efet w=15225 l=12325
+ ad=0 pd=0 as=1.25309e+09 ps=252300 
M2691 N1003 N1002 GND GND efet w=26100 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2692 Vdd Vdd N1007 GND efet w=9425 l=35525
+ ad=0 pd=0 as=-1.15197e+08 ps=791700 
M2693 N1007 N1006 GND GND efet w=34800 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2694 GND N1013 N1002 GND efet w=57275 l=12325
+ ad=0 pd=0 as=2.48535e+08 ps=823600 
M2695 GND N1015 N1006 GND efet w=64525 l=12325
+ ad=0 pd=0 as=-6.49232e+08 ps=667000 
M2696 Vdd Vdd S00689 GND efet w=8700 l=11600
+ ad=0 pd=0 as=-2.12098e+09 ps=252300 
M2697 S00687 Vdd Vdd GND efet w=8700 l=17400
+ ad=1.95953e+09 pd=246500 as=0 ps=0 
M2698 N0687 S00687 N0687 GND efet w=68875 l=7250
+ ad=7.38858e+08 pd=1.7458e+06 as=0 ps=0 
M2699 N0687 S00687 Vdd GND efet w=10150 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2700 Vdd S00689 N0689 GND efet w=10150 l=11600
+ ad=0 pd=0 as=2.49416e+08 ps=2.5404e+06 
M2701 N0689 S00689 N0689 GND efet w=55100 l=34075
+ ad=0 pd=0 as=0 ps=0 
M2702 Vdd N0659 D0 GND efet w=47125 l=18125
+ ad=0 pd=0 as=0 ps=0 
M2703 N0687 N0700 GND GND efet w=253750 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2704 GND N0700 N0689 GND efet w=228375 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2705 N0687 N0688 GND GND efet w=98600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2706 GND N0687 N0689 GND efet w=74675 l=5800
+ ad=0 pd=0 as=0 ps=0 
M2707 D0 SC_M22_CLK2 N1015 GND efet w=10150 l=13050
+ ad=0 pd=0 as=1.04074e+09 ps=197200 
M2708 Vdd N0659 D2 GND efet w=47125 l=16675
+ ad=0 pd=0 as=0 ps=0 
M2709 N1000 Vdd Vdd GND efet w=19575 l=42050
+ ad=0 pd=0 as=0 ps=0 
M2710 N0658 LDM_BBL GND GND efet w=14500 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2711 WRITE_ACC_1_ Vdd Vdd GND efet w=6525 l=71775
+ ad=0 pd=0 as=0 ps=0 
M2712 N1004 Vdd Vdd GND efet w=11600 l=30450
+ ad=0 pd=0 as=0 ps=0 
M2713 N1002 Vdd Vdd GND efet w=19575 l=42050
+ ad=0 pd=0 as=0 ps=0 
M2714 N1006 Vdd Vdd GND efet w=20300 l=40600
+ ad=0 pd=0 as=0 ps=0 
M2715 D2 SC_M22_CLK2 N1013 GND efet w=10875 l=13775
+ ad=0 pd=0 as=-1.28629e+09 ps=562600 
M2716 GND N0689 d3 GND efet w=1246275 l=6525
+ ad=0 pd=0 as=-1.95909e+09 ps=440800 
M2717 GND N0658 OPA_IB GND efet w=42050 l=15950
+ ad=0 pd=0 as=-3.12392e+08 ps=1.3137e+06 
M2718 Vdd Vdd N0658 GND efet w=7250 l=69600
+ ad=0 pd=0 as=0 ps=0 
M2719 OPA_IB __X21__CLK2_ GND GND efet w=41325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2720 D1 SC_M22_CLK2 N1014 GND efet w=10875 l=13775
+ ad=0 pd=0 as=-7.24922e+08 ps=690200 
M2721 d3 N0687 Vdd GND efet w=657575 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2722 OPA_IB S00716 OPA_IB GND efet w=37700 l=47850
+ ad=0 pd=0 as=0 ps=0 
M2723 D3 SC_M22_CLK2 N1012 GND efet w=10150 l=11600
+ ad=0 pd=0 as=2.77727e+07 ps=849700 
M2724 Vdd S00716 OPA_IB GND efet w=8700 l=20300
+ ad=0 pd=0 as=0 ps=0 
M2725 D1 N0659 Vdd GND efet w=46400 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2726 D3 N0659 Vdd GND efet w=39875 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2727 Vdd Vdd S00716 GND efet w=7250 l=11600
+ ad=0 pd=0 as=-1.8035e+09 ps=290000 
M2728 N0675 Vdd Vdd GND efet w=7975 l=36250
+ ad=8.95665e+08 pd=179800 as=0 ps=0 
M2729 N0659 Vdd Vdd GND efet w=11600 l=21025
+ ad=-9.85632e+08 pd=562600 as=0 ps=0 
M2730 N0659 N0675 GND GND efet w=53650 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2731 Vdd Vdd N0678 GND efet w=11600 l=37700
+ ad=0 pd=0 as=1.5979e+09 ps=304500 
M2732 GND INC_GROUP_5_ N0546 GND efet w=11600 l=12325
+ ad=0 pd=0 as=1.07648e+09 ps=203000 
M2733 N0701 Vdd Vdd GND efet w=7250 l=20300
+ ad=0 pd=0 as=0 ps=0 
M2734 GND L N0686 GND efet w=57275 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2735 GND L N0701 GND efet w=42775 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2736 Vdd Vdd N0546 GND efet w=13050 l=87000
+ ad=0 pd=0 as=0 ps=0 
M2737 N0546 N0342 GND GND efet w=12325 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2738 GND SUB_GROUP_6_ CY_ADAC GND efet w=14500 l=11600
+ ad=0 pd=0 as=-1.87289e+09 ps=440800 
M2739 GND ADD_GROUP_4_ CY_ADA GND efet w=11600 l=10875
+ ad=0 pd=0 as=2.07096e+09 ps=417600 
M2740 Vdd Vdd N0677 GND efet w=8700 l=34075
+ ad=0 pd=0 as=7.67412e+08 ps=171100 
M2741 N0685 clk1 N0701 GND efet w=21025 l=18850
+ ad=-1.7993e+09 pd=551000 as=0 ps=0 
M2742 CY_1 ADSR N0513 GND efet w=14500 l=11600
+ ad=1.91958e+09 pd=382800 as=0 ps=0 
M2743 S00729 Vdd Vdd GND efet w=5800 l=11600
+ ad=-1.76356e+09 pd=327700 as=0 ps=0 
M2744 S00724 Vdd Vdd GND efet w=6525 l=15225
+ ad=-1.4608e+09 pd=406000 as=0 ps=0 
M2745 CY N0415 N0860 GND efet w=15950 l=10150
+ ad=1.62734e+09 pd=307400 as=0 ps=0 
M2746 N0860 N0403 Vdd GND efet w=13775 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2747 CY_ADAC S00732 CY_ADAC GND efet w=60175 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2748 CY M12 N0470 GND efet w=7975 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2749 N0550 CY_ADA N0470 GND efet w=14500 l=11600
+ ad=-1.67691e+09 pd=1.2934e+06 as=0 ps=0 
M2750 N0470 Vdd Vdd GND efet w=10150 l=34800
+ ad=0 pd=0 as=0 ps=0 
M2751 N0470 N0855 GND GND efet w=41325 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2752 N0513 ADSL CY GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2753 D0 CY_IB CY_1 GND efet w=57275 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2754 GND N0342 CY_ADAC GND efet w=13775 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2755 CY_ADA S00734 CY_ADA GND efet w=79750 l=20300
+ ad=0 pd=0 as=0 ps=0 
M2756 N0861 ADC_CY CY GND efet w=10150 l=13050
+ ad=8.64127e+08 pd=200100 as=0 ps=0 
M2757 GND CY N0855 GND efet w=59450 l=11600
+ ad=0 pd=0 as=8.17873e+08 ps=171100 
M2758 N0855 Vdd Vdd GND efet w=10150 l=33350
+ ad=0 pd=0 as=0 ps=0 
M2759 N0846 ADSR CY GND efet w=7250 l=11600
+ ad=9.8397e+08 pd=223300 as=0 ps=0 
M2760 CY_ADAC S00732 Vdd GND efet w=6525 l=48575
+ ad=0 pd=0 as=0 ps=0 
M2761 GND N0342 CY_ADA GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2762 GND READ_ACC_3_ ACC_ADA GND efet w=14500 l=11600
+ ad=0 pd=0 as=4.92425e+08 ps=948300 
M2763 GND N0342 ACC_ADA GND efet w=15225 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2764 GND WRITE_CARRY_2_ ADC_CY GND efet w=13775 l=10875
+ ad=0 pd=0 as=3.7889e+08 ps=791700 
M2765 GND WRITE_ACC_1_ ADD_ACC GND efet w=15225 l=11600
+ ad=0 pd=0 as=1.24722e+09 ps=1.189e+06 
M2766 N0678 clk1 GND GND efet w=22475 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2767 N0686 clk1 N0675 GND efet w=46400 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2768 GND N0678 N0677 GND efet w=29000 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2769 GND N0699 N0678 GND efet w=24650 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2770 N0701 N0702 N0699 GND efet w=10150 l=11600
+ ad=0 pd=0 as=6.85415e+08 ps=153700 
M2771 N0676 N0677 Vdd GND efet w=41325 l=14500
+ ad=-3.95612e+08 pd=3.2074e+06 as=0 ps=0 
M2772 N0678 N0685 GND GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2773 GND N0678 N0676 GND efet w=45675 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2774 GND N0477 ADC_CY GND efet w=13050 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2775 GND N0477 ADD_ACC GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2776 ADD_ACC Vdd Vdd GND efet w=10150 l=65250
+ ad=0 pd=0 as=0 ps=0 
M2777 Vdd S00734 CY_ADA GND efet w=5800 l=58000
+ ad=0 pd=0 as=0 ps=0 
M2778 ADC_CY Vdd Vdd GND efet w=8700 l=79750
+ ad=0 pd=0 as=0 ps=0 
M2779 S00734 Vdd Vdd GND efet w=7250 l=11600
+ ad=-1.23583e+09 pd=394400 as=0 ps=0 
M2780 S00732 Vdd Vdd GND efet w=7975 l=10150
+ ad=-1.70889e+09 pd=321900 as=0 ps=0 
M2781 L clk1 N0707 GND efet w=10875 l=13050
+ ad=0 pd=0 as=8.6623e+08 ps=208800 
M2782 N0675 clk2 N0684 GND efet w=44950 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2783 N0684 N0685 GND GND efet w=56550 l=8700
+ ad=0 pd=0 as=0 ps=0 
M2784 N0705 N0707 GND GND efet w=59450 l=9425
+ ad=-1.92335e+09 pd=452400 as=0 ps=0 
M2785 N0705 L N0706 GND efet w=126150 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2786 GND POC N0705 GND efet w=60175 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2787 N0706 N0702 GND GND efet w=96425 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2788 N0705 Vdd Vdd GND efet w=15225 l=27550
+ ad=0 pd=0 as=0 ps=0 
M2789 GND N0705 N0704 GND efet w=37700 l=15950
+ ad=0 pd=0 as=1.08699e+09 ps=232000 
M2790 GND M12 N0550 GND efet w=10150 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2791 N0550 N0546 Vdd GND efet w=9425 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2792 GND N0452 CY_1 GND efet w=53650 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2793 CY_1 Vdd Vdd GND efet w=6525 l=29000
+ ad=0 pd=0 as=0 ps=0 
M2794 N0855 N0854 N0452 GND efet w=8700 l=10150
+ ad=0 pd=0 as=8.70435e+08 ps=197200 
M2795 N0550 CY_ADAC N0855 GND efet w=15950 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2796 GND SUB_GROUP_6_ N0937 GND efet w=13050 l=11600
+ ad=0 pd=0 as=-1.86237e+09 ps=542300 
M2797 N0937 M12 GND GND efet w=18125 l=9425
+ ad=0 pd=0 as=0 ps=0 
M2798 N0704 Vdd Vdd GND efet w=9425 l=38425
+ ad=0 pd=0 as=0 ps=0 
M2799 N0700 N0704 Vdd GND efet w=65975 l=12325
+ ad=-9.41381e+08 pd=4.5269e+06 as=0 ps=0 
M2800 GND M12 SUB_GROUP_6_ GND efet w=13775 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2801 N0886 N0550 N0894 GND efet w=59450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2802 N0548 N0550 N0549 GND efet w=61625 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2803 GND N0878 N0846 GND efet w=60900 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2804 Vdd Vdd N0350 GND efet w=7250 l=50750
+ ad=0 pd=0 as=-1.05712e+09 ps=661200 
M2805 GND N0849 N0346 GND efet w=58725 l=12325
+ ad=0 pd=0 as=-1.65217e+08 ps=1.6733e+06 
M2806 N0856 N0854 N0849 GND efet w=7975 l=12325
+ ad=7.75823e+08 pd=156600 as=9.65047e+08 ps=191400 
M2807 N0346 Vdd Vdd GND efet w=6525 l=32625
+ ad=0 pd=0 as=0 ps=0 
M2808 N0870 ACC_ADAC N0856 GND efet w=14500 l=13050
+ ad=-8.15573e+07 pd=806200 as=0 ps=0 
M2809 N0846 N0874 Vdd GND efet w=13050 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2810 N0894 N0870 GND GND efet w=44225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2811 GND CY_1 N0803 GND efet w=14500 l=17400
+ ad=0 pd=0 as=1.19001e+09 ps=272600 
M2812 N0745 N0725 GND GND efet w=29000 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2813 Vdd Vdd S00761 GND efet w=6525 l=11600
+ ad=0 pd=0 as=-2.00955e+09 ps=278400 
M2814 S00757 Vdd Vdd GND efet w=8700 l=13050
+ ad=1.9343e+09 pd=237800 as=0 ps=0 
M2815 GND _COM N0717 GND efet w=77575 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2816 Vdd S00761 N0745 GND efet w=5800 l=27550
+ ad=0 pd=0 as=0 ps=0 
M2817 N0725 clk1 N0724 GND efet w=15950 l=10150
+ ad=2.01419e+09 pd=406000 as=0 ps=0 
M2818 N0724 N0284 GND GND efet w=27550 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2819 N0284 clk2 A32 GND efet w=14500 l=11600
+ ad=5.90802e+08 pd=130500 as=1.43268e+09 ps=2.0387e+06 
M2820 Vdd Vdd N0724 GND efet w=8700 l=40600
+ ad=0 pd=0 as=0 ps=0 
M2821 N0288 A32 GND GND efet w=23200 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2822 GND DAA N0802 GND efet w=13050 l=11600
+ ad=0 pd=0 as=1.33298e+09 ps=278400 
M2823 N0818 N0803 GND GND efet w=28275 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2824 N0378 DAA N0818 GND efet w=29000 l=11600
+ ad=1.52011e+09 pd=310300 as=0 ps=0 
M2825 GND O_IB N0378 GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2826 N0350 KBP GND GND efet w=17400 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2827 N0856 Vdd Vdd GND efet w=10150 l=37700
+ ad=0 pd=0 as=0 ps=0 
M2828 N0803 N0356 N0819 GND efet w=28275 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2829 Vdd N0746 A32 GND efet w=38425 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2830 A32 N0727 GND GND efet w=39150 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2831 N0746 S00778 N0746 GND efet w=68150 l=6525
+ ad=1.36242e+09 pd=261000 as=0 ps=0 
M2832 N0746 N0727 GND GND efet w=34800 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2833 Vdd Vdd S00778 GND efet w=5800 l=13050
+ ad=0 pd=0 as=-2.04109e+09 ps=263900 
M2834 Vdd S00778 N0746 GND efet w=7250 l=26100
+ ad=0 pd=0 as=0 ps=0 
M2835 Vdd Vdd N0766 GND efet w=8700 l=43500
+ ad=0 pd=0 as=1.71354e+09 ps=391500 
M2836 Vdd Vdd N0751 GND efet w=7975 l=45675
+ ad=0 pd=0 as=1.75349e+09 ps=342200 
M2837 DCL_0 Vdd Vdd GND efet w=7250 l=44950
+ ad=1.81025e+09 pd=417600 as=0 ps=0 
M2838 GND N0348 N0819 GND efet w=34800 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2839 N0819 N0347 GND GND efet w=37700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2840 N0803 Vdd Vdd GND efet w=5800 l=50750
+ ad=0 pd=0 as=0 ps=0 
M2841 N0403 Vdd Vdd GND efet w=6525 l=33350
+ ad=0 pd=0 as=0 ps=0 
M2842 N0802 Vdd Vdd GND efet w=6525 l=70325
+ ad=0 pd=0 as=0 ps=0 
M2843 N0354 Vdd Vdd GND efet w=7250 l=46400
+ ad=-1.98432e+09 pd=484300 as=0 ps=0 
M2844 N0363 Vdd Vdd GND efet w=9425 l=50025
+ ad=-3.12832e+08 pd=762700 as=0 ps=0 
M2845 N0370 Vdd Vdd GND efet w=7975 l=42775
+ ad=-1.44818e+09 pd=582900 as=0 ps=0 
M2846 Vdd Vdd N0345 GND efet w=7975 l=51475
+ ad=0 pd=0 as=1.81255e+08 ps=887400 
M2847 N0378 Vdd Vdd GND efet w=7250 l=47850
+ ad=0 pd=0 as=0 ps=0 
M2848 N0377 N0378 N0376 GND efet w=34075 l=12325
+ ad=-5.81952e+08 pd=678600 as=0 ps=0 
M2849 GND N0346 ACC_0 GND efet w=21750 l=11600
+ ad=0 pd=0 as=-4.80592e+08 ps=1.6211e+06 
M2850 CY_1 ADSL ACC_0 GND efet w=7250 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2851 GND ACC_0 N0856 GND efet w=61625 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2852 GND M12 N0870 GND efet w=13050 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2853 N0471 Vdd Vdd GND efet w=9425 l=36975
+ ad=0 pd=0 as=0 ps=0 
M2854 N0346 ACB_IB D0 GND efet w=43500 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2855 ACC_0 Vdd Vdd GND efet w=8700 l=44950
+ ad=0 pd=0 as=0 ps=0 
M2856 GND N0846 ADD_0 GND efet w=42775 l=10875
+ ad=0 pd=0 as=1.42638e+09 ps=1.8096e+06 
M2857 ACC_0 M12 N0471 GND efet w=7250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2858 N0846 ADD_ACC ACC_0 GND efet w=10150 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2859 GND N0878 N0874 GND efet w=12325 l=13775
+ ad=0 pd=0 as=5.95007e+08 ps=145000 
M2860 N0878 N0887 N0886 GND efet w=60900 l=12325
+ ad=1.18371e+09 pd=240700 as=0 ps=0 
M2861 N0548 N0870 GND GND efet w=62350 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2862 N0549 N0887 GND GND efet w=50025 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2863 GND N0856 N0471 GND efet w=36250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2864 N0874 Vdd Vdd GND efet w=5800 l=59450
+ ad=0 pd=0 as=0 ps=0 
M2865 N0549 N0870 N0911 GND efet w=68875 l=17400
+ ad=0 pd=0 as=1.54113e+09 ps=333500 
M2866 N0911 N0887 N0548 GND efet w=55825 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2867 _TMP_0 N0940 GND GND efet w=22475 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2868 GND N0705 N0700 GND efet w=95700 l=8700
+ ad=0 pd=0 as=0 ps=0 
M2869 _TMP_0 N0937 N0887 GND efet w=13775 l=10875
+ ad=0 pd=0 as=4.52478e+08 ps=933800 
M2870 Vdd N0939 _TMP_0 GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2871 Vdd Vdd N0911 GND efet w=5800 l=66700
+ ad=0 pd=0 as=0 ps=0 
M2872 N0847 ADSR ACC_0 GND efet w=10150 l=11600
+ ad=9.98687e+08 pd=217500 as=0 ps=0 
M2873 N0878 Vdd Vdd GND efet w=7250 l=53650
+ ad=0 pd=0 as=0 ps=0 
M2874 N0898 N0553 N0878 GND efet w=36250 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2875 GND N0870 N0898 GND efet w=35525 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2876 N0898 N0550 GND GND efet w=43500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2877 GND N0887 N0898 GND efet w=35525 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2878 N0915 N0911 GND GND efet w=11600 l=11600
+ ad=4.66755e+08 pd=116000 as=0 ps=0 
M2879 Vdd Vdd N0915 GND efet w=7250 l=63075
+ ad=0 pd=0 as=0 ps=0 
M2880 D0 ADD_IB N0846 GND efet w=40600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2881 N0870 ACC_ADA N0471 GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2882 N0940 Vdd Vdd GND efet w=6525 l=45675
+ ad=9.6715e+08 pd=194300 as=0 ps=0 
M2883 GND N0939 N0940 GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2884 TMP_0 SUB_GROUP_6_ N0887 GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2885 TMP_0 N0940 Vdd GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2886 GND N0939 TMP_0 GND efet w=23200 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2887 Vdd M12 N0604 GND efet w=7250 l=11600
+ ad=0 pd=0 as=1.0071e+09 ps=211700 
M2888 N0553 N0915 GND GND efet w=20300 l=10150
+ ad=1.34394e+09 pd=1.0933e+06 as=0 ps=0 
M2889 D0 N0964 N0604 GND efet w=12325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2890 GND N0604 N0939 GND efet w=42050 l=13775
+ ad=0 pd=0 as=1.12273e+09 ps=237800 
M2891 N0939 S00762 N0939 GND efet w=51475 l=19575
+ ad=0 pd=0 as=0 ps=0 
M2892 N0939 S00762 Vdd GND efet w=5800 l=47850
+ ad=0 pd=0 as=0 ps=0 
M2893 Vdd N0911 N0553 GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2894 GND N0884 N0847 GND efet w=63075 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2895 Vdd S00764 ACC_ADAC GND efet w=5800 l=45675
+ ad=0 pd=0 as=0 ps=0 
M2896 ACC_ADAC S00764 ACC_ADAC GND efet w=79025 l=5075
+ ad=0 pd=0 as=0 ps=0 
M2897 ADD_0 Vdd Vdd GND efet w=8700 l=46400
+ ad=0 pd=0 as=0 ps=0 
M2898 Vdd Vdd N0377 GND efet w=8700 l=43500
+ ad=0 pd=0 as=0 ps=0 
M2899 GND DCL_0 N0751 GND efet w=35525 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2900 N0766 N0351 GND GND efet w=22475 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2901 GND DCL_0 N0716 GND efet w=47850 l=10150
+ ad=0 pd=0 as=-6.3872e+08 ps=684400 
M2902 N0751 N0766 N0767 GND efet w=12325 l=12325
+ ad=0 pd=0 as=1.55165e+09 ps=350900 
M2903 DCL_0 POC GND GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2904 GND N0350 N0376 GND efet w=37700 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2905 GND N0767 DCL_0 GND efet w=50750 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2906 N0345 N0350 GND GND efet w=17400 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2907 N0354 N0350 GND GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2908 GND N0350 N0363 GND efet w=17400 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2909 N0370 N0350 GND GND efet w=18125 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2910 Vdd Vdd N0371 GND efet w=5800 l=59450
+ ad=0 pd=0 as=-1.87499e+09 ps=466900 
M2911 GND N0847 ADD_0 GND efet w=39875 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2912 N0847 ADD_IB D1 GND efet w=39875 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2913 Vdd Vdd S00764 GND efet w=5800 l=11600
+ ad=0 pd=0 as=-1.95068e+09 ps=298700 
M2914 N0847 N0875 Vdd GND efet w=15950 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2915 Vdd Vdd S00767 GND efet w=9425 l=10875
+ ad=0 pd=0 as=-1.74674e+09 ps=333500 
M2916 D1 ACB_IB N0347 GND efet w=39875 l=11600
+ ad=0 pd=0 as=1.13929e+07 ps=1.7516e+06 
M2917 N0871 ACC_ADAC N0472 GND efet w=14500 l=13050
+ ad=-1.6623e+06 pd=843900 as=0 ps=0 
M2918 N0888 N0553 N0895 GND efet w=57275 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2919 N0895 N0871 GND GND efet w=58000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2920 N0875 N0889 N0888 GND efet w=60175 l=11600
+ ad=9.86073e+08 pd=240700 as=0 ps=0 
M2921 GND N0347 ACC_0 GND efet w=23200 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2922 N0472 Vdd Vdd GND efet w=10875 l=35525
+ ad=0 pd=0 as=0 ps=0 
M2923 N0472 M12 ACC_1 GND efet w=8700 l=11600
+ ad=0 pd=0 as=1.21314e+09 ps=234900 
M2924 N0472 N0857 GND GND efet w=36975 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2925 N0846 ADSL ACC_1 GND efet w=8700 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2926 GND N0875 N0884 GND efet w=12325 l=10875
+ ad=0 pd=0 as=9.94482e+08 ps=200100 
M2927 N0551 N0553 N0552 GND efet w=60900 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2928 N0551 N0871 GND GND efet w=65975 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2929 N0552 N0889 GND GND efet w=48575 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2930 N0370 N0371 GND GND efet w=17400 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2931 N0371 N0346 GND GND efet w=14500 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2932 Vdd Vdd N0364 GND efet w=6525 l=68875
+ ad=0 pd=0 as=-1.83084e+09 ps=519100 
M2933 N0726 N0285 GND GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2934 N0285 clk2 A22 GND efet w=13775 l=12325
+ ad=5.67675e+08 pd=127600 as=0 ps=0 
M2935 N0727 clk1 N0726 GND efet w=14500 l=11600
+ ad=2.00158e+09 pd=408900 as=0 ps=0 
M2936 Vdd Vdd N0726 GND efet w=7975 l=37700
+ ad=0 pd=0 as=0 ps=0 
M2937 GND DCL_1 N0716 GND efet w=49300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2938 N0371 N0351 N0767 GND efet w=12325 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2939 N0912 N0889 N0551 GND efet w=57275 l=13775
+ ad=1.22786e+09 pd=292900 as=0 ps=0 
M2940 N0552 N0871 N0912 GND efet w=67425 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2941 N0912 S00767 N0912 GND efet w=50025 l=23200
+ ad=0 pd=0 as=0 ps=0 
M2942 S00762 Vdd Vdd GND efet w=8700 l=11600
+ ad=-1.99063e+09 pd=281300 as=0 ps=0 
M2943 GND N0342 N0964 GND efet w=23925 l=13775
+ ad=0 pd=0 as=-1.40193e+09 ps=556800 
M2944 N0964 Vdd Vdd GND efet w=10875 l=35525
+ ad=0 pd=0 as=0 ps=0 
M2945 GND N0871 N0899 GND efet w=34800 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2946 GND ACC_1 N0857 GND efet w=59450 l=11600
+ ad=0 pd=0 as=8.1577e+08 ps=168200 
M2947 N0847 ADD_ACC ACC_1 GND efet w=8700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2948 N0884 Vdd Vdd GND efet w=10150 l=47125
+ ad=0 pd=0 as=0 ps=0 
M2949 N0857 Vdd Vdd GND efet w=10150 l=33350
+ ad=0 pd=0 as=0 ps=0 
M2950 N0848 ADSR ACC_1 GND efet w=7975 l=13775
+ ad=1.14586e+09 pd=252300 as=0 ps=0 
M2951 N0347 Vdd Vdd GND efet w=7250 l=33350
+ ad=0 pd=0 as=0 ps=0 
M2952 GND N0850 N0347 GND efet w=58000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2953 N0857 N0854 N0850 GND efet w=8700 l=11600
+ ad=0 pd=0 as=9.12485e+08 ps=188500 
M2954 Vdd M12 N0871 GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2955 N0875 Vdd Vdd GND efet w=8700 l=65250
+ ad=0 pd=0 as=0 ps=0 
M2956 N0899 N0556 N0875 GND efet w=35525 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2957 N0899 N0553 GND GND efet w=43500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2958 GND N0889 N0899 GND efet w=36250 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2959 N0871 ACC_ADA N0857 GND efet w=15950 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2960 N0345 N0346 GND GND efet w=18125 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2961 GND N0346 N0354 GND efet w=14500 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2962 GND N0346 N0363 GND efet w=19575 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2963 N0288 A22 GND GND efet w=23200 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2964 GND N0765 DCL_1 GND efet w=39150 l=11600
+ ad=0 pd=0 as=1.6021e+09 ps=365400 
M2965 GND N0346 N0376 GND efet w=36250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2966 GND N0879 N0848 GND efet w=60900 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2967 Vdd S00767 N0912 GND efet w=5800 l=51475
+ ad=0 pd=0 as=0 ps=0 
M2968 TMP_1 N0937 N0889 GND efet w=14500 l=11600
+ ad=0 pd=0 as=3.15815e+08 ps=916400 
M2969 _TMP_1 N0942 GND GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2970 N0672 D2 GND GND efet w=57275 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2971 d2 POC GND GND efet w=29725 l=13775
+ ad=4.60888e+08 pd=829400 as=0 ps=0 
M2972 Vdd Vdd N0672 GND efet w=10875 l=40600
+ ad=0 pd=0 as=0 ps=0 
M2973 S00765 Vdd Vdd GND efet w=7250 l=15950
+ ad=-2.02006e+09 pd=266800 as=0 ps=0 
M2974 S00766 Vdd Vdd GND efet w=7250 l=15225
+ ad=-2.06842e+09 pd=269700 as=0 ps=0 
M2975 N0690 S00765 N0690 GND efet w=71050 l=9425
+ ad=1.20561e+09 pd=1.7313e+06 as=0 ps=0 
M2976 Vdd S00766 N0692 GND efet w=10150 l=12325
+ ad=0 pd=0 as=4.78588e+08 ps=2.4563e+06 
M2977 N0690 S00765 Vdd GND efet w=12325 l=18125
+ ad=0 pd=0 as=0 ps=0 
M2978 Vdd N0941 _TMP_1 GND efet w=13775 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2979 N0691 N0702 N0672 GND efet w=27550 l=12325
+ ad=-1.26947e+09 pd=585800 as=0 ps=0 
M2980 N0942 Vdd Vdd GND efet w=6525 l=47125
+ ad=9.69252e+08 pd=200100 as=0 ps=0 
M2981 N0916 N0912 GND GND efet w=13050 l=10150
+ ad=4.64653e+08 pd=116000 as=0 ps=0 
M2982 Vdd Vdd N0916 GND efet w=7250 l=63075
+ ad=0 pd=0 as=0 ps=0 
M2983 GND N0941 N0942 GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2984 N0692 S00766 N0692 GND efet w=41325 l=47850
+ ad=0 pd=0 as=0 ps=0 
M2985 Vdd M12 N0605 GND efet w=7975 l=10150
+ ad=0 pd=0 as=9.77663e+08 ps=208800 
M2986 TMP_1 N0942 Vdd GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2987 _TMP_1 SUB_GROUP_6_ N0889 GND efet w=18125 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2988 GND N0941 TMP_1 GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2989 N0690 N0700 GND GND efet w=262450 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2990 D1 N0964 N0605 GND efet w=12325 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2991 N0556 N0916 GND GND efet w=20300 l=10150
+ ad=1.2304e+09 pd=1.073e+06 as=0 ps=0 
M2992 N0692 N0700 GND GND efet w=228375 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2993 GND N0605 N0941 GND efet w=41325 l=18125
+ ad=0 pd=0 as=1.10802e+09 ps=217500 
M2994 Vdd N0912 N0556 GND efet w=14500 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2995 N0941 S00781 N0941 GND efet w=50025 l=20300
+ ad=0 pd=0 as=0 ps=0 
M2996 N0941 S00781 Vdd GND efet w=5800 l=43500
+ ad=0 pd=0 as=0 ps=0 
M2997 GND N0851 N0348 GND efet w=56550 l=11600
+ ad=0 pd=0 as=1.92208e+08 ps=1.7429e+06 
M2998 N0858 N0854 N0851 GND efet w=7250 l=13050
+ ad=7.7372e+08 pd=156600 as=9.251e+08 ps=185600 
M2999 N0348 Vdd Vdd GND efet w=8700 l=29000
+ ad=0 pd=0 as=0 ps=0 
M3000 Vdd N0747 A22 GND efet w=41325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3001 A22 N0729 GND GND efet w=37700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3002 GND POC DCL_1 GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3003 DCL_1 Vdd Vdd GND efet w=7250 l=49300
+ ad=0 pd=0 as=0 ps=0 
M3004 N0364 N0351 N0765 GND efet w=12325 l=15225
+ ad=0 pd=0 as=-1.7993e+09 ps=542300 
M3005 GND N0364 N0363 GND efet w=17400 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3006 GND N0347 N0345 GND efet w=24650 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3007 N0354 N0347 GND GND efet w=13775 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3008 N0364 N0347 GND GND efet w=14500 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3009 N0872 ACC_ADAC N0858 GND efet w=15225 l=12325
+ ad=-2.03502e+08 pd=841000 as=0 ps=0 
M3010 N0848 N0876 Vdd GND efet w=13775 l=15225
+ ad=0 pd=0 as=0 ps=0 
M3011 N0858 Vdd Vdd GND efet w=10150 l=41325
+ ad=0 pd=0 as=0 ps=0 
M3012 GND N0347 N0370 GND efet w=18850 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3013 GND N0347 N0376 GND efet w=36250 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3014 GND DCL_1 N0750 GND efet w=23200 l=11600
+ ad=0 pd=0 as=9.9238e+08 ps=194300 
M3015 N0750 Vdd Vdd GND efet w=7250 l=52200
+ ad=0 pd=0 as=0 ps=0 
M3016 N0747 S00800 N0747 GND efet w=69600 l=5800
+ ad=1.33719e+09 pd=263900 as=0 ps=0 
M3017 N0747 N0729 GND GND efet w=32625 l=15225
+ ad=0 pd=0 as=0 ps=0 
M3018 Vdd Vdd S00800 GND efet w=6525 l=13775
+ ad=0 pd=0 as=2.14455e+09 ps=255200 
M3019 Vdd S00800 N0747 GND efet w=5800 l=24650
+ ad=0 pd=0 as=0 ps=0 
M3020 N0750 N0766 N0765 GND efet w=10150 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3021 Vdd Vdd N0355 GND efet w=6525 l=73225
+ ad=0 pd=0 as=-1.80561e+09 ps=493000 
M3022 N0355 N0351 N0768 GND efet w=10150 l=10150
+ ad=0 pd=0 as=-1.73833e+09 ps=507500 
M3023 N0354 N0355 GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3024 N0355 N0348 GND GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3025 GND N0348 ACC_0 GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3026 N0847 ADSL ACC_2 GND efet w=7250 l=14500
+ ad=0 pd=0 as=1.20473e+09 ps=252300 
M3027 GND ACC_2 N0858 GND efet w=64525 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3028 N0473 Vdd Vdd GND efet w=12325 l=36975
+ ad=0 pd=0 as=0 ps=0 
M3029 GND N0848 ADD_0 GND efet w=42775 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3030 N0348 ACB_IB D2 GND efet w=39150 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3031 N0848 ADD_ACC ACC_2 GND efet w=7975 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3032 ACC_2 M12 N0473 GND efet w=7975 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3033 GND N0858 N0473 GND efet w=36250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3034 N0890 N0556 N0896 GND efet w=59450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3035 N0896 N0872 GND GND efet w=60900 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3036 N0879 N0891 N0890 GND efet w=65250 l=10875
+ ad=1.10592e+09 pd=243600 as=0 ps=0 
M3037 N0554 N0872 GND GND efet w=64525 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3038 GND N0879 N0876 GND efet w=10150 l=12325
+ ad=0 pd=0 as=6.93825e+08 ps=147900 
M3039 GND M12 N0872 GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3040 N0514 ADSR ACC_2 GND efet w=9425 l=12325
+ ad=1.14586e+09 pd=252300 as=0 ps=0 
M3041 N0555 N0891 GND GND efet w=52925 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3042 N0555 N0872 N0913 GND efet w=68150 l=14500
+ ad=0 pd=0 as=1.37504e+09 ps=319000 
M3043 N0913 N0891 N0554 GND efet w=56550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3044 N0876 Vdd Vdd GND efet w=8700 l=65975
+ ad=0 pd=0 as=0 ps=0 
M3045 D2 ADD_IB N0848 GND efet w=42775 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3046 N0872 ACC_ADA N0473 GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3047 N0879 Vdd Vdd GND efet w=9425 l=57275
+ ad=0 pd=0 as=0 ps=0 
M3048 GND DCL_2 N0716 GND efet w=43500 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3049 N0728 N0286 GND GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3050 N0729 clk1 N0728 GND efet w=13775 l=12325
+ ad=1.99317e+09 pd=397300 as=0 ps=0 
M3051 N0286 clk2 A12 GND efet w=15950 l=11600
+ ad=6.2234e+08 pd=136300 as=6.40921e+08 ps=3.4829e+06 
M3052 GND N0768 DCL_2 GND efet w=42050 l=10150
+ ad=0 pd=0 as=1.98686e+09 ps=406000 
M3053 GND N0348 N0345 GND efet w=18850 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3054 GND N0348 N0363 GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3055 GND N0348 N0370 GND efet w=19575 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3056 GND N0348 N0376 GND efet w=36250 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3057 N0900 N0559 N0879 GND efet w=34800 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3058 GND N0872 N0900 GND efet w=36250 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3059 N0900 N0556 GND GND efet w=43500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3060 GND N0891 N0900 GND efet w=40600 l=13050
+ ad=0 pd=0 as=0 ps=0 
M3061 ACC_ADA S00803 ACC_ADA GND efet w=81200 l=4350
+ ad=0 pd=0 as=0 ps=0 
M3062 N0554 N0556 N0555 GND efet w=60900 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3063 GND N0691 N0690 GND efet w=97875 l=9425
+ ad=0 pd=0 as=0 ps=0 
M3064 D2 N0964 N0606 GND efet w=19575 l=17400
+ ad=0 pd=0 as=1.70723e+09 ps=333500 
M3065 GND N0690 N0692 GND efet w=73950 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3066 S00781 Vdd Vdd GND efet w=9425 l=12325
+ ad=-1.94647e+09 pd=275500 as=0 ps=0 
M3067 Vdd Vdd N0913 GND efet w=5800 l=58000
+ ad=0 pd=0 as=0 ps=0 
M3068 _TMP_2 N0944 GND GND efet w=22475 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3069 _TMP_2 N0937 N0891 GND efet w=15950 l=10875
+ ad=0 pd=0 as=3.76788e+08 ps=945400 
M3070 Vdd N0943 _TMP_2 GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M3071 GND N0692 d2 GND efet w=1202775 l=7250
+ ad=0 pd=0 as=0 ps=0 
M3072 N0606 M12 Vdd GND efet w=8700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3073 N0665 N0676 GND GND efet w=26100 l=13050
+ ad=1.37714e+09 pd=269700 as=0 ps=0 
M3074 N0917 N0913 GND GND efet w=13050 l=10875
+ ad=5.25625e+08 pd=116000 as=0 ps=0 
M3075 Vdd Vdd N0917 GND efet w=5800 l=63800
+ ad=0 pd=0 as=0 ps=0 
M3076 N0559 N0917 GND GND efet w=20300 l=11600
+ ad=1.27245e+09 pd=1.1107e+06 as=0 ps=0 
M3077 Vdd N0913 N0559 GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3078 Vdd Vdd S00804 GND efet w=5800 l=11600
+ ad=0 pd=0 as=-1.86448e+09 ps=298700 
M3079 N0944 Vdd Vdd GND efet w=7975 l=44225
+ ad=1.04074e+09 pd=208800 as=0 ps=0 
M3080 GND N0943 N0944 GND efet w=13775 l=15225
+ ad=0 pd=0 as=0 ps=0 
M3081 TMP_2 N0944 Vdd GND efet w=15950 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3082 GND N0943 TMP_2 GND efet w=19575 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3083 TMP_2 SUB_GROUP_6_ N0891 GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3084 d2 N0690 Vdd GND efet w=640175 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3085 Vdd Vdd N0665 GND efet w=11600 l=52200
+ ad=0 pd=0 as=0 ps=0 
M3086 N0665 N0666 GND GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M3087 N0943 S00801 Vdd GND efet w=8700 l=53650
+ ad=1.24678e+09 pd=220400 as=0 ps=0 
M3088 Vdd Vdd N0349 GND efet w=6525 l=61625
+ ad=0 pd=0 as=-1.78458e+09 ps=513300 
M3089 Vdd S00803 ACC_ADA GND efet w=6525 l=45675
+ ad=0 pd=0 as=0 ps=0 
M3090 Vdd Vdd N0728 GND efet w=7250 l=38425
+ ad=0 pd=0 as=0 ps=0 
M3091 N0288 A12 GND GND efet w=22475 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3092 DCL_2 Vdd Vdd GND efet w=8700 l=43500
+ ad=0 pd=0 as=0 ps=0 
M3093 N0749 Vdd Vdd GND efet w=7250 l=43500
+ ad=1.21104e+09 pd=240700 as=0 ps=0 
M3094 Vdd N0748 A12 GND efet w=39150 l=13050
+ ad=0 pd=0 as=0 ps=0 
M3095 GND POC DCL_2 GND efet w=26100 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3096 GND DCL_2 N0749 GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3097 A12 N0731 GND GND efet w=38425 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3098 N0748 S00814 N0748 GND efet w=68150 l=5800
+ ad=8.76743e+08 pd=174000 as=0 ps=0 
M3099 N0748 N0731 GND GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3100 Vdd Vdd S00814 GND efet w=5800 l=12325
+ ad=0 pd=0 as=-2.11888e+09 ps=263900 
M3101 N0768 N0766 N0749 GND efet w=9425 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3102 GND N0349 N0345 GND efet w=19575 l=13050
+ ad=0 pd=0 as=0 ps=0 
M3103 N0354 N0356 GND GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3104 N0349 N0356 GND GND efet w=11600 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3105 GND N0514 ADD_0 GND efet w=41325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3106 GND N0356 N0363 GND efet w=17400 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3107 GND N0356 N0370 GND efet w=19575 l=15225
+ ad=0 pd=0 as=0 ps=0 
M3108 GND N0356 N0376 GND efet w=33350 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3109 Vdd S00814 N0748 GND efet w=5800 l=26100
+ ad=0 pd=0 as=0 ps=0 
M3110 N0514 ADD_IB D3 GND efet w=40600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3111 Vdd Vdd S00803 GND efet w=5800 l=10150
+ ad=0 pd=0 as=-1.8813e+09 ps=319000 
M3112 N0514 N0877 Vdd GND efet w=19575 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3113 D3 ACB_IB N0356 GND efet w=40600 l=11600
+ ad=0 pd=0 as=-1.61594e+09 ps=1.4529e+06 
M3114 N0873 ACC_ADAC N0474 GND efet w=15950 l=13775
+ ad=1.2659e+08 pd=855500 as=0 ps=0 
M3115 GND N0377 N0358 GND efet w=64525 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3116 GND N0345 N0358 GND efet w=72500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3117 N0358 N0354 GND GND efet w=66700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3118 GND N0363 N0358 GND efet w=74675 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3119 N0358 N0370 GND GND efet w=60175 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3120 N0358 Vdd Vdd GND efet w=6525 l=65975
+ ad=0 pd=0 as=0 ps=0 
M3121 N0714 S00818 N0714 GND efet w=76850 l=7250
+ ad=-1.30521e+09 pd=545200 as=0 ps=0 
M3122 N0714 N0749 GND GND efet w=45675 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3123 N0731 clk1 N0730 GND efet w=13775 l=10150
+ ad=1.99107e+09 pd=394400 as=0 ps=0 
M3124 N0730 N0287 GND GND efet w=29000 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3125 Vdd Vdd N0730 GND efet w=7975 l=39150
+ ad=0 pd=0 as=0 ps=0 
M3126 N0287 clk2 N0288 GND efet w=13050 l=11600
+ ad=5.90802e+08 pd=127600 as=0 ps=0 
M3127 GND _COM N0714 GND efet w=45675 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3128 Vdd Vdd S00818 GND efet w=7975 l=12325
+ ad=0 pd=0 as=-2.01586e+09 ps=269700 
M3129 Vdd S00818 N0714 GND efet w=10150 l=24650
+ ad=0 pd=0 as=0 ps=0 
M3130 N0366 Vdd Vdd GND efet w=5800 l=66700
+ ad=0 pd=0 as=0 ps=0 
M3131 Vdd Vdd N0288 GND efet w=8700 l=34800
+ ad=0 pd=0 as=0 ps=0 
M3132 N0715 S00825 N0715 GND efet w=76850 l=10150
+ ad=-7.71177e+08 pd=684400 as=0 ps=0 
M3133 N0715 N0750 GND GND efet w=44950 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3134 Vdd N0714 cm_ram3 GND efet w=142100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3135 N0734 N0714 GND GND efet w=47850 l=18850
+ ad=-6.53437e+08 pd=658300 as=0 ps=0 
M3136 GND _COM N0715 GND efet w=43500 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3137 N0366 N0354 GND GND efet w=61625 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3138 GND N0363 N0366 GND efet w=59450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3139 N0366 N0370 GND GND efet w=60900 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3140 GND N0377 N0366 GND efet w=59450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3141 GND N0403 N0358 GND efet w=60900 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3142 GND N0356 ACC_0 GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3143 N0474 Vdd Vdd GND efet w=10875 l=35525
+ ad=0 pd=0 as=0 ps=0 
M3144 N0356 N0852 GND GND efet w=53650 l=13050
+ ad=0 pd=0 as=0 ps=0 
M3145 N0356 Vdd Vdd GND efet w=8700 l=34800
+ ad=0 pd=0 as=0 ps=0 
M3146 N0366 TCS GND GND efet w=60175 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3147 Vdd Vdd S00825 GND efet w=7975 l=12325
+ ad=0 pd=0 as=-2.01165e+09 ps=269700 
M3148 Vdd N0715 cm_ram2 GND efet w=141375 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3149 Vdd Vdd N0734 GND efet w=8700 l=20300
+ ad=0 pd=0 as=0 ps=0 
M3150 Vdd Vdd N0735 GND efet w=9425 l=19575
+ ad=0 pd=0 as=-7.29127e+08 ps=669900 
M3151 GND N0715 N0735 GND efet w=40600 l=13050
+ ad=0 pd=0 as=0 ps=0 
M3152 Vdd S00825 N0715 GND efet w=10150 l=24650
+ ad=0 pd=0 as=0 ps=0 
M3153 N0359 Vdd Vdd GND efet w=6525 l=61625
+ ad=0 pd=0 as=0 ps=0 
M3154 GND N0345 N0359 GND efet w=61625 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3155 N0357 Vdd Vdd GND efet w=6525 l=68150
+ ad=0 pd=0 as=0 ps=0 
M3156 N0716 S00833 N0716 GND efet w=79025 l=6525
+ ad=0 pd=0 as=0 ps=0 
M3157 cm_ram2 N0735 GND GND efet w=263900 l=14500
+ ad=0 pd=0 as=0 ps=0 
M3158 cm_ram3 N0734 GND GND efet w=263900 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3159 GND _COM N0713 GND efet w=43500 l=13050
+ ad=0 pd=0 as=-5.14672e+08 ps=733700 
M3160 N0716 _COM GND GND efet w=59450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3161 N0713 S00834 N0713 GND efet w=75400 l=5800
+ ad=0 pd=0 as=0 ps=0 
M3162 S00834 Vdd Vdd GND efet w=7975 l=12325
+ ad=1.8544e+09 pd=269700 as=0 ps=0 
M3163 N0713 N0751 GND GND efet w=47125 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3164 N0359 N0370 GND GND efet w=65975 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3165 GND N0377 N0359 GND efet w=60175 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3166 D2 N0415 N0366 GND efet w=49300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3167 D3 N0415 N0358 GND efet w=49300 l=14500
+ ad=0 pd=0 as=0 ps=0 
M3168 N0359 TCS GND GND efet w=59450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3169 Vdd Vdd S00833 GND efet w=7975 l=12325
+ ad=0 pd=0 as=-2.02847e+09 ps=284200 
M3170 Vdd S00833 N0716 GND efet w=10875 l=23925
+ ad=0 pd=0 as=0 ps=0 
M3171 N0713 S00834 Vdd GND efet w=9425 l=22475
+ ad=0 pd=0 as=0 ps=0 
M3172 GND N0345 N0357 GND efet w=62350 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3173 GND N0363 N0357 GND efet w=63800 l=15950
+ ad=0 pd=0 as=0 ps=0 
M3174 GND N0377 N0357 GND efet w=60175 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3175 D1 N0415 N0359 GND efet w=50750 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3176 D0 N0415 N0357 GND efet w=55825 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3177 N0474 M12 ACC_3 GND efet w=8700 l=11600
+ ad=0 pd=0 as=1.18791e+09 ps=243600 
M3178 N0474 N0859 GND GND efet w=36250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3179 N0848 ADSL ACC_3 GND efet w=8700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3180 GND N0885 N0514 GND efet w=65975 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3181 GND N0606 N0943 GND efet w=41325 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3182 N0897 N0873 GND GND efet w=60175 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3183 GND N0877 N0885 GND efet w=13775 l=10150
+ ad=0 pd=0 as=9.39817e+08 ps=208800 
M3184 N0892 N0559 N0897 GND efet w=56550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3185 N0877 N0893 N0892 GND efet w=65250 l=10150
+ ad=9.69252e+08 pd=258100 as=0 ps=0 
M3186 N0557 N0873 GND GND efet w=76125 l=19575
+ ad=0 pd=0 as=0 ps=0 
M3187 GND N0893 N0558 GND efet w=61625 l=28275
+ ad=0 pd=0 as=0 ps=0 
M3188 GND ACC_3 N0859 GND efet w=58725 l=13775
+ ad=0 pd=0 as=8.17873e+08 ps=165300 
M3189 N0514 ADD_ACC ACC_3 GND efet w=9425 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3190 N0859 Vdd Vdd GND efet w=9425 l=35525
+ ad=0 pd=0 as=0 ps=0 
M3191 N0514 ADSL N0513 GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3192 N0859 N0854 N0852 GND efet w=7250 l=13050
+ ad=0 pd=0 as=1.37924e+09 ps=278400 
M3193 N0513 ADSR ACC_3 GND efet w=13050 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3194 N0914 N0893 N0557 GND efet w=55825 l=12325
+ ad=1.42129e+09 pd=313200 as=0 ps=0 
M3195 GND N0873 N0901 GND efet w=35525 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3196 N0885 Vdd Vdd GND efet w=9425 l=54375
+ ad=0 pd=0 as=0 ps=0 
M3197 Vdd M12 N0873 GND efet w=13775 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3198 N0901 N0861 N0877 GND efet w=37700 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3199 N0877 Vdd Vdd GND efet w=7975 l=64525
+ ad=0 pd=0 as=0 ps=0 
M3200 N0873 ACC_ADA N0859 GND efet w=15950 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3201 N0558 N0873 N0914 GND efet w=65975 l=16675
+ ad=0 pd=0 as=0 ps=0 
M3202 N0901 N0559 GND GND efet w=43500 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3203 GND N0893 N0901 GND efet w=37700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3204 N0557 N0559 N0558 GND efet w=58000 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3205 N0943 S00801 N0943 GND efet w=46400 l=21025
+ ad=0 pd=0 as=0 ps=0 
M3206 N0914 S00804 N0914 GND efet w=57275 l=34075
+ ad=0 pd=0 as=0 ps=0 
M3207 S00801 Vdd Vdd GND efet w=12325 l=13050
+ ad=-1.94437e+09 pd=287100 as=0 ps=0 
M3208 D2 N0666 GND GND efet w=49300 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3209 Vdd N0665 D2 GND efet w=39875 l=15225
+ ad=0 pd=0 as=0 ps=0 
M3210 Vdd S00804 N0914 GND efet w=5075 l=52200
+ ad=0 pd=0 as=0 ps=0 
M3211 Vdd Vdd N0666 GND efet w=10150 l=39150
+ ad=0 pd=0 as=1.43391e+09 ps=252300 
M3212 _TMP_3 N0946 GND GND efet w=21025 l=13050
+ ad=0 pd=0 as=0 ps=0 
M3213 N0666 d2 GND GND efet w=71050 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3214 _TMP_3 SUB_GROUP_6_ N0893 GND efet w=14500 l=11600
+ ad=0 pd=0 as=5.44988e+08 ps=928000 
M3215 N0666 N0676 GND GND efet w=44950 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3216 Vdd N0945 _TMP_3 GND efet w=13775 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3217 N0918 N0914 GND GND efet w=12325 l=12325
+ ad=5.44548e+08 pd=121800 as=0 ps=0 
M3218 Vdd Vdd N0918 GND efet w=5800 l=63800
+ ad=0 pd=0 as=0 ps=0 
M3219 N0861 N0918 GND GND efet w=18850 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3220 N0946 Vdd Vdd GND efet w=8700 l=43500
+ ad=9.86073e+08 pd=197200 as=0 ps=0 
M3221 GND N0945 N0946 GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3222 Vdd M12 N0607 GND efet w=9425 l=8700
+ ad=0 pd=0 as=7.77925e+08 ps=165300 
M3223 TMP_3 N0937 N0893 GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3224 TMP_3 N0946 Vdd GND efet w=13775 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3225 Vdd N0914 N0861 GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3226 Vdd Vdd S00817 GND efet w=6525 l=9425
+ ad=0 pd=0 as=-1.95488e+09 ps=316100 
M3227 GND N0945 TMP_3 GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3228 D3 N0964 N0607 GND efet w=14500 l=14500
+ ad=0 pd=0 as=0 ps=0 
M3229 N0945 S00817 N0945 GND efet w=68150 l=5800
+ ad=1.14376e+09 pd=226200 as=0 ps=0 
M3230 GND N0607 N0945 GND efet w=38425 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3231 d0 GND GND GND efet w=116000 l=13050
+ ad=-1.7993e+09 pd=513300 as=0 ps=0 
M3232 N0854 S00828 N0854 GND efet w=57275 l=17400
+ ad=0 pd=0 as=0 ps=0 
M3233 GND N0403 N0357 GND efet w=60175 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3234 Vdd Vdd S00819 GND efet w=7250 l=9425
+ ad=0 pd=0 as=-1.76986e+09 ps=356700 
M3235 N0945 S00817 Vdd GND efet w=5800 l=40600
+ ad=0 pd=0 as=0 ps=0 
M3236 N0937 S00819 N0937 GND efet w=66700 l=5800
+ ad=0 pd=0 as=0 ps=0 
M3237 N0670 d0 GND GND efet w=71775 l=12325
+ ad=1.18581e+09 pd=237800 as=0 ps=0 
M3238 GND N0670 D0 GND efet w=49300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3239 GND N0670 N0669 GND efet w=13775 l=11600
+ ad=0 pd=0 as=1.50329e+09 ps=310300 
M3240 d1 GND GND GND efet w=114550 l=14500
+ ad=-1.52808e+09 pd=516200 as=0 ps=0 
M3241 N0854 S00828 Vdd GND efet w=7250 l=52200
+ ad=0 pd=0 as=0 ps=0 
M3242 Vdd Vdd S00828 GND efet w=8700 l=13050
+ ad=0 pd=0 as=-1.7152e+09 ps=316100 
M3243 N0670 N0676 GND GND efet w=51475 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3244 GND N0676 N0669 GND efet w=25375 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3245 D0 N0669 Vdd GND efet w=38425 l=13050
+ ad=0 pd=0 as=0 ps=0 
M3246 N0670 Vdd Vdd GND efet w=10150 l=36975
+ ad=0 pd=0 as=0 ps=0 
M3247 N0669 Vdd Vdd GND efet w=5800 l=50750
+ ad=0 pd=0 as=0 ps=0 
M3248 GND D0 N0674 GND efet w=57275 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3249 N0674 Vdd Vdd GND efet w=13050 l=39150
+ ad=0 pd=0 as=0 ps=0 
M3250 N0674 N0702 N0697 GND efet w=27550 l=11600
+ ad=0 pd=0 as=-1.79509e+09 ps=481400 
M3251 GND N0697 N0696 GND efet w=99325 l=10875
+ ad=0 pd=0 as=5.11788e+08 ps=1.7893e+06 
M3252 d0 N0696 Vdd GND efet w=666275 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3253 N0733 N0713 GND GND efet w=55100 l=14500
+ ad=-6.68155e+08 pd=658300 as=0 ps=0 
M3254 Vdd N0713 cm_ram1 GND efet w=142100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3255 Vdd N0716 cm_ram0 GND efet w=142100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3256 Vdd Vdd N0733 GND efet w=7250 l=23200
+ ad=0 pd=0 as=0 ps=0 
M3257 Vdd Vdd N0736 GND efet w=8700 l=21750
+ ad=0 pd=0 as=-6.87077e+08 ps=652500 
M3258 GND N0716 N0736 GND efet w=43500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3259 cm_ram1 N0733 GND GND efet w=261725 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3260 cm_ram0 N0736 GND GND efet w=256650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3261 GND N0698 d0 GND efet w=1218725 l=6525
+ ad=0 pd=0 as=0 ps=0 
M3262 N0696 N0700 GND GND efet w=247950 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3263 Vdd Vdd S00835 GND efet w=9425 l=12325
+ ad=0 pd=0 as=-1.97801e+09 ps=275500 
M3264 Vdd S00835 N0696 GND efet w=10875 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3265 N0696 S00835 N0696 GND efet w=78300 l=5800
+ ad=0 pd=0 as=0 ps=0 
M3266 GND N0696 N0698 GND efet w=81925 l=12325
+ ad=0 pd=0 as=-5.54469e+07 ps=2.4824e+06 
M3267 N0698 N0700 GND GND efet w=229100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3268 Vdd S00839 N0698 GND efet w=10150 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3269 N0698 S00839 N0698 GND efet w=58000 l=34800
+ ad=0 pd=0 as=0 ps=0 
M3270 Vdd Vdd S00839 GND efet w=10150 l=13050
+ ad=0 pd=0 as=-2.05791e+09 ps=261000 
M3271 N0668 d1 GND GND efet w=66700 l=13050
+ ad=1.20473e+09 pd=243600 as=0 ps=0 
M3272 N0937 S00819 Vdd GND efet w=6525 l=33350
+ ad=0 pd=0 as=0 ps=0 
M3273 GND GND d2 GND efet w=99325 l=15225
+ ad=0 pd=0 as=0 ps=0 
M3274 GND N0668 D1 GND efet w=49300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3275 N0667 N0668 GND GND efet w=16675 l=10875
+ ad=1.07858e+09 pd=223300 as=0 ps=0 
M3276 GND N0676 N0667 GND efet w=26825 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3277 N0668 N0676 GND GND efet w=44225 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3278 Vdd Vdd N0667 GND efet w=6525 l=55825
+ ad=0 pd=0 as=0 ps=0 
M3279 D1 N0667 Vdd GND efet w=39150 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3280 N0668 Vdd Vdd GND efet w=8700 l=35525
+ ad=0 pd=0 as=0 ps=0 
M3281 GND D1 N0673 GND efet w=50750 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3282 N0673 N0702 N0694 GND efet w=27550 l=12325
+ ad=0 pd=0 as=-1.84766e+09 ps=478500 
M3283 N0673 Vdd Vdd GND efet w=10875 l=36975
+ ad=0 pd=0 as=0 ps=0 
M3284 D3 N0664 GND GND efet w=49300 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3285 Vdd N0663 D3 GND efet w=39875 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3286 GND POC d3 GND efet w=29000 l=14500
+ ad=0 pd=0 as=0 ps=0 
M3287 Vdd N0693 d1 GND efet w=681500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3288 d0 POC GND GND efet w=33350 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3289 GND N0694 N0693 GND efet w=99325 l=10875
+ ad=0 pd=0 as=1.23715e+09 ps=1.8357e+06 
M3290 N0693 N0700 GND GND efet w=257375 l=19575
+ ad=0 pd=0 as=0 ps=0 
M3291 Vdd Vdd S00836 GND efet w=7250 l=11600
+ ad=0 pd=0 as=2.14455e+09 ps=263900 
M3292 Vdd S00836 N0693 GND efet w=9425 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3293 GND N0695 d1 GND efet w=1217275 l=6525
+ ad=0 pd=0 as=0 ps=0 
M3294 N0693 S00836 N0693 GND efet w=75400 l=7250
+ ad=0 pd=0 as=0 ps=0 
M3295 Vdd Vdd N0663 GND efet w=9425 l=49300
+ ad=0 pd=0 as=-2.37142e+08 ps=791700 
M3296 Vdd Vdd N0664 GND efet w=8700 l=36250
+ ad=0 pd=0 as=3.19777e+07 ps=800400 
M3297 GND N0676 N0664 GND efet w=56550 l=14500
+ ad=0 pd=0 as=0 ps=0 
M3298 GND N0693 N0695 GND efet w=75400 l=13050
+ ad=0 pd=0 as=5.22741e+08 ps=2.494e+06 
M3299 N0695 N0700 GND GND efet w=229825 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3300 Vdd S00840 N0695 GND efet w=10150 l=14500
+ ad=0 pd=0 as=0 ps=0 
M3301 N0695 S00840 N0695 GND efet w=56550 l=37700
+ ad=0 pd=0 as=0 ps=0 
M3302 Vdd Vdd S00840 GND efet w=7250 l=13775
+ ad=0 pd=0 as=2.11932e+09 ps=261000 
M3303 GND N0664 N0663 GND efet w=23200 l=15950
+ ad=0 pd=0 as=0 ps=0 
M3304 N0663 N0676 GND GND efet w=23925 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3305 GND d3 N0664 GND efet w=86275 l=15225
+ ad=0 pd=0 as=0 ps=0 
M3306 d3 GND GND GND efet w=124700 l=13050
+ ad=0 pd=0 as=0 ps=0 
M3307 d1 POC GND GND efet w=30450 l=10875
+ ad=0 pd=0 as=0 ps=0 
C0 S00042 gnd! 33.7fF ;**FLOATING
C1 S00040 gnd! 73.8fF ;**FLOATING
C2 S00034 gnd! 29.1fF ;**FLOATING
C3 S00033 gnd! 4.4fF ;**FLOATING
C4 S00022 gnd! 7.6fF ;**FLOATING
C5 S00021 gnd! 26.0fF ;**FLOATING
C6 S00020 gnd! 62.4fF ;**FLOATING
C7 S00017 gnd! 17.9fF ;**FLOATING
C8 S00016 gnd! 13.8fF ;**FLOATING
C9 S00026 gnd! 31.4fF ;**FLOATING
C10 S00018 gnd! 30.1fF ;**FLOATING
C11 S00011 gnd! 195.8fF ;**FLOATING
C12 S00010 gnd! 221.7fF ;**FLOATING
C13 S00009 gnd! 54.9fF ;**FLOATING
C14 S00008 gnd! 55.7fF ;**FLOATING
C15 S00007 gnd! 55.5fF ;**FLOATING
C16 S00006 gnd! 55.5fF ;**FLOATING
C17 S00840 gnd! 115.8fF
C18 N0695 gnd! 1031.5fF
C19 S00836 gnd! 118.8fF
C20 N0693 gnd! 883.0fF
C21 N0694 gnd! 139.2fF
C22 N0673 gnd! 93.1fF
C23 N0667 gnd! 130.9fF
C24 N0663 gnd! 285.7fF
C25 N0664 gnd! 410.6fF
C26 N0668 gnd! 225.1fF
C27 S00839 gnd! 122.2fF
C28 S00835 gnd! 129.5fF
C29 N0698 gnd! 1030.5fF
C30 cm_ram0 gnd! 677.7fF
C31 cm_ram1 gnd! 548.8fF
C32 N0736 gnd! 255.5fF
C33 N0733 gnd! 239.8fF
C34 N0696 gnd! 886.8fF
C35 N0697 gnd! 164.7fF
C36 N0674 gnd! 86.4fF
C37 N0669 gnd! 162.8fF
C38 N0670 gnd! 244.9fF
C39 S00819 gnd! 135.1fF
C40 S00828 gnd! 148.5fF
C41 d1 gnd! 2381.2fF
C42 d0 gnd! 2381.0fF
C43 S00817 gnd! 124.4fF
C44 N0607 gnd! 76.7fF
C45 TMP_3 gnd! 104.1fF
C46 N0918 gnd! 50.4fF
C47 N0945 gnd! 180.4fF
C48 _TMP_3 gnd! 114.5fF
C49 N0946 gnd! 81.7fF
C50 N0914 gnd! 269.7fF
C51 N0901 gnd! 116.2fF
C52 N0558 gnd! 175.7fF
C53 N0893 gnd! 379.8fF
C54 N0557 gnd! 104.3fF
C55 N0892 gnd! 65.4fF
C56 N0897 gnd! 51.7fF
C57 N0859 gnd! 431.5fF
C58 S00834 gnd! 103.9fF
C59 N0713 gnd! 451.9fF
C60 S00833 gnd! 126.2fF
C61 N0357 gnd! 532.5fF
C62 N0359 gnd! 367.5fF
C63 cm_ram2 gnd! 343.4fF
C64 cm_ram3 gnd! 445.2fF
C65 N0852 gnd! 112.3fF
C66 N0735 gnd! 254.2fF
C67 N0734 gnd! 240.3fF
C68 S00825 gnd! 129.3fF
C69 N0366 gnd! 398.9fF
C70 N0715 gnd! 532.8fF
C71 N0730 gnd! 62.2fF
C72 N0287 gnd! 44.9fF
C73 S00818 gnd! 129.1fF
C74 N0714 gnd! 594.1fF
C75 N0358 gnd! 441.3fF
C76 ACC_3 gnd! 196.5fF
C77 N0873 gnd! 464.2fF
C78 N0877 gnd! 218.6fF
C79 N0474 gnd! 267.2fF
C80 S00814 gnd! 122.7fF
C81 N0731 gnd! 120.2fF
C82 N0748 gnd! 173.3fF
C83 N0749 gnd! 161.3fF
C84 N0349 gnd! 164.6fF
C85 N0666 gnd! 224.5fF
C86 S00801 gnd! 133.1fF
C87 S00804 gnd! 128.9fF
C88 TMP_2 gnd! 112.2fF
C89 N0917 gnd! 53.8fF
C90 N0665 gnd! 159.5fF
C91 N0943 gnd! 157.6fF
C92 _TMP_2 gnd! 110.6fF
C93 N0944 gnd! 82.7fF
C94 N0606 gnd! 157.1fF
C95 N0913 gnd! 231.5fF
C96 N0885 gnd! 86.1fF
C97 S00803 gnd! 127.0fF
C98 N0728 gnd! 66.2fF
C99 DCL_2 gnd! 180.3fF
C100 N0286 gnd! 46.7fF
C101 N0559 gnd! 126.7fF
C102 N0900 gnd! 116.6fF
C103 N0555 gnd! 182.2fF
C104 N0514 gnd! 923.0fF
C105 N0891 gnd! 411.5fF
C106 N0554 gnd! 130.5fF
C107 N0890 gnd! 64.3fF
C108 N0896 gnd! 51.5fF
C109 N0473 gnd! 292.0fF
C110 N0768 gnd! 206.7fF
C111 N0355 gnd! 175.3fF
C112 S00800 gnd! 118.6fF
C113 N0750 gnd! 223.5fF
C114 ACC_2 gnd! 202.4fF
C115 N0872 gnd! 535.3fF
C116 N0729 gnd! 119.4fF
C117 N0747 gnd! 174.5fF
C118 N0858 gnd! 351.6fF
C119 N0876 gnd! 61.6fF
C120 N0851 gnd! 90.2fF
C121 S00781 gnd! 143.3fF
C122 N0605 gnd! 84.6fF
C123 N0691 gnd! 176.5fF
C124 N0692 gnd! 1069.5fF
C125 N0916 gnd! 50.8fF
C126 N0690 gnd! 967.5fF
C127 S00766 gnd! 121.2fF
C128 S00765 gnd! 131.6fF
C129 N0672 gnd! 113.1fF
C130 N0941 gnd! 166.0fF
C131 _TMP_1 gnd! 153.5fF
C132 TMP_1 gnd! 114.0fF
C133 N0364 gnd! 193.9fF
C134 N0765 gnd! 163.9fF
C135 N0879 gnd! 207.0fF
C136 N0850 gnd! 97.8fF
C137 N0848 gnd! 1097.4fF
C138 N0556 gnd! 340.0fF
C139 N0899 gnd! 115.7fF
C140 N0942 gnd! 80.8fF
C141 d2 gnd! 2347.4fF
C142 S00767 gnd! 140.4fF
C143 DCL_1 gnd! 197.8fF
C144 N0726 gnd! 69.0fF
C145 N0552 gnd! 169.2fF
C146 N0857 gnd! 391.7fF
C147 ACC_1 gnd! 196.7fF
C148 N0889 gnd! 400.6fF
C149 N0551 gnd! 118.0fF
C150 N0888 gnd! 59.3fF
C151 N0895 gnd! 47.9fF
C152 N0912 gnd! 284.2fF
C153 N0871 gnd! 517.3fF
C154 N0472 gnd! 259.2fF
C155 N0875 gnd! 218.5fF
C156 N0371 gnd! 207.8fF
C157 N0285 gnd! 45.2fF
C158 N0716 gnd! 710.6fF
C159 N0767 gnd! 132.2fF
C160 S00764 gnd! 123.7fF
C161 N0884 gnd! 86.9fF
C162 S00762 gnd! 141.1fF
C163 N0964 gnd! 323.2fF
C164 N0604 gnd! 90.9fF
C165 TMP_0 gnd! 124.3fF
C166 N0915 gnd! 50.5fF
C167 N0911 gnd! 221.6fF
C168 N0471 gnd! 291.6fF
C169 N0847 gnd! 1017.6fF
C170 N0553 gnd! 346.3fF
C171 N0898 gnd! 104.7fF
C172 N0939 gnd! 168.6fF
C173 _TMP_0 gnd! 109.4fF
C174 N0940 gnd! 76.7fF
C175 N0549 gnd! 174.9fF
C176 N0887 gnd! 402.7fF
C177 ACC_0 gnd! 988.3fF
C178 N0376 gnd! 386.9fF
C179 N0370 gnd! 382.7fF
C180 N0363 gnd! 441.0fF
C181 N0354 gnd! 333.1fF
C182 N0345 gnd! 526.8fF
C183 N0377 gnd! 358.7fF
C184 N0751 gnd! 323.5fF
C185 N0766 gnd! 251.4fF
C186 N0347 gnd! 606.7fF
C187 N0348 gnd! 636.5fF
C188 S00778 gnd! 125.5fF
C189 N0727 gnd! 121.7fF
C190 N0746 gnd! 189.4fF
C191 DCL_0 gnd! 259.2fF
C192 N0819 gnd! 124.9fF
C193 N0356 gnd! 575.9fF
C194 N0350 gnd! 288.7fF
C195 N0378 gnd! 118.3fF
C196 N0818 gnd! 21.0fF
C197 N0724 gnd! 72.1fF
C198 N0284 gnd! 48.3fF
C199 N0346 gnd! 569.3fF
C200 N0849 gnd! 91.6fF
C201 N0856 gnd! 382.3fF
C202 N0878 gnd! 198.7fF
C203 N0870 gnd! 503.5fF
C204 N0548 gnd! 116.7fF
C205 N0886 gnd! 54.5fF
C206 N0874 gnd! 60.7fF
C207 N0894 gnd! 36.2fF
C208 N0452 gnd! 97.6fF
C209 N0937 gnd! 441.1fF
C210 N0704 gnd! 98.3fF
C211 N0706 gnd! 96.3fF
C212 N0705 gnd! 351.1fF
C213 N0707 gnd! 56.3fF
C214 N0684 gnd! 43.1fF
C215 N0676 gnd! 1685.7fF
C216 N0685 gnd! 175.9fF
C217 N0677 gnd! 78.3fF
C218 N0699 gnd! 57.8fF
C219 N0846 gnd! 1078.2fF
C220 N0861 gnd! 248.0fF
C221 S00734 gnd! 168.9fF
C222 N0855 gnd! 417.7fF
C223 N0550 gnd! 251.6fF
C224 N0470 gnd! 297.5fF
C225 ADC_CY gnd! 347.9fF
C226 S00732 gnd! 139.6fF
C227 CY gnd! 262.0fF
C228 N0860 gnd! 36.8fF
C229 N0513 gnd! 400.6fF
C230 ACC_ADA gnd! 598.9fF
C231 CY_ADAC gnd! 238.4fF
C232 N0686 gnd! 35.5fF
C233 CY_ADA gnd! 235.6fF
C234 ADD_ACC gnd! 571.8fF
C235 N0546 gnd! 127.3fF
C236 N0701 gnd! 150.1fF
C237 N0678 gnd! 181.6fF
C238 N0675 gnd! 224.1fF
C239 S00716 gnd! 132.4fF
C240 d3 gnd! 2687.2fF
C241 N0658 gnd! 119.4fF
C242 N0659 gnd! 291.4fF
C243 N0689 gnd! 1074.4fF
C244 N0700 gnd! 1750.5fF
C245 S00689 gnd! 119.4fF
C246 N0687 gnd! 913.4fF
C247 S00687 gnd! 112.7fF
C248 N1015 gnd! 63.6fF
C249 N1013 gnd! 160.3fF
C250 N1014 gnd! 188.6fF
C251 N0688 gnd! 260.4fF
C252 N0671 gnd! 147.2fF
C253 N1006 gnd! 233.2fF
C254 N1007 gnd! 266.6fF
C255 S00676 gnd! 119.3fF
C256 N0702 gnd! 1096.7fF
C257 N1012 gnd! 227.3fF
C258 ACC_ADAC gnd! 550.7fF
C259 N0854 gnd! 430.0fF
C260 N0515 gnd! 49.8fF
C261 ADSR gnd! 490.9fF
C262 N0490 gnd! 84.0fF
C263 S00724 gnd! 151.4fF
C264 S00729 gnd! 136.5fF
C265 ADSL gnd! 603.7fF
C266 CY_IB gnd! 238.6fF
C267 N0502 gnd! 71.2fF
C268 S00709 gnd! 138.8fF
C269 SUB_GROUP_6_ gnd! 1134.8fF
C270 ADD_IB gnd! 696.1fF
C271 ACB_IB gnd! 851.3fF
C272 N0445 gnd! 90.8fF
C273 INC_GROUP_5_ gnd! 391.7fF
C274 N0448 gnd! 215.5fF
C275 S00761 gnd! 126.0fF
C276 S00757 gnd! 107.6fF
C277 N0725 gnd! 121.7fF
C278 N0745 gnd! 218.8fF
C279 N0803 gnd! 154.9fF
C280 N0403 gnd! 739.5fF
C281 N0802 gnd! 99.7fF
C282 N0425 gnd! 40.2fF
C283 N0421 gnd! 77.8fF
C284 N0422 gnd! 41.8fF
C285 N0853 gnd! 238.6fF
C286 S00731 gnd! 173.2fF
C287 N0433 gnd! 47.2fF
C288 N0722 gnd! 67.9fF
C289 N0283 gnd! 46.1fF
C290 N0431 gnd! 84.7fF
C291 N0430 gnd! 63.1fF
C292 N0340 gnd! 113.9fF
C293 S00740 gnd! 121.4fF
C294 N0723 gnd! 121.4fF
C295 N0744 gnd! 182.5fF
C296 N0423 gnd! 237.3fF
C297 N0342 gnd! 1079.7fF
C298 N0446 gnd! 213.1fF
C299 READ_ACC_3_ gnd! 543.5fF
C300 ADD_GROUP_4_ gnd! 433.0fF
C301 N0442 gnd! 172.0fF
C302 WRITE_CARRY_2_ gnd! 663.0fF
C303 N0336 gnd! 24.6fF
C304 N0335 gnd! 23.3fF
C305 N0332 gnd! 263.1fF
C306 N0330 gnd! 21.0fF
C307 N0331 gnd! 112.3fF
C308 N0328 gnd! 137.8fF
C309 N0369 gnd! 48.6fF
C310 N0720 gnd! 69.6fF
C311 N0282 gnd! 49.8fF
C312 N0360 gnd! 61.0fF
C313 N0337 gnd! 175.6fF
C314 WRITE_ACC_1_ gnd! 702.0fF
C315 N0351 gnd! 922.3fF
C316 N0353 gnd! 61.4fF
C317 __X21__CLK2_ gnd! 950.6fF
C318 N1004 gnd! 217.6fF
C319 N0512 gnd! 52.6fF
C320 S00725 gnd! 119.2fF
C321 N0721 gnd! 120.2fF
C322 N0743 gnd! 207.7fF
C323 N0380 gnd! 48.7fF
C324 S00699 gnd! 132.9fF
C325 N0383 gnd! 26.1fF
C326 N0718 gnd! 70.0fF
C327 N0281 gnd! 48.3fF
C328 S00710 gnd! 116.0fF
C329 N0288 gnd! 573.3fF
C330 N0719 gnd! 117.2fF
C331 N0742 gnd! 190.3fF
C332 N0375 gnd! 156.4fF
C333 N0800 gnd! 20.0fF
C334 _COM gnd! 1060.5fF
C335 N0805 gnd! 516.1fF
C336 N0801 gnd! 394.9fF
C337 N0798 gnd! 53.8fF
C338 N0797 gnd! 96.2fF
C339 OPA_1 gnd! 986.3fF
C340 N0507 gnd! 46.3fF
C341 N0415 gnd! 655.1fF
C342 N0408 gnd! 45.8fF
C343 N0407 gnd! 47.7fF
C344 N0414 gnd! 41.6fF
C345 N0782 gnd! 274.2fF
C346 S00690 gnd! 120.4fF
C347 N0784 gnd! 64.9fF
C348 N0799 gnd! 73.2fF
C349 N0398 gnd! 116.1fF
C350 S00685 gnd! 156.7fF
C351 _OPA_1 gnd! 630.5fF
C352 CY_1 gnd! 1198.5fF
C353 N1005 gnd! 318.1fF
C354 N1002 gnd! 276.6fF
C355 N0501 gnd! 56.6fF
C356 _OPA_2 gnd! 767.8fF
C357 N1000 gnd! 278.6fF
C358 N1001 gnd! 324.8fF
C359 N1003 gnd! 344.8fF
C360 N0483 gnd! 33.2fF
C361 OPA_2 gnd! 752.4fF
C362 N0486 gnd! 207.9fF
C363 N0481 gnd! 106.2fF
C364 ADD_0 gnd! 813.2fF
C365 _OPA_3 gnd! 771.3fF
C366 N0487 gnd! 119.0fF
C367 N0478 gnd! 216.8fF
C368 N0329 gnd! 442.0fF
C369 N0741 gnd! 184.5fF
C370 N0432 gnd! 386.4fF
C371 N0456 gnd! 100.7fF
C372 N0404 gnd! 38.7fF
C373 N0739 gnd! 116.9fF
C374 N0296 gnd! 104.7fF
C375 N0280 gnd! 77.7fF
C376 S00678 gnd! 115.1fF
C377 N0297 gnd! 173.7fF
C378 N0405 gnd! 52.0fF
C379 N0413 gnd! 93.5fF
C380 N0419 gnd! 152.9fF
C381 N0482 gnd! 18.5fF
C382 N0479 gnd! 58.7fF
C383 N0480 gnd! 67.9fF
C384 N0477 gnd! 416.5fF
C385 __X31__CLK2_ gnd! 998.0fF
C386 ADM gnd! 278.0fF
C387 SBM gnd! 298.2fF
C388 CLB gnd! 252.3fF
C389 CLC gnd! 228.2fF
C390 OPA_3 gnd! 818.3fF
C391 OPA_IB gnd! 671.1fF
C392 N0997 gnd! 290.5fF
C393 IAC gnd! 276.7fF
C394 DAC gnd! 252.8fF
C395 CMC gnd! 312.2fF
C396 CMA gnd! 350.7fF
C397 RAL gnd! 365.2fF
C398 RAR gnd! 351.2fF
C399 IOW gnd! 302.0fF
C400 TCC gnd! 279.9fF
C401 STC gnd! 269.5fF
C402 DAA gnd! 765.5fF
C403 TCS gnd! 949.4fF
C404 KBP gnd! 688.9fF
C405 DCL gnd! 221.2fF
C406 O_IB gnd! 592.9fF
C407 N0418 gnd! 26.5fF
C408 N0399 gnd! 50.6fF
C409 N0476 gnd! 75.4fF
C410 _I_O gnd! 871.9fF
C411 _OPE gnd! 622.0fF
C412 N0412 gnd! 25.2fF
C413 N0417 gnd! 27.1fF
C414 N0397 gnd! 100.6fF
C415 N0327 gnd! 217.7fF
C416 _SRC gnd! 253.2fF
C417 N0516 gnd! 26.5fF
C418 N0510 gnd! 75.9fF
C419 N0493 gnd! 52.1fF
C420 N0769 gnd! 66.5fF
C421 OPR_0 gnd! 472.4fF
C422 OPA_0 gnd! 1180.5fF
C423 N0367 gnd! 15.8fF
C424 _OPR_0 gnd! 749.1fF
C425 N0352 gnd! 80.4fF
C426 N0999 gnd! 424.4fF
C427 N0996 gnd! 380.4fF
C428 N1008 gnd! 95.0fF
C429 N0998 gnd! 304.2fF
C430 N1010 gnd! 159.1fF
C431 N1009 gnd! 200.5fF
C432 N1011 gnd! 228.9fF
C433 SC_M12_CLK2 gnd! 150.6fF
C434 N0992 gnd! 263.8fF
C435 N0993 gnd! 309.4fF
C436 N0368 gnd! 164.6fF
C437 OPR_1 gnd! 756.7fF
C438 N0994 gnd! 243.2fF
C439 N0995 gnd! 482.1fF
C440 _OPR_1 gnd! 892.6fF
C441 OPR_2 gnd! 876.2fF
C442 JUN2_JMS2 gnd! 470.1fF
C443 N0362 gnd! 43.7fF
C444 N0361 gnd! 62.9fF
C445 N0372 gnd! 137.9fF
C446 N0373 gnd! 153.3fF
C447 N0523 gnd! 243.9fF
C448 N0660 gnd! 79.5fF
C449 N0644 gnd! 16.8fF
C450 N0661 gnd! 25.9fF
C451 N0662 gnd! 30.3fF
C452 L gnd! 942.2fF
C453 N0631 gnd! 23.1fF
C454 N0629 gnd! 100.4fF
C455 JCN gnd! 319.7fF
C456 _OPR_2 gnd! 851.2fF
C457 ISZ gnd! 326.7fF
C458 FIN_FIM gnd! 253.0fF
C459 N0587 gnd! 338.7fF
C460 FIM_SRC gnd! 251.5fF
C461 N0343 gnd! 163.8fF
C462 OPR_3 gnd! 880.1fF
C463 LDM_BBL gnd! 547.6fF
C464 ADD gnd! 458.5fF
C465 SUB gnd! 485.2fF
C466 LD gnd! 477.0fF
C467 XCH gnd! 572.5fF
C468 IOR gnd! 763.8fF
C469 N0681 gnd! 22.1fF
C470 N0703 gnd! 143.0fF
C471 N0643 gnd! 113.3fF
C472 N0680 gnd! 28.0fF
C473 N0679 gnd! 84.8fF
C474 N0630 gnd! 118.6fF
C475 N0623 gnd! 38.9fF
C476 N0682 gnd! 241.4fF
C477 N0683 gnd! 252.6fF
C478 N0618 gnd! 180.9fF
C479 N0654 gnd! 62.7fF
C480 N0651 gnd! 17.7fF
C481 N0650 gnd! 43.5fF
C482 N0579 gnd! 17.7fF
C483 N0567 gnd! 25.2fF
C484 N0628 gnd! 284.6fF
C485 INC_ISZ gnd! 602.2fF
C486 N0575 gnd! 67.3fF
C487 N0576 gnd! 17.7fF
C488 N0563 gnd! 18.1fF
C489 INC_ISZ_XCH gnd! 388.4fF
C490 N0568 gnd! 203.9fF
C491 _OPR_3 gnd! 821.3fF
C492 OPE gnd! 322.3fF
C493 IO gnd! 306.4fF
C494 N0603 gnd! 73.3fF
C495 N0590 gnd! 111.4fF
C496 N0611 gnd! 71.5fF
C497 N0596 gnd! 72.1fF
C498 N0562 gnd! 60.6fF
C499 N0656 gnd! 51.5fF
C500 N0564 gnd! 223.7fF
C501 N0597 gnd! 22.1fF
C502 N0612 gnd! 62.4fF
C503 N0636 gnd! 409.6fF
C504 N0614 gnd! 37.2fF
C505 N0640 gnd! 35.5fF
C506 _OPA_0 gnd! 1766.9fF
C507 N0639 gnd! 72.1fF
C508 N0602 gnd! 131.8fF
C509 N0627 gnd! 68.4fF
C510 S00627 gnd! 148.5fF
C511 S00620 gnd! 147.3fF
C512 N0621 gnd! 113.5fF
C513 N0622 gnd! 233.4fF
C514 N0626 gnd! 395.6fF
C515 N0652 gnd! 24.4fF
C516 N0547 gnd! 201.8fF
C517 N0595 gnd! 17.7fF
C518 N0527 gnd! 21.0fF
C519 N0468 gnd! 116.9fF
C520 BBL gnd! 290.3fF
C521 N0589 gnd! 15.6fF
C522 N0594 gnd! 21.9fF
C523 FIN_FIM_SRC_JIN gnd! 745.7fF
C524 INC_ISZ_ADD_SUB_XCH_LD gnd! 720.9fF
C525 N0580 gnd! 414.3fF
C526 N0608 gnd! 96.3fF
C527 N0615 gnd! 101.6fF
C528 S00624 gnd! 138.2fF
C529 N0578 gnd! 251.7fF
C530 N0649 gnd! 160.5fF
C531 N0655 gnd! 166.4fF
C532 N0653 gnd! 76.1fF
C533 N0641 gnd! 39.5fF
C534 N0642 gnd! 219.8fF
C535 N0638 gnd! 27.5fF
C536 N0633 gnd! 63.1fF
C537 N0637 gnd! 234.6fF
C538 REG_RFSH_2 gnd! 102.6fF
C539 N0624 gnd! 24.2fF
C540 N0588 gnd! 99.0fF
C541 N0460 gnd! 80.4fF
C542 N0484 gnd! 21.9fF
C543 N0485 gnd! 22.1fF
C544 JMS gnd! 336.9fF
C545 N0525 gnd! 15.8fF
C546 N0526 gnd! 156.4fF
C547 N0528 gnd! 93.0fF
C548 N0429 gnd! 15.8fF
C549 N0428 gnd! 84.1fF
C550 N0495 gnd! 21.4fF
C551 N0524 gnd! 319.7fF
C552 N0496 gnd! 29.6fF
C553 N0601 gnd! 24.6fF
C554 N0585 gnd! 24.4fF
C555 N0625 gnd! 74.3fF
C556 N0609 gnd! 39.9fF
C557 N0467 gnd! 245.6fF
C558 DC gnd! 902.4fF
C559 N0592 gnd! 108.8fF
C560 N0509 gnd! 22.5fF
C561 N0506 gnd! 58.0fF
C562 N0494 gnd! 110.3fF
C563 N0520 gnd! 22.5fF
C564 CLK2_JMS_DC_M22_BBL_M22_X12_X22__ gnd! 254.7fF
C565 N0593 gnd! 67.5fF
C566 N0586 gnd! 70.6fF
C567 N0572 gnd! 24.0fF
C568 N0610 gnd! 367.8fF
C569 N0600 gnd! 456.2fF
C570 N0573 gnd! 38.5fF
C571 SC_A12_CLK2 gnd! 283.5fF
C572 N0566 gnd! 65.8fF
C573 N0571 gnd! 452.7fF
C574 N0521 gnd! 49.1fF
C575 N0505 gnd! 51.7fF
C576 N0511 gnd! 139.2fF
C577 _INH gnd! 341.6fF
C578 N0344 gnd! 131.4fF
C579 S00654 gnd! 115.0fF
C580 N0338 gnd! 24.2fF
C581 N0339 gnd! 190.9fF
C582 N0341 gnd! 28.8fF
C583 N0334 gnd! 25.4fF
C584 N0333 gnd! 26.5fF
C585 _CN gnd! 598.4fF
C586 N0438 gnd! 83.2fF
C587 N0441 gnd! 35.3fF
C588 N0447 gnd! 129.8fF
C589 POC gnd! 4638.9fF
C590 N0451 gnd! 55.3fF
C591 N0435 gnd! 170.3fF
C592 N0443 gnd! 88.4fF
C593 N0522 gnd! 134.8fF
C594 N0517 gnd! 81.5fF
C595 S00628 gnd! 110.1fF
C596 N0437 gnd! 51.1fF
C597 N0436 gnd! 257.8fF
C598 INH gnd! 401.6fF
C599 N0321 gnd! 22.1fF
C600 N0324 gnd! 21.0fF
C601 N0319 gnd! 21.9fF
C602 N0320 gnd! 25.9fF
C603 JCN_ISZ gnd! 818.8fF
C604 N0322 gnd! 333.0fF
C605 JIN_FIN gnd! 893.9fF
C606 SC gnd! 2123.3fF
C607 N0323 gnd! 67.3fF
C608 N0309 gnd! 22.1fF
C609 N0308 gnd! 48.6fF
C610 N0450 gnd! 71.1fF
C611 JUN_JMS gnd! 926.0fF
C612 N0310 gnd! 242.7fF
C613 X22 gnd! 1737.1fF
C614 S00612 gnd! 122.4fF
C615 S00613 gnd! 136.7fF
C616 N0449 gnd! 292.1fF
C617 ADDR_PTR_0 gnd! 203.3fF
C618 REG_RFSH_1 gnd! 108.1fF
C619 N0574 gnd! 244.8fF
C620 REG_RFSH_0 gnd! 102.6fF
C621 SC_A22 gnd! 658.2fF
C622 SC_M22_CLK2 gnd! 806.3fF
C623 S00585 gnd! 169.7fF
C624 S00584 gnd! 170.1fF
C625 S00583 gnd! 172.8fF
C626 S00582 gnd! 171.6fF
C627 S00581 gnd! 171.1fF
C628 S00580 gnd! 170.5fF
C629 N0582 gnd! 449.5fF
C630 N0465 gnd! 22.5fF
C631 S00601 gnd! 165.6fF
C632 N0466 gnd! 231.0fF
C633 N0491 gnd! 23.1fF
C634 S00600 gnd! 164.5fF
C635 S00599 gnd! 166.1fF
C636 X12 gnd! 2666.8fF
C637 S00598 gnd! 171.9fF
C638 N0420 gnd! 202.1fF
C639 N0458 gnd! 60.4fF
C640 N0492 gnd! 50.5fF
C641 N0401 gnd! 193.2fF
C642 N0279 gnd! 80.3fF
C643 N0709 gnd! 32.6fF
C644 N0278 gnd! 68.3fF
C645 M22 gnd! 2059.7fF
C646 M12 gnd! 4535.7fF
C647 N0365 gnd! 221.2fF
C648 N0379 gnd! 162.4fF
C649 N0459 gnd! 318.6fF
C650 N0457 gnd! 52.1fF
C651 ADDR_PTR_1 gnd! 209.4fF
C652 N0464 gnd! 182.2fF
C653 N0475 gnd! 192.1fF
C654 S00579 gnd! 170.4fF
C655 S00578 gnd! 173.5fF
C656 N0560 gnd! 359.6fF
C657 N0409 gnd! 230.7fF
C658 N0402 gnd! 145.3fF
C659 X32 gnd! 2478.4fF
C660 S00609 gnd! 123.0fF
C661 N0708 gnd! 171.4fF
C662 N0710 gnd! 110.6fF
C663 N0416 gnd! 49.1fF
C664 N0374 gnd! 50.7fF
C665 N0384 gnd! 48.8fF
C666 N0400 gnd! 247.5fF
C667 __FIN_X12_ gnd! 418.5fF
C668 N0508 gnd! 22.7fF
C669 N0617 gnd! 349.0fF
C670 N0561 gnd! 362.4fF
C671 N0504 gnd! 60.1fF
C672 __INH__X32_CLK2 gnd! 267.2fF
C673 N0518 gnd! 22.9fF
C674 N0440 gnd! 235.1fF
C675 N0427 gnd! 230.5fF
C676 N0519 gnd! 49.1fF
C677 N0542 gnd! 423.0fF
C678 N0577 gnd! 134.0fF
C679 N0541 gnd! 398.7fF
C680 N0646 gnd! 258.0fF
C681 N0833 gnd! 160.9fF
C682 ___SC__JIN_FIN__CLK1_M11_X21_INH_ gnd! 444.5fF
C683 N0732 gnd! 119.7fF
C684 __POC_CLK2_X12_X32__INH gnd! 393.8fF
C685 N0411 gnd! 235.2fF
C686 N0382 gnd! 249.4fF
C687 N0820 gnd! 107.1fF
C688 N0804 gnd! 116.1fF
C689 N0783 gnd! 139.7fF
C690 N0304 gnd! 432.7fF
C691 N0539 gnd! 187.1fF
C692 N0503 gnd! 52.4fF
C693 ADDR_RFSH_0 gnd! 284.3fF
C694 S00564 gnd! 131.0fF
C695 N0540 gnd! 160.0fF
C696 N0613 gnd! 354.5fF
C697 N0648 gnd! 312.9fF
C698 N0635 gnd! 301.3fF
C699 N0983 gnd! 130.5fF
C700 S00557 gnd! 133.5fF
C701 N0620 gnd! 289.2fF
C702 N0599 gnd! 292.4fF
C703 N0974 gnd! 129.5fF
C704 N0965 gnd! 130.6fF
C705 N0584 gnd! 280.9fF
C706 N0570 gnd! 284.1fF
C707 N0955 gnd! 128.5fF
C708 N0938 gnd! 126.0fF
C709 N0462 gnd! 22.9fF
C710 N0488 gnd! 22.5fF
C711 N0463 gnd! 253.5fF
C712 N0454 gnd! 69.0fF
C713 N0489 gnd! 56.0fF
C714 N0845 gnd! 17.5fF
C715 N0832 gnd! 17.2fF
C716 N0817 gnd! 18.5fF
C717 PC3_8 gnd! 36.7fF
C718 PC2_8 gnd! 36.6fF
C719 N0796 gnd! 16.8fF
C720 N0326 gnd! 652.1fF
C721 N0317 gnd! 56.9fF
C722 N0711 gnd! 123.2fF
C723 N0316 gnd! 55.3fF
C724 N0300 gnd! 349.0fF
C725 A12 gnd! 2975.7fF
C726 N0737 gnd! 489.7fF
C727 cm_rom gnd! 696.8fF
C728 A22 gnd! 2968.8fF
C729 N0712 gnd! 97.1fF
C730 N0315 gnd! 50.5fF
C731 A32 gnd! 2627.4fF
C732 N0318 gnd! 565.4fF
C733 PC1_8 gnd! 35.3fF
C734 PC0_8 gnd! 35.1fF
C735 N0844 gnd! 16.4fF
C736 PC3_4 gnd! 36.5fF
C737 N0455 gnd! 332.1fF
C738 CLK2_SC_A12_M12_ gnd! 950.3fF
C739 N0545 gnd! 277.9fF
C740 N0530 gnd! 209.3fF
C741 N0928 gnd! 125.6fF
C742 N0919 gnd! 126.3fF
C743 N0453 gnd! 53.2fF
C744 ADDR_RFSH_1 gnd! 323.5fF
C745 N0902 gnd! 132.2fF
C746 __POC__CLK2_SC_A32_X12_ gnd! 775.4fF
C747 N0991 gnd! 13.9fF
C748 N0982 gnd! 16.0fF
C749 N0973 gnd! 14.7fF
C750 R15_3 gnd! 41.1fF
C751 R13_3 gnd! 38.2fF
C752 N0963 gnd! 17.7fF
C753 N0954 gnd! 17.9fF
C754 R11_3 gnd! 37.4fF
C755 R9_3 gnd! 36.0fF
C756 N0990 gnd! 15.8fF
C757 R14_3 gnd! 38.6fF
C758 clk1 gnd! 5962.6fF
C759 N0989 gnd! 12.6fF
C760 N0981 gnd! 15.6fF
C761 N0972 gnd! 16.4fF
C762 N0936 gnd! 18.5fF
C763 N0927 gnd! 17.7fF
C764 N0461 gnd! 184.3fF
C765 N0469 gnd! 199.3fF
C766 R7_3 gnd! 35.6fF
C767 R5_3 gnd! 34.9fF
C768 R12_3 gnd! 38.1fF
C769 R10_3 gnd! 36.7fF
C770 R8_3 gnd! 36.4fF
C771 N0962 gnd! 15.3fF
C772 N0953 gnd! 16.8fF
C773 N0910 gnd! 16.2fF
C774 R3_3 gnd! 35.8fF
C775 R1_3 gnd! 36.0fF
C776 R6_3 gnd! 35.6fF
C777 N0980 gnd! 16.0fF
C778 N0971 gnd! 16.0fF
C779 R14_2 gnd! 38.5fF
C780 R12_2 gnd! 36.5fF
C781 N0961 gnd! 17.9fF
C782 N0952 gnd! 17.2fF
C783 N0935 gnd! 16.8fF
C784 N0926 gnd! 17.0fF
C785 R4_3 gnd! 38.4fF
C786 R10_2 gnd! 36.3fF
C787 R8_2 gnd! 35.7fF
C788 N0988 gnd! 13.7fF
C789 R15_2 gnd! 38.8fF
C790 clk2 gnd! 7223.1fF
C791 N0987 gnd! 12.6fF
C792 N0979 gnd! 17.9fF
C793 N0970 gnd! 15.3fF
C794 R13_2 gnd! 34.2fF
C795 R2_3 gnd! 34.5fF
C796 N0934 gnd! 17.9fF
C797 N0925 gnd! 16.6fF
C798 N0909 gnd! 16.2fF
C799 N0869 gnd! 494.8fF
C800 N0843 gnd! 17.0fF
C801 N0831 gnd! 16.2fF
C802 N0773 gnd! 350.3fF
C803 N0816 gnd! 16.4fF
C804 PC2_4 gnd! 37.0fF
C805 PC1_4 gnd! 35.6fF
C806 N0795 gnd! 16.8fF
C807 N0314 gnd! 57.2fF
C808 N0396 gnd! 310.4fF
C809 N0395 gnd! 365.1fF
C810 PC0_4 gnd! 35.2fF
C811 N0777 gnd! 348.6fF
C812 N0815 gnd! 17.9fF
C813 N0830 gnd! 17.5fF
C814 PC3_0 gnd! 36.5fF
C815 PC2_0 gnd! 35.5fF
C816 N0794 gnd! 18.1fF
C817 PC1_0 gnd! 34.8fF
C818 N0842 gnd! 17.2fF
C819 PC0_0 gnd! 36.0fF
C820 PC3_1 gnd! 35.7fF
C821 N0537 gnd! 421.5fF
C822 N0538 gnd! 452.0fF
C823 N0883 gnd! 466.5fF
C824 R0_3 gnd! 36.6fF
C825 R6_2 gnd! 36.0fF
C826 R4_2 gnd! 36.3fF
C827 R11_2 gnd! 36.4fF
C828 N0960 gnd! 16.8fF
C829 N0951 gnd! 16.2fF
C830 R9_2 gnd! 35.0fF
C831 N0908 gnd! 16.4fF
C832 R2_2 gnd! 36.2fF
C833 R0_2 gnd! 36.0fF
C834 R7_2 gnd! 35.3fF
C835 N0978 gnd! 17.9fF
C836 N0969 gnd! 13.7fF
C837 R15_1 gnd! 41.7fF
C838 R13_1 gnd! 35.7fF
C839 N0986 gnd! 13.2fF
C840 N0959 gnd! 18.3fF
C841 N0950 gnd! 15.1fF
C842 N0933 gnd! 16.6fF
C843 N0924 gnd! 16.6fF
C844 R5_2 gnd! 34.8fF
C845 N0882 gnd! 479.6fF
C846 R3_2 gnd! 36.8fF
C847 R11_1 gnd! 36.9fF
C848 R9_1 gnd! 34.4fF
C849 R14_1 gnd! 39.5fF
C850 N0932 gnd! 17.7fF
C851 N0907 gnd! 16.4fF
C852 R1_2 gnd! 34.7fF
C853 N0923 gnd! 16.2fF
C854 R7_1 gnd! 36.8fF
C855 R5_1 gnd! 34.9fF
C856 N0977 gnd! 17.5fF
C857 N0985 gnd! 12.4fF
C858 R12_1 gnd! 34.4fF
C859 N0968 gnd! 13.7fF
C860 R10_1 gnd! 37.8fF
C861 N0976 gnd! 17.7fF
C862 N0967 gnd! 12.8fF
C863 N0958 gnd! 17.5fF
C864 N0906 gnd! 16.6fF
C865 R3_1 gnd! 35.8fF
C866 R1_1 gnd! 36.1fF
C867 N0949 gnd! 16.6fF
C868 R8_1 gnd! 34.0fF
C869 R6_1 gnd! 36.2fF
C870 R14_0 gnd! 41.2fF
C871 R12_0 gnd! 37.3fF
C872 N0647 gnd! 331.2fF
C873 N0634 gnd! 323.7fF
C874 N0931 gnd! 17.0fF
C875 N0922 gnd! 16.8fF
C876 R4_1 gnd! 35.3fF
C877 N0957 gnd! 16.8fF
C878 N0948 gnd! 13.5fF
C879 R10_0 gnd! 39.6fF
C880 R8_0 gnd! 34.9fF
C881 N0619 gnd! 312.4fF
C882 N0598 gnd! 322.5fF
C883 N0984 gnd! 12.0fF
C884 R15_0 gnd! 39.3fF
C885 R13_0 gnd! 39.6fF
C886 N0975 gnd! 13.0fF
C887 N0966 gnd! 12.6fF
C888 N0657 gnd! 342.5fF
C889 R2_1 gnd! 35.2fF
C890 N0930 gnd! 16.8fF
C891 N0921 gnd! 16.4fF
C892 N0905 gnd! 16.4fF
C893 N0536 gnd! 424.2fF
C894 N0500 gnd! 107.0fF
C895 N0865 gnd! 218.7fF
C896 N0829 gnd! 18.9fF
C897 N0814 gnd! 19.1fF
C898 PC2_1 gnd! 34.6fF
C899 PC1_1 gnd! 34.7fF
C900 N0841 gnd! 16.8fF
C901 N0828 gnd! 18.7fF
C902 N0793 gnd! 16.2fF
C903 PC0_1 gnd! 35.6fF
C904 N0813 gnd! 20.4fF
C905 PC3_5 gnd! 37.1fF
C906 PC2_5 gnd! 35.8fF
C907 N0792 gnd! 18.1fF
C908 PC1_5 gnd! 32.9fF
C909 PC0_5 gnd! 35.4fF
C910 N0840 gnd! 17.9fF
C911 PC3_9 gnd! 36.4fF
C912 N0868 gnd! 493.1fF
C913 N0867 gnd! 491.2fF
C914 N0881 gnd! 468.6fF
C915 N0864 gnd! 232.2fF
C916 N0535 gnd! 454.1fF
C917 N0499 gnd! 110.0fF
C918 N0839 gnd! 18.1fF
C919 N0827 gnd! 18.3fF
C920 N0812 gnd! 19.6fF
C921 PC2_9 gnd! 35.7fF
C922 N0781 gnd! 351.3fF
C923 N0780 gnd! 349.7fF
C924 PC1_9 gnd! 32.8fF
C925 N0826 gnd! 20.0fF
C926 N0811 gnd! 18.3fF
C927 PC0_9 gnd! 36.0fF
C928 N0791 gnd! 16.0fF
C929 N0776 gnd! 353.6fF
C930 N0772 gnd! 343.3fF
C931 PC3_10 gnd! 35.8fF
C932 PC2_10 gnd! 34.1fF
C933 N0790 gnd! 17.5fF
C934 PC1_10 gnd! 35.2fF
C935 PC0_10 gnd! 36.8fF
C936 N0838 gnd! 17.7fF
C937 PC3_6 gnd! 35.2fF
C938 R0_1 gnd! 36.1fF
C939 R6_0 gnd! 37.7fF
C940 R4_0 gnd! 35.5fF
C941 N0904 gnd! 17.7fF
C942 R2_0 gnd! 37.3fF
C943 R0_0 gnd! 36.1fF
C944 N0583 gnd! 308.3fF
C945 N0569 gnd! 309.3fF
C946 N0544 gnd! 308.0fF
C947 N0529 gnd! 311.0fF
C948 R11_0 gnd! 40.5fF
C949 N0645 gnd! 330.8fF
C950 N0632 gnd! 328.6fF
C951 N0956 gnd! 13.7fF
C952 N0947 gnd! 13.0fF
C953 R9_0 gnd! 37.8fF
C954 R7_0 gnd! 39.8fF
C955 N0616 gnd! 318.2fF
C956 N0591 gnd! 327.3fF
C957 N0929 gnd! 16.8fF
C958 N0920 gnd! 13.5fF
C959 R5_0 gnd! 36.0fF
C960 N0581 gnd! 314.4fF
C961 R3_0 gnd! 39.2fF
C962 N0565 gnd! 318.7fF
C963 R1_0 gnd! 39.5fF
C964 N0903 gnd! 14.1fF
C965 N0880 gnd! 474.2fF
C966 WRAB0 gnd! 628.7fF
C967 N0533 gnd! 422.6fF
C968 N0837 gnd! 18.7fF
C969 N0825 gnd! 18.7fF
C970 N0810 gnd! 16.4fF
C971 PC2_6 gnd! 34.6fF
C972 PC1_6 gnd! 35.4fF
C973 N0534 gnd! 435.9fF
C974 N0498 gnd! 106.3fF
C975 N0824 gnd! 19.8fF
C976 N0809 gnd! 17.7fF
C977 PC0_6 gnd! 37.2fF
C978 N0789 gnd! 15.3fF
C979 N0771 gnd! 345.5fF
C980 PC3_2 gnd! 35.4fF
C981 PC2_2 gnd! 34.2fF
C982 N0863 gnd! 221.4fF
C983 N0788 gnd! 17.2fF
C984 PC1_2 gnd! 35.0fF
C985 PC0_2 gnd! 37.6fF
C986 N0836 gnd! 18.9fF
C987 PC3_3 gnd! 34.5fF
C988 N0532 gnd! 423.4fF
C989 RRAB0 gnd! 1005.1fF
C990 N0835 gnd! 18.3fF
C991 N0823 gnd! 19.1fF
C992 N0808 gnd! 18.7fF
C993 PC2_3 gnd! 34.1fF
C994 N0497 gnd! 105.2fF
C995 N0531 gnd! 456.7fF
C996 RRAB1 gnd! 797.7fF
C997 N0862 gnd! 240.2fF
C998 N0866 gnd! 478.0fF
C999 WRAB1 gnd! 702.9fF
C1000 N0543 gnd! 318.8fF
C1001 SC_A22_M22_CLK2 gnd! 720.5fF
C1002 PC1_3 gnd! 34.7fF
C1003 N0822 gnd! 20.2fF
C1004 N0807 gnd! 18.7fF
C1005 N0787 gnd! 15.3fF
C1006 PC0_3 gnd! 37.5fF
C1007 PC3_7 gnd! 36.4fF
C1008 PC2_7 gnd! 35.2fF
C1009 N0439 gnd! 416.0fF
C1010 N0426 gnd! 426.9fF
C1011 N0786 gnd! 17.0fF
C1012 PC1_7 gnd! 35.4fF
C1013 PC0_7 gnd! 38.4fF
C1014 N0410 gnd! 435.3fF
C1015 N0381 gnd! 431.9fF
C1016 N0834 gnd! 17.7fF
C1017 __INH__X11_X31_CLK1 gnd! 818.5fF
C1018 PC3_11 gnd! 32.4fF
C1019 N0444 gnd! 442.3fF
C1020 N0821 gnd! 13.9fF
C1021 N0806 gnd! 17.7fF
C1022 PC2_11 gnd! 38.9fF
C1023 PC1_11 gnd! 32.7fF
C1024 N0434 gnd! 431.3fF
C1025 N0424 gnd! 436.3fF
C1026 N0306 gnd! 182.9fF
C1027 N0717 gnd! 1210.7fF
C1028 N0295 gnd! 624.9fF
C1029 N0307 gnd! 265.5fF
C1030 N0764 gnd! 402.1fF
C1031 N0760 gnd! 121.1fF
C1032 N0752 gnd! 138.7fF
C1033 N0759 gnd! 95.7fF
C1034 N0394 gnd! 338.0fF
C1035 N0294 gnd! 182.3fF
C1036 N0305 gnd! 154.2fF
C1037 N0292 gnd! 298.0fF
C1038 N0393 gnd! 344.6fF
C1039 N0391 gnd! 319.9fF
C1040 N0392 gnd! 357.8fF
C1041 N0390 gnd! 313.5fF
C1042 N0389 gnd! 356.5fF
C1043 N0775 gnd! 355.7fF
C1044 N0779 gnd! 355.0fF
C1045 N0778 gnd! 351.1fF
C1046 WADB0 gnd! 495.9fF
C1047 N0774 gnd! 354.1fF
C1048 WADB1 gnd! 458.2fF
C1049 N0299 gnd! 12.6fF
C1050 N0303 gnd! 16.8fF
C1051 N0313 gnd! 9.5fF
C1052 N0291 gnd! 313.5fF
C1053 N0757 gnd! 92.7fF
C1054 N0763 gnd! 396.4fF
C1055 N0293 gnd! 254.2fF
C1056 N0758 gnd! 126.3fF
C1057 N0762 gnd! 402.2fF
C1058 N0756 gnd! 125.1fF
C1059 N0298 gnd! 240.2fF
C1060 N0388 gnd! 331.5fF
C1061 N0755 gnd! 97.1fF
C1062 S00536 gnd! 100.1fF
C1063 N0738 gnd! 771.5fF
C1064 S00531 gnd! 101.1fF
C1065 sync gnd! 1675.4fF
C1066 N0740 gnd! 1009.7fF
C1067 N0302 gnd! 148.4fF
C1068 N0312 gnd! 168.7fF
C1069 N0290 gnd! 276.0fF
C1070 N0387 gnd! 342.7fF
C1071 RADB0 gnd! 390.7fF
C1072 N0325 gnd! 510.6fF
C1073 N0311 gnd! 116.4fF
C1074 N0289 gnd! 217.2fF
C1075 N0753 gnd! 101.1fF
C1076 WADB2 gnd! 287.4fF
C1077 RADB2 gnd! 578.1fF
C1078 RADB1 gnd! 345.9fF
C1079 N0386 gnd! 353.2fF
C1080 Vdd gnd! 57604.7fF
C1081 N0761 gnd! 417.2fF
C1082 N0785 gnd! 16.0fF
C1083 PC0_11 gnd! 38.6fF
C1084 N0406 gnd! 440.4fF
C1085 N0385 gnd! 337.2fF
C1086 N0770 gnd! 353.6fF
C1087 N0301 gnd! 269.8fF
C1088 N0754 gnd! 123.5fF
C1089 M12_M22_CLK1__M11_M12_ gnd! 1062.7fF
C1090 D3 gnd! 3103.8fF
C1091 D2 gnd! 3244.2fF
C1092 D1 gnd! 3804.4fF
C1093 D0 gnd! 3749.5fF
C1094 test gnd! 1379.0fF
C1095 reset gnd! 1288.8fF
