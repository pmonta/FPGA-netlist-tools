* SPICE3 file created from 4001.ext - technology: nmos

.option scale=0.01u

M1000 clk2 GND GND GND efet w=9720 l=720
+ ad=6.90624e+07 pd=154800 as=2.09344e+09 ps=3.9312e+06 
M1001 clk1 GND GND GND efet w=9720 l=720
+ ad=4.71456e+07 pd=118320 as=0 ps=0 
M1002 d2 GND d2 GND efet w=17700 l=11220
+ ad=1.4963e+08 pd=299520 as=0 ps=0 
M1003 d3 GND d3 GND efet w=17880 l=11520
+ ad=1.91736e+08 pd=409920 as=0 ps=0 
M1004 sync GND GND GND efet w=9120 l=720
+ ad=1.04342e+08 pd=261840 as=0 ps=0 
M1005 GND diff_33840_166200# d3 GND efet w=93360 l=360
+ ad=0 pd=0 as=0 ps=0 
M1006 GND diff_49440_166200# d2 GND efet w=93240 l=360
+ ad=0 pd=0 as=0 ps=0 
M1007 Vdd diff_35520_136680# d3 GND efet w=43140 l=1020
+ ad=6.95491e+08 pd=1.52592e+06 as=0 ps=0 
M1008 GND diff_64920_166200# d1 GND efet w=93240 l=360
+ ad=0 pd=0 as=1.48781e+08 ps=303600 
M1009 GND diff_80400_166200# d0 GND efet w=93240 l=360
+ ad=0 pd=0 as=1.47384e+08 ps=301680 
M1010 GND diff_243360_174240# diff_243720_169800# GND efet w=35640 l=600
+ ad=0 pd=0 as=9.29232e+07 ps=147600 
M1011 GND clk1 diff_261360_171960# GND efet w=2520 l=720
+ ad=0 pd=0 as=4.4784e+06 ps=9120 
M1012 GND sync diff_243360_174240# GND efet w=7680 l=720
+ ad=0 pd=0 as=2.94048e+07 ps=60720 
M1013 diff_280200_173280# diff_275160_168600# GND GND efet w=2760 l=600
+ ad=5.2992e+06 pd=18240 as=0 ps=0 
M1014 diff_264960_142800# diff_280200_173280# GND GND efet w=4080 l=600
+ ad=7.632e+06 pd=20400 as=0 ps=0 
M1015 GND diff_243360_174240# diff_274320_171480# GND efet w=4080 l=600
+ ad=0 pd=0 as=3.9168e+06 ps=10080 
M1016 diff_261360_171960# Vdd Vdd GND efet w=720 l=960
+ ad=0 pd=0 as=0 ps=0 
M1017 diff_243360_174240# diff_266400_168600# GND GND efet w=4680 l=720
+ ad=0 pd=0 as=0 ps=0 
M1018 GND diff_100320_170280# diff_100800_168600# GND efet w=61920 l=720
+ ad=0 pd=0 as=1.94112e+08 ps=277920 
M1019 Vdd diff_165720_170280# diff_100800_168600# GND efet w=64320 l=720
+ ad=0 pd=0 as=0 ps=0 
M1020 diff_100800_168600# diff_100440_168000# diff_100800_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1021 diff_100800_168600# diff_100440_168000# diff_102840_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1022 diff_100800_168600# diff_100440_168000# diff_104880_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1023 diff_100800_168600# diff_100440_168000# diff_106920_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1024 diff_100800_168600# diff_100440_168000# diff_108960_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1025 diff_100800_168600# diff_100440_168000# diff_111000_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1026 diff_100800_168600# diff_100440_168000# diff_113040_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1027 diff_100800_168600# diff_100440_168000# diff_115080_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1028 diff_100800_168600# diff_100440_168000# diff_117120_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1029 diff_100800_168600# diff_100440_168000# diff_119160_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1030 diff_100800_168600# diff_100440_168000# diff_121200_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1031 diff_100800_168600# diff_100440_168000# diff_123240_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1032 diff_100800_168600# diff_100440_168000# diff_125280_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1033 diff_100800_168600# diff_100440_168000# diff_127320_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1034 diff_100800_168600# diff_100440_168000# diff_129360_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1035 diff_100800_168600# diff_100440_168000# diff_131400_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1036 diff_100800_168600# diff_100440_168000# diff_133440_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1037 diff_100800_168600# diff_100440_168000# diff_135480_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1038 diff_100800_168600# diff_100440_168000# diff_137520_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1039 diff_100800_168600# diff_100440_168000# diff_139560_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1040 diff_100800_168600# diff_100440_168000# diff_141600_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1041 diff_100800_168600# diff_100440_168000# diff_143640_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1042 diff_100800_168600# diff_100440_168000# diff_145680_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1043 diff_100800_168600# diff_100440_168000# diff_147720_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1044 diff_100800_168600# diff_100440_168000# diff_149760_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1045 diff_100800_168600# diff_100440_168000# diff_151800_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1046 diff_100800_168600# diff_100440_168000# diff_153840_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1047 diff_100800_168600# diff_100440_168000# diff_155880_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1048 diff_100800_168600# diff_100440_168000# diff_157920_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1049 diff_100800_168600# diff_100440_168000# diff_159960_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1050 diff_100800_168600# diff_100440_168000# diff_162000_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1051 diff_100800_168600# diff_100440_168000# diff_164040_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1052 diff_100800_168600# diff_100440_168000# diff_166080_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1053 diff_100800_168600# diff_100440_168000# diff_168120_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1054 diff_100800_168600# diff_100440_168000# diff_170160_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1055 diff_100800_168600# diff_100440_168000# diff_172200_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1056 diff_100800_168600# diff_100440_168000# diff_174240_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1057 diff_100800_168600# diff_100440_168000# diff_176280_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1058 diff_100800_168600# diff_100440_168000# diff_178320_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1059 diff_100800_168600# diff_100440_168000# diff_180360_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1060 diff_100800_168600# diff_100440_168000# diff_182400_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1061 diff_100800_168600# diff_100440_168000# diff_184440_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1062 diff_100800_168600# diff_100440_168000# diff_186480_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1063 diff_100800_168600# diff_100440_168000# diff_188520_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1064 diff_100800_168600# diff_100440_168000# diff_190560_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1065 diff_100800_168600# diff_100440_168000# diff_192600_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1066 diff_100800_168600# diff_100440_168000# diff_194640_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1067 diff_100800_168600# diff_100440_168000# diff_196680_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1068 diff_100800_168600# diff_100440_168000# diff_198720_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1069 diff_100800_168600# diff_100440_168000# diff_200760_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1070 diff_100800_168600# diff_100440_168000# diff_202800_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1071 diff_100800_168600# diff_100440_168000# diff_204840_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1072 diff_100800_168600# diff_100440_168000# diff_206880_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1073 diff_100800_168600# diff_100440_168000# diff_208920_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1074 diff_100800_168600# diff_100440_168000# diff_210960_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1075 diff_100800_168600# diff_100440_168000# diff_213000_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1076 diff_100800_168600# diff_100440_168000# diff_215040_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1077 diff_100800_168600# diff_100440_168000# diff_217080_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1078 diff_100800_168600# diff_100440_168000# diff_219120_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1079 diff_100800_168600# diff_100440_168000# diff_221160_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1080 diff_100800_168600# diff_100440_168000# diff_223200_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1081 diff_100800_168600# diff_100440_168000# diff_225240_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1082 diff_100800_168600# diff_100440_168000# diff_227280_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1083 diff_100800_168600# diff_100440_168000# diff_229320_166320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1084 diff_236760_167400# diff_236160_42720# diff_100440_168000# GND efet w=8940 l=720
+ ad=3.62016e+07 pd=68880 as=9.5616e+06 ps=23040 
M1085 Vdd Vdd diff_36600_150480# GND efet w=960 l=960
+ ad=0 pd=0 as=2.4912e+06 ps=7200 
M1086 Vdd Vdd diff_42840_150720# GND efet w=840 l=1080
+ ad=0 pd=0 as=1.9872e+06 ps=6720 
M1087 diff_36600_150480# diff_36600_150480# diff_36600_150480# GND efet w=180 l=360
+ ad=0 pd=0 as=0 ps=0 
M1088 Vdd diff_36600_150480# diff_35520_136680# GND efet w=840 l=720
+ ad=0 pd=0 as=3.02544e+07 ps=65040 
M1089 Vdd diff_42840_150720# diff_33840_166200# GND efet w=840 l=720
+ ad=0 pd=0 as=3.69504e+07 ps=76800 
M1090 diff_42840_150720# diff_42840_150720# diff_42840_150720# GND efet w=180 l=480
+ ad=0 pd=0 as=0 ps=0 
M1091 Vdd diff_51000_136680# d2 GND efet w=42960 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1092 diff_36600_150480# diff_36600_150480# diff_36600_150480# GND efet w=120 l=360
+ ad=0 pd=0 as=0 ps=0 
M1093 diff_35520_136680# diff_36600_150480# diff_35520_136680# GND efet w=4260 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1094 diff_42840_150720# diff_42840_150720# diff_42840_150720# GND efet w=120 l=600
+ ad=0 pd=0 as=0 ps=0 
M1095 Vdd Vdd diff_52080_150360# GND efet w=720 l=960
+ ad=0 pd=0 as=2.1312e+06 ps=7440 
M1096 Vdd Vdd diff_58320_150600# GND efet w=960 l=1080
+ ad=0 pd=0 as=2.2032e+06 ps=7920 
M1097 diff_52080_150360# diff_52080_150360# diff_52080_150360# GND efet w=240 l=300
+ ad=0 pd=0 as=0 ps=0 
M1098 Vdd diff_52080_150360# diff_51000_136680# GND efet w=840 l=720
+ ad=0 pd=0 as=3.02688e+07 ps=65040 
M1099 Vdd diff_58320_150600# diff_49440_166200# GND efet w=840 l=720
+ ad=0 pd=0 as=3.75696e+07 ps=77040 
M1100 diff_58320_150600# diff_58320_150600# diff_58320_150600# GND efet w=360 l=420
+ ad=0 pd=0 as=0 ps=0 
M1101 diff_52080_150360# diff_52080_150360# diff_52080_150360# GND efet w=120 l=480
+ ad=0 pd=0 as=0 ps=0 
M1102 diff_33840_166200# diff_42840_150720# diff_33840_166200# GND efet w=5700 l=660
+ ad=0 pd=0 as=0 ps=0 
M1103 diff_51000_136680# diff_52080_150360# diff_51000_136680# GND efet w=4380 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1104 diff_58320_150600# diff_58320_150600# diff_58320_150600# GND efet w=120 l=720
+ ad=0 pd=0 as=0 ps=0 
M1105 Vdd diff_66480_136560# d1 GND efet w=43080 l=720
+ ad=0 pd=0 as=0 ps=0 
M1106 Vdd Vdd diff_67320_150600# GND efet w=840 l=1080
+ ad=0 pd=0 as=1.7712e+06 ps=6480 
M1107 Vdd Vdd diff_73800_150600# GND efet w=840 l=1080
+ ad=0 pd=0 as=1.9152e+06 ps=6240 
M1108 Vdd diff_82080_136560# d0 GND efet w=42840 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1109 Vdd diff_67320_150600# diff_66480_136560# GND efet w=720 l=720
+ ad=0 pd=0 as=3.05568e+07 ps=69600 
M1110 diff_67320_150600# diff_67320_150600# diff_67320_150600# GND efet w=240 l=480
+ ad=0 pd=0 as=0 ps=0 
M1111 diff_49440_166200# diff_58320_150600# diff_49440_166200# GND efet w=5700 l=660
+ ad=0 pd=0 as=0 ps=0 
M1112 Vdd diff_73800_150600# diff_64920_166200# GND efet w=780 l=780
+ ad=0 pd=0 as=3.65616e+07 ps=76560 
M1113 diff_73800_150600# diff_73800_150600# diff_73800_150600# GND efet w=120 l=180
+ ad=0 pd=0 as=0 ps=0 
M1114 diff_67320_150600# diff_67320_150600# diff_67320_150600# GND efet w=120 l=480
+ ad=0 pd=0 as=0 ps=0 
M1115 diff_73800_150600# diff_73800_150600# diff_73800_150600# GND efet w=60 l=180
+ ad=0 pd=0 as=0 ps=0 
M1116 Vdd Vdd diff_83160_150480# GND efet w=840 l=960
+ ad=0 pd=0 as=2.1744e+06 ps=6720 
M1117 Vdd Vdd diff_88680_154680# GND efet w=840 l=960
+ ad=0 pd=0 as=1.7856e+06 ps=6000 
M1118 diff_83160_150480# diff_83160_150480# diff_83160_150480# GND efet w=60 l=180
+ ad=0 pd=0 as=0 ps=0 
M1119 Vdd diff_83160_150480# diff_82080_136560# GND efet w=720 l=720
+ ad=0 pd=0 as=3.0456e+07 ps=64800 
M1120 Vdd diff_88680_154680# diff_80400_166200# GND efet w=720 l=720
+ ad=0 pd=0 as=3.71952e+07 ps=74880 
M1121 diff_88680_154680# diff_88680_154680# diff_88680_154680# GND efet w=120 l=180
+ ad=0 pd=0 as=0 ps=0 
M1122 diff_100800_166320# diff_100440_165720# diff_100800_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1123 diff_102840_166320# diff_100440_165720# diff_102840_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1124 diff_104880_166320# diff_100440_165720# diff_104880_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1125 diff_106920_166320# diff_100440_165720# diff_106920_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1126 diff_108960_166320# diff_100440_165720# diff_108960_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1127 diff_111000_166320# diff_100440_165720# diff_111000_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1128 diff_113040_166320# diff_100440_165720# diff_113040_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1129 diff_115080_166320# diff_100440_165720# diff_115080_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1130 diff_117120_166320# diff_100440_165720# diff_117120_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1131 diff_119160_166320# diff_100440_165720# diff_119160_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1132 diff_121200_166320# diff_100440_165720# diff_121200_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1133 diff_123240_166320# diff_100440_165720# diff_123240_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1134 diff_125280_166320# diff_100440_165720# diff_125280_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1135 diff_127320_166320# diff_100440_165720# diff_127320_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1136 diff_129360_166320# diff_100440_165720# diff_129360_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1137 diff_131400_166320# diff_100440_165720# diff_131400_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1138 diff_133440_166320# diff_100440_165720# diff_133440_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1139 diff_135480_166320# diff_100440_165720# diff_135480_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1140 diff_137520_166320# diff_100440_165720# diff_137520_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1141 diff_139560_166320# diff_100440_165720# diff_139560_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1142 diff_141600_166320# diff_100440_165720# diff_141600_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1143 diff_143640_166320# diff_100440_165720# diff_143640_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1144 diff_145680_166320# diff_100440_165720# diff_145680_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1145 diff_147720_166320# diff_100440_165720# diff_147720_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1146 diff_149760_166320# diff_100440_165720# diff_149760_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1147 diff_151800_166320# diff_100440_165720# diff_151800_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1148 diff_153840_166320# diff_100440_165720# diff_153840_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1149 diff_155880_166320# diff_100440_165720# diff_155880_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1150 diff_157920_166320# diff_100440_165720# diff_157920_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1151 diff_159960_166320# diff_100440_165720# diff_159960_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1152 diff_162000_166320# diff_100440_165720# diff_162000_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1153 diff_164040_166320# diff_100440_165720# diff_164040_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1154 diff_166080_166320# diff_100440_165720# diff_166080_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1155 diff_168120_166320# diff_100440_165720# diff_168120_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1156 diff_170160_166320# diff_100440_165720# diff_170160_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1157 diff_172200_166320# diff_100440_165720# diff_172200_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1158 diff_174240_166320# diff_100440_165720# diff_174240_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1159 diff_176280_166320# diff_100440_165720# diff_176280_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1160 diff_178320_166320# diff_100440_165720# diff_178320_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1161 diff_180360_166320# diff_100440_165720# diff_180360_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1162 diff_182400_166320# diff_100440_165720# diff_182400_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1163 diff_184440_166320# diff_100440_165720# diff_184440_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1164 diff_186480_166320# diff_100440_165720# diff_186480_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1165 diff_188520_166320# diff_100440_165720# diff_188520_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1166 diff_190560_166320# diff_100440_165720# diff_190560_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1167 diff_192600_166320# diff_100440_165720# diff_192600_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1168 diff_194640_166320# diff_100440_165720# diff_194640_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1169 diff_196680_166320# diff_100440_165720# diff_196680_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1170 diff_198720_166320# diff_100440_165720# diff_198720_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1171 diff_200760_166320# diff_100440_165720# diff_200760_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1172 diff_202800_166320# diff_100440_165720# diff_202800_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1173 diff_204840_166320# diff_100440_165720# diff_204840_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1174 diff_206880_166320# diff_100440_165720# diff_206880_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1175 diff_208920_166320# diff_100440_165720# diff_208920_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1176 diff_210960_166320# diff_100440_165720# diff_210960_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1177 diff_213000_166320# diff_100440_165720# diff_213000_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1178 diff_215040_166320# diff_100440_165720# diff_215040_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1179 diff_217080_166320# diff_100440_165720# diff_217080_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1180 diff_219120_166320# diff_100440_165720# diff_219120_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1181 diff_221160_166320# diff_100440_165720# diff_221160_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1182 diff_223200_166320# diff_100440_165720# diff_223200_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1183 diff_225240_166320# diff_100440_165720# diff_225240_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1184 diff_227280_166320# diff_100440_165720# diff_227280_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1185 diff_229320_166320# diff_100440_165720# diff_229320_164160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1186 diff_100440_168000# Vdd Vdd GND efet w=600 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1187 diff_100800_164160# diff_100440_163560# diff_100800_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1188 diff_102840_164160# diff_100440_163560# diff_102840_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1189 diff_104880_164160# diff_100440_163560# diff_104880_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1190 diff_106920_164160# diff_100440_163560# diff_106920_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1191 diff_108960_164160# diff_100440_163560# diff_108960_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1192 diff_111000_164160# diff_100440_163560# diff_111000_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1193 diff_113040_164160# diff_100440_163560# diff_113040_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1194 diff_115080_164160# diff_100440_163560# diff_115080_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1195 diff_117120_164160# diff_100440_163560# diff_117120_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1196 diff_119160_164160# diff_100440_163560# diff_119160_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1197 diff_121200_164160# diff_100440_163560# diff_121200_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1198 diff_123240_164160# diff_100440_163560# diff_123240_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1199 diff_125280_164160# diff_100440_163560# diff_125280_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1200 diff_127320_164160# diff_100440_163560# diff_127320_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1201 diff_129360_164160# diff_100440_163560# diff_129360_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1202 diff_131400_164160# diff_100440_163560# diff_131400_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1203 diff_133440_164160# diff_100440_163560# diff_133440_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1204 diff_135480_164160# diff_100440_163560# diff_135480_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1205 diff_137520_164160# diff_100440_163560# diff_137520_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1206 diff_139560_164160# diff_100440_163560# diff_139560_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1207 diff_141600_164160# diff_100440_163560# diff_141600_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1208 diff_143640_164160# diff_100440_163560# diff_143640_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1209 diff_145680_164160# diff_100440_163560# diff_145680_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1210 diff_147720_164160# diff_100440_163560# diff_147720_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1211 diff_149760_164160# diff_100440_163560# diff_149760_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1212 diff_151800_164160# diff_100440_163560# diff_151800_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1213 diff_153840_164160# diff_100440_163560# diff_153840_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1214 diff_155880_164160# diff_100440_163560# diff_155880_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1215 diff_157920_164160# diff_100440_163560# diff_157920_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1216 diff_159960_164160# diff_100440_163560# diff_159960_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1217 diff_162000_164160# diff_100440_163560# diff_162000_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1218 diff_164040_164160# diff_100440_163560# diff_164040_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1219 diff_166080_164160# diff_100440_163560# diff_166080_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1220 diff_168120_164160# diff_100440_163560# diff_168120_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1221 diff_170160_164160# diff_100440_163560# diff_170160_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1222 diff_172200_164160# diff_100440_163560# diff_172200_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1223 diff_174240_164160# diff_100440_163560# diff_174240_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1224 diff_176280_164160# diff_100440_163560# diff_176280_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1225 diff_178320_164160# diff_100440_163560# diff_178320_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1226 diff_180360_164160# diff_100440_163560# diff_180360_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1227 diff_182400_164160# diff_100440_163560# diff_182400_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1228 diff_184440_164160# diff_100440_163560# diff_184440_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1229 diff_186480_164160# diff_100440_163560# diff_186480_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1230 diff_188520_164160# diff_100440_163560# diff_188520_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1231 diff_190560_164160# diff_100440_163560# diff_190560_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1232 diff_192600_164160# diff_100440_163560# diff_192600_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1233 diff_194640_164160# diff_100440_163560# diff_194640_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1234 diff_196680_164160# diff_100440_163560# diff_196680_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1235 diff_198720_164160# diff_100440_163560# diff_198720_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1236 diff_200760_164160# diff_100440_163560# diff_200760_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1237 diff_202800_164160# diff_100440_163560# diff_202800_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1238 diff_204840_164160# diff_100440_163560# diff_204840_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1239 diff_206880_164160# diff_100440_163560# diff_206880_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1240 diff_208920_164160# diff_100440_163560# diff_208920_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1241 diff_210960_164160# diff_100440_163560# diff_210960_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1242 diff_213000_164160# diff_100440_163560# diff_213000_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1243 diff_215040_164160# diff_100440_163560# diff_215040_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1244 diff_217080_164160# diff_100440_163560# diff_217080_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1245 diff_219120_164160# diff_100440_163560# diff_219120_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1246 diff_221160_164160# diff_100440_163560# diff_221160_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1247 diff_223200_164160# diff_100440_163560# diff_223200_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1248 diff_225240_164160# diff_100440_163560# diff_225240_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1249 diff_227280_164160# diff_100440_163560# diff_227280_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1250 diff_229320_164160# diff_100440_163560# diff_229320_161880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1251 Vdd Vdd diff_100440_161280# GND efet w=600 l=1200
+ ad=0 pd=0 as=8.5104e+06 ps=25920 
M1252 diff_100800_161880# diff_100440_161280# diff_100800_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1253 diff_102840_161880# diff_100440_161280# diff_102840_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1254 diff_104880_161880# diff_100440_161280# diff_104880_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1255 diff_106920_161880# diff_100440_161280# diff_106920_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1256 diff_108960_161880# diff_100440_161280# diff_108960_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1257 diff_111000_161880# diff_100440_161280# diff_111000_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1258 diff_113040_161880# diff_100440_161280# diff_113040_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1259 diff_115080_161880# diff_100440_161280# diff_115080_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1260 diff_117120_161880# diff_100440_161280# diff_117120_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1261 diff_119160_161880# diff_100440_161280# diff_119160_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1262 diff_121200_161880# diff_100440_161280# diff_121200_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1263 diff_123240_161880# diff_100440_161280# diff_123240_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1264 diff_125280_161880# diff_100440_161280# diff_125280_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1265 diff_127320_161880# diff_100440_161280# diff_127320_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1266 diff_129360_161880# diff_100440_161280# diff_129360_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1267 diff_131400_161880# diff_100440_161280# diff_131400_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1268 diff_133440_161880# diff_100440_161280# diff_133440_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1269 diff_135480_161880# diff_100440_161280# diff_135480_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1270 diff_137520_161880# diff_100440_161280# diff_137520_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1271 diff_139560_161880# diff_100440_161280# diff_139560_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1272 diff_141600_161880# diff_100440_161280# diff_141600_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1273 diff_143640_161880# diff_100440_161280# diff_143640_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1274 diff_145680_161880# diff_100440_161280# diff_145680_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1275 diff_147720_161880# diff_100440_161280# diff_147720_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1276 diff_149760_161880# diff_100440_161280# diff_149760_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1277 diff_151800_161880# diff_100440_161280# diff_151800_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1278 diff_153840_161880# diff_100440_161280# diff_153840_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1279 diff_155880_161880# diff_100440_161280# diff_155880_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1280 diff_157920_161880# diff_100440_161280# diff_157920_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1281 diff_159960_161880# diff_100440_161280# diff_159960_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1282 diff_162000_161880# diff_100440_161280# diff_162000_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1283 diff_164040_161880# diff_100440_161280# diff_164040_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1284 diff_166080_161880# diff_100440_161280# diff_166080_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1285 diff_168120_161880# diff_100440_161280# diff_168120_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1286 diff_170160_161880# diff_100440_161280# diff_170160_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1287 diff_172200_161880# diff_100440_161280# diff_172200_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1288 diff_174240_161880# diff_100440_161280# diff_174240_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1289 diff_176280_161880# diff_100440_161280# diff_176280_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1290 diff_178320_161880# diff_100440_161280# diff_178320_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1291 diff_180360_161880# diff_100440_161280# diff_180360_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1292 diff_182400_161880# diff_100440_161280# diff_182400_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1293 diff_184440_161880# diff_100440_161280# diff_184440_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1294 diff_186480_161880# diff_100440_161280# diff_186480_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1295 diff_188520_161880# diff_100440_161280# diff_188520_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1296 diff_190560_161880# diff_100440_161280# diff_190560_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1297 diff_192600_161880# diff_100440_161280# diff_192600_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1298 diff_194640_161880# diff_100440_161280# diff_194640_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1299 diff_196680_161880# diff_100440_161280# diff_196680_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1300 diff_198720_161880# diff_100440_161280# diff_198720_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1301 diff_200760_161880# diff_100440_161280# diff_200760_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1302 diff_202800_161880# diff_100440_161280# diff_202800_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1303 diff_204840_161880# diff_100440_161280# diff_204840_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1304 diff_206880_161880# diff_100440_161280# diff_206880_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1305 diff_208920_161880# diff_100440_161280# diff_208920_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1306 diff_210960_161880# diff_100440_161280# diff_210960_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1307 diff_213000_161880# diff_100440_161280# diff_213000_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1308 diff_215040_161880# diff_100440_161280# diff_215040_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1309 diff_217080_161880# diff_100440_161280# diff_217080_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1310 diff_219120_161880# diff_100440_161280# diff_219120_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1311 diff_221160_161880# diff_100440_161280# diff_221160_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1312 diff_223200_161880# diff_100440_161280# diff_223200_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1313 diff_225240_161880# diff_100440_161280# diff_225240_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1314 diff_227280_161880# diff_100440_161280# diff_227280_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1315 diff_229320_161880# diff_100440_161280# diff_229320_159720# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1316 diff_100440_161280# diff_238440_42720# diff_236760_167400# GND efet w=7440 l=600
+ ad=0 pd=0 as=0 ps=0 
M1317 diff_236760_167400# diff_241320_99600# diff_100440_165720# GND efet w=8280 l=720
+ ad=0 pd=0 as=1.08e+07 ps=22320 
M1318 diff_100440_165720# Vdd Vdd GND efet w=720 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1319 Vdd Vdd diff_100440_163560# GND efet w=720 l=1200
+ ad=0 pd=0 as=9.4176e+06 ps=24720 
M1320 diff_100800_159720# diff_100440_159120# diff_100800_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1321 diff_102840_159720# diff_100440_159120# diff_102840_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1322 diff_104880_159720# diff_100440_159120# diff_104880_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1323 diff_106920_159720# diff_100440_159120# diff_106920_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1324 diff_108960_159720# diff_100440_159120# diff_108960_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1325 diff_111000_159720# diff_100440_159120# diff_111000_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1326 diff_113040_159720# diff_100440_159120# diff_113040_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1327 diff_115080_159720# diff_100440_159120# diff_115080_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1328 diff_117120_159720# diff_100440_159120# diff_117120_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1329 diff_119160_159720# diff_100440_159120# diff_119160_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1330 diff_121200_159720# diff_100440_159120# diff_121200_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1331 diff_123240_159720# diff_100440_159120# diff_123240_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1332 diff_125280_159720# diff_100440_159120# diff_125280_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1333 diff_127320_159720# diff_100440_159120# diff_127320_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1334 diff_129360_159720# diff_100440_159120# diff_129360_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1335 diff_131400_159720# diff_100440_159120# diff_131400_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1336 diff_133440_159720# diff_100440_159120# diff_133440_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1337 diff_135480_159720# diff_100440_159120# diff_135480_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1338 diff_137520_159720# diff_100440_159120# diff_137520_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1339 diff_139560_159720# diff_100440_159120# diff_139560_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1340 diff_141600_159720# diff_100440_159120# diff_141600_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1341 diff_143640_159720# diff_100440_159120# diff_143640_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1342 diff_145680_159720# diff_100440_159120# diff_145680_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1343 diff_147720_159720# diff_100440_159120# diff_147720_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1344 diff_149760_159720# diff_100440_159120# diff_149760_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1345 diff_151800_159720# diff_100440_159120# diff_151800_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1346 diff_153840_159720# diff_100440_159120# diff_153840_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1347 diff_155880_159720# diff_100440_159120# diff_155880_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1348 diff_157920_159720# diff_100440_159120# diff_157920_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1349 diff_159960_159720# diff_100440_159120# diff_159960_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1350 diff_162000_159720# diff_100440_159120# diff_162000_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1351 diff_164040_159720# diff_100440_159120# diff_164040_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1352 diff_166080_159720# diff_100440_159120# diff_166080_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1353 diff_168120_159720# diff_100440_159120# diff_168120_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1354 diff_170160_159720# diff_100440_159120# diff_170160_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1355 diff_172200_159720# diff_100440_159120# diff_172200_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1356 diff_174240_159720# diff_100440_159120# diff_174240_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1357 diff_176280_159720# diff_100440_159120# diff_176280_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1358 diff_178320_159720# diff_100440_159120# diff_178320_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1359 diff_180360_159720# diff_100440_159120# diff_180360_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1360 diff_182400_159720# diff_100440_159120# diff_182400_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1361 diff_184440_159720# diff_100440_159120# diff_184440_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1362 diff_186480_159720# diff_100440_159120# diff_186480_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1363 diff_188520_159720# diff_100440_159120# diff_188520_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1364 diff_190560_159720# diff_100440_159120# diff_190560_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1365 diff_192600_159720# diff_100440_159120# diff_192600_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1366 diff_194640_159720# diff_100440_159120# diff_194640_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1367 diff_196680_159720# diff_100440_159120# diff_196680_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1368 diff_198720_159720# diff_100440_159120# diff_198720_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1369 diff_200760_159720# diff_100440_159120# diff_200760_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1370 diff_202800_159720# diff_100440_159120# diff_202800_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1371 diff_204840_159720# diff_100440_159120# diff_204840_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1372 diff_206880_159720# diff_100440_159120# diff_206880_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1373 diff_208920_159720# diff_100440_159120# diff_208920_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1374 diff_210960_159720# diff_100440_159120# diff_210960_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1375 diff_213000_159720# diff_100440_159120# diff_213000_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1376 diff_215040_159720# diff_100440_159120# diff_215040_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1377 diff_217080_159720# diff_100440_159120# diff_217080_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1378 diff_219120_159720# diff_100440_159120# diff_219120_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1379 diff_221160_159720# diff_100440_159120# diff_221160_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1380 diff_223200_159720# diff_100440_159120# diff_223200_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1381 diff_225240_159720# diff_100440_159120# diff_225240_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1382 diff_227280_159720# diff_100440_159120# diff_227280_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1383 diff_229320_159720# diff_100440_159120# diff_229320_157440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1384 diff_236760_158520# diff_236160_42720# diff_100440_159120# GND efet w=8760 l=660
+ ad=3.8232e+07 pd=73200 as=8.8992e+06 ps=22560 
M1385 diff_100440_163560# diff_243120_97920# diff_236760_167400# GND efet w=7920 l=600
+ ad=0 pd=0 as=0 ps=0 
M1386 diff_100800_157440# diff_100440_156840# diff_100800_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1387 diff_102840_157440# diff_100440_156840# diff_102840_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1388 diff_104880_157440# diff_100440_156840# diff_104880_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1389 diff_106920_157440# diff_100440_156840# diff_106920_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1390 diff_108960_157440# diff_100440_156840# diff_108960_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1391 diff_111000_157440# diff_100440_156840# diff_111000_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1392 diff_113040_157440# diff_100440_156840# diff_113040_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1393 diff_115080_157440# diff_100440_156840# diff_115080_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1394 diff_117120_157440# diff_100440_156840# diff_117120_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1395 diff_119160_157440# diff_100440_156840# diff_119160_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1396 diff_121200_157440# diff_100440_156840# diff_121200_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1397 diff_123240_157440# diff_100440_156840# diff_123240_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1398 diff_125280_157440# diff_100440_156840# diff_125280_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1399 diff_127320_157440# diff_100440_156840# diff_127320_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1400 diff_129360_157440# diff_100440_156840# diff_129360_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1401 diff_131400_157440# diff_100440_156840# diff_131400_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1402 diff_133440_157440# diff_100440_156840# diff_133440_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1403 diff_135480_157440# diff_100440_156840# diff_135480_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1404 diff_137520_157440# diff_100440_156840# diff_137520_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1405 diff_139560_157440# diff_100440_156840# diff_139560_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1406 diff_141600_157440# diff_100440_156840# diff_141600_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1407 diff_143640_157440# diff_100440_156840# diff_143640_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1408 diff_145680_157440# diff_100440_156840# diff_145680_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1409 diff_147720_157440# diff_100440_156840# diff_147720_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1410 diff_149760_157440# diff_100440_156840# diff_149760_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1411 diff_151800_157440# diff_100440_156840# diff_151800_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1412 diff_153840_157440# diff_100440_156840# diff_153840_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1413 diff_155880_157440# diff_100440_156840# diff_155880_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1414 diff_157920_157440# diff_100440_156840# diff_157920_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1415 diff_159960_157440# diff_100440_156840# diff_159960_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1416 diff_162000_157440# diff_100440_156840# diff_162000_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1417 diff_164040_157440# diff_100440_156840# diff_164040_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1418 diff_166080_157440# diff_100440_156840# diff_166080_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1419 diff_168120_157440# diff_100440_156840# diff_168120_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1420 diff_170160_157440# diff_100440_156840# diff_170160_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1421 diff_172200_157440# diff_100440_156840# diff_172200_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1422 diff_174240_157440# diff_100440_156840# diff_174240_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1423 diff_176280_157440# diff_100440_156840# diff_176280_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1424 diff_178320_157440# diff_100440_156840# diff_178320_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1425 diff_180360_157440# diff_100440_156840# diff_180360_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1426 diff_182400_157440# diff_100440_156840# diff_182400_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1427 diff_184440_157440# diff_100440_156840# diff_184440_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1428 diff_186480_157440# diff_100440_156840# diff_186480_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1429 diff_188520_157440# diff_100440_156840# diff_188520_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1430 diff_190560_157440# diff_100440_156840# diff_190560_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1431 diff_192600_157440# diff_100440_156840# diff_192600_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1432 diff_194640_157440# diff_100440_156840# diff_194640_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1433 diff_196680_157440# diff_100440_156840# diff_196680_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1434 diff_198720_157440# diff_100440_156840# diff_198720_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1435 diff_200760_157440# diff_100440_156840# diff_200760_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1436 diff_202800_157440# diff_100440_156840# diff_202800_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1437 diff_204840_157440# diff_100440_156840# diff_204840_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1438 diff_206880_157440# diff_100440_156840# diff_206880_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1439 diff_208920_157440# diff_100440_156840# diff_208920_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1440 diff_210960_157440# diff_100440_156840# diff_210960_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1441 diff_213000_157440# diff_100440_156840# diff_213000_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1442 diff_215040_157440# diff_100440_156840# diff_215040_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1443 diff_217080_157440# diff_100440_156840# diff_217080_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1444 diff_219120_157440# diff_100440_156840# diff_219120_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1445 diff_221160_157440# diff_100440_156840# diff_221160_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1446 diff_223200_157440# diff_100440_156840# diff_223200_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1447 diff_225240_157440# diff_100440_156840# diff_225240_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1448 diff_227280_157440# diff_100440_156840# diff_227280_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1449 diff_229320_157440# diff_100440_156840# diff_229320_155280# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1450 diff_83160_150480# diff_83160_150480# diff_83160_150480# GND efet w=60 l=180
+ ad=0 pd=0 as=0 ps=0 
M1451 diff_35520_136680# diff_33840_166200# GND GND efet w=9720 l=720
+ ad=0 pd=0 as=0 ps=0 
M1452 diff_33840_166200# diff_40800_144840# GND GND efet w=18720 l=720
+ ad=0 pd=0 as=0 ps=0 
M1453 diff_66480_136560# diff_67320_150600# diff_66480_136560# GND efet w=6120 l=360
+ ad=0 pd=0 as=0 ps=0 
M1454 diff_64920_166200# diff_73800_150600# diff_64920_166200# GND efet w=5700 l=780
+ ad=0 pd=0 as=0 ps=0 
M1455 GND diff_18960_80400# diff_35520_136680# GND efet w=18960 l=720
+ ad=0 pd=0 as=0 ps=0 
M1456 diff_51000_136680# diff_49440_166200# GND GND efet w=9720 l=720
+ ad=0 pd=0 as=0 ps=0 
M1457 diff_49440_166200# diff_56280_144840# GND GND efet w=18840 l=720
+ ad=0 pd=0 as=0 ps=0 
M1458 diff_82080_136560# diff_83160_150480# diff_82080_136560# GND efet w=4260 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1459 diff_88680_154680# diff_88680_154680# diff_88680_154680# GND efet w=60 l=180
+ ad=0 pd=0 as=0 ps=0 
M1460 diff_100440_159120# Vdd Vdd GND efet w=600 l=1320
+ ad=0 pd=0 as=0 ps=0 
M1461 diff_100800_155280# diff_100440_154680# diff_100800_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1462 diff_102840_155280# diff_100440_154680# diff_102840_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1463 diff_104880_155280# diff_100440_154680# diff_104880_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1464 diff_106920_155280# diff_100440_154680# diff_106920_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1465 diff_108960_155280# diff_100440_154680# diff_108960_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1466 diff_111000_155280# diff_100440_154680# diff_111000_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1467 diff_113040_155280# diff_100440_154680# diff_113040_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1468 diff_115080_155280# diff_100440_154680# diff_115080_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1469 diff_117120_155280# diff_100440_154680# diff_117120_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1470 diff_119160_155280# diff_100440_154680# diff_119160_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1471 diff_121200_155280# diff_100440_154680# diff_121200_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1472 diff_123240_155280# diff_100440_154680# diff_123240_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1473 diff_125280_155280# diff_100440_154680# diff_125280_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1474 diff_127320_155280# diff_100440_154680# diff_127320_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1475 diff_129360_155280# diff_100440_154680# diff_129360_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1476 diff_131400_155280# diff_100440_154680# diff_131400_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1477 diff_133440_155280# diff_100440_154680# diff_133440_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1478 diff_135480_155280# diff_100440_154680# diff_135480_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1479 diff_137520_155280# diff_100440_154680# diff_137520_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1480 diff_139560_155280# diff_100440_154680# diff_139560_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1481 diff_141600_155280# diff_100440_154680# diff_141600_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1482 diff_143640_155280# diff_100440_154680# diff_143640_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1483 diff_145680_155280# diff_100440_154680# diff_145680_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1484 diff_147720_155280# diff_100440_154680# diff_147720_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1485 diff_149760_155280# diff_100440_154680# diff_149760_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1486 diff_151800_155280# diff_100440_154680# diff_151800_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1487 diff_153840_155280# diff_100440_154680# diff_153840_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1488 diff_155880_155280# diff_100440_154680# diff_155880_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1489 diff_157920_155280# diff_100440_154680# diff_157920_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1490 diff_159960_155280# diff_100440_154680# diff_159960_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1491 diff_162000_155280# diff_100440_154680# diff_162000_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1492 diff_164040_155280# diff_100440_154680# diff_164040_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1493 diff_166080_155280# diff_100440_154680# diff_166080_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1494 diff_168120_155280# diff_100440_154680# diff_168120_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1495 diff_170160_155280# diff_100440_154680# diff_170160_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1496 diff_172200_155280# diff_100440_154680# diff_172200_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1497 diff_174240_155280# diff_100440_154680# diff_174240_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1498 diff_176280_155280# diff_100440_154680# diff_176280_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1499 diff_178320_155280# diff_100440_154680# diff_178320_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1500 diff_180360_155280# diff_100440_154680# diff_180360_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1501 diff_182400_155280# diff_100440_154680# diff_182400_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1502 diff_184440_155280# diff_100440_154680# diff_184440_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1503 diff_186480_155280# diff_100440_154680# diff_186480_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1504 diff_188520_155280# diff_100440_154680# diff_188520_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1505 diff_190560_155280# diff_100440_154680# diff_190560_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1506 diff_192600_155280# diff_100440_154680# diff_192600_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1507 diff_194640_155280# diff_100440_154680# diff_194640_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1508 diff_196680_155280# diff_100440_154680# diff_196680_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1509 diff_198720_155280# diff_100440_154680# diff_198720_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1510 diff_200760_155280# diff_100440_154680# diff_200760_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1511 diff_202800_155280# diff_100440_154680# diff_202800_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1512 diff_204840_155280# diff_100440_154680# diff_204840_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1513 diff_206880_155280# diff_100440_154680# diff_206880_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1514 diff_208920_155280# diff_100440_154680# diff_208920_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1515 diff_210960_155280# diff_100440_154680# diff_210960_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1516 diff_213000_155280# diff_100440_154680# diff_213000_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1517 diff_215040_155280# diff_100440_154680# diff_215040_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1518 diff_217080_155280# diff_100440_154680# diff_217080_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1519 diff_219120_155280# diff_100440_154680# diff_219120_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1520 diff_221160_155280# diff_100440_154680# diff_221160_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1521 diff_223200_155280# diff_100440_154680# diff_223200_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1522 diff_225240_155280# diff_100440_154680# diff_225240_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1523 diff_227280_155280# diff_100440_154680# diff_227280_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1524 diff_229320_155280# diff_100440_154680# diff_229320_153000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1525 diff_80400_166200# diff_88680_154680# diff_80400_166200# GND efet w=5040 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1526 Vdd Vdd diff_100440_152400# GND efet w=600 l=1320
+ ad=0 pd=0 as=8.5104e+06 ps=25920 
M1527 diff_100800_153000# diff_100440_152400# diff_100800_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1528 diff_102840_153000# diff_100440_152400# diff_102840_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1529 diff_104880_153000# diff_100440_152400# diff_104880_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1530 diff_106920_153000# diff_100440_152400# diff_106920_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1531 diff_108960_153000# diff_100440_152400# diff_108960_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1532 diff_111000_153000# diff_100440_152400# diff_111000_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1533 diff_113040_153000# diff_100440_152400# diff_113040_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1534 diff_115080_153000# diff_100440_152400# diff_115080_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1535 diff_117120_153000# diff_100440_152400# diff_117120_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1536 diff_119160_153000# diff_100440_152400# diff_119160_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1537 diff_121200_153000# diff_100440_152400# diff_121200_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1538 diff_123240_153000# diff_100440_152400# diff_123240_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1539 diff_125280_153000# diff_100440_152400# diff_125280_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1540 diff_127320_153000# diff_100440_152400# diff_127320_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1541 diff_129360_153000# diff_100440_152400# diff_129360_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1542 diff_131400_153000# diff_100440_152400# diff_131400_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1543 diff_133440_153000# diff_100440_152400# diff_133440_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1544 diff_135480_153000# diff_100440_152400# diff_135480_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1545 diff_137520_153000# diff_100440_152400# diff_137520_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1546 diff_139560_153000# diff_100440_152400# diff_139560_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1547 diff_141600_153000# diff_100440_152400# diff_141600_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1548 diff_143640_153000# diff_100440_152400# diff_143640_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1549 diff_145680_153000# diff_100440_152400# diff_145680_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1550 diff_147720_153000# diff_100440_152400# diff_147720_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1551 diff_149760_153000# diff_100440_152400# diff_149760_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1552 diff_151800_153000# diff_100440_152400# diff_151800_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1553 diff_153840_153000# diff_100440_152400# diff_153840_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1554 diff_155880_153000# diff_100440_152400# diff_155880_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1555 diff_157920_153000# diff_100440_152400# diff_157920_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1556 diff_159960_153000# diff_100440_152400# diff_159960_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1557 diff_162000_153000# diff_100440_152400# diff_162000_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1558 diff_164040_153000# diff_100440_152400# diff_164040_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1559 diff_166080_153000# diff_100440_152400# diff_166080_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1560 diff_168120_153000# diff_100440_152400# diff_168120_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1561 diff_170160_153000# diff_100440_152400# diff_170160_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1562 diff_172200_153000# diff_100440_152400# diff_172200_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1563 diff_174240_153000# diff_100440_152400# diff_174240_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1564 diff_176280_153000# diff_100440_152400# diff_176280_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1565 diff_178320_153000# diff_100440_152400# diff_178320_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1566 diff_180360_153000# diff_100440_152400# diff_180360_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1567 diff_182400_153000# diff_100440_152400# diff_182400_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1568 diff_184440_153000# diff_100440_152400# diff_184440_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1569 diff_186480_153000# diff_100440_152400# diff_186480_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1570 diff_188520_153000# diff_100440_152400# diff_188520_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1571 diff_190560_153000# diff_100440_152400# diff_190560_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1572 diff_192600_153000# diff_100440_152400# diff_192600_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1573 diff_194640_153000# diff_100440_152400# diff_194640_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1574 diff_196680_153000# diff_100440_152400# diff_196680_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1575 diff_198720_153000# diff_100440_152400# diff_198720_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1576 diff_200760_153000# diff_100440_152400# diff_200760_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1577 diff_202800_153000# diff_100440_152400# diff_202800_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1578 diff_204840_153000# diff_100440_152400# diff_204840_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1579 diff_206880_153000# diff_100440_152400# diff_206880_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1580 diff_208920_153000# diff_100440_152400# diff_208920_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1581 diff_210960_153000# diff_100440_152400# diff_210960_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1582 diff_213000_153000# diff_100440_152400# diff_213000_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1583 diff_215040_153000# diff_100440_152400# diff_215040_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1584 diff_217080_153000# diff_100440_152400# diff_217080_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1585 diff_219120_153000# diff_100440_152400# diff_219120_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1586 diff_221160_153000# diff_100440_152400# diff_221160_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1587 diff_223200_153000# diff_100440_152400# diff_223200_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1588 diff_225240_153000# diff_100440_152400# diff_225240_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1589 diff_227280_153000# diff_100440_152400# diff_227280_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1590 diff_229320_153000# diff_100440_152400# diff_229320_150840# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1591 diff_100440_152400# diff_238440_42720# diff_236760_158520# GND efet w=7440 l=600
+ ad=0 pd=0 as=0 ps=0 
M1592 diff_236760_158520# diff_241320_99600# diff_100440_156840# GND efet w=8460 l=660
+ ad=0 pd=0 as=1.1232e+07 ps=22320 
M1593 diff_100440_156840# Vdd Vdd GND efet w=720 l=1440
+ ad=0 pd=0 as=0 ps=0 
M1594 Vdd Vdd diff_100440_154680# GND efet w=720 l=1320
+ ad=0 pd=0 as=9.4176e+06 ps=24720 
M1595 diff_100800_150840# diff_100440_150240# diff_100800_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1596 diff_102840_150840# diff_100440_150240# diff_102840_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1597 diff_104880_150840# diff_100440_150240# diff_104880_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1598 diff_106920_150840# diff_100440_150240# diff_106920_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1599 diff_108960_150840# diff_100440_150240# diff_108960_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1600 diff_111000_150840# diff_100440_150240# diff_111000_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1601 diff_113040_150840# diff_100440_150240# diff_113040_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1602 diff_115080_150840# diff_100440_150240# diff_115080_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1603 diff_117120_150840# diff_100440_150240# diff_117120_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1604 diff_119160_150840# diff_100440_150240# diff_119160_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1605 diff_121200_150840# diff_100440_150240# diff_121200_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1606 diff_123240_150840# diff_100440_150240# diff_123240_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1607 diff_125280_150840# diff_100440_150240# diff_125280_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1608 diff_127320_150840# diff_100440_150240# diff_127320_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1609 diff_129360_150840# diff_100440_150240# diff_129360_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1610 diff_131400_150840# diff_100440_150240# diff_131400_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1611 diff_133440_150840# diff_100440_150240# diff_133440_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1612 diff_135480_150840# diff_100440_150240# diff_135480_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1613 diff_137520_150840# diff_100440_150240# diff_137520_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1614 diff_139560_150840# diff_100440_150240# diff_139560_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1615 diff_141600_150840# diff_100440_150240# diff_141600_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1616 diff_143640_150840# diff_100440_150240# diff_143640_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1617 diff_145680_150840# diff_100440_150240# diff_145680_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1618 diff_147720_150840# diff_100440_150240# diff_147720_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1619 diff_149760_150840# diff_100440_150240# diff_149760_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1620 diff_151800_150840# diff_100440_150240# diff_151800_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1621 diff_153840_150840# diff_100440_150240# diff_153840_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1622 diff_155880_150840# diff_100440_150240# diff_155880_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1623 diff_157920_150840# diff_100440_150240# diff_157920_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1624 diff_159960_150840# diff_100440_150240# diff_159960_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1625 diff_162000_150840# diff_100440_150240# diff_162000_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1626 diff_164040_150840# diff_100440_150240# diff_164040_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1627 diff_166080_150840# diff_100440_150240# diff_166080_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1628 diff_168120_150840# diff_100440_150240# diff_168120_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1629 diff_170160_150840# diff_100440_150240# diff_170160_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1630 diff_172200_150840# diff_100440_150240# diff_172200_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1631 diff_174240_150840# diff_100440_150240# diff_174240_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1632 diff_176280_150840# diff_100440_150240# diff_176280_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1633 diff_178320_150840# diff_100440_150240# diff_178320_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1634 diff_180360_150840# diff_100440_150240# diff_180360_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1635 diff_182400_150840# diff_100440_150240# diff_182400_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1636 diff_184440_150840# diff_100440_150240# diff_184440_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1637 diff_186480_150840# diff_100440_150240# diff_186480_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1638 diff_188520_150840# diff_100440_150240# diff_188520_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1639 diff_190560_150840# diff_100440_150240# diff_190560_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1640 diff_192600_150840# diff_100440_150240# diff_192600_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1641 diff_194640_150840# diff_100440_150240# diff_194640_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1642 diff_196680_150840# diff_100440_150240# diff_196680_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1643 diff_198720_150840# diff_100440_150240# diff_198720_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1644 diff_200760_150840# diff_100440_150240# diff_200760_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1645 diff_202800_150840# diff_100440_150240# diff_202800_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1646 diff_204840_150840# diff_100440_150240# diff_204840_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1647 diff_206880_150840# diff_100440_150240# diff_206880_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1648 diff_208920_150840# diff_100440_150240# diff_208920_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1649 diff_210960_150840# diff_100440_150240# diff_210960_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1650 diff_213000_150840# diff_100440_150240# diff_213000_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1651 diff_215040_150840# diff_100440_150240# diff_215040_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1652 diff_217080_150840# diff_100440_150240# diff_217080_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1653 diff_219120_150840# diff_100440_150240# diff_219120_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1654 diff_221160_150840# diff_100440_150240# diff_221160_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1655 diff_223200_150840# diff_100440_150240# diff_223200_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1656 diff_225240_150840# diff_100440_150240# diff_225240_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1657 diff_227280_150840# diff_100440_150240# diff_227280_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1658 diff_229320_150840# diff_100440_150240# diff_229320_148560# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1659 diff_33840_166200# diff_18960_80400# GND GND efet w=19080 l=720
+ ad=0 pd=0 as=0 ps=0 
M1660 GND diff_18960_80400# diff_51000_136680# GND efet w=18960 l=720
+ ad=0 pd=0 as=0 ps=0 
M1661 diff_66480_136560# diff_64920_166200# GND GND efet w=9720 l=720
+ ad=0 pd=0 as=0 ps=0 
M1662 diff_64920_166200# diff_71880_144840# GND GND efet w=18840 l=720
+ ad=0 pd=0 as=0 ps=0 
M1663 diff_49440_166200# diff_18960_80400# GND GND efet w=19080 l=720
+ ad=0 pd=0 as=0 ps=0 
M1664 GND diff_18960_80400# diff_66480_136560# GND efet w=19080 l=720
+ ad=0 pd=0 as=0 ps=0 
M1665 diff_82080_136560# diff_80400_166200# GND GND efet w=9720 l=720
+ ad=0 pd=0 as=0 ps=0 
M1666 diff_80400_166200# diff_87360_144840# GND GND efet w=18840 l=720
+ ad=0 pd=0 as=0 ps=0 
M1667 diff_236760_149400# diff_236160_42720# diff_100440_150240# GND efet w=8820 l=720
+ ad=3.86208e+07 pd=71760 as=9.4176e+06 ps=23040 
M1668 diff_100440_154680# diff_243120_97920# diff_236760_158520# GND efet w=7920 l=600
+ ad=0 pd=0 as=0 ps=0 
M1669 diff_243720_169800# diff_248880_85320# diff_236760_158520# GND efet w=15480 l=720
+ ad=0 pd=0 as=0 ps=0 
M1670 diff_236760_167400# diff_250560_91920# diff_243720_169800# GND efet w=16080 l=720
+ ad=0 pd=0 as=0 ps=0 
M1671 diff_243360_174240# Vdd Vdd GND efet w=720 l=1440
+ ad=0 pd=0 as=0 ps=0 
M1672 diff_275160_168600# diff_275160_168600# diff_275160_168600# GND efet w=120 l=180
+ ad=8.5968e+06 pd=23280 as=0 ps=0 
M1673 diff_274320_171480# diff_266400_142200# diff_274320_170280# GND efet w=4080 l=600
+ ad=0 pd=0 as=4.3776e+06 ps=12000 
M1674 diff_275160_168600# diff_275160_168600# diff_275160_168600# GND efet w=60 l=120
+ ad=0 pd=0 as=0 ps=0 
M1675 GND diff_268200_169080# diff_266400_168600# GND efet w=2280 l=600
+ ad=0 pd=0 as=7.4304e+06 ps=21600 
M1676 diff_274320_170280# diff_264960_151920# diff_275160_168600# GND efet w=4200 l=600
+ ad=0 pd=0 as=0 ps=0 
M1677 diff_266400_168600# diff_266400_168600# diff_266400_168600# GND efet w=120 l=120
+ ad=0 pd=0 as=0 ps=0 
M1678 GND d3 diff_282840_108600# GND efet w=16200 l=600
+ ad=0 pd=0 as=1.82592e+07 ps=35520 
M1679 diff_266400_168600# Vdd Vdd GND efet w=660 l=3840
+ ad=0 pd=0 as=0 ps=0 
M1680 diff_268200_169080# diff_268200_169080# diff_268200_169080# GND efet w=180 l=420
+ ad=1.44e+06 pd=5040 as=0 ps=0 
M1681 Vdd Vdd Vdd GND efet w=60 l=120
+ ad=0 pd=0 as=0 ps=0 
M1682 Vdd Vdd Vdd GND efet w=120 l=240
+ ad=0 pd=0 as=0 ps=0 
M1683 diff_268200_169080# diff_268200_169080# diff_268200_169080# GND efet w=120 l=300
+ ad=0 pd=0 as=0 ps=0 
M1684 Vdd Vdd diff_275160_168600# GND efet w=720 l=3240
+ ad=0 pd=0 as=0 ps=0 
M1685 diff_280200_173280# Vdd Vdd GND efet w=600 l=2160
+ ad=0 pd=0 as=0 ps=0 
M1686 diff_264960_142800# Vdd Vdd GND efet w=720 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1687 diff_282840_108600# Vdd Vdd GND efet w=960 l=1560
+ ad=0 pd=0 as=0 ps=0 
M1688 diff_268200_169080# diff_261360_171960# diff_271080_135600# GND efet w=1200 l=720
+ ad=0 pd=0 as=1.58256e+07 ps=36240 
M1689 diff_282840_127320# Vdd Vdd GND efet w=960 l=1560
+ ad=1.20096e+07 pd=19680 as=0 ps=0 
M1690 GND diff_282840_108600# diff_282840_127320# GND efet w=4560 l=600
+ ad=0 pd=0 as=0 ps=0 
M1691 diff_266400_168600# diff_264960_151920# GND GND efet w=1560 l=600
+ ad=0 pd=0 as=0 ps=0 
M1692 sync clk2 diff_276720_158280# GND efet w=1200 l=600
+ ad=0 pd=0 as=1.5264e+06 ps=5280 
M1693 diff_276720_158280# diff_276720_158280# diff_276720_158280# GND efet w=120 l=120
+ ad=0 pd=0 as=0 ps=0 
M1694 diff_276720_158280# diff_276720_158280# diff_276720_158280# GND efet w=60 l=180
+ ad=0 pd=0 as=0 ps=0 
M1695 GND diff_264960_151920# diff_165720_170280# GND efet w=29400 l=600
+ ad=0 pd=0 as=5.22864e+07 ps=106320 
M1696 diff_165720_170280# diff_259200_153240# diff_165720_170280# GND efet w=5520 l=1680
+ ad=0 pd=0 as=0 ps=0 
M1697 diff_165720_170280# diff_259200_153240# Vdd GND efet w=1560 l=600
+ ad=0 pd=0 as=0 ps=0 
M1698 diff_64920_166200# diff_18960_80400# GND GND efet w=18960 l=720
+ ad=0 pd=0 as=0 ps=0 
M1699 GND diff_18960_80400# diff_82080_136560# GND efet w=18960 l=720
+ ad=0 pd=0 as=0 ps=0 
M1700 diff_100800_148560# diff_100440_147960# diff_100800_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1701 diff_102840_148560# diff_100440_147960# diff_102840_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1702 diff_104880_148560# diff_100440_147960# diff_104880_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1703 diff_106920_148560# diff_100440_147960# diff_106920_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1704 diff_108960_148560# diff_100440_147960# diff_108960_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1705 diff_111000_148560# diff_100440_147960# diff_111000_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1706 diff_113040_148560# diff_100440_147960# diff_113040_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1707 diff_115080_148560# diff_100440_147960# diff_115080_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1708 diff_117120_148560# diff_100440_147960# diff_117120_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1709 diff_119160_148560# diff_100440_147960# diff_119160_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1710 diff_121200_148560# diff_100440_147960# diff_121200_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1711 diff_123240_148560# diff_100440_147960# diff_123240_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1712 diff_125280_148560# diff_100440_147960# diff_125280_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1713 diff_127320_148560# diff_100440_147960# diff_127320_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1714 diff_129360_148560# diff_100440_147960# diff_129360_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1715 diff_131400_148560# diff_100440_147960# diff_131400_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1716 diff_133440_148560# diff_100440_147960# diff_133440_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1717 diff_135480_148560# diff_100440_147960# diff_135480_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1718 diff_137520_148560# diff_100440_147960# diff_137520_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1719 diff_139560_148560# diff_100440_147960# diff_139560_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1720 diff_141600_148560# diff_100440_147960# diff_141600_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1721 diff_143640_148560# diff_100440_147960# diff_143640_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1722 diff_145680_148560# diff_100440_147960# diff_145680_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1723 diff_147720_148560# diff_100440_147960# diff_147720_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1724 diff_149760_148560# diff_100440_147960# diff_149760_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1725 diff_151800_148560# diff_100440_147960# diff_151800_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1726 diff_153840_148560# diff_100440_147960# diff_153840_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1727 diff_155880_148560# diff_100440_147960# diff_155880_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1728 diff_157920_148560# diff_100440_147960# diff_157920_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1729 diff_159960_148560# diff_100440_147960# diff_159960_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1730 diff_162000_148560# diff_100440_147960# diff_162000_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1731 diff_164040_148560# diff_100440_147960# diff_164040_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1732 diff_166080_148560# diff_100440_147960# diff_166080_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1733 diff_168120_148560# diff_100440_147960# diff_168120_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1734 diff_170160_148560# diff_100440_147960# diff_170160_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1735 diff_172200_148560# diff_100440_147960# diff_172200_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1736 diff_174240_148560# diff_100440_147960# diff_174240_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1737 diff_176280_148560# diff_100440_147960# diff_176280_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1738 diff_178320_148560# diff_100440_147960# diff_178320_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1739 diff_180360_148560# diff_100440_147960# diff_180360_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1740 diff_182400_148560# diff_100440_147960# diff_182400_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1741 diff_184440_148560# diff_100440_147960# diff_184440_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1742 diff_186480_148560# diff_100440_147960# diff_186480_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1743 diff_188520_148560# diff_100440_147960# diff_188520_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1744 diff_190560_148560# diff_100440_147960# diff_190560_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1745 diff_192600_148560# diff_100440_147960# diff_192600_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1746 diff_194640_148560# diff_100440_147960# diff_194640_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1747 diff_196680_148560# diff_100440_147960# diff_196680_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1748 diff_198720_148560# diff_100440_147960# diff_198720_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1749 diff_200760_148560# diff_100440_147960# diff_200760_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1750 diff_202800_148560# diff_100440_147960# diff_202800_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1751 diff_204840_148560# diff_100440_147960# diff_204840_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1752 diff_206880_148560# diff_100440_147960# diff_206880_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1753 diff_208920_148560# diff_100440_147960# diff_208920_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1754 diff_210960_148560# diff_100440_147960# diff_210960_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1755 diff_213000_148560# diff_100440_147960# diff_213000_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1756 diff_215040_148560# diff_100440_147960# diff_215040_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1757 diff_217080_148560# diff_100440_147960# diff_217080_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1758 diff_219120_148560# diff_100440_147960# diff_219120_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1759 diff_221160_148560# diff_100440_147960# diff_221160_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1760 diff_223200_148560# diff_100440_147960# diff_223200_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1761 diff_225240_148560# diff_100440_147960# diff_225240_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1762 diff_227280_148560# diff_100440_147960# diff_227280_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1763 diff_229320_148560# diff_100440_147960# diff_229320_146400# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1764 diff_100440_150240# Vdd Vdd GND efet w=600 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1765 diff_100800_146400# diff_100440_145800# diff_100800_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1766 diff_102840_146400# diff_100440_145800# diff_102840_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1767 diff_104880_146400# diff_100440_145800# diff_104880_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1768 diff_106920_146400# diff_100440_145800# diff_106920_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1769 diff_108960_146400# diff_100440_145800# diff_108960_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1770 diff_111000_146400# diff_100440_145800# diff_111000_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1771 diff_113040_146400# diff_100440_145800# diff_113040_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1772 diff_115080_146400# diff_100440_145800# diff_115080_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1773 diff_117120_146400# diff_100440_145800# diff_117120_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1774 diff_119160_146400# diff_100440_145800# diff_119160_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1775 diff_121200_146400# diff_100440_145800# diff_121200_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1776 diff_123240_146400# diff_100440_145800# diff_123240_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1777 diff_125280_146400# diff_100440_145800# diff_125280_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1778 diff_127320_146400# diff_100440_145800# diff_127320_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1779 diff_129360_146400# diff_100440_145800# diff_129360_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1780 diff_131400_146400# diff_100440_145800# diff_131400_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1781 diff_133440_146400# diff_100440_145800# diff_133440_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1782 diff_135480_146400# diff_100440_145800# diff_135480_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1783 diff_137520_146400# diff_100440_145800# diff_137520_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1784 diff_139560_146400# diff_100440_145800# diff_139560_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1785 diff_141600_146400# diff_100440_145800# diff_141600_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1786 diff_143640_146400# diff_100440_145800# diff_143640_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1787 diff_145680_146400# diff_100440_145800# diff_145680_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1788 diff_147720_146400# diff_100440_145800# diff_147720_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1789 diff_149760_146400# diff_100440_145800# diff_149760_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1790 diff_151800_146400# diff_100440_145800# diff_151800_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1791 diff_153840_146400# diff_100440_145800# diff_153840_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1792 diff_155880_146400# diff_100440_145800# diff_155880_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1793 diff_157920_146400# diff_100440_145800# diff_157920_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1794 diff_159960_146400# diff_100440_145800# diff_159960_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1795 diff_162000_146400# diff_100440_145800# diff_162000_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1796 diff_164040_146400# diff_100440_145800# diff_164040_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1797 diff_166080_146400# diff_100440_145800# diff_166080_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1798 diff_168120_146400# diff_100440_145800# diff_168120_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1799 diff_170160_146400# diff_100440_145800# diff_170160_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1800 diff_172200_146400# diff_100440_145800# diff_172200_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1801 diff_174240_146400# diff_100440_145800# diff_174240_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1802 diff_176280_146400# diff_100440_145800# diff_176280_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1803 diff_178320_146400# diff_100440_145800# diff_178320_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1804 diff_180360_146400# diff_100440_145800# diff_180360_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1805 diff_182400_146400# diff_100440_145800# diff_182400_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1806 diff_184440_146400# diff_100440_145800# diff_184440_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1807 diff_186480_146400# diff_100440_145800# diff_186480_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1808 diff_188520_146400# diff_100440_145800# diff_188520_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1809 diff_190560_146400# diff_100440_145800# diff_190560_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1810 diff_192600_146400# diff_100440_145800# diff_192600_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1811 diff_194640_146400# diff_100440_145800# diff_194640_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1812 diff_196680_146400# diff_100440_145800# diff_196680_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1813 diff_198720_146400# diff_100440_145800# diff_198720_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1814 diff_200760_146400# diff_100440_145800# diff_200760_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1815 diff_202800_146400# diff_100440_145800# diff_202800_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1816 diff_204840_146400# diff_100440_145800# diff_204840_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1817 diff_206880_146400# diff_100440_145800# diff_206880_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1818 diff_208920_146400# diff_100440_145800# diff_208920_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1819 diff_210960_146400# diff_100440_145800# diff_210960_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1820 diff_213000_146400# diff_100440_145800# diff_213000_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1821 diff_215040_146400# diff_100440_145800# diff_215040_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1822 diff_217080_146400# diff_100440_145800# diff_217080_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1823 diff_219120_146400# diff_100440_145800# diff_219120_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1824 diff_221160_146400# diff_100440_145800# diff_221160_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1825 diff_223200_146400# diff_100440_145800# diff_223200_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1826 diff_225240_146400# diff_100440_145800# diff_225240_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1827 diff_227280_146400# diff_100440_145800# diff_227280_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1828 diff_229320_146400# diff_100440_145800# diff_229320_144120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1829 Vdd Vdd diff_100440_143520# GND efet w=600 l=1320
+ ad=0 pd=0 as=8.5104e+06 ps=25920 
M1830 diff_100800_144120# diff_100440_143520# diff_100800_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1831 diff_102840_144120# diff_100440_143520# diff_102840_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1832 diff_104880_144120# diff_100440_143520# diff_104880_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1833 diff_106920_144120# diff_100440_143520# diff_106920_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1834 diff_108960_144120# diff_100440_143520# diff_108960_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1835 diff_111000_144120# diff_100440_143520# diff_111000_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1836 diff_113040_144120# diff_100440_143520# diff_113040_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1837 diff_115080_144120# diff_100440_143520# diff_115080_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1838 diff_117120_144120# diff_100440_143520# diff_117120_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1839 diff_119160_144120# diff_100440_143520# diff_119160_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1840 diff_121200_144120# diff_100440_143520# diff_121200_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1841 diff_123240_144120# diff_100440_143520# diff_123240_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1842 diff_125280_144120# diff_100440_143520# diff_125280_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1843 diff_127320_144120# diff_100440_143520# diff_127320_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1844 diff_129360_144120# diff_100440_143520# diff_129360_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1845 diff_131400_144120# diff_100440_143520# diff_131400_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1846 diff_133440_144120# diff_100440_143520# diff_133440_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1847 diff_135480_144120# diff_100440_143520# diff_135480_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1848 diff_137520_144120# diff_100440_143520# diff_137520_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1849 diff_139560_144120# diff_100440_143520# diff_139560_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1850 diff_141600_144120# diff_100440_143520# diff_141600_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1851 diff_143640_144120# diff_100440_143520# diff_143640_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1852 diff_145680_144120# diff_100440_143520# diff_145680_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1853 diff_147720_144120# diff_100440_143520# diff_147720_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1854 diff_149760_144120# diff_100440_143520# diff_149760_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1855 diff_151800_144120# diff_100440_143520# diff_151800_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1856 diff_153840_144120# diff_100440_143520# diff_153840_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1857 diff_155880_144120# diff_100440_143520# diff_155880_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1858 diff_157920_144120# diff_100440_143520# diff_157920_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1859 diff_159960_144120# diff_100440_143520# diff_159960_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1860 diff_162000_144120# diff_100440_143520# diff_162000_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1861 diff_164040_144120# diff_100440_143520# diff_164040_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1862 diff_166080_144120# diff_100440_143520# diff_166080_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1863 diff_168120_144120# diff_100440_143520# diff_168120_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1864 diff_170160_144120# diff_100440_143520# diff_170160_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1865 diff_172200_144120# diff_100440_143520# diff_172200_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1866 diff_174240_144120# diff_100440_143520# diff_174240_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1867 diff_176280_144120# diff_100440_143520# diff_176280_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1868 diff_178320_144120# diff_100440_143520# diff_178320_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1869 diff_180360_144120# diff_100440_143520# diff_180360_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1870 diff_182400_144120# diff_100440_143520# diff_182400_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1871 diff_184440_144120# diff_100440_143520# diff_184440_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1872 diff_186480_144120# diff_100440_143520# diff_186480_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1873 diff_188520_144120# diff_100440_143520# diff_188520_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1874 diff_190560_144120# diff_100440_143520# diff_190560_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1875 diff_192600_144120# diff_100440_143520# diff_192600_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1876 diff_194640_144120# diff_100440_143520# diff_194640_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1877 diff_196680_144120# diff_100440_143520# diff_196680_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1878 diff_198720_144120# diff_100440_143520# diff_198720_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1879 diff_200760_144120# diff_100440_143520# diff_200760_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1880 diff_202800_144120# diff_100440_143520# diff_202800_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1881 diff_204840_144120# diff_100440_143520# diff_204840_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1882 diff_206880_144120# diff_100440_143520# diff_206880_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1883 diff_208920_144120# diff_100440_143520# diff_208920_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1884 diff_210960_144120# diff_100440_143520# diff_210960_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1885 diff_213000_144120# diff_100440_143520# diff_213000_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1886 diff_215040_144120# diff_100440_143520# diff_215040_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1887 diff_217080_144120# diff_100440_143520# diff_217080_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1888 diff_219120_144120# diff_100440_143520# diff_219120_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1889 diff_221160_144120# diff_100440_143520# diff_221160_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1890 diff_223200_144120# diff_100440_143520# diff_223200_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1891 diff_225240_144120# diff_100440_143520# diff_225240_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1892 diff_227280_144120# diff_100440_143520# diff_227280_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1893 diff_229320_144120# diff_100440_143520# diff_229320_141960# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1894 diff_80400_166200# diff_18960_80400# GND GND efet w=19080 l=720
+ ad=0 pd=0 as=0 ps=0 
M1895 diff_100440_143520# diff_238440_42720# diff_236760_149400# GND efet w=7440 l=600
+ ad=0 pd=0 as=0 ps=0 
M1896 diff_236760_149400# diff_241320_99600# diff_100440_147960# GND efet w=8400 l=600
+ ad=0 pd=0 as=1.15488e+07 ps=22800 
M1897 diff_100440_147960# Vdd Vdd GND efet w=720 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1898 Vdd Vdd diff_100440_145800# GND efet w=720 l=1200
+ ad=0 pd=0 as=9.4176e+06 ps=24720 
M1899 diff_100800_141960# diff_100440_141360# diff_100800_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1900 diff_102840_141960# diff_100440_141360# diff_102840_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1901 diff_104880_141960# diff_100440_141360# diff_104880_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1902 diff_106920_141960# diff_100440_141360# diff_106920_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1903 diff_108960_141960# diff_100440_141360# diff_108960_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1904 diff_111000_141960# diff_100440_141360# diff_111000_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1905 diff_113040_141960# diff_100440_141360# diff_113040_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1906 diff_115080_141960# diff_100440_141360# diff_115080_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1907 diff_117120_141960# diff_100440_141360# diff_117120_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1908 diff_119160_141960# diff_100440_141360# diff_119160_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1909 diff_121200_141960# diff_100440_141360# diff_121200_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1910 diff_123240_141960# diff_100440_141360# diff_123240_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1911 diff_125280_141960# diff_100440_141360# diff_125280_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1912 diff_127320_141960# diff_100440_141360# diff_127320_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1913 diff_129360_141960# diff_100440_141360# diff_129360_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1914 diff_131400_141960# diff_100440_141360# diff_131400_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1915 diff_133440_141960# diff_100440_141360# diff_133440_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1916 diff_135480_141960# diff_100440_141360# diff_135480_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1917 diff_137520_141960# diff_100440_141360# diff_137520_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1918 diff_139560_141960# diff_100440_141360# diff_139560_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1919 diff_141600_141960# diff_100440_141360# diff_141600_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1920 diff_143640_141960# diff_100440_141360# diff_143640_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1921 diff_145680_141960# diff_100440_141360# diff_145680_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1922 diff_147720_141960# diff_100440_141360# diff_147720_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1923 diff_149760_141960# diff_100440_141360# diff_149760_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1924 diff_151800_141960# diff_100440_141360# diff_151800_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1925 diff_153840_141960# diff_100440_141360# diff_153840_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1926 diff_155880_141960# diff_100440_141360# diff_155880_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1927 diff_157920_141960# diff_100440_141360# diff_157920_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1928 diff_159960_141960# diff_100440_141360# diff_159960_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1929 diff_162000_141960# diff_100440_141360# diff_162000_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1930 diff_164040_141960# diff_100440_141360# diff_164040_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1931 diff_166080_141960# diff_100440_141360# diff_166080_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1932 diff_168120_141960# diff_100440_141360# diff_168120_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1933 diff_170160_141960# diff_100440_141360# diff_170160_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1934 diff_172200_141960# diff_100440_141360# diff_172200_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1935 diff_174240_141960# diff_100440_141360# diff_174240_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1936 diff_176280_141960# diff_100440_141360# diff_176280_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1937 diff_178320_141960# diff_100440_141360# diff_178320_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1938 diff_180360_141960# diff_100440_141360# diff_180360_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1939 diff_182400_141960# diff_100440_141360# diff_182400_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1940 diff_184440_141960# diff_100440_141360# diff_184440_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1941 diff_186480_141960# diff_100440_141360# diff_186480_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1942 diff_188520_141960# diff_100440_141360# diff_188520_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1943 diff_190560_141960# diff_100440_141360# diff_190560_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1944 diff_192600_141960# diff_100440_141360# diff_192600_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1945 diff_194640_141960# diff_100440_141360# diff_194640_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1946 diff_196680_141960# diff_100440_141360# diff_196680_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1947 diff_198720_141960# diff_100440_141360# diff_198720_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1948 diff_200760_141960# diff_100440_141360# diff_200760_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1949 diff_202800_141960# diff_100440_141360# diff_202800_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1950 diff_204840_141960# diff_100440_141360# diff_204840_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1951 diff_206880_141960# diff_100440_141360# diff_206880_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1952 diff_208920_141960# diff_100440_141360# diff_208920_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1953 diff_210960_141960# diff_100440_141360# diff_210960_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1954 diff_213000_141960# diff_100440_141360# diff_213000_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1955 diff_215040_141960# diff_100440_141360# diff_215040_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1956 diff_217080_141960# diff_100440_141360# diff_217080_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1957 diff_219120_141960# diff_100440_141360# diff_219120_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1958 diff_221160_141960# diff_100440_141360# diff_221160_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1959 diff_223200_141960# diff_100440_141360# diff_223200_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1960 diff_225240_141960# diff_100440_141360# diff_225240_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1961 diff_227280_141960# diff_100440_141360# diff_227280_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1962 diff_229320_141960# diff_100440_141360# diff_229320_139680# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M1963 diff_236760_140760# diff_236160_42720# diff_100440_141360# GND efet w=8640 l=600
+ ad=3.82608e+07 pd=72960 as=9.6768e+06 ps=23040 
M1964 diff_100440_145800# diff_243120_97920# diff_236760_149400# GND efet w=7920 l=600
+ ad=0 pd=0 as=0 ps=0 
M1965 diff_100800_139680# diff_100440_139080# diff_100800_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1966 diff_102840_139680# diff_100440_139080# diff_102840_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1967 diff_104880_139680# diff_100440_139080# diff_104880_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1968 diff_106920_139680# diff_100440_139080# diff_106920_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1969 diff_108960_139680# diff_100440_139080# diff_108960_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1970 diff_111000_139680# diff_100440_139080# diff_111000_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1971 diff_113040_139680# diff_100440_139080# diff_113040_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1972 diff_115080_139680# diff_100440_139080# diff_115080_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1973 diff_117120_139680# diff_100440_139080# diff_117120_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1974 diff_119160_139680# diff_100440_139080# diff_119160_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1975 diff_121200_139680# diff_100440_139080# diff_121200_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1976 diff_123240_139680# diff_100440_139080# diff_123240_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1977 diff_125280_139680# diff_100440_139080# diff_125280_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1978 diff_127320_139680# diff_100440_139080# diff_127320_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1979 diff_129360_139680# diff_100440_139080# diff_129360_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1980 diff_131400_139680# diff_100440_139080# diff_131400_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1981 diff_133440_139680# diff_100440_139080# diff_133440_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1982 diff_135480_139680# diff_100440_139080# diff_135480_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1983 diff_137520_139680# diff_100440_139080# diff_137520_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1984 diff_139560_139680# diff_100440_139080# diff_139560_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1985 diff_141600_139680# diff_100440_139080# diff_141600_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1986 diff_143640_139680# diff_100440_139080# diff_143640_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1987 diff_145680_139680# diff_100440_139080# diff_145680_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1988 diff_147720_139680# diff_100440_139080# diff_147720_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1989 diff_149760_139680# diff_100440_139080# diff_149760_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1990 diff_151800_139680# diff_100440_139080# diff_151800_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1991 diff_153840_139680# diff_100440_139080# diff_153840_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1992 diff_155880_139680# diff_100440_139080# diff_155880_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1993 diff_157920_139680# diff_100440_139080# diff_157920_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1994 diff_159960_139680# diff_100440_139080# diff_159960_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1995 diff_162000_139680# diff_100440_139080# diff_162000_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1996 diff_164040_139680# diff_100440_139080# diff_164040_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1997 diff_166080_139680# diff_100440_139080# diff_166080_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1998 diff_168120_139680# diff_100440_139080# diff_168120_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M1999 diff_170160_139680# diff_100440_139080# diff_170160_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2000 diff_172200_139680# diff_100440_139080# diff_172200_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2001 diff_174240_139680# diff_100440_139080# diff_174240_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2002 diff_176280_139680# diff_100440_139080# diff_176280_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2003 diff_178320_139680# diff_100440_139080# diff_178320_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2004 diff_180360_139680# diff_100440_139080# diff_180360_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2005 diff_182400_139680# diff_100440_139080# diff_182400_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2006 diff_184440_139680# diff_100440_139080# diff_184440_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2007 diff_186480_139680# diff_100440_139080# diff_186480_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2008 diff_188520_139680# diff_100440_139080# diff_188520_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2009 diff_190560_139680# diff_100440_139080# diff_190560_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2010 diff_192600_139680# diff_100440_139080# diff_192600_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2011 diff_194640_139680# diff_100440_139080# diff_194640_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2012 diff_196680_139680# diff_100440_139080# diff_196680_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2013 diff_198720_139680# diff_100440_139080# diff_198720_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2014 diff_200760_139680# diff_100440_139080# diff_200760_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2015 diff_202800_139680# diff_100440_139080# diff_202800_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2016 diff_204840_139680# diff_100440_139080# diff_204840_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2017 diff_206880_139680# diff_100440_139080# diff_206880_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2018 diff_208920_139680# diff_100440_139080# diff_208920_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2019 diff_210960_139680# diff_100440_139080# diff_210960_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2020 diff_213000_139680# diff_100440_139080# diff_213000_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2021 diff_215040_139680# diff_100440_139080# diff_215040_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2022 diff_217080_139680# diff_100440_139080# diff_217080_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2023 diff_219120_139680# diff_100440_139080# diff_219120_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2024 diff_221160_139680# diff_100440_139080# diff_221160_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2025 diff_223200_139680# diff_100440_139080# diff_223200_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2026 diff_225240_139680# diff_100440_139080# diff_225240_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2027 diff_227280_139680# diff_100440_139080# diff_227280_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2028 diff_229320_139680# diff_100440_139080# diff_229320_137520# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2029 diff_100440_141360# Vdd Vdd GND efet w=600 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2030 diff_100800_137520# diff_100440_136920# diff_100800_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2031 diff_102840_137520# diff_100440_136920# diff_102840_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2032 diff_104880_137520# diff_100440_136920# diff_104880_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2033 diff_106920_137520# diff_100440_136920# diff_106920_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2034 diff_108960_137520# diff_100440_136920# diff_108960_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2035 diff_111000_137520# diff_100440_136920# diff_111000_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2036 diff_113040_137520# diff_100440_136920# diff_113040_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2037 diff_115080_137520# diff_100440_136920# diff_115080_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2038 diff_117120_137520# diff_100440_136920# diff_117120_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2039 diff_119160_137520# diff_100440_136920# diff_119160_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2040 diff_121200_137520# diff_100440_136920# diff_121200_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2041 diff_123240_137520# diff_100440_136920# diff_123240_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2042 diff_125280_137520# diff_100440_136920# diff_125280_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2043 diff_127320_137520# diff_100440_136920# diff_127320_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2044 diff_129360_137520# diff_100440_136920# diff_129360_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2045 diff_131400_137520# diff_100440_136920# diff_131400_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2046 diff_133440_137520# diff_100440_136920# diff_133440_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2047 diff_135480_137520# diff_100440_136920# diff_135480_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2048 diff_137520_137520# diff_100440_136920# diff_137520_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2049 diff_139560_137520# diff_100440_136920# diff_139560_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2050 diff_141600_137520# diff_100440_136920# diff_141600_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2051 diff_143640_137520# diff_100440_136920# diff_143640_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2052 diff_145680_137520# diff_100440_136920# diff_145680_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2053 diff_147720_137520# diff_100440_136920# diff_147720_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2054 diff_149760_137520# diff_100440_136920# diff_149760_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2055 diff_151800_137520# diff_100440_136920# diff_151800_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2056 diff_153840_137520# diff_100440_136920# diff_153840_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2057 diff_155880_137520# diff_100440_136920# diff_155880_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2058 diff_157920_137520# diff_100440_136920# diff_157920_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2059 diff_159960_137520# diff_100440_136920# diff_159960_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2060 diff_162000_137520# diff_100440_136920# diff_162000_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2061 diff_164040_137520# diff_100440_136920# diff_164040_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2062 diff_166080_137520# diff_100440_136920# diff_166080_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2063 diff_168120_137520# diff_100440_136920# diff_168120_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2064 diff_170160_137520# diff_100440_136920# diff_170160_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2065 diff_172200_137520# diff_100440_136920# diff_172200_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2066 diff_174240_137520# diff_100440_136920# diff_174240_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2067 diff_176280_137520# diff_100440_136920# diff_176280_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2068 diff_178320_137520# diff_100440_136920# diff_178320_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2069 diff_180360_137520# diff_100440_136920# diff_180360_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2070 diff_182400_137520# diff_100440_136920# diff_182400_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2071 diff_184440_137520# diff_100440_136920# diff_184440_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2072 diff_186480_137520# diff_100440_136920# diff_186480_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2073 diff_188520_137520# diff_100440_136920# diff_188520_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2074 diff_190560_137520# diff_100440_136920# diff_190560_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2075 diff_192600_137520# diff_100440_136920# diff_192600_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2076 diff_194640_137520# diff_100440_136920# diff_194640_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2077 diff_196680_137520# diff_100440_136920# diff_196680_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2078 diff_198720_137520# diff_100440_136920# diff_198720_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2079 diff_200760_137520# diff_100440_136920# diff_200760_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2080 diff_202800_137520# diff_100440_136920# diff_202800_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2081 diff_204840_137520# diff_100440_136920# diff_204840_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2082 diff_206880_137520# diff_100440_136920# diff_206880_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2083 diff_208920_137520# diff_100440_136920# diff_208920_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2084 diff_210960_137520# diff_100440_136920# diff_210960_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2085 diff_213000_137520# diff_100440_136920# diff_213000_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2086 diff_215040_137520# diff_100440_136920# diff_215040_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2087 diff_217080_137520# diff_100440_136920# diff_217080_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2088 diff_219120_137520# diff_100440_136920# diff_219120_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2089 diff_221160_137520# diff_100440_136920# diff_221160_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2090 diff_223200_137520# diff_100440_136920# diff_223200_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2091 diff_225240_137520# diff_100440_136920# diff_225240_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2092 diff_227280_137520# diff_100440_136920# diff_227280_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2093 diff_229320_137520# diff_100440_136920# diff_229320_135240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2094 d3 clk2 diff_33360_134640# GND efet w=1200 l=720
+ ad=0 pd=0 as=1.008e+06 ps=4080 
M2095 d2 clk2 diff_48840_134640# GND efet w=1200 l=720
+ ad=0 pd=0 as=1.008e+06 ps=4080 
M2096 d1 clk2 diff_64440_134640# GND efet w=1200 l=720
+ ad=0 pd=0 as=1.008e+06 ps=4080 
M2097 d0 clk2 diff_79920_134640# GND efet w=1200 l=720
+ ad=0 pd=0 as=1.008e+06 ps=4080 
M2098 Vdd Vdd diff_100440_134640# GND efet w=600 l=1320
+ ad=0 pd=0 as=8.5104e+06 ps=25920 
M2099 diff_33360_134640# diff_15480_82200# diff_33360_127800# GND efet w=1200 l=720
+ ad=0 pd=0 as=1.64736e+07 ps=35520 
M2100 diff_48840_134640# diff_15480_82200# diff_48840_127680# GND efet w=1200 l=720
+ ad=0 pd=0 as=1.61136e+07 ps=35280 
M2101 diff_64440_134640# diff_15480_82200# diff_64440_127680# GND efet w=1200 l=720
+ ad=0 pd=0 as=1.66896e+07 ps=35280 
M2102 diff_79920_134640# diff_15480_82200# diff_79920_127680# GND efet w=1200 l=720
+ ad=0 pd=0 as=1.65888e+07 ps=35760 
M2103 diff_100800_135240# diff_100440_134640# diff_100800_132000# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2104 diff_102840_135240# diff_100440_134640# diff_102480_126360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2105 diff_104880_135240# diff_100440_134640# diff_104880_132240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2106 diff_106920_135240# diff_100440_134640# diff_106920_128160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2107 diff_108960_135240# diff_100440_134640# diff_108960_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2108 diff_111000_135240# diff_100440_134640# diff_111000_126240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2109 diff_113040_135240# diff_100440_134640# diff_113040_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2110 diff_115080_135240# diff_100440_134640# diff_115080_128160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2111 diff_117120_135240# diff_100440_134640# diff_117120_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2112 diff_119160_135240# diff_100440_134640# diff_119160_126240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2113 diff_121200_135240# diff_100440_134640# diff_121200_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2114 diff_123240_135240# diff_100440_134640# diff_123240_128160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2115 diff_125280_135240# diff_100440_134640# diff_125280_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2116 diff_127320_135240# diff_100440_134640# diff_127320_126240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2117 diff_129360_135240# diff_100440_134640# diff_129360_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2118 diff_131400_135240# diff_100440_134640# diff_131400_128160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2119 diff_133440_135240# diff_100440_134640# diff_133440_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2120 diff_135480_135240# diff_100440_134640# diff_135480_126240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2121 diff_137520_135240# diff_100440_134640# diff_137520_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2122 diff_139560_135240# diff_100440_134640# diff_139560_128160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2123 diff_141600_135240# diff_100440_134640# diff_141600_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2124 diff_143640_135240# diff_100440_134640# diff_143640_126240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2125 diff_145680_135240# diff_100440_134640# diff_145680_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2126 diff_147720_135240# diff_100440_134640# diff_147720_128160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2127 diff_149760_135240# diff_100440_134640# diff_149760_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2128 diff_151800_135240# diff_100440_134640# diff_151800_126240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2129 diff_153840_135240# diff_100440_134640# diff_153840_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2130 diff_155880_135240# diff_100440_134640# diff_155880_128160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2131 diff_157920_135240# diff_100440_134640# diff_157920_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2132 diff_159960_135240# diff_100440_134640# diff_159960_126240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2133 diff_162000_135240# diff_100440_134640# diff_162000_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2134 diff_164040_135240# diff_100440_134640# diff_164040_128160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2135 diff_166080_135240# diff_100440_134640# diff_166080_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2136 diff_168120_135240# diff_100440_134640# diff_168120_126240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2137 diff_170160_135240# diff_100440_134640# diff_170160_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2138 diff_172200_135240# diff_100440_134640# diff_172200_128160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2139 diff_174240_135240# diff_100440_134640# diff_174240_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2140 diff_176280_135240# diff_100440_134640# diff_176280_126240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2141 diff_178320_135240# diff_100440_134640# diff_178320_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2142 diff_180360_135240# diff_100440_134640# diff_180360_128160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2143 diff_182400_135240# diff_100440_134640# diff_182400_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2144 diff_184440_135240# diff_100440_134640# diff_184440_126240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2145 diff_186480_135240# diff_100440_134640# diff_186480_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2146 diff_188520_135240# diff_100440_134640# diff_188520_128160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2147 diff_190560_135240# diff_100440_134640# diff_190560_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2148 diff_192600_135240# diff_100440_134640# diff_192600_126240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2149 diff_194640_135240# diff_100440_134640# diff_194640_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2150 diff_196680_135240# diff_100440_134640# diff_196680_128160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2151 diff_198720_135240# diff_100440_134640# diff_198720_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2152 diff_200760_135240# diff_100440_134640# diff_200760_126240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2153 diff_202800_135240# diff_100440_134640# diff_202800_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2154 diff_204840_135240# diff_100440_134640# diff_204840_128160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2155 diff_206880_135240# diff_100440_134640# diff_206880_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2156 diff_208920_135240# diff_100440_134640# diff_208920_126240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2157 diff_210960_135240# diff_100440_134640# diff_210960_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2158 diff_213000_135240# diff_100440_134640# diff_213000_128160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2159 diff_215040_135240# diff_100440_134640# diff_215040_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2160 diff_217080_135240# diff_100440_134640# diff_217080_126240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2161 diff_219120_135240# diff_100440_134640# diff_219120_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2162 diff_221160_135240# diff_100440_134640# diff_221160_128160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2163 diff_223200_135240# diff_100440_134640# diff_223200_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2164 diff_225240_135240# diff_100440_134640# diff_225240_126240# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2165 diff_227280_135240# diff_100440_134640# diff_227280_132120# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2166 diff_229320_135240# diff_100440_134640# diff_229320_128160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M2167 diff_28080_131640# diff_15480_82200# GND GND efet w=1800 l=720
+ ad=2.5776e+06 pd=7200 as=0 ps=0 
M2168 diff_33360_127800# diff_33360_127800# diff_33360_127800# GND efet w=360 l=360
+ ad=0 pd=0 as=0 ps=0 
M2169 Vdd Vdd diff_28080_131640# GND efet w=420 l=4140
+ ad=0 pd=0 as=0 ps=0 
M2170 GND GND sync GND efet w=11580 l=780
+ ad=0 pd=0 as=0 ps=0 
M2171 diff_33600_117000# diff_33360_127800# GND GND efet w=7680 l=720
+ ad=7.5168e+06 pd=22080 as=0 ps=0 
M2172 diff_48840_127680# diff_48840_127680# diff_48840_127680# GND efet w=360 l=360
+ ad=0 pd=0 as=0 ps=0 
M2173 diff_33360_127800# diff_33360_127800# diff_33360_127800# GND efet w=240 l=240
+ ad=0 pd=0 as=0 ps=0 
M2174 GND diff_33600_117000# diff_35520_129960# GND efet w=5040 l=600
+ ad=0 pd=0 as=1.3752e+07 ps=34560 
M2175 diff_35520_129960# diff_28080_131640# diff_33360_127800# GND efet w=1200 l=720
+ ad=0 pd=0 as=0 ps=0 
M2176 diff_49200_117000# diff_48840_127680# GND GND efet w=7680 l=720
+ ad=7.4448e+06 pd=22080 as=0 ps=0 
M2177 diff_64440_127680# diff_64440_127680# diff_64440_127680# GND efet w=240 l=240
+ ad=0 pd=0 as=0 ps=0 
M2178 diff_48840_127680# diff_48840_127680# diff_48840_127680# GND efet w=240 l=240
+ ad=0 pd=0 as=0 ps=0 
M2179 GND diff_49200_117000# diff_50880_129960# GND efet w=5040 l=600
+ ad=0 pd=0 as=1.37664e+07 ps=34320 
M2180 diff_50880_129960# diff_28080_131640# diff_48840_127680# GND efet w=1200 l=720
+ ad=0 pd=0 as=0 ps=0 
M2181 diff_64680_117000# diff_64440_127680# GND GND efet w=7560 l=720
+ ad=7.9488e+06 pd=21840 as=0 ps=0 
M2182 diff_100440_134640# diff_238440_42720# diff_236760_140760# GND efet w=7440 l=600
+ ad=0 pd=0 as=0 ps=0 
M2183 diff_236760_140760# diff_241320_99600# diff_100440_139080# GND efet w=8520 l=600
+ ad=0 pd=0 as=1.14768e+07 ps=22800 
M2184 diff_100440_139080# Vdd Vdd GND efet w=720 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2185 Vdd Vdd diff_100440_136920# GND efet w=720 l=1320
+ ad=0 pd=0 as=9.4176e+06 ps=24720 
M2186 diff_79920_127680# diff_79920_127680# diff_79920_127680# GND efet w=360 l=360
+ ad=0 pd=0 as=0 ps=0 
M2187 diff_64440_127680# diff_64440_127680# diff_64440_127680# GND efet w=120 l=120
+ ad=0 pd=0 as=0 ps=0 
M2188 GND diff_64680_117000# diff_66600_129960# GND efet w=5040 l=720
+ ad=0 pd=0 as=1.34208e+07 ps=34080 
M2189 diff_66600_129960# diff_28080_131640# diff_64440_127680# GND efet w=1200 l=720
+ ad=0 pd=0 as=0 ps=0 
M2190 diff_80160_117000# diff_79920_127680# GND GND efet w=7680 l=720
+ ad=7.4448e+06 pd=21840 as=0 ps=0 
M2191 diff_79920_127680# diff_79920_127680# diff_79920_127680# GND efet w=240 l=240
+ ad=0 pd=0 as=0 ps=0 
M2192 GND diff_80160_117000# diff_82080_129960# GND efet w=5040 l=600
+ ad=0 pd=0 as=1.368e+07 ps=34320 
M2193 diff_82080_129960# diff_28080_131640# diff_79920_127680# GND efet w=1200 l=720
+ ad=0 pd=0 as=0 ps=0 
M2194 diff_33360_127800# cl GND GND efet w=3600 l=720
+ ad=0 pd=0 as=0 ps=0 
M2195 GND cl diff_33360_127800# GND efet w=3600 l=840
+ ad=0 pd=0 as=0 ps=0 
M2196 diff_33360_127800# diff_26040_78600# GND GND efet w=4740 l=780
+ ad=0 pd=0 as=0 ps=0 
M2197 diff_33600_117000# Vdd Vdd GND efet w=600 l=1560
+ ad=0 pd=0 as=0 ps=0 
M2198 diff_35520_129960# Vdd Vdd GND efet w=600 l=1440
+ ad=0 pd=0 as=0 ps=0 
M2199 Vdd Vdd Vdd GND efet w=240 l=240
+ ad=0 pd=0 as=0 ps=0 
M2200 Vdd Vdd Vdd GND efet w=180 l=240
+ ad=0 pd=0 as=0 ps=0 
M2201 diff_48840_127680# cl GND GND efet w=3600 l=720
+ ad=0 pd=0 as=0 ps=0 
M2202 GND cl diff_48840_127680# GND efet w=3600 l=840
+ ad=0 pd=0 as=0 ps=0 
M2203 GND diff_100800_132000# diff_99720_123600# GND efet w=2880 l=600
+ ad=0 pd=0 as=7.92e+06 ps=19440 
M2204 diff_103320_126720# diff_102480_126360# GND GND efet w=4620 l=720
+ ad=3.6864e+06 pd=10560 as=0 ps=0 
M2205 GND diff_104880_132240# diff_103680_120240# GND efet w=3960 l=600
+ ad=0 pd=0 as=7.5456e+06 ps=19200 
M2206 diff_107520_128400# diff_106920_128160# GND GND efet w=3960 l=600
+ ad=6.408e+06 pd=18720 as=0 ps=0 
M2207 GND diff_108960_132120# diff_107400_118080# GND efet w=3540 l=720
+ ad=0 pd=0 as=6.6816e+06 ps=17520 
M2208 GND diff_113040_132120# diff_111600_120120# GND efet w=3960 l=600
+ ad=0 pd=0 as=7.5888e+06 ps=19680 
M2209 diff_115680_128400# diff_115080_128160# GND GND efet w=3960 l=600
+ ad=6.6096e+06 pd=18720 as=0 ps=0 
M2210 diff_111600_126600# diff_111000_126240# GND GND efet w=3540 l=660
+ ad=3.2976e+06 pd=9360 as=0 ps=0 
M2211 GND diff_117120_132120# diff_115560_118080# GND efet w=3540 l=720
+ ad=0 pd=0 as=6.7392e+06 ps=17520 
M2212 GND diff_121200_132120# diff_119760_120240# GND efet w=3960 l=600
+ ad=0 pd=0 as=7.7616e+06 ps=19680 
M2213 diff_123840_128400# diff_123240_128160# GND GND efet w=3960 l=600
+ ad=6.552e+06 pd=18720 as=0 ps=0 
M2214 diff_119760_126600# diff_119160_126240# GND GND efet w=3540 l=660
+ ad=3.2976e+06 pd=9360 as=0 ps=0 
M2215 GND diff_125280_132120# diff_123600_118080# GND efet w=3540 l=720
+ ad=0 pd=0 as=7.056e+06 ps=17760 
M2216 GND diff_129360_132120# diff_127800_120240# GND efet w=3960 l=600
+ ad=0 pd=0 as=7.9488e+06 ps=19680 
M2217 diff_132000_128400# diff_131400_128160# GND GND efet w=3960 l=600
+ ad=6.8688e+06 pd=18960 as=0 ps=0 
M2218 diff_127920_126600# diff_127320_126240# GND GND efet w=3540 l=660
+ ad=3.2976e+06 pd=9360 as=0 ps=0 
M2219 GND diff_133440_132120# diff_131760_118080# GND efet w=3540 l=720
+ ad=0 pd=0 as=7.1136e+06 ps=17760 
M2220 GND diff_137520_132120# diff_135960_120120# GND efet w=3960 l=600
+ ad=0 pd=0 as=8.1504e+06 ps=20160 
M2221 diff_140160_128400# diff_139560_128160# GND GND efet w=3960 l=600
+ ad=5.9616e+06 pd=18480 as=0 ps=0 
M2222 diff_136080_126600# diff_135480_126240# GND GND efet w=3540 l=660
+ ad=3.2976e+06 pd=9360 as=0 ps=0 
M2223 GND diff_141600_132120# diff_140040_118080# GND efet w=3540 l=720
+ ad=0 pd=0 as=6.3072e+06 ps=17280 
M2224 GND diff_145680_132120# diff_144240_120240# GND efet w=3960 l=600
+ ad=0 pd=0 as=7.2e+06 ps=19200 
M2225 diff_148320_128400# diff_147720_128160# GND GND efet w=3960 l=600
+ ad=6.2064e+06 pd=18480 as=0 ps=0 
M2226 diff_144240_126600# diff_143640_126240# GND GND efet w=3540 l=660
+ ad=3.2976e+06 pd=9360 as=0 ps=0 
M2227 GND diff_149760_132120# diff_148200_118080# GND efet w=3540 l=720
+ ad=0 pd=0 as=6.3648e+06 ps=17280 
M2228 GND diff_153840_132120# diff_152400_120240# GND efet w=3960 l=600
+ ad=0 pd=0 as=7.3872e+06 ps=19440 
M2229 diff_156480_128400# diff_155880_128160# GND GND efet w=3960 l=600
+ ad=5.9616e+06 pd=18480 as=0 ps=0 
M2230 diff_152400_126600# diff_151800_126240# GND GND efet w=3540 l=660
+ ad=3.2976e+06 pd=9360 as=0 ps=0 
M2231 GND diff_157920_132120# diff_156360_118080# GND efet w=3540 l=720
+ ad=0 pd=0 as=6.3072e+06 ps=17280 
M2232 GND diff_162000_132120# diff_160560_120240# GND efet w=3960 l=600
+ ad=0 pd=0 as=7.2e+06 ps=19200 
M2233 diff_164640_128400# diff_164040_128160# GND GND efet w=3960 l=600
+ ad=6.2496e+06 pd=18480 as=0 ps=0 
M2234 diff_160560_126600# diff_159960_126240# GND GND efet w=3540 l=660
+ ad=3.2976e+06 pd=9360 as=0 ps=0 
M2235 GND diff_166080_132120# diff_164520_118080# GND efet w=3540 l=720
+ ad=0 pd=0 as=6.3648e+06 ps=17280 
M2236 GND diff_170160_132120# diff_168720_120240# GND efet w=3960 l=600
+ ad=0 pd=0 as=7.3872e+06 ps=19440 
M2237 diff_172800_128400# diff_172200_128160# GND GND efet w=3960 l=600
+ ad=6.3648e+06 pd=18720 as=0 ps=0 
M2238 diff_168720_126600# diff_168120_126240# GND GND efet w=3540 l=660
+ ad=3.2976e+06 pd=9360 as=0 ps=0 
M2239 GND diff_174240_132120# diff_172800_118080# GND efet w=3540 l=720
+ ad=0 pd=0 as=6.6816e+06 ps=17520 
M2240 GND diff_178320_132120# diff_177000_120240# GND efet w=3960 l=600
+ ad=0 pd=0 as=7.5744e+06 ps=19440 
M2241 diff_180960_128400# diff_180360_128160# GND GND efet w=3960 l=600
+ ad=6.6384e+06 pd=18720 as=0 ps=0 
M2242 diff_176880_126600# diff_176280_126240# GND GND efet w=3540 l=660
+ ad=3.2976e+06 pd=9360 as=0 ps=0 
M2243 GND diff_182400_132120# diff_180960_118080# GND efet w=3540 l=720
+ ad=0 pd=0 as=6.7392e+06 ps=17520 
M2244 GND diff_186480_132120# diff_185160_120240# GND efet w=3960 l=600
+ ad=0 pd=0 as=7.7616e+06 ps=19680 
M2245 diff_189120_128400# diff_188520_128160# GND GND efet w=3960 l=600
+ ad=6.3504e+06 pd=18720 as=0 ps=0 
M2246 diff_185040_126600# diff_184440_126240# GND GND efet w=3540 l=660
+ ad=3.2976e+06 pd=9360 as=0 ps=0 
M2247 GND diff_190560_132120# diff_189000_118080# GND efet w=3540 l=720
+ ad=0 pd=0 as=6.6816e+06 ps=17520 
M2248 GND diff_194640_132120# diff_193200_120240# GND efet w=3960 l=600
+ ad=0 pd=0 as=7.5744e+06 ps=19440 
M2249 diff_197280_128400# diff_196680_128160# GND GND efet w=3960 l=600
+ ad=6.6096e+06 pd=18720 as=0 ps=0 
M2250 diff_193200_126600# diff_192600_126240# GND GND efet w=3540 l=660
+ ad=3.2976e+06 pd=9360 as=0 ps=0 
M2251 GND diff_198720_132120# diff_197160_118080# GND efet w=3540 l=720
+ ad=0 pd=0 as=6.7392e+06 ps=17520 
M2252 GND diff_202800_132120# diff_201360_120240# GND efet w=3960 l=600
+ ad=0 pd=0 as=7.7616e+06 ps=19680 
M2253 diff_205440_128400# diff_204840_128160# GND GND efet w=3960 l=600
+ ad=6.3504e+06 pd=18720 as=0 ps=0 
M2254 diff_201360_126600# diff_200760_126240# GND GND efet w=3540 l=660
+ ad=3.2976e+06 pd=9360 as=0 ps=0 
M2255 GND diff_206880_132120# diff_205320_118080# GND efet w=3540 l=720
+ ad=0 pd=0 as=6.6816e+06 ps=17520 
M2256 GND diff_210960_132120# diff_209520_120240# GND efet w=3960 l=600
+ ad=0 pd=0 as=7.5744e+06 ps=19440 
M2257 diff_213600_128400# diff_213000_128160# GND GND efet w=3960 l=600
+ ad=6.6096e+06 pd=18720 as=0 ps=0 
M2258 diff_209520_126600# diff_208920_126240# GND GND efet w=3540 l=660
+ ad=3.2976e+06 pd=9360 as=0 ps=0 
M2259 GND diff_215040_132120# diff_213480_118080# GND efet w=3540 l=720
+ ad=0 pd=0 as=6.7392e+06 ps=17520 
M2260 GND diff_219120_132120# diff_217680_120240# GND efet w=3960 l=600
+ ad=0 pd=0 as=7.7616e+06 ps=19680 
M2261 diff_221760_128400# diff_221160_128160# GND GND efet w=3960 l=600
+ ad=6.1776e+06 pd=18240 as=0 ps=0 
M2262 diff_217680_126600# diff_217080_126240# GND GND efet w=3540 l=660
+ ad=3.2976e+06 pd=9360 as=0 ps=0 
M2263 GND diff_223200_132120# diff_221760_118080# GND efet w=3540 l=720
+ ad=0 pd=0 as=6.5952e+06 ps=17280 
M2264 GND diff_227280_132120# diff_225960_120240# GND efet w=3960 l=600
+ ad=0 pd=0 as=7.3584e+06 ps=19200 
M2265 diff_229920_128400# diff_229320_128160# GND GND efet w=3960 l=600
+ ad=8.0352e+06 pd=24960 as=0 ps=0 
M2266 diff_225840_126600# diff_225240_126240# GND GND efet w=3540 l=660
+ ad=3.2976e+06 pd=9360 as=0 ps=0 
M2267 diff_48840_127680# diff_26040_78600# GND GND efet w=4620 l=780
+ ad=0 pd=0 as=0 ps=0 
M2268 diff_49200_117000# Vdd Vdd GND efet w=600 l=1560
+ ad=0 pd=0 as=0 ps=0 
M2269 diff_50880_129960# Vdd Vdd GND efet w=600 l=1440
+ ad=0 pd=0 as=0 ps=0 
M2270 Vdd Vdd Vdd GND efet w=240 l=240
+ ad=0 pd=0 as=0 ps=0 
M2271 Vdd Vdd Vdd GND efet w=120 l=240
+ ad=0 pd=0 as=0 ps=0 
M2272 diff_64440_127680# cl GND GND efet w=3600 l=720
+ ad=0 pd=0 as=0 ps=0 
M2273 GND cl diff_64440_127680# GND efet w=3600 l=840
+ ad=0 pd=0 as=0 ps=0 
M2274 diff_64440_127680# diff_26040_78600# GND GND efet w=4860 l=780
+ ad=0 pd=0 as=0 ps=0 
M2275 diff_64680_117000# Vdd Vdd GND efet w=600 l=1560
+ ad=0 pd=0 as=0 ps=0 
M2276 diff_66600_129960# Vdd Vdd GND efet w=600 l=1440
+ ad=0 pd=0 as=0 ps=0 
M2277 Vdd Vdd Vdd GND efet w=120 l=120
+ ad=0 pd=0 as=0 ps=0 
M2278 Vdd Vdd Vdd GND efet w=120 l=120
+ ad=0 pd=0 as=0 ps=0 
M2279 diff_79920_127680# cl GND GND efet w=3600 l=720
+ ad=0 pd=0 as=0 ps=0 
M2280 GND cl diff_79920_127680# GND efet w=3600 l=840
+ ad=0 pd=0 as=0 ps=0 
M2281 diff_79920_127680# diff_26040_78600# GND GND efet w=4860 l=780
+ ad=0 pd=0 as=0 ps=0 
M2282 diff_99960_121680# diff_104880_84600# diff_103320_126720# GND efet w=3120 l=720
+ ad=2.03184e+07 pd=48000 as=0 ps=0 
M2283 diff_107760_120720# diff_104880_84600# diff_111600_126600# GND efet w=3000 l=600
+ ad=1.69056e+07 pd=40800 as=0 ps=0 
M2284 diff_115920_120720# diff_104880_84600# diff_119760_126600# GND efet w=3000 l=600
+ ad=1.7568e+07 pd=45840 as=0 ps=0 
M2285 diff_123960_120840# diff_104880_84600# diff_127920_126600# GND efet w=3000 l=600
+ ad=1.62e+07 pd=40320 as=0 ps=0 
M2286 diff_132120_120840# diff_104880_84600# diff_136080_126600# GND efet w=3000 l=600
+ ad=1.79712e+07 pd=46800 as=0 ps=0 
M2287 diff_140400_120600# diff_104880_84600# diff_144240_126600# GND efet w=3000 l=600
+ ad=1.74384e+07 pd=41280 as=0 ps=0 
M2288 diff_148560_120600# diff_104880_84600# diff_152400_126600# GND efet w=3000 l=600
+ ad=1.8576e+07 pd=47040 as=0 ps=0 
M2289 diff_156720_120600# diff_104880_84600# diff_160560_126600# GND efet w=3000 l=600
+ ad=1.74384e+07 pd=41280 as=0 ps=0 
M2290 diff_164880_120600# diff_104880_84600# diff_168720_126600# GND efet w=3000 l=600
+ ad=1.82016e+07 pd=46320 as=0 ps=0 
M2291 diff_173160_120720# diff_104880_84600# diff_176880_126600# GND efet w=3000 l=600
+ ad=1.69344e+07 pd=40800 as=0 ps=0 
M2292 diff_181320_120720# diff_104880_84600# diff_185040_126600# GND efet w=3000 l=600
+ ad=1.8e+07 pd=46080 as=0 ps=0 
M2293 diff_189360_120720# diff_104880_84600# diff_193200_126600# GND efet w=3000 l=600
+ ad=1.68768e+07 pd=40800 as=0 ps=0 
M2294 diff_197520_120720# diff_104880_84600# diff_201360_126600# GND efet w=3000 l=600
+ ad=1.8e+07 pd=46320 as=0 ps=0 
M2295 diff_205680_120720# diff_104880_84600# diff_209520_126600# GND efet w=3000 l=600
+ ad=1.68768e+07 pd=40800 as=0 ps=0 
M2296 diff_213840_120720# diff_104880_84600# diff_217680_126600# GND efet w=3000 l=600
+ ad=1.82304e+07 pd=46560 as=0 ps=0 
M2297 diff_222120_120600# diff_104880_84600# diff_225840_126600# GND efet w=3000 l=600
+ ad=1.77984e+07 pd=42480 as=0 ps=0 
M2298 diff_100440_136920# diff_243120_97920# diff_236760_140760# GND efet w=7920 l=600
+ ad=0 pd=0 as=0 ps=0 
M2299 diff_243720_169800# diff_245160_97920# diff_236760_140760# GND efet w=15480 l=720
+ ad=0 pd=0 as=0 ps=0 
M2300 diff_236760_149400# diff_246960_91200# diff_243720_169800# GND efet w=15480 l=720
+ ad=0 pd=0 as=0 ps=0 
M2301 diff_99960_121680# diff_99480_122520# diff_99720_123600# GND efet w=4080 l=600
+ ad=0 pd=0 as=0 ps=0 
M2302 diff_80160_117000# Vdd Vdd GND efet w=600 l=1560
+ ad=0 pd=0 as=0 ps=0 
M2303 diff_82080_129960# Vdd Vdd GND efet w=600 l=1440
+ ad=0 pd=0 as=0 ps=0 
M2304 diff_132000_128400# diff_99480_122520# diff_132120_120840# GND efet w=3420 l=600
+ ad=0 pd=0 as=0 ps=0 
M2305 diff_123840_128400# diff_99480_122520# diff_123960_120840# GND efet w=3120 l=660
+ ad=0 pd=0 as=0 ps=0 
M2306 diff_140160_128400# diff_99480_122520# diff_140400_120600# GND efet w=3120 l=660
+ ad=0 pd=0 as=0 ps=0 
M2307 diff_148320_128400# diff_99480_122520# diff_148560_120600# GND efet w=3240 l=600
+ ad=0 pd=0 as=0 ps=0 
M2308 diff_156480_128400# diff_99480_122520# diff_156720_120600# GND efet w=3120 l=660
+ ad=0 pd=0 as=0 ps=0 
M2309 diff_107520_128400# diff_99480_122520# diff_107760_120720# GND efet w=3060 l=660
+ ad=0 pd=0 as=0 ps=0 
M2310 diff_115680_128400# diff_99480_122520# diff_115920_120720# GND efet w=3120 l=660
+ ad=0 pd=0 as=0 ps=0 
M2311 diff_164640_128400# diff_99480_122520# diff_164880_120600# GND efet w=3120 l=660
+ ad=0 pd=0 as=0 ps=0 
M2312 diff_189120_128400# diff_99480_122520# diff_189360_120720# GND efet w=3060 l=660
+ ad=0 pd=0 as=0 ps=0 
M2313 diff_197280_128400# diff_99480_122520# diff_197520_120720# GND efet w=3120 l=660
+ ad=0 pd=0 as=0 ps=0 
M2314 diff_205440_128400# diff_99480_122520# diff_205680_120720# GND efet w=3060 l=660
+ ad=0 pd=0 as=0 ps=0 
M2315 diff_213600_128400# diff_99480_122520# diff_213840_120720# GND efet w=3120 l=660
+ ad=0 pd=0 as=0 ps=0 
M2316 Vdd Vdd Vdd GND efet w=120 l=120
+ ad=0 pd=0 as=0 ps=0 
M2317 Vdd Vdd Vdd GND efet w=120 l=120
+ ad=0 pd=0 as=0 ps=0 
M2318 diff_103680_120240# diff_103320_91920# diff_99960_121680# GND efet w=2880 l=600
+ ad=0 pd=0 as=0 ps=0 
M2319 diff_111600_120120# diff_103320_91920# diff_107760_120720# GND efet w=3420 l=660
+ ad=0 pd=0 as=0 ps=0 
M2320 diff_119760_120240# diff_103320_91920# diff_115920_120720# GND efet w=3360 l=840
+ ad=0 pd=0 as=0 ps=0 
M2321 diff_127800_120240# diff_103320_91920# diff_123960_120840# GND efet w=3360 l=780
+ ad=0 pd=0 as=0 ps=0 
M2322 diff_135960_120120# diff_103320_91920# diff_132120_120840# GND efet w=3480 l=600
+ ad=0 pd=0 as=0 ps=0 
M2323 diff_144240_120240# diff_103320_91920# diff_140400_120600# GND efet w=3360 l=780
+ ad=0 pd=0 as=0 ps=0 
M2324 diff_152400_120240# diff_103320_91920# diff_148560_120600# GND efet w=3420 l=840
+ ad=0 pd=0 as=0 ps=0 
M2325 diff_172800_128400# diff_99480_122520# diff_173160_120720# GND efet w=3000 l=600
+ ad=0 pd=0 as=0 ps=0 
M2326 diff_180960_128400# diff_99480_122520# diff_181320_120720# GND efet w=3060 l=660
+ ad=0 pd=0 as=0 ps=0 
M2327 diff_160560_120240# diff_103320_91920# diff_156720_120600# GND efet w=3360 l=780
+ ad=0 pd=0 as=0 ps=0 
M2328 diff_168720_120240# diff_103320_91920# diff_164880_120600# GND efet w=3360 l=840
+ ad=0 pd=0 as=0 ps=0 
M2329 diff_177000_120240# diff_103320_91920# diff_173160_120720# GND efet w=3300 l=780
+ ad=0 pd=0 as=0 ps=0 
M2330 diff_185160_120240# diff_103320_91920# diff_181320_120720# GND efet w=3300 l=780
+ ad=0 pd=0 as=0 ps=0 
M2331 diff_193200_120240# diff_103320_91920# diff_189360_120720# GND efet w=3360 l=840
+ ad=0 pd=0 as=0 ps=0 
M2332 diff_201360_120240# diff_103320_91920# diff_197520_120720# GND efet w=3360 l=840
+ ad=0 pd=0 as=0 ps=0 
M2333 diff_221760_128400# diff_99480_122520# diff_222120_120600# GND efet w=2880 l=600
+ ad=0 pd=0 as=0 ps=0 
M2334 diff_209520_120240# diff_103320_91920# diff_205680_120720# GND efet w=3360 l=840
+ ad=0 pd=0 as=0 ps=0 
M2335 diff_217680_120240# diff_103320_91920# diff_213840_120720# GND efet w=3360 l=840
+ ad=0 pd=0 as=0 ps=0 
M2336 diff_225960_120240# diff_103320_91920# diff_222120_120600# GND efet w=3180 l=780
+ ad=0 pd=0 as=0 ps=0 
M2337 GND diff_33600_117000# diff_33720_108720# GND efet w=5640 l=600
+ ad=0 pd=0 as=1.11456e+07 ps=25920 
M2338 GND diff_49200_117000# diff_49320_108720# GND efet w=5640 l=600
+ ad=0 pd=0 as=1.11744e+07 ps=25440 
M2339 Vdd Vdd diff_33720_108720# GND efet w=720 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2340 GND diff_64680_117000# diff_64800_108720# GND efet w=5640 l=600
+ ad=0 pd=0 as=1.17072e+07 ps=25920 
M2341 diff_33720_108720# diff_33720_108720# diff_33720_108720# GND efet w=180 l=180
+ ad=0 pd=0 as=0 ps=0 
M2342 diff_33720_108720# diff_33720_108720# diff_33720_108720# GND efet w=360 l=360
+ ad=0 pd=0 as=0 ps=0 
M2343 Vdd Vdd diff_49320_108720# GND efet w=720 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2344 GND diff_80160_117000# diff_80280_108720# GND efet w=5640 l=600
+ ad=0 pd=0 as=1.17216e+07 ps=26640 
M2345 diff_49320_108720# diff_49320_108720# diff_49320_108720# GND efet w=360 l=420
+ ad=0 pd=0 as=0 ps=0 
M2346 Vdd Vdd diff_64800_108720# GND efet w=720 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2347 diff_107400_118080# diff_106320_94080# diff_99960_121680# GND efet w=3120 l=600
+ ad=0 pd=0 as=0 ps=0 
M2348 diff_115560_118080# diff_106320_94080# diff_107760_120720# GND efet w=3120 l=600
+ ad=0 pd=0 as=0 ps=0 
M2349 diff_123600_118080# diff_106320_94080# diff_115920_120720# GND efet w=3120 l=600
+ ad=0 pd=0 as=0 ps=0 
M2350 diff_131760_118080# diff_106320_94080# diff_123960_120840# GND efet w=3120 l=600
+ ad=0 pd=0 as=0 ps=0 
M2351 diff_140040_118080# diff_106320_94080# diff_132120_120840# GND efet w=3120 l=600
+ ad=0 pd=0 as=0 ps=0 
M2352 diff_148200_118080# diff_106320_94080# diff_140400_120600# GND efet w=3120 l=600
+ ad=0 pd=0 as=0 ps=0 
M2353 diff_156360_118080# diff_106320_94080# diff_148560_120600# GND efet w=3120 l=600
+ ad=0 pd=0 as=0 ps=0 
M2354 diff_164520_118080# diff_106320_94080# diff_156720_120600# GND efet w=3120 l=600
+ ad=0 pd=0 as=0 ps=0 
M2355 diff_172800_118080# diff_106320_94080# diff_164880_120600# GND efet w=3120 l=600
+ ad=0 pd=0 as=0 ps=0 
M2356 diff_180960_118080# diff_106320_94080# diff_173160_120720# GND efet w=3120 l=600
+ ad=0 pd=0 as=0 ps=0 
M2357 diff_189000_118080# diff_106320_94080# diff_181320_120720# GND efet w=3120 l=600
+ ad=0 pd=0 as=0 ps=0 
M2358 diff_197160_118080# diff_106320_94080# diff_189360_120720# GND efet w=3120 l=600
+ ad=0 pd=0 as=0 ps=0 
M2359 diff_205320_118080# diff_106320_94080# diff_197520_120720# GND efet w=3120 l=600
+ ad=0 pd=0 as=0 ps=0 
M2360 diff_213480_118080# diff_106320_94080# diff_205680_120720# GND efet w=3120 l=600
+ ad=0 pd=0 as=0 ps=0 
M2361 diff_221760_118080# diff_106320_94080# diff_213840_120720# GND efet w=3000 l=600
+ ad=0 pd=0 as=0 ps=0 
M2362 diff_229920_128400# diff_106320_94080# diff_222120_120600# GND efet w=4620 l=660
+ ad=0 pd=0 as=0 ps=0 
M2363 diff_64800_108720# diff_64800_108720# diff_64800_108720# GND efet w=480 l=480
+ ad=0 pd=0 as=0 ps=0 
M2364 diff_80280_108720# diff_80280_108720# diff_80280_108720# GND efet w=240 l=240
+ ad=0 pd=0 as=0 ps=0 
M2365 Vdd Vdd diff_80280_108720# GND efet w=720 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2366 diff_80280_108720# diff_80280_108720# diff_80280_108720# GND efet w=420 l=420
+ ad=0 pd=0 as=0 ps=0 
M2367 diff_99960_121680# diff_101160_115320# diff_101640_96840# GND efet w=4080 l=720
+ ad=0 pd=0 as=3.5424e+07 ps=69120 
M2368 diff_107760_120720# diff_112440_115320# diff_101640_96840# GND efet w=4080 l=600
+ ad=0 pd=0 as=0 ps=0 
M2369 diff_123960_120840# diff_112440_115320# diff_118080_98520# GND efet w=4080 l=600
+ ad=0 pd=0 as=3.32496e+07 ps=65520 
M2370 diff_140400_120600# diff_112440_115320# diff_134280_112200# GND efet w=4080 l=600
+ ad=0 pd=0 as=3.72672e+07 ps=70080 
M2371 diff_156720_120600# diff_112440_115320# diff_150720_98400# GND efet w=4080 l=600
+ ad=0 pd=0 as=3.76704e+07 ps=69360 
M2372 diff_173160_120720# diff_112440_115320# diff_167040_98400# GND efet w=4080 l=600
+ ad=0 pd=0 as=3.45888e+07 ps=66000 
M2373 diff_189360_120720# diff_112440_115320# diff_183480_98400# GND efet w=4080 l=600
+ ad=0 pd=0 as=3.38544e+07 ps=63600 
M2374 diff_205680_120720# diff_112440_115320# diff_199680_98400# GND efet w=4080 l=600
+ ad=0 pd=0 as=3.75264e+07 ps=71520 
M2375 diff_222120_120600# diff_112440_115320# diff_216000_98520# GND efet w=3480 l=600
+ ad=0 pd=0 as=2.96208e+07 ps=57600 
M2376 Vdd diff_33720_108720# io3 GND efet w=17640 l=720
+ ad=0 pd=0 as=1.00282e+08 ps=193920 
M2377 d3 GND d3 GND efet w=17700 l=11220
+ ad=0 pd=0 as=0 ps=0 
M2378 GND diff_33600_117000# io3 GND efet w=18060 l=840
+ ad=0 pd=0 as=0 ps=0 
M2379 Vdd diff_49320_108720# io2 GND efet w=17760 l=720
+ ad=0 pd=0 as=9.5328e+07 ps=192720 
M2380 io2 GND io2 GND efet w=17580 l=10740
+ ad=0 pd=0 as=0 ps=0 
M2381 GND diff_49200_117000# io2 GND efet w=18060 l=840
+ ad=0 pd=0 as=0 ps=0 
M2382 Vdd diff_64800_108720# io1 GND efet w=17760 l=720
+ ad=0 pd=0 as=9.19152e+07 ps=185280 
M2383 GND diff_64680_117000# io1 GND efet w=18060 l=840
+ ad=0 pd=0 as=0 ps=0 
M2384 Vdd diff_80280_108720# io0 GND efet w=17640 l=720
+ ad=0 pd=0 as=9.51552e+07 ps=193680 
M2385 diff_49680_96720# diff_40680_69240# diff_40800_144840# GND efet w=2280 l=720
+ ad=8.9424e+06 pd=23040 as=1.25136e+07 ps=32640 
M2386 diff_54360_101760# diff_44640_90240# diff_49680_96720# GND efet w=2280 l=720
+ ad=1.09008e+07 pd=24480 as=0 ps=0 
M2387 diff_64800_96720# diff_40680_69240# diff_56280_144840# GND efet w=2280 l=720
+ ad=9.6048e+06 pd=24000 as=1.00656e+07 ps=26160 
M2388 diff_68280_103440# diff_44640_90240# diff_64800_96720# GND efet w=2280 l=720
+ ad=1.02528e+07 pd=21600 as=0 ps=0 
M2389 io1 GND io1 GND efet w=16740 l=12540
+ ad=0 pd=0 as=0 ps=0 
M2390 io3 GND io3 GND efet w=14940 l=7020
+ ad=0 pd=0 as=0 ps=0 
M2391 diff_49680_96720# diff_41160_86760# io3 GND efet w=2160 l=600
+ ad=0 pd=0 as=0 ps=0 
M2392 GND diff_80160_117000# io0 GND efet w=18060 l=840
+ ad=0 pd=0 as=0 ps=0 
M2393 diff_115920_120720# diff_101160_115320# diff_118080_98520# GND efet w=3960 l=720
+ ad=0 pd=0 as=0 ps=0 
M2394 diff_132120_120840# diff_101160_115320# diff_134280_112200# GND efet w=4080 l=720
+ ad=0 pd=0 as=0 ps=0 
M2395 diff_148560_120600# diff_101160_115320# diff_150720_98400# GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2396 diff_164880_120600# diff_101160_115320# diff_167040_98400# GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2397 diff_181320_120720# diff_101160_115320# diff_183480_98400# GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2398 diff_197520_120720# diff_101160_115320# diff_199680_98400# GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2399 diff_213840_120720# diff_101160_115320# diff_216000_98520# GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2400 diff_90120_96840# diff_40680_69240# diff_87360_144840# GND efet w=2160 l=720
+ ad=1.53504e+07 pd=40320 as=2.8224e+06 ps=6960 
M2401 diff_96720_108360# diff_44640_90240# diff_90120_96840# GND efet w=2160 l=720
+ ad=7.2432e+06 pd=16080 as=0 ps=0 
M2402 diff_80280_96720# diff_40680_69240# diff_71880_144840# GND efet w=2280 l=720
+ ad=1.0368e+07 pd=26400 as=8.8704e+06 ps=23280 
M2403 diff_82920_103920# diff_44640_90240# diff_80280_96720# GND efet w=2280 l=720
+ ad=1.6344e+07 pd=34320 as=0 ps=0 
M2404 io0 GND io0 GND efet w=17760 l=12960
+ ad=0 pd=0 as=0 ps=0 
M2405 io3 GND io3 GND efet w=2820 l=3420
+ ad=0 pd=0 as=0 ps=0 
M2406 GND diff_41160_86760# diff_44640_90240# GND efet w=1680 l=720
+ ad=0 pd=0 as=1.30464e+07 ps=42720 
M2407 diff_49440_88920# io3 GND GND efet w=3480 l=720
+ ad=8.352e+06 pd=18240 as=0 ps=0 
M2408 GND io3 diff_49440_88920# GND efet w=3480 l=720
+ ad=0 pd=0 as=0 ps=0 
M2409 diff_64800_96720# diff_41160_86760# io2 GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2410 diff_118080_98520# diff_56400_47520# diff_99960_108720# GND efet w=2280 l=600
+ ad=0 pd=0 as=1.57968e+07 ps=33120 
M2411 diff_96720_108360# diff_99960_108720# GND GND efet w=5040 l=600
+ ad=0 pd=0 as=0 ps=0 
M2412 diff_99960_108720# diff_99960_108720# diff_99960_108720# GND efet w=120 l=120
+ ad=0 pd=0 as=0 ps=0 
M2413 diff_96720_108360# Vdd Vdd GND efet w=960 l=2520
+ ad=0 pd=0 as=0 ps=0 
M2414 diff_99960_108720# diff_99960_108720# diff_99960_108720# GND efet w=120 l=240
+ ad=0 pd=0 as=0 ps=0 
M2415 diff_150720_98400# diff_56400_47520# diff_134400_100800# GND efet w=2400 l=600
+ ad=0 pd=0 as=1.4976e+07 ps=31680 
M2416 diff_183480_98400# diff_56400_47520# diff_167040_100800# GND efet w=2160 l=600
+ ad=0 pd=0 as=1.81296e+07 ps=33360 
M2417 Vdd Vdd Vdd GND efet w=240 l=300
+ ad=0 pd=0 as=0 ps=0 
M2418 Vdd Vdd Vdd GND efet w=240 l=300
+ ad=0 pd=0 as=0 ps=0 
M2419 diff_44640_90240# diff_44640_90240# diff_44640_90240# GND efet w=240 l=600
+ ad=0 pd=0 as=0 ps=0 
M2420 Vdd Vdd Vdd GND efet w=120 l=720
+ ad=0 pd=0 as=0 ps=0 
M2421 Vdd Vdd diff_118080_98520# GND efet w=660 l=6480
+ ad=0 pd=0 as=0 ps=0 
M2422 Vdd Vdd diff_101640_96840# GND efet w=600 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2423 Vdd Vdd Vdd GND efet w=120 l=540
+ ad=0 pd=0 as=0 ps=0 
M2424 diff_134400_100800# diff_134400_100800# diff_134400_100800# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M2425 diff_134400_100800# diff_134400_100800# diff_134400_100800# GND efet w=120 l=240
+ ad=0 pd=0 as=0 ps=0 
M2426 diff_150720_98400# Vdd Vdd GND efet w=600 l=6480
+ ad=0 pd=0 as=0 ps=0 
M2427 Vdd Vdd diff_82920_103920# GND efet w=840 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2428 Vdd Vdd Vdd GND efet w=120 l=480
+ ad=0 pd=0 as=0 ps=0 
M2429 Vdd Vdd diff_134280_112200# GND efet w=600 l=6480
+ ad=0 pd=0 as=0 ps=0 
M2430 Vdd Vdd Vdd GND efet w=240 l=480
+ ad=0 pd=0 as=0 ps=0 
M2431 diff_82920_103920# diff_134400_100800# GND GND efet w=4200 l=720
+ ad=0 pd=0 as=0 ps=0 
M2432 diff_167040_98400# Vdd Vdd GND efet w=660 l=6780
+ ad=0 pd=0 as=0 ps=0 
M2433 Vdd Vdd diff_68280_103440# GND efet w=840 l=3960
+ ad=0 pd=0 as=0 ps=0 
M2434 diff_216000_98520# diff_56400_47520# diff_199680_100800# GND efet w=2400 l=720
+ ad=0 pd=0 as=1.74096e+07 ps=32160 
M2435 diff_183480_98400# Vdd Vdd GND efet w=540 l=6660
+ ad=0 pd=0 as=0 ps=0 
M2436 diff_68280_103440# diff_167040_100800# GND GND efet w=5040 l=600
+ ad=0 pd=0 as=0 ps=0 
M2437 Vdd Vdd Vdd GND efet w=120 l=300
+ ad=0 pd=0 as=0 ps=0 
M2438 diff_134400_100800# diff_62400_47520# diff_134280_112200# GND efet w=2280 l=600
+ ad=0 pd=0 as=0 ps=0 
M2439 diff_199680_98400# Vdd Vdd GND efet w=780 l=6780
+ ad=0 pd=0 as=0 ps=0 
M2440 diff_167040_100800# diff_62400_47520# diff_167040_98400# GND efet w=2400 l=600
+ ad=0 pd=0 as=0 ps=0 
M2441 diff_199680_100800# diff_62400_47520# diff_199680_98400# GND efet w=2400 l=600
+ ad=0 pd=0 as=0 ps=0 
M2442 Vdd Vdd diff_54360_101760# GND efet w=840 l=2520
+ ad=0 pd=0 as=0 ps=0 
M2443 diff_216000_98520# Vdd Vdd GND efet w=720 l=7080
+ ad=0 pd=0 as=0 ps=0 
M2444 diff_54360_101760# diff_199680_100800# GND GND efet w=4080 l=600
+ ad=0 pd=0 as=0 ps=0 
M2445 Vdd Vdd diff_44640_90240# GND efet w=720 l=4440
+ ad=0 pd=0 as=0 ps=0 
M2446 diff_44640_90240# diff_44640_90240# diff_44640_90240# GND efet w=180 l=660
+ ad=0 pd=0 as=0 ps=0 
M2447 diff_99960_108720# diff_62400_47520# diff_101640_96840# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2448 io3 Vdd Vdd GND efet w=840 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2449 diff_56760_85560# diff_56760_85560# diff_56760_85560# GND efet w=180 l=360
+ ad=2.0016e+06 pd=7680 as=0 ps=0 
M2450 diff_41160_86760# diff_41160_86760# diff_41160_86760# GND efet w=60 l=180
+ ad=1.86192e+07 pd=54720 as=0 ps=0 
M2451 diff_41160_86760# diff_41160_86760# diff_41160_86760# GND efet w=60 l=120
+ ad=0 pd=0 as=0 ps=0 
M2452 diff_56760_85560# diff_56760_85560# diff_56760_85560# GND efet w=180 l=540
+ ad=0 pd=0 as=0 ps=0 
M2453 diff_41160_86760# diff_41160_86760# diff_41160_86760# GND efet w=120 l=360
+ ad=0 pd=0 as=0 ps=0 
M2454 diff_64680_88800# io2 GND GND efet w=3480 l=720
+ ad=8.4384e+06 pd=18480 as=0 ps=0 
M2455 GND io2 diff_64680_88800# GND efet w=3480 l=720
+ ad=0 pd=0 as=0 ps=0 
M2456 diff_80280_96720# diff_41160_86760# io1 GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2457 diff_90120_96840# diff_41160_86760# io0 GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2458 io2 Vdd Vdd GND efet w=840 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2459 diff_56760_85560# Vdd Vdd GND efet w=720 l=720
+ ad=0 pd=0 as=0 ps=0 
M2460 diff_41160_86760# clk1 diff_41160_85320# GND efet w=1080 l=720
+ ad=0 pd=0 as=2.8944e+06 ps=11040 
M2461 diff_41160_85320# diff_41160_85320# diff_41160_85320# GND efet w=180 l=420
+ ad=0 pd=0 as=0 ps=0 
M2462 GND diff_41160_85320# diff_44640_90240# GND efet w=3660 l=660
+ ad=0 pd=0 as=0 ps=0 
M2463 Vdd Vdd diff_49440_88920# GND efet w=720 l=2160
+ ad=0 pd=0 as=0 ps=0 
M2464 diff_41160_85320# diff_41160_85320# diff_41160_85320# GND efet w=180 l=240
+ ad=0 pd=0 as=0 ps=0 
M2465 Vdd Vdd Vdd GND efet w=120 l=360
+ ad=0 pd=0 as=0 ps=0 
M2466 Vdd diff_56760_85560# diff_41160_86760# GND efet w=900 l=2160
+ ad=0 pd=0 as=0 ps=0 
M2467 Vdd Vdd diff_48120_80160# GND efet w=720 l=1440
+ ad=0 pd=0 as=8.2224e+06 ps=22080 
M2468 diff_41160_86760# diff_56760_85560# diff_41160_86760# GND efet w=4680 l=300
+ ad=0 pd=0 as=0 ps=0 
M2469 diff_80160_88800# io1 GND GND efet w=3480 l=720
+ ad=8.352e+06 pd=18240 as=0 ps=0 
M2470 GND io1 diff_80160_88800# GND efet w=3480 l=720
+ ad=0 pd=0 as=0 ps=0 
M2471 diff_118080_98520# diff_101400_96240# diff_115920_90840# GND efet w=3960 l=720
+ ad=0 pd=0 as=1.69344e+07 ps=45360 
M2472 diff_134280_112200# diff_101400_96240# diff_132120_90480# GND efet w=3900 l=660
+ ad=0 pd=0 as=1.71504e+07 ps=46080 
M2473 diff_216000_98520# diff_101400_96240# diff_213840_90840# GND efet w=4080 l=720
+ ad=0 pd=0 as=1.7136e+07 ps=45840 
M2474 diff_150720_98400# diff_101400_96240# diff_148560_90720# GND efet w=3960 l=600
+ ad=0 pd=0 as=1.78848e+07 ps=46320 
M2475 diff_167040_98400# diff_101400_96240# diff_164880_90840# GND efet w=3960 l=600
+ ad=0 pd=0 as=1.7568e+07 ps=45840 
M2476 diff_101640_96840# diff_101400_96240# diff_99960_89640# GND efet w=4080 l=720
+ ad=0 pd=0 as=1.96128e+07 ps=47280 
M2477 diff_101640_96840# diff_112440_96360# diff_107760_90720# GND efet w=4080 l=600
+ ad=0 pd=0 as=1.62864e+07 ps=40320 
M2478 diff_118080_98520# diff_112440_96360# diff_123960_90720# GND efet w=4080 l=600
+ ad=0 pd=0 as=1.55808e+07 ps=39840 
M2479 diff_134280_112200# diff_112440_96360# diff_140400_90720# GND efet w=4080 l=600
+ ad=0 pd=0 as=1.68192e+07 ps=40800 
M2480 diff_150720_98400# diff_112440_96360# diff_156720_90720# GND efet w=4080 l=600
+ ad=0 pd=0 as=1.68192e+07 ps=40800 
M2481 diff_183480_98400# diff_101400_96240# diff_181320_90840# GND efet w=3960 l=600
+ ad=0 pd=0 as=1.73664e+07 ps=45600 
M2482 diff_167040_98400# diff_112440_96360# diff_173160_90720# GND efet w=4080 l=600
+ ad=0 pd=0 as=1.63152e+07 ps=40320 
M2483 diff_199680_98400# diff_101400_96240# diff_197520_90840# GND efet w=3960 l=600
+ ad=0 pd=0 as=1.73088e+07 ps=45600 
M2484 diff_183480_98400# diff_112440_96360# diff_189360_90720# GND efet w=4080 l=600
+ ad=0 pd=0 as=1.62576e+07 ps=40320 
M2485 diff_199680_98400# diff_112440_96360# diff_205680_90720# GND efet w=4080 l=600
+ ad=0 pd=0 as=1.62576e+07 ps=40320 
M2486 diff_216000_98520# diff_112440_96360# diff_222120_90720# GND efet w=3480 l=480
+ ad=0 pd=0 as=1.70496e+07 ps=41760 
M2487 diff_229920_82920# diff_106320_94080# diff_222120_90720# GND efet w=4380 l=660
+ ad=8.5968e+06 pd=24960 as=0 ps=0 
M2488 diff_99960_89640# diff_106320_94080# diff_107400_92760# GND efet w=3120 l=600
+ ad=0 pd=0 as=7.0704e+06 ps=17760 
M2489 diff_107760_90720# diff_106320_94080# diff_115560_92760# GND efet w=3120 l=600
+ ad=0 pd=0 as=7.128e+06 ps=17760 
M2490 diff_115920_90840# diff_106320_94080# diff_123600_92640# GND efet w=3120 l=600
+ ad=0 pd=0 as=7.4448e+06 ps=18000 
M2491 diff_123960_90720# diff_106320_94080# diff_131760_92640# GND efet w=3120 l=600
+ ad=0 pd=0 as=7.5024e+06 ps=18000 
M2492 diff_132120_90480# diff_106320_94080# diff_140040_92880# GND efet w=3120 l=600
+ ad=0 pd=0 as=6.696e+06 ps=17520 
M2493 diff_140400_90720# diff_106320_94080# diff_148200_92880# GND efet w=3120 l=600
+ ad=0 pd=0 as=6.7536e+06 ps=17520 
M2494 diff_148560_90720# diff_106320_94080# diff_156360_92880# GND efet w=3120 l=600
+ ad=0 pd=0 as=6.696e+06 ps=17520 
M2495 diff_156720_90720# diff_106320_94080# diff_164520_92880# GND efet w=3120 l=600
+ ad=0 pd=0 as=6.7536e+06 ps=17520 
M2496 diff_164880_90840# diff_106320_94080# diff_172800_92760# GND efet w=3120 l=600
+ ad=0 pd=0 as=7.0704e+06 ps=17760 
M2497 diff_173160_90720# diff_106320_94080# diff_180960_92760# GND efet w=3120 l=600
+ ad=0 pd=0 as=7.128e+06 ps=17760 
M2498 diff_181320_90840# diff_106320_94080# diff_189000_92760# GND efet w=3120 l=600
+ ad=0 pd=0 as=7.0704e+06 ps=17760 
M2499 diff_189360_90720# diff_106320_94080# diff_197160_92760# GND efet w=3120 l=600
+ ad=0 pd=0 as=7.128e+06 ps=17760 
M2500 diff_197520_90840# diff_106320_94080# diff_205320_92760# GND efet w=3120 l=600
+ ad=0 pd=0 as=7.0704e+06 ps=17760 
M2501 diff_205680_90720# diff_106320_94080# diff_213480_92760# GND efet w=3120 l=600
+ ad=0 pd=0 as=7.128e+06 ps=17760 
M2502 diff_213840_90840# diff_106320_94080# diff_221760_92760# GND efet w=3000 l=600
+ ad=0 pd=0 as=6.9696e+06 ps=17520 
M2503 io1 Vdd Vdd GND efet w=840 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2504 diff_89880_88800# io0 GND GND efet w=3480 l=720
+ ad=8.4384e+06 pd=18480 as=0 ps=0 
M2505 GND io0 diff_89880_88800# GND efet w=3480 l=720
+ ad=0 pd=0 as=0 ps=0 
M2506 io0 Vdd Vdd GND efet w=840 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2507 Vdd Vdd diff_64680_88800# GND efet w=720 l=2280
+ ad=0 pd=0 as=0 ps=0 
M2508 Vdd Vdd diff_80160_88800# GND efet w=720 l=2160
+ ad=0 pd=0 as=0 ps=0 
M2509 Vdd Vdd diff_89880_88800# GND efet w=720 l=2040
+ ad=0 pd=0 as=0 ps=0 
M2510 GND diff_49680_79800# diff_48120_80160# GND efet w=6120 l=720
+ ad=0 pd=0 as=0 ps=0 
M2511 diff_48120_80160# diff_40680_69240# diff_44760_77160# GND efet w=1200 l=720
+ ad=0 pd=0 as=1.6704e+06 ps=5280 
M2512 diff_107760_90720# diff_103320_91920# diff_111600_90720# GND efet w=3420 l=660
+ ad=0 pd=0 as=7.9056e+06 ps=19920 
M2513 diff_115920_90840# diff_103320_91920# diff_119760_90720# GND efet w=3360 l=840
+ ad=0 pd=0 as=8.0784e+06 ps=19920 
M2514 diff_132120_90480# diff_103320_91920# diff_135960_90600# GND efet w=3480 l=600
+ ad=0 pd=0 as=8.4672e+06 ps=20400 
M2515 diff_123960_90720# diff_103320_91920# diff_127800_90600# GND efet w=3360 l=780
+ ad=0 pd=0 as=8.2656e+06 ps=19920 
M2516 diff_140400_90720# diff_103320_91920# diff_144240_90840# GND efet w=3360 l=780
+ ad=0 pd=0 as=7.5168e+06 ps=19440 
M2517 diff_148560_90720# diff_103320_91920# diff_152400_90840# GND efet w=3420 l=840
+ ad=0 pd=0 as=7.704e+06 ps=19680 
M2518 diff_156720_90720# diff_103320_91920# diff_160560_90840# GND efet w=3360 l=780
+ ad=0 pd=0 as=7.5168e+06 ps=19440 
M2519 diff_164880_90840# diff_103320_91920# diff_168720_90840# GND efet w=3360 l=840
+ ad=0 pd=0 as=7.704e+06 ps=19680 
M2520 diff_173160_90720# diff_103320_91920# diff_177000_90720# GND efet w=3300 l=780
+ ad=0 pd=0 as=7.8912e+06 ps=19680 
M2521 diff_189360_90720# diff_103320_91920# diff_193200_90720# GND efet w=3360 l=840
+ ad=0 pd=0 as=7.8912e+06 ps=19680 
M2522 diff_181320_90840# diff_103320_91920# diff_185160_90720# GND efet w=3300 l=780
+ ad=0 pd=0 as=8.0784e+06 ps=19920 
M2523 diff_197520_90840# diff_103320_91920# diff_201360_90720# GND efet w=3360 l=840
+ ad=0 pd=0 as=8.0784e+06 ps=19920 
M2524 diff_205680_90720# diff_103320_91920# diff_209520_90720# GND efet w=3360 l=840
+ ad=0 pd=0 as=7.8912e+06 ps=19680 
M2525 diff_213840_90840# diff_103320_91920# diff_217680_90720# GND efet w=3360 l=840
+ ad=0 pd=0 as=8.0784e+06 ps=19920 
M2526 diff_222120_90720# diff_103320_91920# diff_225960_90720# GND efet w=3240 l=840
+ ad=0 pd=0 as=7.6464e+06 ps=19440 
M2527 diff_41160_86760# diff_41160_86760# diff_41160_86760# GND efet w=120 l=120
+ ad=0 pd=0 as=0 ps=0 
M2528 diff_99960_89640# diff_103320_91920# diff_103680_90360# GND efet w=2880 l=600
+ ad=0 pd=0 as=7.8336e+06 ps=19440 
M2529 diff_107760_90720# diff_99480_122520# diff_107520_82680# GND efet w=3060 l=660
+ ad=0 pd=0 as=6.7104e+06 ps=18960 
M2530 diff_115920_90840# diff_99480_122520# diff_115680_82920# GND efet w=3120 l=660
+ ad=0 pd=0 as=6.912e+06 ps=18960 
M2531 diff_132120_90480# diff_99480_122520# diff_132000_82920# GND efet w=3420 l=600
+ ad=0 pd=0 as=7.1712e+06 ps=19200 
M2532 diff_123960_90720# diff_99480_122520# diff_123840_82920# GND efet w=3120 l=660
+ ad=0 pd=0 as=6.8544e+06 ps=18960 
M2533 diff_140400_90720# diff_99480_122520# diff_140160_82920# GND efet w=3120 l=660
+ ad=0 pd=0 as=6.264e+06 ps=18720 
M2534 diff_148560_90720# diff_99480_122520# diff_148320_82920# GND efet w=3240 l=600
+ ad=0 pd=0 as=6.5088e+06 ps=18720 
M2535 diff_156720_90720# diff_99480_122520# diff_156480_82920# GND efet w=3120 l=660
+ ad=0 pd=0 as=6.264e+06 ps=18720 
M2536 diff_164880_90840# diff_99480_122520# diff_164640_82920# GND efet w=3120 l=660
+ ad=0 pd=0 as=6.552e+06 ps=18720 
M2537 diff_173160_90720# diff_99480_122520# diff_172800_82920# GND efet w=3000 l=600
+ ad=0 pd=0 as=6.6672e+06 ps=18960 
M2538 diff_181320_90840# diff_99480_122520# diff_180960_82920# GND efet w=3060 l=660
+ ad=0 pd=0 as=6.9408e+06 ps=18960 
M2539 diff_189360_90720# diff_99480_122520# diff_189120_82920# GND efet w=3060 l=660
+ ad=0 pd=0 as=6.6528e+06 ps=18960 
M2540 diff_197520_90840# diff_99480_122520# diff_197280_82920# GND efet w=3120 l=660
+ ad=0 pd=0 as=6.912e+06 ps=18960 
M2541 diff_205680_90720# diff_99480_122520# diff_205440_82920# GND efet w=3060 l=660
+ ad=0 pd=0 as=6.6528e+06 ps=18960 
M2542 diff_213840_90840# diff_99480_122520# diff_213600_82920# GND efet w=3120 l=660
+ ad=0 pd=0 as=6.912e+06 ps=18960 
M2543 diff_222120_90720# diff_99480_122520# diff_221760_82920# GND efet w=2880 l=600
+ ad=0 pd=0 as=6.4656e+06 ps=18480 
M2544 diff_99960_89640# diff_99480_122520# diff_99720_83640# GND efet w=3840 l=480
+ ad=0 pd=0 as=8.3952e+06 ps=19440 
M2545 diff_103320_85080# diff_102480_84960# GND GND efet w=4680 l=720
+ ad=3.6432e+06 pd=10560 as=0 ps=0 
M2546 diff_41160_86760# diff_41160_86760# diff_41160_86760# GND efet w=60 l=180
+ ad=0 pd=0 as=0 ps=0 
M2547 GND diff_44760_77160# diff_18960_80400# GND efet w=9120 l=720
+ ad=0 pd=0 as=5.35104e+07 ps=118080 
M2548 diff_18960_80400# diff_42120_72840# Vdd GND efet w=8340 l=660
+ ad=0 pd=0 as=0 ps=0 
M2549 diff_55800_76560# diff_40920_47640# diff_53640_77640# GND efet w=3600 l=720
+ ad=8.64e+06 pd=22800 as=8.4528e+06 ps=22080 
M2550 diff_53640_77640# diff_33960_53280# diff_49680_79800# GND efet w=3960 l=720
+ ad=0 pd=0 as=6.0192e+06 ps=15120 
M2551 GND diff_100800_77520# diff_99720_83640# GND efet w=2880 l=600
+ ad=0 pd=0 as=0 ps=0 
M2552 diff_99960_89640# diff_104880_84600# diff_103320_85080# GND efet w=3120 l=600
+ ad=0 pd=0 as=0 ps=0 
M2553 GND diff_108960_77520# diff_107400_92760# GND efet w=3540 l=780
+ ad=0 pd=0 as=0 ps=0 
M2554 diff_111600_84960# diff_111000_77520# GND GND efet w=3600 l=720
+ ad=3.3264e+06 pd=9360 as=0 ps=0 
M2555 diff_107760_90720# diff_104880_84600# diff_111600_84960# GND efet w=3000 l=600
+ ad=0 pd=0 as=0 ps=0 
M2556 GND diff_117120_77520# diff_115560_92760# GND efet w=3540 l=780
+ ad=0 pd=0 as=0 ps=0 
M2557 diff_119760_84960# diff_119160_77520# GND GND efet w=3600 l=720
+ ad=3.3264e+06 pd=9360 as=0 ps=0 
M2558 diff_115920_90840# diff_104880_84600# diff_119760_84960# GND efet w=3000 l=600
+ ad=0 pd=0 as=0 ps=0 
M2559 GND diff_125280_77520# diff_123600_92640# GND efet w=3540 l=780
+ ad=0 pd=0 as=0 ps=0 
M2560 diff_127920_84960# diff_127320_77520# GND GND efet w=3600 l=720
+ ad=3.3264e+06 pd=9360 as=0 ps=0 
M2561 diff_123960_90720# diff_104880_84600# diff_127920_84960# GND efet w=3000 l=600
+ ad=0 pd=0 as=0 ps=0 
M2562 GND diff_133440_77520# diff_131760_92640# GND efet w=3540 l=780
+ ad=0 pd=0 as=0 ps=0 
M2563 diff_136080_84960# diff_135480_77520# GND GND efet w=3600 l=720
+ ad=3.3264e+06 pd=9360 as=0 ps=0 
M2564 diff_132120_90480# diff_104880_84600# diff_136080_84960# GND efet w=3000 l=600
+ ad=0 pd=0 as=0 ps=0 
M2565 GND diff_141600_77520# diff_140040_92880# GND efet w=3540 l=780
+ ad=0 pd=0 as=0 ps=0 
M2566 diff_144240_84960# diff_143640_77520# GND GND efet w=3600 l=720
+ ad=3.3264e+06 pd=9360 as=0 ps=0 
M2567 diff_140400_90720# diff_104880_84600# diff_144240_84960# GND efet w=3000 l=600
+ ad=0 pd=0 as=0 ps=0 
M2568 GND diff_149760_77520# diff_148200_92880# GND efet w=3540 l=780
+ ad=0 pd=0 as=0 ps=0 
M2569 diff_152400_84960# diff_151800_77520# GND GND efet w=3600 l=720
+ ad=3.3264e+06 pd=9360 as=0 ps=0 
M2570 diff_148560_90720# diff_104880_84600# diff_152400_84960# GND efet w=3000 l=600
+ ad=0 pd=0 as=0 ps=0 
M2571 GND diff_157920_77520# diff_156360_92880# GND efet w=3540 l=780
+ ad=0 pd=0 as=0 ps=0 
M2572 diff_160560_84960# diff_159960_77520# GND GND efet w=3600 l=720
+ ad=3.3264e+06 pd=9360 as=0 ps=0 
M2573 diff_156720_90720# diff_104880_84600# diff_160560_84960# GND efet w=3000 l=600
+ ad=0 pd=0 as=0 ps=0 
M2574 GND diff_166080_77520# diff_164520_92880# GND efet w=3540 l=780
+ ad=0 pd=0 as=0 ps=0 
M2575 diff_168720_84960# diff_168120_77520# GND GND efet w=3600 l=720
+ ad=3.3264e+06 pd=9360 as=0 ps=0 
M2576 diff_164880_90840# diff_104880_84600# diff_168720_84960# GND efet w=3000 l=600
+ ad=0 pd=0 as=0 ps=0 
M2577 GND diff_174240_77520# diff_172800_92760# GND efet w=3540 l=780
+ ad=0 pd=0 as=0 ps=0 
M2578 diff_176880_84960# diff_176280_77520# GND GND efet w=3600 l=720
+ ad=3.3264e+06 pd=9360 as=0 ps=0 
M2579 diff_173160_90720# diff_104880_84600# diff_176880_84960# GND efet w=3000 l=600
+ ad=0 pd=0 as=0 ps=0 
M2580 GND diff_182400_77520# diff_180960_92760# GND efet w=3540 l=780
+ ad=0 pd=0 as=0 ps=0 
M2581 diff_185040_84960# diff_184440_77520# GND GND efet w=3600 l=720
+ ad=3.3264e+06 pd=9360 as=0 ps=0 
M2582 diff_181320_90840# diff_104880_84600# diff_185040_84960# GND efet w=3000 l=600
+ ad=0 pd=0 as=0 ps=0 
M2583 GND diff_190560_77520# diff_189000_92760# GND efet w=3540 l=780
+ ad=0 pd=0 as=0 ps=0 
M2584 diff_193200_84960# diff_192600_77520# GND GND efet w=3600 l=720
+ ad=3.3264e+06 pd=9360 as=0 ps=0 
M2585 diff_189360_90720# diff_104880_84600# diff_193200_84960# GND efet w=3000 l=600
+ ad=0 pd=0 as=0 ps=0 
M2586 GND diff_198720_77520# diff_197160_92760# GND efet w=3540 l=780
+ ad=0 pd=0 as=0 ps=0 
M2587 diff_201360_84960# diff_200760_77520# GND GND efet w=3600 l=720
+ ad=3.3264e+06 pd=9360 as=0 ps=0 
M2588 diff_197520_90840# diff_104880_84600# diff_201360_84960# GND efet w=3000 l=600
+ ad=0 pd=0 as=0 ps=0 
M2589 GND diff_206880_77520# diff_205320_92760# GND efet w=3540 l=780
+ ad=0 pd=0 as=0 ps=0 
M2590 diff_209520_84960# diff_208920_77520# GND GND efet w=3600 l=720
+ ad=3.3264e+06 pd=9360 as=0 ps=0 
M2591 diff_205680_90720# diff_104880_84600# diff_209520_84960# GND efet w=3000 l=600
+ ad=0 pd=0 as=0 ps=0 
M2592 GND diff_215040_77520# diff_213480_92760# GND efet w=3540 l=780
+ ad=0 pd=0 as=0 ps=0 
M2593 diff_217680_84960# diff_217080_77520# GND GND efet w=3600 l=720
+ ad=3.3264e+06 pd=9360 as=0 ps=0 
M2594 diff_213840_90840# diff_104880_84600# diff_217680_84960# GND efet w=3000 l=600
+ ad=0 pd=0 as=0 ps=0 
M2595 GND diff_223200_77520# diff_221760_92760# GND efet w=3540 l=780
+ ad=0 pd=0 as=0 ps=0 
M2596 diff_225840_84960# diff_225240_77520# GND GND efet w=3600 l=720
+ ad=3.3264e+06 pd=9360 as=0 ps=0 
M2597 diff_222120_90720# diff_104880_84600# diff_225840_84960# GND efet w=3000 l=600
+ ad=0 pd=0 as=0 ps=0 
M2598 diff_259200_153240# Vdd Vdd GND efet w=1320 l=720
+ ad=1.5696e+06 pd=5760 as=0 ps=0 
M2599 diff_259200_153240# diff_259200_153240# diff_259200_153240# GND efet w=180 l=540
+ ad=0 pd=0 as=0 ps=0 
M2600 diff_259200_153240# diff_259200_153240# diff_259200_153240# GND efet w=180 l=180
+ ad=0 pd=0 as=0 ps=0 
M2601 Vdd Vdd Vdd GND efet w=60 l=180
+ ad=0 pd=0 as=0 ps=0 
M2602 GND diff_276720_158280# diff_264960_151920# GND efet w=8040 l=600
+ ad=0 pd=0 as=1.30896e+07 ps=25200 
M2603 Vdd Vdd diff_264960_151920# GND efet w=840 l=1680
+ ad=0 pd=0 as=0 ps=0 
M2604 Vdd Vdd Vdd GND efet w=60 l=120
+ ad=0 pd=0 as=0 ps=0 
M2605 GND d2 diff_281280_100320# GND efet w=19560 l=600
+ ad=0 pd=0 as=2.04336e+07 ps=39600 
M2606 diff_281280_100320# Vdd Vdd GND efet w=840 l=1680
+ ad=0 pd=0 as=0 ps=0 
M2607 diff_264960_151920# clk1 diff_276840_154080# GND efet w=1320 l=600
+ ad=0 pd=0 as=1.6848e+06 ps=5520 
M2608 Vdd Vdd diff_281280_113400# GND efet w=840 l=1680
+ ad=0 pd=0 as=1.09296e+07 ps=22800 
M2609 diff_276840_154080# diff_276840_154080# diff_276840_154080# GND efet w=180 l=180
+ ad=0 pd=0 as=0 ps=0 
M2610 GND diff_276840_154080# diff_271080_135600# GND efet w=4440 l=600
+ ad=0 pd=0 as=0 ps=0 
M2611 Vdd Vdd diff_271080_135600# GND efet w=960 l=1920
+ ad=0 pd=0 as=0 ps=0 
M2612 Vdd Vdd Vdd GND efet w=240 l=480
+ ad=0 pd=0 as=0 ps=0 
M2613 Vdd Vdd Vdd GND efet w=240 l=300
+ ad=0 pd=0 as=0 ps=0 
M2614 diff_271080_135600# clk2 diff_276840_149760# GND efet w=1200 l=600
+ ad=0 pd=0 as=1.3824e+06 ps=4800 
M2615 diff_100320_170280# diff_258960_146400# Vdd GND efet w=1560 l=600
+ ad=3.87072e+07 pd=73920 as=0 ps=0 
M2616 GND diff_264960_142800# diff_100320_170280# GND efet w=29640 l=600
+ ad=0 pd=0 as=0 ps=0 
M2617 diff_100320_170280# diff_258960_146400# diff_100320_170280# GND efet w=4080 l=480
+ ad=0 pd=0 as=0 ps=0 
M2618 diff_258960_146400# Vdd Vdd GND efet w=1200 l=600
+ ad=1.7424e+06 pd=6000 as=0 ps=0 
M2619 diff_258960_146400# diff_258960_146400# diff_258960_146400# GND efet w=120 l=480
+ ad=0 pd=0 as=0 ps=0 
M2620 diff_258960_146400# diff_258960_146400# diff_258960_146400# GND efet w=180 l=180
+ ad=0 pd=0 as=0 ps=0 
M2621 diff_276840_149760# diff_276840_149760# diff_276840_149760# GND efet w=120 l=240
+ ad=0 pd=0 as=0 ps=0 
M2622 GND diff_276840_149760# diff_266400_142200# GND efet w=4440 l=720
+ ad=0 pd=0 as=1.56816e+07 ps=33600 
M2623 Vdd Vdd diff_266400_142200# GND efet w=840 l=1800
+ ad=0 pd=0 as=0 ps=0 
M2624 Vdd Vdd Vdd GND efet w=60 l=180
+ ad=0 pd=0 as=0 ps=0 
M2625 GND diff_281280_100320# diff_281280_113400# GND efet w=4440 l=600
+ ad=0 pd=0 as=0 ps=0 
M2626 diff_266400_142200# clk1 diff_276720_145680# GND efet w=1440 l=600
+ ad=0 pd=0 as=1.6704e+06 ps=5280 
M2627 GND diff_276720_145680# diff_272280_84480# GND efet w=4440 l=600
+ ad=0 pd=0 as=1.13616e+07 ps=22560 
M2628 Vdd Vdd diff_272280_84480# GND efet w=840 l=1680
+ ad=0 pd=0 as=0 ps=0 
M2629 Vdd Vdd Vdd GND efet w=120 l=120
+ ad=0 pd=0 as=0 ps=0 
M2630 Vdd Vdd Vdd GND efet w=120 l=180
+ ad=0 pd=0 as=0 ps=0 
M2631 GND diff_266400_142200# diff_262680_141120# GND efet w=1320 l=600
+ ad=0 pd=0 as=4.824e+06 ps=13920 
M2632 diff_262680_141120# Vdd Vdd GND efet w=720 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2633 diff_260520_137280# Vdd Vdd GND efet w=720 l=1800
+ ad=7.1568e+06 pd=17520 as=0 ps=0 
M2634 diff_270840_139200# diff_266400_142200# diff_260160_136800# GND efet w=1560 l=600
+ ad=2.8368e+06 pd=8880 as=5.1552e+06 ps=13680 
M2635 diff_260520_137280# diff_260160_136800# GND GND efet w=6120 l=600
+ ad=0 pd=0 as=0 ps=0 
M2636 diff_260160_136800# diff_260160_136800# diff_260160_136800# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M2637 diff_260160_136800# diff_260160_136800# diff_260160_136800# GND efet w=180 l=180
+ ad=0 pd=0 as=0 ps=0 
M2638 diff_270840_139200# diff_261360_171960# diff_271080_135600# GND efet w=1320 l=600
+ ad=0 pd=0 as=0 ps=0 
M2639 diff_260160_136800# diff_262680_141120# GND GND efet w=1200 l=600
+ ad=0 pd=0 as=0 ps=0 
M2640 diff_273840_127440# diff_271080_135600# diff_252600_124320# GND efet w=2040 l=600
+ ad=5.688e+06 pd=13680 as=2.9088e+06 ps=6960 
M2641 diff_277440_130800# clk2 diff_273840_127440# GND efet w=2040 l=600
+ ad=9.9216e+06 pd=16320 as=0 ps=0 
M2642 GND diff_256800_128160# diff_112440_115320# GND efet w=14040 l=600
+ ad=0 pd=0 as=1.95408e+07 ps=39600 
M2643 diff_273840_127440# diff_272280_84480# diff_256800_128160# GND efet w=1920 l=600
+ ad=0 pd=0 as=2.5056e+06 ps=6480 
M2644 GND diff_41160_86760# diff_53640_77640# GND efet w=2700 l=780
+ ad=0 pd=0 as=0 ps=0 
M2645 diff_55800_76560# diff_56400_47520# GND GND efet w=3720 l=720
+ ad=0 pd=0 as=0 ps=0 
M2646 GND diff_62400_47520# diff_55800_76560# GND efet w=3600 l=720
+ ad=0 pd=0 as=0 ps=0 
M2647 diff_82560_78240# d3 GND GND efet w=3660 l=660
+ ad=8.8704e+06 pd=21120 as=0 ps=0 
M2648 GND diff_70080_67920# diff_69600_78240# GND efet w=2160 l=720
+ ad=0 pd=0 as=3.4272e+06 ps=8160 
M2649 GND diff_69600_78240# diff_15480_82200# GND efet w=1680 l=720
+ ad=0 pd=0 as=2.32992e+07 ps=73680 
M2650 diff_81600_78720# clk2 diff_70080_67920# GND efet w=1080 l=720
+ ad=1.0368e+06 pd=4080 as=3.4272e+06 ps=11040 
M2651 Vdd diff_82560_78240# diff_81600_78720# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M2652 diff_82560_78240# Vdd Vdd GND efet w=720 l=3360
+ ad=0 pd=0 as=0 ps=0 
M2653 GND diff_69480_55680# diff_82560_78240# GND efet w=1800 l=720
+ ad=0 pd=0 as=0 ps=0 
M2654 GND diff_91920_42120# diff_82560_78240# GND efet w=1800 l=720
+ ad=0 pd=0 as=0 ps=0 
M2655 GND diff_104880_77520# diff_103680_90360# GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2656 diff_107520_82680# diff_106920_77520# GND GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2657 GND diff_113040_77520# diff_111600_90720# GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2658 diff_115680_82920# diff_115080_77520# GND GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2659 GND diff_121200_77520# diff_119760_90720# GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2660 diff_123840_82920# diff_123240_77520# GND GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2661 GND diff_129360_77520# diff_127800_90600# GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2662 diff_132000_82920# diff_131400_77520# GND GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2663 GND diff_137520_77520# diff_135960_90600# GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2664 diff_140160_82920# diff_139560_77520# GND GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2665 GND diff_145680_77520# diff_144240_90840# GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2666 diff_148320_82920# diff_147720_77520# GND GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2667 GND diff_153840_77520# diff_152400_90840# GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2668 diff_156480_82920# diff_155880_77520# GND GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2669 GND diff_162000_77520# diff_160560_90840# GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2670 diff_164640_82920# diff_164040_77520# GND GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2671 GND diff_170160_77520# diff_168720_90840# GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2672 diff_172800_82920# diff_172200_77520# GND GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2673 GND diff_178320_77520# diff_177000_90720# GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2674 diff_180960_82920# diff_180360_77520# GND GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2675 GND diff_186480_77520# diff_185160_90720# GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2676 diff_189120_82920# diff_188520_77520# GND GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2677 GND diff_194640_77520# diff_193200_90720# GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2678 diff_197280_82920# diff_196680_77520# GND GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2679 GND diff_202800_77520# diff_201360_90720# GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2680 diff_205440_82920# diff_204840_77520# GND GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2681 GND diff_210960_77520# diff_209520_90720# GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2682 diff_213600_82920# diff_213000_77520# GND GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2683 GND diff_219120_77520# diff_217680_90720# GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2684 diff_221760_82920# diff_221160_77520# GND GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2685 GND diff_227280_77520# diff_225960_90720# GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2686 diff_229920_82920# diff_229320_77520# GND GND efet w=3960 l=600
+ ad=0 pd=0 as=0 ps=0 
M2687 GND diff_48120_80160# diff_49800_71520# GND efet w=4860 l=660
+ ad=0 pd=0 as=3.9024e+06 ps=12480 
M2688 diff_49800_71520# diff_40680_69240# diff_42120_72840# GND efet w=1080 l=600
+ ad=0 pd=0 as=3.1248e+06 ps=10080 
M2689 diff_49800_71520# Vdd Vdd GND efet w=720 l=1560
+ ad=0 pd=0 as=0 ps=0 
M2690 Vdd Vdd Vdd GND efet w=120 l=480
+ ad=0 pd=0 as=0 ps=0 
M2691 Vdd Vdd Vdd GND efet w=180 l=480
+ ad=0 pd=0 as=0 ps=0 
M2692 Vdd Vdd diff_49680_79800# GND efet w=720 l=6720
+ ad=0 pd=0 as=0 ps=0 
M2693 Vdd Vdd Vdd GND efet w=180 l=360
+ ad=0 pd=0 as=0 ps=0 
M2694 Vdd Vdd Vdd GND efet w=180 l=540
+ ad=0 pd=0 as=0 ps=0 
M2695 diff_26040_78600# Vdd Vdd GND efet w=960 l=1800
+ ad=9.5184e+06 pd=21360 as=0 ps=0 
M2696 diff_40680_69240# diff_48000_61440# Vdd GND efet w=840 l=840
+ ad=9.8352e+06 pd=24000 as=0 ps=0 
M2697 diff_40680_69240# diff_48000_61440# diff_40680_69240# GND efet w=4620 l=2340
+ ad=0 pd=0 as=0 ps=0 
M2698 diff_48000_61440# Vdd Vdd GND efet w=840 l=720
+ ad=1.8e+06 pd=5760 as=0 ps=0 
M2699 Vdd Vdd diff_33960_53280# GND efet w=840 l=1800
+ ad=0 pd=0 as=1.39104e+07 ps=29280 
M2700 diff_26040_78600# diff_33960_53280# GND GND efet w=8640 l=720
+ ad=0 pd=0 as=0 ps=0 
M2701 GND clk2 diff_40680_69240# GND efet w=4560 l=720
+ ad=0 pd=0 as=0 ps=0 
M2702 Vdd Vdd Vdd GND efet w=300 l=360
+ ad=0 pd=0 as=0 ps=0 
M2703 reset GND reset GND efet w=18240 l=11280
+ ad=3.5784e+07 pd=87360 as=0 ps=0 
M2704 diff_33960_53280# reset GND GND efet w=14460 l=660
+ ad=0 pd=0 as=0 ps=0 
M2705 Vdd Vdd Vdd GND efet w=180 l=240
+ ad=0 pd=0 as=0 ps=0 
M2706 sync clk2 diff_28440_46560# GND efet w=1200 l=720
+ ad=0 pd=0 as=1.8144e+06 ps=6000 
M2707 diff_28440_46560# diff_28440_46560# diff_28440_46560# GND efet w=240 l=420
+ ad=0 pd=0 as=0 ps=0 
M2708 diff_28440_46560# diff_28440_46560# diff_28440_46560# GND efet w=120 l=480
+ ad=0 pd=0 as=0 ps=0 
M2709 GND diff_28440_46560# diff_28920_45720# GND efet w=4020 l=660
+ ad=0 pd=0 as=1.11456e+07 ps=29520 
M2710 Vdd Vdd Vdd GND efet w=60 l=180
+ ad=0 pd=0 as=0 ps=0 
M2711 Vdd Vdd diff_40920_47640# GND efet w=900 l=3540
+ ad=0 pd=0 as=3.7584e+06 ps=10080 
M2712 Vdd Vdd diff_49080_50040# GND efet w=840 l=6480
+ ad=0 pd=0 as=4.1904e+06 ps=9840 
M2713 diff_15480_82200# diff_69480_76200# GND GND efet w=1680 l=720
+ ad=0 pd=0 as=0 ps=0 
M2714 diff_15480_82200# Vdd Vdd GND efet w=720 l=3360
+ ad=0 pd=0 as=0 ps=0 
M2715 Vdd Vdd Vdd GND efet w=120 l=360
+ ad=0 pd=0 as=0 ps=0 
M2716 Vdd Vdd Vdd GND efet w=120 l=240
+ ad=0 pd=0 as=0 ps=0 
M2717 diff_69600_78240# Vdd Vdd GND efet w=720 l=5040
+ ad=0 pd=0 as=0 ps=0 
M2718 diff_70080_67920# diff_33840_37560# GND GND efet w=1200 l=720
+ ad=0 pd=0 as=0 ps=0 
M2719 diff_70080_67920# diff_70080_67920# diff_70080_67920# GND efet w=180 l=180
+ ad=0 pd=0 as=0 ps=0 
M2720 diff_70080_67920# diff_70080_67920# diff_70080_67920# GND efet w=60 l=180
+ ad=0 pd=0 as=0 ps=0 
M2721 diff_90480_76920# Vdd Vdd GND efet w=720 l=5160
+ ad=5.8464e+06 pd=17520 as=0 ps=0 
M2722 GND d3 diff_90480_76920# GND efet w=2880 l=660
+ ad=0 pd=0 as=0 ps=0 
M2723 diff_100800_77520# diff_100440_76920# diff_100800_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2724 diff_102480_84960# diff_100440_76920# diff_102840_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2725 diff_104880_77520# diff_100440_76920# diff_104880_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2726 diff_106920_77520# diff_100440_76920# diff_106920_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2727 diff_108960_77520# diff_100440_76920# diff_108960_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2728 diff_111000_77520# diff_100440_76920# diff_111000_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2729 diff_113040_77520# diff_100440_76920# diff_113040_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2730 diff_115080_77520# diff_100440_76920# diff_115080_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2731 diff_117120_77520# diff_100440_76920# diff_117120_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2732 diff_119160_77520# diff_100440_76920# diff_119160_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2733 diff_121200_77520# diff_100440_76920# diff_121200_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2734 diff_123240_77520# diff_100440_76920# diff_123240_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2735 diff_125280_77520# diff_100440_76920# diff_125280_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2736 diff_127320_77520# diff_100440_76920# diff_127320_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2737 diff_129360_77520# diff_100440_76920# diff_129360_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2738 diff_131400_77520# diff_100440_76920# diff_131400_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2739 diff_133440_77520# diff_100440_76920# diff_133440_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2740 diff_135480_77520# diff_100440_76920# diff_135480_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2741 diff_137520_77520# diff_100440_76920# diff_137520_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2742 diff_139560_77520# diff_100440_76920# diff_139560_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2743 diff_141600_77520# diff_100440_76920# diff_141600_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2744 diff_143640_77520# diff_100440_76920# diff_143640_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2745 diff_145680_77520# diff_100440_76920# diff_145680_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2746 diff_147720_77520# diff_100440_76920# diff_147720_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2747 diff_149760_77520# diff_100440_76920# diff_149760_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2748 diff_151800_77520# diff_100440_76920# diff_151800_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2749 diff_153840_77520# diff_100440_76920# diff_153840_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2750 diff_155880_77520# diff_100440_76920# diff_155880_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2751 diff_157920_77520# diff_100440_76920# diff_157920_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2752 diff_159960_77520# diff_100440_76920# diff_159960_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2753 diff_162000_77520# diff_100440_76920# diff_162000_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2754 diff_164040_77520# diff_100440_76920# diff_164040_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2755 diff_166080_77520# diff_100440_76920# diff_166080_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2756 diff_168120_77520# diff_100440_76920# diff_168120_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2757 diff_170160_77520# diff_100440_76920# diff_170160_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2758 diff_172200_77520# diff_100440_76920# diff_172200_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2759 diff_174240_77520# diff_100440_76920# diff_174240_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2760 diff_176280_77520# diff_100440_76920# diff_176280_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2761 diff_178320_77520# diff_100440_76920# diff_178320_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2762 diff_180360_77520# diff_100440_76920# diff_180360_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2763 diff_182400_77520# diff_100440_76920# diff_182400_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2764 diff_184440_77520# diff_100440_76920# diff_184440_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2765 diff_186480_77520# diff_100440_76920# diff_186480_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2766 diff_188520_77520# diff_100440_76920# diff_188520_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2767 diff_190560_77520# diff_100440_76920# diff_190560_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2768 diff_192600_77520# diff_100440_76920# diff_192600_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2769 diff_194640_77520# diff_100440_76920# diff_194640_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2770 diff_196680_77520# diff_100440_76920# diff_196680_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2771 diff_198720_77520# diff_100440_76920# diff_198720_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2772 diff_200760_77520# diff_100440_76920# diff_200760_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2773 diff_202800_77520# diff_100440_76920# diff_202800_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2774 diff_204840_77520# diff_100440_76920# diff_204840_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2775 diff_206880_77520# diff_100440_76920# diff_206880_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2776 diff_208920_77520# diff_100440_76920# diff_208920_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2777 diff_210960_77520# diff_100440_76920# diff_210960_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2778 diff_213000_77520# diff_100440_76920# diff_213000_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2779 diff_215040_77520# diff_100440_76920# diff_215040_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2780 diff_217080_77520# diff_100440_76920# diff_217080_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2781 diff_219120_77520# diff_100440_76920# diff_219120_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2782 diff_221160_77520# diff_100440_76920# diff_221160_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2783 diff_223200_77520# diff_100440_76920# diff_223200_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2784 diff_225240_77520# diff_100440_76920# diff_225240_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2785 diff_227280_77520# diff_100440_76920# diff_227280_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2786 diff_229320_77520# diff_100440_76920# diff_229320_75240# GND efet w=1080 l=720
+ ad=1.1376e+06 pd=4320 as=1.6848e+06 ps=5280 
M2787 GND diff_252600_124320# diff_243120_97920# GND efet w=12240 l=600
+ ad=0 pd=0 as=1.69776e+07 ps=33120 
M2788 Vdd Vdd diff_112440_115320# GND efet w=720 l=1440
+ ad=0 pd=0 as=0 ps=0 
M2789 Vdd Vdd diff_243120_97920# GND efet w=720 l=1440
+ ad=0 pd=0 as=0 ps=0 
M2790 diff_273840_122880# diff_272280_84480# diff_253080_120120# GND efet w=1920 l=600
+ ad=5.8752e+06 pd=13920 as=2.736e+06 ps=6720 
M2791 Vdd Vdd diff_112440_96360# GND efet w=720 l=1440
+ ad=0 pd=0 as=1.77552e+07 ps=32160 
M2792 diff_112440_96360# diff_253080_120120# GND GND efet w=12240 l=600
+ ad=0 pd=0 as=0 ps=0 
M2793 GND diff_253080_117840# diff_236160_42720# GND efet w=12240 l=600
+ ad=0 pd=0 as=2.0016e+07 ps=33120 
M2794 Vdd Vdd diff_236160_42720# GND efet w=720 l=1440
+ ad=0 pd=0 as=0 ps=0 
M2795 Vdd Vdd diff_238440_42720# GND efet w=720 l=1440
+ ad=0 pd=0 as=1.99008e+07 ps=32640 
M2796 diff_277440_130800# Vdd Vdd GND efet w=840 l=3360
+ ad=0 pd=0 as=0 ps=0 
M2797 diff_281880_129240# diff_281280_113400# diff_277440_130800# GND efet w=3600 l=600
+ ad=3.456e+06 pd=9120 as=0 ps=0 
M2798 GND diff_282840_127320# diff_281880_129240# GND efet w=3600 l=600
+ ad=0 pd=0 as=0 ps=0 
M2799 Vdd Vdd Vdd GND efet w=120 l=240
+ ad=0 pd=0 as=0 ps=0 
M2800 Vdd Vdd Vdd GND efet w=120 l=240
+ ad=0 pd=0 as=0 ps=0 
M2801 Vdd Vdd diff_277440_118920# GND efet w=840 l=3360
+ ad=0 pd=0 as=1.1808e+07 ps=21120 
M2802 diff_273840_122880# diff_271080_135600# diff_253080_117840# GND efet w=2160 l=600
+ ad=0 pd=0 as=3.3408e+06 ps=7440 
M2803 diff_277440_118920# clk2 diff_273840_122880# GND efet w=2160 l=600
+ ad=0 pd=0 as=0 ps=0 
M2804 diff_284160_122760# diff_282840_127320# diff_277440_118920# GND efet w=3480 l=600
+ ad=3.3408e+06 pd=8880 as=0 ps=0 
M2805 GND diff_281280_100320# diff_284160_122760# GND efet w=3480 l=600
+ ad=0 pd=0 as=0 ps=0 
M2806 GND diff_282840_108600# diff_281880_113640# GND efet w=3600 l=600
+ ad=0 pd=0 as=9.8784e+06 ps=19920 
M2807 diff_273840_111480# diff_271080_135600# diff_253080_113280# GND efet w=1920 l=600
+ ad=5.6592e+06 pd=13680 as=2.736e+06 ps=6720 
M2808 diff_277440_115320# clk2 diff_273840_111480# GND efet w=1920 l=600
+ ad=8.9568e+06 pd=15360 as=0 ps=0 
M2809 diff_238440_42720# diff_253080_113280# GND GND efet w=12240 l=600
+ ad=0 pd=0 as=0 ps=0 
M2810 GND diff_253200_111120# diff_101160_115320# GND efet w=12240 l=600
+ ad=0 pd=0 as=1.88064e+07 ps=32400 
M2811 diff_273840_111480# diff_272280_84480# diff_253200_111120# GND efet w=2040 l=600
+ ad=0 pd=0 as=2.9088e+06 ps=6960 
M2812 Vdd Vdd diff_101160_115320# GND efet w=720 l=1440
+ ad=0 pd=0 as=0 ps=0 
M2813 diff_273840_107760# diff_272280_84480# diff_253080_105840# GND efet w=1920 l=600
+ ad=5.5008e+06 pd=13440 as=2.736e+06 ps=6720 
M2814 Vdd Vdd diff_101400_96240# GND efet w=720 l=1440
+ ad=0 pd=0 as=1.90944e+07 ps=32400 
M2815 diff_101400_96240# diff_253080_105840# GND GND efet w=12240 l=600
+ ad=0 pd=0 as=0 ps=0 
M2816 GND diff_253080_103560# diff_241320_99600# GND efet w=12240 l=600
+ ad=0 pd=0 as=1.94256e+07 ps=32400 
M2817 Vdd Vdd diff_241320_99600# GND efet w=720 l=1440
+ ad=0 pd=0 as=0 ps=0 
M2818 Vdd Vdd diff_246960_91200# GND efet w=720 l=1440
+ ad=0 pd=0 as=1.9512e+07 ps=32640 
M2819 diff_246960_91200# diff_253080_99120# GND GND efet w=12240 l=600
+ ad=0 pd=0 as=0 ps=0 
M2820 GND diff_253080_96840# diff_103320_91920# GND efet w=12240 l=600
+ ad=0 pd=0 as=1.85184e+07 ps=32640 
M2821 diff_277440_115320# Vdd Vdd GND efet w=720 l=3360
+ ad=0 pd=0 as=0 ps=0 
M2822 diff_281880_113640# diff_281280_113400# diff_277440_115320# GND efet w=3600 l=600
+ ad=0 pd=0 as=0 ps=0 
M2823 diff_286560_112440# diff_281280_100320# diff_277440_104040# GND efet w=3720 l=600
+ ad=4.0176e+06 pd=9600 as=1.18656e+07 ps=21600 
M2824 GND diff_282840_108600# diff_286560_112440# GND efet w=3720 l=600
+ ad=0 pd=0 as=0 ps=0 
M2825 Vdd Vdd Vdd GND efet w=180 l=420
+ ad=0 pd=0 as=0 ps=0 
M2826 Vdd Vdd Vdd GND efet w=180 l=420
+ ad=0 pd=0 as=0 ps=0 
M2827 Vdd Vdd diff_277440_104040# GND efet w=720 l=3360
+ ad=0 pd=0 as=0 ps=0 
M2828 diff_273840_107760# diff_271080_135600# diff_253080_103560# GND efet w=1920 l=600
+ ad=0 pd=0 as=2.736e+06 ps=6720 
M2829 diff_277440_104040# clk2 diff_273840_107760# GND efet w=1920 l=600
+ ad=0 pd=0 as=0 ps=0 
M2830 diff_273840_96480# diff_271080_135600# diff_253080_99120# GND efet w=2040 l=600
+ ad=5.8464e+06 pd=13920 as=2.9088e+06 ps=6960 
M2831 diff_277440_100200# clk2 diff_273840_96480# GND efet w=2040 l=600
+ ad=1.188e+07 pd=21600 as=0 ps=0 
M2832 d1 GND d1 GND efet w=17760 l=11160
+ ad=0 pd=0 as=0 ps=0 
M2833 GND diff_282840_108600# diff_283200_107520# GND efet w=6360 l=600
+ ad=0 pd=0 as=6.1056e+06 ps=14640 
M2834 diff_283200_107520# diff_281280_100320# diff_283200_105600# GND efet w=6360 l=600
+ ad=0 pd=0 as=1.92528e+07 ps=35040 
M2835 diff_91920_42120# diff_281280_100320# diff_284880_99240# GND efet w=4680 l=600
+ ad=2.85696e+07 pd=60000 as=4.4928e+06 ps=11280 
M2836 diff_273840_96480# diff_272280_84480# diff_253080_96840# GND efet w=2040 l=600
+ ad=0 pd=0 as=2.9088e+06 ps=6960 
M2837 Vdd Vdd diff_103320_91920# GND efet w=600 l=1440
+ ad=0 pd=0 as=0 ps=0 
M2838 Vdd Vdd diff_106320_94080# GND efet w=600 l=1440
+ ad=0 pd=0 as=1.764e+07 ps=32400 
M2839 diff_273840_92640# diff_272280_84480# diff_252960_91560# GND efet w=2160 l=600
+ ad=6.0048e+06 pd=14160 as=3.0816e+06 ps=7200 
M2840 diff_106320_94080# diff_252960_91560# GND GND efet w=12120 l=600
+ ad=0 pd=0 as=0 ps=0 
M2841 GND diff_252960_89400# diff_245160_97920# GND efet w=12120 l=600
+ ad=0 pd=0 as=1.96272e+07 ps=32400 
M2842 Vdd Vdd diff_245160_97920# GND efet w=840 l=1440
+ ad=0 pd=0 as=0 ps=0 
M2843 Vdd Vdd Vdd GND efet w=600 l=480
+ ad=0 pd=0 as=0 ps=0 
M2844 diff_100800_75240# diff_100440_74640# diff_100800_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2845 diff_102840_75240# diff_100440_74640# diff_102840_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2846 diff_104880_75240# diff_100440_74640# diff_104880_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2847 diff_106920_75240# diff_100440_74640# diff_106920_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2848 diff_108960_75240# diff_100440_74640# diff_108960_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2849 diff_111000_75240# diff_100440_74640# diff_111000_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2850 diff_113040_75240# diff_100440_74640# diff_113040_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2851 diff_115080_75240# diff_100440_74640# diff_115080_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2852 diff_117120_75240# diff_100440_74640# diff_117120_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2853 diff_119160_75240# diff_100440_74640# diff_119160_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2854 diff_121200_75240# diff_100440_74640# diff_121200_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2855 diff_123240_75240# diff_100440_74640# diff_123240_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2856 diff_125280_75240# diff_100440_74640# diff_125280_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2857 diff_127320_75240# diff_100440_74640# diff_127320_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2858 diff_129360_75240# diff_100440_74640# diff_129360_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2859 diff_131400_75240# diff_100440_74640# diff_131400_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2860 diff_133440_75240# diff_100440_74640# diff_133440_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2861 diff_135480_75240# diff_100440_74640# diff_135480_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2862 diff_137520_75240# diff_100440_74640# diff_137520_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2863 diff_139560_75240# diff_100440_74640# diff_139560_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2864 diff_141600_75240# diff_100440_74640# diff_141600_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2865 diff_143640_75240# diff_100440_74640# diff_143640_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2866 diff_145680_75240# diff_100440_74640# diff_145680_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2867 diff_147720_75240# diff_100440_74640# diff_147720_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2868 diff_149760_75240# diff_100440_74640# diff_149760_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2869 diff_151800_75240# diff_100440_74640# diff_151800_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2870 diff_153840_75240# diff_100440_74640# diff_153840_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2871 diff_155880_75240# diff_100440_74640# diff_155880_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2872 diff_157920_75240# diff_100440_74640# diff_157920_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2873 diff_159960_75240# diff_100440_74640# diff_159960_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2874 diff_162000_75240# diff_100440_74640# diff_162000_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2875 diff_164040_75240# diff_100440_74640# diff_164040_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2876 diff_166080_75240# diff_100440_74640# diff_166080_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2877 diff_168120_75240# diff_100440_74640# diff_168120_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2878 diff_170160_75240# diff_100440_74640# diff_170160_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2879 diff_172200_75240# diff_100440_74640# diff_172200_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2880 diff_174240_75240# diff_100440_74640# diff_174240_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2881 diff_176280_75240# diff_100440_74640# diff_176280_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2882 diff_178320_75240# diff_100440_74640# diff_178320_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2883 diff_180360_75240# diff_100440_74640# diff_180360_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2884 diff_182400_75240# diff_100440_74640# diff_182400_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2885 diff_184440_75240# diff_100440_74640# diff_184440_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2886 diff_186480_75240# diff_100440_74640# diff_186480_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2887 diff_188520_75240# diff_100440_74640# diff_188520_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2888 diff_190560_75240# diff_100440_74640# diff_190560_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2889 diff_192600_75240# diff_100440_74640# diff_192600_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2890 diff_194640_75240# diff_100440_74640# diff_194640_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2891 diff_196680_75240# diff_100440_74640# diff_196680_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2892 diff_198720_75240# diff_100440_74640# diff_198720_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2893 diff_200760_75240# diff_100440_74640# diff_200760_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2894 diff_202800_75240# diff_100440_74640# diff_202800_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2895 diff_204840_75240# diff_100440_74640# diff_204840_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2896 diff_206880_75240# diff_100440_74640# diff_206880_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2897 diff_208920_75240# diff_100440_74640# diff_208920_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2898 diff_210960_75240# diff_100440_74640# diff_210960_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2899 diff_213000_75240# diff_100440_74640# diff_213000_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2900 diff_215040_75240# diff_100440_74640# diff_215040_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2901 diff_217080_75240# diff_100440_74640# diff_217080_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2902 diff_219120_75240# diff_100440_74640# diff_219120_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2903 diff_221160_75240# diff_100440_74640# diff_221160_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2904 diff_223200_75240# diff_100440_74640# diff_223200_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2905 diff_225240_75240# diff_100440_74640# diff_225240_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2906 diff_227280_75240# diff_100440_74640# diff_227280_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2907 diff_229320_75240# diff_100440_74640# diff_229320_73080# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2908 diff_100440_76920# Vdd Vdd GND efet w=600 l=1320
+ ad=9.4032e+06 pd=26160 as=0 ps=0 
M2909 Vdd Vdd Vdd GND efet w=240 l=600
+ ad=0 pd=0 as=0 ps=0 
M2910 Vdd Vdd Vdd GND efet w=120 l=480
+ ad=0 pd=0 as=0 ps=0 
M2911 diff_86640_69120# Vdd Vdd GND efet w=720 l=5040
+ ad=6.2064e+06 pd=14880 as=0 ps=0 
M2912 diff_41160_86760# diff_84000_37560# GND GND efet w=2160 l=600
+ ad=0 pd=0 as=0 ps=0 
M2913 GND diff_86640_69120# diff_41160_86760# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2914 diff_100800_73080# diff_100440_72480# diff_100800_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2915 diff_102840_73080# diff_100440_72480# diff_102840_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2916 diff_104880_73080# diff_100440_72480# diff_104880_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2917 diff_106920_73080# diff_100440_72480# diff_106920_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2918 diff_108960_73080# diff_100440_72480# diff_108960_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2919 diff_111000_73080# diff_100440_72480# diff_111000_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2920 diff_113040_73080# diff_100440_72480# diff_113040_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2921 diff_115080_73080# diff_100440_72480# diff_115080_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2922 diff_117120_73080# diff_100440_72480# diff_117120_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2923 diff_119160_73080# diff_100440_72480# diff_119160_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2924 diff_121200_73080# diff_100440_72480# diff_121200_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2925 diff_123240_73080# diff_100440_72480# diff_123240_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2926 diff_125280_73080# diff_100440_72480# diff_125280_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2927 diff_127320_73080# diff_100440_72480# diff_127320_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2928 diff_129360_73080# diff_100440_72480# diff_129360_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2929 diff_131400_73080# diff_100440_72480# diff_131400_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2930 diff_133440_73080# diff_100440_72480# diff_133440_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2931 diff_135480_73080# diff_100440_72480# diff_135480_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2932 diff_137520_73080# diff_100440_72480# diff_137520_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2933 diff_139560_73080# diff_100440_72480# diff_139560_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2934 diff_141600_73080# diff_100440_72480# diff_141600_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2935 diff_143640_73080# diff_100440_72480# diff_143640_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2936 diff_145680_73080# diff_100440_72480# diff_145680_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2937 diff_147720_73080# diff_100440_72480# diff_147720_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2938 diff_149760_73080# diff_100440_72480# diff_149760_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2939 diff_151800_73080# diff_100440_72480# diff_151800_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2940 diff_153840_73080# diff_100440_72480# diff_153840_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2941 diff_155880_73080# diff_100440_72480# diff_155880_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2942 diff_157920_73080# diff_100440_72480# diff_157920_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2943 diff_159960_73080# diff_100440_72480# diff_159960_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2944 diff_162000_73080# diff_100440_72480# diff_162000_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2945 diff_164040_73080# diff_100440_72480# diff_164040_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2946 diff_166080_73080# diff_100440_72480# diff_166080_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2947 diff_168120_73080# diff_100440_72480# diff_168120_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2948 diff_170160_73080# diff_100440_72480# diff_170160_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2949 diff_172200_73080# diff_100440_72480# diff_172200_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2950 diff_174240_73080# diff_100440_72480# diff_174240_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2951 diff_176280_73080# diff_100440_72480# diff_176280_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2952 diff_178320_73080# diff_100440_72480# diff_178320_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2953 diff_180360_73080# diff_100440_72480# diff_180360_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2954 diff_182400_73080# diff_100440_72480# diff_182400_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2955 diff_184440_73080# diff_100440_72480# diff_184440_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2956 diff_186480_73080# diff_100440_72480# diff_186480_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2957 diff_188520_73080# diff_100440_72480# diff_188520_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2958 diff_190560_73080# diff_100440_72480# diff_190560_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2959 diff_192600_73080# diff_100440_72480# diff_192600_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2960 diff_194640_73080# diff_100440_72480# diff_194640_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2961 diff_196680_73080# diff_100440_72480# diff_196680_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2962 diff_198720_73080# diff_100440_72480# diff_198720_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2963 diff_200760_73080# diff_100440_72480# diff_200760_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2964 diff_202800_73080# diff_100440_72480# diff_202800_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2965 diff_204840_73080# diff_100440_72480# diff_204840_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2966 diff_206880_73080# diff_100440_72480# diff_206880_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2967 diff_208920_73080# diff_100440_72480# diff_208920_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2968 diff_210960_73080# diff_100440_72480# diff_210960_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2969 diff_213000_73080# diff_100440_72480# diff_213000_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2970 diff_215040_73080# diff_100440_72480# diff_215040_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2971 diff_217080_73080# diff_100440_72480# diff_217080_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2972 diff_219120_73080# diff_100440_72480# diff_219120_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2973 diff_221160_73080# diff_100440_72480# diff_221160_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2974 diff_223200_73080# diff_100440_72480# diff_223200_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2975 diff_225240_73080# diff_100440_72480# diff_225240_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2976 diff_227280_73080# diff_100440_72480# diff_227280_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2977 diff_229320_73080# diff_100440_72480# diff_229320_70800# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M2978 Vdd Vdd diff_100440_70200# GND efet w=600 l=1200
+ ad=0 pd=0 as=8.7264e+06 ps=22800 
M2979 diff_236760_69600# diff_236160_42720# diff_100440_70200# GND efet w=8640 l=600
+ ad=3.64608e+07 pd=72720 as=0 ps=0 
M2980 diff_86640_69120# diff_86640_69120# diff_86640_69120# GND efet w=180 l=240
+ ad=0 pd=0 as=0 ps=0 
M2981 diff_86640_69120# diff_86640_69120# diff_86640_69120# GND efet w=240 l=240
+ ad=0 pd=0 as=0 ps=0 
M2982 GND diff_90480_65640# diff_86640_69120# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M2983 diff_100800_70800# diff_100440_70200# diff_100800_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2984 diff_102840_70800# diff_100440_70200# diff_102840_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2985 diff_104880_70800# diff_100440_70200# diff_104880_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2986 diff_106920_70800# diff_100440_70200# diff_106920_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2987 diff_108960_70800# diff_100440_70200# diff_108960_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2988 diff_111000_70800# diff_100440_70200# diff_111000_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2989 diff_113040_70800# diff_100440_70200# diff_113040_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2990 diff_115080_70800# diff_100440_70200# diff_115080_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2991 diff_117120_70800# diff_100440_70200# diff_117120_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2992 diff_119160_70800# diff_100440_70200# diff_119160_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2993 diff_121200_70800# diff_100440_70200# diff_121200_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2994 diff_123240_70800# diff_100440_70200# diff_123240_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2995 diff_125280_70800# diff_100440_70200# diff_125280_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2996 diff_127320_70800# diff_100440_70200# diff_127320_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2997 diff_129360_70800# diff_100440_70200# diff_129360_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2998 diff_131400_70800# diff_100440_70200# diff_131400_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M2999 diff_133440_70800# diff_100440_70200# diff_133440_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3000 diff_135480_70800# diff_100440_70200# diff_135480_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3001 diff_137520_70800# diff_100440_70200# diff_137520_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3002 diff_139560_70800# diff_100440_70200# diff_139560_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3003 diff_141600_70800# diff_100440_70200# diff_141600_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3004 diff_143640_70800# diff_100440_70200# diff_143640_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3005 diff_145680_70800# diff_100440_70200# diff_145680_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3006 diff_147720_70800# diff_100440_70200# diff_147720_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3007 diff_149760_70800# diff_100440_70200# diff_149760_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3008 diff_151800_70800# diff_100440_70200# diff_151800_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3009 diff_153840_70800# diff_100440_70200# diff_153840_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3010 diff_155880_70800# diff_100440_70200# diff_155880_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3011 diff_157920_70800# diff_100440_70200# diff_157920_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3012 diff_159960_70800# diff_100440_70200# diff_159960_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3013 diff_162000_70800# diff_100440_70200# diff_162000_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3014 diff_164040_70800# diff_100440_70200# diff_164040_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3015 diff_166080_70800# diff_100440_70200# diff_166080_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3016 diff_168120_70800# diff_100440_70200# diff_168120_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3017 diff_170160_70800# diff_100440_70200# diff_170160_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3018 diff_172200_70800# diff_100440_70200# diff_172200_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3019 diff_174240_70800# diff_100440_70200# diff_174240_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3020 diff_176280_70800# diff_100440_70200# diff_176280_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3021 diff_178320_70800# diff_100440_70200# diff_178320_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3022 diff_180360_70800# diff_100440_70200# diff_180360_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3023 diff_182400_70800# diff_100440_70200# diff_182400_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3024 diff_184440_70800# diff_100440_70200# diff_184440_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3025 diff_186480_70800# diff_100440_70200# diff_186480_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3026 diff_188520_70800# diff_100440_70200# diff_188520_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3027 diff_190560_70800# diff_100440_70200# diff_190560_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3028 diff_192600_70800# diff_100440_70200# diff_192600_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3029 diff_194640_70800# diff_100440_70200# diff_194640_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3030 diff_196680_70800# diff_100440_70200# diff_196680_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3031 diff_198720_70800# diff_100440_70200# diff_198720_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3032 diff_200760_70800# diff_100440_70200# diff_200760_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3033 diff_202800_70800# diff_100440_70200# diff_202800_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3034 diff_204840_70800# diff_100440_70200# diff_204840_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3035 diff_206880_70800# diff_100440_70200# diff_206880_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3036 diff_208920_70800# diff_100440_70200# diff_208920_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3037 diff_210960_70800# diff_100440_70200# diff_210960_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3038 diff_213000_70800# diff_100440_70200# diff_213000_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3039 diff_215040_70800# diff_100440_70200# diff_215040_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3040 diff_217080_70800# diff_100440_70200# diff_217080_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3041 diff_219120_70800# diff_100440_70200# diff_219120_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3042 diff_221160_70800# diff_100440_70200# diff_221160_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3043 diff_223200_70800# diff_100440_70200# diff_223200_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3044 diff_225240_70800# diff_100440_70200# diff_225240_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3045 diff_227280_70800# diff_100440_70200# diff_227280_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3046 diff_229320_70800# diff_100440_70200# diff_229320_68640# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3047 diff_100440_76920# diff_238440_42720# diff_236760_69600# GND efet w=7440 l=600
+ ad=0 pd=0 as=0 ps=0 
M3048 diff_100440_74640# Vdd Vdd GND efet w=720 l=1320
+ ad=1.0368e+07 pd=24960 as=0 ps=0 
M3049 Vdd Vdd diff_100440_72480# GND efet w=720 l=1080
+ ad=0 pd=0 as=1.05264e+07 ps=22560 
M3050 diff_236760_69600# diff_241320_99600# diff_100440_72480# GND efet w=8520 l=600
+ ad=0 pd=0 as=0 ps=0 
M3051 diff_100800_68640# diff_100440_68040# diff_100800_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3052 diff_102840_68640# diff_100440_68040# diff_102840_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3053 diff_104880_68640# diff_100440_68040# diff_104880_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3054 diff_106920_68640# diff_100440_68040# diff_106920_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3055 diff_108960_68640# diff_100440_68040# diff_108960_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3056 diff_111000_68640# diff_100440_68040# diff_111000_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3057 diff_113040_68640# diff_100440_68040# diff_113040_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3058 diff_115080_68640# diff_100440_68040# diff_115080_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3059 diff_117120_68640# diff_100440_68040# diff_117120_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3060 diff_119160_68640# diff_100440_68040# diff_119160_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3061 diff_121200_68640# diff_100440_68040# diff_121200_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3062 diff_123240_68640# diff_100440_68040# diff_123240_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3063 diff_125280_68640# diff_100440_68040# diff_125280_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3064 diff_127320_68640# diff_100440_68040# diff_127320_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3065 diff_129360_68640# diff_100440_68040# diff_129360_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3066 diff_131400_68640# diff_100440_68040# diff_131400_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3067 diff_133440_68640# diff_100440_68040# diff_133440_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3068 diff_135480_68640# diff_100440_68040# diff_135480_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3069 diff_137520_68640# diff_100440_68040# diff_137520_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3070 diff_139560_68640# diff_100440_68040# diff_139560_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3071 diff_141600_68640# diff_100440_68040# diff_141600_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3072 diff_143640_68640# diff_100440_68040# diff_143640_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3073 diff_145680_68640# diff_100440_68040# diff_145680_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3074 diff_147720_68640# diff_100440_68040# diff_147720_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3075 diff_149760_68640# diff_100440_68040# diff_149760_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3076 diff_151800_68640# diff_100440_68040# diff_151800_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3077 diff_153840_68640# diff_100440_68040# diff_153840_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3078 diff_155880_68640# diff_100440_68040# diff_155880_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3079 diff_157920_68640# diff_100440_68040# diff_157920_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3080 diff_159960_68640# diff_100440_68040# diff_159960_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3081 diff_162000_68640# diff_100440_68040# diff_162000_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3082 diff_164040_68640# diff_100440_68040# diff_164040_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3083 diff_166080_68640# diff_100440_68040# diff_166080_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3084 diff_168120_68640# diff_100440_68040# diff_168120_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3085 diff_170160_68640# diff_100440_68040# diff_170160_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3086 diff_172200_68640# diff_100440_68040# diff_172200_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3087 diff_174240_68640# diff_100440_68040# diff_174240_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3088 diff_176280_68640# diff_100440_68040# diff_176280_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3089 diff_178320_68640# diff_100440_68040# diff_178320_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3090 diff_180360_68640# diff_100440_68040# diff_180360_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3091 diff_182400_68640# diff_100440_68040# diff_182400_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3092 diff_184440_68640# diff_100440_68040# diff_184440_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3093 diff_186480_68640# diff_100440_68040# diff_186480_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3094 diff_188520_68640# diff_100440_68040# diff_188520_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3095 diff_190560_68640# diff_100440_68040# diff_190560_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3096 diff_192600_68640# diff_100440_68040# diff_192600_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3097 diff_194640_68640# diff_100440_68040# diff_194640_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3098 diff_196680_68640# diff_100440_68040# diff_196680_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3099 diff_198720_68640# diff_100440_68040# diff_198720_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3100 diff_200760_68640# diff_100440_68040# diff_200760_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3101 diff_202800_68640# diff_100440_68040# diff_202800_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3102 diff_204840_68640# diff_100440_68040# diff_204840_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3103 diff_206880_68640# diff_100440_68040# diff_206880_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3104 diff_208920_68640# diff_100440_68040# diff_208920_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3105 diff_210960_68640# diff_100440_68040# diff_210960_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3106 diff_213000_68640# diff_100440_68040# diff_213000_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3107 diff_215040_68640# diff_100440_68040# diff_215040_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3108 diff_217080_68640# diff_100440_68040# diff_217080_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3109 diff_219120_68640# diff_100440_68040# diff_219120_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3110 diff_221160_68640# diff_100440_68040# diff_221160_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3111 diff_223200_68640# diff_100440_68040# diff_223200_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3112 diff_225240_68640# diff_100440_68040# diff_225240_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3113 diff_227280_68640# diff_100440_68040# diff_227280_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3114 diff_229320_68640# diff_100440_68040# diff_229320_66360# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3115 diff_100440_74640# diff_243120_97920# diff_236760_69600# GND efet w=7920 l=600
+ ad=0 pd=0 as=0 ps=0 
M3116 diff_236760_60720# diff_236160_42720# diff_100440_61320# GND efet w=8820 l=720
+ ad=4.0536e+07 pd=72000 as=8.4672e+06 ps=22800 
M3117 diff_89160_65640# clk2 Vdd GND efet w=1200 l=720
+ ad=720000 pd=3600 as=0 ps=0 
M3118 diff_90480_65640# diff_89760_63840# diff_89160_65640# GND efet w=1200 l=720
+ ad=4.608e+06 pd=10080 as=0 ps=0 
M3119 GND diff_33840_37560# diff_90480_65640# GND efet w=1200 l=720
+ ad=0 pd=0 as=0 ps=0 
M3120 diff_100800_66360# diff_100440_65760# diff_100800_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3121 diff_102840_66360# diff_100440_65760# diff_102840_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3122 diff_104880_66360# diff_100440_65760# diff_104880_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3123 diff_106920_66360# diff_100440_65760# diff_106920_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3124 diff_108960_66360# diff_100440_65760# diff_108960_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3125 diff_111000_66360# diff_100440_65760# diff_111000_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3126 diff_113040_66360# diff_100440_65760# diff_113040_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3127 diff_115080_66360# diff_100440_65760# diff_115080_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3128 diff_117120_66360# diff_100440_65760# diff_117120_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3129 diff_119160_66360# diff_100440_65760# diff_119160_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3130 diff_121200_66360# diff_100440_65760# diff_121200_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3131 diff_123240_66360# diff_100440_65760# diff_123240_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3132 diff_125280_66360# diff_100440_65760# diff_125280_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3133 diff_127320_66360# diff_100440_65760# diff_127320_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3134 diff_129360_66360# diff_100440_65760# diff_129360_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3135 diff_131400_66360# diff_100440_65760# diff_131400_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3136 diff_133440_66360# diff_100440_65760# diff_133440_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3137 diff_135480_66360# diff_100440_65760# diff_135480_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3138 diff_137520_66360# diff_100440_65760# diff_137520_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3139 diff_139560_66360# diff_100440_65760# diff_139560_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3140 diff_141600_66360# diff_100440_65760# diff_141600_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3141 diff_143640_66360# diff_100440_65760# diff_143640_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3142 diff_145680_66360# diff_100440_65760# diff_145680_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3143 diff_147720_66360# diff_100440_65760# diff_147720_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3144 diff_149760_66360# diff_100440_65760# diff_149760_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3145 diff_151800_66360# diff_100440_65760# diff_151800_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3146 diff_153840_66360# diff_100440_65760# diff_153840_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3147 diff_155880_66360# diff_100440_65760# diff_155880_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3148 diff_157920_66360# diff_100440_65760# diff_157920_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3149 diff_159960_66360# diff_100440_65760# diff_159960_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3150 diff_162000_66360# diff_100440_65760# diff_162000_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3151 diff_164040_66360# diff_100440_65760# diff_164040_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3152 diff_166080_66360# diff_100440_65760# diff_166080_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3153 diff_168120_66360# diff_100440_65760# diff_168120_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3154 diff_170160_66360# diff_100440_65760# diff_170160_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3155 diff_172200_66360# diff_100440_65760# diff_172200_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3156 diff_174240_66360# diff_100440_65760# diff_174240_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3157 diff_176280_66360# diff_100440_65760# diff_176280_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3158 diff_178320_66360# diff_100440_65760# diff_178320_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3159 diff_180360_66360# diff_100440_65760# diff_180360_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3160 diff_182400_66360# diff_100440_65760# diff_182400_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3161 diff_184440_66360# diff_100440_65760# diff_184440_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3162 diff_186480_66360# diff_100440_65760# diff_186480_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3163 diff_188520_66360# diff_100440_65760# diff_188520_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3164 diff_190560_66360# diff_100440_65760# diff_190560_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3165 diff_192600_66360# diff_100440_65760# diff_192600_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3166 diff_194640_66360# diff_100440_65760# diff_194640_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3167 diff_196680_66360# diff_100440_65760# diff_196680_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3168 diff_198720_66360# diff_100440_65760# diff_198720_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3169 diff_200760_66360# diff_100440_65760# diff_200760_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3170 diff_202800_66360# diff_100440_65760# diff_202800_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3171 diff_204840_66360# diff_100440_65760# diff_204840_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3172 diff_206880_66360# diff_100440_65760# diff_206880_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3173 diff_208920_66360# diff_100440_65760# diff_208920_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3174 diff_210960_66360# diff_100440_65760# diff_210960_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3175 diff_213000_66360# diff_100440_65760# diff_213000_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3176 diff_215040_66360# diff_100440_65760# diff_215040_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3177 diff_217080_66360# diff_100440_65760# diff_217080_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3178 diff_219120_66360# diff_100440_65760# diff_219120_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3179 diff_221160_66360# diff_100440_65760# diff_221160_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3180 diff_223200_66360# diff_100440_65760# diff_223200_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3181 diff_225240_66360# diff_100440_65760# diff_225240_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3182 diff_227280_66360# diff_100440_65760# diff_227280_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3183 diff_229320_66360# diff_100440_65760# diff_229320_64200# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3184 diff_100440_68040# Vdd Vdd GND efet w=600 l=1320
+ ad=9.4032e+06 pd=26160 as=0 ps=0 
M3185 diff_69480_76200# diff_74640_62520# GND GND efet w=1200 l=720
+ ad=2.4768e+06 pd=6960 as=0 ps=0 
M3186 Vdd Vdd diff_69480_76200# GND efet w=780 l=5100
+ ad=0 pd=0 as=0 ps=0 
M3187 diff_56400_47520# diff_56400_47520# diff_56400_47520# GND efet w=300 l=360
+ ad=1.12032e+07 pd=25680 as=0 ps=0 
M3188 diff_56400_47520# diff_56400_47520# diff_56400_47520# GND efet w=300 l=420
+ ad=0 pd=0 as=0 ps=0 
M3189 Vdd Vdd diff_56400_47520# GND efet w=960 l=1680
+ ad=0 pd=0 as=0 ps=0 
M3190 diff_100800_64200# diff_100440_63600# diff_100800_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3191 diff_102840_64200# diff_100440_63600# diff_102840_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3192 diff_104880_64200# diff_100440_63600# diff_104880_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3193 diff_106920_64200# diff_100440_63600# diff_106920_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3194 diff_108960_64200# diff_100440_63600# diff_108960_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3195 diff_111000_64200# diff_100440_63600# diff_111000_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3196 diff_113040_64200# diff_100440_63600# diff_113040_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3197 diff_115080_64200# diff_100440_63600# diff_115080_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3198 diff_117120_64200# diff_100440_63600# diff_117120_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3199 diff_119160_64200# diff_100440_63600# diff_119160_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3200 diff_121200_64200# diff_100440_63600# diff_121200_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3201 diff_123240_64200# diff_100440_63600# diff_123240_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3202 diff_125280_64200# diff_100440_63600# diff_125280_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3203 diff_127320_64200# diff_100440_63600# diff_127320_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3204 diff_129360_64200# diff_100440_63600# diff_129360_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3205 diff_131400_64200# diff_100440_63600# diff_131400_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3206 diff_133440_64200# diff_100440_63600# diff_133440_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3207 diff_135480_64200# diff_100440_63600# diff_135480_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3208 diff_137520_64200# diff_100440_63600# diff_137520_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3209 diff_139560_64200# diff_100440_63600# diff_139560_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3210 diff_141600_64200# diff_100440_63600# diff_141600_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3211 diff_143640_64200# diff_100440_63600# diff_143640_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3212 diff_145680_64200# diff_100440_63600# diff_145680_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3213 diff_147720_64200# diff_100440_63600# diff_147720_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3214 diff_149760_64200# diff_100440_63600# diff_149760_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3215 diff_151800_64200# diff_100440_63600# diff_151800_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3216 diff_153840_64200# diff_100440_63600# diff_153840_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3217 diff_155880_64200# diff_100440_63600# diff_155880_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3218 diff_157920_64200# diff_100440_63600# diff_157920_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3219 diff_159960_64200# diff_100440_63600# diff_159960_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3220 diff_162000_64200# diff_100440_63600# diff_162000_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3221 diff_164040_64200# diff_100440_63600# diff_164040_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3222 diff_166080_64200# diff_100440_63600# diff_166080_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3223 diff_168120_64200# diff_100440_63600# diff_168120_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3224 diff_170160_64200# diff_100440_63600# diff_170160_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3225 diff_172200_64200# diff_100440_63600# diff_172200_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3226 diff_174240_64200# diff_100440_63600# diff_174240_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3227 diff_176280_64200# diff_100440_63600# diff_176280_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3228 diff_178320_64200# diff_100440_63600# diff_178320_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3229 diff_180360_64200# diff_100440_63600# diff_180360_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3230 diff_182400_64200# diff_100440_63600# diff_182400_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3231 diff_184440_64200# diff_100440_63600# diff_184440_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3232 diff_186480_64200# diff_100440_63600# diff_186480_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3233 diff_188520_64200# diff_100440_63600# diff_188520_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3234 diff_190560_64200# diff_100440_63600# diff_190560_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3235 diff_192600_64200# diff_100440_63600# diff_192600_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3236 diff_194640_64200# diff_100440_63600# diff_194640_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3237 diff_196680_64200# diff_100440_63600# diff_196680_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3238 diff_198720_64200# diff_100440_63600# diff_198720_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3239 diff_200760_64200# diff_100440_63600# diff_200760_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3240 diff_202800_64200# diff_100440_63600# diff_202800_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3241 diff_204840_64200# diff_100440_63600# diff_204840_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3242 diff_206880_64200# diff_100440_63600# diff_206880_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3243 diff_208920_64200# diff_100440_63600# diff_208920_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3244 diff_210960_64200# diff_100440_63600# diff_210960_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3245 diff_213000_64200# diff_100440_63600# diff_213000_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3246 diff_215040_64200# diff_100440_63600# diff_215040_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3247 diff_217080_64200# diff_100440_63600# diff_217080_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3248 diff_219120_64200# diff_100440_63600# diff_219120_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3249 diff_221160_64200# diff_100440_63600# diff_221160_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3250 diff_223200_64200# diff_100440_63600# diff_223200_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3251 diff_225240_64200# diff_100440_63600# diff_225240_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3252 diff_227280_64200# diff_100440_63600# diff_227280_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3253 diff_229320_64200# diff_100440_63600# diff_229320_61920# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3254 Vdd Vdd diff_100440_61320# GND efet w=600 l=1200
+ ad=0 pd=0 as=0 ps=0 
M3255 Vdd Vdd diff_62400_47520# GND efet w=960 l=1680
+ ad=0 pd=0 as=8.5104e+06 ps=18960 
M3256 Vdd Vdd Vdd GND efet w=420 l=420
+ ad=0 pd=0 as=0 ps=0 
M3257 Vdd Vdd diff_69480_55680# GND efet w=720 l=6360
+ ad=0 pd=0 as=8.6256e+06 ps=20880 
M3258 diff_69480_55680# cm diff_69480_49320# GND efet w=7800 l=720
+ ad=0 pd=0 as=7.1424e+06 ps=17280 
M3259 diff_40440_47040# diff_33840_37560# Vdd GND efet w=1320 l=600
+ ad=2.5344e+06 pd=6480 as=0 ps=0 
M3260 diff_47520_50040# clk2 diff_40440_47040# GND efet w=1320 l=720
+ ad=1.1088e+06 pd=4320 as=0 ps=0 
M3261 diff_49080_50040# diff_47880_47040# diff_47520_50040# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M3262 Vdd Vdd diff_69120_48720# GND efet w=840 l=5040
+ ad=0 pd=0 as=1.02096e+07 ps=22080 
M3263 Vdd Vdd diff_75600_45480# GND efet w=720 l=5040
+ ad=0 pd=0 as=4.7808e+06 ps=12960 
M3264 Vdd Vdd Vdd GND efet w=360 l=360
+ ad=0 pd=0 as=0 ps=0 
M3265 diff_89760_63840# Vdd Vdd GND efet w=720 l=3480
+ ad=6.3792e+06 pd=16320 as=0 ps=0 
M3266 GND diff_69480_55680# diff_89760_63840# GND efet w=1800 l=720
+ ad=0 pd=0 as=0 ps=0 
M3267 diff_89760_63840# diff_90480_76920# GND GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M3268 GND diff_91920_42120# diff_89760_63840# GND efet w=1800 l=720
+ ad=0 pd=0 as=0 ps=0 
M3269 diff_100800_61920# diff_100440_61320# diff_100800_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3270 diff_102840_61920# diff_100440_61320# diff_102840_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3271 diff_104880_61920# diff_100440_61320# diff_104880_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3272 diff_106920_61920# diff_100440_61320# diff_106920_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3273 diff_108960_61920# diff_100440_61320# diff_108960_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3274 diff_111000_61920# diff_100440_61320# diff_111000_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3275 diff_113040_61920# diff_100440_61320# diff_113040_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3276 diff_115080_61920# diff_100440_61320# diff_115080_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3277 diff_117120_61920# diff_100440_61320# diff_117120_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3278 diff_119160_61920# diff_100440_61320# diff_119160_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3279 diff_121200_61920# diff_100440_61320# diff_121200_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3280 diff_123240_61920# diff_100440_61320# diff_123240_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3281 diff_125280_61920# diff_100440_61320# diff_125280_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3282 diff_127320_61920# diff_100440_61320# diff_127320_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3283 diff_129360_61920# diff_100440_61320# diff_129360_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3284 diff_131400_61920# diff_100440_61320# diff_131400_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3285 diff_133440_61920# diff_100440_61320# diff_133440_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3286 diff_135480_61920# diff_100440_61320# diff_135480_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3287 diff_137520_61920# diff_100440_61320# diff_137520_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3288 diff_139560_61920# diff_100440_61320# diff_139560_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3289 diff_141600_61920# diff_100440_61320# diff_141600_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3290 diff_143640_61920# diff_100440_61320# diff_143640_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3291 diff_145680_61920# diff_100440_61320# diff_145680_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3292 diff_147720_61920# diff_100440_61320# diff_147720_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3293 diff_149760_61920# diff_100440_61320# diff_149760_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3294 diff_151800_61920# diff_100440_61320# diff_151800_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3295 diff_153840_61920# diff_100440_61320# diff_153840_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3296 diff_155880_61920# diff_100440_61320# diff_155880_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3297 diff_157920_61920# diff_100440_61320# diff_157920_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3298 diff_159960_61920# diff_100440_61320# diff_159960_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3299 diff_162000_61920# diff_100440_61320# diff_162000_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3300 diff_164040_61920# diff_100440_61320# diff_164040_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3301 diff_166080_61920# diff_100440_61320# diff_166080_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3302 diff_168120_61920# diff_100440_61320# diff_168120_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3303 diff_170160_61920# diff_100440_61320# diff_170160_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3304 diff_172200_61920# diff_100440_61320# diff_172200_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3305 diff_174240_61920# diff_100440_61320# diff_174240_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3306 diff_176280_61920# diff_100440_61320# diff_176280_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3307 diff_178320_61920# diff_100440_61320# diff_178320_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3308 diff_180360_61920# diff_100440_61320# diff_180360_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3309 diff_182400_61920# diff_100440_61320# diff_182400_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3310 diff_184440_61920# diff_100440_61320# diff_184440_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3311 diff_186480_61920# diff_100440_61320# diff_186480_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3312 diff_188520_61920# diff_100440_61320# diff_188520_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3313 diff_190560_61920# diff_100440_61320# diff_190560_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3314 diff_192600_61920# diff_100440_61320# diff_192600_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3315 diff_194640_61920# diff_100440_61320# diff_194640_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3316 diff_196680_61920# diff_100440_61320# diff_196680_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3317 diff_198720_61920# diff_100440_61320# diff_198720_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3318 diff_200760_61920# diff_100440_61320# diff_200760_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3319 diff_202800_61920# diff_100440_61320# diff_202800_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3320 diff_204840_61920# diff_100440_61320# diff_204840_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3321 diff_206880_61920# diff_100440_61320# diff_206880_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3322 diff_208920_61920# diff_100440_61320# diff_208920_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3323 diff_210960_61920# diff_100440_61320# diff_210960_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3324 diff_213000_61920# diff_100440_61320# diff_213000_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3325 diff_215040_61920# diff_100440_61320# diff_215040_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3326 diff_217080_61920# diff_100440_61320# diff_217080_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3327 diff_219120_61920# diff_100440_61320# diff_219120_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3328 diff_221160_61920# diff_100440_61320# diff_221160_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3329 diff_223200_61920# diff_100440_61320# diff_223200_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3330 diff_225240_61920# diff_100440_61320# diff_225240_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3331 diff_227280_61920# diff_100440_61320# diff_227280_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3332 diff_229320_61920# diff_100440_61320# diff_229320_59760# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3333 Vdd Vdd diff_81000_51000# GND efet w=720 l=5160
+ ad=0 pd=0 as=6.4368e+06 ps=17280 
M3334 diff_100440_68040# diff_238440_42720# diff_236760_60720# GND efet w=7440 l=600
+ ad=0 pd=0 as=0 ps=0 
M3335 diff_100440_65760# Vdd Vdd GND efet w=720 l=1200
+ ad=1.0368e+07 pd=24960 as=0 ps=0 
M3336 Vdd Vdd diff_100440_63600# GND efet w=720 l=1080
+ ad=0 pd=0 as=1.05984e+07 ps=22560 
M3337 diff_236760_60720# diff_241320_99600# diff_100440_63600# GND efet w=8400 l=600
+ ad=0 pd=0 as=0 ps=0 
M3338 diff_100800_59760# diff_100440_59160# diff_100800_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3339 diff_102840_59760# diff_100440_59160# diff_102840_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3340 diff_104880_59760# diff_100440_59160# diff_104880_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3341 diff_106920_59760# diff_100440_59160# diff_106920_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3342 diff_108960_59760# diff_100440_59160# diff_108960_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3343 diff_111000_59760# diff_100440_59160# diff_111000_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3344 diff_113040_59760# diff_100440_59160# diff_113040_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3345 diff_115080_59760# diff_100440_59160# diff_115080_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3346 diff_117120_59760# diff_100440_59160# diff_117120_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3347 diff_119160_59760# diff_100440_59160# diff_119160_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3348 diff_121200_59760# diff_100440_59160# diff_121200_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3349 diff_123240_59760# diff_100440_59160# diff_123240_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3350 diff_125280_59760# diff_100440_59160# diff_125280_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3351 diff_127320_59760# diff_100440_59160# diff_127320_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3352 diff_129360_59760# diff_100440_59160# diff_129360_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3353 diff_131400_59760# diff_100440_59160# diff_131400_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3354 diff_133440_59760# diff_100440_59160# diff_133440_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3355 diff_135480_59760# diff_100440_59160# diff_135480_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3356 diff_137520_59760# diff_100440_59160# diff_137520_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3357 diff_139560_59760# diff_100440_59160# diff_139560_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3358 diff_141600_59760# diff_100440_59160# diff_141600_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3359 diff_143640_59760# diff_100440_59160# diff_143640_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3360 diff_145680_59760# diff_100440_59160# diff_145680_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3361 diff_147720_59760# diff_100440_59160# diff_147720_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3362 diff_149760_59760# diff_100440_59160# diff_149760_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3363 diff_151800_59760# diff_100440_59160# diff_151800_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3364 diff_153840_59760# diff_100440_59160# diff_153840_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3365 diff_155880_59760# diff_100440_59160# diff_155880_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3366 diff_157920_59760# diff_100440_59160# diff_157920_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3367 diff_159960_59760# diff_100440_59160# diff_159960_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3368 diff_162000_59760# diff_100440_59160# diff_162000_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3369 diff_164040_59760# diff_100440_59160# diff_164040_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3370 diff_166080_59760# diff_100440_59160# diff_166080_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3371 diff_168120_59760# diff_100440_59160# diff_168120_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3372 diff_170160_59760# diff_100440_59160# diff_170160_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3373 diff_172200_59760# diff_100440_59160# diff_172200_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3374 diff_174240_59760# diff_100440_59160# diff_174240_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3375 diff_176280_59760# diff_100440_59160# diff_176280_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3376 diff_178320_59760# diff_100440_59160# diff_178320_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3377 diff_180360_59760# diff_100440_59160# diff_180360_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3378 diff_182400_59760# diff_100440_59160# diff_182400_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3379 diff_184440_59760# diff_100440_59160# diff_184440_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3380 diff_186480_59760# diff_100440_59160# diff_186480_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3381 diff_188520_59760# diff_100440_59160# diff_188520_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3382 diff_190560_59760# diff_100440_59160# diff_190560_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3383 diff_192600_59760# diff_100440_59160# diff_192600_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3384 diff_194640_59760# diff_100440_59160# diff_194640_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3385 diff_196680_59760# diff_100440_59160# diff_196680_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3386 diff_198720_59760# diff_100440_59160# diff_198720_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3387 diff_200760_59760# diff_100440_59160# diff_200760_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3388 diff_202800_59760# diff_100440_59160# diff_202800_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3389 diff_204840_59760# diff_100440_59160# diff_204840_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3390 diff_206880_59760# diff_100440_59160# diff_206880_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3391 diff_208920_59760# diff_100440_59160# diff_208920_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3392 diff_210960_59760# diff_100440_59160# diff_210960_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3393 diff_213000_59760# diff_100440_59160# diff_213000_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3394 diff_215040_59760# diff_100440_59160# diff_215040_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3395 diff_217080_59760# diff_100440_59160# diff_217080_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3396 diff_219120_59760# diff_100440_59160# diff_219120_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3397 diff_221160_59760# diff_100440_59160# diff_221160_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3398 diff_223200_59760# diff_100440_59160# diff_223200_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3399 diff_225240_59760# diff_100440_59160# diff_225240_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3400 diff_227280_59760# diff_100440_59160# diff_227280_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3401 diff_229320_59760# diff_100440_59160# diff_229320_57480# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3402 diff_100440_65760# diff_243120_97920# diff_236760_60720# GND efet w=7920 l=600
+ ad=0 pd=0 as=0 ps=0 
M3403 diff_250800_43080# diff_245160_97920# diff_236760_69600# GND efet w=15480 l=720
+ ad=7.18272e+07 pd=112560 as=0 ps=0 
M3404 diff_236760_60720# diff_246960_91200# diff_250800_43080# GND efet w=15480 l=720
+ ad=0 pd=0 as=0 ps=0 
M3405 diff_236760_51960# diff_236160_42720# diff_100440_52440# GND efet w=8760 l=660
+ ad=3.6432e+07 pd=72960 as=7.9488e+06 ps=22320 
M3406 diff_100800_57480# diff_100440_56880# diff_100800_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3407 diff_102840_57480# diff_100440_56880# diff_102840_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3408 diff_104880_57480# diff_100440_56880# diff_104880_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3409 diff_106920_57480# diff_100440_56880# diff_106920_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3410 diff_108960_57480# diff_100440_56880# diff_108960_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3411 diff_111000_57480# diff_100440_56880# diff_111000_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3412 diff_113040_57480# diff_100440_56880# diff_113040_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3413 diff_115080_57480# diff_100440_56880# diff_115080_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3414 diff_117120_57480# diff_100440_56880# diff_117120_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3415 diff_119160_57480# diff_100440_56880# diff_119160_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3416 diff_121200_57480# diff_100440_56880# diff_121200_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3417 diff_123240_57480# diff_100440_56880# diff_123240_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3418 diff_125280_57480# diff_100440_56880# diff_125280_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3419 diff_127320_57480# diff_100440_56880# diff_127320_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3420 diff_129360_57480# diff_100440_56880# diff_129360_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3421 diff_131400_57480# diff_100440_56880# diff_131400_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3422 diff_133440_57480# diff_100440_56880# diff_133440_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3423 diff_135480_57480# diff_100440_56880# diff_135480_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3424 diff_137520_57480# diff_100440_56880# diff_137520_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3425 diff_139560_57480# diff_100440_56880# diff_139560_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3426 diff_141600_57480# diff_100440_56880# diff_141600_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3427 diff_143640_57480# diff_100440_56880# diff_143640_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3428 diff_145680_57480# diff_100440_56880# diff_145680_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3429 diff_147720_57480# diff_100440_56880# diff_147720_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3430 diff_149760_57480# diff_100440_56880# diff_149760_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3431 diff_151800_57480# diff_100440_56880# diff_151800_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3432 diff_153840_57480# diff_100440_56880# diff_153840_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3433 diff_155880_57480# diff_100440_56880# diff_155880_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3434 diff_157920_57480# diff_100440_56880# diff_157920_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3435 diff_159960_57480# diff_100440_56880# diff_159960_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3436 diff_162000_57480# diff_100440_56880# diff_162000_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3437 diff_164040_57480# diff_100440_56880# diff_164040_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3438 diff_166080_57480# diff_100440_56880# diff_166080_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3439 diff_168120_57480# diff_100440_56880# diff_168120_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3440 diff_170160_57480# diff_100440_56880# diff_170160_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3441 diff_172200_57480# diff_100440_56880# diff_172200_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3442 diff_174240_57480# diff_100440_56880# diff_174240_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3443 diff_176280_57480# diff_100440_56880# diff_176280_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3444 diff_178320_57480# diff_100440_56880# diff_178320_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3445 diff_180360_57480# diff_100440_56880# diff_180360_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3446 diff_182400_57480# diff_100440_56880# diff_182400_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3447 diff_184440_57480# diff_100440_56880# diff_184440_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3448 diff_186480_57480# diff_100440_56880# diff_186480_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3449 diff_188520_57480# diff_100440_56880# diff_188520_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3450 diff_190560_57480# diff_100440_56880# diff_190560_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3451 diff_192600_57480# diff_100440_56880# diff_192600_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3452 diff_194640_57480# diff_100440_56880# diff_194640_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3453 diff_196680_57480# diff_100440_56880# diff_196680_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3454 diff_198720_57480# diff_100440_56880# diff_198720_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3455 diff_200760_57480# diff_100440_56880# diff_200760_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3456 diff_202800_57480# diff_100440_56880# diff_202800_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3457 diff_204840_57480# diff_100440_56880# diff_204840_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3458 diff_206880_57480# diff_100440_56880# diff_206880_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3459 diff_208920_57480# diff_100440_56880# diff_208920_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3460 diff_210960_57480# diff_100440_56880# diff_210960_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3461 diff_213000_57480# diff_100440_56880# diff_213000_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3462 diff_215040_57480# diff_100440_56880# diff_215040_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3463 diff_217080_57480# diff_100440_56880# diff_217080_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3464 diff_219120_57480# diff_100440_56880# diff_219120_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3465 diff_221160_57480# diff_100440_56880# diff_221160_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3466 diff_223200_57480# diff_100440_56880# diff_223200_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3467 diff_225240_57480# diff_100440_56880# diff_225240_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3468 diff_227280_57480# diff_100440_56880# diff_227280_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3469 diff_229320_57480# diff_100440_56880# diff_229320_55320# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3470 diff_100440_59160# Vdd Vdd GND efet w=600 l=1320
+ ad=9.4032e+06 pd=26160 as=0 ps=0 
M3471 diff_77640_48840# Vdd Vdd GND efet w=780 l=8700
+ ad=3.6288e+06 pd=10800 as=0 ps=0 
M3472 diff_100800_55320# diff_100440_54720# diff_100800_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3473 diff_102840_55320# diff_100440_54720# diff_102840_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3474 diff_104880_55320# diff_100440_54720# diff_104880_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3475 diff_106920_55320# diff_100440_54720# diff_106920_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3476 diff_108960_55320# diff_100440_54720# diff_108960_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3477 diff_111000_55320# diff_100440_54720# diff_111000_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3478 diff_113040_55320# diff_100440_54720# diff_113040_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3479 diff_115080_55320# diff_100440_54720# diff_115080_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3480 diff_117120_55320# diff_100440_54720# diff_117120_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3481 diff_119160_55320# diff_100440_54720# diff_119160_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3482 diff_121200_55320# diff_100440_54720# diff_121200_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3483 diff_123240_55320# diff_100440_54720# diff_123240_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3484 diff_125280_55320# diff_100440_54720# diff_125280_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3485 diff_127320_55320# diff_100440_54720# diff_127320_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3486 diff_129360_55320# diff_100440_54720# diff_129360_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3487 diff_131400_55320# diff_100440_54720# diff_131400_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3488 diff_133440_55320# diff_100440_54720# diff_133440_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3489 diff_135480_55320# diff_100440_54720# diff_135480_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3490 diff_137520_55320# diff_100440_54720# diff_137520_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3491 diff_139560_55320# diff_100440_54720# diff_139560_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3492 diff_141600_55320# diff_100440_54720# diff_141600_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3493 diff_143640_55320# diff_100440_54720# diff_143640_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3494 diff_145680_55320# diff_100440_54720# diff_145680_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3495 diff_147720_55320# diff_100440_54720# diff_147720_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3496 diff_149760_55320# diff_100440_54720# diff_149760_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3497 diff_151800_55320# diff_100440_54720# diff_151800_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3498 diff_153840_55320# diff_100440_54720# diff_153840_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3499 diff_155880_55320# diff_100440_54720# diff_155880_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3500 diff_157920_55320# diff_100440_54720# diff_157920_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3501 diff_159960_55320# diff_100440_54720# diff_159960_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3502 diff_162000_55320# diff_100440_54720# diff_162000_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3503 diff_164040_55320# diff_100440_54720# diff_164040_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3504 diff_166080_55320# diff_100440_54720# diff_166080_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3505 diff_168120_55320# diff_100440_54720# diff_168120_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3506 diff_170160_55320# diff_100440_54720# diff_170160_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3507 diff_172200_55320# diff_100440_54720# diff_172200_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3508 diff_174240_55320# diff_100440_54720# diff_174240_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3509 diff_176280_55320# diff_100440_54720# diff_176280_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3510 diff_178320_55320# diff_100440_54720# diff_178320_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3511 diff_180360_55320# diff_100440_54720# diff_180360_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3512 diff_182400_55320# diff_100440_54720# diff_182400_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3513 diff_184440_55320# diff_100440_54720# diff_184440_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3514 diff_186480_55320# diff_100440_54720# diff_186480_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3515 diff_188520_55320# diff_100440_54720# diff_188520_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3516 diff_190560_55320# diff_100440_54720# diff_190560_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3517 diff_192600_55320# diff_100440_54720# diff_192600_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3518 diff_194640_55320# diff_100440_54720# diff_194640_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3519 diff_196680_55320# diff_100440_54720# diff_196680_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3520 diff_198720_55320# diff_100440_54720# diff_198720_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3521 diff_200760_55320# diff_100440_54720# diff_200760_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3522 diff_202800_55320# diff_100440_54720# diff_202800_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3523 diff_204840_55320# diff_100440_54720# diff_204840_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3524 diff_206880_55320# diff_100440_54720# diff_206880_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3525 diff_208920_55320# diff_100440_54720# diff_208920_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3526 diff_210960_55320# diff_100440_54720# diff_210960_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3527 diff_213000_55320# diff_100440_54720# diff_213000_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3528 diff_215040_55320# diff_100440_54720# diff_215040_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3529 diff_217080_55320# diff_100440_54720# diff_217080_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3530 diff_219120_55320# diff_100440_54720# diff_219120_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3531 diff_221160_55320# diff_100440_54720# diff_221160_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3532 diff_223200_55320# diff_100440_54720# diff_223200_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3533 diff_225240_55320# diff_100440_54720# diff_225240_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3534 diff_227280_55320# diff_100440_54720# diff_227280_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3535 diff_229320_55320# diff_100440_54720# diff_229320_53040# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3536 diff_40920_47640# diff_40440_47040# GND GND efet w=3240 l=720
+ ad=0 pd=0 as=0 ps=0 
M3537 diff_49080_50040# diff_49680_49200# diff_50040_48000# GND efet w=1920 l=720
+ ad=0 pd=0 as=3.096e+06 ps=8880 
M3538 diff_78000_44640# diff_77640_48840# diff_69120_48720# GND efet w=1320 l=720
+ ad=8.7552e+06 pd=19680 as=0 ps=0 
M3539 diff_49680_49200# diff_81000_51000# diff_78000_44640# GND efet w=1320 l=720
+ ad=1.04688e+07 pd=24000 as=0 ps=0 
M3540 diff_50040_48000# cm GND GND efet w=3360 l=720
+ ad=0 pd=0 as=0 ps=0 
M3541 diff_69480_49320# diff_69120_48720# diff_69480_47880# GND efet w=3000 l=720
+ ad=0 pd=0 as=2.3184e+06 ps=8400 
M3542 diff_69120_48720# diff_69120_48720# diff_69120_48720# GND efet w=120 l=120
+ ad=0 pd=0 as=0 ps=0 
M3543 diff_69120_48720# diff_69120_48720# diff_69120_48720# GND efet w=180 l=300
+ ad=0 pd=0 as=0 ps=0 
M3544 diff_69480_47880# diff_69120_47280# GND GND efet w=3480 l=660
+ ad=0 pd=0 as=0 ps=0 
M3545 diff_56400_47520# diff_55080_45480# GND GND efet w=4560 l=720
+ ad=0 pd=0 as=0 ps=0 
M3546 diff_62400_47520# diff_62160_46920# GND GND efet w=4560 l=720
+ ad=0 pd=0 as=0 ps=0 
M3547 diff_33840_37560# diff_32160_39840# GND GND efet w=2040 l=720
+ ad=8.856e+06 pd=20400 as=0 ps=0 
M3548 diff_38280_37560# diff_36720_39840# GND GND efet w=1920 l=720
+ ad=7.488e+06 pd=19200 as=0 ps=0 
M3549 diff_42960_37560# diff_41400_39840# GND GND efet w=2040 l=720
+ ad=6.8544e+06 pd=18720 as=0 ps=0 
M3550 diff_32160_39840# clk1 diff_28920_45720# GND efet w=1080 l=720
+ ad=1.3824e+06 pd=5520 as=0 ps=0 
M3551 diff_32160_39840# diff_32160_39840# diff_32160_39840# GND efet w=120 l=540
+ ad=0 pd=0 as=0 ps=0 
M3552 diff_32160_39840# diff_32160_39840# diff_32160_39840# GND efet w=180 l=240
+ ad=0 pd=0 as=0 ps=0 
M3553 diff_36720_39840# clk2 diff_33840_37560# GND efet w=1200 l=720
+ ad=1.4832e+06 pd=5280 as=0 ps=0 
M3554 diff_36720_39840# diff_36720_39840# diff_36720_39840# GND efet w=180 l=300
+ ad=0 pd=0 as=0 ps=0 
M3555 diff_36720_39840# diff_36720_39840# diff_36720_39840# GND efet w=60 l=120
+ ad=0 pd=0 as=0 ps=0 
M3556 diff_41400_39840# clk1 diff_38280_37560# GND efet w=1200 l=720
+ ad=1.4256e+06 pd=5520 as=0 ps=0 
M3557 diff_41400_39840# diff_41400_39840# diff_41400_39840# GND efet w=240 l=420
+ ad=0 pd=0 as=0 ps=0 
M3558 GND diff_75600_45480# diff_69120_48720# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M3559 diff_47400_37560# diff_45960_39840# GND GND efet w=1920 l=720
+ ad=7.4016e+06 pd=19200 as=0 ps=0 
M3560 diff_47880_47040# diff_50640_39840# GND GND efet w=2040 l=720
+ ad=8.5824e+06 pd=21120 as=0 ps=0 
M3561 diff_55080_45480# diff_55080_39840# GND GND efet w=1920 l=720
+ ad=8.7408e+06 pd=21120 as=0 ps=0 
M3562 diff_61320_37560# diff_59760_39840# GND GND efet w=2040 l=720
+ ad=6.8544e+06 pd=18720 as=0 ps=0 
M3563 diff_62160_46920# diff_64320_39840# GND GND efet w=1920 l=720
+ ad=8.5392e+06 pd=21120 as=0 ps=0 
M3564 diff_75600_45480# diff_78000_44640# GND GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M3565 diff_77640_48840# diff_77640_48840# diff_77640_48840# GND efet w=60 l=180
+ ad=0 pd=0 as=0 ps=0 
M3566 diff_81000_51000# diff_77640_48840# GND GND efet w=1200 l=720
+ ad=0 pd=0 as=0 ps=0 
M3567 diff_77640_48840# diff_77640_48840# diff_77640_48840# GND efet w=120 l=120
+ ad=0 pd=0 as=0 ps=0 
M3568 diff_78000_44640# diff_78000_44640# diff_78000_44640# GND efet w=180 l=540
+ ad=0 pd=0 as=0 ps=0 
M3569 diff_78000_44640# diff_78000_44640# diff_78000_44640# GND efet w=180 l=420
+ ad=0 pd=0 as=0 ps=0 
M3570 diff_90480_46440# clk2 diff_77640_48840# GND efet w=2280 l=720
+ ad=2.8944e+06 pd=7920 as=0 ps=0 
M3571 diff_92280_45840# diff_74640_62520# diff_90480_46440# GND efet w=2880 l=720
+ ad=9.3024e+06 pd=19920 as=0 ps=0 
M3572 Vdd Vdd diff_100440_52440# GND efet w=600 l=1320
+ ad=0 pd=0 as=0 ps=0 
M3573 diff_100800_53040# diff_100440_52440# diff_100800_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3574 diff_102840_53040# diff_100440_52440# diff_102840_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3575 diff_104880_53040# diff_100440_52440# diff_104880_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3576 diff_106920_53040# diff_100440_52440# diff_106920_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3577 diff_108960_53040# diff_100440_52440# diff_108960_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3578 diff_111000_53040# diff_100440_52440# diff_111000_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3579 diff_113040_53040# diff_100440_52440# diff_113040_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3580 diff_115080_53040# diff_100440_52440# diff_115080_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3581 diff_117120_53040# diff_100440_52440# diff_117120_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3582 diff_119160_53040# diff_100440_52440# diff_119160_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3583 diff_121200_53040# diff_100440_52440# diff_121200_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3584 diff_123240_53040# diff_100440_52440# diff_123240_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3585 diff_125280_53040# diff_100440_52440# diff_125280_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3586 diff_127320_53040# diff_100440_52440# diff_127320_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3587 diff_129360_53040# diff_100440_52440# diff_129360_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3588 diff_131400_53040# diff_100440_52440# diff_131400_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3589 diff_133440_53040# diff_100440_52440# diff_133440_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3590 diff_135480_53040# diff_100440_52440# diff_135480_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3591 diff_137520_53040# diff_100440_52440# diff_137520_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3592 diff_139560_53040# diff_100440_52440# diff_139560_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3593 diff_141600_53040# diff_100440_52440# diff_141600_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3594 diff_143640_53040# diff_100440_52440# diff_143640_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3595 diff_145680_53040# diff_100440_52440# diff_145680_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3596 diff_147720_53040# diff_100440_52440# diff_147720_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3597 diff_149760_53040# diff_100440_52440# diff_149760_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3598 diff_151800_53040# diff_100440_52440# diff_151800_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3599 diff_153840_53040# diff_100440_52440# diff_153840_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3600 diff_155880_53040# diff_100440_52440# diff_155880_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3601 diff_157920_53040# diff_100440_52440# diff_157920_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3602 diff_159960_53040# diff_100440_52440# diff_159960_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3603 diff_162000_53040# diff_100440_52440# diff_162000_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3604 diff_164040_53040# diff_100440_52440# diff_164040_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3605 diff_166080_53040# diff_100440_52440# diff_166080_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3606 diff_168120_53040# diff_100440_52440# diff_168120_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3607 diff_170160_53040# diff_100440_52440# diff_170160_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3608 diff_172200_53040# diff_100440_52440# diff_172200_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3609 diff_174240_53040# diff_100440_52440# diff_174240_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3610 diff_176280_53040# diff_100440_52440# diff_176280_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3611 diff_178320_53040# diff_100440_52440# diff_178320_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3612 diff_180360_53040# diff_100440_52440# diff_180360_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3613 diff_182400_53040# diff_100440_52440# diff_182400_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3614 diff_184440_53040# diff_100440_52440# diff_184440_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3615 diff_186480_53040# diff_100440_52440# diff_186480_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3616 diff_188520_53040# diff_100440_52440# diff_188520_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3617 diff_190560_53040# diff_100440_52440# diff_190560_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3618 diff_192600_53040# diff_100440_52440# diff_192600_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3619 diff_194640_53040# diff_100440_52440# diff_194640_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3620 diff_196680_53040# diff_100440_52440# diff_196680_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3621 diff_198720_53040# diff_100440_52440# diff_198720_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3622 diff_200760_53040# diff_100440_52440# diff_200760_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3623 diff_202800_53040# diff_100440_52440# diff_202800_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3624 diff_204840_53040# diff_100440_52440# diff_204840_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3625 diff_206880_53040# diff_100440_52440# diff_206880_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3626 diff_208920_53040# diff_100440_52440# diff_208920_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3627 diff_210960_53040# diff_100440_52440# diff_210960_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3628 diff_213000_53040# diff_100440_52440# diff_213000_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3629 diff_215040_53040# diff_100440_52440# diff_215040_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3630 diff_217080_53040# diff_100440_52440# diff_217080_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3631 diff_219120_53040# diff_100440_52440# diff_219120_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3632 diff_221160_53040# diff_100440_52440# diff_221160_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3633 diff_223200_53040# diff_100440_52440# diff_223200_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3634 diff_225240_53040# diff_100440_52440# diff_225240_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3635 diff_227280_53040# diff_100440_52440# diff_227280_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3636 diff_229320_53040# diff_100440_52440# diff_229320_50880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3637 diff_100440_59160# diff_238440_42720# diff_236760_51960# GND efet w=7440 l=600
+ ad=0 pd=0 as=0 ps=0 
M3638 diff_100440_56880# Vdd Vdd GND efet w=720 l=1320
+ ad=1.0368e+07 pd=24960 as=0 ps=0 
M3639 Vdd Vdd diff_100440_54720# GND efet w=720 l=1440
+ ad=0 pd=0 as=1.02816e+07 ps=22080 
M3640 diff_236760_51960# diff_241320_99600# diff_100440_54720# GND efet w=8460 l=660
+ ad=0 pd=0 as=0 ps=0 
M3641 diff_100800_50880# diff_100440_50280# diff_100800_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3642 diff_102840_50880# diff_100440_50280# diff_102840_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3643 diff_104880_50880# diff_100440_50280# diff_104880_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3644 diff_106920_50880# diff_100440_50280# diff_106920_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3645 diff_108960_50880# diff_100440_50280# diff_108960_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3646 diff_111000_50880# diff_100440_50280# diff_111000_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3647 diff_113040_50880# diff_100440_50280# diff_113040_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3648 diff_115080_50880# diff_100440_50280# diff_115080_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3649 diff_117120_50880# diff_100440_50280# diff_117120_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3650 diff_119160_50880# diff_100440_50280# diff_119160_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3651 diff_121200_50880# diff_100440_50280# diff_121200_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3652 diff_123240_50880# diff_100440_50280# diff_123240_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3653 diff_125280_50880# diff_100440_50280# diff_125280_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3654 diff_127320_50880# diff_100440_50280# diff_127320_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3655 diff_129360_50880# diff_100440_50280# diff_129360_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3656 diff_131400_50880# diff_100440_50280# diff_131400_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3657 diff_133440_50880# diff_100440_50280# diff_133440_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3658 diff_135480_50880# diff_100440_50280# diff_135480_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3659 diff_137520_50880# diff_100440_50280# diff_137520_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3660 diff_139560_50880# diff_100440_50280# diff_139560_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3661 diff_141600_50880# diff_100440_50280# diff_141600_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3662 diff_143640_50880# diff_100440_50280# diff_143640_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3663 diff_145680_50880# diff_100440_50280# diff_145680_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3664 diff_147720_50880# diff_100440_50280# diff_147720_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3665 diff_149760_50880# diff_100440_50280# diff_149760_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3666 diff_151800_50880# diff_100440_50280# diff_151800_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3667 diff_153840_50880# diff_100440_50280# diff_153840_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3668 diff_155880_50880# diff_100440_50280# diff_155880_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3669 diff_157920_50880# diff_100440_50280# diff_157920_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3670 diff_159960_50880# diff_100440_50280# diff_159960_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3671 diff_162000_50880# diff_100440_50280# diff_162000_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3672 diff_164040_50880# diff_100440_50280# diff_164040_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3673 diff_166080_50880# diff_100440_50280# diff_166080_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3674 diff_168120_50880# diff_100440_50280# diff_168120_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3675 diff_170160_50880# diff_100440_50280# diff_170160_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3676 diff_172200_50880# diff_100440_50280# diff_172200_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3677 diff_174240_50880# diff_100440_50280# diff_174240_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3678 diff_176280_50880# diff_100440_50280# diff_176280_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3679 diff_178320_50880# diff_100440_50280# diff_178320_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3680 diff_180360_50880# diff_100440_50280# diff_180360_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3681 diff_182400_50880# diff_100440_50280# diff_182400_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3682 diff_184440_50880# diff_100440_50280# diff_184440_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3683 diff_186480_50880# diff_100440_50280# diff_186480_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3684 diff_188520_50880# diff_100440_50280# diff_188520_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3685 diff_190560_50880# diff_100440_50280# diff_190560_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3686 diff_192600_50880# diff_100440_50280# diff_192600_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3687 diff_194640_50880# diff_100440_50280# diff_194640_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3688 diff_196680_50880# diff_100440_50280# diff_196680_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3689 diff_198720_50880# diff_100440_50280# diff_198720_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3690 diff_200760_50880# diff_100440_50280# diff_200760_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3691 diff_202800_50880# diff_100440_50280# diff_202800_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3692 diff_204840_50880# diff_100440_50280# diff_204840_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3693 diff_206880_50880# diff_100440_50280# diff_206880_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3694 diff_208920_50880# diff_100440_50280# diff_208920_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3695 diff_210960_50880# diff_100440_50280# diff_210960_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3696 diff_213000_50880# diff_100440_50280# diff_213000_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3697 diff_215040_50880# diff_100440_50280# diff_215040_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3698 diff_217080_50880# diff_100440_50280# diff_217080_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3699 diff_219120_50880# diff_100440_50280# diff_219120_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3700 diff_221160_50880# diff_100440_50280# diff_221160_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3701 diff_223200_50880# diff_100440_50280# diff_223200_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3702 diff_225240_50880# diff_100440_50280# diff_225240_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3703 diff_227280_50880# diff_100440_50280# diff_227280_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3704 diff_229320_50880# diff_100440_50280# diff_229320_48600# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3705 diff_100440_56880# diff_243120_97920# diff_236760_51960# GND efet w=7920 l=600
+ ad=0 pd=0 as=0 ps=0 
M3706 Vdd Vdd Vdd GND efet w=540 l=780
+ ad=0 pd=0 as=0 ps=0 
M3707 Vdd Vdd diff_248880_85320# GND efet w=720 l=1440
+ ad=0 pd=0 as=2.42928e+07 ps=42240 
M3708 diff_277440_100200# Vdd Vdd GND efet w=720 l=3240
+ ad=0 pd=0 as=0 ps=0 
M3709 diff_284880_99240# diff_277920_48600# diff_284880_97680# GND efet w=4680 l=600
+ ad=0 pd=0 as=4.4928e+06 ps=11280 
M3710 Vdd Vdd Vdd GND efet w=240 l=480
+ ad=0 pd=0 as=0 ps=0 
M3711 Vdd Vdd Vdd GND efet w=180 l=420
+ ad=0 pd=0 as=0 ps=0 
M3712 Vdd Vdd diff_277440_88920# GND efet w=720 l=3240
+ ad=0 pd=0 as=9.7776e+06 ps=16080 
M3713 diff_284880_97680# diff_273240_54960# GND GND efet w=4680 l=600
+ ad=0 pd=0 as=0 ps=0 
M3714 diff_273840_92640# diff_271080_135600# diff_252960_89400# GND efet w=2040 l=600
+ ad=0 pd=0 as=3.1536e+06 ps=7200 
M3715 diff_277440_88920# clk2 diff_273840_92640# GND efet w=2040 l=600
+ ad=0 pd=0 as=0 ps=0 
M3716 diff_281880_88920# diff_273840_55200# diff_277440_88920# GND efet w=3720 l=600
+ ad=9.6048e+06 pd=19920 as=0 ps=0 
M3717 diff_273840_81360# diff_271080_135600# diff_259800_65640# GND efet w=2040 l=600
+ ad=5.8464e+06 pd=13920 as=2.9088e+06 ps=6960 
M3718 diff_277440_85200# clk2 diff_273840_81360# GND efet w=2040 l=600
+ ad=1.15632e+07 pd=21120 as=0 ps=0 
M3719 Vdd Vdd diff_104880_84600# GND efet w=720 l=1320
+ ad=0 pd=0 as=1.81152e+07 ps=32400 
M3720 Vdd Vdd diff_99480_122520# GND efet w=720 l=1320
+ ad=0 pd=0 as=2.10816e+07 ps=32880 
M3721 Vdd Vdd diff_250560_91920# GND efet w=840 l=1320
+ ad=0 pd=0 as=1.99008e+07 ps=32640 
M3722 diff_273840_81360# diff_272280_84480# diff_261720_78960# GND efet w=2040 l=600
+ ad=0 pd=0 as=2.9088e+06 ps=6960 
M3723 GND diff_259800_65640# diff_248880_85320# GND efet w=12360 l=600
+ ad=0 pd=0 as=0 ps=0 
M3724 diff_104880_84600# diff_261720_78960# GND GND efet w=12360 l=600
+ ad=0 pd=0 as=0 ps=0 
M3725 GND diff_266520_78960# diff_99480_122520# GND efet w=12360 l=600
+ ad=0 pd=0 as=0 ps=0 
M3726 diff_250560_91920# diff_268680_78960# GND GND efet w=12360 l=600
+ ad=0 pd=0 as=0 ps=0 
M3727 diff_273840_77640# diff_272280_84480# diff_266520_78960# GND efet w=2040 l=600
+ ad=6.0336e+06 pd=14160 as=2.9088e+06 ps=6960 
M3728 diff_277440_85200# Vdd Vdd GND efet w=720 l=3360
+ ad=0 pd=0 as=0 ps=0 
M3729 Vdd Vdd Vdd GND efet w=300 l=660
+ ad=0 pd=0 as=0 ps=0 
M3730 Vdd Vdd Vdd GND efet w=120 l=480
+ ad=0 pd=0 as=0 ps=0 
M3731 Vdd Vdd diff_277440_73800# GND efet w=720 l=3240
+ ad=0 pd=0 as=1.0152e+07 ps=16080 
M3732 diff_286560_90000# diff_273240_54960# diff_277440_100200# GND efet w=3840 l=600
+ ad=3.6864e+06 pd=9600 as=0 ps=0 
M3733 GND diff_275160_45240# diff_286560_90000# GND efet w=3840 l=600
+ ad=0 pd=0 as=0 ps=0 
M3734 d0 GND d0 GND efet w=17940 l=11220
+ ad=0 pd=0 as=0 ps=0 
M3735 GND diff_275160_45240# diff_281880_88920# GND efet w=3600 l=600
+ ad=0 pd=0 as=0 ps=0 
M3736 diff_284160_79920# diff_277920_48600# diff_277440_85200# GND efet w=3600 l=600
+ ad=3.456e+06 pd=9120 as=0 ps=0 
M3737 GND diff_273240_54960# diff_284160_79920# GND efet w=3600 l=600
+ ad=0 pd=0 as=0 ps=0 
M3738 diff_273840_77640# diff_271080_135600# diff_268680_78960# GND efet w=2160 l=600
+ ad=0 pd=0 as=3.312e+06 ps=7440 
M3739 diff_277440_73800# clk2 diff_273840_77640# GND efet w=2160 l=600
+ ad=0 pd=0 as=0 ps=0 
M3740 diff_281880_73800# diff_273840_55200# diff_277440_73800# GND efet w=3840 l=600
+ ad=3.6864e+06 pd=9600 as=0 ps=0 
M3741 GND diff_277920_48600# diff_281880_73800# GND efet w=3840 l=600
+ ad=0 pd=0 as=0 ps=0 
M3742 Vdd Vdd Vdd GND efet w=240 l=420
+ ad=0 pd=0 as=0 ps=0 
M3743 Vdd Vdd Vdd GND efet w=240 l=480
+ ad=0 pd=0 as=0 ps=0 
M3744 diff_273240_54960# Vdd Vdd GND efet w=1080 l=1680
+ ad=1.73808e+07 pd=33840 as=0 ps=0 
M3745 GND diff_243360_174240# diff_250800_43080# GND efet w=30120 l=600
+ ad=0 pd=0 as=0 ps=0 
M3746 diff_236760_43080# diff_236160_42720# diff_100440_43560# GND efet w=8940 l=720
+ ad=3.79584e+07 pd=69120 as=8.6112e+06 ps=22800 
M3747 diff_100800_48600# diff_100440_48000# diff_100800_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3748 diff_102840_48600# diff_100440_48000# diff_102840_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3749 diff_104880_48600# diff_100440_48000# diff_104880_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3750 diff_106920_48600# diff_100440_48000# diff_106920_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3751 diff_108960_48600# diff_100440_48000# diff_108960_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3752 diff_111000_48600# diff_100440_48000# diff_111000_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3753 diff_113040_48600# diff_100440_48000# diff_113040_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3754 diff_115080_48600# diff_100440_48000# diff_115080_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3755 diff_117120_48600# diff_100440_48000# diff_117120_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3756 diff_119160_48600# diff_100440_48000# diff_119160_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3757 diff_121200_48600# diff_100440_48000# diff_121200_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3758 diff_123240_48600# diff_100440_48000# diff_123240_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3759 diff_125280_48600# diff_100440_48000# diff_125280_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3760 diff_127320_48600# diff_100440_48000# diff_127320_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3761 diff_129360_48600# diff_100440_48000# diff_129360_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3762 diff_131400_48600# diff_100440_48000# diff_131400_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3763 diff_133440_48600# diff_100440_48000# diff_133440_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3764 diff_135480_48600# diff_100440_48000# diff_135480_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3765 diff_137520_48600# diff_100440_48000# diff_137520_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3766 diff_139560_48600# diff_100440_48000# diff_139560_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3767 diff_141600_48600# diff_100440_48000# diff_141600_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3768 diff_143640_48600# diff_100440_48000# diff_143640_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3769 diff_145680_48600# diff_100440_48000# diff_145680_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3770 diff_147720_48600# diff_100440_48000# diff_147720_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3771 diff_149760_48600# diff_100440_48000# diff_149760_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3772 diff_151800_48600# diff_100440_48000# diff_151800_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3773 diff_153840_48600# diff_100440_48000# diff_153840_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3774 diff_155880_48600# diff_100440_48000# diff_155880_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3775 diff_157920_48600# diff_100440_48000# diff_157920_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3776 diff_159960_48600# diff_100440_48000# diff_159960_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3777 diff_162000_48600# diff_100440_48000# diff_162000_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3778 diff_164040_48600# diff_100440_48000# diff_164040_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3779 diff_166080_48600# diff_100440_48000# diff_166080_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3780 diff_168120_48600# diff_100440_48000# diff_168120_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3781 diff_170160_48600# diff_100440_48000# diff_170160_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3782 diff_172200_48600# diff_100440_48000# diff_172200_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3783 diff_174240_48600# diff_100440_48000# diff_174240_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3784 diff_176280_48600# diff_100440_48000# diff_176280_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3785 diff_178320_48600# diff_100440_48000# diff_178320_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3786 diff_180360_48600# diff_100440_48000# diff_180360_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3787 diff_182400_48600# diff_100440_48000# diff_182400_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3788 diff_184440_48600# diff_100440_48000# diff_184440_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3789 diff_186480_48600# diff_100440_48000# diff_186480_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3790 diff_188520_48600# diff_100440_48000# diff_188520_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3791 diff_190560_48600# diff_100440_48000# diff_190560_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3792 diff_192600_48600# diff_100440_48000# diff_192600_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3793 diff_194640_48600# diff_100440_48000# diff_194640_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3794 diff_196680_48600# diff_100440_48000# diff_196680_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3795 diff_198720_48600# diff_100440_48000# diff_198720_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3796 diff_200760_48600# diff_100440_48000# diff_200760_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3797 diff_202800_48600# diff_100440_48000# diff_202800_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3798 diff_204840_48600# diff_100440_48000# diff_204840_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3799 diff_206880_48600# diff_100440_48000# diff_206880_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3800 diff_208920_48600# diff_100440_48000# diff_208920_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3801 diff_210960_48600# diff_100440_48000# diff_210960_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3802 diff_213000_48600# diff_100440_48000# diff_213000_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3803 diff_215040_48600# diff_100440_48000# diff_215040_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3804 diff_217080_48600# diff_100440_48000# diff_217080_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3805 diff_219120_48600# diff_100440_48000# diff_219120_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3806 diff_221160_48600# diff_100440_48000# diff_221160_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3807 diff_223200_48600# diff_100440_48000# diff_223200_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3808 diff_225240_48600# diff_100440_48000# diff_225240_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3809 diff_227280_48600# diff_100440_48000# diff_227280_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3810 diff_229320_48600# diff_100440_48000# diff_229320_46440# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.5552e+06 ps=5040 
M3811 diff_100440_50280# Vdd Vdd GND efet w=600 l=1200
+ ad=9.4032e+06 pd=26160 as=0 ps=0 
M3812 GND cm diff_92280_45840# GND efet w=6720 l=720
+ ad=0 pd=0 as=0 ps=0 
M3813 diff_69120_47280# clk1 GND GND efet w=2040 l=720
+ ad=8.3088e+06 pd=20640 as=0 ps=0 
M3814 diff_74880_37560# diff_73320_39840# GND GND efet w=1920 l=720
+ ad=7.488e+06 pd=19200 as=0 ps=0 
M3815 diff_79560_37560# diff_78000_39840# GND GND efet w=2040 l=720
+ ad=6.8544e+06 pd=18720 as=0 ps=0 
M3816 diff_41400_39840# diff_41400_39840# diff_41400_39840# GND efet w=120 l=180
+ ad=0 pd=0 as=0 ps=0 
M3817 diff_45960_39840# clk2 diff_42960_37560# GND efet w=1200 l=720
+ ad=1.3824e+06 pd=4800 as=0 ps=0 
M3818 diff_45960_39840# diff_45960_39840# diff_45960_39840# GND efet w=120 l=180
+ ad=0 pd=0 as=0 ps=0 
M3819 diff_50640_39840# clk1 diff_47400_37560# GND efet w=1200 l=720
+ ad=1.2816e+06 pd=5280 as=0 ps=0 
M3820 diff_50640_39840# diff_50640_39840# diff_50640_39840# GND efet w=240 l=420
+ ad=0 pd=0 as=0 ps=0 
M3821 diff_50640_39840# diff_50640_39840# diff_50640_39840# GND efet w=120 l=180
+ ad=0 pd=0 as=0 ps=0 
M3822 diff_55080_39840# clk2 diff_47880_47040# GND efet w=1200 l=720
+ ad=1.4832e+06 pd=5280 as=0 ps=0 
M3823 diff_55080_39840# diff_55080_39840# diff_55080_39840# GND efet w=180 l=300
+ ad=0 pd=0 as=0 ps=0 
M3824 diff_55080_39840# diff_55080_39840# diff_55080_39840# GND efet w=60 l=120
+ ad=0 pd=0 as=0 ps=0 
M3825 diff_59760_39840# clk1 diff_55080_45480# GND efet w=1200 l=720
+ ad=1.4256e+06 pd=5520 as=0 ps=0 
M3826 diff_59760_39840# diff_59760_39840# diff_59760_39840# GND efet w=240 l=420
+ ad=0 pd=0 as=0 ps=0 
M3827 diff_59760_39840# diff_59760_39840# diff_59760_39840# GND efet w=120 l=180
+ ad=0 pd=0 as=0 ps=0 
M3828 diff_64320_39840# clk2 diff_61320_37560# GND efet w=1200 l=720
+ ad=1.3824e+06 pd=4800 as=0 ps=0 
M3829 diff_64320_39840# diff_64320_39840# diff_64320_39840# GND efet w=120 l=180
+ ad=0 pd=0 as=0 ps=0 
M3830 clk1 clk1 diff_62160_46920# GND efet w=1020 l=900
+ ad=0 pd=0 as=0 ps=0 
M3831 clk1 clk1 clk1 GND efet w=240 l=480
+ ad=0 pd=0 as=0 ps=0 
M3832 clk1 clk1 clk1 GND efet w=180 l=240
+ ad=0 pd=0 as=0 ps=0 
M3833 diff_73320_39840# clk2 diff_69120_47280# GND efet w=1200 l=720
+ ad=1.4832e+06 pd=5280 as=0 ps=0 
M3834 diff_73320_39840# diff_73320_39840# diff_73320_39840# GND efet w=180 l=300
+ ad=0 pd=0 as=0 ps=0 
M3835 diff_73320_39840# diff_73320_39840# diff_73320_39840# GND efet w=60 l=120
+ ad=0 pd=0 as=0 ps=0 
M3836 diff_78000_39840# clk1 diff_74880_37560# GND efet w=1200 l=720
+ ad=1.4256e+06 pd=5520 as=0 ps=0 
M3837 diff_78000_39840# diff_78000_39840# diff_78000_39840# GND efet w=240 l=420
+ ad=0 pd=0 as=0 ps=0 
M3838 diff_84000_37560# diff_82560_39840# GND GND efet w=1920 l=720
+ ad=8.2944e+06 pd=20880 as=0 ps=0 
M3839 diff_74640_62520# diff_87240_39840# GND GND efet w=2040 l=600
+ ad=7.5456e+06 pd=19920 as=0 ps=0 
M3840 diff_100800_46440# diff_100440_45840# diff_100800_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3841 diff_102840_46440# diff_100440_45840# diff_102840_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3842 diff_104880_46440# diff_100440_45840# diff_104880_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3843 diff_106920_46440# diff_100440_45840# diff_106920_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3844 diff_108960_46440# diff_100440_45840# diff_108960_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3845 diff_111000_46440# diff_100440_45840# diff_111000_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3846 diff_113040_46440# diff_100440_45840# diff_113040_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3847 diff_115080_46440# diff_100440_45840# diff_115080_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3848 diff_117120_46440# diff_100440_45840# diff_117120_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3849 diff_119160_46440# diff_100440_45840# diff_119160_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3850 diff_121200_46440# diff_100440_45840# diff_121200_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3851 diff_123240_46440# diff_100440_45840# diff_123240_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3852 diff_125280_46440# diff_100440_45840# diff_125280_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3853 diff_127320_46440# diff_100440_45840# diff_127320_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3854 diff_129360_46440# diff_100440_45840# diff_129360_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3855 diff_131400_46440# diff_100440_45840# diff_131400_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3856 diff_133440_46440# diff_100440_45840# diff_133440_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3857 diff_135480_46440# diff_100440_45840# diff_135480_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3858 diff_137520_46440# diff_100440_45840# diff_137520_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3859 diff_139560_46440# diff_100440_45840# diff_139560_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3860 diff_141600_46440# diff_100440_45840# diff_141600_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3861 diff_143640_46440# diff_100440_45840# diff_143640_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3862 diff_145680_46440# diff_100440_45840# diff_145680_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3863 diff_147720_46440# diff_100440_45840# diff_147720_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3864 diff_149760_46440# diff_100440_45840# diff_149760_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3865 diff_151800_46440# diff_100440_45840# diff_151800_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3866 diff_153840_46440# diff_100440_45840# diff_153840_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3867 diff_155880_46440# diff_100440_45840# diff_155880_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3868 diff_157920_46440# diff_100440_45840# diff_157920_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3869 diff_159960_46440# diff_100440_45840# diff_159960_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3870 diff_162000_46440# diff_100440_45840# diff_162000_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3871 diff_164040_46440# diff_100440_45840# diff_164040_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3872 diff_166080_46440# diff_100440_45840# diff_166080_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3873 diff_168120_46440# diff_100440_45840# diff_168120_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3874 diff_170160_46440# diff_100440_45840# diff_170160_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3875 diff_172200_46440# diff_100440_45840# diff_172200_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3876 diff_174240_46440# diff_100440_45840# diff_174240_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3877 diff_176280_46440# diff_100440_45840# diff_176280_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3878 diff_178320_46440# diff_100440_45840# diff_178320_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3879 diff_180360_46440# diff_100440_45840# diff_180360_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3880 diff_182400_46440# diff_100440_45840# diff_182400_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3881 diff_184440_46440# diff_100440_45840# diff_184440_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3882 diff_186480_46440# diff_100440_45840# diff_186480_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3883 diff_188520_46440# diff_100440_45840# diff_188520_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3884 diff_190560_46440# diff_100440_45840# diff_190560_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3885 diff_192600_46440# diff_100440_45840# diff_192600_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3886 diff_194640_46440# diff_100440_45840# diff_194640_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3887 diff_196680_46440# diff_100440_45840# diff_196680_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3888 diff_198720_46440# diff_100440_45840# diff_198720_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3889 diff_200760_46440# diff_100440_45840# diff_200760_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3890 diff_202800_46440# diff_100440_45840# diff_202800_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3891 diff_204840_46440# diff_100440_45840# diff_204840_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3892 diff_206880_46440# diff_100440_45840# diff_206880_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3893 diff_208920_46440# diff_100440_45840# diff_208920_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3894 diff_210960_46440# diff_100440_45840# diff_210960_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3895 diff_213000_46440# diff_100440_45840# diff_213000_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3896 diff_215040_46440# diff_100440_45840# diff_215040_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3897 diff_217080_46440# diff_100440_45840# diff_217080_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3898 diff_219120_46440# diff_100440_45840# diff_219120_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3899 diff_221160_46440# diff_100440_45840# diff_221160_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3900 diff_223200_46440# diff_100440_45840# diff_223200_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3901 diff_225240_46440# diff_100440_45840# diff_225240_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3902 diff_227280_46440# diff_100440_45840# diff_227280_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3903 diff_229320_46440# diff_100440_45840# diff_229320_44160# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.6848e+06 ps=5280 
M3904 diff_78000_39840# diff_78000_39840# diff_78000_39840# GND efet w=120 l=180
+ ad=0 pd=0 as=0 ps=0 
M3905 diff_82560_39840# clk2 diff_79560_37560# GND efet w=1200 l=720
+ ad=1.3824e+06 pd=4800 as=0 ps=0 
M3906 diff_82560_39840# diff_82560_39840# diff_82560_39840# GND efet w=120 l=180
+ ad=0 pd=0 as=0 ps=0 
M3907 diff_87240_39840# clk1 diff_84000_37560# GND efet w=1200 l=720
+ ad=1.3104e+06 pd=5520 as=0 ps=0 
M3908 diff_87240_39840# diff_87240_39840# diff_87240_39840# GND efet w=240 l=300
+ ad=0 pd=0 as=0 ps=0 
M3909 diff_87240_39840# diff_87240_39840# diff_87240_39840# GND efet w=120 l=180
+ ad=0 pd=0 as=0 ps=0 
M3910 Vdd Vdd diff_28920_45720# GND efet w=780 l=3540
+ ad=0 pd=0 as=0 ps=0 
M3911 diff_33840_37560# Vdd Vdd GND efet w=720 l=3480
+ ad=0 pd=0 as=0 ps=0 
M3912 Vdd Vdd diff_38280_37560# GND efet w=780 l=3660
+ ad=0 pd=0 as=0 ps=0 
M3913 diff_42960_37560# Vdd Vdd GND efet w=720 l=3360
+ ad=0 pd=0 as=0 ps=0 
M3914 Vdd Vdd diff_47400_37560# GND efet w=780 l=3780
+ ad=0 pd=0 as=0 ps=0 
M3915 diff_47880_47040# Vdd Vdd GND efet w=720 l=3360
+ ad=0 pd=0 as=0 ps=0 
M3916 Vdd Vdd diff_55080_45480# GND efet w=780 l=3660
+ ad=0 pd=0 as=0 ps=0 
M3917 diff_61320_37560# Vdd Vdd GND efet w=720 l=3360
+ ad=0 pd=0 as=0 ps=0 
M3918 Vdd Vdd diff_62160_46920# GND efet w=780 l=3780
+ ad=0 pd=0 as=0 ps=0 
M3919 diff_69120_47280# Vdd Vdd GND efet w=720 l=3480
+ ad=0 pd=0 as=0 ps=0 
M3920 Vdd Vdd diff_74880_37560# GND efet w=780 l=3660
+ ad=0 pd=0 as=0 ps=0 
M3921 diff_79560_37560# Vdd Vdd GND efet w=720 l=3360
+ ad=0 pd=0 as=0 ps=0 
M3922 Vdd Vdd diff_84000_37560# GND efet w=780 l=3780
+ ad=0 pd=0 as=0 ps=0 
M3923 diff_74640_62520# Vdd Vdd GND efet w=720 l=3360
+ ad=0 pd=0 as=0 ps=0 
M3924 cl GND GND GND efet w=9840 l=720
+ ad=4.0968e+07 pd=96720 as=0 ps=0 
M3925 Vdd Vdd diff_100440_43560# GND efet w=600 l=1200
+ ad=0 pd=0 as=0 ps=0 
M3926 diff_100800_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=1.94515e+08 ps=277680 
M3927 diff_102840_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3928 diff_104880_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3929 diff_106920_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3930 diff_108960_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3931 diff_111000_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3932 diff_113040_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3933 diff_115080_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3934 diff_117120_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3935 diff_119160_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3936 diff_121200_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3937 diff_123240_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3938 diff_125280_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3939 diff_127320_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3940 diff_129360_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3941 diff_131400_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3942 diff_133440_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3943 diff_135480_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3944 diff_137520_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3945 diff_139560_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3946 diff_141600_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3947 diff_143640_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3948 diff_145680_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3949 diff_147720_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3950 diff_149760_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3951 diff_151800_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3952 diff_153840_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3953 diff_155880_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3954 diff_157920_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3955 diff_159960_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3956 diff_162000_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3957 diff_164040_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3958 diff_166080_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3959 diff_168120_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3960 diff_170160_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3961 diff_172200_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3962 diff_174240_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3963 diff_176280_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3964 diff_178320_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3965 diff_180360_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3966 diff_182400_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3967 diff_184440_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3968 diff_186480_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3969 diff_188520_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3970 diff_190560_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3971 diff_192600_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3972 diff_194640_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3973 diff_196680_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3974 diff_198720_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3975 diff_200760_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3976 diff_202800_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3977 diff_204840_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3978 diff_206880_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3979 diff_208920_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3980 diff_210960_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3981 diff_213000_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3982 diff_215040_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3983 diff_217080_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3984 diff_219120_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3985 diff_221160_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3986 diff_223200_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3987 diff_225240_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3988 diff_227280_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3989 diff_229320_44160# diff_100440_43560# diff_100800_41880# GND efet w=1080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3990 diff_100440_50280# diff_238440_42720# diff_236760_43080# GND efet w=7440 l=600
+ ad=0 pd=0 as=0 ps=0 
M3991 diff_100440_48000# Vdd Vdd GND efet w=720 l=1200
+ ad=1.0368e+07 pd=24960 as=0 ps=0 
M3992 Vdd Vdd diff_100440_45840# GND efet w=720 l=1200
+ ad=0 pd=0 as=9.8496e+06 ps=22080 
M3993 diff_236760_43080# diff_241320_99600# diff_100440_45840# GND efet w=8280 l=720
+ ad=0 pd=0 as=0 ps=0 
M3994 diff_100440_48000# diff_243120_97920# diff_236760_43080# GND efet w=7920 l=600
+ ad=0 pd=0 as=0 ps=0 
M3995 diff_250800_43080# diff_248880_85320# diff_236760_51960# GND efet w=15480 l=720
+ ad=0 pd=0 as=0 ps=0 
M3996 diff_236760_43080# diff_250560_91920# diff_250800_43080# GND efet w=16200 l=720
+ ad=0 pd=0 as=0 ps=0 
M3997 diff_273240_54960# d0 GND GND efet w=17160 l=600
+ ad=0 pd=0 as=0 ps=0 
M3998 diff_285960_61200# diff_273240_54960# diff_95160_43680# GND efet w=8280 l=600
+ ad=8.3088e+06 pd=18720 as=3.30624e+07 ps=70320 
M3999 diff_283200_105600# diff_275160_45240# diff_285960_61200# GND efet w=8400 l=600
+ ad=0 pd=0 as=0 ps=0 
M4000 diff_273840_55200# diff_273240_54960# GND GND efet w=4440 l=600
+ ad=7.2432e+06 pd=15360 as=0 ps=0 
M4001 diff_273840_55200# Vdd Vdd GND efet w=720 l=1680
+ ad=0 pd=0 as=0 ps=0 
M4002 diff_277920_48600# Vdd Vdd GND efet w=960 l=1680
+ ad=5.8032e+06 pd=12480 as=0 ps=0 
M4003 Vdd Vdd diff_275160_45240# GND efet w=720 l=1800
+ ad=0 pd=0 as=2.15712e+07 ps=51840 
M4004 GND diff_275160_45240# diff_277920_48600# GND efet w=4440 l=600
+ ad=0 pd=0 as=0 ps=0 
M4005 diff_275160_45240# d1 GND GND efet w=17160 l=600
+ ad=0 pd=0 as=0 ps=0 
M4006 GND diff_95160_43680# diff_49680_49200# GND efet w=1920 l=720
+ ad=0 pd=0 as=0 ps=0 
M4007 diff_100800_41880# diff_100320_170280# GND GND efet w=61920 l=720
+ ad=0 pd=0 as=0 ps=0 
M4008 diff_100800_41880# diff_165720_170280# Vdd GND efet w=64320 l=720
+ ad=0 pd=0 as=0 ps=0 
M4009 Vdd Vdd Vdd GND efet w=300 l=480
+ ad=0 pd=0 as=0 ps=0 
M4010 Vdd Vdd Vdd GND efet w=240 l=660
+ ad=0 pd=0 as=0 ps=0 
M4011 Vdd Vdd diff_49680_49200# GND efet w=840 l=3360
+ ad=0 pd=0 as=0 ps=0 
M4012 Vdd Vdd Vdd GND efet w=60 l=180
+ ad=0 pd=0 as=0 ps=0 
M4013 Vdd Vdd Vdd GND efet w=240 l=300
+ ad=0 pd=0 as=0 ps=0 
M4014 diff_91920_42120# Vdd Vdd GND efet w=780 l=4140
+ ad=0 pd=0 as=0 ps=0 
M4015 Vdd Vdd diff_95160_43680# GND efet w=900 l=3420
+ ad=0 pd=0 as=0 ps=0 
M4016 cm GND GND GND efet w=9960 l=720
+ ad=3.51504e+07 pd=77040 as=0 ps=0 
C0 metal_182880_18480# gnd! 5.9fF ;**FLOATING
C1 metal_181080_18840# gnd! 7.5fF ;**FLOATING
C2 metal_170880_15600# gnd! 7.1fF ;**FLOATING
C3 metal_170280_15600# gnd! 3.0fF ;**FLOATING
C4 metal_172920_17880# gnd! 21.1fF ;**FLOATING
C5 metal_165720_16680# gnd! 8.3fF ;**FLOATING
C6 metal_179400_15720# gnd! 10.6fF ;**FLOATING
C7 metal_178320_18480# gnd! 5.9fF ;**FLOATING
C8 metal_164880_16320# gnd! 18.4fF ;**FLOATING
C9 metal_41160_16320# gnd! 18.8fF ;**FLOATING
C10 metal_36120_17040# gnd! 39.8fF ;**FLOATING
C11 metal_31200_17280# gnd! 41.6fF ;**FLOATING
C12 metal_26520_18120# gnd! 37.8fF ;**FLOATING
C13 diff_262200_6960# gnd! 3003.1fF ;**FLOATING
C14 diff_285960_61200# gnd! 101.8fF
C15 diff_100800_41880# gnd! 2735.9fF
C16 diff_95160_43680# gnd! 992.1fF
C17 diff_229320_44160# gnd! 26.2fF
C18 diff_227280_44160# gnd! 26.2fF
C19 diff_225240_44160# gnd! 26.2fF
C20 diff_223200_44160# gnd! 26.2fF
C21 diff_221160_44160# gnd! 26.2fF
C22 diff_219120_44160# gnd! 26.2fF
C23 diff_217080_44160# gnd! 26.2fF
C24 diff_215040_44160# gnd! 26.2fF
C25 diff_213000_44160# gnd! 26.2fF
C26 diff_210960_44160# gnd! 26.2fF
C27 diff_208920_44160# gnd! 26.2fF
C28 diff_206880_44160# gnd! 26.2fF
C29 diff_204840_44160# gnd! 26.2fF
C30 diff_202800_44160# gnd! 26.2fF
C31 diff_200760_44160# gnd! 26.2fF
C32 diff_198720_44160# gnd! 26.2fF
C33 diff_196680_44160# gnd! 26.2fF
C34 diff_194640_44160# gnd! 26.2fF
C35 diff_192600_44160# gnd! 26.2fF
C36 diff_190560_44160# gnd! 26.2fF
C37 diff_188520_44160# gnd! 26.2fF
C38 diff_186480_44160# gnd! 26.2fF
C39 diff_184440_44160# gnd! 26.2fF
C40 diff_182400_44160# gnd! 26.2fF
C41 diff_180360_44160# gnd! 26.2fF
C42 diff_178320_44160# gnd! 26.2fF
C43 diff_176280_44160# gnd! 26.2fF
C44 diff_174240_44160# gnd! 26.2fF
C45 diff_172200_44160# gnd! 26.2fF
C46 diff_170160_44160# gnd! 26.2fF
C47 diff_168120_44160# gnd! 26.2fF
C48 diff_166080_44160# gnd! 26.2fF
C49 diff_164040_44160# gnd! 26.2fF
C50 diff_162000_44160# gnd! 26.2fF
C51 diff_159960_44160# gnd! 26.2fF
C52 diff_157920_44160# gnd! 26.2fF
C53 diff_155880_44160# gnd! 26.2fF
C54 diff_153840_44160# gnd! 26.2fF
C55 diff_151800_44160# gnd! 26.2fF
C56 diff_149760_44160# gnd! 26.2fF
C57 diff_147720_44160# gnd! 26.2fF
C58 diff_145680_44160# gnd! 26.2fF
C59 diff_143640_44160# gnd! 26.2fF
C60 diff_141600_44160# gnd! 26.2fF
C61 diff_139560_44160# gnd! 26.2fF
C62 diff_137520_44160# gnd! 26.2fF
C63 diff_135480_44160# gnd! 26.2fF
C64 diff_133440_44160# gnd! 26.2fF
C65 diff_131400_44160# gnd! 26.2fF
C66 diff_129360_44160# gnd! 26.2fF
C67 diff_127320_44160# gnd! 26.2fF
C68 diff_125280_44160# gnd! 26.2fF
C69 diff_123240_44160# gnd! 26.2fF
C70 diff_121200_44160# gnd! 26.2fF
C71 diff_119160_44160# gnd! 26.2fF
C72 diff_117120_44160# gnd! 26.2fF
C73 diff_115080_44160# gnd! 26.2fF
C74 diff_113040_44160# gnd! 26.2fF
C75 diff_111000_44160# gnd! 26.2fF
C76 diff_108960_44160# gnd! 26.2fF
C77 diff_106920_44160# gnd! 26.2fF
C78 diff_104880_44160# gnd! 26.2fF
C79 diff_102840_44160# gnd! 26.2fF
C80 diff_100800_44160# gnd! 26.2fF
C81 diff_100440_45840# gnd! 631.7fF
C82 diff_229320_46440# gnd! 24.7fF
C83 diff_227280_46440# gnd! 24.7fF
C84 diff_225240_46440# gnd! 24.7fF
C85 diff_223200_46440# gnd! 24.7fF
C86 diff_221160_46440# gnd! 24.7fF
C87 diff_219120_46440# gnd! 24.7fF
C88 diff_217080_46440# gnd! 24.7fF
C89 diff_215040_46440# gnd! 24.7fF
C90 diff_213000_46440# gnd! 24.7fF
C91 diff_210960_46440# gnd! 24.7fF
C92 diff_208920_46440# gnd! 24.7fF
C93 diff_206880_46440# gnd! 24.7fF
C94 diff_204840_46440# gnd! 24.7fF
C95 diff_202800_46440# gnd! 24.7fF
C96 diff_200760_46440# gnd! 24.7fF
C97 diff_198720_46440# gnd! 24.7fF
C98 diff_196680_46440# gnd! 24.7fF
C99 diff_194640_46440# gnd! 24.7fF
C100 diff_192600_46440# gnd! 24.7fF
C101 diff_190560_46440# gnd! 24.7fF
C102 diff_188520_46440# gnd! 24.7fF
C103 diff_186480_46440# gnd! 24.7fF
C104 diff_184440_46440# gnd! 24.7fF
C105 diff_182400_46440# gnd! 24.7fF
C106 diff_180360_46440# gnd! 24.7fF
C107 diff_178320_46440# gnd! 24.7fF
C108 diff_176280_46440# gnd! 24.7fF
C109 diff_174240_46440# gnd! 24.7fF
C110 diff_172200_46440# gnd! 24.7fF
C111 diff_170160_46440# gnd! 24.7fF
C112 diff_168120_46440# gnd! 24.7fF
C113 diff_166080_46440# gnd! 24.7fF
C114 diff_164040_46440# gnd! 24.7fF
C115 diff_162000_46440# gnd! 24.7fF
C116 diff_159960_46440# gnd! 24.7fF
C117 diff_157920_46440# gnd! 24.7fF
C118 diff_155880_46440# gnd! 24.7fF
C119 diff_153840_46440# gnd! 24.7fF
C120 diff_151800_46440# gnd! 24.7fF
C121 diff_149760_46440# gnd! 24.7fF
C122 diff_147720_46440# gnd! 24.7fF
C123 diff_145680_46440# gnd! 24.7fF
C124 diff_143640_46440# gnd! 24.7fF
C125 diff_141600_46440# gnd! 24.7fF
C126 diff_139560_46440# gnd! 24.7fF
C127 diff_137520_46440# gnd! 24.7fF
C128 diff_135480_46440# gnd! 24.7fF
C129 diff_133440_46440# gnd! 24.7fF
C130 diff_131400_46440# gnd! 24.7fF
C131 diff_129360_46440# gnd! 24.7fF
C132 diff_127320_46440# gnd! 24.7fF
C133 diff_125280_46440# gnd! 24.7fF
C134 diff_123240_46440# gnd! 24.7fF
C135 diff_121200_46440# gnd! 24.7fF
C136 diff_119160_46440# gnd! 24.7fF
C137 diff_117120_46440# gnd! 24.7fF
C138 diff_115080_46440# gnd! 24.7fF
C139 diff_113040_46440# gnd! 24.7fF
C140 diff_111000_46440# gnd! 24.7fF
C141 diff_108960_46440# gnd! 24.7fF
C142 diff_106920_46440# gnd! 24.7fF
C143 diff_104880_46440# gnd! 24.7fF
C144 diff_102840_46440# gnd! 24.7fF
C145 diff_79560_37560# gnd! 87.3fF
C146 diff_74880_37560# gnd! 94.1fF
C147 diff_87240_39840# gnd! 37.8fF
C148 diff_82560_39840# gnd! 41.1fF
C149 diff_78000_39840# gnd! 42.1fF
C150 diff_73320_39840# gnd! 42.2fF
C151 diff_100800_46440# gnd! 24.7fF
C152 diff_100440_48000# gnd! 653.0fF
C153 diff_229320_48600# gnd! 26.2fF
C154 diff_227280_48600# gnd! 26.2fF
C155 diff_225240_48600# gnd! 26.2fF
C156 diff_223200_48600# gnd! 26.2fF
C157 diff_221160_48600# gnd! 26.2fF
C158 diff_219120_48600# gnd! 26.2fF
C159 diff_217080_48600# gnd! 26.2fF
C160 diff_215040_48600# gnd! 26.2fF
C161 diff_213000_48600# gnd! 26.2fF
C162 diff_210960_48600# gnd! 26.2fF
C163 diff_208920_48600# gnd! 26.2fF
C164 diff_206880_48600# gnd! 26.2fF
C165 diff_204840_48600# gnd! 26.2fF
C166 diff_202800_48600# gnd! 26.2fF
C167 diff_200760_48600# gnd! 26.2fF
C168 diff_198720_48600# gnd! 26.2fF
C169 diff_196680_48600# gnd! 26.2fF
C170 diff_194640_48600# gnd! 26.2fF
C171 diff_192600_48600# gnd! 26.2fF
C172 diff_190560_48600# gnd! 26.2fF
C173 diff_188520_48600# gnd! 26.2fF
C174 diff_186480_48600# gnd! 26.2fF
C175 diff_184440_48600# gnd! 26.2fF
C176 diff_182400_48600# gnd! 26.2fF
C177 diff_180360_48600# gnd! 26.2fF
C178 diff_178320_48600# gnd! 26.2fF
C179 diff_176280_48600# gnd! 26.2fF
C180 diff_174240_48600# gnd! 26.2fF
C181 diff_172200_48600# gnd! 26.2fF
C182 diff_170160_48600# gnd! 26.2fF
C183 diff_168120_48600# gnd! 26.2fF
C184 diff_166080_48600# gnd! 26.2fF
C185 diff_164040_48600# gnd! 26.2fF
C186 diff_162000_48600# gnd! 26.2fF
C187 diff_159960_48600# gnd! 26.2fF
C188 diff_157920_48600# gnd! 26.2fF
C189 diff_155880_48600# gnd! 26.2fF
C190 diff_153840_48600# gnd! 26.2fF
C191 diff_151800_48600# gnd! 26.2fF
C192 diff_149760_48600# gnd! 26.2fF
C193 diff_147720_48600# gnd! 26.2fF
C194 diff_145680_48600# gnd! 26.2fF
C195 diff_143640_48600# gnd! 26.2fF
C196 diff_141600_48600# gnd! 26.2fF
C197 diff_139560_48600# gnd! 26.2fF
C198 diff_137520_48600# gnd! 26.2fF
C199 diff_135480_48600# gnd! 26.2fF
C200 diff_133440_48600# gnd! 26.2fF
C201 diff_131400_48600# gnd! 26.2fF
C202 diff_129360_48600# gnd! 26.2fF
C203 diff_127320_48600# gnd! 26.2fF
C204 diff_125280_48600# gnd! 26.2fF
C205 diff_123240_48600# gnd! 26.2fF
C206 diff_121200_48600# gnd! 26.2fF
C207 diff_119160_48600# gnd! 26.2fF
C208 diff_117120_48600# gnd! 26.2fF
C209 diff_115080_48600# gnd! 26.2fF
C210 diff_113040_48600# gnd! 26.2fF
C211 diff_111000_48600# gnd! 26.2fF
C212 diff_108960_48600# gnd! 26.2fF
C213 diff_106920_48600# gnd! 26.2fF
C214 diff_104880_48600# gnd! 26.2fF
C215 diff_102840_48600# gnd! 26.2fF
C216 diff_100800_48600# gnd! 26.2fF
C217 diff_236760_43080# gnd! 519.2fF
C218 diff_100440_43560# gnd! 598.0fF
C219 diff_281880_73800# gnd! 46.5fF
C220 diff_277440_73800# gnd! 117.6fF
C221 diff_284160_79920# gnd! 43.7fF
C222 diff_286560_90000# gnd! 46.5fF
C223 diff_273840_77640# gnd! 92.4fF
C224 diff_268680_78960# gnd! 113.8fF
C225 diff_266520_78960# gnd! 110.7fF
C226 diff_261720_78960# gnd! 122.4fF
C227 diff_277440_85200# gnd! 164.5fF
C228 diff_273840_81360# gnd! 90.0fF
C229 diff_259800_65640# gnd! 138.3fF
C230 diff_281880_88920# gnd! 145.9fF
C231 diff_277440_88920# gnd! 113.9fF
C232 diff_273840_55200# gnd! 217.4fF
C233 diff_275160_45240# gnd! 542.6fF
C234 diff_273240_54960# gnd! 457.7fF
C235 diff_284880_97680# gnd! 56.2fF
C236 diff_277920_48600# gnd! 326.9fF
C237 diff_284880_99240# gnd! 56.2fF
C238 diff_100440_50280# gnd! 622.9fF
C239 diff_229320_50880# gnd! 24.7fF
C240 diff_227280_50880# gnd! 24.7fF
C241 diff_225240_50880# gnd! 24.7fF
C242 diff_223200_50880# gnd! 24.7fF
C243 diff_221160_50880# gnd! 24.7fF
C244 diff_219120_50880# gnd! 24.7fF
C245 diff_217080_50880# gnd! 24.7fF
C246 diff_215040_50880# gnd! 24.7fF
C247 diff_213000_50880# gnd! 24.7fF
C248 diff_210960_50880# gnd! 24.7fF
C249 diff_208920_50880# gnd! 24.7fF
C250 diff_206880_50880# gnd! 24.7fF
C251 diff_204840_50880# gnd! 24.7fF
C252 diff_202800_50880# gnd! 24.7fF
C253 diff_200760_50880# gnd! 24.7fF
C254 diff_198720_50880# gnd! 24.7fF
C255 diff_196680_50880# gnd! 24.7fF
C256 diff_194640_50880# gnd! 24.7fF
C257 diff_192600_50880# gnd! 24.7fF
C258 diff_190560_50880# gnd! 24.7fF
C259 diff_188520_50880# gnd! 24.7fF
C260 diff_186480_50880# gnd! 24.7fF
C261 diff_184440_50880# gnd! 24.7fF
C262 diff_182400_50880# gnd! 24.7fF
C263 diff_180360_50880# gnd! 24.7fF
C264 diff_178320_50880# gnd! 24.7fF
C265 diff_176280_50880# gnd! 24.7fF
C266 diff_174240_50880# gnd! 24.7fF
C267 diff_172200_50880# gnd! 24.7fF
C268 diff_170160_50880# gnd! 24.7fF
C269 diff_168120_50880# gnd! 24.7fF
C270 diff_166080_50880# gnd! 24.7fF
C271 diff_164040_50880# gnd! 24.7fF
C272 diff_162000_50880# gnd! 24.7fF
C273 diff_159960_50880# gnd! 24.7fF
C274 diff_157920_50880# gnd! 24.7fF
C275 diff_155880_50880# gnd! 24.7fF
C276 diff_153840_50880# gnd! 24.7fF
C277 diff_151800_50880# gnd! 24.7fF
C278 diff_149760_50880# gnd! 24.7fF
C279 diff_147720_50880# gnd! 24.7fF
C280 diff_145680_50880# gnd! 24.7fF
C281 diff_143640_50880# gnd! 24.7fF
C282 diff_141600_50880# gnd! 24.7fF
C283 diff_139560_50880# gnd! 24.7fF
C284 diff_137520_50880# gnd! 24.7fF
C285 diff_135480_50880# gnd! 24.7fF
C286 diff_133440_50880# gnd! 24.7fF
C287 diff_131400_50880# gnd! 24.7fF
C288 diff_129360_50880# gnd! 24.7fF
C289 diff_127320_50880# gnd! 24.7fF
C290 diff_125280_50880# gnd! 24.7fF
C291 diff_123240_50880# gnd! 24.7fF
C292 diff_121200_50880# gnd! 24.7fF
C293 diff_119160_50880# gnd! 24.7fF
C294 diff_117120_50880# gnd! 24.7fF
C295 diff_115080_50880# gnd! 24.7fF
C296 diff_113040_50880# gnd! 24.7fF
C297 diff_111000_50880# gnd! 24.7fF
C298 diff_108960_50880# gnd! 24.7fF
C299 diff_106920_50880# gnd! 24.7fF
C300 diff_104880_50880# gnd! 24.7fF
C301 diff_102840_50880# gnd! 24.7fF
C302 diff_100800_50880# gnd! 24.7fF
C303 diff_229320_53040# gnd! 26.2fF
C304 diff_227280_53040# gnd! 26.2fF
C305 diff_225240_53040# gnd! 26.2fF
C306 diff_223200_53040# gnd! 26.2fF
C307 diff_221160_53040# gnd! 26.2fF
C308 diff_219120_53040# gnd! 26.2fF
C309 diff_217080_53040# gnd! 26.2fF
C310 diff_215040_53040# gnd! 26.2fF
C311 diff_213000_53040# gnd! 26.2fF
C312 diff_210960_53040# gnd! 26.2fF
C313 diff_208920_53040# gnd! 26.2fF
C314 diff_206880_53040# gnd! 26.2fF
C315 diff_204840_53040# gnd! 26.2fF
C316 diff_202800_53040# gnd! 26.2fF
C317 diff_200760_53040# gnd! 26.2fF
C318 diff_198720_53040# gnd! 26.2fF
C319 diff_196680_53040# gnd! 26.2fF
C320 diff_194640_53040# gnd! 26.2fF
C321 diff_192600_53040# gnd! 26.2fF
C322 diff_190560_53040# gnd! 26.2fF
C323 diff_188520_53040# gnd! 26.2fF
C324 diff_186480_53040# gnd! 26.2fF
C325 diff_184440_53040# gnd! 26.2fF
C326 diff_182400_53040# gnd! 26.2fF
C327 diff_180360_53040# gnd! 26.2fF
C328 diff_178320_53040# gnd! 26.2fF
C329 diff_176280_53040# gnd! 26.2fF
C330 diff_174240_53040# gnd! 26.2fF
C331 diff_172200_53040# gnd! 26.2fF
C332 diff_170160_53040# gnd! 26.2fF
C333 diff_168120_53040# gnd! 26.2fF
C334 diff_166080_53040# gnd! 26.2fF
C335 diff_164040_53040# gnd! 26.2fF
C336 diff_162000_53040# gnd! 26.2fF
C337 diff_159960_53040# gnd! 26.2fF
C338 diff_157920_53040# gnd! 26.2fF
C339 diff_155880_53040# gnd! 26.2fF
C340 diff_153840_53040# gnd! 26.2fF
C341 diff_151800_53040# gnd! 26.2fF
C342 diff_149760_53040# gnd! 26.2fF
C343 diff_147720_53040# gnd! 26.2fF
C344 diff_145680_53040# gnd! 26.2fF
C345 diff_143640_53040# gnd! 26.2fF
C346 diff_141600_53040# gnd! 26.2fF
C347 diff_139560_53040# gnd! 26.2fF
C348 diff_137520_53040# gnd! 26.2fF
C349 diff_135480_53040# gnd! 26.2fF
C350 diff_133440_53040# gnd! 26.2fF
C351 diff_131400_53040# gnd! 26.2fF
C352 diff_129360_53040# gnd! 26.2fF
C353 diff_127320_53040# gnd! 26.2fF
C354 diff_125280_53040# gnd! 26.2fF
C355 diff_123240_53040# gnd! 26.2fF
C356 diff_121200_53040# gnd! 26.2fF
C357 diff_119160_53040# gnd! 26.2fF
C358 diff_117120_53040# gnd! 26.2fF
C359 diff_115080_53040# gnd! 26.2fF
C360 diff_113040_53040# gnd! 26.2fF
C361 diff_111000_53040# gnd! 26.2fF
C362 diff_108960_53040# gnd! 26.2fF
C363 diff_106920_53040# gnd! 26.2fF
C364 diff_104880_53040# gnd! 26.2fF
C365 diff_102840_53040# gnd! 26.2fF
C366 diff_92280_45840# gnd! 112.9fF
C367 diff_90480_46440# gnd! 36.9fF
C368 diff_61320_37560# gnd! 87.3fF
C369 diff_47400_37560# gnd! 93.2fF
C370 diff_64320_39840# gnd! 41.5fF
C371 diff_59760_39840# gnd! 41.7fF
C372 diff_55080_39840# gnd! 42.6fF
C373 diff_50640_39840# gnd! 40.0fF
C374 diff_45960_39840# gnd! 41.5fF
C375 diff_42960_37560# gnd! 87.3fF
C376 diff_38280_37560# gnd! 94.1fF
C377 diff_41400_39840# gnd! 41.7fF
C378 diff_36720_39840# gnd! 42.6fF
C379 diff_32160_39840# gnd! 40.9fF
C380 diff_62160_46920# gnd! 145.3fF
C381 diff_55080_45480# gnd! 153.6fF
C382 diff_69120_47280# gnd! 138.8fF
C383 diff_69480_47880# gnd! 31.6fF
C384 diff_50040_48000# gnd! 39.8fF
C385 diff_78000_44640# gnd! 140.2fF
C386 diff_28920_45720# gnd! 141.0fF
C387 diff_81000_51000# gnd! 108.7fF
C388 diff_100800_53040# gnd! 26.2fF
C389 diff_100440_54720# gnd! 636.7fF
C390 diff_229320_55320# gnd! 24.7fF
C391 diff_227280_55320# gnd! 24.7fF
C392 diff_225240_55320# gnd! 24.7fF
C393 diff_223200_55320# gnd! 24.7fF
C394 diff_221160_55320# gnd! 24.7fF
C395 diff_219120_55320# gnd! 24.7fF
C396 diff_217080_55320# gnd! 24.7fF
C397 diff_215040_55320# gnd! 24.7fF
C398 diff_213000_55320# gnd! 24.7fF
C399 diff_210960_55320# gnd! 24.7fF
C400 diff_208920_55320# gnd! 24.7fF
C401 diff_206880_55320# gnd! 24.7fF
C402 diff_204840_55320# gnd! 24.7fF
C403 diff_202800_55320# gnd! 24.7fF
C404 diff_200760_55320# gnd! 24.7fF
C405 diff_198720_55320# gnd! 24.7fF
C406 diff_196680_55320# gnd! 24.7fF
C407 diff_194640_55320# gnd! 24.7fF
C408 diff_192600_55320# gnd! 24.7fF
C409 diff_190560_55320# gnd! 24.7fF
C410 diff_188520_55320# gnd! 24.7fF
C411 diff_186480_55320# gnd! 24.7fF
C412 diff_184440_55320# gnd! 24.7fF
C413 diff_182400_55320# gnd! 24.7fF
C414 diff_180360_55320# gnd! 24.7fF
C415 diff_178320_55320# gnd! 24.7fF
C416 diff_176280_55320# gnd! 24.7fF
C417 diff_174240_55320# gnd! 24.7fF
C418 diff_172200_55320# gnd! 24.7fF
C419 diff_170160_55320# gnd! 24.7fF
C420 diff_168120_55320# gnd! 24.7fF
C421 diff_166080_55320# gnd! 24.7fF
C422 diff_164040_55320# gnd! 24.7fF
C423 diff_162000_55320# gnd! 24.7fF
C424 diff_159960_55320# gnd! 24.7fF
C425 diff_157920_55320# gnd! 24.7fF
C426 diff_155880_55320# gnd! 24.7fF
C427 diff_153840_55320# gnd! 24.7fF
C428 diff_151800_55320# gnd! 24.7fF
C429 diff_149760_55320# gnd! 24.7fF
C430 diff_147720_55320# gnd! 24.7fF
C431 diff_145680_55320# gnd! 24.7fF
C432 diff_143640_55320# gnd! 24.7fF
C433 diff_141600_55320# gnd! 24.7fF
C434 diff_139560_55320# gnd! 24.7fF
C435 diff_137520_55320# gnd! 24.7fF
C436 diff_135480_55320# gnd! 24.7fF
C437 diff_133440_55320# gnd! 24.7fF
C438 diff_131400_55320# gnd! 24.7fF
C439 diff_129360_55320# gnd! 24.7fF
C440 diff_127320_55320# gnd! 24.7fF
C441 diff_125280_55320# gnd! 24.7fF
C442 diff_123240_55320# gnd! 24.7fF
C443 diff_121200_55320# gnd! 24.7fF
C444 diff_119160_55320# gnd! 24.7fF
C445 diff_117120_55320# gnd! 24.7fF
C446 diff_115080_55320# gnd! 24.7fF
C447 diff_113040_55320# gnd! 24.7fF
C448 diff_111000_55320# gnd! 24.7fF
C449 diff_108960_55320# gnd! 24.7fF
C450 diff_106920_55320# gnd! 24.7fF
C451 diff_104880_55320# gnd! 24.7fF
C452 diff_102840_55320# gnd! 24.7fF
C453 diff_100800_55320# gnd! 24.7fF
C454 diff_100440_56880# gnd! 652.0fF
C455 diff_229320_57480# gnd! 26.2fF
C456 diff_227280_57480# gnd! 26.2fF
C457 diff_225240_57480# gnd! 26.2fF
C458 diff_223200_57480# gnd! 26.2fF
C459 diff_221160_57480# gnd! 26.2fF
C460 diff_219120_57480# gnd! 26.2fF
C461 diff_217080_57480# gnd! 26.2fF
C462 diff_215040_57480# gnd! 26.2fF
C463 diff_213000_57480# gnd! 26.2fF
C464 diff_210960_57480# gnd! 26.2fF
C465 diff_208920_57480# gnd! 26.2fF
C466 diff_206880_57480# gnd! 26.2fF
C467 diff_204840_57480# gnd! 26.2fF
C468 diff_202800_57480# gnd! 26.2fF
C469 diff_200760_57480# gnd! 26.2fF
C470 diff_198720_57480# gnd! 26.2fF
C471 diff_196680_57480# gnd! 26.2fF
C472 diff_194640_57480# gnd! 26.2fF
C473 diff_192600_57480# gnd! 26.2fF
C474 diff_190560_57480# gnd! 26.2fF
C475 diff_188520_57480# gnd! 26.2fF
C476 diff_186480_57480# gnd! 26.2fF
C477 diff_184440_57480# gnd! 26.2fF
C478 diff_182400_57480# gnd! 26.2fF
C479 diff_180360_57480# gnd! 26.2fF
C480 diff_178320_57480# gnd! 26.2fF
C481 diff_176280_57480# gnd! 26.2fF
C482 diff_174240_57480# gnd! 26.2fF
C483 diff_172200_57480# gnd! 26.2fF
C484 diff_170160_57480# gnd! 26.2fF
C485 diff_168120_57480# gnd! 26.2fF
C486 diff_166080_57480# gnd! 26.2fF
C487 diff_164040_57480# gnd! 26.2fF
C488 diff_162000_57480# gnd! 26.2fF
C489 diff_159960_57480# gnd! 26.2fF
C490 diff_157920_57480# gnd! 26.2fF
C491 diff_155880_57480# gnd! 26.2fF
C492 diff_153840_57480# gnd! 26.2fF
C493 diff_151800_57480# gnd! 26.2fF
C494 diff_149760_57480# gnd! 26.2fF
C495 diff_147720_57480# gnd! 26.2fF
C496 diff_145680_57480# gnd! 26.2fF
C497 diff_143640_57480# gnd! 26.2fF
C498 diff_141600_57480# gnd! 26.2fF
C499 diff_139560_57480# gnd! 26.2fF
C500 diff_137520_57480# gnd! 26.2fF
C501 diff_135480_57480# gnd! 26.2fF
C502 diff_133440_57480# gnd! 26.2fF
C503 diff_131400_57480# gnd! 26.2fF
C504 diff_129360_57480# gnd! 26.2fF
C505 diff_127320_57480# gnd! 26.2fF
C506 diff_125280_57480# gnd! 26.2fF
C507 diff_123240_57480# gnd! 26.2fF
C508 diff_121200_57480# gnd! 26.2fF
C509 diff_119160_57480# gnd! 26.2fF
C510 diff_117120_57480# gnd! 26.2fF
C511 diff_115080_57480# gnd! 26.2fF
C512 diff_113040_57480# gnd! 26.2fF
C513 diff_111000_57480# gnd! 26.2fF
C514 diff_108960_57480# gnd! 26.2fF
C515 diff_106920_57480# gnd! 26.2fF
C516 diff_104880_57480# gnd! 26.2fF
C517 diff_102840_57480# gnd! 26.2fF
C518 diff_100800_57480# gnd! 26.2fF
C519 diff_236760_51960# gnd! 482.7fF
C520 diff_100440_52440# gnd! 592.4fF
C521 diff_250800_43080# gnd! 973.1fF
C522 diff_100440_59160# gnd! 621.9fF
C523 diff_229320_59760# gnd! 24.7fF
C524 diff_227280_59760# gnd! 24.7fF
C525 diff_225240_59760# gnd! 24.7fF
C526 diff_223200_59760# gnd! 24.7fF
C527 diff_221160_59760# gnd! 24.7fF
C528 diff_219120_59760# gnd! 24.7fF
C529 diff_217080_59760# gnd! 24.7fF
C530 diff_215040_59760# gnd! 24.7fF
C531 diff_213000_59760# gnd! 24.7fF
C532 diff_210960_59760# gnd! 24.7fF
C533 diff_208920_59760# gnd! 24.7fF
C534 diff_206880_59760# gnd! 24.7fF
C535 diff_204840_59760# gnd! 24.7fF
C536 diff_202800_59760# gnd! 24.7fF
C537 diff_200760_59760# gnd! 24.7fF
C538 diff_198720_59760# gnd! 24.7fF
C539 diff_196680_59760# gnd! 24.7fF
C540 diff_194640_59760# gnd! 24.7fF
C541 diff_192600_59760# gnd! 24.7fF
C542 diff_190560_59760# gnd! 24.7fF
C543 diff_188520_59760# gnd! 24.7fF
C544 diff_186480_59760# gnd! 24.7fF
C545 diff_184440_59760# gnd! 24.7fF
C546 diff_182400_59760# gnd! 24.7fF
C547 diff_180360_59760# gnd! 24.7fF
C548 diff_178320_59760# gnd! 24.7fF
C549 diff_176280_59760# gnd! 24.7fF
C550 diff_174240_59760# gnd! 24.7fF
C551 diff_172200_59760# gnd! 24.7fF
C552 diff_170160_59760# gnd! 24.7fF
C553 diff_168120_59760# gnd! 24.7fF
C554 diff_166080_59760# gnd! 24.7fF
C555 diff_164040_59760# gnd! 24.7fF
C556 diff_162000_59760# gnd! 24.7fF
C557 diff_159960_59760# gnd! 24.7fF
C558 diff_157920_59760# gnd! 24.7fF
C559 diff_155880_59760# gnd! 24.7fF
C560 diff_153840_59760# gnd! 24.7fF
C561 diff_151800_59760# gnd! 24.7fF
C562 diff_149760_59760# gnd! 24.7fF
C563 diff_147720_59760# gnd! 24.7fF
C564 diff_145680_59760# gnd! 24.7fF
C565 diff_143640_59760# gnd! 24.7fF
C566 diff_141600_59760# gnd! 24.7fF
C567 diff_139560_59760# gnd! 24.7fF
C568 diff_137520_59760# gnd! 24.7fF
C569 diff_135480_59760# gnd! 24.7fF
C570 diff_133440_59760# gnd! 24.7fF
C571 diff_131400_59760# gnd! 24.7fF
C572 diff_129360_59760# gnd! 24.7fF
C573 diff_127320_59760# gnd! 24.7fF
C574 diff_125280_59760# gnd! 24.7fF
C575 diff_123240_59760# gnd! 24.7fF
C576 diff_121200_59760# gnd! 24.7fF
C577 diff_119160_59760# gnd! 24.7fF
C578 diff_117120_59760# gnd! 24.7fF
C579 diff_115080_59760# gnd! 24.7fF
C580 diff_113040_59760# gnd! 24.7fF
C581 diff_111000_59760# gnd! 24.7fF
C582 diff_108960_59760# gnd! 24.7fF
C583 diff_106920_59760# gnd! 24.7fF
C584 diff_104880_59760# gnd! 24.7fF
C585 diff_102840_59760# gnd! 24.7fF
C586 diff_77640_48840# gnd! 105.8fF
C587 diff_69120_48720# gnd! 146.6fF
C588 diff_75600_45480# gnd! 104.1fF
C589 diff_100800_59760# gnd! 24.7fF
C590 diff_69480_49320# gnd! 88.7fF
C591 diff_47520_50040# gnd! 15.4fF
C592 diff_40440_47040# gnd! 67.7fF
C593 diff_49080_50040# gnd! 51.7fF
C594 diff_47880_47040# gnd! 150.8fF
C595 diff_49680_49200# gnd! 357.1fF
C596 cm gnd! 1310.0fF
C597 diff_236760_60720# gnd! 544.8fF
C598 diff_229320_61920# gnd! 26.2fF
C599 diff_227280_61920# gnd! 26.2fF
C600 diff_225240_61920# gnd! 26.2fF
C601 diff_223200_61920# gnd! 26.2fF
C602 diff_221160_61920# gnd! 26.2fF
C603 diff_219120_61920# gnd! 26.2fF
C604 diff_217080_61920# gnd! 26.2fF
C605 diff_215040_61920# gnd! 26.2fF
C606 diff_213000_61920# gnd! 26.2fF
C607 diff_210960_61920# gnd! 26.2fF
C608 diff_208920_61920# gnd! 26.2fF
C609 diff_206880_61920# gnd! 26.2fF
C610 diff_204840_61920# gnd! 26.2fF
C611 diff_202800_61920# gnd! 26.2fF
C612 diff_200760_61920# gnd! 26.2fF
C613 diff_198720_61920# gnd! 26.2fF
C614 diff_196680_61920# gnd! 26.2fF
C615 diff_194640_61920# gnd! 26.2fF
C616 diff_192600_61920# gnd! 26.2fF
C617 diff_190560_61920# gnd! 26.2fF
C618 diff_188520_61920# gnd! 26.2fF
C619 diff_186480_61920# gnd! 26.2fF
C620 diff_184440_61920# gnd! 26.2fF
C621 diff_182400_61920# gnd! 26.2fF
C622 diff_180360_61920# gnd! 26.2fF
C623 diff_178320_61920# gnd! 26.2fF
C624 diff_176280_61920# gnd! 26.2fF
C625 diff_174240_61920# gnd! 26.2fF
C626 diff_172200_61920# gnd! 26.2fF
C627 diff_170160_61920# gnd! 26.2fF
C628 diff_168120_61920# gnd! 26.2fF
C629 diff_166080_61920# gnd! 26.2fF
C630 diff_164040_61920# gnd! 26.2fF
C631 diff_162000_61920# gnd! 26.2fF
C632 diff_159960_61920# gnd! 26.2fF
C633 diff_157920_61920# gnd! 26.2fF
C634 diff_155880_61920# gnd! 26.2fF
C635 diff_153840_61920# gnd! 26.2fF
C636 diff_151800_61920# gnd! 26.2fF
C637 diff_149760_61920# gnd! 26.2fF
C638 diff_147720_61920# gnd! 26.2fF
C639 diff_145680_61920# gnd! 26.2fF
C640 diff_143640_61920# gnd! 26.2fF
C641 diff_141600_61920# gnd! 26.2fF
C642 diff_139560_61920# gnd! 26.2fF
C643 diff_137520_61920# gnd! 26.2fF
C644 diff_135480_61920# gnd! 26.2fF
C645 diff_133440_61920# gnd! 26.2fF
C646 diff_131400_61920# gnd! 26.2fF
C647 diff_129360_61920# gnd! 26.2fF
C648 diff_127320_61920# gnd! 26.2fF
C649 diff_125280_61920# gnd! 26.2fF
C650 diff_123240_61920# gnd! 26.2fF
C651 diff_121200_61920# gnd! 26.2fF
C652 diff_119160_61920# gnd! 26.2fF
C653 diff_117120_61920# gnd! 26.2fF
C654 diff_115080_61920# gnd! 26.2fF
C655 diff_113040_61920# gnd! 26.2fF
C656 diff_111000_61920# gnd! 26.2fF
C657 diff_108960_61920# gnd! 26.2fF
C658 diff_106920_61920# gnd! 26.2fF
C659 diff_104880_61920# gnd! 26.2fF
C660 diff_102840_61920# gnd! 26.2fF
C661 diff_100800_61920# gnd! 26.2fF
C662 diff_100440_63600# gnd! 641.1fF
C663 diff_229320_64200# gnd! 24.7fF
C664 diff_227280_64200# gnd! 24.7fF
C665 diff_225240_64200# gnd! 24.7fF
C666 diff_223200_64200# gnd! 24.7fF
C667 diff_221160_64200# gnd! 24.7fF
C668 diff_219120_64200# gnd! 24.7fF
C669 diff_217080_64200# gnd! 24.7fF
C670 diff_215040_64200# gnd! 24.7fF
C671 diff_213000_64200# gnd! 24.7fF
C672 diff_210960_64200# gnd! 24.7fF
C673 diff_208920_64200# gnd! 24.7fF
C674 diff_206880_64200# gnd! 24.7fF
C675 diff_204840_64200# gnd! 24.7fF
C676 diff_202800_64200# gnd! 24.7fF
C677 diff_200760_64200# gnd! 24.7fF
C678 diff_198720_64200# gnd! 24.7fF
C679 diff_196680_64200# gnd! 24.7fF
C680 diff_194640_64200# gnd! 24.7fF
C681 diff_192600_64200# gnd! 24.7fF
C682 diff_190560_64200# gnd! 24.7fF
C683 diff_188520_64200# gnd! 24.7fF
C684 diff_186480_64200# gnd! 24.7fF
C685 diff_184440_64200# gnd! 24.7fF
C686 diff_182400_64200# gnd! 24.7fF
C687 diff_180360_64200# gnd! 24.7fF
C688 diff_178320_64200# gnd! 24.7fF
C689 diff_176280_64200# gnd! 24.7fF
C690 diff_174240_64200# gnd! 24.7fF
C691 diff_172200_64200# gnd! 24.7fF
C692 diff_170160_64200# gnd! 24.7fF
C693 diff_168120_64200# gnd! 24.7fF
C694 diff_166080_64200# gnd! 24.7fF
C695 diff_164040_64200# gnd! 24.7fF
C696 diff_162000_64200# gnd! 24.7fF
C697 diff_159960_64200# gnd! 24.7fF
C698 diff_157920_64200# gnd! 24.7fF
C699 diff_155880_64200# gnd! 24.7fF
C700 diff_153840_64200# gnd! 24.7fF
C701 diff_151800_64200# gnd! 24.7fF
C702 diff_149760_64200# gnd! 24.7fF
C703 diff_147720_64200# gnd! 24.7fF
C704 diff_145680_64200# gnd! 24.7fF
C705 diff_143640_64200# gnd! 24.7fF
C706 diff_141600_64200# gnd! 24.7fF
C707 diff_139560_64200# gnd! 24.7fF
C708 diff_137520_64200# gnd! 24.7fF
C709 diff_135480_64200# gnd! 24.7fF
C710 diff_133440_64200# gnd! 24.7fF
C711 diff_131400_64200# gnd! 24.7fF
C712 diff_129360_64200# gnd! 24.7fF
C713 diff_127320_64200# gnd! 24.7fF
C714 diff_125280_64200# gnd! 24.7fF
C715 diff_123240_64200# gnd! 24.7fF
C716 diff_121200_64200# gnd! 24.7fF
C717 diff_119160_64200# gnd! 24.7fF
C718 diff_117120_64200# gnd! 24.7fF
C719 diff_115080_64200# gnd! 24.7fF
C720 diff_113040_64200# gnd! 24.7fF
C721 diff_111000_64200# gnd! 24.7fF
C722 diff_108960_64200# gnd! 24.7fF
C723 diff_106920_64200# gnd! 24.7fF
C724 diff_104880_64200# gnd! 24.7fF
C725 diff_102840_64200# gnd! 24.7fF
C726 diff_100800_64200# gnd! 24.7fF
C727 diff_74640_62520# gnd! 237.2fF
C728 diff_100440_65760# gnd! 652.7fF
C729 diff_229320_66360# gnd! 26.2fF
C730 diff_227280_66360# gnd! 26.2fF
C731 diff_225240_66360# gnd! 26.2fF
C732 diff_223200_66360# gnd! 26.2fF
C733 diff_221160_66360# gnd! 26.2fF
C734 diff_219120_66360# gnd! 26.2fF
C735 diff_217080_66360# gnd! 26.2fF
C736 diff_215040_66360# gnd! 26.2fF
C737 diff_213000_66360# gnd! 26.2fF
C738 diff_210960_66360# gnd! 26.2fF
C739 diff_208920_66360# gnd! 26.2fF
C740 diff_206880_66360# gnd! 26.2fF
C741 diff_204840_66360# gnd! 26.2fF
C742 diff_202800_66360# gnd! 26.2fF
C743 diff_200760_66360# gnd! 26.2fF
C744 diff_198720_66360# gnd! 26.2fF
C745 diff_196680_66360# gnd! 26.2fF
C746 diff_194640_66360# gnd! 26.2fF
C747 diff_192600_66360# gnd! 26.2fF
C748 diff_190560_66360# gnd! 26.2fF
C749 diff_188520_66360# gnd! 26.2fF
C750 diff_186480_66360# gnd! 26.2fF
C751 diff_184440_66360# gnd! 26.2fF
C752 diff_182400_66360# gnd! 26.2fF
C753 diff_180360_66360# gnd! 26.2fF
C754 diff_178320_66360# gnd! 26.2fF
C755 diff_176280_66360# gnd! 26.2fF
C756 diff_174240_66360# gnd! 26.2fF
C757 diff_172200_66360# gnd! 26.2fF
C758 diff_170160_66360# gnd! 26.2fF
C759 diff_168120_66360# gnd! 26.2fF
C760 diff_166080_66360# gnd! 26.2fF
C761 diff_164040_66360# gnd! 26.2fF
C762 diff_162000_66360# gnd! 26.2fF
C763 diff_159960_66360# gnd! 26.2fF
C764 diff_157920_66360# gnd! 26.2fF
C765 diff_155880_66360# gnd! 26.2fF
C766 diff_153840_66360# gnd! 26.2fF
C767 diff_151800_66360# gnd! 26.2fF
C768 diff_149760_66360# gnd! 26.2fF
C769 diff_147720_66360# gnd! 26.2fF
C770 diff_145680_66360# gnd! 26.2fF
C771 diff_143640_66360# gnd! 26.2fF
C772 diff_141600_66360# gnd! 26.2fF
C773 diff_139560_66360# gnd! 26.2fF
C774 diff_137520_66360# gnd! 26.2fF
C775 diff_135480_66360# gnd! 26.2fF
C776 diff_133440_66360# gnd! 26.2fF
C777 diff_131400_66360# gnd! 26.2fF
C778 diff_129360_66360# gnd! 26.2fF
C779 diff_127320_66360# gnd! 26.2fF
C780 diff_125280_66360# gnd! 26.2fF
C781 diff_123240_66360# gnd! 26.2fF
C782 diff_121200_66360# gnd! 26.2fF
C783 diff_119160_66360# gnd! 26.2fF
C784 diff_117120_66360# gnd! 26.2fF
C785 diff_115080_66360# gnd! 26.2fF
C786 diff_113040_66360# gnd! 26.2fF
C787 diff_111000_66360# gnd! 26.2fF
C788 diff_108960_66360# gnd! 26.2fF
C789 diff_106920_66360# gnd! 26.2fF
C790 diff_104880_66360# gnd! 26.2fF
C791 diff_102840_66360# gnd! 26.2fF
C792 diff_89160_65640# gnd! 10.8fF
C793 diff_89760_63840# gnd! 124.6fF
C794 diff_100800_66360# gnd! 26.2fF
C795 diff_100440_61320# gnd! 597.6fF
C796 diff_100440_68040# gnd! 622.9fF
C797 diff_229320_68640# gnd! 24.7fF
C798 diff_227280_68640# gnd! 24.7fF
C799 diff_225240_68640# gnd! 24.7fF
C800 diff_223200_68640# gnd! 24.7fF
C801 diff_221160_68640# gnd! 24.7fF
C802 diff_219120_68640# gnd! 24.7fF
C803 diff_217080_68640# gnd! 24.7fF
C804 diff_215040_68640# gnd! 24.7fF
C805 diff_213000_68640# gnd! 24.7fF
C806 diff_210960_68640# gnd! 24.7fF
C807 diff_208920_68640# gnd! 24.7fF
C808 diff_206880_68640# gnd! 24.7fF
C809 diff_204840_68640# gnd! 24.7fF
C810 diff_202800_68640# gnd! 24.7fF
C811 diff_200760_68640# gnd! 24.7fF
C812 diff_198720_68640# gnd! 24.7fF
C813 diff_196680_68640# gnd! 24.7fF
C814 diff_194640_68640# gnd! 24.7fF
C815 diff_192600_68640# gnd! 24.7fF
C816 diff_190560_68640# gnd! 24.7fF
C817 diff_188520_68640# gnd! 24.7fF
C818 diff_186480_68640# gnd! 24.7fF
C819 diff_184440_68640# gnd! 24.7fF
C820 diff_182400_68640# gnd! 24.7fF
C821 diff_180360_68640# gnd! 24.7fF
C822 diff_178320_68640# gnd! 24.7fF
C823 diff_176280_68640# gnd! 24.7fF
C824 diff_174240_68640# gnd! 24.7fF
C825 diff_172200_68640# gnd! 24.7fF
C826 diff_170160_68640# gnd! 24.7fF
C827 diff_168120_68640# gnd! 24.7fF
C828 diff_166080_68640# gnd! 24.7fF
C829 diff_164040_68640# gnd! 24.7fF
C830 diff_162000_68640# gnd! 24.7fF
C831 diff_159960_68640# gnd! 24.7fF
C832 diff_157920_68640# gnd! 24.7fF
C833 diff_155880_68640# gnd! 24.7fF
C834 diff_153840_68640# gnd! 24.7fF
C835 diff_151800_68640# gnd! 24.7fF
C836 diff_149760_68640# gnd! 24.7fF
C837 diff_147720_68640# gnd! 24.7fF
C838 diff_145680_68640# gnd! 24.7fF
C839 diff_143640_68640# gnd! 24.7fF
C840 diff_141600_68640# gnd! 24.7fF
C841 diff_139560_68640# gnd! 24.7fF
C842 diff_137520_68640# gnd! 24.7fF
C843 diff_135480_68640# gnd! 24.7fF
C844 diff_133440_68640# gnd! 24.7fF
C845 diff_131400_68640# gnd! 24.7fF
C846 diff_129360_68640# gnd! 24.7fF
C847 diff_127320_68640# gnd! 24.7fF
C848 diff_125280_68640# gnd! 24.7fF
C849 diff_123240_68640# gnd! 24.7fF
C850 diff_121200_68640# gnd! 24.7fF
C851 diff_119160_68640# gnd! 24.7fF
C852 diff_117120_68640# gnd! 24.7fF
C853 diff_115080_68640# gnd! 24.7fF
C854 diff_113040_68640# gnd! 24.7fF
C855 diff_111000_68640# gnd! 24.7fF
C856 diff_108960_68640# gnd! 24.7fF
C857 diff_106920_68640# gnd! 24.7fF
C858 diff_104880_68640# gnd! 24.7fF
C859 diff_102840_68640# gnd! 24.7fF
C860 diff_100800_68640# gnd! 24.7fF
C861 diff_236760_69600# gnd! 481.1fF
C862 diff_229320_70800# gnd! 26.2fF
C863 diff_227280_70800# gnd! 26.2fF
C864 diff_225240_70800# gnd! 26.2fF
C865 diff_223200_70800# gnd! 26.2fF
C866 diff_221160_70800# gnd! 26.2fF
C867 diff_219120_70800# gnd! 26.2fF
C868 diff_217080_70800# gnd! 26.2fF
C869 diff_215040_70800# gnd! 26.2fF
C870 diff_213000_70800# gnd! 26.2fF
C871 diff_210960_70800# gnd! 26.2fF
C872 diff_208920_70800# gnd! 26.2fF
C873 diff_206880_70800# gnd! 26.2fF
C874 diff_204840_70800# gnd! 26.2fF
C875 diff_202800_70800# gnd! 26.2fF
C876 diff_200760_70800# gnd! 26.2fF
C877 diff_198720_70800# gnd! 26.2fF
C878 diff_196680_70800# gnd! 26.2fF
C879 diff_194640_70800# gnd! 26.2fF
C880 diff_192600_70800# gnd! 26.2fF
C881 diff_190560_70800# gnd! 26.2fF
C882 diff_188520_70800# gnd! 26.2fF
C883 diff_186480_70800# gnd! 26.2fF
C884 diff_184440_70800# gnd! 26.2fF
C885 diff_182400_70800# gnd! 26.2fF
C886 diff_180360_70800# gnd! 26.2fF
C887 diff_178320_70800# gnd! 26.2fF
C888 diff_176280_70800# gnd! 26.2fF
C889 diff_174240_70800# gnd! 26.2fF
C890 diff_172200_70800# gnd! 26.2fF
C891 diff_170160_70800# gnd! 26.2fF
C892 diff_168120_70800# gnd! 26.2fF
C893 diff_166080_70800# gnd! 26.2fF
C894 diff_164040_70800# gnd! 26.2fF
C895 diff_162000_70800# gnd! 26.2fF
C896 diff_159960_70800# gnd! 26.2fF
C897 diff_157920_70800# gnd! 26.2fF
C898 diff_155880_70800# gnd! 26.2fF
C899 diff_153840_70800# gnd! 26.2fF
C900 diff_151800_70800# gnd! 26.2fF
C901 diff_149760_70800# gnd! 26.2fF
C902 diff_147720_70800# gnd! 26.2fF
C903 diff_145680_70800# gnd! 26.2fF
C904 diff_143640_70800# gnd! 26.2fF
C905 diff_141600_70800# gnd! 26.2fF
C906 diff_139560_70800# gnd! 26.2fF
C907 diff_137520_70800# gnd! 26.2fF
C908 diff_135480_70800# gnd! 26.2fF
C909 diff_133440_70800# gnd! 26.2fF
C910 diff_131400_70800# gnd! 26.2fF
C911 diff_129360_70800# gnd! 26.2fF
C912 diff_127320_70800# gnd! 26.2fF
C913 diff_125280_70800# gnd! 26.2fF
C914 diff_123240_70800# gnd! 26.2fF
C915 diff_121200_70800# gnd! 26.2fF
C916 diff_119160_70800# gnd! 26.2fF
C917 diff_117120_70800# gnd! 26.2fF
C918 diff_115080_70800# gnd! 26.2fF
C919 diff_113040_70800# gnd! 26.2fF
C920 diff_111000_70800# gnd! 26.2fF
C921 diff_108960_70800# gnd! 26.2fF
C922 diff_106920_70800# gnd! 26.2fF
C923 diff_104880_70800# gnd! 26.2fF
C924 diff_102840_70800# gnd! 26.2fF
C925 diff_90480_65640# gnd! 78.3fF
C926 diff_100800_70800# gnd! 26.2fF
C927 diff_100440_72480# gnd! 639.6fF
C928 diff_229320_73080# gnd! 24.7fF
C929 diff_227280_73080# gnd! 24.7fF
C930 diff_225240_73080# gnd! 24.7fF
C931 diff_223200_73080# gnd! 24.7fF
C932 diff_221160_73080# gnd! 24.7fF
C933 diff_219120_73080# gnd! 24.7fF
C934 diff_217080_73080# gnd! 24.7fF
C935 diff_215040_73080# gnd! 24.7fF
C936 diff_213000_73080# gnd! 24.7fF
C937 diff_210960_73080# gnd! 24.7fF
C938 diff_208920_73080# gnd! 24.7fF
C939 diff_206880_73080# gnd! 24.7fF
C940 diff_204840_73080# gnd! 24.7fF
C941 diff_202800_73080# gnd! 24.7fF
C942 diff_200760_73080# gnd! 24.7fF
C943 diff_198720_73080# gnd! 24.7fF
C944 diff_196680_73080# gnd! 24.7fF
C945 diff_194640_73080# gnd! 24.7fF
C946 diff_192600_73080# gnd! 24.7fF
C947 diff_190560_73080# gnd! 24.7fF
C948 diff_188520_73080# gnd! 24.7fF
C949 diff_186480_73080# gnd! 24.7fF
C950 diff_184440_73080# gnd! 24.7fF
C951 diff_182400_73080# gnd! 24.7fF
C952 diff_180360_73080# gnd! 24.7fF
C953 diff_178320_73080# gnd! 24.7fF
C954 diff_176280_73080# gnd! 24.7fF
C955 diff_174240_73080# gnd! 24.7fF
C956 diff_172200_73080# gnd! 24.7fF
C957 diff_170160_73080# gnd! 24.7fF
C958 diff_168120_73080# gnd! 24.7fF
C959 diff_166080_73080# gnd! 24.7fF
C960 diff_164040_73080# gnd! 24.7fF
C961 diff_162000_73080# gnd! 24.7fF
C962 diff_159960_73080# gnd! 24.7fF
C963 diff_157920_73080# gnd! 24.7fF
C964 diff_155880_73080# gnd! 24.7fF
C965 diff_153840_73080# gnd! 24.7fF
C966 diff_151800_73080# gnd! 24.7fF
C967 diff_149760_73080# gnd! 24.7fF
C968 diff_147720_73080# gnd! 24.7fF
C969 diff_145680_73080# gnd! 24.7fF
C970 diff_143640_73080# gnd! 24.7fF
C971 diff_141600_73080# gnd! 24.7fF
C972 diff_139560_73080# gnd! 24.7fF
C973 diff_137520_73080# gnd! 24.7fF
C974 diff_135480_73080# gnd! 24.7fF
C975 diff_133440_73080# gnd! 24.7fF
C976 diff_131400_73080# gnd! 24.7fF
C977 diff_129360_73080# gnd! 24.7fF
C978 diff_127320_73080# gnd! 24.7fF
C979 diff_125280_73080# gnd! 24.7fF
C980 diff_123240_73080# gnd! 24.7fF
C981 diff_121200_73080# gnd! 24.7fF
C982 diff_119160_73080# gnd! 24.7fF
C983 diff_117120_73080# gnd! 24.7fF
C984 diff_115080_73080# gnd! 24.7fF
C985 diff_113040_73080# gnd! 24.7fF
C986 diff_111000_73080# gnd! 24.7fF
C987 diff_108960_73080# gnd! 24.7fF
C988 diff_106920_73080# gnd! 24.7fF
C989 diff_104880_73080# gnd! 24.7fF
C990 diff_102840_73080# gnd! 24.7fF
C991 diff_100800_73080# gnd! 24.7fF
C992 diff_100440_74640# gnd! 652.7fF
C993 diff_229320_75240# gnd! 26.2fF
C994 diff_227280_75240# gnd! 26.2fF
C995 diff_225240_75240# gnd! 26.2fF
C996 diff_223200_75240# gnd! 26.2fF
C997 diff_221160_75240# gnd! 26.2fF
C998 diff_219120_75240# gnd! 26.2fF
C999 diff_217080_75240# gnd! 26.2fF
C1000 diff_215040_75240# gnd! 26.2fF
C1001 diff_213000_75240# gnd! 26.2fF
C1002 diff_210960_75240# gnd! 26.2fF
C1003 diff_208920_75240# gnd! 26.2fF
C1004 diff_206880_75240# gnd! 26.2fF
C1005 diff_204840_75240# gnd! 26.2fF
C1006 diff_202800_75240# gnd! 26.2fF
C1007 diff_200760_75240# gnd! 26.2fF
C1008 diff_198720_75240# gnd! 26.2fF
C1009 diff_196680_75240# gnd! 26.2fF
C1010 diff_194640_75240# gnd! 26.2fF
C1011 diff_192600_75240# gnd! 26.2fF
C1012 diff_190560_75240# gnd! 26.2fF
C1013 diff_188520_75240# gnd! 26.2fF
C1014 diff_186480_75240# gnd! 26.2fF
C1015 diff_184440_75240# gnd! 26.2fF
C1016 diff_182400_75240# gnd! 26.2fF
C1017 diff_180360_75240# gnd! 26.2fF
C1018 diff_178320_75240# gnd! 26.2fF
C1019 diff_176280_75240# gnd! 26.2fF
C1020 diff_174240_75240# gnd! 26.2fF
C1021 diff_172200_75240# gnd! 26.2fF
C1022 diff_170160_75240# gnd! 26.2fF
C1023 diff_168120_75240# gnd! 26.2fF
C1024 diff_166080_75240# gnd! 26.2fF
C1025 diff_164040_75240# gnd! 26.2fF
C1026 diff_162000_75240# gnd! 26.2fF
C1027 diff_159960_75240# gnd! 26.2fF
C1028 diff_157920_75240# gnd! 26.2fF
C1029 diff_155880_75240# gnd! 26.2fF
C1030 diff_153840_75240# gnd! 26.2fF
C1031 diff_151800_75240# gnd! 26.2fF
C1032 diff_149760_75240# gnd! 26.2fF
C1033 diff_147720_75240# gnd! 26.2fF
C1034 diff_145680_75240# gnd! 26.2fF
C1035 diff_143640_75240# gnd! 26.2fF
C1036 diff_141600_75240# gnd! 26.2fF
C1037 diff_139560_75240# gnd! 26.2fF
C1038 diff_137520_75240# gnd! 26.2fF
C1039 diff_135480_75240# gnd! 26.2fF
C1040 diff_133440_75240# gnd! 26.2fF
C1041 diff_131400_75240# gnd! 26.2fF
C1042 diff_129360_75240# gnd! 26.2fF
C1043 diff_127320_75240# gnd! 26.2fF
C1044 diff_125280_75240# gnd! 26.2fF
C1045 diff_123240_75240# gnd! 26.2fF
C1046 diff_121200_75240# gnd! 26.2fF
C1047 diff_119160_75240# gnd! 26.2fF
C1048 diff_117120_75240# gnd! 26.2fF
C1049 diff_115080_75240# gnd! 26.2fF
C1050 diff_113040_75240# gnd! 26.2fF
C1051 diff_111000_75240# gnd! 26.2fF
C1052 diff_108960_75240# gnd! 26.2fF
C1053 diff_106920_75240# gnd! 26.2fF
C1054 diff_104880_75240# gnd! 26.2fF
C1055 diff_102840_75240# gnd! 26.2fF
C1056 diff_100800_75240# gnd! 26.2fF
C1057 diff_86640_69120# gnd! 97.8fF
C1058 diff_84000_37560# gnd! 212.4fF
C1059 diff_100440_70200# gnd! 600.3fF
C1060 diff_252960_89400# gnd! 107.9fF
C1061 diff_273840_92640# gnd! 91.8fF
C1062 diff_252960_91560# gnd! 106.8fF
C1063 diff_283200_105600# gnd! 373.6fF
C1064 diff_283200_107520# gnd! 75.7fF
C1065 diff_277440_100200# gnd! 185.6fF
C1066 diff_273840_96480# gnd! 92.6fF
C1067 diff_286560_112440# gnd! 49.8fF
C1068 diff_277440_104040# gnd! 182.7fF
C1069 diff_253080_96840# gnd! 101.7fF
C1070 diff_253080_99120# gnd! 109.8fF
C1071 diff_253080_103560# gnd! 104.8fF
C1072 diff_273840_107760# gnd! 86.6fF
C1073 diff_253080_105840# gnd! 104.0fF
C1074 diff_253200_111120# gnd! 101.9fF
C1075 diff_277440_115320# gnd! 104.9fF
C1076 diff_273840_111480# gnd! 85.9fF
C1077 diff_253080_113280# gnd! 108.9fF
C1078 diff_281880_113640# gnd! 148.5fF
C1079 diff_284160_122760# gnd! 42.3fF
C1080 diff_277440_118920# gnd! 165.5fF
C1081 diff_281880_129240# gnd! 43.7fF
C1082 diff_253080_117840# gnd! 114.0fF
C1083 diff_273840_122880# gnd! 91.0fF
C1084 diff_253080_120120# gnd! 107.1fF
C1085 diff_100440_76920# gnd! 622.9fF
C1086 diff_90480_76920# gnd! 128.8fF
C1087 diff_28440_46560# gnd! 58.9fF
C1088 diff_33840_37560# gnd! 430.5fF
C1089 reset gnd! 1008.9fF
C1090 diff_48000_61440# gnd! 91.6fF
C1091 diff_49800_71520# gnd! 51.5fF
C1092 diff_69480_76200# gnd! 135.1fF
C1093 diff_229320_77520# gnd! 41.3fF
C1094 diff_227280_77520# gnd! 41.9fF
C1095 diff_221160_77520# gnd! 41.3fF
C1096 diff_219120_77520# gnd! 41.9fF
C1097 diff_213000_77520# gnd! 41.3fF
C1098 diff_210960_77520# gnd! 41.9fF
C1099 diff_204840_77520# gnd! 41.3fF
C1100 diff_202800_77520# gnd! 41.9fF
C1101 diff_196680_77520# gnd! 41.3fF
C1102 diff_194640_77520# gnd! 41.9fF
C1103 diff_188520_77520# gnd! 41.3fF
C1104 diff_186480_77520# gnd! 41.9fF
C1105 diff_180360_77520# gnd! 41.3fF
C1106 diff_178320_77520# gnd! 41.9fF
C1107 diff_172200_77520# gnd! 41.3fF
C1108 diff_170160_77520# gnd! 41.9fF
C1109 diff_164040_77520# gnd! 41.3fF
C1110 diff_162000_77520# gnd! 41.9fF
C1111 diff_155880_77520# gnd! 41.3fF
C1112 diff_153840_77520# gnd! 41.9fF
C1113 diff_147720_77520# gnd! 41.3fF
C1114 diff_145680_77520# gnd! 41.9fF
C1115 diff_139560_77520# gnd! 41.3fF
C1116 diff_137520_77520# gnd! 41.9fF
C1117 diff_131400_77520# gnd! 41.3fF
C1118 diff_129360_77520# gnd! 41.9fF
C1119 diff_123240_77520# gnd! 41.3fF
C1120 diff_121200_77520# gnd! 41.9fF
C1121 diff_115080_77520# gnd! 41.3fF
C1122 diff_113040_77520# gnd! 41.9fF
C1123 diff_106920_77520# gnd! 40.3fF
C1124 diff_104880_77520# gnd! 41.1fF
C1125 diff_81600_78720# gnd! 14.4fF
C1126 diff_69600_78240# gnd! 69.5fF
C1127 diff_70080_67920# gnd! 147.1fF
C1128 diff_69480_55680# gnd! 265.6fF
C1129 diff_91920_42120# gnd! 1212.7fF
C1130 diff_82560_78240# gnd! 167.2fF
C1131 diff_277440_130800# gnd! 115.5fF
C1132 diff_273840_127440# gnd! 89.4fF
C1133 diff_252600_124320# gnd! 141.7fF
C1134 diff_256800_128160# gnd! 88.2fF
C1135 diff_270840_139200# gnd! 37.2fF
C1136 diff_260520_137280# gnd! 92.6fF
C1137 diff_260160_136800# gnd! 97.9fF
C1138 diff_262680_141120# gnd! 91.0fF
C1139 diff_272280_84480# gnd! 365.9fF
C1140 diff_276720_145680# gnd! 49.5fF
C1141 diff_258960_146400# gnd! 78.8fF
C1142 diff_281280_113400# gnd! 303.0fF
C1143 diff_276840_149760# gnd! 49.5fF
C1144 diff_276840_154080# gnd! 48.3fF
C1145 diff_225240_77520# gnd! 53.1fF
C1146 diff_223200_77520# gnd! 53.0fF
C1147 diff_225840_84960# gnd! 42.5fF
C1148 diff_217080_77520# gnd! 53.1fF
C1149 diff_215040_77520# gnd! 53.0fF
C1150 diff_217680_84960# gnd! 42.5fF
C1151 diff_208920_77520# gnd! 53.1fF
C1152 diff_206880_77520# gnd! 53.0fF
C1153 diff_209520_84960# gnd! 42.5fF
C1154 diff_200760_77520# gnd! 53.1fF
C1155 diff_198720_77520# gnd! 53.0fF
C1156 diff_201360_84960# gnd! 42.5fF
C1157 diff_192600_77520# gnd! 53.1fF
C1158 diff_190560_77520# gnd! 53.0fF
C1159 diff_193200_84960# gnd! 42.5fF
C1160 diff_184440_77520# gnd! 53.1fF
C1161 diff_182400_77520# gnd! 53.0fF
C1162 diff_185040_84960# gnd! 42.5fF
C1163 diff_176280_77520# gnd! 53.1fF
C1164 diff_174240_77520# gnd! 53.0fF
C1165 diff_176880_84960# gnd! 42.5fF
C1166 diff_168120_77520# gnd! 53.1fF
C1167 diff_166080_77520# gnd! 53.0fF
C1168 diff_168720_84960# gnd! 42.5fF
C1169 diff_159960_77520# gnd! 53.1fF
C1170 diff_157920_77520# gnd! 53.0fF
C1171 diff_160560_84960# gnd! 42.5fF
C1172 diff_151800_77520# gnd! 53.1fF
C1173 diff_149760_77520# gnd! 53.0fF
C1174 diff_152400_84960# gnd! 42.5fF
C1175 diff_143640_77520# gnd! 53.1fF
C1176 diff_141600_77520# gnd! 53.0fF
C1177 diff_144240_84960# gnd! 42.5fF
C1178 diff_135480_77520# gnd! 53.1fF
C1179 diff_133440_77520# gnd! 53.0fF
C1180 diff_136080_84960# gnd! 42.5fF
C1181 diff_127320_77520# gnd! 53.1fF
C1182 diff_125280_77520# gnd! 53.0fF
C1183 diff_127920_84960# gnd! 42.5fF
C1184 diff_119160_77520# gnd! 53.1fF
C1185 diff_117120_77520# gnd! 53.0fF
C1186 diff_119760_84960# gnd! 42.5fF
C1187 diff_111000_77520# gnd! 53.1fF
C1188 diff_108960_77520# gnd! 53.0fF
C1189 diff_111600_84960# gnd! 42.5fF
C1190 diff_55800_76560# gnd! 136.6fF
C1191 diff_42120_72840# gnd! 98.6fF
C1192 diff_53640_77640# gnd! 127.9fF
C1193 diff_33960_53280# gnd! 392.4fF
C1194 diff_40920_47640# gnd! 209.4fF
C1195 diff_100800_77520# gnd! 47.9fF
C1196 diff_103320_85080# gnd! 46.8fF
C1197 diff_102480_84960# gnd! 55.4fF
C1198 diff_99720_83640# gnd! 103.4fF
C1199 diff_221760_82920# gnd! 109.8fF
C1200 diff_205440_82920# gnd! 112.1fF
C1201 diff_189120_82920# gnd! 112.1fF
C1202 diff_172800_82920# gnd! 112.3fF
C1203 diff_156480_82920# gnd! 108.0fF
C1204 diff_140160_82920# gnd! 108.0fF
C1205 diff_123840_82920# gnd! 114.1fF
C1206 diff_107520_82680# gnd! 112.7fF
C1207 diff_213600_82920# gnd! 114.7fF
C1208 diff_225960_90720# gnd! 122.5fF
C1209 diff_197280_82920# gnd! 114.7fF
C1210 diff_217680_90720# gnd! 127.3fF
C1211 diff_209520_90720# gnd! 125.2fF
C1212 diff_201360_90720# gnd! 127.3fF
C1213 diff_180960_82920# gnd! 115.0fF
C1214 diff_193200_90720# gnd! 125.2fF
C1215 diff_185160_90720# gnd! 127.3fF
C1216 diff_164640_82920# gnd! 110.9fF
C1217 diff_177000_90720# gnd! 125.2fF
C1218 diff_168720_90840# gnd! 123.3fF
C1219 diff_148320_82920# gnd! 110.4fF
C1220 diff_160560_90840# gnd! 121.2fF
C1221 diff_152400_90840# gnd! 123.3fF
C1222 diff_132000_82920# gnd! 117.5fF
C1223 diff_144240_90840# gnd! 121.2fF
C1224 diff_115680_82920# gnd! 114.7fF
C1225 diff_127800_90600# gnd! 129.2fF
C1226 diff_119760_90720# gnd! 127.3fF
C1227 diff_103680_90360# gnd! 124.5fF
C1228 diff_135960_90600# gnd! 129.6fF
C1229 diff_111600_90720# gnd! 125.6fF
C1230 diff_221760_92760# gnd! 111.9fF
C1231 diff_213480_92760# gnd! 113.7fF
C1232 diff_205320_92760# gnd! 113.1fF
C1233 diff_197160_92760# gnd! 113.7fF
C1234 diff_189000_92760# gnd! 113.1fF
C1235 diff_180960_92760# gnd! 113.7fF
C1236 diff_172800_92760# gnd! 113.1fF
C1237 diff_164520_92880# gnd! 109.7fF
C1238 diff_156360_92880# gnd! 109.2fF
C1239 diff_148200_92880# gnd! 109.7fF
C1240 diff_140040_92880# gnd! 109.2fF
C1241 diff_131760_92640# gnd! 116.6fF
C1242 diff_123600_92640# gnd! 117.1fF
C1243 diff_44760_77160# gnd! 78.1fF
C1244 diff_49680_79800# gnd! 136.7fF
C1245 diff_89880_88800# gnd! 111.5fF
C1246 diff_115560_92760# gnd! 113.7fF
C1247 diff_107400_92760# gnd! 113.1fF
C1248 diff_229920_82920# gnd! 137.1fF
C1249 diff_205680_90720# gnd! 259.2fF
C1250 diff_189360_90720# gnd! 259.6fF
C1251 diff_173160_90720# gnd! 260.2fF
C1252 diff_156720_90720# gnd! 264.9fF
C1253 diff_140400_90720# gnd! 263.6fF
C1254 diff_123960_90720# gnd! 250.6fF
C1255 diff_107760_90720# gnd! 257.7fF
C1256 diff_99960_89640# gnd! 314.6fF
C1257 diff_222120_90720# gnd! 265.1fF
C1258 diff_213840_90840# gnd! 288.9fF
C1259 diff_197520_90840# gnd! 287.2fF
C1260 diff_181320_90840# gnd! 289.6fF
C1261 diff_164880_90840# gnd! 289.1fF
C1262 diff_148560_90720# gnd! 293.2fF
C1263 diff_132120_90480# gnd! 285.3fF
C1264 diff_115920_90840# gnd! 282.6fF
C1265 diff_112440_96360# gnd! 757.2fF
C1266 diff_80160_88800# gnd! 110.4fF
C1267 diff_48120_80160# gnd! 151.9fF
C1268 diff_64680_88800# gnd! 111.5fF
C1269 diff_41160_85320# gnd! 61.3fF
C1270 diff_56760_85560# gnd! 100.9fF
C1271 diff_101400_96240# gnd! 823.9fF
C1272 diff_199680_100800# gnd! 296.7fF
C1273 diff_167040_100800# gnd! 331.5fF
C1274 diff_62400_47520# gnd! 849.3fF
C1275 diff_134400_100800# gnd! 290.6fF
C1276 diff_99960_108720# gnd! 267.7fF
C1277 diff_49440_88920# gnd! 110.4fF
C1278 diff_82920_103920# gnd! 391.8fF
C1279 diff_80280_96720# gnd! 130.1fF
C1280 diff_96720_108360# gnd! 107.7fF
C1281 diff_90120_96840# gnd! 193.8fF
C1282 diff_216000_98520# gnd! 470.1fF
C1283 diff_199680_98400# gnd! 559.2fF
C1284 diff_56400_47520# gnd! 986.9fF
C1285 diff_183480_98400# gnd! 529.8fF
C1286 diff_167040_98400# gnd! 532.3fF
C1287 diff_150720_98400# gnd! 574.9fF
C1288 diff_134280_112200# gnd! 548.7fF
C1289 diff_118080_98520# gnd! 507.2fF
C1290 diff_41160_86760# gnd! 680.4fF
C1291 diff_68280_103440# gnd! 407.4fF
C1292 diff_64800_96720# gnd! 120.0fF
C1293 diff_54360_101760# gnd! 558.4fF
C1294 diff_49680_96720# gnd! 112.5fF
C1295 io0 gnd! 2887.2fF
C1296 diff_44640_90240# gnd! 452.9fF
C1297 diff_40680_69240# gnd! 589.3fF
C1298 io1 gnd! 2793.0fF
C1299 io2 gnd! 2636.2fF
C1300 io3 gnd! 2527.4fF
C1301 diff_101640_96840# gnd! 534.7fF
C1302 diff_101160_115320# gnd! 800.4fF
C1303 diff_80280_108720# gnd! 222.6fF
C1304 diff_64800_108720# gnd! 221.8fF
C1305 diff_49320_108720# gnd! 216.4fF
C1306 diff_33720_108720# gnd! 216.7fF
C1307 diff_106320_94080# gnd! 1157.4fF
C1308 diff_103320_91920# gnd! 1257.7fF
C1309 diff_99480_122520# gnd! 1372.5fF
C1310 diff_222120_120600# gnd! 269.5fF
C1311 diff_225840_126600# gnd! 42.2fF
C1312 diff_213840_120720# gnd! 294.8fF
C1313 diff_221760_118080# gnd! 105.1fF
C1314 diff_217680_126600# gnd! 42.2fF
C1315 diff_205680_120720# gnd! 257.9fF
C1316 diff_213480_118080# gnd! 106.6fF
C1317 diff_209520_126600# gnd! 42.2fF
C1318 diff_197520_120720# gnd! 291.9fF
C1319 diff_205320_118080# gnd! 106.2fF
C1320 diff_201360_126600# gnd! 42.2fF
C1321 diff_189360_120720# gnd! 257.9fF
C1322 diff_197160_118080# gnd! 106.6fF
C1323 diff_193200_126600# gnd! 42.2fF
C1324 diff_181320_120720# gnd! 290.2fF
C1325 diff_189000_118080# gnd! 106.2fF
C1326 diff_185040_126600# gnd! 42.2fF
C1327 diff_173160_120720# gnd! 258.3fF
C1328 diff_180960_118080# gnd! 106.6fF
C1329 diff_176880_126600# gnd! 42.2fF
C1330 diff_164880_120600# gnd! 292.5fF
C1331 diff_172800_118080# gnd! 106.2fF
C1332 diff_168720_126600# gnd! 42.2fF
C1333 diff_156720_120600# gnd! 264.0fF
C1334 diff_164520_118080# gnd! 102.6fF
C1335 diff_160560_126600# gnd! 42.2fF
C1336 diff_148560_120600# gnd! 296.4fF
C1337 diff_156360_118080# gnd! 102.2fF
C1338 diff_152400_126600# gnd! 42.2fF
C1339 diff_140400_120600# gnd! 264.0fF
C1340 diff_148200_118080# gnd! 102.6fF
C1341 diff_144240_126600# gnd! 42.2fF
C1342 diff_132120_120840# gnd! 290.3fF
C1343 diff_140040_118080# gnd! 102.2fF
C1344 diff_136080_126600# gnd! 42.2fF
C1345 diff_123960_120840# gnd! 250.3fF
C1346 diff_131760_118080# gnd! 107.6fF
C1347 diff_127920_126600# gnd! 42.2fF
C1348 diff_115920_120720# gnd! 285.7fF
C1349 diff_123600_118080# gnd! 110.2fF
C1350 diff_119760_126600# gnd! 42.2fF
C1351 diff_107760_120720# gnd! 258.2fF
C1352 diff_115560_118080# gnd! 106.6fF
C1353 diff_111600_126600# gnd! 42.2fF
C1354 diff_107400_118080# gnd! 106.2fF
C1355 diff_99960_121680# gnd! 312.8fF
C1356 diff_103320_126720# gnd! 47.3fF
C1357 diff_104880_84600# gnd! 1606.5fF
C1358 diff_229920_128400# gnd! 131.7fF
C1359 diff_225960_120240# gnd! 117.6fF
C1360 diff_221760_128400# gnd! 103.0fF
C1361 diff_217680_120240# gnd! 122.4fF
C1362 diff_213600_128400# gnd! 108.7fF
C1363 diff_209520_120240# gnd! 120.2fF
C1364 diff_205440_128400# gnd! 105.2fF
C1365 diff_201360_120240# gnd! 122.4fF
C1366 diff_197280_128400# gnd! 108.7fF
C1367 diff_193200_120240# gnd! 120.2fF
C1368 diff_189120_128400# gnd! 105.2fF
C1369 diff_185160_120240# gnd! 122.4fF
C1370 diff_180960_128400# gnd! 109.0fF
C1371 diff_177000_120240# gnd! 120.2fF
C1372 diff_172800_128400# gnd! 105.4fF
C1373 diff_168720_120240# gnd! 118.5fF
C1374 diff_164640_128400# gnd! 104.8fF
C1375 diff_160560_120240# gnd! 116.2fF
C1376 diff_156480_128400# gnd! 101.1fF
C1377 diff_152400_120240# gnd! 118.5fF
C1378 diff_148320_128400# gnd! 104.1fF
C1379 diff_144240_120240# gnd! 116.2fF
C1380 diff_140160_128400# gnd! 101.1fF
C1381 diff_135960_120120# gnd! 126.8fF
C1382 diff_132000_128400# gnd! 111.6fF
C1383 diff_127800_120240# gnd! 124.1fF
C1384 diff_123840_128400# gnd! 107.2fF
C1385 diff_119760_120240# gnd! 122.4fF
C1386 diff_115680_128400# gnd! 109.0fF
C1387 diff_111600_120120# gnd! 120.5fF
C1388 diff_107520_128400# gnd! 105.8fF
C1389 diff_103680_120240# gnd! 119.6fF
C1390 diff_112440_115320# gnd! 787.8fF
C1391 diff_26040_78600# gnd! 665.5fF
C1392 cl gnd! 1717.2fF
C1393 diff_99720_123600# gnd! 98.6fF
C1394 diff_82080_129960# gnd! 206.4fF
C1395 diff_93600_128280# gnd! 24.3fF ;**FLOATING
C1396 diff_66600_129960# gnd! 203.3fF
C1397 diff_80160_117000# gnd! 309.1fF
C1398 diff_229320_128160# gnd! 42.9fF
C1399 diff_227280_132120# gnd! 43.5fF
C1400 diff_225240_126240# gnd! 54.6fF
C1401 diff_223200_132120# gnd! 54.5fF
C1402 diff_221160_128160# gnd! 42.9fF
C1403 diff_219120_132120# gnd! 43.5fF
C1404 diff_217080_126240# gnd! 54.6fF
C1405 diff_215040_132120# gnd! 54.5fF
C1406 diff_213000_128160# gnd! 42.9fF
C1407 diff_210960_132120# gnd! 43.5fF
C1408 diff_208920_126240# gnd! 54.6fF
C1409 diff_206880_132120# gnd! 54.5fF
C1410 diff_204840_128160# gnd! 42.9fF
C1411 diff_202800_132120# gnd! 43.5fF
C1412 diff_200760_126240# gnd! 54.6fF
C1413 diff_198720_132120# gnd! 54.5fF
C1414 diff_196680_128160# gnd! 42.9fF
C1415 diff_194640_132120# gnd! 43.5fF
C1416 diff_192600_126240# gnd! 54.6fF
C1417 diff_190560_132120# gnd! 54.5fF
C1418 diff_188520_128160# gnd! 42.9fF
C1419 diff_186480_132120# gnd! 43.5fF
C1420 diff_184440_126240# gnd! 54.6fF
C1421 diff_182400_132120# gnd! 54.5fF
C1422 diff_180360_128160# gnd! 42.9fF
C1423 diff_178320_132120# gnd! 43.5fF
C1424 diff_176280_126240# gnd! 54.6fF
C1425 diff_174240_132120# gnd! 54.5fF
C1426 diff_172200_128160# gnd! 42.9fF
C1427 diff_170160_132120# gnd! 43.5fF
C1428 diff_168120_126240# gnd! 54.6fF
C1429 diff_166080_132120# gnd! 54.5fF
C1430 diff_164040_128160# gnd! 42.9fF
C1431 diff_162000_132120# gnd! 43.5fF
C1432 diff_159960_126240# gnd! 54.6fF
C1433 diff_157920_132120# gnd! 54.5fF
C1434 diff_155880_128160# gnd! 42.9fF
C1435 diff_153840_132120# gnd! 43.5fF
C1436 diff_151800_126240# gnd! 54.6fF
C1437 diff_149760_132120# gnd! 54.5fF
C1438 diff_147720_128160# gnd! 42.9fF
C1439 diff_145680_132120# gnd! 43.5fF
C1440 diff_143640_126240# gnd! 54.6fF
C1441 diff_141600_132120# gnd! 54.5fF
C1442 diff_139560_128160# gnd! 42.9fF
C1443 diff_137520_132120# gnd! 43.5fF
C1444 diff_135480_126240# gnd! 54.6fF
C1445 diff_133440_132120# gnd! 54.5fF
C1446 diff_131400_128160# gnd! 42.9fF
C1447 diff_129360_132120# gnd! 43.5fF
C1448 diff_127320_126240# gnd! 54.6fF
C1449 diff_125280_132120# gnd! 54.5fF
C1450 diff_123240_128160# gnd! 42.9fF
C1451 diff_121200_132120# gnd! 43.5fF
C1452 diff_119160_126240# gnd! 54.6fF
C1453 diff_117120_132120# gnd! 54.5fF
C1454 diff_115080_128160# gnd! 42.9fF
C1455 diff_113040_132120# gnd! 43.5fF
C1456 diff_111000_126240# gnd! 54.6fF
C1457 diff_108960_132120# gnd! 54.5fF
C1458 diff_106920_128160# gnd! 41.8fF
C1459 diff_104880_132240# gnd! 42.6fF
C1460 diff_102480_126360# gnd! 56.9fF
C1461 diff_79920_127680# gnd! 305.3fF
C1462 diff_50880_129960# gnd! 206.6fF
C1463 diff_64680_117000# gnd! 318.7fF
C1464 diff_64440_127680# gnd! 304.3fF
C1465 diff_35520_129960# gnd! 207.4fF
C1466 diff_49200_117000# gnd! 308.5fF
C1467 diff_48840_127680# gnd! 297.6fF
C1468 diff_33600_117000# gnd! 309.9fF
C1469 diff_33360_127800# gnd! 303.1fF
C1470 diff_28080_131640# gnd! 278.2fF
C1471 diff_100800_132000# gnd! 50.4fF
C1472 diff_100440_134640# gnd! 613.8fF
C1473 diff_229320_135240# gnd! 26.2fF
C1474 diff_227280_135240# gnd! 26.2fF
C1475 diff_225240_135240# gnd! 26.2fF
C1476 diff_223200_135240# gnd! 26.2fF
C1477 diff_221160_135240# gnd! 26.2fF
C1478 diff_219120_135240# gnd! 26.2fF
C1479 diff_217080_135240# gnd! 26.2fF
C1480 diff_215040_135240# gnd! 26.2fF
C1481 diff_213000_135240# gnd! 26.2fF
C1482 diff_210960_135240# gnd! 26.2fF
C1483 diff_208920_135240# gnd! 26.2fF
C1484 diff_206880_135240# gnd! 26.2fF
C1485 diff_204840_135240# gnd! 26.2fF
C1486 diff_202800_135240# gnd! 26.2fF
C1487 diff_200760_135240# gnd! 26.2fF
C1488 diff_198720_135240# gnd! 26.2fF
C1489 diff_196680_135240# gnd! 26.2fF
C1490 diff_194640_135240# gnd! 26.2fF
C1491 diff_192600_135240# gnd! 26.2fF
C1492 diff_190560_135240# gnd! 26.2fF
C1493 diff_188520_135240# gnd! 26.2fF
C1494 diff_186480_135240# gnd! 26.2fF
C1495 diff_184440_135240# gnd! 26.2fF
C1496 diff_182400_135240# gnd! 26.2fF
C1497 diff_180360_135240# gnd! 26.2fF
C1498 diff_178320_135240# gnd! 26.2fF
C1499 diff_176280_135240# gnd! 26.2fF
C1500 diff_174240_135240# gnd! 26.2fF
C1501 diff_172200_135240# gnd! 26.2fF
C1502 diff_170160_135240# gnd! 26.2fF
C1503 diff_168120_135240# gnd! 26.2fF
C1504 diff_166080_135240# gnd! 26.2fF
C1505 diff_164040_135240# gnd! 26.2fF
C1506 diff_162000_135240# gnd! 26.2fF
C1507 diff_159960_135240# gnd! 26.2fF
C1508 diff_157920_135240# gnd! 26.2fF
C1509 diff_155880_135240# gnd! 26.2fF
C1510 diff_153840_135240# gnd! 26.2fF
C1511 diff_151800_135240# gnd! 26.2fF
C1512 diff_149760_135240# gnd! 26.2fF
C1513 diff_147720_135240# gnd! 26.2fF
C1514 diff_145680_135240# gnd! 26.2fF
C1515 diff_143640_135240# gnd! 26.2fF
C1516 diff_141600_135240# gnd! 26.2fF
C1517 diff_139560_135240# gnd! 26.2fF
C1518 diff_137520_135240# gnd! 26.2fF
C1519 diff_135480_135240# gnd! 26.2fF
C1520 diff_133440_135240# gnd! 26.2fF
C1521 diff_131400_135240# gnd! 26.2fF
C1522 diff_129360_135240# gnd! 26.2fF
C1523 diff_127320_135240# gnd! 26.2fF
C1524 diff_125280_135240# gnd! 26.2fF
C1525 diff_123240_135240# gnd! 26.2fF
C1526 diff_121200_135240# gnd! 26.2fF
C1527 diff_119160_135240# gnd! 26.2fF
C1528 diff_117120_135240# gnd! 26.2fF
C1529 diff_115080_135240# gnd! 26.2fF
C1530 diff_113040_135240# gnd! 26.2fF
C1531 diff_111000_135240# gnd! 26.2fF
C1532 diff_108960_135240# gnd! 26.2fF
C1533 diff_106920_135240# gnd! 26.2fF
C1534 diff_104880_135240# gnd! 26.2fF
C1535 diff_102840_135240# gnd! 26.2fF
C1536 diff_79920_134640# gnd! 14.2fF
C1537 diff_64440_134640# gnd! 14.2fF
C1538 diff_48840_134640# gnd! 14.2fF
C1539 diff_33360_134640# gnd! 14.2fF
C1540 diff_15480_82200# gnd! 792.9fF
C1541 diff_100800_135240# gnd! 26.2fF
C1542 diff_100440_136920# gnd! 644.8fF
C1543 diff_229320_137520# gnd! 24.7fF
C1544 diff_227280_137520# gnd! 24.7fF
C1545 diff_225240_137520# gnd! 24.7fF
C1546 diff_223200_137520# gnd! 24.7fF
C1547 diff_221160_137520# gnd! 24.7fF
C1548 diff_219120_137520# gnd! 24.7fF
C1549 diff_217080_137520# gnd! 24.7fF
C1550 diff_215040_137520# gnd! 24.7fF
C1551 diff_213000_137520# gnd! 24.7fF
C1552 diff_210960_137520# gnd! 24.7fF
C1553 diff_208920_137520# gnd! 24.7fF
C1554 diff_206880_137520# gnd! 24.7fF
C1555 diff_204840_137520# gnd! 24.7fF
C1556 diff_202800_137520# gnd! 24.7fF
C1557 diff_200760_137520# gnd! 24.7fF
C1558 diff_198720_137520# gnd! 24.7fF
C1559 diff_196680_137520# gnd! 24.7fF
C1560 diff_194640_137520# gnd! 24.7fF
C1561 diff_192600_137520# gnd! 24.7fF
C1562 diff_190560_137520# gnd! 24.7fF
C1563 diff_188520_137520# gnd! 24.7fF
C1564 diff_186480_137520# gnd! 24.7fF
C1565 diff_184440_137520# gnd! 24.7fF
C1566 diff_182400_137520# gnd! 24.7fF
C1567 diff_180360_137520# gnd! 24.7fF
C1568 diff_178320_137520# gnd! 24.7fF
C1569 diff_176280_137520# gnd! 24.7fF
C1570 diff_174240_137520# gnd! 24.7fF
C1571 diff_172200_137520# gnd! 24.7fF
C1572 diff_170160_137520# gnd! 24.7fF
C1573 diff_168120_137520# gnd! 24.7fF
C1574 diff_166080_137520# gnd! 24.7fF
C1575 diff_164040_137520# gnd! 24.7fF
C1576 diff_162000_137520# gnd! 24.7fF
C1577 diff_159960_137520# gnd! 24.7fF
C1578 diff_157920_137520# gnd! 24.7fF
C1579 diff_155880_137520# gnd! 24.7fF
C1580 diff_153840_137520# gnd! 24.7fF
C1581 diff_151800_137520# gnd! 24.7fF
C1582 diff_149760_137520# gnd! 24.7fF
C1583 diff_147720_137520# gnd! 24.7fF
C1584 diff_145680_137520# gnd! 24.7fF
C1585 diff_143640_137520# gnd! 24.7fF
C1586 diff_141600_137520# gnd! 24.7fF
C1587 diff_139560_137520# gnd! 24.7fF
C1588 diff_137520_137520# gnd! 24.7fF
C1589 diff_135480_137520# gnd! 24.7fF
C1590 diff_133440_137520# gnd! 24.7fF
C1591 diff_131400_137520# gnd! 24.7fF
C1592 diff_129360_137520# gnd! 24.7fF
C1593 diff_127320_137520# gnd! 24.7fF
C1594 diff_125280_137520# gnd! 24.7fF
C1595 diff_123240_137520# gnd! 24.7fF
C1596 diff_121200_137520# gnd! 24.7fF
C1597 diff_119160_137520# gnd! 24.7fF
C1598 diff_117120_137520# gnd! 24.7fF
C1599 diff_115080_137520# gnd! 24.7fF
C1600 diff_113040_137520# gnd! 24.7fF
C1601 diff_111000_137520# gnd! 24.7fF
C1602 diff_108960_137520# gnd! 24.7fF
C1603 diff_106920_137520# gnd! 24.7fF
C1604 diff_104880_137520# gnd! 24.7fF
C1605 diff_102840_137520# gnd! 24.7fF
C1606 diff_100800_137520# gnd! 24.7fF
C1607 diff_100440_139080# gnd! 649.5fF
C1608 diff_236760_140760# gnd! 500.4fF
C1609 diff_229320_139680# gnd! 26.2fF
C1610 diff_227280_139680# gnd! 26.2fF
C1611 diff_225240_139680# gnd! 26.2fF
C1612 diff_223200_139680# gnd! 26.2fF
C1613 diff_221160_139680# gnd! 26.2fF
C1614 diff_219120_139680# gnd! 26.2fF
C1615 diff_217080_139680# gnd! 26.2fF
C1616 diff_215040_139680# gnd! 26.2fF
C1617 diff_213000_139680# gnd! 26.2fF
C1618 diff_210960_139680# gnd! 26.2fF
C1619 diff_208920_139680# gnd! 26.2fF
C1620 diff_206880_139680# gnd! 26.2fF
C1621 diff_204840_139680# gnd! 26.2fF
C1622 diff_202800_139680# gnd! 26.2fF
C1623 diff_200760_139680# gnd! 26.2fF
C1624 diff_198720_139680# gnd! 26.2fF
C1625 diff_196680_139680# gnd! 26.2fF
C1626 diff_194640_139680# gnd! 26.2fF
C1627 diff_192600_139680# gnd! 26.2fF
C1628 diff_190560_139680# gnd! 26.2fF
C1629 diff_188520_139680# gnd! 26.2fF
C1630 diff_186480_139680# gnd! 26.2fF
C1631 diff_184440_139680# gnd! 26.2fF
C1632 diff_182400_139680# gnd! 26.2fF
C1633 diff_180360_139680# gnd! 26.2fF
C1634 diff_178320_139680# gnd! 26.2fF
C1635 diff_176280_139680# gnd! 26.2fF
C1636 diff_174240_139680# gnd! 26.2fF
C1637 diff_172200_139680# gnd! 26.2fF
C1638 diff_170160_139680# gnd! 26.2fF
C1639 diff_168120_139680# gnd! 26.2fF
C1640 diff_166080_139680# gnd! 26.2fF
C1641 diff_164040_139680# gnd! 26.2fF
C1642 diff_162000_139680# gnd! 26.2fF
C1643 diff_159960_139680# gnd! 26.2fF
C1644 diff_157920_139680# gnd! 26.2fF
C1645 diff_155880_139680# gnd! 26.2fF
C1646 diff_153840_139680# gnd! 26.2fF
C1647 diff_151800_139680# gnd! 26.2fF
C1648 diff_149760_139680# gnd! 26.2fF
C1649 diff_147720_139680# gnd! 26.2fF
C1650 diff_145680_139680# gnd! 26.2fF
C1651 diff_143640_139680# gnd! 26.2fF
C1652 diff_141600_139680# gnd! 26.2fF
C1653 diff_139560_139680# gnd! 26.2fF
C1654 diff_137520_139680# gnd! 26.2fF
C1655 diff_135480_139680# gnd! 26.2fF
C1656 diff_133440_139680# gnd! 26.2fF
C1657 diff_131400_139680# gnd! 26.2fF
C1658 diff_129360_139680# gnd! 26.2fF
C1659 diff_127320_139680# gnd! 26.2fF
C1660 diff_125280_139680# gnd! 26.2fF
C1661 diff_123240_139680# gnd! 26.2fF
C1662 diff_121200_139680# gnd! 26.2fF
C1663 diff_119160_139680# gnd! 26.2fF
C1664 diff_117120_139680# gnd! 26.2fF
C1665 diff_115080_139680# gnd! 26.2fF
C1666 diff_113040_139680# gnd! 26.2fF
C1667 diff_111000_139680# gnd! 26.2fF
C1668 diff_108960_139680# gnd! 26.2fF
C1669 diff_106920_139680# gnd! 26.2fF
C1670 diff_104880_139680# gnd! 26.2fF
C1671 diff_102840_139680# gnd! 26.2fF
C1672 diff_100800_139680# gnd! 26.2fF
C1673 diff_100440_141360# gnd! 609.5fF
C1674 diff_229320_141960# gnd! 24.7fF
C1675 diff_227280_141960# gnd! 24.7fF
C1676 diff_225240_141960# gnd! 24.7fF
C1677 diff_223200_141960# gnd! 24.7fF
C1678 diff_221160_141960# gnd! 24.7fF
C1679 diff_219120_141960# gnd! 24.7fF
C1680 diff_217080_141960# gnd! 24.7fF
C1681 diff_215040_141960# gnd! 24.7fF
C1682 diff_213000_141960# gnd! 24.7fF
C1683 diff_210960_141960# gnd! 24.7fF
C1684 diff_208920_141960# gnd! 24.7fF
C1685 diff_206880_141960# gnd! 24.7fF
C1686 diff_204840_141960# gnd! 24.7fF
C1687 diff_202800_141960# gnd! 24.7fF
C1688 diff_200760_141960# gnd! 24.7fF
C1689 diff_198720_141960# gnd! 24.7fF
C1690 diff_196680_141960# gnd! 24.7fF
C1691 diff_194640_141960# gnd! 24.7fF
C1692 diff_192600_141960# gnd! 24.7fF
C1693 diff_190560_141960# gnd! 24.7fF
C1694 diff_188520_141960# gnd! 24.7fF
C1695 diff_186480_141960# gnd! 24.7fF
C1696 diff_184440_141960# gnd! 24.7fF
C1697 diff_182400_141960# gnd! 24.7fF
C1698 diff_180360_141960# gnd! 24.7fF
C1699 diff_178320_141960# gnd! 24.7fF
C1700 diff_176280_141960# gnd! 24.7fF
C1701 diff_174240_141960# gnd! 24.7fF
C1702 diff_172200_141960# gnd! 24.7fF
C1703 diff_170160_141960# gnd! 24.7fF
C1704 diff_168120_141960# gnd! 24.7fF
C1705 diff_166080_141960# gnd! 24.7fF
C1706 diff_164040_141960# gnd! 24.7fF
C1707 diff_162000_141960# gnd! 24.7fF
C1708 diff_159960_141960# gnd! 24.7fF
C1709 diff_157920_141960# gnd! 24.7fF
C1710 diff_155880_141960# gnd! 24.7fF
C1711 diff_153840_141960# gnd! 24.7fF
C1712 diff_151800_141960# gnd! 24.7fF
C1713 diff_149760_141960# gnd! 24.7fF
C1714 diff_147720_141960# gnd! 24.7fF
C1715 diff_145680_141960# gnd! 24.7fF
C1716 diff_143640_141960# gnd! 24.7fF
C1717 diff_141600_141960# gnd! 24.7fF
C1718 diff_139560_141960# gnd! 24.7fF
C1719 diff_137520_141960# gnd! 24.7fF
C1720 diff_135480_141960# gnd! 24.7fF
C1721 diff_133440_141960# gnd! 24.7fF
C1722 diff_131400_141960# gnd! 24.7fF
C1723 diff_129360_141960# gnd! 24.7fF
C1724 diff_127320_141960# gnd! 24.7fF
C1725 diff_125280_141960# gnd! 24.7fF
C1726 diff_123240_141960# gnd! 24.7fF
C1727 diff_121200_141960# gnd! 24.7fF
C1728 diff_119160_141960# gnd! 24.7fF
C1729 diff_117120_141960# gnd! 24.7fF
C1730 diff_115080_141960# gnd! 24.7fF
C1731 diff_113040_141960# gnd! 24.7fF
C1732 diff_111000_141960# gnd! 24.7fF
C1733 diff_108960_141960# gnd! 24.7fF
C1734 diff_106920_141960# gnd! 24.7fF
C1735 diff_104880_141960# gnd! 24.7fF
C1736 diff_102840_141960# gnd! 24.7fF
C1737 diff_100800_141960# gnd! 24.7fF
C1738 diff_100440_143520# gnd! 614.5fF
C1739 diff_229320_144120# gnd! 26.2fF
C1740 diff_227280_144120# gnd! 26.2fF
C1741 diff_225240_144120# gnd! 26.2fF
C1742 diff_223200_144120# gnd! 26.2fF
C1743 diff_221160_144120# gnd! 26.2fF
C1744 diff_219120_144120# gnd! 26.2fF
C1745 diff_217080_144120# gnd! 26.2fF
C1746 diff_215040_144120# gnd! 26.2fF
C1747 diff_213000_144120# gnd! 26.2fF
C1748 diff_210960_144120# gnd! 26.2fF
C1749 diff_208920_144120# gnd! 26.2fF
C1750 diff_206880_144120# gnd! 26.2fF
C1751 diff_204840_144120# gnd! 26.2fF
C1752 diff_202800_144120# gnd! 26.2fF
C1753 diff_200760_144120# gnd! 26.2fF
C1754 diff_198720_144120# gnd! 26.2fF
C1755 diff_196680_144120# gnd! 26.2fF
C1756 diff_194640_144120# gnd! 26.2fF
C1757 diff_192600_144120# gnd! 26.2fF
C1758 diff_190560_144120# gnd! 26.2fF
C1759 diff_188520_144120# gnd! 26.2fF
C1760 diff_186480_144120# gnd! 26.2fF
C1761 diff_184440_144120# gnd! 26.2fF
C1762 diff_182400_144120# gnd! 26.2fF
C1763 diff_180360_144120# gnd! 26.2fF
C1764 diff_178320_144120# gnd! 26.2fF
C1765 diff_176280_144120# gnd! 26.2fF
C1766 diff_174240_144120# gnd! 26.2fF
C1767 diff_172200_144120# gnd! 26.2fF
C1768 diff_170160_144120# gnd! 26.2fF
C1769 diff_168120_144120# gnd! 26.2fF
C1770 diff_166080_144120# gnd! 26.2fF
C1771 diff_164040_144120# gnd! 26.2fF
C1772 diff_162000_144120# gnd! 26.2fF
C1773 diff_159960_144120# gnd! 26.2fF
C1774 diff_157920_144120# gnd! 26.2fF
C1775 diff_155880_144120# gnd! 26.2fF
C1776 diff_153840_144120# gnd! 26.2fF
C1777 diff_151800_144120# gnd! 26.2fF
C1778 diff_149760_144120# gnd! 26.2fF
C1779 diff_147720_144120# gnd! 26.2fF
C1780 diff_145680_144120# gnd! 26.2fF
C1781 diff_143640_144120# gnd! 26.2fF
C1782 diff_141600_144120# gnd! 26.2fF
C1783 diff_139560_144120# gnd! 26.2fF
C1784 diff_137520_144120# gnd! 26.2fF
C1785 diff_135480_144120# gnd! 26.2fF
C1786 diff_133440_144120# gnd! 26.2fF
C1787 diff_131400_144120# gnd! 26.2fF
C1788 diff_129360_144120# gnd! 26.2fF
C1789 diff_127320_144120# gnd! 26.2fF
C1790 diff_125280_144120# gnd! 26.2fF
C1791 diff_123240_144120# gnd! 26.2fF
C1792 diff_121200_144120# gnd! 26.2fF
C1793 diff_119160_144120# gnd! 26.2fF
C1794 diff_117120_144120# gnd! 26.2fF
C1795 diff_115080_144120# gnd! 26.2fF
C1796 diff_113040_144120# gnd! 26.2fF
C1797 diff_111000_144120# gnd! 26.2fF
C1798 diff_108960_144120# gnd! 26.2fF
C1799 diff_106920_144120# gnd! 26.2fF
C1800 diff_104880_144120# gnd! 26.2fF
C1801 diff_102840_144120# gnd! 26.2fF
C1802 diff_100800_144120# gnd! 26.2fF
C1803 diff_100440_145800# gnd! 646.1fF
C1804 diff_229320_146400# gnd! 24.7fF
C1805 diff_227280_146400# gnd! 24.7fF
C1806 diff_225240_146400# gnd! 24.7fF
C1807 diff_223200_146400# gnd! 24.7fF
C1808 diff_221160_146400# gnd! 24.7fF
C1809 diff_219120_146400# gnd! 24.7fF
C1810 diff_217080_146400# gnd! 24.7fF
C1811 diff_215040_146400# gnd! 24.7fF
C1812 diff_213000_146400# gnd! 24.7fF
C1813 diff_210960_146400# gnd! 24.7fF
C1814 diff_208920_146400# gnd! 24.7fF
C1815 diff_206880_146400# gnd! 24.7fF
C1816 diff_204840_146400# gnd! 24.7fF
C1817 diff_202800_146400# gnd! 24.7fF
C1818 diff_200760_146400# gnd! 24.7fF
C1819 diff_198720_146400# gnd! 24.7fF
C1820 diff_196680_146400# gnd! 24.7fF
C1821 diff_194640_146400# gnd! 24.7fF
C1822 diff_192600_146400# gnd! 24.7fF
C1823 diff_190560_146400# gnd! 24.7fF
C1824 diff_188520_146400# gnd! 24.7fF
C1825 diff_186480_146400# gnd! 24.7fF
C1826 diff_184440_146400# gnd! 24.7fF
C1827 diff_182400_146400# gnd! 24.7fF
C1828 diff_180360_146400# gnd! 24.7fF
C1829 diff_178320_146400# gnd! 24.7fF
C1830 diff_176280_146400# gnd! 24.7fF
C1831 diff_174240_146400# gnd! 24.7fF
C1832 diff_172200_146400# gnd! 24.7fF
C1833 diff_170160_146400# gnd! 24.7fF
C1834 diff_168120_146400# gnd! 24.7fF
C1835 diff_166080_146400# gnd! 24.7fF
C1836 diff_164040_146400# gnd! 24.7fF
C1837 diff_162000_146400# gnd! 24.7fF
C1838 diff_159960_146400# gnd! 24.7fF
C1839 diff_157920_146400# gnd! 24.7fF
C1840 diff_155880_146400# gnd! 24.7fF
C1841 diff_153840_146400# gnd! 24.7fF
C1842 diff_151800_146400# gnd! 24.7fF
C1843 diff_149760_146400# gnd! 24.7fF
C1844 diff_147720_146400# gnd! 24.7fF
C1845 diff_145680_146400# gnd! 24.7fF
C1846 diff_143640_146400# gnd! 24.7fF
C1847 diff_141600_146400# gnd! 24.7fF
C1848 diff_139560_146400# gnd! 24.7fF
C1849 diff_137520_146400# gnd! 24.7fF
C1850 diff_135480_146400# gnd! 24.7fF
C1851 diff_133440_146400# gnd! 24.7fF
C1852 diff_131400_146400# gnd! 24.7fF
C1853 diff_129360_146400# gnd! 24.7fF
C1854 diff_127320_146400# gnd! 24.7fF
C1855 diff_125280_146400# gnd! 24.7fF
C1856 diff_123240_146400# gnd! 24.7fF
C1857 diff_121200_146400# gnd! 24.7fF
C1858 diff_119160_146400# gnd! 24.7fF
C1859 diff_117120_146400# gnd! 24.7fF
C1860 diff_115080_146400# gnd! 24.7fF
C1861 diff_113040_146400# gnd! 24.7fF
C1862 diff_111000_146400# gnd! 24.7fF
C1863 diff_108960_146400# gnd! 24.7fF
C1864 diff_106920_146400# gnd! 24.7fF
C1865 diff_104880_146400# gnd! 24.7fF
C1866 diff_102840_146400# gnd! 24.7fF
C1867 diff_100800_146400# gnd! 24.7fF
C1868 diff_100440_147960# gnd! 650.3fF
C1869 diff_245160_97920# gnd! 624.8fF
C1870 diff_246960_91200# gnd! 639.2fF
C1871 diff_259200_153240# gnd! 78.7fF
C1872 diff_281280_100320# gnd! 664.5fF
C1873 diff_276720_158280# gnd! 54.0fF
C1874 diff_271080_135600# gnd! 535.5fF
C1875 diff_282840_127320# gnd! 309.1fF
C1876 diff_282840_108600# gnd! 573.8fF
C1877 diff_268200_169080# gnd! 53.5fF
C1878 diff_264960_151920# gnd! 381.4fF
C1879 diff_274320_170280# gnd! 55.8fF
C1880 diff_266400_142200# gnd! 332.6fF
C1881 diff_274320_171480# gnd! 49.2fF
C1882 diff_236760_149400# gnd! 529.2fF
C1883 diff_229320_148560# gnd! 26.2fF
C1884 diff_227280_148560# gnd! 26.2fF
C1885 diff_225240_148560# gnd! 26.2fF
C1886 diff_223200_148560# gnd! 26.2fF
C1887 diff_221160_148560# gnd! 26.2fF
C1888 diff_219120_148560# gnd! 26.2fF
C1889 diff_217080_148560# gnd! 26.2fF
C1890 diff_215040_148560# gnd! 26.2fF
C1891 diff_213000_148560# gnd! 26.2fF
C1892 diff_210960_148560# gnd! 26.2fF
C1893 diff_208920_148560# gnd! 26.2fF
C1894 diff_206880_148560# gnd! 26.2fF
C1895 diff_204840_148560# gnd! 26.2fF
C1896 diff_202800_148560# gnd! 26.2fF
C1897 diff_200760_148560# gnd! 26.2fF
C1898 diff_198720_148560# gnd! 26.2fF
C1899 diff_196680_148560# gnd! 26.2fF
C1900 diff_194640_148560# gnd! 26.2fF
C1901 diff_192600_148560# gnd! 26.2fF
C1902 diff_190560_148560# gnd! 26.2fF
C1903 diff_188520_148560# gnd! 26.2fF
C1904 diff_186480_148560# gnd! 26.2fF
C1905 diff_184440_148560# gnd! 26.2fF
C1906 diff_182400_148560# gnd! 26.2fF
C1907 diff_180360_148560# gnd! 26.2fF
C1908 diff_178320_148560# gnd! 26.2fF
C1909 diff_176280_148560# gnd! 26.2fF
C1910 diff_174240_148560# gnd! 26.2fF
C1911 diff_172200_148560# gnd! 26.2fF
C1912 diff_170160_148560# gnd! 26.2fF
C1913 diff_168120_148560# gnd! 26.2fF
C1914 diff_166080_148560# gnd! 26.2fF
C1915 diff_164040_148560# gnd! 26.2fF
C1916 diff_162000_148560# gnd! 26.2fF
C1917 diff_159960_148560# gnd! 26.2fF
C1918 diff_157920_148560# gnd! 26.2fF
C1919 diff_155880_148560# gnd! 26.2fF
C1920 diff_153840_148560# gnd! 26.2fF
C1921 diff_151800_148560# gnd! 26.2fF
C1922 diff_149760_148560# gnd! 26.2fF
C1923 diff_147720_148560# gnd! 26.2fF
C1924 diff_145680_148560# gnd! 26.2fF
C1925 diff_143640_148560# gnd! 26.2fF
C1926 diff_141600_148560# gnd! 26.2fF
C1927 diff_139560_148560# gnd! 26.2fF
C1928 diff_137520_148560# gnd! 26.2fF
C1929 diff_135480_148560# gnd! 26.2fF
C1930 diff_133440_148560# gnd! 26.2fF
C1931 diff_131400_148560# gnd! 26.2fF
C1932 diff_129360_148560# gnd! 26.2fF
C1933 diff_127320_148560# gnd! 26.2fF
C1934 diff_125280_148560# gnd! 26.2fF
C1935 diff_123240_148560# gnd! 26.2fF
C1936 diff_121200_148560# gnd! 26.2fF
C1937 diff_119160_148560# gnd! 26.2fF
C1938 diff_117120_148560# gnd! 26.2fF
C1939 diff_115080_148560# gnd! 26.2fF
C1940 diff_113040_148560# gnd! 26.2fF
C1941 diff_111000_148560# gnd! 26.2fF
C1942 diff_108960_148560# gnd! 26.2fF
C1943 diff_106920_148560# gnd! 26.2fF
C1944 diff_104880_148560# gnd! 26.2fF
C1945 diff_102840_148560# gnd! 26.2fF
C1946 diff_87360_144840# gnd! 235.4fF
C1947 diff_100800_148560# gnd! 26.2fF
C1948 diff_71880_144840# gnd! 309.7fF
C1949 diff_100440_150240# gnd! 606.7fF
C1950 diff_229320_150840# gnd! 24.7fF
C1951 diff_227280_150840# gnd! 24.7fF
C1952 diff_225240_150840# gnd! 24.7fF
C1953 diff_223200_150840# gnd! 24.7fF
C1954 diff_221160_150840# gnd! 24.7fF
C1955 diff_219120_150840# gnd! 24.7fF
C1956 diff_217080_150840# gnd! 24.7fF
C1957 diff_215040_150840# gnd! 24.7fF
C1958 diff_213000_150840# gnd! 24.7fF
C1959 diff_210960_150840# gnd! 24.7fF
C1960 diff_208920_150840# gnd! 24.7fF
C1961 diff_206880_150840# gnd! 24.7fF
C1962 diff_204840_150840# gnd! 24.7fF
C1963 diff_202800_150840# gnd! 24.7fF
C1964 diff_200760_150840# gnd! 24.7fF
C1965 diff_198720_150840# gnd! 24.7fF
C1966 diff_196680_150840# gnd! 24.7fF
C1967 diff_194640_150840# gnd! 24.7fF
C1968 diff_192600_150840# gnd! 24.7fF
C1969 diff_190560_150840# gnd! 24.7fF
C1970 diff_188520_150840# gnd! 24.7fF
C1971 diff_186480_150840# gnd! 24.7fF
C1972 diff_184440_150840# gnd! 24.7fF
C1973 diff_182400_150840# gnd! 24.7fF
C1974 diff_180360_150840# gnd! 24.7fF
C1975 diff_178320_150840# gnd! 24.7fF
C1976 diff_176280_150840# gnd! 24.7fF
C1977 diff_174240_150840# gnd! 24.7fF
C1978 diff_172200_150840# gnd! 24.7fF
C1979 diff_170160_150840# gnd! 24.7fF
C1980 diff_168120_150840# gnd! 24.7fF
C1981 diff_166080_150840# gnd! 24.7fF
C1982 diff_164040_150840# gnd! 24.7fF
C1983 diff_162000_150840# gnd! 24.7fF
C1984 diff_159960_150840# gnd! 24.7fF
C1985 diff_157920_150840# gnd! 24.7fF
C1986 diff_155880_150840# gnd! 24.7fF
C1987 diff_153840_150840# gnd! 24.7fF
C1988 diff_151800_150840# gnd! 24.7fF
C1989 diff_149760_150840# gnd! 24.7fF
C1990 diff_147720_150840# gnd! 24.7fF
C1991 diff_145680_150840# gnd! 24.7fF
C1992 diff_143640_150840# gnd! 24.7fF
C1993 diff_141600_150840# gnd! 24.7fF
C1994 diff_139560_150840# gnd! 24.7fF
C1995 diff_137520_150840# gnd! 24.7fF
C1996 diff_135480_150840# gnd! 24.7fF
C1997 diff_133440_150840# gnd! 24.7fF
C1998 diff_131400_150840# gnd! 24.7fF
C1999 diff_129360_150840# gnd! 24.7fF
C2000 diff_127320_150840# gnd! 24.7fF
C2001 diff_125280_150840# gnd! 24.7fF
C2002 diff_123240_150840# gnd! 24.7fF
C2003 diff_121200_150840# gnd! 24.7fF
C2004 diff_119160_150840# gnd! 24.7fF
C2005 diff_117120_150840# gnd! 24.7fF
C2006 diff_115080_150840# gnd! 24.7fF
C2007 diff_113040_150840# gnd! 24.7fF
C2008 diff_111000_150840# gnd! 24.7fF
C2009 diff_108960_150840# gnd! 24.7fF
C2010 diff_106920_150840# gnd! 24.7fF
C2011 diff_104880_150840# gnd! 24.7fF
C2012 diff_102840_150840# gnd! 24.7fF
C2013 diff_100800_150840# gnd! 24.7fF
C2014 diff_100440_152400# gnd! 614.7fF
C2015 diff_229320_153000# gnd! 26.2fF
C2016 diff_227280_153000# gnd! 26.2fF
C2017 diff_225240_153000# gnd! 26.2fF
C2018 diff_223200_153000# gnd! 26.2fF
C2019 diff_221160_153000# gnd! 26.2fF
C2020 diff_219120_153000# gnd! 26.2fF
C2021 diff_217080_153000# gnd! 26.2fF
C2022 diff_215040_153000# gnd! 26.2fF
C2023 diff_213000_153000# gnd! 26.2fF
C2024 diff_210960_153000# gnd! 26.2fF
C2025 diff_208920_153000# gnd! 26.2fF
C2026 diff_206880_153000# gnd! 26.2fF
C2027 diff_204840_153000# gnd! 26.2fF
C2028 diff_202800_153000# gnd! 26.2fF
C2029 diff_200760_153000# gnd! 26.2fF
C2030 diff_198720_153000# gnd! 26.2fF
C2031 diff_196680_153000# gnd! 26.2fF
C2032 diff_194640_153000# gnd! 26.2fF
C2033 diff_192600_153000# gnd! 26.2fF
C2034 diff_190560_153000# gnd! 26.2fF
C2035 diff_188520_153000# gnd! 26.2fF
C2036 diff_186480_153000# gnd! 26.2fF
C2037 diff_184440_153000# gnd! 26.2fF
C2038 diff_182400_153000# gnd! 26.2fF
C2039 diff_180360_153000# gnd! 26.2fF
C2040 diff_178320_153000# gnd! 26.2fF
C2041 diff_176280_153000# gnd! 26.2fF
C2042 diff_174240_153000# gnd! 26.2fF
C2043 diff_172200_153000# gnd! 26.2fF
C2044 diff_170160_153000# gnd! 26.2fF
C2045 diff_168120_153000# gnd! 26.2fF
C2046 diff_166080_153000# gnd! 26.2fF
C2047 diff_164040_153000# gnd! 26.2fF
C2048 diff_162000_153000# gnd! 26.2fF
C2049 diff_159960_153000# gnd! 26.2fF
C2050 diff_157920_153000# gnd! 26.2fF
C2051 diff_155880_153000# gnd! 26.2fF
C2052 diff_153840_153000# gnd! 26.2fF
C2053 diff_151800_153000# gnd! 26.2fF
C2054 diff_149760_153000# gnd! 26.2fF
C2055 diff_147720_153000# gnd! 26.2fF
C2056 diff_145680_153000# gnd! 26.2fF
C2057 diff_143640_153000# gnd! 26.2fF
C2058 diff_141600_153000# gnd! 26.2fF
C2059 diff_139560_153000# gnd! 26.2fF
C2060 diff_137520_153000# gnd! 26.2fF
C2061 diff_135480_153000# gnd! 26.2fF
C2062 diff_133440_153000# gnd! 26.2fF
C2063 diff_131400_153000# gnd! 26.2fF
C2064 diff_129360_153000# gnd! 26.2fF
C2065 diff_127320_153000# gnd! 26.2fF
C2066 diff_125280_153000# gnd! 26.2fF
C2067 diff_123240_153000# gnd! 26.2fF
C2068 diff_121200_153000# gnd! 26.2fF
C2069 diff_119160_153000# gnd! 26.2fF
C2070 diff_117120_153000# gnd! 26.2fF
C2071 diff_115080_153000# gnd! 26.2fF
C2072 diff_113040_153000# gnd! 26.2fF
C2073 diff_111000_153000# gnd! 26.2fF
C2074 diff_108960_153000# gnd! 26.2fF
C2075 diff_106920_153000# gnd! 26.2fF
C2076 diff_104880_153000# gnd! 26.2fF
C2077 diff_102840_153000# gnd! 26.2fF
C2078 diff_100800_153000# gnd! 26.2fF
C2079 diff_100440_154680# gnd! 645.4fF
C2080 diff_229320_155280# gnd! 24.7fF
C2081 diff_227280_155280# gnd! 24.7fF
C2082 diff_225240_155280# gnd! 24.7fF
C2083 diff_223200_155280# gnd! 24.7fF
C2084 diff_221160_155280# gnd! 24.7fF
C2085 diff_219120_155280# gnd! 24.7fF
C2086 diff_217080_155280# gnd! 24.7fF
C2087 diff_215040_155280# gnd! 24.7fF
C2088 diff_213000_155280# gnd! 24.7fF
C2089 diff_210960_155280# gnd! 24.7fF
C2090 diff_208920_155280# gnd! 24.7fF
C2091 diff_206880_155280# gnd! 24.7fF
C2092 diff_204840_155280# gnd! 24.7fF
C2093 diff_202800_155280# gnd! 24.7fF
C2094 diff_200760_155280# gnd! 24.7fF
C2095 diff_198720_155280# gnd! 24.7fF
C2096 diff_196680_155280# gnd! 24.7fF
C2097 diff_194640_155280# gnd! 24.7fF
C2098 diff_192600_155280# gnd! 24.7fF
C2099 diff_190560_155280# gnd! 24.7fF
C2100 diff_188520_155280# gnd! 24.7fF
C2101 diff_186480_155280# gnd! 24.7fF
C2102 diff_184440_155280# gnd! 24.7fF
C2103 diff_182400_155280# gnd! 24.7fF
C2104 diff_180360_155280# gnd! 24.7fF
C2105 diff_178320_155280# gnd! 24.7fF
C2106 diff_176280_155280# gnd! 24.7fF
C2107 diff_174240_155280# gnd! 24.7fF
C2108 diff_172200_155280# gnd! 24.7fF
C2109 diff_170160_155280# gnd! 24.7fF
C2110 diff_168120_155280# gnd! 24.7fF
C2111 diff_166080_155280# gnd! 24.7fF
C2112 diff_164040_155280# gnd! 24.7fF
C2113 diff_162000_155280# gnd! 24.7fF
C2114 diff_159960_155280# gnd! 24.7fF
C2115 diff_157920_155280# gnd! 24.7fF
C2116 diff_155880_155280# gnd! 24.7fF
C2117 diff_153840_155280# gnd! 24.7fF
C2118 diff_151800_155280# gnd! 24.7fF
C2119 diff_149760_155280# gnd! 24.7fF
C2120 diff_147720_155280# gnd! 24.7fF
C2121 diff_145680_155280# gnd! 24.7fF
C2122 diff_143640_155280# gnd! 24.7fF
C2123 diff_141600_155280# gnd! 24.7fF
C2124 diff_139560_155280# gnd! 24.7fF
C2125 diff_137520_155280# gnd! 24.7fF
C2126 diff_135480_155280# gnd! 24.7fF
C2127 diff_133440_155280# gnd! 24.7fF
C2128 diff_131400_155280# gnd! 24.7fF
C2129 diff_129360_155280# gnd! 24.7fF
C2130 diff_127320_155280# gnd! 24.7fF
C2131 diff_125280_155280# gnd! 24.7fF
C2132 diff_123240_155280# gnd! 24.7fF
C2133 diff_121200_155280# gnd! 24.7fF
C2134 diff_119160_155280# gnd! 24.7fF
C2135 diff_117120_155280# gnd! 24.7fF
C2136 diff_115080_155280# gnd! 24.7fF
C2137 diff_113040_155280# gnd! 24.7fF
C2138 diff_111000_155280# gnd! 24.7fF
C2139 diff_108960_155280# gnd! 24.7fF
C2140 diff_106920_155280# gnd! 24.7fF
C2141 diff_104880_155280# gnd! 24.7fF
C2142 diff_102840_155280# gnd! 24.7fF
C2143 diff_100800_155280# gnd! 24.7fF
C2144 diff_56280_144840# gnd! 324.8fF
C2145 diff_40800_144840# gnd! 356.5fF
C2146 diff_100440_156840# gnd! 646.5fF
C2147 diff_236760_158520# gnd! 505.2fF
C2148 diff_229320_157440# gnd! 26.2fF
C2149 diff_227280_157440# gnd! 26.2fF
C2150 diff_225240_157440# gnd! 26.2fF
C2151 diff_223200_157440# gnd! 26.2fF
C2152 diff_221160_157440# gnd! 26.2fF
C2153 diff_219120_157440# gnd! 26.2fF
C2154 diff_217080_157440# gnd! 26.2fF
C2155 diff_215040_157440# gnd! 26.2fF
C2156 diff_213000_157440# gnd! 26.2fF
C2157 diff_210960_157440# gnd! 26.2fF
C2158 diff_208920_157440# gnd! 26.2fF
C2159 diff_206880_157440# gnd! 26.2fF
C2160 diff_204840_157440# gnd! 26.2fF
C2161 diff_202800_157440# gnd! 26.2fF
C2162 diff_200760_157440# gnd! 26.2fF
C2163 diff_198720_157440# gnd! 26.2fF
C2164 diff_196680_157440# gnd! 26.2fF
C2165 diff_194640_157440# gnd! 26.2fF
C2166 diff_192600_157440# gnd! 26.2fF
C2167 diff_190560_157440# gnd! 26.2fF
C2168 diff_188520_157440# gnd! 26.2fF
C2169 diff_186480_157440# gnd! 26.2fF
C2170 diff_184440_157440# gnd! 26.2fF
C2171 diff_182400_157440# gnd! 26.2fF
C2172 diff_180360_157440# gnd! 26.2fF
C2173 diff_178320_157440# gnd! 26.2fF
C2174 diff_176280_157440# gnd! 26.2fF
C2175 diff_174240_157440# gnd! 26.2fF
C2176 diff_172200_157440# gnd! 26.2fF
C2177 diff_170160_157440# gnd! 26.2fF
C2178 diff_168120_157440# gnd! 26.2fF
C2179 diff_166080_157440# gnd! 26.2fF
C2180 diff_164040_157440# gnd! 26.2fF
C2181 diff_162000_157440# gnd! 26.2fF
C2182 diff_159960_157440# gnd! 26.2fF
C2183 diff_157920_157440# gnd! 26.2fF
C2184 diff_155880_157440# gnd! 26.2fF
C2185 diff_153840_157440# gnd! 26.2fF
C2186 diff_151800_157440# gnd! 26.2fF
C2187 diff_149760_157440# gnd! 26.2fF
C2188 diff_147720_157440# gnd! 26.2fF
C2189 diff_145680_157440# gnd! 26.2fF
C2190 diff_143640_157440# gnd! 26.2fF
C2191 diff_141600_157440# gnd! 26.2fF
C2192 diff_139560_157440# gnd! 26.2fF
C2193 diff_137520_157440# gnd! 26.2fF
C2194 diff_135480_157440# gnd! 26.2fF
C2195 diff_133440_157440# gnd! 26.2fF
C2196 diff_131400_157440# gnd! 26.2fF
C2197 diff_129360_157440# gnd! 26.2fF
C2198 diff_127320_157440# gnd! 26.2fF
C2199 diff_125280_157440# gnd! 26.2fF
C2200 diff_123240_157440# gnd! 26.2fF
C2201 diff_121200_157440# gnd! 26.2fF
C2202 diff_119160_157440# gnd! 26.2fF
C2203 diff_117120_157440# gnd! 26.2fF
C2204 diff_115080_157440# gnd! 26.2fF
C2205 diff_113040_157440# gnd! 26.2fF
C2206 diff_111000_157440# gnd! 26.2fF
C2207 diff_108960_157440# gnd! 26.2fF
C2208 diff_106920_157440# gnd! 26.2fF
C2209 diff_104880_157440# gnd! 26.2fF
C2210 diff_102840_157440# gnd! 26.2fF
C2211 diff_100800_157440# gnd! 26.2fF
C2212 diff_100440_159120# gnd! 600.9fF
C2213 diff_229320_159720# gnd! 24.7fF
C2214 diff_227280_159720# gnd! 24.7fF
C2215 diff_225240_159720# gnd! 24.7fF
C2216 diff_223200_159720# gnd! 24.7fF
C2217 diff_221160_159720# gnd! 24.7fF
C2218 diff_219120_159720# gnd! 24.7fF
C2219 diff_217080_159720# gnd! 24.7fF
C2220 diff_215040_159720# gnd! 24.7fF
C2221 diff_213000_159720# gnd! 24.7fF
C2222 diff_210960_159720# gnd! 24.7fF
C2223 diff_208920_159720# gnd! 24.7fF
C2224 diff_206880_159720# gnd! 24.7fF
C2225 diff_204840_159720# gnd! 24.7fF
C2226 diff_202800_159720# gnd! 24.7fF
C2227 diff_200760_159720# gnd! 24.7fF
C2228 diff_198720_159720# gnd! 24.7fF
C2229 diff_196680_159720# gnd! 24.7fF
C2230 diff_194640_159720# gnd! 24.7fF
C2231 diff_192600_159720# gnd! 24.7fF
C2232 diff_190560_159720# gnd! 24.7fF
C2233 diff_188520_159720# gnd! 24.7fF
C2234 diff_186480_159720# gnd! 24.7fF
C2235 diff_184440_159720# gnd! 24.7fF
C2236 diff_182400_159720# gnd! 24.7fF
C2237 diff_180360_159720# gnd! 24.7fF
C2238 diff_178320_159720# gnd! 24.7fF
C2239 diff_176280_159720# gnd! 24.7fF
C2240 diff_174240_159720# gnd! 24.7fF
C2241 diff_172200_159720# gnd! 24.7fF
C2242 diff_170160_159720# gnd! 24.7fF
C2243 diff_168120_159720# gnd! 24.7fF
C2244 diff_166080_159720# gnd! 24.7fF
C2245 diff_164040_159720# gnd! 24.7fF
C2246 diff_162000_159720# gnd! 24.7fF
C2247 diff_159960_159720# gnd! 24.7fF
C2248 diff_157920_159720# gnd! 24.7fF
C2249 diff_155880_159720# gnd! 24.7fF
C2250 diff_153840_159720# gnd! 24.7fF
C2251 diff_151800_159720# gnd! 24.7fF
C2252 diff_149760_159720# gnd! 24.7fF
C2253 diff_147720_159720# gnd! 24.7fF
C2254 diff_145680_159720# gnd! 24.7fF
C2255 diff_143640_159720# gnd! 24.7fF
C2256 diff_141600_159720# gnd! 24.7fF
C2257 diff_139560_159720# gnd! 24.7fF
C2258 diff_137520_159720# gnd! 24.7fF
C2259 diff_135480_159720# gnd! 24.7fF
C2260 diff_133440_159720# gnd! 24.7fF
C2261 diff_131400_159720# gnd! 24.7fF
C2262 diff_129360_159720# gnd! 24.7fF
C2263 diff_127320_159720# gnd! 24.7fF
C2264 diff_125280_159720# gnd! 24.7fF
C2265 diff_123240_159720# gnd! 24.7fF
C2266 diff_121200_159720# gnd! 24.7fF
C2267 diff_119160_159720# gnd! 24.7fF
C2268 diff_117120_159720# gnd! 24.7fF
C2269 diff_115080_159720# gnd! 24.7fF
C2270 diff_113040_159720# gnd! 24.7fF
C2271 diff_111000_159720# gnd! 24.7fF
C2272 diff_108960_159720# gnd! 24.7fF
C2273 diff_106920_159720# gnd! 24.7fF
C2274 diff_104880_159720# gnd! 24.7fF
C2275 diff_102840_159720# gnd! 24.7fF
C2276 diff_100800_159720# gnd! 24.7fF
C2277 diff_100440_161280# gnd! 613.3fF
C2278 diff_229320_161880# gnd! 26.2fF
C2279 diff_227280_161880# gnd! 26.2fF
C2280 diff_225240_161880# gnd! 26.2fF
C2281 diff_223200_161880# gnd! 26.2fF
C2282 diff_221160_161880# gnd! 26.2fF
C2283 diff_219120_161880# gnd! 26.2fF
C2284 diff_217080_161880# gnd! 26.2fF
C2285 diff_215040_161880# gnd! 26.2fF
C2286 diff_213000_161880# gnd! 26.2fF
C2287 diff_210960_161880# gnd! 26.2fF
C2288 diff_208920_161880# gnd! 26.2fF
C2289 diff_206880_161880# gnd! 26.2fF
C2290 diff_204840_161880# gnd! 26.2fF
C2291 diff_202800_161880# gnd! 26.2fF
C2292 diff_200760_161880# gnd! 26.2fF
C2293 diff_198720_161880# gnd! 26.2fF
C2294 diff_196680_161880# gnd! 26.2fF
C2295 diff_194640_161880# gnd! 26.2fF
C2296 diff_192600_161880# gnd! 26.2fF
C2297 diff_190560_161880# gnd! 26.2fF
C2298 diff_188520_161880# gnd! 26.2fF
C2299 diff_186480_161880# gnd! 26.2fF
C2300 diff_184440_161880# gnd! 26.2fF
C2301 diff_182400_161880# gnd! 26.2fF
C2302 diff_180360_161880# gnd! 26.2fF
C2303 diff_178320_161880# gnd! 26.2fF
C2304 diff_176280_161880# gnd! 26.2fF
C2305 diff_174240_161880# gnd! 26.2fF
C2306 diff_172200_161880# gnd! 26.2fF
C2307 diff_170160_161880# gnd! 26.2fF
C2308 diff_168120_161880# gnd! 26.2fF
C2309 diff_166080_161880# gnd! 26.2fF
C2310 diff_164040_161880# gnd! 26.2fF
C2311 diff_162000_161880# gnd! 26.2fF
C2312 diff_159960_161880# gnd! 26.2fF
C2313 diff_157920_161880# gnd! 26.2fF
C2314 diff_155880_161880# gnd! 26.2fF
C2315 diff_153840_161880# gnd! 26.2fF
C2316 diff_151800_161880# gnd! 26.2fF
C2317 diff_149760_161880# gnd! 26.2fF
C2318 diff_147720_161880# gnd! 26.2fF
C2319 diff_145680_161880# gnd! 26.2fF
C2320 diff_143640_161880# gnd! 26.2fF
C2321 diff_141600_161880# gnd! 26.2fF
C2322 diff_139560_161880# gnd! 26.2fF
C2323 diff_137520_161880# gnd! 26.2fF
C2324 diff_135480_161880# gnd! 26.2fF
C2325 diff_133440_161880# gnd! 26.2fF
C2326 diff_131400_161880# gnd! 26.2fF
C2327 diff_129360_161880# gnd! 26.2fF
C2328 diff_127320_161880# gnd! 26.2fF
C2329 diff_125280_161880# gnd! 26.2fF
C2330 diff_123240_161880# gnd! 26.2fF
C2331 diff_121200_161880# gnd! 26.2fF
C2332 diff_119160_161880# gnd! 26.2fF
C2333 diff_117120_161880# gnd! 26.2fF
C2334 diff_115080_161880# gnd! 26.2fF
C2335 diff_113040_161880# gnd! 26.2fF
C2336 diff_111000_161880# gnd! 26.2fF
C2337 diff_108960_161880# gnd! 26.2fF
C2338 diff_106920_161880# gnd! 26.2fF
C2339 diff_104880_161880# gnd! 26.2fF
C2340 diff_102840_161880# gnd! 26.2fF
C2341 diff_100800_161880# gnd! 26.2fF
C2342 diff_100440_163560# gnd! 644.8fF
C2343 diff_229320_164160# gnd! 24.7fF
C2344 diff_227280_164160# gnd! 24.7fF
C2345 diff_225240_164160# gnd! 24.7fF
C2346 diff_223200_164160# gnd! 24.7fF
C2347 diff_221160_164160# gnd! 24.7fF
C2348 diff_219120_164160# gnd! 24.7fF
C2349 diff_217080_164160# gnd! 24.7fF
C2350 diff_215040_164160# gnd! 24.7fF
C2351 diff_213000_164160# gnd! 24.7fF
C2352 diff_210960_164160# gnd! 24.7fF
C2353 diff_208920_164160# gnd! 24.7fF
C2354 diff_206880_164160# gnd! 24.7fF
C2355 diff_204840_164160# gnd! 24.7fF
C2356 diff_202800_164160# gnd! 24.7fF
C2357 diff_200760_164160# gnd! 24.7fF
C2358 diff_198720_164160# gnd! 24.7fF
C2359 diff_196680_164160# gnd! 24.7fF
C2360 diff_194640_164160# gnd! 24.7fF
C2361 diff_192600_164160# gnd! 24.7fF
C2362 diff_190560_164160# gnd! 24.7fF
C2363 diff_188520_164160# gnd! 24.7fF
C2364 diff_186480_164160# gnd! 24.7fF
C2365 diff_184440_164160# gnd! 24.7fF
C2366 diff_182400_164160# gnd! 24.7fF
C2367 diff_180360_164160# gnd! 24.7fF
C2368 diff_178320_164160# gnd! 24.7fF
C2369 diff_176280_164160# gnd! 24.7fF
C2370 diff_174240_164160# gnd! 24.7fF
C2371 diff_172200_164160# gnd! 24.7fF
C2372 diff_170160_164160# gnd! 24.7fF
C2373 diff_168120_164160# gnd! 24.7fF
C2374 diff_166080_164160# gnd! 24.7fF
C2375 diff_164040_164160# gnd! 24.7fF
C2376 diff_162000_164160# gnd! 24.7fF
C2377 diff_159960_164160# gnd! 24.7fF
C2378 diff_157920_164160# gnd! 24.7fF
C2379 diff_155880_164160# gnd! 24.7fF
C2380 diff_153840_164160# gnd! 24.7fF
C2381 diff_151800_164160# gnd! 24.7fF
C2382 diff_149760_164160# gnd! 24.7fF
C2383 diff_147720_164160# gnd! 24.7fF
C2384 diff_145680_164160# gnd! 24.7fF
C2385 diff_143640_164160# gnd! 24.7fF
C2386 diff_141600_164160# gnd! 24.7fF
C2387 diff_139560_164160# gnd! 24.7fF
C2388 diff_137520_164160# gnd! 24.7fF
C2389 diff_135480_164160# gnd! 24.7fF
C2390 diff_133440_164160# gnd! 24.7fF
C2391 diff_131400_164160# gnd! 24.7fF
C2392 diff_129360_164160# gnd! 24.7fF
C2393 diff_127320_164160# gnd! 24.7fF
C2394 diff_125280_164160# gnd! 24.7fF
C2395 diff_123240_164160# gnd! 24.7fF
C2396 diff_121200_164160# gnd! 24.7fF
C2397 diff_119160_164160# gnd! 24.7fF
C2398 diff_117120_164160# gnd! 24.7fF
C2399 diff_115080_164160# gnd! 24.7fF
C2400 diff_113040_164160# gnd! 24.7fF
C2401 diff_111000_164160# gnd! 24.7fF
C2402 diff_108960_164160# gnd! 24.7fF
C2403 diff_106920_164160# gnd! 24.7fF
C2404 diff_104880_164160# gnd! 24.7fF
C2405 diff_102840_164160# gnd! 24.7fF
C2406 diff_100800_164160# gnd! 24.7fF
C2407 diff_88680_154680# gnd! 88.0fF
C2408 diff_83160_150480# gnd! 90.3fF
C2409 diff_82080_136560# gnd! 612.4fF
C2410 diff_73800_150600# gnd! 88.4fF
C2411 diff_67320_150600# gnd! 97.3fF
C2412 diff_66480_136560# gnd! 604.0fF
C2413 diff_18960_80400# gnd! 1890.3fF
C2414 diff_58320_150600# gnd! 94.7fF
C2415 diff_52080_150360# gnd! 89.9fF
C2416 diff_51000_136680# gnd! 615.1fF
C2417 diff_42840_150720# gnd! 90.8fF
C2418 diff_36600_150480# gnd! 94.2fF
C2419 diff_100440_165720# gnd! 642.3fF
C2420 diff_250560_91920# gnd! 844.5fF
C2421 diff_248880_85320# gnd! 854.9fF
C2422 diff_236760_167400# gnd! 499.8fF
C2423 diff_229320_166320# gnd! 26.2fF
C2424 diff_227280_166320# gnd! 26.2fF
C2425 diff_225240_166320# gnd! 26.2fF
C2426 diff_223200_166320# gnd! 26.2fF
C2427 diff_221160_166320# gnd! 26.2fF
C2428 diff_219120_166320# gnd! 26.2fF
C2429 diff_217080_166320# gnd! 26.2fF
C2430 diff_215040_166320# gnd! 26.2fF
C2431 diff_213000_166320# gnd! 26.2fF
C2432 diff_210960_166320# gnd! 26.2fF
C2433 diff_208920_166320# gnd! 26.2fF
C2434 diff_206880_166320# gnd! 26.2fF
C2435 diff_204840_166320# gnd! 26.2fF
C2436 diff_202800_166320# gnd! 26.2fF
C2437 diff_200760_166320# gnd! 26.2fF
C2438 diff_198720_166320# gnd! 26.2fF
C2439 diff_196680_166320# gnd! 26.2fF
C2440 diff_194640_166320# gnd! 26.2fF
C2441 diff_192600_166320# gnd! 26.2fF
C2442 diff_190560_166320# gnd! 26.2fF
C2443 diff_188520_166320# gnd! 26.2fF
C2444 diff_186480_166320# gnd! 26.2fF
C2445 diff_184440_166320# gnd! 26.2fF
C2446 diff_182400_166320# gnd! 26.2fF
C2447 diff_180360_166320# gnd! 26.2fF
C2448 diff_178320_166320# gnd! 26.2fF
C2449 diff_176280_166320# gnd! 26.2fF
C2450 diff_174240_166320# gnd! 26.2fF
C2451 diff_172200_166320# gnd! 26.2fF
C2452 diff_170160_166320# gnd! 26.2fF
C2453 diff_168120_166320# gnd! 26.2fF
C2454 diff_166080_166320# gnd! 26.2fF
C2455 diff_164040_166320# gnd! 26.2fF
C2456 diff_162000_166320# gnd! 26.2fF
C2457 diff_159960_166320# gnd! 26.2fF
C2458 diff_157920_166320# gnd! 26.2fF
C2459 diff_155880_166320# gnd! 26.2fF
C2460 diff_153840_166320# gnd! 26.2fF
C2461 diff_151800_166320# gnd! 26.2fF
C2462 diff_149760_166320# gnd! 26.2fF
C2463 diff_147720_166320# gnd! 26.2fF
C2464 diff_145680_166320# gnd! 26.2fF
C2465 diff_143640_166320# gnd! 26.2fF
C2466 diff_141600_166320# gnd! 26.2fF
C2467 diff_139560_166320# gnd! 26.2fF
C2468 diff_137520_166320# gnd! 26.2fF
C2469 diff_135480_166320# gnd! 26.2fF
C2470 diff_133440_166320# gnd! 26.2fF
C2471 diff_131400_166320# gnd! 26.2fF
C2472 diff_129360_166320# gnd! 26.2fF
C2473 diff_127320_166320# gnd! 26.2fF
C2474 diff_125280_166320# gnd! 26.2fF
C2475 diff_123240_166320# gnd! 26.2fF
C2476 diff_121200_166320# gnd! 26.2fF
C2477 diff_119160_166320# gnd! 26.2fF
C2478 diff_117120_166320# gnd! 26.2fF
C2479 diff_115080_166320# gnd! 26.2fF
C2480 diff_113040_166320# gnd! 26.2fF
C2481 diff_111000_166320# gnd! 26.2fF
C2482 diff_108960_166320# gnd! 26.2fF
C2483 diff_106920_166320# gnd! 26.2fF
C2484 diff_104880_166320# gnd! 26.2fF
C2485 diff_102840_166320# gnd! 26.2fF
C2486 diff_100800_166320# gnd! 26.2fF
C2487 diff_100440_168000# gnd! 607.3fF
C2488 diff_243120_97920# gnd! 701.5fF
C2489 diff_241320_99600# gnd! 740.5fF
C2490 diff_238440_42720# gnd! 721.5fF
C2491 diff_236160_42720# gnd! 748.2fF
C2492 diff_100800_168600# gnd! 2732.1fF
C2493 diff_165720_170280# gnd! 1786.5fF
C2494 diff_266400_168600# gnd! 153.5fF
C2495 diff_264960_142800# gnd! 296.5fF
C2496 diff_261360_171960# gnd! 236.2fF
C2497 diff_243720_169800# gnd! 1171.5fF
C2498 diff_100320_170280# gnd! 1986.6fF
C2499 diff_243360_174240# gnd! 1155.5fF
C2500 diff_275160_168600# gnd! 129.0fF
C2501 diff_280200_173280# gnd! 101.5fF
C2502 diff_80400_166200# gnd! 965.5fF
C2503 diff_64920_166200# gnd! 967.9fF
C2504 Vdd gnd! 19277.9fF
C2505 diff_35520_136680# gnd! 615.1fF
C2506 diff_49440_166200# gnd! 978.3fF
C2507 diff_33840_166200# gnd! 977.5fF
C2508 d0 gnd! 3375.1fF
C2509 d1 gnd! 3489.1fF
C2510 d3 gnd! 4191.8fF
C2511 sync gnd! 2776.3fF
C2512 d2 gnd! 3420.1fF
C2513 clk1 gnd! 2695.6fF
C2514 clk2 gnd! 3523.0fF
