* SPICE3 file created from 6502.ext - technology: nmos

.option scale=2u

M1000 nmi GND GND GND efet w=52 l=8
+ ad=4427 pd=1102 as=1.6652e+06 ps=281796 
M1001 GND nmi n_1392 GND efet w=70 l=7
+ ad=0 pd=0 as=820 ps=206 
M1002 n_1392 n_1392 Vdd GND dfet w=9 l=12
+ ad=2118 pd=670 as=0 ps=0 
M1003 GND pipeT4out n_1703 GND efet w=110 l=7
+ ad=0 pd=0 as=1351 ps=352 
M1004 n_468 n_16 n_1703 GND efet w=59 l=7
+ ad=886 pd=306 as=0 ps=0 
M1005 GND pipeT4out n_395 GND efet w=124 l=7
+ ad=0 pd=0 as=820 ps=244 
M1006 GND pipeT5out n_1615 GND efet w=117 l=7
+ ad=0 pd=0 as=1117 ps=318 
M1007 n_1615 notRdy0 n_468 GND efet w=74 l=7
+ ad=0 pd=0 as=0 ps=0 
M1008 n_378 n_18 GND GND efet w=66 l=6
+ ad=1274 pd=348 as=0 ps=0 
M1009 Vdd n_468 n_468 GND dfet w=10 l=17
+ ad=0 pd=0 as=404 ps=104 
M1010 n_395 notRdy0 n_472 GND efet w=48 l=6
+ ad=0 pd=0 as=1079 ps=284 
M1011 GND n_378 _t5 GND efet w=73 l=6
+ ad=0 pd=0 as=1001 ps=238 
M1012 pipeT5out cclk n_378 GND efet w=12 l=9
+ ad=191 pd=76 as=0 ps=0 
M1013 GND n_1392 n_284 GND efet w=37 l=7
+ ad=0 pd=0 as=517 ps=138 
M1014 GND NMIP n_645 GND efet w=43 l=6
+ ad=0 pd=0 as=796 ps=278 
M1015 n_891 cclk GND GND efet w=46 l=7
+ ad=472 pd=128 as=0 ps=0 
M1016 n_468 cp1 n_18 GND efet w=12 l=8
+ ad=0 pd=0 as=320 ps=102 
M1017 pipeT4out cclk n_188 GND efet w=12 l=8
+ ad=251 pd=92 as=1730 ps=456 
M1018 n_472 n_16 n_1366 GND efet w=55 l=7
+ ad=0 pd=0 as=1107 ps=278 
M1019 GND pipeT3out n_1366 GND efet w=110 l=7
+ ad=0 pd=0 as=0 ps=0 
M1020 n_378 n_378 Vdd GND dfet w=10 l=17
+ ad=930 pd=288 as=0 ps=0 
M1021 GND n_1357 n_378 GND efet w=47 l=7
+ ad=0 pd=0 as=0 ps=0 
M1022 NMIP n_284 n_891 GND efet w=48 l=7
+ ad=961 pd=280 as=0 ps=0 
M1023 n_284 n_284 Vdd GND dfet w=10 l=12
+ ad=991 pd=306 as=0 ps=0 
M1024 GND nNMIP NMIP GND efet w=25 l=7
+ ad=0 pd=0 as=0 ps=0 
M1025 nNMIP NMIP GND GND efet w=25 l=6
+ ad=725 pd=218 as=0 ps=0 
M1026 n_346 n_1392 nNMIP GND efet w=47 l=7
+ ad=235 pd=104 as=0 ps=0 
M1027 GND cclk n_346 GND efet w=47 l=6
+ ad=0 pd=0 as=0 ps=0 
M1028 irq GND GND GND efet w=51 l=8
+ ad=4660 pd=1162 as=0 ps=0 
M1029 Vdd n_472 n_472 GND dfet w=10 l=16
+ ad=0 pd=0 as=390 ps=100 
M1030 _t5 _t5 Vdd GND dfet w=10 l=6
+ ad=20517 pd=6238 as=0 ps=0 
M1031 n_645 n_645 Vdd GND dfet w=9 l=10
+ ad=6071 pd=2006 as=0 ps=0 
M1032 NMIP NMIP Vdd GND dfet w=7 l=14
+ ad=1419 pd=468 as=0 ps=0 
M1033 nNMIP nNMIP Vdd GND dfet w=10 l=16
+ ad=804 pd=222 as=0 ps=0 
M1034 GND irq n_1599 GND efet w=62 l=6
+ ad=0 pd=0 as=850 ps=210 
M1035 n_881 cclk GND GND efet w=53 l=6
+ ad=808 pd=172 as=0 ps=0 
M1036 n_538 n_1599 GND GND efet w=33 l=6
+ ad=583 pd=146 as=0 ps=0 
M1037 GND n_807 n_330 GND efet w=24 l=7
+ ad=0 pd=0 as=1391 ps=324 
M1038 n_431 n_1599 n_807 GND efet w=58 l=6
+ ad=650 pd=172 as=970 ps=244 
M1039 n_1599 n_1599 Vdd GND dfet w=11 l=13
+ ad=2239 pd=704 as=0 ps=0 
M1040 n_538 n_538 Vdd GND dfet w=10 l=12
+ ad=741 pd=224 as=0 ps=0 
M1041 n_881 n_538 n_330 GND efet w=54 l=6
+ ad=0 pd=0 as=0 ps=0 
M1042 GND n_330 n_807 GND efet w=33 l=7
+ ad=0 pd=0 as=0 ps=0 
M1043 GND cclk n_431 GND efet w=46 l=7
+ ad=0 pd=0 as=0 ps=0 
M1044 n_806 GND GND GND efet w=46 l=8
+ ad=3480 pd=272 as=0 ps=0 
M1045 n_807 n_807 Vdd GND dfet w=9 l=14
+ ad=770 pd=244 as=0 ps=0 
M1046 GND IRQP nIRQP GND efet w=42 l=6
+ ad=0 pd=0 as=1104 ps=240 
M1047 n_330 n_330 Vdd GND dfet w=10 l=14
+ ad=625 pd=196 as=0 ps=0 
M1048 IRQP cp1 n_330 GND efet w=12 l=8
+ ad=136 pd=70 as=0 ps=0 
M1049 GND IRQP nIRQP GND efet w=48 l=7
+ ad=0 pd=0 as=0 ps=0 
M1050 nIRQP nIRQP Vdd GND dfet w=11 l=10
+ ad=5075 pd=1750 as=0 ps=0 
M1051 clk1out n_1417 GND GND efet w=104 l=6
+ ad=12284 pd=1634 as=0 ps=0 
M1052 GND n_1417 clk1out GND efet w=221 l=6
+ ad=0 pd=0 as=0 ps=0 
M1053 clk1out n_1417 GND GND efet w=221 l=7
+ ad=0 pd=0 as=0 ps=0 
M1054 GND n_1417 clk1out GND efet w=221 l=6
+ ad=0 pd=0 as=0 ps=0 
M1055 clk1out n_1417 GND GND efet w=221 l=6
+ ad=0 pd=0 as=0 ps=0 
M1056 GND n_747 n_1417 GND efet w=226 l=7
+ ad=0 pd=0 as=3742 ps=524 
M1057 GND n_670 n_747 GND efet w=276 l=7
+ ad=0 pd=0 as=4486 ps=612 
M1058 GND GND rdy GND efet w=51 l=7
+ ad=0 pd=0 as=4872 ps=1250 
M1059 GND rdy n_958 GND efet w=149 l=8
+ ad=0 pd=0 as=1524 ps=410 
M1060 rdy rdy Vdd GND dfet w=10 l=16
+ ad=2328 pd=682 as=0 ps=0 
M1061 n_420 n_865 GND GND efet w=54 l=7
+ ad=893 pd=296 as=0 ps=0 
M1062 n_47 cp1 n_420 GND efet w=13 l=7
+ ad=153 pd=64 as=0 ps=0 
M1063 n_1449 n_958 GND GND efet w=118 l=6
+ ad=1196 pd=356 as=0 ps=0 
M1064 n_865 cclk n_958 GND efet w=13 l=8
+ ad=173 pd=64 as=0 ps=0 
M1065 GND n_47 n_603 GND efet w=50 l=7
+ ad=0 pd=0 as=561 ps=162 
M1066 clk1out n_747 Vdd GND dfet w=68 l=7
+ ad=0 pd=0 as=568855 ps=107108 
M1067 n_1417 n_670 Vdd GND dfet w=25 l=8
+ ad=0 pd=0 as=0 ps=0 
M1068 Vdd n_747 n_747 GND dfet w=26 l=8
+ ad=0 pd=0 as=2832 ps=816 
M1069 n_420 n_420 Vdd GND dfet w=10 l=17
+ ad=475 pd=108 as=0 ps=0 
M1070 n_958 n_958 Vdd GND dfet w=9 l=6
+ ad=1625 pd=528 as=0 ps=0 
M1071 n_603 n_603 Vdd GND dfet w=10 l=17
+ ad=5483 pd=1802 as=0 ps=0 
M1072 clk2out n_135 GND GND efet w=332 l=7
+ ad=10493 pd=1504 as=0 ps=0 
M1073 GND GND res GND efet w=78 l=7
+ ad=0 pd=0 as=5344 ps=1320 
M1074 n_312 res GND GND efet w=78 l=6
+ ad=963 pd=278 as=0 ps=0 
M1075 Vdd n_1449 n_1449 GND dfet w=16 l=7
+ ad=0 pd=0 as=8170 ps=2998 
M1076 GND n_312 n_995 GND efet w=32 l=6
+ ad=0 pd=0 as=587 ps=156 
M1077 n_886 cclk GND GND efet w=47 l=6
+ ad=235 pd=104 as=0 ps=0 
M1078 n_975 n_995 n_886 GND efet w=47 l=7
+ ad=767 pd=192 as=0 ps=0 
M1079 GND n_854 n_975 GND efet w=25 l=6
+ ad=0 pd=0 as=0 ps=0 
M1080 n_854 n_975 GND GND efet w=25 l=6
+ ad=981 pd=314 as=0 ps=0 
M1081 n_742 n_312 n_854 GND efet w=47 l=6
+ ad=235 pd=104 as=0 ps=0 
M1082 GND cclk n_742 GND efet w=47 l=7
+ ad=0 pd=0 as=0 ps=0 
M1083 GND n_1395 Reset0 GND efet w=78 l=7
+ ad=0 pd=0 as=1666 ps=418 
M1084 n_1395 cp1 n_854 GND efet w=12 l=8
+ ad=161 pd=62 as=0 ps=0 
M1085 n_312 n_312 Vdd GND dfet w=10 l=12
+ ad=1617 pd=538 as=0 ps=0 
M1086 n_995 n_995 Vdd GND dfet w=11 l=12
+ ad=1216 pd=386 as=0 ps=0 
M1087 n_975 n_975 Vdd GND dfet w=9 l=14
+ ad=646 pd=192 as=0 ps=0 
M1088 n_854 n_854 Vdd GND dfet w=9 l=14
+ ad=1439 pd=486 as=0 ps=0 
M1089 Reset0 n_1395 GND GND efet w=71 l=7
+ ad=0 pd=0 as=0 ps=0 
M1090 GND n_519 n_670 GND efet w=88 l=7
+ ad=0 pd=0 as=2095 ps=486 
M1091 Vdd Reset0 Reset0 GND dfet w=10 l=9
+ ad=0 pd=0 as=14236 ps=4882 
M1092 n_670 n_670 Vdd GND dfet w=25 l=7
+ ad=3856 pd=1154 as=0 ps=0 
M1093 GND n_519 n_670 GND efet w=85 l=9
+ ad=0 pd=0 as=0 ps=0 
M1094 clk2out n_135 GND GND efet w=236 l=7
+ ad=0 pd=0 as=0 ps=0 
M1095 GND n_135 clk2out GND efet w=236 l=6
+ ad=0 pd=0 as=0 ps=0 
M1096 clk2out n_135 GND GND efet w=236 l=8
+ ad=0 pd=0 as=0 ps=0 
M1097 Vdd n_127 clk2out GND dfet w=67 l=7
+ ad=0 pd=0 as=0 ps=0 
M1098 n_135 n_519 Vdd GND dfet w=24 l=7
+ ad=2286 pd=512 as=0 ps=0 
M1099 GND n_127 n_135 GND efet w=222 l=6
+ ad=0 pd=0 as=0 ps=0 
M1100 n_127 cp1 GND GND efet w=126 l=7
+ ad=3045 pd=648 as=0 ps=0 
M1101 GND n_519 n_127 GND efet w=226 l=6
+ ad=0 pd=0 as=0 ps=0 
M1102 GND clk0 n_519 GND efet w=280 l=6
+ ad=0 pd=0 as=2799 ps=644 
M1103 GND GND so GND efet w=46 l=7
+ ad=0 pd=0 as=6079 ps=1468 
M1104 clk0 GND GND GND efet w=55 l=7
+ ad=8528 pd=1926 as=0 ps=0 
M1105 n_127 n_127 Vdd GND dfet w=25 l=8
+ ad=3702 pd=1134 as=0 ps=0 
M1106 n_519 n_519 Vdd GND dfet w=25 l=7
+ ad=5789 pd=1744 as=0 ps=0 
M1107 n_1650 cp1 n_94 GND efet w=12 l=8
+ ad=1479 pd=346 as=222 ps=78 
M1108 so so Vdd GND dfet w=10 l=16
+ ad=2070 pd=662 as=0 ps=0 
M1109 n_1069 n_1024 GND GND efet w=30 l=7
+ ad=1358 pd=336 as=0 ps=0 
M1110 n_1069 n_1069 Vdd GND dfet w=10 l=13
+ ad=4549 pd=1504 as=0 ps=0 
M1111 GND n_1274 n_1069 GND efet w=63 l=7
+ ad=0 pd=0 as=0 ps=0 
M1112 n_1024 cclk n_1699 GND efet w=12 l=7
+ ad=1654 pd=462 as=140 ps=74 
M1113 n_913 n_1699 GND GND efet w=44 l=6
+ ad=743 pd=232 as=0 ps=0 
M1114 GND n_94 n_1024 GND efet w=63 l=6
+ ad=0 pd=0 as=0 ps=0 
M1115 n_913 cp1 n_1274 GND efet w=12 l=8
+ ad=0 pd=0 as=220 ps=72 
M1116 n_1024 n_1024 Vdd GND dfet w=10 l=14
+ ad=701 pd=222 as=0 ps=0 
M1117 GND so n_1650 GND efet w=123 l=7
+ ad=0 pd=0 as=0 ps=0 
M1118 Vdd op_sty_cpy_mem op_sty_cpy_mem GND dfet w=9 l=19
+ ad=0 pd=0 as=2542 ps=746 
M1119 Vdd _t4 _t4 GND dfet w=9 l=6
+ ad=0 pd=0 as=18491 ps=6132 
M1120 n_472 cp1 n_1606 GND efet w=12 l=8
+ ad=0 pd=0 as=185 ps=80 
M1121 Vdd n_188 n_188 GND dfet w=10 l=13
+ ad=0 pd=0 as=1409 ps=416 
M1122 _t4 n_188 GND GND efet w=96 l=7
+ ad=611 pd=206 as=0 ps=0 
M1123 n_188 n_1606 GND GND efet w=74 l=6
+ ad=0 pd=0 as=0 ps=0 
M1124 Vdd op_T2_abs_y op_T2_abs_y GND dfet w=9 l=19
+ ad=0 pd=0 as=795 ps=204 
M1125 Vdd op_T3_ind_y op_T3_ind_y GND dfet w=9 l=18
+ ad=0 pd=0 as=1128 ps=338 
M1126 Vdd x_op_T0_tya x_op_T0_tya GND dfet w=9 l=19
+ ad=0 pd=0 as=862 ps=216 
M1127 Vdd op_T0_iny_dey op_T0_iny_dey GND dfet w=10 l=19
+ ad=0 pd=0 as=808 ps=224 
M1128 Vdd op_xy op_xy GND dfet w=9 l=19
+ ad=0 pd=0 as=2026 ps=600 
M1129 Vdd op_T0_cpy_iny op_T0_cpy_iny GND dfet w=9 l=19
+ ad=0 pd=0 as=795 ps=228 
M1130 Vdd op_T2_idx_x_xy op_T2_idx_x_xy GND dfet w=10 l=19
+ ad=0 pd=0 as=2345 ps=710 
M1131 Vdd x_op_T0_txa x_op_T0_txa GND dfet w=10 l=19
+ ad=0 pd=0 as=765 ps=204 
M1132 Vdd op_T0_cpx_inx op_T0_cpx_inx GND dfet w=9 l=18
+ ad=0 pd=0 as=777 ps=202 
M1133 Vdd op_T2_ind_x op_T2_ind_x GND dfet w=10 l=19
+ ad=0 pd=0 as=839 ps=234 
M1134 Vdd op_T0_dex op_T0_dex GND dfet w=9 l=19
+ ad=0 pd=0 as=777 ps=226 
M1135 Vdd op_T0_txs op_T0_txs GND dfet w=9 l=19
+ ad=0 pd=0 as=1952 ps=628 
M1136 Vdd op_from_x op_from_x GND dfet w=10 l=19
+ ad=0 pd=0 as=2502 ps=808 
M1137 Vdd op_T__dex op_T__dex GND dfet w=9 l=18
+ ad=0 pd=0 as=605 ps=180 
M1138 Vdd op_T0_ldx_tax_tsx op_T0_ldx_tax_tsx GND dfet w=11 l=19
+ ad=0 pd=0 as=862 ps=256 
M1139 Vdd op_T0_tsx op_T0_tsx GND dfet w=10 l=19
+ ad=0 pd=0 as=1472 ps=446 
M1140 Vdd op_T0_ldy_mem op_T0_ldy_mem GND dfet w=9 l=19
+ ad=0 pd=0 as=878 ps=238 
M1141 Vdd op_T__inx op_T__inx GND dfet w=9 l=19
+ ad=0 pd=0 as=767 ps=224 
M1142 Vdd op_T__iny_dey op_T__iny_dey GND dfet w=9 l=19
+ ad=0 pd=0 as=699 ps=212 
M1143 Vdd op_T0_tay_ldy_not_idx op_T0_tay_ldy_not_idx GND dfet w=9 l=19
+ ad=0 pd=0 as=864 ps=256 
M1144 Vdd op_T5_brk op_T5_brk GND dfet w=10 l=19
+ ad=0 pd=0 as=1275 ps=352 
M1145 Vdd op_T0_jsr op_T0_jsr GND dfet w=10 l=19
+ ad=0 pd=0 as=2036 ps=634 
M1146 Vdd op_T4_rts op_T4_rts GND dfet w=10 l=19
+ ad=0 pd=0 as=743 ps=192 
M1147 Vdd op_T5_rti op_T5_rti GND dfet w=9 l=19
+ ad=0 pd=0 as=4773 ps=1708 
M1148 Vdd op_T0_php_pha op_T0_php_pha GND dfet w=10 l=19
+ ad=0 pd=0 as=785 ps=216 
M1149 Vdd op_T3_plp_pla op_T3_plp_pla GND dfet w=9 l=19
+ ad=0 pd=0 as=836 ps=226 
M1150 Vdd op_T2 op_T2 GND dfet w=10 l=19
+ ad=0 pd=0 as=4990 ps=1666 
M1151 Vdd op_ror op_ror GND dfet w=11 l=19
+ ad=0 pd=0 as=2130 ps=656 
M1152 Vdd op_jmp op_jmp GND dfet w=9 l=19
+ ad=0 pd=0 as=1886 ps=594 
M1153 Vdd op_T0_eor op_T0_eor GND dfet w=10 l=19
+ ad=0 pd=0 as=2670 ps=900 
M1154 Vdd op_T0_ora op_T0_ora GND dfet w=9 l=19
+ ad=0 pd=0 as=2308 ps=698 
M1155 Vdd op_T2_abs op_T2_abs GND dfet w=10 l=19
+ ad=0 pd=0 as=1987 ps=628 
M1156 Vdd op_T0 op_T0 GND dfet w=9 l=19
+ ad=0 pd=0 as=1077 ps=308 
M1157 Vdd op_T2_ADL_ADD op_T2_ADL_ADD GND dfet w=9 l=19
+ ad=0 pd=0 as=1881 ps=602 
M1158 Vdd op_T3_stack_bit_jmp op_T3_stack_bit_jmp GND dfet w=10 l=19
+ ad=0 pd=0 as=803 ps=214 
M1159 Vdd op_T2_stack op_T2_stack GND dfet w=9 l=19
+ ad=0 pd=0 as=1898 ps=590 
M1160 Vdd op_T4_rti op_T4_rti GND dfet w=10 l=19
+ ad=0 pd=0 as=717 ps=196 
M1161 Vdd op_T4_brk_jsr op_T4_brk_jsr GND dfet w=10 l=19
+ ad=0 pd=0 as=830 ps=236 
M1162 Vdd op_T4_ind_y op_T4_ind_y GND dfet w=9 l=19
+ ad=0 pd=0 as=946 ps=282 
M1163 Vdd op_T3_ind_x op_T3_ind_x GND dfet w=10 l=19
+ ad=0 pd=0 as=1171 ps=402 
M1164 Vdd op_T3_abs_idx op_T3_abs_idx GND dfet w=9 l=19
+ ad=0 pd=0 as=958 ps=278 
M1165 Vdd op_T2_ind_y op_T2_ind_y GND dfet w=9 l=18
+ ad=0 pd=0 as=1021 ps=292 
M1166 Vdd op_inc_nop op_inc_nop GND dfet w=9 l=19
+ ad=0 pd=0 as=1199 ps=310 
M1167 Vdd op_plp_pla op_plp_pla GND dfet w=10 l=19
+ ad=0 pd=0 as=946 ps=290 
M1168 Vdd x_op_T3_ind_y x_op_T3_ind_y GND dfet w=9 l=18
+ ad=0 pd=0 as=828 ps=226 
M1169 Vdd op_T4_ind_x op_T4_ind_x GND dfet w=9 l=19
+ ad=0 pd=0 as=1896 ps=628 
M1170 Vdd op_T2_jsr op_T2_jsr GND dfet w=9 l=19
+ ad=0 pd=0 as=2351 ps=756 
M1171 Vdd op_rti_rts op_rti_rts GND dfet w=9 l=19
+ ad=0 pd=0 as=2456 ps=754 
M1172 Vdd op_T0_cmp op_T0_cmp GND dfet w=9 l=19
+ ad=0 pd=0 as=849 ps=236 
M1173 Vdd op_T0_cpx_cpy_inx_iny op_T0_cpx_cpy_inx_iny GND dfet w=9 l=19
+ ad=0 pd=0 as=896 ps=264 
M1174 Vdd op_T0_adc_sbc op_T0_adc_sbc GND dfet w=9 l=19
+ ad=0 pd=0 as=3638 ps=1278 
M1175 Vdd op_T3_jmp op_T3_jmp GND dfet w=9 l=19
+ ad=0 pd=0 as=838 ps=232 
M1176 Vdd op_T0_sbc op_T0_sbc GND dfet w=9 l=19
+ ad=0 pd=0 as=5052 ps=1690 
M1177 Vdd op_rol_ror op_rol_ror GND dfet w=10 l=19
+ ad=0 pd=0 as=1142 ps=324 
M1178 Vdd op_T5_jsr op_T5_jsr GND dfet w=10 l=19
+ ad=0 pd=0 as=2713 ps=926 
M1179 op_shift op_shift Vdd GND dfet w=10 l=19
+ ad=1861 pd=568 as=0 ps=0 
M1180 Vdd op_T0_tya op_T0_tya GND dfet w=9 l=18
+ ad=0 pd=0 as=870 ps=230 
M1181 Vdd op_T2_stack_access op_T2_stack_access GND dfet w=10 l=19
+ ad=0 pd=0 as=1628 ps=544 
M1182 Vdd op_T__adc_sbc op_T__adc_sbc GND dfet w=10 l=18
+ ad=0 pd=0 as=1099 ps=336 
M1183 GND n_1357 n_188 GND efet w=48 l=6
+ ad=0 pd=0 as=0 ps=0 
M1184 GND pipeT3out n_1456 GND efet w=127 l=7
+ ad=0 pd=0 as=783 ps=246 
M1185 Vdd op_T__ora_and_eor_adc op_T__ora_and_eor_adc GND dfet w=8 l=19
+ ad=0 pd=0 as=1440 ps=486 
M1186 Vdd op_T0_txa op_T0_txa GND dfet w=9 l=19
+ ad=0 pd=0 as=850 ps=222 
M1187 Vdd op_T__shift_a op_T__shift_a GND dfet w=9 l=18
+ ad=0 pd=0 as=850 ps=246 
M1188 Vdd op_T0_lda op_T0_lda GND dfet w=10 l=19
+ ad=0 pd=0 as=1105 ps=302 
M1189 Vdd op_T0_pla op_T0_pla GND dfet w=10 l=19
+ ad=0 pd=0 as=830 ps=228 
M1190 Vdd op_T0_tay op_T0_tay GND dfet w=9 l=19
+ ad=0 pd=0 as=834 ps=222 
M1191 Vdd op_T0_acc op_T0_acc GND dfet w=10 l=18
+ ad=0 pd=0 as=985 ps=278 
M1192 Vdd op_T0_tax op_T0_tax GND dfet w=9 l=19
+ ad=0 pd=0 as=923 ps=236 
M1193 Vdd op_T0_shift_a op_T0_shift_a GND dfet w=9 l=19
+ ad=0 pd=0 as=2109 ps=678 
M1194 Vdd op_T0_and op_T0_and GND dfet w=9 l=19
+ ad=0 pd=0 as=977 ps=262 
M1195 Vdd op_T5_ind_y op_T5_ind_y GND dfet w=9 l=19
+ ad=0 pd=0 as=911 ps=256 
M1196 Vdd op_T0_bit op_T0_bit GND dfet w=9 l=19
+ ad=0 pd=0 as=1153 ps=332 
M1197 Vdd op_T4_abs_idx op_T4_abs_idx GND dfet w=10 l=18
+ ad=0 pd=0 as=1128 ps=320 
M1198 Vdd op_branch_done op_branch_done GND dfet w=9 l=18
+ ad=0 pd=0 as=4883 ps=1638 
M1199 Vdd op_T0_shift_right_a op_T0_shift_right_a GND dfet w=9 l=18
+ ad=0 pd=0 as=904 ps=252 
M1200 Vdd op_T2_pha op_T2_pha GND dfet w=10 l=18
+ ad=0 pd=0 as=1736 ps=568 
M1201 Vdd op_T2_brk op_T2_brk GND dfet w=9 l=19
+ ad=0 pd=0 as=782 ps=214 
M1202 op_branch_done n_603 GND GND efet w=18 l=7
+ ad=1375 pd=352 as=0 ps=0 
M1203 Vdd op_shift_right op_shift_right GND dfet w=9 l=19
+ ad=0 pd=0 as=1047 ps=298 
M1204 Vdd op_sta_cmp op_sta_cmp GND dfet w=9 l=18
+ ad=0 pd=0 as=2343 ps=760 
M1205 Vdd op_T3_jsr op_T3_jsr GND dfet w=10 l=19
+ ad=0 pd=0 as=927 ps=252 
M1206 Vdd op_T2_zp_zp_idx op_T2_zp_zp_idx GND dfet w=9 l=19
+ ad=0 pd=0 as=1888 ps=558 
M1207 n_913 n_913 Vdd GND dfet w=10 l=16
+ ad=575 pd=160 as=0 ps=0 
M1208 cp1 n_1105 GND GND efet w=198 l=7
+ ad=36125 pd=5694 as=0 ps=0 
M1209 GND n_1105 cp1 GND efet w=200 l=7
+ ad=0 pd=0 as=0 ps=0 
M1210 cp1 n_1105 GND GND efet w=198 l=8
+ ad=0 pd=0 as=0 ps=0 
M1211 GND n_1105 cp1 GND efet w=200 l=6
+ ad=0 pd=0 as=0 ps=0 
M1212 cp1 n_1105 GND GND efet w=198 l=8
+ ad=0 pd=0 as=0 ps=0 
M1213 Vdd n_1399 cp1 GND dfet w=68 l=7
+ ad=0 pd=0 as=0 ps=0 
M1214 n_1650 n_1650 Vdd GND dfet w=10 l=7
+ ad=285 pd=108 as=0 ps=0 
M1215 n_1105 n_1715 Vdd GND dfet w=24 l=6
+ ad=2597 pd=550 as=0 ps=0 
M1216 GND n_1399 n_1105 GND efet w=222 l=7
+ ad=0 pd=0 as=0 ps=0 
M1217 n_1399 n_1715 GND GND efet w=98 l=7
+ ad=2339 pd=520 as=0 ps=0 
M1218 GND n_1715 n_1399 GND efet w=185 l=6
+ ad=0 pd=0 as=0 ps=0 
M1219 GND n_358 n_1715 GND efet w=155 l=6
+ ad=0 pd=0 as=2655 ps=522 
M1220 Vdd n_1399 n_1399 GND dfet w=25 l=7
+ ad=0 pd=0 as=2893 ps=846 
M1221 Vdd n_1715 n_1715 GND dfet w=25 l=7
+ ad=0 pd=0 as=4571 ps=1442 
M1222 GND n_1467 cclk GND efet w=247 l=6
+ ad=0 pd=0 as=60259 ps=9520 
M1223 cclk n_1467 GND GND efet w=247 l=6
+ ad=0 pd=0 as=0 ps=0 
M1224 GND n_1467 cclk GND efet w=247 l=6
+ ad=0 pd=0 as=0 ps=0 
M1225 cclk n_1467 GND GND efet w=247 l=6
+ ad=0 pd=0 as=0 ps=0 
M1226 Vdd n_1129 cclk GND dfet w=68 l=8
+ ad=0 pd=0 as=0 ps=0 
M1227 n_1467 n_358 Vdd GND dfet w=25 l=6
+ ad=2780 pd=562 as=0 ps=0 
M1228 GND n_1129 n_1467 GND efet w=220 l=7
+ ad=0 pd=0 as=0 ps=0 
M1229 n_1129 n_358 GND GND efet w=39 l=6
+ ad=2724 pd=552 as=0 ps=0 
M1230 n_1129 cp1 GND GND efet w=112 l=6
+ ad=0 pd=0 as=0 ps=0 
M1231 GND n_358 n_1129 GND efet w=177 l=6
+ ad=0 pd=0 as=0 ps=0 
M1232 n_358 clk0 GND GND efet w=284 l=7
+ ad=2116 pd=412 as=0 ps=0 
M1233 n_358 n_358 Vdd GND dfet w=25 l=6
+ ad=4785 pd=1654 as=0 ps=0 
M1234 Vdd n_1129 n_1129 GND dfet w=25 l=7
+ ad=0 pd=0 as=4008 ps=1172 
M1235 rw n_102 Vdd GND efet w=139 l=7
+ ad=15066 pd=2234 as=0 ps=0 
M1236 Vdd n_102 rw GND efet w=139 l=6
+ ad=0 pd=0 as=0 ps=0 
M1237 GND GND clk0 GND efet w=47 l=8
+ ad=0 pd=0 as=0 ps=0 
M1238 rw n_102 Vdd GND efet w=138 l=6
+ ad=0 pd=0 as=0 ps=0 
M1239 Vdd n_102 rw GND efet w=138 l=7
+ ad=0 pd=0 as=0 ps=0 
M1240 rw n_102 Vdd GND efet w=138 l=7
+ ad=0 pd=0 as=0 ps=0 
M1241 Vdd n_102 rw GND efet w=138 l=7
+ ad=0 pd=0 as=0 ps=0 
M1242 rw n_102 Vdd GND efet w=155 l=6
+ ad=0 pd=0 as=0 ps=0 
M1243 n_633 cclk n_1059 GND efet w=10 l=16
+ ad=414 pd=98 as=1121 ps=240 
M1244 rw n_1696 GND GND efet w=151 l=7
+ ad=0 pd=0 as=0 ps=0 
M1245 GND n_1696 rw GND efet w=151 l=7
+ ad=0 pd=0 as=0 ps=0 
M1246 rw n_1696 GND GND efet w=151 l=6
+ ad=0 pd=0 as=0 ps=0 
M1247 GND n_1696 rw GND efet w=151 l=7
+ ad=0 pd=0 as=0 ps=0 
M1248 rw n_1696 GND GND efet w=213 l=6
+ ad=0 pd=0 as=0 ps=0 
M1249 GND n_400 n_102 GND efet w=123 l=8
+ ad=0 pd=0 as=1206 ps=302 
M1250 GND GND cclk GND efet w=55 l=6
+ ad=0 pd=0 as=0 ps=0 
M1251 Vdd op_T2_abs_access op_T2_abs_access GND dfet w=9 l=19
+ ad=0 pd=0 as=6070 ps=1986 
M1252 Vdd op_T2_branch op_T2_branch GND dfet w=9 l=18
+ ad=0 pd=0 as=1603 ps=504 
M1253 op_T2_ind op_T2_ind Vdd GND dfet w=10 l=19
+ ad=1216 pd=364 as=0 ps=0 
M1254 Vdd op_T4 op_T4 GND dfet w=9 l=19
+ ad=0 pd=0 as=895 ps=238 
M1255 op_T5_rts op_T5_rts Vdd GND dfet w=10 l=19
+ ad=6231 pd=2100 as=0 ps=0 
M1256 Vdd op_T0_brk_rti op_T0_brk_rti GND dfet w=9 l=19
+ ad=0 pd=0 as=997 ps=266 
M1257 Vdd op_T5_ind_x op_T5_ind_x GND dfet w=9 l=19
+ ad=0 pd=0 as=1127 ps=316 
M1258 Vdd op_T3 op_T3 GND dfet w=9 l=19
+ ad=0 pd=0 as=912 ps=252 
M1259 Vdd x_op_T3_abs_idx x_op_T3_abs_idx GND dfet w=9 l=19
+ ad=0 pd=0 as=869 ps=224 
M1260 Vdd op_T0_jmp op_T0_jmp GND dfet w=9 l=19
+ ad=0 pd=0 as=957 ps=276 
M1261 Vdd op_brk_rti op_brk_rti GND dfet w=9 l=19
+ ad=0 pd=0 as=827 ps=220 
M1262 Vdd x_op_jmp x_op_jmp GND dfet w=10 l=19
+ ad=0 pd=0 as=1180 ps=334 
M1263 Vdd diff_2598_3600# n_9 GND dfet w=10 l=19
+ ad=0 pd=0 as=258 ps=66 
M1264 Vdd op_T3_abs_idx_ind op_T3_abs_idx_ind GND dfet w=10 l=18
+ ad=0 pd=0 as=835 ps=252 
M1265 Vdd x_op_T4_ind_y x_op_T4_ind_y GND dfet w=9 l=19
+ ad=0 pd=0 as=1076 ps=324 
M1266 Vdd op_T3_branch op_T3_branch GND dfet w=9 l=18
+ ad=0 pd=0 as=1994 ps=644 
M1267 Vdd op_jsr op_jsr GND dfet w=9 l=19
+ ad=0 pd=0 as=745 ps=216 
M1268 Vdd op_push_pull op_push_pull GND dfet w=9 l=19
+ ad=0 pd=0 as=2361 ps=820 
M1269 Vdd op_T4_brk op_T4_brk GND dfet w=9 l=19
+ ad=0 pd=0 as=1642 ps=492 
M1270 Vdd op_T2_php_pha op_T2_php_pha GND dfet w=9 l=19
+ ad=0 pd=0 as=1520 ps=436 
M1271 Vdd n_173 n_173 GND dfet w=9 l=19
+ ad=0 pd=0 as=369 ps=82 
M1272 Vdd xx_op_T5_jsr xx_op_T5_jsr GND dfet w=9 l=18
+ ad=0 pd=0 as=753 ps=194 
M1273 Vdd op_T2_jmp_abs op_T2_jmp_abs GND dfet w=9 l=19
+ ad=0 pd=0 as=752 ps=194 
M1274 Vdd op_store op_store GND dfet w=10 l=19
+ ad=0 pd=0 as=978 ps=280 
M1275 Vdd op_T2_php op_T2_php GND dfet w=8 l=19
+ ad=0 pd=0 as=876 ps=242 
M1276 Vdd op_T4_jmp op_T4_jmp GND dfet w=10 l=19
+ ad=0 pd=0 as=2893 ps=950 
M1277 Vdd op_T5_rti_rts op_T5_rti_rts GND dfet w=9 l=19
+ ad=0 pd=0 as=827 ps=228 
M1278 Vdd op_lsr_ror_dec_inc op_lsr_ror_dec_inc GND dfet w=9 l=19
+ ad=0 pd=0 as=736 ps=190 
M1279 Vdd op_T0_cli_sei op_T0_cli_sei GND dfet w=9 l=19
+ ad=0 pd=0 as=696 ps=194 
M1280 Vdd op_T__bit op_T__bit GND dfet w=9 l=19
+ ad=0 pd=0 as=3287 ps=1068 
M1281 Vdd op_T3_mem_zp_idx op_T3_mem_zp_idx GND dfet w=10 l=19
+ ad=0 pd=0 as=926 ps=240 
M1282 n_834 n_402 GND GND efet w=71 l=7
+ ad=535 pd=170 as=0 ps=0 
M1283 n_102 n_834 Vdd GND dfet w=17 l=7
+ ad=0 pd=0 as=0 ps=0 
M1284 Vdd x_op_T0_bit x_op_T0_bit GND dfet w=9 l=19
+ ad=0 pd=0 as=1840 ps=574 
M1285 Vdd x_op_T3_plp_pla x_op_T3_plp_pla GND dfet w=9 l=19
+ ad=0 pd=0 as=781 ps=220 
M1286 GND _t5 op_T5_brk GND efet w=15 l=6
+ ad=0 pd=0 as=2366 ps=590 
M1287 GND _t5 op_T5_rti GND efet w=15 l=6
+ ad=0 pd=0 as=2064 ps=520 
M1288 GND _t5 op_T5_jsr GND efet w=14 l=7
+ ad=0 pd=0 as=2221 ps=572 
M1289 op_T2_abs_access op_push_pull GND GND efet w=14 l=6
+ ad=968 pd=238 as=0 ps=0 
M1290 op_T3_abs_idx_ind op_push_pull GND GND efet w=13 l=6
+ ad=1084 pd=262 as=0 ps=0 
M1291 Vdd op_asl_rol op_asl_rol GND dfet w=9 l=19
+ ad=0 pd=0 as=1439 ps=434 
M1292 Vdd n_1363 n_1363 GND dfet w=9 l=19
+ ad=0 pd=0 as=450 ps=110 
M1293 Vdd op_T0_clc_sec op_T0_clc_sec GND dfet w=9 l=19
+ ad=0 pd=0 as=1804 ps=554 
M1294 Vdd x_op_T__adc_sbc x_op_T__adc_sbc GND dfet w=10 l=19
+ ad=0 pd=0 as=3508 ps=1150 
M1295 Vdd x_op_T4_rti x_op_T4_rti GND dfet w=9 l=19
+ ad=0 pd=0 as=838 ps=216 
M1296 Vdd op_T0_plp op_T0_plp GND dfet w=9 l=19
+ ad=0 pd=0 as=803 ps=226 
M1297 Vdd op_T__cpx_cpy_abs op_T__cpx_cpy_abs GND dfet w=9 l=19
+ ad=0 pd=0 as=635 ps=176 
M1298 Vdd op_T__cmp op_T__cmp GND dfet w=10 l=19
+ ad=0 pd=0 as=736 ps=220 
M1299 Vdd op_T__cpx_cpy_imm_zp op_T__cpx_cpy_imm_zp GND dfet w=9 l=19
+ ad=0 pd=0 as=726 ps=202 
M1300 Vdd op_T0_cld_sed op_T0_cld_sed GND dfet w=9 l=19
+ ad=0 pd=0 as=729 ps=190 
M1301 Vdd op_T3_mem_abs op_T3_mem_abs GND dfet w=9 l=19
+ ad=0 pd=0 as=940 ps=236 
M1302 Vdd op_T5_mem_ind_idx op_T5_mem_ind_idx GND dfet w=9 l=18
+ ad=0 pd=0 as=945 ps=246 
M1303 Vdd op_T__asl_rol_a op_T__asl_rol_a GND dfet w=9 l=18
+ ad=0 pd=0 as=782 ps=242 
M1304 Vdd x_op_push_pull x_op_push_pull GND dfet w=10 l=20
+ ad=0 pd=0 as=1705 ps=578 
M1305 Vdd nop_branch_bit6 nop_branch_bit6 GND dfet w=10 l=20
+ ad=0 pd=0 as=5185 ps=1658 
M1306 Vdd op_T2_mem_zp op_T2_mem_zp GND dfet w=10 l=20
+ ad=0 pd=0 as=909 ps=276 
M1307 Vdd nop_branch_bit7 nop_branch_bit7 GND dfet w=10 l=15
+ ad=0 pd=0 as=5191 ps=1648 
M1308 Vdd op_implied op_implied GND dfet w=9 l=18
+ ad=0 pd=0 as=1471 ps=442 
M1309 Vdd op_T4_mem_abs_idx op_T4_mem_abs_idx GND dfet w=10 l=19
+ ad=0 pd=0 as=924 ps=250 
M1310 Vdd op_clv op_clv GND dfet w=10 l=19
+ ad=0 pd=0 as=2622 ps=810 
M1311 n_1696 n_400 Vdd GND dfet w=20 l=6
+ ad=1693 pd=376 as=0 ps=0 
M1312 GND n_834 n_1696 GND efet w=141 l=7
+ ad=0 pd=0 as=0 ps=0 
M1313 Vdd n_834 n_834 GND dfet w=10 l=12
+ ad=0 pd=0 as=2355 ps=680 
M1314 n_400 n_400 Vdd GND dfet w=10 l=10
+ ad=1700 pd=472 as=0 ps=0 
M1315 n_402 cp1 notRnWprepad GND efet w=13 l=7
+ ad=240 pd=76 as=2954 ps=702 
M1316 GND _t5 op_T5_ind_y GND efet w=14 l=7
+ ad=0 pd=0 as=1259 ps=322 
M1317 GND n_678 _t3 GND efet w=68 l=6
+ ad=0 pd=0 as=962 ps=280 
M1318 op_T4_rts _t4 GND GND efet w=14 l=6
+ ad=2337 pd=586 as=0 ps=0 
M1319 op_T4_brk_jsr _t4 GND GND efet w=14 l=6
+ ad=2135 pd=560 as=0 ps=0 
M1320 op_T4_rti _t4 GND GND efet w=14 l=6
+ ad=2064 pd=520 as=0 ps=0 
M1321 op_T4_ind_y _t4 GND GND efet w=14 l=6
+ ad=1264 pd=322 as=0 ps=0 
M1322 op_T4_ind_x _t4 GND GND efet w=15 l=6
+ ad=1638 pd=420 as=0 ps=0 
M1323 GND _t5 op_T5_rts GND efet w=14 l=6
+ ad=0 pd=0 as=2359 ps=620 
M1324 GND _t5 op_T5_ind_x GND efet w=14 l=6
+ ad=0 pd=0 as=1495 ps=382 
M1325 GND _t5 op_T5_rti_rts GND efet w=14 l=7
+ ad=0 pd=0 as=2095 ps=540 
M1326 GND _t5 xx_op_T5_jsr GND efet w=13 l=7
+ ad=0 pd=0 as=2207 ps=570 
M1327 op_T4_abs_idx _t4 GND GND efet w=14 l=6
+ ad=1113 pd=306 as=0 ps=0 
M1328 op_T4 _t4 GND GND efet w=14 l=6
+ ad=495 pd=128 as=0 ps=0 
M1329 x_op_T4_ind_y _t4 GND GND efet w=13 l=6
+ ad=1400 pd=372 as=0 ps=0 
M1330 GND _t5 op_T5_mem_ind_idx GND efet w=13 l=7
+ ad=0 pd=0 as=1232 ps=318 
M1331 GND x_op_push_pull op_implied GND efet w=21 l=7
+ ad=0 pd=0 as=1161 ps=276 
M1332 GND n_834 n_400 GND efet w=36 l=7
+ ad=0 pd=0 as=432 ps=146 
M1333 Vdd notir1 notir1 GND dfet w=10 l=7
+ ad=0 pd=0 as=20581 ps=6616 
M1334 GND ir1 n_1133 GND efet w=65 l=7
+ ad=0 pd=0 as=1183 ps=298 
M1335 n_119 cclk notir1 GND efet w=12 l=7
+ ad=560 pd=158 as=762 ps=208 
M1336 notir1 ir1 GND GND efet w=63 l=7
+ ad=0 pd=0 as=0 ps=0 
M1337 op_T4_brk _t4 GND GND efet w=14 l=6
+ ad=2285 pd=580 as=0 ps=0 
M1338 op_T4_jmp _t4 GND GND efet w=14 l=6
+ ad=2214 pd=568 as=0 ps=0 
M1339 x_op_T4_rti _t4 GND GND efet w=14 l=6
+ ad=1984 pd=508 as=0 ps=0 
M1340 n_1456 notRdy0 n_428 GND efet w=47 l=7
+ ad=0 pd=0 as=1266 ps=298 
M1341 pipeT3out cclk n_678 GND efet w=12 l=8
+ ad=225 pd=80 as=1614 ps=420 
M1342 _t3 _t3 Vdd GND dfet w=11 l=7
+ ad=18716 pd=5952 as=0 ps=0 
M1343 GND _t3 op_T3_ind_y GND efet w=14 l=6
+ ad=0 pd=0 as=1427 ps=376 
M1344 GND _t3 op_T3_plp_pla GND efet w=14 l=6
+ ad=0 pd=0 as=1999 ps=498 
M1345 op_T4_mem_abs_idx _t4 GND GND efet w=14 l=6
+ ad=1166 pd=306 as=0 ps=0 
M1346 n_428 n_16 n_1558 GND efet w=51 l=6
+ ad=0 pd=0 as=991 ps=278 
M1347 GND pipeT2out n_1558 GND efet w=110 l=6
+ ad=0 pd=0 as=0 ps=0 
M1348 Vdd n_428 n_428 GND dfet w=9 l=16
+ ad=0 pd=0 as=306 ps=84 
M1349 Vdd n_678 n_678 GND dfet w=10 l=12
+ ad=0 pd=0 as=1112 ps=352 
M1350 GND n_1357 n_678 GND efet w=32 l=7
+ ad=0 pd=0 as=0 ps=0 
M1351 GND _t3 op_T3_stack_bit_jmp GND efet w=14 l=6
+ ad=0 pd=0 as=1276 ps=324 
M1352 GND _t3 op_T3_ind_x GND efet w=14 l=6
+ ad=0 pd=0 as=1643 ps=436 
M1353 GND _t3 op_T3_abs_idx GND efet w=13 l=6
+ ad=0 pd=0 as=1013 ps=258 
M1354 op_T2_abs_y _t2 GND GND efet w=14 l=6
+ ad=1296 pd=328 as=0 ps=0 
M1355 op_T2_idx_x_xy _t2 GND GND efet w=14 l=6
+ ad=1181 pd=310 as=0 ps=0 
M1356 op_T2_ind_x _t2 GND GND efet w=15 l=6
+ ad=1702 pd=440 as=0 ps=0 
M1357 op_T2 _t2 GND GND efet w=16 l=6
+ ad=539 pd=134 as=0 ps=0 
M1358 GND _t3 x_op_T3_ind_y GND efet w=15 l=7
+ ad=0 pd=0 as=1335 ps=332 
M1359 GND _t3 op_T3_jmp GND efet w=14 l=7
+ ad=0 pd=0 as=2033 ps=518 
M1360 GND _t3 op_T3_jsr GND efet w=14 l=6
+ ad=0 pd=0 as=2433 ps=630 
M1361 op_T2_abs _t2 GND GND efet w=15 l=6
+ ad=1420 pd=376 as=0 ps=0 
M1362 op_T2_ADL_ADD _t2 GND GND efet w=15 l=6
+ ad=901 pd=244 as=0 ps=0 
M1363 op_T2_stack _t2 GND GND efet w=15 l=6
+ ad=1686 pd=436 as=0 ps=0 
M1364 op_T2_ind_y _t2 GND GND efet w=15 l=6
+ ad=1462 pd=366 as=0 ps=0 
M1365 GND _t3 op_T3 GND efet w=15 l=6
+ ad=0 pd=0 as=663 ps=168 
M1366 GND _t3 op_T3_abs_idx_ind GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1367 GND _t3 x_op_T3_abs_idx GND efet w=14 l=6
+ ad=0 pd=0 as=1074 ps=266 
M1368 GND _t3 op_T3_branch GND efet w=14 l=6
+ ad=0 pd=0 as=1421 ps=378 
M1369 n_1133 n_1133 Vdd GND dfet w=9 l=8
+ ad=1000 pd=306 as=0 ps=0 
M1370 n_678 n_644 GND GND efet w=61 l=6
+ ad=0 pd=0 as=0 ps=0 
M1371 n_644 cp1 n_428 GND efet w=13 l=9
+ ad=247 pd=102 as=0 ps=0 
M1372 GND n_1575 _t2 GND efet w=76 l=6
+ ad=0 pd=0 as=920 ps=228 
M1373 GND pipeT2out n_12 GND efet w=124 l=7
+ ad=0 pd=0 as=586 ps=222 
M1374 n_1575 cclk pipeT2out GND efet w=12 l=8
+ ad=1062 pd=300 as=320 ps=92 
M1375 _t2 _t2 Vdd GND dfet w=10 l=7
+ ad=18572 pd=6192 as=0 ps=0 
M1376 op_T2_jsr _t2 GND GND efet w=13 l=6
+ ad=2237 pd=574 as=0 ps=0 
M1377 op_T2_stack_access _t2 GND GND efet w=14 l=6
+ ad=1631 pd=436 as=0 ps=0 
M1378 op_T2_pha _t2 GND GND efet w=14 l=6
+ ad=1967 pd=516 as=0 ps=0 
M1379 op_T2_brk _t2 GND GND efet w=14 l=6
+ ad=2199 pd=568 as=0 ps=0 
M1380 op_T2_branch _t2 GND GND efet w=14 l=6
+ ad=1398 pd=356 as=0 ps=0 
M1381 op_T2_zp_zp_idx _t2 GND GND efet w=14 l=6
+ ad=998 pd=256 as=0 ps=0 
M1382 GND _t3 x_op_T3_plp_pla GND efet w=15 l=6
+ ad=0 pd=0 as=1914 ps=502 
M1383 GND _t3 op_T3_mem_zp_idx GND efet w=15 l=6
+ ad=0 pd=0 as=1074 ps=268 
M1384 op_T2_ind _t2 GND GND efet w=14 l=6
+ ad=1260 pd=322 as=0 ps=0 
M1385 op_T2_abs_access _t2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1386 GND _t3 op_T3_mem_abs GND efet w=14 l=7
+ ad=0 pd=0 as=1294 ps=326 
M1387 GND ir0 op_implied GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1388 GND n_1133 irline3 GND efet w=84 l=7
+ ad=0 pd=0 as=892 ps=238 
M1389 n_1133 ir0 GND GND efet w=70 l=5
+ ad=0 pd=0 as=0 ps=0 
M1390 ir1 ir1 Vdd GND dfet w=11 l=12
+ ad=1631 pd=456 as=0 ps=0 
M1391 GND n_119 ir1 GND efet w=77 l=7
+ ad=0 pd=0 as=798 ps=244 
M1392 n_237 fetch n_119 GND efet w=22 l=8
+ ad=110 pd=54 as=0 ps=0 
M1393 n_1641 cp1 n_237 GND efet w=22 l=7
+ ad=1074 pd=302 as=0 ps=0 
M1394 op_T2_php _t2 GND GND efet w=14 l=6
+ ad=2193 pd=556 as=0 ps=0 
M1395 op_T2_php_pha _t2 GND GND efet w=14 l=6
+ ad=1780 pd=452 as=0 ps=0 
M1396 op_T2_jmp_abs _t2 GND GND efet w=14 l=6
+ ad=2104 pd=524 as=0 ps=0 
M1397 op_T2_mem_zp _t2 GND GND efet w=15 l=6
+ ad=1379 pd=368 as=0 ps=0 
M1398 ir0 ir0 Vdd GND dfet w=10 l=11
+ ad=2975 pd=944 as=0 ps=0 
M1399 ir0 n_310 GND GND efet w=70 l=8
+ ad=988 pd=224 as=0 ps=0 
M1400 GND notir1 op_xy GND efet w=14 l=6
+ ad=0 pd=0 as=1024 ps=260 
M1401 GND notir1 x_op_T0_txa GND efet w=14 l=6
+ ad=0 pd=0 as=1879 ps=464 
M1402 GND notir1 op_T0_dex GND efet w=14 l=6
+ ad=0 pd=0 as=1753 ps=452 
M1403 GND notir1 op_from_x GND efet w=14 l=6
+ ad=0 pd=0 as=1323 ps=360 
M1404 GND notir1 op_T0_txs GND efet w=15 l=6
+ ad=0 pd=0 as=2104 ps=530 
M1405 irline3 irline3 Vdd GND dfet w=13 l=6
+ ad=18753 pd=6276 as=0 ps=0 
M1406 n_724 fetch n_310 GND efet w=23 l=8
+ ad=115 pd=56 as=516 ps=152 
M1407 n_409 cp1 n_724 GND efet w=23 l=7
+ ad=1226 pd=274 as=0 ps=0 
M1408 GND ir0 notir0 GND efet w=66 l=7
+ ad=0 pd=0 as=956 ps=258 
M1409 GND notir1 op_T0_ldx_tax_tsx GND efet w=14 l=6
+ ad=0 pd=0 as=1418 ps=374 
M1410 GND notir1 op_T__dex GND efet w=15 l=6
+ ad=0 pd=0 as=1632 ps=420 
M1411 GND notir1 op_T0_tsx GND efet w=16 l=6
+ ad=0 pd=0 as=1888 ps=466 
M1412 GND notir1 op_ror GND efet w=14 l=6
+ ad=0 pd=0 as=1447 ps=378 
M1413 op_sty_cpy_mem irline3 GND GND efet w=14 l=6
+ ad=1306 pd=328 as=0 ps=0 
M1414 op_T0_iny_dey irline3 GND GND efet w=14 l=6
+ ad=1707 pd=440 as=0 ps=0 
M1415 x_op_T0_tya irline3 GND GND efet w=14 l=6
+ ad=2146 pd=530 as=0 ps=0 
M1416 op_T0_cpy_iny irline3 GND GND efet w=14 l=6
+ ad=1486 pd=380 as=0 ps=0 
M1417 op_T0_cpx_inx irline3 GND GND efet w=14 l=6
+ ad=1393 pd=340 as=0 ps=0 
M1418 GND notir1 op_inc_nop GND efet w=14 l=7
+ ad=0 pd=0 as=1260 ps=320 
M1419 GND notir1 op_rol_ror GND efet w=13 l=6
+ ad=0 pd=0 as=1329 ps=350 
M1420 GND notir1 op_shift GND efet w=15 l=6
+ ad=0 pd=0 as=1141 ps=304 
M1421 GND notir1 op_T__shift_a GND efet w=14 l=6
+ ad=0 pd=0 as=1726 ps=454 
M1422 GND notir1 op_T0_txa GND efet w=14 l=6
+ ad=0 pd=0 as=1830 ps=460 
M1423 op_T__inx irline3 GND GND efet w=15 l=6
+ ad=1993 pd=520 as=0 ps=0 
M1424 op_T__iny_dey irline3 GND GND efet w=14 l=6
+ ad=1816 pd=472 as=0 ps=0 
M1425 op_T0_ldy_mem irline3 GND GND efet w=13 l=6
+ ad=1342 pd=334 as=0 ps=0 
M1426 op_T0_tay_ldy_not_idx irline3 GND GND efet w=14 l=6
+ ad=1483 pd=384 as=0 ps=0 
M1427 op_T0_jsr irline3 GND GND efet w=14 l=6
+ ad=2271 pd=578 as=0 ps=0 
M1428 op_T5_brk irline3 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1429 op_T0_php_pha irline3 GND GND efet w=15 l=6
+ ad=2003 pd=512 as=0 ps=0 
M1430 op_T4_rts irline3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1431 op_T3_plp_pla irline3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1432 op_T5_rti irline3 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1433 op_jmp irline3 GND GND efet w=14 l=6
+ ad=1862 pd=462 as=0 ps=0 
M1434 op_T2_stack irline3 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1435 op_T3_stack_bit_jmp irline3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1436 op_T4_brk_jsr irline3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1437 op_T4_rti irline3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1438 op_plp_pla irline3 GND GND efet w=14 l=6
+ ad=1642 pd=432 as=0 ps=0 
M1439 GND notir1 op_T0_shift_a GND efet w=14 l=6
+ ad=0 pd=0 as=1714 ps=446 
M1440 GND notir1 op_T0_tax GND efet w=14 l=6
+ ad=0 pd=0 as=1548 ps=392 
M1441 GND notir1 op_T0_shift_right_a GND efet w=14 l=6
+ ad=0 pd=0 as=1819 ps=458 
M1442 GND notir1 op_shift_right GND efet w=14 l=6
+ ad=0 pd=0 as=1194 ps=316 
M1443 op_rti_rts irline3 GND GND efet w=14 l=6
+ ad=1925 pd=502 as=0 ps=0 
M1444 op_T2_jsr irline3 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1445 op_T0_cpx_cpy_inx_iny irline3 GND GND efet w=14 l=6
+ ad=1438 pd=380 as=0 ps=0 
M1446 op_T3_jmp irline3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1447 op_T5_jsr irline3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1448 op_T2_stack_access irline3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1449 op_T0_tya irline3 GND GND efet w=14 l=6
+ ad=2038 pd=518 as=0 ps=0 
M1450 op_T0_pla irline3 GND GND efet w=15 l=6
+ ad=1975 pd=512 as=0 ps=0 
M1451 GND notir1 op_lsr_ror_dec_inc GND efet w=14 l=7
+ ad=0 pd=0 as=732 ps=190 
M1452 GND notir1 op_asl_rol GND efet w=14 l=7
+ ad=0 pd=0 as=1113 ps=304 
M1453 GND notir1 op_T__asl_rol_a GND efet w=14 l=6
+ ad=0 pd=0 as=1915 ps=506 
M1454 op_T0_tay irline3 GND GND efet w=14 l=6
+ ad=1541 pd=392 as=0 ps=0 
M1455 op_T0_bit irline3 GND GND efet w=14 l=6
+ ad=1711 pd=448 as=0 ps=0 
M1456 op_branch_done irline3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1457 op_T2_pha irline3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1458 op_T2_brk irline3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1459 op_T3_jsr irline3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1460 op_T2_branch irline3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1461 op_T5_rts irline3 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1462 op_T0_brk_rti irline3 GND GND efet w=14 l=6
+ ad=1912 pd=502 as=0 ps=0 
M1463 op_T0_jmp irline3 GND GND efet w=14 l=6
+ ad=2200 pd=572 as=0 ps=0 
M1464 op_T3_branch irline3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1465 op_brk_rti irline3 GND GND efet w=15 l=6
+ ad=1773 pd=450 as=0 ps=0 
M1466 op_jsr irline3 GND GND efet w=15 l=6
+ ad=2139 pd=562 as=0 ps=0 
M1467 x_op_jmp irline3 GND GND efet w=14 l=6
+ ad=1816 pd=456 as=0 ps=0 
M1468 op_push_pull irline3 GND GND efet w=14 l=6
+ ad=1392 pd=356 as=0 ps=0 
M1469 notir0 notir0 Vdd GND dfet w=10 l=7
+ ad=20026 pd=6376 as=0 ps=0 
M1470 op_T4_brk irline3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1471 op_T2_php irline3 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1472 op_T2_php_pha irline3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1473 op_T4_jmp irline3 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1474 op_T5_rti_rts irline3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1475 xx_op_T5_jsr irline3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1476 op_T2_jmp_abs irline3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1477 x_op_T3_plp_pla irline3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1478 op_T0_cli_sei irline3 GND GND efet w=14 l=6
+ ad=1768 pd=450 as=0 ps=0 
M1479 op_T__bit irline3 GND GND efet w=14 l=6
+ ad=1959 pd=532 as=0 ps=0 
M1480 op_T0_clc_sec irline3 GND GND efet w=14 l=6
+ ad=1899 pd=498 as=0 ps=0 
M1481 x_op_T0_bit irline3 GND GND efet w=14 l=6
+ ad=1551 pd=390 as=0 ps=0 
M1482 op_T0_plp irline3 GND GND efet w=13 l=6
+ ad=1904 pd=506 as=0 ps=0 
M1483 x_op_T4_rti irline3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1484 op_T__cpx_cpy_abs irline3 GND GND efet w=15 l=6
+ ad=1859 pd=486 as=0 ps=0 
M1485 op_T__cpx_cpy_imm_zp irline3 GND GND efet w=15 l=6
+ ad=1657 pd=424 as=0 ps=0 
M1486 GND notir0 op_T3_ind_y GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1487 GND notir0 op_T2_abs_y GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1488 n_1575 n_1575 Vdd GND dfet w=10 l=12
+ ad=1142 pd=376 as=0 ps=0 
M1489 GND notir0 op_T2_ind_x GND efet w=15 l=7
+ ad=0 pd=0 as=0 ps=0 
M1490 x_op_push_pull irline3 GND GND efet w=14 l=6
+ ad=1409 pd=364 as=0 ps=0 
M1491 op_T0_cld_sed irline3 GND GND efet w=14 l=6
+ ad=1815 pd=456 as=0 ps=0 
M1492 op_clv irline3 GND GND efet w=13 l=6
+ ad=1946 pd=486 as=0 ps=0 
M1493 n_310 cclk notir0 GND efet w=13 l=7
+ ad=0 pd=0 as=0 ps=0 
M1494 GND notir0 op_T0_eor GND efet w=15 l=6
+ ad=0 pd=0 as=1250 ps=320 
M1495 GND notir0 op_T0_ora GND efet w=14 l=6
+ ad=0 pd=0 as=1315 ps=330 
M1496 GND notir0 op_T3_ind_x GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1497 GND notir0 op_T4_ind_y GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1498 GND notir0 op_T2_ind_y GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1499 GND notir0 op_T4_ind_x GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1500 GND n_1357 n_1575 GND efet w=47 l=7
+ ad=0 pd=0 as=0 ps=0 
M1501 op_T0_jsr ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1502 op_T5_brk ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1503 op_T0_php_pha ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1504 op_T4_rts ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1505 op_T3_plp_pla ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1506 op_T5_rti ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1507 op_ror ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1508 GND notir0 x_op_T3_ind_y GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1509 GND notir0 op_T0_cmp GND efet w=14 l=7
+ ad=0 pd=0 as=1322 ps=330 
M1510 GND notir0 op_T0_sbc GND efet w=14 l=7
+ ad=0 pd=0 as=1410 ps=374 
M1511 GND notir0 op_T0_adc_sbc GND efet w=14 l=7
+ ad=0 pd=0 as=1088 ps=268 
M1512 GND notir0 op_T__ora_and_eor_adc GND efet w=14 l=7
+ ad=0 pd=0 as=943 ps=272 
M1513 GND notir0 op_T__adc_sbc GND efet w=14 l=7
+ ad=0 pd=0 as=1278 ps=334 
M1514 GND notir0 op_T0_lda GND efet w=15 l=6
+ ad=0 pd=0 as=1264 ps=322 
M1515 GND notir0 op_T0_acc GND efet w=13 l=6
+ ad=0 pd=0 as=895 ps=248 
M1516 GND notir0 op_T0_and GND efet w=14 l=6
+ ad=0 pd=0 as=1034 ps=262 
M1517 GND notir0 op_T5_ind_y GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1518 GND notir0 op_sta_cmp GND efet w=13 l=6
+ ad=0 pd=0 as=1265 ps=322 
M1519 n_12 notRdy0 n_1091 GND efet w=51 l=8
+ ad=0 pd=0 as=1086 ps=244 
M1520 op_T0_eor ir7 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1521 op_jmp ir7 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1522 op_T0_ora ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1523 op_T2_stack ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1524 op_T3_stack_bit_jmp ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1525 op_T4_brk_jsr ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1526 op_T4_rti ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1527 op_plp_pla ir7 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1528 op_rti_rts ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1529 op_T2_jsr ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1530 op_rol_ror ir7 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1531 op_T3_jmp ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1532 op_shift ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1533 op_T5_jsr ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1534 op_T2_stack_access ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1535 op_T__ora_and_eor_adc ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1536 op_T__shift_a ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1537 op_T0_pla ir7 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1538 GND notir0 op_T2_ind GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1539 GND notir0 op_T5_ind_x GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1540 GND notir0 x_op_T4_ind_y GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1541 op_T0_shift_a ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1542 op_T0_bit ir7 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1543 op_T0_and ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1544 op_T2_pha ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1545 op_T0_shift_right_a ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1546 op_shift_right ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1547 op_T2_brk ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1548 op_T3_jsr ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1549 GND notir0 x_op_T__adc_sbc GND efet w=15 l=7
+ ad=0 pd=0 as=2220 ps=590 
M1550 GND notir0 op_T__cmp GND efet w=13 l=7
+ ad=0 pd=0 as=1432 ps=386 
M1551 GND notir0 op_T5_mem_ind_idx GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1552 n_1575 n_1360 GND GND efet w=73 l=7
+ ad=0 pd=0 as=0 ps=0 
M1553 n_1091 n_16 n_363 GND efet w=51 l=6
+ ad=0 pd=0 as=989 ps=256 
M1554 n_1360 cp1 n_1091 GND efet w=12 l=7
+ ad=167 pd=74 as=0 ps=0 
M1555 GND notir7 op_sty_cpy_mem GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1556 GND notir7 op_T0_iny_dey GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1557 GND notir7 x_op_T0_tya GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1558 GND notir7 op_T0_cpy_iny GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1559 GND notir7 op_xy GND efet w=15 l=7
+ ad=0 pd=0 as=0 ps=0 
M1560 GND notir7 x_op_T0_txa GND efet w=15 l=7
+ ad=0 pd=0 as=0 ps=0 
M1561 GND notir7 op_T0_dex GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1562 GND notir7 op_T0_cpx_inx GND efet w=15 l=7
+ ad=0 pd=0 as=0 ps=0 
M1563 GND notir7 op_from_x GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1564 GND notir7 op_T0_txs GND efet w=16 l=6
+ ad=0 pd=0 as=0 ps=0 
M1565 op_T5_rts ir7 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1566 op_T0_brk_rti ir7 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1567 op_T0_jmp ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1568 op_brk_rti ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1569 op_jsr ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1570 x_op_jmp ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1571 op_push_pull ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1572 op_T4_brk ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1573 op_T2_php ir7 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1574 op_T2_php_pha ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1575 op_T4_jmp ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1576 op_T5_rti_rts ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1577 xx_op_T5_jsr ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1578 op_T2_jmp_abs ir7 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1579 x_op_T3_plp_pla ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1580 op_asl_rol ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1581 op_T0_cli_sei ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1582 op_T__bit ir7 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1583 op_T0_clc_sec ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1584 ir7 ir7 Vdd GND dfet w=10 l=6
+ ad=19941 pd=6644 as=0 ps=0 
M1585 GND n_541 ir7 GND efet w=121 l=6
+ ad=0 pd=0 as=1252 ps=296 
M1586 notir7 notir7 Vdd GND dfet w=10 l=7
+ ad=19293 pd=6134 as=0 ps=0 
M1587 GND ir7 notir7 GND efet w=89 l=6
+ ad=0 pd=0 as=1797 ps=404 
M1588 n_1183 fetch n_541 GND efet w=22 l=8
+ ad=110 pd=54 as=468 ps=112 
M1589 n_1605 cp1 n_1183 GND efet w=22 l=8
+ ad=1228 pd=270 as=0 ps=0 
M1590 n_541 cclk notir7 GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M1591 GND notir7 op_T0_ldx_tax_tsx GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1592 GND notir7 op_T__dex GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1593 GND notir7 op_T__inx GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1594 GND notir7 op_T0_tsx GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1595 GND notir7 op_T__iny_dey GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1596 GND notir7 op_T0_ldy_mem GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1597 GND notir7 op_T0_tay_ldy_not_idx GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1598 x_op_T0_bit ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1599 op_T0_plp ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1600 x_op_T4_rti ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1601 op_T__asl_rol_a ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1602 x_op_push_pull ir7 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1603 nop_branch_bit7 ir7 GND GND efet w=31 l=6
+ ad=663 pd=166 as=0 ps=0 
M1604 GND pipeT_SYNC n_363 GND efet w=120 l=6
+ ad=0 pd=0 as=0 ps=0 
M1605 Vdd n_1091 n_1091 GND dfet w=10 l=16
+ ad=0 pd=0 as=326 ps=84 
M1606 op_T0_iny_dey ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1607 op_T0_cpy_iny ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1608 op_T2_ind_x ir4 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1609 x_op_T0_txa ir4 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1610 op_T0_dex ir4 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1611 op_T0_cpx_inx ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1612 GND notir7 op_inc_nop GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1613 op_T__dex ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1614 op_T__inx ir4 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1615 op_T__iny_dey ir4 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1616 op_T0_tay_ldy_not_idx ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1617 op_T0_jsr ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1618 op_T5_brk ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1619 op_T0_php_pha ir4 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1620 op_T4_rts ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1621 op_T3_plp_pla ir4 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1622 op_T5_rti ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1623 op_jmp ir4 GND GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1624 op_T2_abs ir4 GND GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1625 op_T2_stack ir4 GND GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1626 op_T3_stack_bit_jmp ir4 GND GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1627 GND notir7 op_T0_cpx_cpy_inx_iny GND efet w=15 l=7
+ ad=0 pd=0 as=0 ps=0 
M1628 GND notir7 op_T0_cmp GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1629 GND notir7 op_T0_sbc GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1630 GND notir7 op_T0_tya GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1631 GND notir7 op_T0_txa GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1632 GND notir7 op_T0_lda GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1633 GND notir7 op_T0_tay GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1634 GND notir7 op_T0_tax GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1635 GND notir7 op_sta_cmp GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1636 op_T4_brk_jsr ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1637 op_T4_rti ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1638 op_T3_ind_x ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1639 op_plp_pla ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1640 op_T4_ind_x ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1641 op_rti_rts ir4 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1642 op_T2_jsr ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1643 op_T0_cpx_cpy_inx_iny ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1644 op_T3_jmp ir4 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1645 op_T5_jsr ir4 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1646 op_T2_stack_access ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1647 op_T__shift_a ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1648 op_T0_txa ir4 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1649 op_T0_pla ir4 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1650 GND notir7 op_store GND efet w=14 l=6
+ ad=0 pd=0 as=1070 ps=286 
M1651 n_862 cclk pipeT_SYNC GND efet w=12 l=7
+ ad=1833 pd=530 as=190 ps=76 
M1652 op_T0_tay ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1653 op_T0_shift_a ir4 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1654 op_T0_tax ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1655 op_T0_bit ir4 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1656 op_T2_pha ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1657 op_T0_shift_right_a ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1658 op_T2_brk ir4 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1659 op_T3_jsr ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1660 GND notir7 op_T__cmp GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1661 GND notir7 op_T__cpx_cpy_abs GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1662 GND notir7 op_T__cpx_cpy_imm_zp GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1663 GND notir7 op_T0_cld_sed GND efet w=15 l=7
+ ad=0 pd=0 as=0 ps=0 
M1664 GND notir7 op_clv GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1665 op_T5_rts ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1666 op_T0_brk_rti ir4 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1667 op_T0_jmp ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1668 op_T5_ind_x ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1669 op_brk_rti ir4 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1670 op_jsr ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1671 x_op_jmp ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1672 op_push_pull ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1673 op_T4_brk ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1674 op_T2_php ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1675 op_T2_php_pha ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1676 op_T4_jmp ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1677 op_T5_rti_rts ir4 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1678 xx_op_T5_jsr ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1679 op_T2_jmp_abs ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1680 x_op_T3_plp_pla ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1681 op_T__bit ir4 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1682 ir4 ir4 Vdd GND dfet w=10 l=7
+ ad=20206 pd=6646 as=0 ps=0 
M1683 GND n_927 ir4 GND efet w=122 l=6
+ ad=0 pd=0 as=1109 ps=284 
M1684 x_op_T0_bit ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1685 op_T0_plp ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1686 x_op_T4_rti ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1687 op_T__cpx_cpy_abs ir4 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1688 op_T__asl_rol_a ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1689 op_T__cpx_cpy_imm_zp ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1690 x_op_push_pull ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1691 op_T3_mem_abs ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1692 op_T2_mem_zp ir4 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1693 notir4 notir4 Vdd GND dfet w=10 l=6
+ ad=18955 pd=6044 as=0 ps=0 
M1694 GND ir4 notir4 GND efet w=86 l=6
+ ad=0 pd=0 as=1994 ps=414 
M1695 n_703 fetch n_927 GND efet w=24 l=8
+ ad=120 pd=58 as=458 ps=108 
M1696 n_227 cp1 n_703 GND efet w=24 l=8
+ ad=1294 pd=288 as=0 ps=0 
M1697 GND notir4 op_T3_ind_y GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1698 GND notir4 op_T2_abs_y GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1699 GND notir4 x_op_T0_tya GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1700 GND notir4 op_T2_idx_x_xy GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1701 GND notir4 op_T0_txs GND efet w=16 l=6
+ ad=0 pd=0 as=0 ps=0 
M1702 n_927 cclk notir4 GND efet w=12 l=7
+ ad=0 pd=0 as=0 ps=0 
M1703 n_1368 NMIL GND GND efet w=51 l=6
+ ad=1754 pd=486 as=0 ps=0 
M1704 GND n_562 NMIL GND efet w=66 l=6
+ ad=0 pd=0 as=1147 ps=322 
M1705 NMIL NMIL Vdd GND dfet w=10 l=14
+ ad=1405 pd=430 as=0 ps=0 
M1706 GND notRdy0 n_16 GND efet w=55 l=6
+ ad=0 pd=0 as=779 ps=168 
M1707 Vdd n_16 n_16 GND dfet w=10 l=10
+ ad=0 pd=0 as=2630 ps=820 
M1708 NMIL n_882 GND GND efet w=35 l=7
+ ad=0 pd=0 as=0 ps=0 
M1709 n_562 cp1 n_645 GND efet w=12 l=9
+ ad=256 pd=90 as=0 ps=0 
M1710 GND n_645 n_1368 GND efet w=36 l=7
+ ad=0 pd=0 as=0 ps=0 
M1711 n_1368 n_1578 GND GND efet w=44 l=7
+ ad=0 pd=0 as=0 ps=0 
M1712 Vdd n_1368 n_1368 GND dfet w=10 l=10
+ ad=0 pd=0 as=2455 ps=818 
M1713 NMIL cclk n_1252 GND efet w=13 l=7
+ ad=0 pd=0 as=342 ps=94 
M1714 n_1578 pipenVEC GND GND efet w=60 l=8
+ ad=519 pd=128 as=0 ps=0 
M1715 Vdd n_1578 n_1578 GND dfet w=11 l=17
+ ad=0 pd=0 as=798 ps=210 
M1716 n_882 n_1252 GND GND efet w=54 l=7
+ ad=1001 pd=284 as=0 ps=0 
M1717 GND notir4 op_T0_tsx GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1718 GND notir4 op_T4_ind_y GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1719 GND notir4 op_T2_ind_y GND efet w=15 l=7
+ ad=0 pd=0 as=0 ps=0 
M1720 GND notir4 op_T3_abs_idx GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1721 GND notir4 x_op_T3_ind_y GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1722 GND notir4 op_T0_tya GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1723 op_T3_ind_y ir3 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1724 op_T2_ind_x ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1725 op_T0_jsr ir3 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1726 op_T5_brk ir3 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1727 op_T4_rts ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1728 op_T5_rti ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1729 op_T2_ADL_ADD ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1730 op_T4_brk_jsr ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1731 op_T4_rti ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1732 op_T3_ind_x ir3 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1733 op_T4_ind_y ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1734 op_T2_ind_y ir3 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1735 op_T4_ind_x ir3 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1736 GND notir4 op_T4_abs_idx GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1737 GND notir4 op_T5_ind_y GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1738 GND notir4 op_branch_done GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1739 GND notir4 op_T2_branch GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1740 GND notir4 x_op_T4_ind_y GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1741 GND notir4 x_op_T3_abs_idx GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1742 GND notir4 op_T3_branch GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1743 x_op_T3_ind_y ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1744 op_rti_rts ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1745 op_T2_jsr ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1746 op_T5_jsr ir3 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1747 op_T5_ind_y ir3 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1748 op_branch_done ir3 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1749 op_T2_brk ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1750 op_T3_jsr ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1751 op_T2_branch ir3 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1752 op_T2_zp_zp_idx ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1753 GND notir4 op_T0_cli_sei GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1754 GND notir4 op_T0_clc_sec GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1755 GND notir4 op_T3_mem_zp_idx GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1756 GND notir4 op_T0_cld_sed GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1757 GND notir3 op_T2_abs_y GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1758 GND notir3 op_T0_iny_dey GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1759 GND notir3 x_op_T0_tya GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1760 GND notir3 x_op_T0_txa GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1761 GND notir3 op_T0_dex GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1762 GND notir3 op_T0_txs GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1763 op_T2_ind ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1764 op_T5_rts ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1765 op_T0_brk_rti ir3 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1766 op_T5_ind_x ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1767 x_op_T4_ind_y ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1768 op_T3_branch ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1769 op_brk_rti ir3 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1770 op_jsr ir3 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1771 GND notir4 op_T4_mem_abs_idx GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1772 GND notir4 op_clv GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1773 ir3 ir3 Vdd GND dfet w=9 l=7
+ ad=19949 pd=6530 as=0 ps=0 
M1774 op_T4_brk ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1775 op_T5_rti_rts ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1776 xx_op_T5_jsr ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1777 op_T3_mem_zp_idx ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1778 x_op_T4_rti ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1779 op_T__cpx_cpy_imm_zp ir3 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1780 op_T2_mem_zp ir3 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1781 op_T5_mem_ind_idx ir3 GND GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1782 GND n_1620 ir3 GND efet w=128 l=7
+ ad=0 pd=0 as=1297 ps=302 
M1783 GND notir3 op_T__dex GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1784 GND notir3 op_T__inx GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1785 GND notir3 op_T0_tsx GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1786 GND notir3 op_T__iny_dey GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1787 GND notir3 op_T0_php_pha GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1788 GND notir3 op_T3_plp_pla GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1789 GND notir3 op_jmp GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1790 GND notir3 op_T2_abs GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1791 GND notir3 op_T3_abs_idx GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1792 GND notir3 op_plp_pla GND efet w=13 l=7
+ ad=0 pd=0 as=0 ps=0 
M1793 GND notir3 op_T3_jmp GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1794 GND notir3 op_T0_tya GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1795 GND notir3 op_T__shift_a GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1796 GND notir3 op_T0_txa GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1797 GND notir3 op_T0_pla GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1798 op_T3_ind_y ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1799 op_T2_abs_y ir2 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1800 op_T0_iny_dey ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1801 x_op_T0_tya ir2 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1802 op_T2_ind_x ir2 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1803 x_op_T0_txa ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1804 op_T0_dex ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1805 op_T0_txs ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1806 op_T__dex ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1807 op_T__inx ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1808 op_T0_tsx ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1809 op_T__iny_dey ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1810 op_T0_jsr ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1811 op_T5_brk ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1812 op_T0_php_pha ir2 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1813 op_T4_rts ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1814 op_T3_plp_pla ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1815 op_T5_rti ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1816 GND n_597 n_882 GND efet w=71 l=7
+ ad=0 pd=0 as=0 ps=0 
M1817 n_882 n_882 Vdd GND dfet w=9 l=17
+ ad=895 pd=250 as=0 ps=0 
M1818 op_T2_stack ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1819 op_T4_brk_jsr ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1820 op_T4_rti ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1821 op_T3_ind_x ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1822 op_T4_ind_y ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1823 op_T2_ind_y ir2 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1824 op_plp_pla ir2 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1825 op_T4_ind_x ir2 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1826 GND notir3 op_T0_tay GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1827 GND notir3 op_T0_shift_a GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1828 GND notir3 op_T0_tax GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1829 GND notir3 op_T4_abs_idx GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1830 GND notir3 op_T2_pha GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1831 GND notir3 op_T0_shift_right_a GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1832 notir3 notir3 Vdd GND dfet w=9 l=7
+ ad=18731 pd=6008 as=0 ps=0 
M1833 GND ir3 notir3 GND efet w=85 l=7
+ ad=0 pd=0 as=1805 ps=402 
M1834 GND notir3 op_T2_abs_access GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1835 GND notir3 op_T0_jmp GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1836 GND notir3 op_T3_abs_idx_ind GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1837 GND notir3 x_op_T3_abs_idx GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1838 GND notir3 x_op_jmp GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1839 GND notir3 op_push_pull GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1840 x_op_T3_ind_y ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1841 op_rti_rts ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1842 op_T2_jsr ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1843 op_T5_jsr ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1844 op_T2_stack_access ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1845 op_T0_tya ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1846 op_T__shift_a ir2 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1847 op_T0_txa ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1848 op_T0_pla ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1849 op_T0_tay ir2 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1850 op_T0_shift_a ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1851 op_T0_tax ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1852 op_T5_ind_y ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1853 op_branch_done ir2 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1854 op_T2_pha ir2 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1855 op_T0_shift_right_a ir2 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1856 op_T2_brk ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1857 op_T3_jsr ir2 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1858 op_T2_branch ir2 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1859 GND notir3 op_T2_php GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1860 GND notir3 op_T2_php_pha GND efet w=15 l=7
+ ad=0 pd=0 as=0 ps=0 
M1861 GND notir3 op_T4_jmp GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1862 GND notir3 op_T2_jmp_abs GND efet w=15 l=7
+ ad=0 pd=0 as=0 ps=0 
M1863 GND notir3 x_op_T3_plp_pla GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1864 GND notir3 op_T0_cli_sei GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1865 GND notir3 op_T0_clc_sec GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1866 n_1590 fetch n_1620 GND efet w=24 l=8
+ ad=120 pd=58 as=480 ps=112 
M1867 n_1083 cp1 n_1590 GND efet w=24 l=8
+ ad=1078 pd=268 as=0 ps=0 
M1868 n_1620 cclk notir3 GND efet w=11 l=7
+ ad=0 pd=0 as=0 ps=0 
M1869 GND notir3 op_T0_plp GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1870 GND notir3 op_T__cpx_cpy_abs GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1871 GND notir3 op_T__asl_rol_a GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1872 GND notir3 x_op_push_pull GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1873 GND notir3 op_T0_cld_sed GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1874 GND notir3 op_T3_mem_abs GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1875 GND notir3 op_T4_mem_abs_idx GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1876 GND notir3 op_clv GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1877 GND notir3 op_implied GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1878 op_T2_ind ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1879 op_T5_rts ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1880 op_T0_brk_rti ir2 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1881 op_T5_ind_x ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1882 x_op_T4_ind_y ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1883 op_T3_branch ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1884 op_brk_rti ir2 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1885 op_jsr ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1886 op_push_pull ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1887 op_T4_brk ir2 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1888 op_T2_php ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1889 op_T2_php_pha ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1890 op_T5_rti_rts ir2 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1891 xx_op_T5_jsr ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1892 x_op_T3_plp_pla ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1893 op_T0_cli_sei ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1894 op_T0_clc_sec ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1895 op_T0_plp ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1896 x_op_T4_rti ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1897 op_T__asl_rol_a ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1898 x_op_push_pull ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1899 op_T0_cld_sed ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1900 op_T5_mem_ind_idx ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1901 GND notir2 op_sty_cpy_mem GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1902 GND notir2 op_T2_idx_x_xy GND efet w=15 l=7
+ ad=0 pd=0 as=0 ps=0 
M1903 GND notir2 op_T0_ldy_mem GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1904 op_sty_cpy_mem ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1905 x_op_T0_tya ir6 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1906 op_xy ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1907 x_op_T0_txa ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1908 op_from_x ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1909 op_T0_txs ir6 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1910 GND notir2 op_jmp GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1911 GND notir2 op_T2_abs GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1912 GND notir2 op_T3_jmp GND efet w=13 l=7
+ ad=0 pd=0 as=0 ps=0 
M1913 op_clv ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1914 op_implied ir2 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1915 ir2 ir2 Vdd GND dfet w=10 l=7
+ ad=19647 pd=6500 as=0 ps=0 
M1916 GND notir2 op_T0_bit GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1917 GND notir2 op_T2_zp_zp_idx GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1918 op_T0_ldx_tax_tsx ir6 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1919 op_T0_tsx ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1920 op_T0_ldy_mem ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1921 op_T0_tay_ldy_not_idx ir6 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1922 op_T0_jsr ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1923 op_T5_brk ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1924 op_T0_ora ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1925 op_T4_brk_jsr ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1926 op_rol_ror ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1927 op_T2_jsr ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1928 op_shift ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1929 op_T5_jsr ir6 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1930 op_T0_tya ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1931 op_T0_txa ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1932 op_T0_lda ir6 GND GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1933 op_T0_tay ir6 GND GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1934 op_T0_tax ir6 GND GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1935 op_T0_bit ir6 GND GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1936 op_T0_and ir6 GND GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1937 GND notir2 op_T0_jmp GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1938 GND notir2 x_op_jmp GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1939 GND notir2 op_T4_jmp GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1940 GND notir2 op_T2_jmp_abs GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1941 GND notir2 op_T__bit GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1942 GND notir2 op_T3_mem_zp_idx GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1943 op_T2_brk ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1944 op_T3_jsr ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1945 op_sta_cmp ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1946 op_jsr ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1947 GND notir2 x_op_T0_bit GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1948 GND notir2 op_T__cpx_cpy_abs GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1949 GND notir2 op_T3_mem_abs GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1950 GND notir2 op_T2_mem_zp GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1951 GND n_1300 ir2 GND efet w=127 l=7
+ ad=0 pd=0 as=1414 ps=302 
M1952 notir2 notir2 Vdd GND dfet w=10 l=7
+ ad=19135 pd=6072 as=0 ps=0 
M1953 GND ir2 notir2 GND efet w=87 l=7
+ ad=0 pd=0 as=1908 ps=404 
M1954 n_343 fetch n_1300 GND efet w=23 l=8
+ ad=115 pd=56 as=471 ps=112 
M1955 n_571 cp1 n_343 GND efet w=23 l=9
+ ad=1314 pd=284 as=0 ps=0 
M1956 n_1300 cclk notir2 GND efet w=11 l=7
+ ad=0 pd=0 as=0 ps=0 
M1957 op_store ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1958 op_T4_brk ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1959 op_T2_php ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1960 xx_op_T5_jsr ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1961 op_asl_rol ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1962 op_T__bit ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1963 op_T0_clc_sec ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1964 x_op_T0_bit ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1965 op_T0_plp ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1966 op_T__asl_rol_a ir6 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M1967 GND notir6 op_T0_cpy_iny GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1968 GND notir6 op_T0_dex GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1969 GND notir6 op_T0_cpx_inx GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1970 GND notir6 op_T__dex GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1971 GND notir6 op_T__inx GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1972 GND notir6 op_T4_rts GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1973 GND notir6 op_T5_rti GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1974 GND notir6 op_ror GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1975 pipenVEC cclk nVEC GND efet w=11 l=8
+ ad=250 pd=96 as=1085 ps=328 
M1976 n_597 cp1 n_1339 GND efet w=13 l=7
+ ad=151 pd=76 as=793 ps=182 
M1977 n_1368 cp1 n_1149 GND efet w=13 l=7
+ ad=0 pd=0 as=175 ps=78 
M1978 op_sty_cpy_mem ir5 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1979 op_T0_iny_dey ir5 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1980 x_op_T0_tya ir5 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1981 op_T0_cpy_iny ir5 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1982 x_op_T0_txa ir5 GND GND efet w=15 l=7
+ ad=0 pd=0 as=0 ps=0 
M1983 op_T0_dex ir5 GND GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1984 op_from_x ir5 GND GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1985 op_T0_txs ir5 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1986 GND notir6 op_T0_eor GND efet w=15 l=7
+ ad=0 pd=0 as=0 ps=0 
M1987 GND notir6 op_jmp GND efet w=15 l=7
+ ad=0 pd=0 as=0 ps=0 
M1988 GND notir6 op_T4_rti GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M1989 GND notir6 op_inc_nop GND efet w=15 l=7
+ ad=0 pd=0 as=0 ps=0 
M1990 nop_branch_bit6 ir6 GND GND efet w=14 l=6
+ ad=599 pd=172 as=0 ps=0 
M1991 op_clv ir6 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1992 GND notir6 op_rti_rts GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1993 GND notir6 op_T0_cpx_cpy_inx_iny GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1994 GND notir6 op_T0_cmp GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1995 GND notir6 op_T0_sbc GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1996 GND notir6 op_T0_adc_sbc GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M1997 GND notir6 op_T3_jmp GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1998 GND notir6 op_T__adc_sbc GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M1999 GND notir6 op_T0_pla GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M2000 op_T__dex ir5 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M2001 op_T__iny_dey ir5 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2002 op_T5_brk ir5 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2003 op_T0_php_pha ir5 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2004 op_T5_rti ir5 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2005 GND notir6 op_T2_pha GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M2006 GND notir6 op_T0_shift_right_a GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2007 GND notir6 op_shift_right GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M2008 op_T0_eor ir5 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M2009 op_T0_ora ir5 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2010 op_T4_rti ir5 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2011 op_T0_cmp ir5 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2012 op_T0_tya ir5 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2013 op_T0_txa ir5 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2014 GND notir6 op_T5_rts GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2015 GND notir6 op_T0_jmp GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2016 GND notir6 x_op_jmp GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M2017 op_T2_pha ir5 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2018 op_T2_brk ir5 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2019 op_sta_cmp ir5 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2020 GND notir6 op_T4_jmp GND efet w=15 l=7
+ ad=0 pd=0 as=0 ps=0 
M2021 GND notir6 op_T5_rti_rts GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M2022 GND notir6 op_T2_jmp_abs GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M2023 GND notir6 op_lsr_ror_dec_inc GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M2024 GND notir6 op_T0_cli_sei GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M2025 ir6 ir6 Vdd GND dfet w=10 l=7
+ ad=19726 pd=6516 as=0 ps=0 
M2026 GND n_1675 ir6 GND efet w=129 l=7
+ ad=0 pd=0 as=1284 ps=304 
M2027 GND notir6 x_op_T__adc_sbc GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2028 GND notir6 x_op_T4_rti GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2029 GND notir6 op_T__cmp GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2030 GND notir6 op_T__cpx_cpy_abs GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2031 GND notir6 op_T__cpx_cpy_imm_zp GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2032 GND notir6 op_T0_cld_sed GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M2033 op_T0_brk_rti ir5 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M2034 op_brk_rti ir5 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M2035 op_store ir5 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2036 op_T4_brk ir5 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2037 op_T2_php ir5 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M2038 op_T2_php_pha ir5 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2039 op_T2_jmp_abs ir5 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2040 notir6 notir6 Vdd GND dfet w=10 l=7
+ ad=18955 pd=6062 as=0 ps=0 
M2041 GND ir6 notir6 GND efet w=88 l=7
+ ad=0 pd=0 as=1837 ps=420 
M2042 x_op_T4_rti ir5 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2043 op_T__cmp ir5 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M2044 n_1339 n_1339 Vdd GND dfet w=10 l=12
+ ad=330 pd=92 as=0 ps=0 
M2045 GND n_799 n_1339 GND efet w=71 l=7
+ ad=0 pd=0 as=0 ps=0 
M2046 nNMIG cclk n_1693 GND efet w=13 l=7
+ ad=2275 pd=538 as=225 ps=84 
M2047 n_799 cclk nNMIG GND efet w=12 l=7
+ ad=200 pd=86 as=0 ps=0 
M2048 GND notir5 op_T0_cpx_inx GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2049 GND n_1149 nNMIG GND efet w=109 l=7
+ ad=0 pd=0 as=0 ps=0 
M2050 op_T0_cpy_iny clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2051 op_T0_iny_dey clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2052 x_op_T0_tya clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2053 GND notir5 op_T0_ldx_tax_tsx GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M2054 GND notir5 op_T__inx GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2055 GND notir5 op_T0_tsx GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2056 GND notir5 op_T0_ldy_mem GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2057 GND notir5 op_T0_tay_ldy_not_idx GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2058 GND notir5 op_T0_jsr GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M2059 GND notir5 op_T4_rts GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2060 GND notir5 op_T3_plp_pla GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M2061 GND notir5 op_ror GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M2062 x_op_T0_txa clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2063 op_T0_dex clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2064 op_T0_cpx_inx clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2065 op_T0_txs clock1 GND GND efet w=16 l=6
+ ad=0 pd=0 as=0 ps=0 
M2066 op_T0_tay_ldy_not_idx clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2067 GND notir5 op_plp_pla GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2068 GND notir5 op_inc_nop GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2069 GND notir5 op_T2_jsr GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2070 GND notir5 op_T0_sbc GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2071 GND notir5 op_T0_adc_sbc GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2072 GND notir5 op_rol_ror GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M2073 op_T0_ldx_tax_tsx clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2074 op_T0_tsx clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2075 op_T0_ldy_mem clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2076 op_T0_jsr clock1 GND GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M2077 op_T0_php_pha clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2078 op_T0_eor clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2079 op_T0_ora clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2080 op_T0 clock1 GND GND efet w=15 l=6
+ ad=551 pd=136 as=0 ps=0 
M2081 GND notir5 op_T5_jsr GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M2082 GND notir5 op_T__adc_sbc GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M2083 GND notir5 op_T0_pla GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2084 GND notir5 op_T0_lda GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2085 GND notir5 op_T0_tay GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2086 GND notir5 op_T0_tax GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M2087 GND notir5 op_T0_bit GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2088 GND notir5 op_T0_and GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M2089 GND notir5 op_T3_jsr GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M2090 op_T0_cpx_cpy_inx_iny clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2091 op_T0_cmp clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2092 op_T0_sbc clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2093 op_T0_adc_sbc clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2094 op_T0_tya clock1 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M2095 op_T0_txa clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2096 op_T0_pla clock1 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M2097 op_T0_lda clock1 GND GND efet w=15 l=7
+ ad=0 pd=0 as=0 ps=0 
M2098 op_T0_acc clock1 GND GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M2099 op_T0_tay clock1 GND GND efet w=13 l=7
+ ad=0 pd=0 as=0 ps=0 
M2100 op_T0_shift_a clock1 GND GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M2101 op_T0_tax clock1 GND GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M2102 op_T0_bit clock1 GND GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M2103 op_T0_and clock1 GND GND efet w=13 l=7
+ ad=0 pd=0 as=0 ps=0 
M2104 GND notir5 op_T5_rts GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2105 GND notir5 op_jsr GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2106 GND notir5 xx_op_T5_jsr GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M2107 GND notir5 x_op_T3_plp_pla GND efet w=13 l=7
+ ad=0 pd=0 as=0 ps=0 
M2108 GND notir5 op_T__bit GND efet w=13 l=7
+ ad=0 pd=0 as=0 ps=0 
M2109 GND notir5 x_op_T__adc_sbc GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2110 GND notir5 x_op_T0_bit GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2111 GND notir5 op_T0_plp GND efet w=15 l=6
+ ad=0 pd=0 as=0 ps=0 
M2112 n_74 fetch n_1675 GND efet w=23 l=8
+ ad=115 pd=56 as=439 ps=108 
M2113 n_1309 cp1 n_74 GND efet w=23 l=10
+ ad=1258 pd=366 as=0 ps=0 
M2114 n_1675 cclk notir6 GND efet w=13 l=8
+ ad=0 pd=0 as=0 ps=0 
M2115 op_branch_done clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2116 op_T0_shift_right_a clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2117 op_T0_brk_rti clock1 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M2118 op_T0_jmp clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2119 GND notir5 op_clv GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2120 op_T0_cli_sei clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2121 op_T0_clc_sec clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2122 x_op_T0_bit clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2123 op_T0_plp clock1 GND GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M2124 ir5 ir5 Vdd GND dfet w=10 l=7
+ ad=19819 pd=6546 as=0 ps=0 
M2125 op_T0_cld_sed clock1 GND GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2126 GND n_1609 ir5 GND efet w=126 l=7
+ ad=0 pd=0 as=1394 ps=304 
M2127 GND n_1693 n_1312 GND efet w=60 l=6
+ ad=0 pd=0 as=720 ps=232 
M2128 Vdd n_1312 n_1312 GND dfet w=10 l=16
+ ad=0 pd=0 as=1278 ps=354 
M2129 n_1312 n_1291 GND GND efet w=59 l=7
+ ad=0 pd=0 as=0 ps=0 
M2130 nNMIG nNMIG Vdd GND dfet w=10 l=8
+ ad=6478 pd=2174 as=0 ps=0 
M2131 GND n_1312 nNMIG GND efet w=54 l=6
+ ad=0 pd=0 as=0 ps=0 
M2132 GND clock2 op_T__dex GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M2133 GND clock2 op_T__inx GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M2134 GND clock2 op_T__iny_dey GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M2135 brk_done notRdy0 GND GND efet w=86 l=6
+ ad=2025 pd=460 as=0 ps=0 
M2136 n_1291 cp1 brk_done GND efet w=13 l=8
+ ad=234 pd=92 as=0 ps=0 
M2137 Vdd brk_done brk_done GND dfet w=9 l=8
+ ad=0 pd=0 as=12990 ps=4446 
M2138 GND n_861 brk_done GND efet w=96 l=6
+ ad=0 pd=0 as=0 ps=0 
M2139 GND n_1452 n_861 GND efet w=76 l=7
+ ad=0 pd=0 as=1124 ps=296 
M2140 Vdd n_861 n_861 GND dfet w=10 l=12
+ ad=0 pd=0 as=1930 ps=586 
M2141 VEC1 cclk n_1452 GND efet w=12 l=9
+ ad=985 pd=290 as=232 ps=88 
M2142 n_912 VEC1 GND GND efet w=48 l=7
+ ad=434 pd=138 as=0 ps=0 
M2143 n_912 notRdy0 n_1290 GND efet w=39 l=6
+ ad=0 pd=0 as=1366 ps=360 
M2144 Vdd n_1290 n_1290 GND dfet w=10 l=17
+ ad=0 pd=0 as=782 ps=226 
M2145 n_1290 n_1126 GND GND efet w=44 l=6
+ ad=0 pd=0 as=0 ps=0 
M2146 n_1717 op_T2_abs_y GND GND efet w=30 l=7
+ ad=3182 pd=730 as=0 ps=0 
M2147 GND op_T0_iny_dey n_1717 GND efet w=30 l=7
+ ad=0 pd=0 as=0 ps=0 
M2148 n_1717 x_op_T0_tya GND GND efet w=30 l=7
+ ad=0 pd=0 as=0 ps=0 
M2149 GND op_T0_cpy_iny n_1717 GND efet w=30 l=6
+ ad=0 pd=0 as=0 ps=0 
M2150 n_1717 op_T3_ind_y GND GND efet w=31 l=7
+ ad=0 pd=0 as=0 ps=0 
M2151 n_1717 n_1717 Vdd GND dfet w=10 l=15
+ ad=6985 pd=2378 as=0 ps=0 
M2152 n_1303 n_1303 Vdd GND dfet w=10 l=14
+ ad=2706 pd=880 as=0 ps=0 
M2153 n_1303 n_335 n_508 GND efet w=73 l=6
+ ad=1421 pd=362 as=588 ps=200 
M2154 n_508 op_from_x GND GND efet w=82 l=6
+ ad=0 pd=0 as=0 ps=0 
M2155 n_1126 cclk VEC0 GND efet w=12 l=8
+ ad=210 pd=70 as=2021 ps=518 
M2156 n_1290 cp1 n_698 GND efet w=12 l=8
+ ad=0 pd=0 as=170 ps=76 
M2157 n_1397 n_335 n_1303 GND efet w=59 l=6
+ ad=295 pd=128 as=0 ps=0 
M2158 GND op_sty_cpy_mem n_1397 GND efet w=59 l=7
+ ad=0 pd=0 as=0 ps=0 
M2159 n_1604 op_sty_cpy_mem GND GND efet w=59 l=7
+ ad=295 pd=128 as=0 ps=0 
M2160 n_1717 n_335 n_1604 GND efet w=59 l=6
+ ad=0 pd=0 as=0 ps=0 
M2161 n_1106 op_T2_ind_x GND GND efet w=30 l=7
+ ad=3038 pd=700 as=0 ps=0 
M2162 GND x_op_T0_txa n_1106 GND efet w=30 l=6
+ ad=0 pd=0 as=0 ps=0 
M2163 n_1106 op_T0_dex GND GND efet w=30 l=6
+ ad=0 pd=0 as=0 ps=0 
M2164 GND op_T0_cpx_inx n_1106 GND efet w=30 l=7
+ ad=0 pd=0 as=0 ps=0 
M2165 n_1106 n_1106 Vdd GND dfet w=9 l=14
+ ad=7193 pd=2712 as=0 ps=0 
M2166 GND op_T0_txs n_1106 GND efet w=30 l=6
+ ad=0 pd=0 as=0 ps=0 
M2167 Vdd n_1244 n_1244 GND dfet w=10 l=17
+ ad=0 pd=0 as=1121 ps=314 
M2168 n_1351 op_T2_idx_x_xy n_1717 GND efet w=60 l=7
+ ad=497 pd=140 as=0 ps=0 
M2169 GND op_xy n_1351 GND efet w=62 l=6
+ ad=0 pd=0 as=0 ps=0 
M2170 n_1244 op_xy GND GND efet w=34 l=6
+ ad=418 pd=114 as=0 ps=0 
M2171 GND clock2 op_T__ora_and_eor_adc GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2172 GND clock2 op_T__adc_sbc GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M2173 GND clock2 op_T__shift_a GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2174 n_844 op_T0_ldx_tax_tsx GND GND efet w=29 l=6
+ ad=1424 pd=378 as=0 ps=0 
M2175 GND op_T__dex n_844 GND efet w=29 l=5
+ ad=0 pd=0 as=0 ps=0 
M2176 n_844 op_T__inx GND GND efet w=29 l=7
+ ad=0 pd=0 as=0 ps=0 
M2177 GND op_T__iny_dey n_616 GND efet w=29 l=6
+ ad=0 pd=0 as=1384 ps=372 
M2178 n_616 op_T0_ldy_mem GND GND efet w=29 l=6
+ ad=0 pd=0 as=0 ps=0 
M2179 GND op_T0_tay_ldy_not_idx n_616 GND efet w=29 l=6
+ ad=0 pd=0 as=0 ps=0 
M2180 n_1464 op_T0_jsr GND GND efet w=26 l=7
+ ad=2181 pd=504 as=0 ps=0 
M2181 GND op_T5_brk n_1464 GND efet w=26 l=7
+ ad=0 pd=0 as=0 ps=0 
M2182 n_1464 op_T0_php_pha GND GND efet w=26 l=7
+ ad=0 pd=0 as=0 ps=0 
M2183 GND op_T4_rts n_1464 GND efet w=26 l=7
+ ad=0 pd=0 as=0 ps=0 
M2184 n_1464 op_T3_plp_pla GND GND efet w=26 l=7
+ ad=0 pd=0 as=0 ps=0 
M2185 GND op_T5_rti n_1464 GND efet w=26 l=8
+ ad=0 pd=0 as=0 ps=0 
M2186 n_844 n_844 Vdd GND dfet w=9 l=17
+ ad=7505 pd=2780 as=0 ps=0 
M2187 VEC0 notRdy0 GND GND efet w=39 l=6
+ ad=0 pd=0 as=0 ps=0 
M2188 GND n_698 VEC1 GND efet w=61 l=8
+ ad=0 pd=0 as=0 ps=0 
M2189 Vdd VEC1 VEC1 GND dfet w=11 l=11
+ ad=0 pd=0 as=2851 ps=846 
M2190 GND VEC1 nVEC GND efet w=38 l=7
+ ad=0 pd=0 as=0 ps=0 
M2191 Vdd nVEC nVEC GND dfet w=10 l=10
+ ad=0 pd=0 as=9123 ps=3054 
M2192 nVEC VEC0 GND GND efet w=37 l=6
+ ad=0 pd=0 as=0 ps=0 
M2193 n_445 n_862 GND GND efet w=173 l=6
+ ad=884 pd=254 as=0 ps=0 
M2194 n_1103 n_1244 GND GND efet w=58 l=7
+ ad=232 pd=124 as=0 ps=0 
M2195 n_1106 op_T2_idx_x_xy n_1103 GND efet w=58 l=7
+ ad=0 pd=0 as=0 ps=0 
M2196 n_734 n_335 n_1106 GND efet w=59 l=6
+ ad=649 pd=140 as=0 ps=0 
M2197 GND op_from_x n_734 GND efet w=59 l=6
+ ad=0 pd=0 as=0 ps=0 
M2198 Vdd VEC0 VEC0 GND dfet w=10 l=14
+ ad=0 pd=0 as=6005 ps=2088 
M2199 Vdd n_946 n_946 GND dfet w=9 l=13
+ ad=0 pd=0 as=1224 ps=376 
M2200 n_616 n_616 Vdd GND dfet w=8 l=16
+ ad=7828 pd=2838 as=0 ps=0 
M2201 Vdd n_1586 n_1586 GND dfet w=10 l=16
+ ad=0 pd=0 as=7228 ps=2672 
M2202 VEC0 n_689 GND GND efet w=34 l=6
+ ad=0 pd=0 as=0 ps=0 
M2203 n_454 n_844 n_946 GND efet w=60 l=7
+ ad=387 pd=138 as=1142 ps=292 
M2204 GND n_616 n_454 GND efet w=63 l=5
+ ad=0 pd=0 as=0 ps=0 
M2205 n_1586 op_T0_tsx GND GND efet w=31 l=7
+ ad=679 pd=216 as=0 ps=0 
M2206 n_1464 n_1464 Vdd GND dfet w=9 l=17
+ ad=767 pd=206 as=0 ps=0 
M2207 n_1109 n_1464 GND GND efet w=35 l=7
+ ad=1397 pd=372 as=0 ps=0 
M2208 GND op_T5_brk n_689 GND efet w=27 l=7
+ ad=0 pd=0 as=544 ps=174 
M2209 Vdd n_1109 n_1109 GND dfet w=9 l=13
+ ad=0 pd=0 as=3576 ps=1116 
M2210 Vdd n_632 n_632 GND dfet w=9 l=16
+ ad=0 pd=0 as=5801 ps=2108 
M2211 Vdd n_1358 n_1358 GND dfet w=9 l=10
+ ad=0 pd=0 as=5570 ps=2110 
M2212 n_689 n_689 Vdd GND dfet w=10 l=17
+ ad=1409 pd=430 as=0 ps=0 
M2213 n_632 op_T2_stack GND GND efet w=34 l=7
+ ad=1109 pd=352 as=0 ps=0 
M2214 Vdd n_1714 n_1714 GND dfet w=10 l=16
+ ad=0 pd=0 as=1116 ps=342 
M2215 n_445 n_445 Vdd GND dfet w=17 l=6
+ ad=9205 pd=3050 as=0 ps=0 
M2216 n_317 n_445 GND GND efet w=48 l=7
+ ad=455 pd=150 as=0 ps=0 
M2217 n_1714 pipeUNK26 GND GND efet w=59 l=6
+ ad=876 pd=200 as=0 ps=0 
M2218 pipeUNK26 cclk n_132 GND efet w=11 l=8
+ ad=131 pd=56 as=707 ps=224 
M2219 Vdd n_317 n_317 GND dfet w=10 l=10
+ ad=0 pd=0 as=1532 ps=506 
M2220 GND n_445 n_417 GND efet w=73 l=7
+ ad=0 pd=0 as=1512 ps=374 
M2221 Vdd n_317 n_417 GND dfet w=16 l=7
+ ad=0 pd=0 as=0 ps=0 
M2222 n_417 n_445 GND GND efet w=54 l=6
+ ad=0 pd=0 as=0 ps=0 
M2223 sync n_445 GND GND efet w=182 l=7
+ ad=18998 pd=2444 as=0 ps=0 
M2224 Vdd n_417 sync GND efet w=93 l=6
+ ad=0 pd=0 as=0 ps=0 
M2225 Vdd n_417 sync GND efet w=173 l=6
+ ad=0 pd=0 as=0 ps=0 
M2226 GND n_445 sync GND efet w=182 l=6
+ ad=0 pd=0 as=0 ps=0 
M2227 sync n_417 Vdd GND efet w=158 l=6
+ ad=0 pd=0 as=0 ps=0 
M2228 sync n_445 GND GND efet w=182 l=6
+ ad=0 pd=0 as=0 ps=0 
M2229 Vdd n_417 sync GND efet w=133 l=7
+ ad=0 pd=0 as=0 ps=0 
M2230 GND n_445 sync GND efet w=182 l=6
+ ad=0 pd=0 as=0 ps=0 
M2231 sync n_417 Vdd GND efet w=127 l=7
+ ad=0 pd=0 as=0 ps=0 
M2232 GND n_1447 n_1175 GND efet w=50 l=7
+ ad=0 pd=0 as=623 ps=216 
M2233 n_1175 n_1175 Vdd GND dfet w=9 l=17
+ ad=1377 pd=400 as=0 ps=0 
M2234 n_1447 cp1 n_262 GND efet w=11 l=7
+ ad=238 pd=90 as=1499 ps=380 
M2235 Vdd n_169 n_169 GND dfet w=9 l=18
+ ad=0 pd=0 as=398 ps=88 
M2236 pipeUNK29 cclk n_169 GND efet w=12 l=7
+ ad=169 pd=72 as=904 ps=274 
M2237 n_1058 n_1289 n_632 GND efet w=51 l=7
+ ad=306 pd=114 as=0 ps=0 
M2238 GND op_T0_jsr n_1058 GND efet w=51 l=6
+ ad=0 pd=0 as=0 ps=0 
M2239 n_1358 n_1109 GND GND efet w=52 l=6
+ ad=1756 pd=468 as=0 ps=0 
M2240 n_1358 op_T0_txs GND GND efet w=45 l=6
+ ad=0 pd=0 as=0 ps=0 
M2241 GND n_917 n_1358 GND efet w=55 l=6
+ ad=0 pd=0 as=0 ps=0 
M2242 n_267 n_267 Vdd GND dfet w=10 l=15
+ ad=5060 pd=1842 as=0 ps=0 
M2243 n_1175 cclk pipeUNK28 GND efet w=11 l=8
+ ad=0 pd=0 as=163 ps=72 
M2244 GND n_1175 n_267 GND efet w=44 l=7
+ ad=0 pd=0 as=1900 ps=460 
M2245 n_169 n_1624 GND GND efet w=53 l=6
+ ad=0 pd=0 as=0 ps=0 
M2246 GND n_139 n_169 GND efet w=53 l=6
+ ad=0 pd=0 as=0 ps=0 
M2247 n_1189 pipeUNK29 GND GND efet w=100 l=6
+ ad=781 pd=224 as=0 ps=0 
M2248 n_262 n_1714 n_1189 GND efet w=77 l=6
+ ad=0 pd=0 as=0 ps=0 
M2249 n_267 n_544 GND GND efet w=29 l=7
+ ad=0 pd=0 as=0 ps=0 
M2250 n_917 notRdy0 GND GND efet w=27 l=7
+ ad=759 pd=176 as=0 ps=0 
M2251 GND n_383 n_917 GND efet w=27 l=6
+ ad=0 pd=0 as=0 ps=0 
M2252 n_1624 cp1 notRdy0 GND efet w=12 l=7
+ ad=364 pd=124 as=2200 ps=666 
M2253 n_1598 n_1511 n_262 GND efet w=46 l=7
+ ad=509 pd=154 as=0 ps=0 
M2254 GND pipeUNK28 n_1598 GND efet w=69 l=5
+ ad=0 pd=0 as=0 ps=0 
M2255 n_262 n_262 Vdd GND dfet w=10 l=27
+ ad=531 pd=116 as=0 ps=0 
M2256 GND n_785 n_267 GND efet w=41 l=7
+ ad=0 pd=0 as=0 ps=0 
M2257 n_920 cp1 n_785 GND efet w=11 l=6
+ ad=619 pd=190 as=149 ps=58 
M2258 GND pipeUNK29 n_1511 GND efet w=49 l=6
+ ad=0 pd=0 as=423 ps=146 
M2259 n_139 n_139 Vdd GND dfet w=10 l=16
+ ad=1212 pd=382 as=0 ps=0 
M2260 n_1511 n_1511 Vdd GND dfet w=9 l=17
+ ad=1029 pd=294 as=0 ps=0 
M2261 GND pipeUNK27 n_920 GND efet w=44 l=5
+ ad=0 pd=0 as=0 ps=0 
M2262 Vdd n_917 n_917 GND dfet w=10 l=12
+ ad=0 pd=0 as=817 ps=266 
M2263 notRdy0 cp1 n_902 GND efet w=12 l=8
+ ad=0 pd=0 as=149 ps=72 
M2264 n_1109 n_902 GND GND efet w=46 l=6
+ ad=0 pd=0 as=0 ps=0 
M2265 GND n_902 n_1109 GND efet w=35 l=7
+ ad=0 pd=0 as=0 ps=0 
M2266 n_1289 n_1289 Vdd GND dfet w=10 l=17
+ ad=1779 pd=588 as=0 ps=0 
M2267 GND n_902 n_1289 GND efet w=52 l=6
+ ad=0 pd=0 as=764 ps=202 
M2268 n_920 n_920 Vdd GND dfet w=10 l=17
+ ad=459 pd=110 as=0 ps=0 
M2269 op_SRS cclk pipeUNK27 GND efet w=12 l=9
+ ad=713 pd=270 as=171 ps=78 
M2270 GND op_SRS n_139 GND efet w=38 l=7
+ ad=0 pd=0 as=766 ps=192 
M2271 Vdd n_728 n_728 GND dfet w=10 l=16
+ ad=0 pd=0 as=1542 ps=498 
M2272 n_728 VEC0 GND GND efet w=26 l=7
+ ad=665 pd=174 as=0 ps=0 
M2273 sync n_445 GND GND efet w=182 l=5
+ ad=0 pd=0 as=0 ps=0 
M2274 Vdd n_417 sync GND efet w=127 l=6
+ ad=0 pd=0 as=0 ps=0 
M2275 sync n_417 Vdd GND efet w=127 l=7
+ ad=0 pd=0 as=0 ps=0 
M2276 Vdd n_1712 n_1712 GND dfet w=10 l=10
+ ad=0 pd=0 as=941 ps=338 
M2277 Vdd C1x5Reset C1x5Reset GND dfet w=10 l=7
+ ad=0 pd=0 as=8565 ps=2934 
M2278 Vdd n_1087 n_1087 GND dfet w=9 l=7
+ ad=0 pd=0 as=302 ps=110 
M2279 GND nVEC n_1712 GND efet w=37 l=6
+ ad=0 pd=0 as=1534 ps=360 
M2280 n_1712 nNMIG GND GND efet w=37 l=6
+ ad=0 pd=0 as=0 ps=0 
M2281 GND C1x5Reset n_1712 GND efet w=38 l=6
+ ad=0 pd=0 as=0 ps=0 
M2282 GND n_717 C1x5Reset GND efet w=63 l=6
+ ad=0 pd=0 as=873 ps=224 
M2283 Vdd n_717 n_717 GND dfet w=9 l=17
+ ad=0 pd=0 as=1877 ps=630 
M2284 Reset0 cclk pipephi2Reset0x GND efet w=11 l=9
+ ad=0 pd=0 as=161 ps=68 
M2285 n_1087 brk_done GND GND efet w=55 l=6
+ ad=1341 pd=280 as=0 ps=0 
M2286 GND n_717 n_1087 GND efet w=55 l=6
+ ad=0 pd=0 as=0 ps=0 
M2287 n_717 n_1132 GND GND efet w=46 l=6
+ ad=686 pd=202 as=0 ps=0 
M2288 GND pipephi2Reset0x n_717 GND efet w=47 l=6
+ ad=0 pd=0 as=0 ps=0 
M2289 n_1132 cp1 n_1087 GND efet w=11 l=7
+ ad=262 pd=88 as=0 ps=0 
M2290 n_696 n_0_ADL0 GND GND efet w=42 l=6
+ ad=1455 pd=418 as=0 ps=0 
M2291 n_696 n_79 n_911 GND efet w=97 l=7
+ ad=0 pd=0 as=2583 ps=548 
M2292 n_728 cclk pipeVectorA0 GND efet w=11 l=9
+ ad=0 pd=0 as=145 ps=70 
M2293 n_696 n_696 Vdd GND dfet w=9 l=8
+ ad=1699 pd=556 as=0 ps=0 
M2294 n_70 nVEC GND GND efet w=37 l=7
+ ad=845 pd=192 as=0 ps=0 
M2295 GND n_1054 n_70 GND efet w=37 l=7
+ ad=0 pd=0 as=0 ps=0 
M2296 n_1054 C1x5Reset GND GND efet w=37 l=6
+ ad=686 pd=194 as=0 ps=0 
M2297 n_70 n_70 Vdd GND dfet w=10 l=10
+ ad=1152 pd=376 as=0 ps=0 
M2298 n_1712 cclk pipeVectorA2 GND efet w=11 l=9
+ ad=0 pd=0 as=140 ps=66 
M2299 GND op_ror n_544 GND efet w=58 l=7
+ ad=0 pd=0 as=1024 ps=234 
M2300 GND op_T3_stack_bit_jmp n_604 GND efet w=34 l=6
+ ad=0 pd=0 as=2928 ps=818 
M2301 n_604 op_T2_stack GND GND efet w=36 l=6
+ ad=0 pd=0 as=0 ps=0 
M2302 GND op_T0 n_638 GND efet w=35 l=6
+ ad=0 pd=0 as=524 ps=146 
M2303 n_604 op_T4_brk_jsr GND GND efet w=37 l=6
+ ad=0 pd=0 as=0 ps=0 
M2304 GND op_T4_rti n_604 GND efet w=30 l=6
+ ad=0 pd=0 as=0 ps=0 
M2305 n_638 n_638 Vdd GND dfet w=9 l=16
+ ad=886 pd=278 as=0 ps=0 
M2306 n_604 n_604 Vdd GND dfet w=10 l=15
+ ad=7670 pd=2660 as=0 ps=0 
M2307 GND op_T3_ind_x n_604 GND efet w=35 l=5
+ ad=0 pd=0 as=0 ps=0 
M2308 n_1107 op_T3_ind_x GND GND efet w=33 l=5
+ ad=1821 pd=500 as=0 ps=0 
M2309 GND op_T4_ind_y n_1107 GND efet w=34 l=6
+ ad=0 pd=0 as=0 ps=0 
M2310 n_1107 op_T2_ind_y GND GND efet w=33 l=6
+ ad=0 pd=0 as=0 ps=0 
M2311 GND op_T3_abs_idx n_1107 GND efet w=33 l=6
+ ad=0 pd=0 as=0 ps=0 
M2312 n_1107 op_plp_pla GND GND efet w=39 l=5
+ ad=0 pd=0 as=0 ps=0 
M2313 n_1649 op_jmp GND GND efet w=34 l=6
+ ad=2795 pd=766 as=0 ps=0 
M2314 GND op_T2_abs n_1649 GND efet w=46 l=6
+ ad=0 pd=0 as=0 ps=0 
M2315 n_544 n_544 Vdd GND dfet w=10 l=13
+ ad=1561 pd=502 as=0 ps=0 
M2316 n_1118 op_T2_ADL_ADD GND GND efet w=55 l=6
+ ad=330 pd=122 as=0 ps=0 
M2317 n_604 n_638 n_1118 GND efet w=55 l=6
+ ad=0 pd=0 as=0 ps=0 
M2318 Vdd n_1649 n_1649 GND dfet w=10 l=14
+ ad=0 pd=0 as=5807 ps=2160 
M2319 n_1555 op_inc_nop n_1107 GND efet w=53 l=8
+ ad=265 pd=116 as=0 ps=0 
M2320 GND n_440 n_1555 GND efet w=53 l=6
+ ad=0 pd=0 as=0 ps=0 
M2321 n_300 x_op_T3_ind_y GND GND efet w=30 l=6
+ ad=2459 pd=698 as=0 ps=0 
M2322 GND op_rti_rts n_300 GND efet w=33 l=6
+ ad=0 pd=0 as=0 ps=0 
M2323 n_1000 op_T0_adc_sbc GND GND efet w=70 l=6
+ ad=1146 pd=342 as=0 ps=0 
M2324 GND op_T4_ind_x n_300 GND efet w=39 l=6
+ ad=0 pd=0 as=0 ps=0 
M2325 GND op_T2_jsr n_300 GND efet w=40 l=6
+ ad=0 pd=0 as=0 ps=0 
M2326 n_1560 op_T0_cpx_cpy_inx_iny GND GND efet w=26 l=6
+ ad=950 pd=230 as=0 ps=0 
M2327 GND op_T0_cmp n_1560 GND efet w=26 l=6
+ ad=0 pd=0 as=0 ps=0 
M2328 n_1560 n_1055 GND GND efet w=28 l=6
+ ad=0 pd=0 as=0 ps=0 
M2329 Vdd n_1107 n_1107 GND dfet w=10 l=17
+ ad=0 pd=0 as=608 ps=168 
M2330 Vdd n_383 n_383 GND dfet w=10 l=14
+ ad=0 pd=0 as=2291 ps=696 
M2331 n_389 n_1107 GND GND efet w=37 l=6
+ ad=674 pd=188 as=0 ps=0 
M2332 Vdd n_389 n_389 GND dfet w=10 l=13
+ ad=0 pd=0 as=2882 ps=948 
M2333 n_1560 n_1560 Vdd GND dfet w=8 l=15
+ ad=933 pd=304 as=0 ps=0 
M2334 GND op_rol_ror n_1000 GND efet w=53 l=7
+ ad=0 pd=0 as=0 ps=0 
M2335 n_980 op_T3_jmp GND GND efet w=36 l=6
+ ad=709 pd=184 as=0 ps=0 
M2336 n_300 n_300 Vdd GND dfet w=9 l=13
+ ad=2679 pd=1022 as=0 ps=0 
M2337 GND op_T2_jsr n_383 GND efet w=45 l=7
+ ad=0 pd=0 as=589 ps=174 
M2338 GND op_T0_ora n_1145 GND efet w=38 l=6
+ ad=0 pd=0 as=722 ps=256 
M2339 Vdd n_837 n_837 GND dfet w=10 l=17
+ ad=0 pd=0 as=2929 ps=970 
M2340 n_837 op_T0_eor GND GND efet w=40 l=6
+ ad=827 pd=228 as=0 ps=0 
M2341 n_1145 n_1145 Vdd GND dfet w=10 l=14
+ ad=1387 pd=464 as=0 ps=0 
M2342 GND op_rti_rts n_1649 GND efet w=46 l=6
+ ad=0 pd=0 as=0 ps=0 
M2343 Vdd n_480 n_480 GND dfet w=10 l=10
+ ad=0 pd=0 as=1151 ps=366 
M2344 n_480 nNMIG n_1092 GND efet w=79 l=6
+ ad=1226 pd=350 as=1712 ps=394 
M2345 GND nIRQP n_1092 GND efet w=72 l=6
+ ad=0 pd=0 as=0 ps=0 
M2346 n_1092 n_118 GND GND efet w=82 l=6
+ ad=0 pd=0 as=0 ps=0 
M2347 n_1145 notRdy0 GND GND efet w=32 l=5
+ ad=0 pd=0 as=0 ps=0 
M2348 GND op_rti_rts n_1377 GND efet w=38 l=6
+ ad=0 pd=0 as=423 ps=132 
M2349 n_1377 n_1377 Vdd GND dfet w=9 l=17
+ ad=1128 pd=320 as=0 ps=0 
M2350 n_1040 n_383 GND GND efet w=65 l=7
+ ad=1107 pd=278 as=0 ps=0 
M2351 n_1649 n_389 GND GND efet w=30 l=5
+ ad=0 pd=0 as=0 ps=0 
M2352 GND op_T4_ind_x n_1649 GND efet w=31 l=7
+ ad=0 pd=0 as=0 ps=0 
M2353 Vdd n_385 n_385 GND dfet w=9 l=13
+ ad=0 pd=0 as=306 ps=86 
M2354 n_604 notRdy0 GND GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M2355 n_385 n_604 GND GND efet w=51 l=6
+ ad=881 pd=276 as=0 ps=0 
M2356 GND n_1377 n_385 GND efet w=49 l=6
+ ad=0 pd=0 as=0 ps=0 
M2357 GND n_1145 op_ORS GND efet w=44 l=6
+ ad=0 pd=0 as=493 ps=166 
M2358 op_ORS op_ORS Vdd GND dfet w=8 l=9
+ ad=4746 pd=1706 as=0 ps=0 
M2359 n_202 nnT2BR GND GND efet w=46 l=8
+ ad=924 pd=264 as=0 ps=0 
M2360 n_202 n_646 GND GND efet w=46 l=6
+ ad=0 pd=0 as=0 ps=0 
M2361 n_629 n_480 n_202 GND efet w=47 l=7
+ ad=2001 pd=502 as=0 ps=0 
M2362 Vdd n_629 n_629 GND dfet w=10 l=16
+ ad=0 pd=0 as=1448 ps=462 
M2363 n_1040 n_383 GND GND efet w=30 l=7
+ ad=0 pd=0 as=0 ps=0 
M2364 n_782 n_1303 n_1040 GND efet w=94 l=6
+ ad=1741 pd=394 as=0 ps=0 
M2365 Vdd n_782 n_782 GND dfet w=9 l=7
+ ad=0 pd=0 as=512 ps=178 
M2366 n_1649 notRdy0 GND GND efet w=37 l=7
+ ad=0 pd=0 as=0 ps=0 
M2367 GND n_1109 n_1649 GND efet w=43 l=6
+ ad=0 pd=0 as=0 ps=0 
M2368 GND brk_done n_300 GND efet w=50 l=6
+ ad=0 pd=0 as=0 ps=0 
M2369 n_1649 brk_done GND GND efet w=31 l=6
+ ad=0 pd=0 as=0 ps=0 
M2370 GND op_T2_jsr n_1649 GND efet w=36 l=6
+ ad=0 pd=0 as=0 ps=0 
M2371 n_385 cclk pipeUNK30 GND efet w=12 l=7
+ ad=0 pd=0 as=159 ps=66 
M2372 Vdd n_1178 n_1178 GND dfet w=10 l=13
+ ad=0 pd=0 as=3313 ps=1134 
M2373 GND pipeUNK31 n_1178 GND efet w=60 l=6
+ ad=0 pd=0 as=1900 ps=546 
M2374 GND pipeVectorA2 n_815 GND efet w=51 l=7
+ ad=0 pd=0 as=714 ps=204 
M2375 n_1054 n_1054 Vdd GND dfet w=10 l=9
+ ad=698 pd=226 as=0 ps=0 
M2376 Vdd n_0_ADL0 n_0_ADL0 GND dfet w=10 l=17
+ ad=0 pd=0 as=4325 ps=1410 
M2377 GND pipeVectorA0 n_0_ADL0 GND efet w=105 l=7
+ ad=0 pd=0 as=1298 ps=344 
M2378 n_1117 cclk pipeVectorA1 GND efet w=11 l=7
+ ad=801 pd=242 as=149 ps=72 
M2379 n_815 n_815 Vdd GND dfet w=9 l=16
+ ad=1112 pd=280 as=0 ps=0 
M2380 n_1117 n_1117 Vdd GND dfet w=10 l=9
+ ad=390 pd=124 as=0 ps=0 
M2381 n_1117 n_70 GND GND efet w=45 l=6
+ ad=0 pd=0 as=0 ps=0 
M2382 GND pipeVectorA1 n_0_ADL1 GND efet w=94 l=7
+ ad=0 pd=0 as=1034 ps=316 
M2383 Vdd n_0_ADL1 n_0_ADL1 GND dfet w=9 l=16
+ ad=0 pd=0 as=3501 ps=1242 
M2384 Vdd n_0_ADL2 n_0_ADL2 GND dfet w=9 l=15
+ ad=0 pd=0 as=4670 ps=1736 
M2385 GND n_815 n_0_ADL2 GND efet w=51 l=6
+ ad=0 pd=0 as=665 ps=168 
M2386 n_696 cclk n_610 GND efet w=12 l=10
+ ad=0 pd=0 as=220 ps=80 
M2387 n_1101 cclk n_190 GND efet w=12 l=8
+ ad=1182 pd=334 as=178 ps=62 
M2388 n_1717 cclk n_1113 GND efet w=12 l=9
+ ad=0 pd=0 as=123 ps=58 
M2389 Vdd n_582 n_582 GND dfet w=9 l=10
+ ad=0 pd=0 as=1321 ps=400 
M2390 GND n_610 n_582 GND efet w=71 l=6
+ ad=0 pd=0 as=854 ps=200 
M2391 GND cp1 n_43 GND efet w=206 l=7
+ ad=0 pd=0 as=2534 ps=556 
M2392 n_43 n_839 Vdd GND dfet w=42 l=7
+ ad=0 pd=0 as=0 ps=0 
M2393 GND cp1 n_43 GND efet w=126 l=6
+ ad=0 pd=0 as=0 ps=0 
M2394 Vdd n_220 n_220 GND dfet w=9 l=10
+ ad=0 pd=0 as=1298 ps=390 
M2395 GND n_190 n_220 GND efet w=70 l=6
+ ad=0 pd=0 as=823 ps=198 
M2396 n_161 n_1113 GND GND efet w=57 l=6
+ ad=813 pd=214 as=0 ps=0 
M2397 Vdd n_161 n_161 GND dfet w=10 l=12
+ ad=0 pd=0 as=1033 ps=328 
M2398 n_1106 cclk n_1404 GND efet w=12 l=10
+ ad=0 pd=0 as=125 ps=66 
M2399 n_133 n_133 Vdd GND dfet w=8 l=11
+ ad=1097 pd=324 as=0 ps=0 
M2400 GND n_1404 n_133 GND efet w=60 l=5
+ ad=0 pd=0 as=825 ps=230 
M2401 GND cp1 n_1247 GND efet w=104 l=6
+ ad=0 pd=0 as=2764 ps=672 
M2402 testpad_5 n_1127 testpad_5 GND efet w=84 l=73
+ ad=5355 pd=642 as=0 ps=0 
M2403 testpad_1 n_1127 testpad_1 GND efet w=63 l=68
+ ad=2825 pd=328 as=0 ps=0 
M2404 testpad_2 testpad_4 testpad_5 GND efet w=10 l=6
+ ad=8375 pd=516 as=0 ps=0 
M2405 n_1247 cp1 GND GND efet w=209 l=7
+ ad=0 pd=0 as=0 ps=0 
M2406 GND cp1 n_1247 GND efet w=180 l=6
+ ad=0 pd=0 as=0 ps=0 
M2407 n_1247 n_38 Vdd GND dfet w=64 l=7
+ ad=0 pd=0 as=0 ps=0 
M2408 n_839 n_839 Vdd GND dfet w=13 l=7
+ ad=938 pd=282 as=0 ps=0 
M2409 GND cp1 n_839 GND efet w=63 l=7
+ ad=0 pd=0 as=602 ps=172 
M2410 n_1067 n_582 GND GND efet w=25 l=7
+ ad=322 pd=102 as=0 ps=0 
M2411 n_130 n_220 GND GND efet w=26 l=7
+ ad=347 pd=104 as=0 ps=0 
M2412 GND cclk n_161 GND efet w=25 l=6
+ ad=0 pd=0 as=0 ps=0 
M2413 n_133 cclk GND GND efet w=25 l=6
+ ad=0 pd=0 as=0 ps=0 
M2414 n_969 n_161 GND GND efet w=25 l=6
+ ad=343 pd=90 as=0 ps=0 
M2415 n_1067 n_1067 Vdd GND dfet w=10 l=13
+ ad=1495 pd=474 as=0 ps=0 
M2416 Vdd n_582 ADH_ABH GND dfet w=12 l=8
+ ad=0 pd=0 as=1735 ps=378 
M2417 n_130 n_130 Vdd GND dfet w=11 l=14
+ ad=1233 pd=360 as=0 ps=0 
M2418 n_38 cp1 GND GND efet w=55 l=6
+ ad=543 pd=168 as=0 ps=0 
M2419 Vdd n_38 n_38 GND dfet w=14 l=7
+ ad=0 pd=0 as=1139 ps=366 
M2420 GND n_1067 ADH_ABH GND efet w=149 l=6
+ ad=0 pd=0 as=0 ps=0 
M2421 Vdd n_220 ADL_ABL GND dfet w=9 l=8
+ ad=0 pd=0 as=1282 ps=306 
M2422 Vdd n_969 n_969 GND dfet w=10 l=12
+ ad=0 pd=0 as=1187 ps=358 
M2423 testpad_5 diff_237_1656# n_1701 GND efet w=11 l=42
+ ad=0 pd=0 as=1452 ps=242 
M2424 testpad_6 diff_237_1656# n_1701 GND efet w=10 l=6
+ ad=848 pd=128 as=0 ps=0 
M2425 testpad_2 testpad_4 testpad_6 GND efet w=38 l=6
+ ad=0 pd=0 as=0 ps=0 
M2426 GND n_130 ADL_ABL GND efet w=97 l=6
+ ad=0 pd=0 as=0 ps=0 
M2427 Vdd n_161 dpc0_YSB GND dfet w=11 l=8
+ ad=0 pd=0 as=1642 ps=322 
M2428 GND n_133 n_602 GND efet w=25 l=7
+ ad=0 pd=0 as=372 ps=108 
M2429 n_602 n_602 Vdd GND dfet w=10 l=11
+ ad=1133 pd=386 as=0 ps=0 
M2430 Vdd n_133 dpc2_XSB GND dfet w=10 l=8
+ ad=0 pd=0 as=1756 ps=362 
M2431 dpc0_YSB n_1247 GND GND efet w=74 l=6
+ ad=0 pd=0 as=0 ps=0 
M2432 GND n_969 dpc0_YSB GND efet w=77 l=6
+ ad=0 pd=0 as=0 ps=0 
M2433 dpc2_XSB n_602 GND GND efet w=92 l=6
+ ad=0 pd=0 as=0 ps=0 
M2434 GND n_1247 dpc2_XSB GND efet w=91 l=5
+ ad=0 pd=0 as=0 ps=0 
M2435 ab0 n_1100 GND GND efet w=443 l=7
+ ad=14563 pd=2238 as=0 ps=0 
M2436 ab0 n_1100 GND GND efet w=352 l=6
+ ad=0 pd=0 as=0 ps=0 
M2437 ab0 n_1100 GND GND efet w=170 l=7
+ ad=0 pd=0 as=0 ps=0 
M2438 Vdd n_855 ab0 GND efet w=68 l=7
+ ad=0 pd=0 as=0 ps=0 
M2439 Vdd n_855 ab0 GND efet w=239 l=6
+ ad=0 pd=0 as=0 ps=0 
M2440 GND n_1660 n_855 GND efet w=126 l=7
+ ad=0 pd=0 as=1564 ps=378 
M2441 Vdd n_855 ab0 GND efet w=238 l=6
+ ad=0 pd=0 as=0 ps=0 
M2442 Vdd n_855 ab0 GND efet w=240 l=7
+ ad=0 pd=0 as=0 ps=0 
M2443 n_1660 abl0 GND GND efet w=36 l=8
+ ad=466 pd=140 as=0 ps=0 
M2444 n_1660 n_1660 Vdd GND dfet w=10 l=10
+ ad=1792 pd=532 as=0 ps=0 
M2445 GND abl0 n_1100 GND efet w=154 l=7
+ ad=0 pd=0 as=1503 ps=400 
M2446 n_855 abl0 Vdd GND dfet w=18 l=7
+ ad=0 pd=0 as=0 ps=0 
M2447 n_1100 n_1660 Vdd GND dfet w=21 l=7
+ ad=0 pd=0 as=0 ps=0 
M2448 n_629 n_50 GND GND efet w=40 l=7
+ ad=0 pd=0 as=0 ps=0 
M2449 n_50 cp1 INTG GND efet w=12 l=9
+ ad=141 pd=60 as=1383 ps=372 
M2450 Vdd n_152 n_152 GND dfet w=9 l=12
+ ad=0 pd=0 as=1577 ps=530 
M2451 n_152 n_1002 GND GND efet w=29 l=6
+ ad=1244 pd=284 as=0 ps=0 
M2452 n_1178 pipeUNK30 GND GND efet w=54 l=6
+ ad=0 pd=0 as=0 ps=0 
M2453 n_389 cclk pipeUNK31 GND efet w=11 l=7
+ ad=0 pd=0 as=185 ps=76 
M2454 n_1178 pipeUNK32 GND GND efet w=54 l=6
+ ad=0 pd=0 as=0 ps=0 
M2455 GND pipeUNK33 n_1178 GND efet w=50 l=6
+ ad=0 pd=0 as=0 ps=0 
M2456 n_1081 cclk pipeUNK32 GND efet w=12 l=7
+ ad=1011 pd=292 as=279 ps=68 
M2457 n_473 cclk pipeUNK33 GND efet w=13 l=7
+ ad=1040 pd=258 as=206 ps=84 
M2458 Vdd n_1081 n_1081 GND dfet w=9 l=13
+ ad=0 pd=0 as=2885 ps=1060 
M2459 n_1081 n_1560 GND GND efet w=38 l=6
+ ad=0 pd=0 as=0 ps=0 
M2460 n_300 n_389 GND GND efet w=31 l=7
+ ad=0 pd=0 as=0 ps=0 
M2461 Vdd n_1130 n_1130 GND dfet w=10 l=13
+ ad=0 pd=0 as=5560 ps=1964 
M2462 n_1130 n_1109 GND GND efet w=30 l=7
+ ad=2255 pd=636 as=0 ps=0 
M2463 GND n_1258 n_1130 GND efet w=42 l=6
+ ad=0 pd=0 as=0 ps=0 
M2464 n_1130 n_862 GND GND efet w=29 l=6
+ ad=0 pd=0 as=0 ps=0 
M2465 GND n_192 n_1130 GND efet w=28 l=7
+ ad=0 pd=0 as=0 ps=0 
M2466 n_847 n_300 GND GND efet w=37 l=6
+ ad=717 pd=202 as=0 ps=0 
M2467 GND op_T2 n_152 GND efet w=41 l=6
+ ad=0 pd=0 as=0 ps=0 
M2468 n_256 op_T5_rti GND GND efet w=31 l=6
+ ad=2295 pd=680 as=0 ps=0 
M2469 n_152 n_952 GND GND efet w=28 l=7
+ ad=0 pd=0 as=0 ps=0 
M2470 GND n_630 n_152 GND efet w=45 l=6
+ ad=0 pd=0 as=0 ps=0 
M2471 Vdd op_EORS op_EORS GND dfet w=10 l=17
+ ad=0 pd=0 as=2936 ps=918 
M2472 op_EORS n_837 GND GND efet w=37 l=6
+ ad=756 pd=202 as=0 ps=0 
M2473 n_372 notRdy0 GND GND efet w=29 l=7
+ ad=346 pd=98 as=0 ps=0 
M2474 n_372 n_372 Vdd GND dfet w=10 l=12
+ ad=988 pd=312 as=0 ps=0 
M2475 n_847 n_847 Vdd GND dfet w=9 l=11
+ ad=774 pd=238 as=0 ps=0 
M2476 n_1408 n_1044 n_1000 GND efet w=56 l=6
+ ad=472 pd=144 as=0 ps=0 
M2477 n_980 n_980 Vdd GND dfet w=9 l=16
+ ad=2157 pd=696 as=0 ps=0 
M2478 Vdd n_1408 n_1408 GND dfet w=9 l=17
+ ad=0 pd=0 as=1787 ps=594 
M2479 n_104 n_847 GND GND efet w=35 l=7
+ ad=3147 pd=778 as=0 ps=0 
M2480 n_1130 n_1002 GND GND efet w=33 l=6
+ ad=0 pd=0 as=0 ps=0 
M2481 n_1365 n_862 GND GND efet w=40 l=5
+ ad=240 pd=92 as=0 ps=0 
M2482 n_1085 notRdy0 n_1365 GND efet w=40 l=7
+ ad=1360 pd=364 as=0 ps=0 
M2483 n_911 n_877 GND GND efet w=22 l=7
+ ad=0 pd=0 as=0 ps=0 
M2484 GND n_1343 n_911 GND efet w=97 l=6
+ ad=0 pd=0 as=0 ps=0 
M2485 n_911 n_877 GND GND efet w=61 l=6
+ ad=0 pd=0 as=0 ps=0 
M2486 n_1172 n_372 n_1085 GND efet w=55 l=6
+ ad=1249 pd=248 as=0 ps=0 
M2487 n_405 BRtaken n_1172 GND efet w=55 l=7
+ ad=550 pd=130 as=0 ps=0 
M2488 GND nnT2BR n_405 GND efet w=55 l=7
+ ad=0 pd=0 as=0 ps=0 
M2489 n_1343 n_152 GND GND efet w=30 l=7
+ ad=677 pd=196 as=0 ps=0 
M2490 GND notRdy0 n_1343 GND efet w=30 l=6
+ ad=0 pd=0 as=0 ps=0 
M2491 Vdd n_1085 n_1085 GND dfet w=9 l=17
+ ad=0 pd=0 as=849 ps=260 
M2492 n_79 n_236 GND GND efet w=91 l=6
+ ad=1160 pd=304 as=0 ps=0 
M2493 GND n_646 n_1172 GND efet w=36 l=7
+ ad=0 pd=0 as=0 ps=0 
M2494 n_1343 n_1343 Vdd GND dfet w=8 l=12
+ ad=989 pd=290 as=0 ps=0 
M2495 n_629 cclk n_760 GND efet w=11 l=9
+ ad=0 pd=0 as=371 ps=112 
M2496 D1x1 D1x1 Vdd GND dfet w=9 l=8
+ ad=8548 pd=3088 as=0 ps=0 
M2497 Vdd n_1594 n_1594 GND dfet w=9 l=13
+ ad=0 pd=0 as=1029 ps=366 
M2498 GND n_1358 n_396 GND efet w=29 l=7
+ ad=0 pd=0 as=544 ps=188 
M2499 INTG brk_done GND GND efet w=25 l=5
+ ad=0 pd=0 as=0 ps=0 
M2500 GND n_760 INTG GND efet w=44 l=6
+ ad=0 pd=0 as=0 ps=0 
M2501 D1x1 C1x5Reset GND GND efet w=62 l=5
+ ad=1529 pd=352 as=0 ps=0 
M2502 GND INTG D1x1 GND efet w=64 l=7
+ ad=0 pd=0 as=0 ps=0 
M2503 n_79 n_79 Vdd GND dfet w=10 l=9
+ ad=1454 pd=442 as=0 ps=0 
M2504 n_656 n_779 n_1594 GND efet w=54 l=7
+ ad=270 pd=118 as=760 ps=256 
M2505 GND n_604 n_656 GND efet w=54 l=7
+ ad=0 pd=0 as=0 ps=0 
M2506 n_795 n_1649 GND GND efet w=29 l=7
+ ad=529 pd=196 as=0 ps=0 
M2507 Vdd n_795 n_795 GND dfet w=9 l=12
+ ad=0 pd=0 as=707 ps=238 
M2508 n_396 n_396 Vdd GND dfet w=10 l=11
+ ad=485 pd=142 as=0 ps=0 
M2509 n_616 cclk n_460 GND efet w=12 l=9
+ ad=0 pd=0 as=140 ps=76 
M2510 n_844 cclk n_459 GND efet w=13 l=9
+ ad=0 pd=0 as=148 ps=78 
M2511 n_1586 cclk n_621 GND efet w=11 l=9
+ ad=0 pd=0 as=159 ps=76 
M2512 n_632 cclk n_339 GND efet w=12 l=10
+ ad=0 pd=0 as=155 ps=58 
M2513 n_1358 cclk n_521 GND efet w=13 l=10
+ ad=0 pd=0 as=148 ps=70 
M2514 INTG INTG Vdd GND dfet w=10 l=16
+ ad=2288 pd=794 as=0 ps=0 
M2515 n_1304 op_T0_sbc GND GND efet w=47 l=6
+ ad=796 pd=184 as=0 ps=0 
M2516 GND n_673 n_1304 GND efet w=39 l=7
+ ad=0 pd=0 as=0 ps=0 
M2517 n_1304 n_1304 Vdd GND dfet w=10 l=13
+ ad=1448 pd=476 as=0 ps=0 
M2518 n_605 n_1081 GND GND efet w=81 l=6
+ ad=1768 pd=522 as=0 ps=0 
M2519 GND op_T0_sbc n_605 GND efet w=81 l=6
+ ad=0 pd=0 as=0 ps=0 
M2520 GND clock2 op_T__bit GND efet w=13 l=7
+ ad=0 pd=0 as=0 ps=0 
M2521 GND clock2 x_op_T__adc_sbc GND efet w=15 l=8
+ ad=0 pd=0 as=0 ps=0 
M2522 GND clock2 op_T__cmp GND efet w=13 l=7
+ ad=0 pd=0 as=0 ps=0 
M2523 GND clock2 op_T__cpx_cpy_abs GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M2524 GND clock2 op_T__asl_rol_a GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M2525 notir5 notir5 Vdd GND dfet w=10 l=6
+ ad=22059 pd=7174 as=0 ps=0 
M2526 GND ir5 notir5 GND efet w=93 l=7
+ ad=0 pd=0 as=2097 ps=464 
M2527 GND clock2 op_T__cpx_cpy_imm_zp GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M2528 n_1378 fetch n_1609 GND efet w=23 l=8
+ ad=115 pd=56 as=435 ps=108 
M2529 n_928 cp1 n_1378 GND efet w=23 l=10
+ ad=1603 pd=390 as=0 ps=0 
M2530 n_1609 cclk notir5 GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M2531 n_1455 op_T0_tya GND GND efet w=37 l=7
+ ad=2536 pd=626 as=0 ps=0 
M2532 n_1455 n_1455 Vdd GND dfet w=9 l=17
+ ad=7631 pd=2644 as=0 ps=0 
M2533 n_1455 op_T__shift_a GND GND efet w=38 l=7
+ ad=0 pd=0 as=0 ps=0 
M2534 GND op_T0_txa n_1455 GND efet w=30 l=7
+ ad=0 pd=0 as=0 ps=0 
M2535 n_1455 op_T0_pla GND GND efet w=29 l=7
+ ad=0 pd=0 as=0 ps=0 
M2536 GND op_T0_lda n_1455 GND efet w=29 l=7
+ ad=0 pd=0 as=0 ps=0 
M2537 n_1563 op_T0_acc GND GND efet w=51 l=7
+ ad=253 pd=112 as=0 ps=0 
M2538 n_11 n_397 n_1563 GND efet w=51 l=7
+ ad=2067 pd=628 as=0 ps=0 
M2539 GND op_T0_tay n_11 GND efet w=35 l=6
+ ad=0 pd=0 as=0 ps=0 
M2540 n_11 op_T0_shift_a GND GND efet w=40 l=5
+ ad=0 pd=0 as=0 ps=0 
M2541 GND op_T__adc_sbc n_1455 GND efet w=35 l=7
+ ad=0 pd=0 as=0 ps=0 
M2542 GND op_T__ora_and_eor_adc n_1455 GND efet w=31 l=7
+ ad=0 pd=0 as=0 ps=0 
M2543 GND op_T0_lda n_397 GND efet w=33 l=6
+ ad=0 pd=0 as=641 ps=176 
M2544 GND op_T0_tax n_11 GND efet w=42 l=7
+ ad=0 pd=0 as=0 ps=0 
M2545 n_669 op_T0_bit GND GND efet w=42 l=7
+ ad=525 pd=176 as=0 ps=0 
M2546 Vdd n_397 n_397 GND dfet w=9 l=13
+ ad=0 pd=0 as=814 ps=224 
M2547 Vdd n_1090 n_1090 GND dfet w=9 l=12
+ ad=0 pd=0 as=5604 ps=2082 
M2548 n_1681 n_440 n_905 GND efet w=52 l=7
+ ad=273 pd=114 as=560 ps=164 
M2549 GND op_shift n_1681 GND efet w=52 l=7
+ ad=0 pd=0 as=0 ps=0 
M2550 Vdd n_384 n_384 GND dfet w=9 l=13
+ ad=0 pd=0 as=1135 ps=342 
M2551 Vdd n_1412 n_1412 GND dfet w=9 l=12
+ ad=0 pd=0 as=633 ps=198 
M2552 GND n_1222 n_1090 GND efet w=37 l=7
+ ad=0 pd=0 as=1411 ps=400 
M2553 n_1090 op_T2_stack_access GND GND efet w=39 l=7
+ ad=0 pd=0 as=0 ps=0 
M2554 n_1222 n_1225 GND GND efet w=43 l=7
+ ad=727 pd=228 as=0 ps=0 
M2555 n_905 n_905 Vdd GND dfet w=10 l=16
+ ad=652 pd=180 as=0 ps=0 
M2556 GND op_T0_and n_669 GND efet w=30 l=7
+ ad=0 pd=0 as=0 ps=0 
M2557 n_595 op_T4_abs_idx GND GND efet w=53 l=7
+ ad=760 pd=194 as=0 ps=0 
M2558 GND op_T5_ind_y n_595 GND efet w=37 l=6
+ ad=0 pd=0 as=0 ps=0 
M2559 nop_branch_done op_branch_done GND GND efet w=37 l=7
+ ad=505 pd=164 as=0 ps=0 
M2560 n_11 n_11 Vdd GND dfet w=9 l=16
+ ad=6988 pd=2392 as=0 ps=0 
M2561 n_669 n_669 Vdd GND dfet w=9 l=16
+ ad=908 pd=262 as=0 ps=0 
M2562 n_595 n_595 Vdd GND dfet w=9 l=13
+ ad=1423 pd=454 as=0 ps=0 
M2563 GND n_1412 n_384 GND efet w=34 l=6
+ ad=0 pd=0 as=2542 ps=590 
M2564 Vdd op_ANDS op_ANDS GND dfet w=10 l=16
+ ad=0 pd=0 as=6913 ps=2392 
M2565 nop_branch_done nop_branch_done Vdd GND dfet w=10 l=16
+ ad=872 pd=240 as=0 ps=0 
M2566 n_366 op_T0_shift_right_a GND GND efet w=49 l=6
+ ad=944 pd=264 as=0 ps=0 
M2567 n_1012 n_440 n_366 GND efet w=56 l=6
+ ad=362 pd=138 as=0 ps=0 
M2568 GND op_shift_right n_1012 GND efet w=59 l=6
+ ad=0 pd=0 as=0 ps=0 
M2569 n_824 op_T2_brk GND GND efet w=36 l=6
+ ad=1286 pd=358 as=0 ps=0 
M2570 GND op_T3_jsr n_824 GND efet w=40 l=7
+ ad=0 pd=0 as=0 ps=0 
M2571 GND op_ANDS n_11 GND efet w=39 l=6
+ ad=0 pd=0 as=0 ps=0 
M2572 Vdd n_1037 n_1037 GND dfet w=9 l=16
+ ad=0 pd=0 as=6831 ps=2252 
M2573 Vdd n_366 n_366 GND dfet w=10 l=11
+ ad=0 pd=0 as=676 ps=218 
M2574 n_1222 n_1222 Vdd GND dfet w=10 l=12
+ ad=795 pd=228 as=0 ps=0 
M2575 GND n_946 n_384 GND efet w=28 l=7
+ ad=0 pd=0 as=0 ps=0 
M2576 GND n_1455 n_1412 GND efet w=43 l=6
+ ad=0 pd=0 as=586 ps=152 
M2577 n_1347 op_T0_shift_a GND GND efet w=46 l=7
+ ad=2959 pd=798 as=0 ps=0 
M2578 GND n_905 n_979 GND efet w=27 l=6
+ ad=0 pd=0 as=452 ps=134 
M2579 n_979 n_979 Vdd GND dfet w=9 l=17
+ ad=704 pd=202 as=0 ps=0 
M2580 Vdd n_473 n_473 GND dfet w=9 l=13
+ ad=0 pd=0 as=1776 ps=662 
M2581 n_1004 n_1408 GND GND efet w=71 l=6
+ ad=389 pd=154 as=0 ps=0 
M2582 n_473 n_980 n_1004 GND efet w=71 l=6
+ ad=0 pd=0 as=0 ps=0 
M2583 n_1347 n_979 GND GND efet w=29 l=7
+ ad=0 pd=0 as=0 ps=0 
M2584 GND op_T5_jsr n_1219 GND efet w=26 l=6
+ ad=0 pd=0 as=400 ps=106 
M2585 n_1347 n_782 GND GND efet w=28 l=7
+ ad=0 pd=0 as=0 ps=0 
M2586 GND n_1219 n_1002 GND efet w=45 l=6
+ ad=0 pd=0 as=645 ps=168 
M2587 n_1219 n_1219 Vdd GND dfet w=10 l=17
+ ad=836 pd=236 as=0 ps=0 
M2588 n_1347 n_862 GND GND efet w=36 l=7
+ ad=0 pd=0 as=0 ps=0 
M2589 n_384 n_1258 GND GND efet w=39 l=7
+ ad=0 pd=0 as=0 ps=0 
M2590 GND n_550 n_1347 GND efet w=35 l=6
+ ad=0 pd=0 as=0 ps=0 
M2591 n_384 op_ANDS GND GND efet w=17 l=6
+ ad=0 pd=0 as=0 ps=0 
M2592 GND op_ANDS n_550 GND efet w=38 l=6
+ ad=0 pd=0 as=1004 ps=252 
M2593 n_384 op_ANDS GND GND efet w=20 l=7
+ ad=0 pd=0 as=0 ps=0 
M2594 n_1347 n_1347 Vdd GND dfet w=8 l=13
+ ad=5510 pd=1920 as=0 ps=0 
M2595 Vdd n_506 n_506 GND dfet w=8 l=11
+ ad=0 pd=0 as=5964 ps=2028 
M2596 GND n_669 op_ANDS GND efet w=51 l=7
+ ad=0 pd=0 as=689 ps=208 
M2597 GND n_192 n_506 GND efet w=38 l=6
+ ad=0 pd=0 as=1143 ps=352 
M2598 GND n_1258 n_813 GND efet w=36 l=7
+ ad=0 pd=0 as=822 ps=232 
M2599 n_1002 n_1002 Vdd GND dfet w=9 l=10
+ ad=3455 pd=1176 as=0 ps=0 
M2600 Vdd n_673 n_673 GND dfet w=10 l=13
+ ad=0 pd=0 as=1142 ps=336 
M2601 n_1053 op_T0_adc_sbc n_673 GND efet w=66 l=6
+ ad=474 pd=170 as=539 ps=170 
M2602 GND n_1002 n_605 GND efet w=36 l=6
+ ad=0 pd=0 as=0 ps=0 
M2603 n_605 n_1002 GND GND efet w=31 l=6
+ ad=0 pd=0 as=0 ps=0 
M2604 n_779 n_1440 n_605 GND efet w=62 l=6
+ ad=867 pd=250 as=0 ps=0 
M2605 GND Pout3 n_1053 GND efet w=59 l=6
+ ad=0 pd=0 as=0 ps=0 
M2606 Vdd n_25 n_25 GND dfet w=9 l=12
+ ad=0 pd=0 as=4084 ps=1362 
M2607 n_25 n_192 GND GND efet w=44 l=6
+ ad=898 pd=224 as=0 ps=0 
M2608 Vdd n_1440 n_1440 GND dfet w=9 l=12
+ ad=0 pd=0 as=1068 ps=338 
M2609 n_779 n_779 Vdd GND dfet w=8 l=15
+ ad=4280 pd=1396 as=0 ps=0 
M2610 GND n_384 n_550 GND efet w=32 l=7
+ ad=0 pd=0 as=0 ps=0 
M2611 n_885 n_384 GND GND efet w=46 l=7
+ ad=555 pd=196 as=0 ps=0 
M2612 n_813 n_440 GND GND efet w=35 l=7
+ ad=0 pd=0 as=0 ps=0 
M2613 GND n_595 n_992 GND efet w=33 l=6
+ ad=0 pd=0 as=549 ps=156 
M2614 n_239 n_595 GND GND efet w=49 l=7
+ ad=245 pd=108 as=0 ps=0 
M2615 n_192 nop_branch_done n_239 GND efet w=49 l=7
+ ad=776 pd=206 as=0 ps=0 
M2616 GND n_992 n_46 GND efet w=45 l=6
+ ad=0 pd=0 as=934 ps=250 
M2617 n_813 n_813 Vdd GND dfet w=10 l=18
+ ad=1306 pd=340 as=0 ps=0 
M2618 n_992 n_992 Vdd GND dfet w=10 l=13
+ ad=810 pd=240 as=0 ps=0 
M2619 Vdd n_1101 n_1101 GND dfet w=9 l=11
+ ad=0 pd=0 as=5873 ps=1936 
M2620 n_192 n_192 Vdd GND dfet w=9 l=13
+ ad=4832 pd=1650 as=0 ps=0 
M2621 Vdd n_46 n_46 GND dfet w=9 l=17
+ ad=0 pd=0 as=1200 ps=372 
M2622 GND notRdy0 n_46 GND efet w=51 l=7
+ ad=0 pd=0 as=0 ps=0 
M2623 n_550 n_550 Vdd GND dfet w=8 l=13
+ ad=994 pd=312 as=0 ps=0 
M2624 n_885 n_885 Vdd GND dfet w=9 l=11
+ ad=4576 pd=1528 as=0 ps=0 
M2625 n_1508 n_813 n_1101 GND efet w=86 l=7
+ ad=821 pd=228 as=0 ps=0 
M2626 GND n_334 n_118 GND efet w=43 l=7
+ ad=0 pd=0 as=623 ps=170 
M2627 n_1688 n_1304 GND GND efet w=31 l=7
+ ad=867 pd=242 as=0 ps=0 
M2628 n_118 n_118 Vdd GND dfet w=10 l=10
+ ad=1109 pd=354 as=0 ps=0 
M2629 n_1688 n_1688 Vdd GND dfet w=9 l=12
+ ad=2773 pd=920 as=0 ps=0 
M2630 n_1440 notRdy0 GND GND efet w=36 l=6
+ ad=278 pd=84 as=0 ps=0 
M2631 n_25 n_256 GND GND efet w=28 l=7
+ ad=0 pd=0 as=0 ps=0 
M2632 n_51 Pout3 GND GND efet w=62 l=6
+ ad=310 pd=134 as=0 ps=0 
M2633 n_29 op_T0_sbc n_51 GND efet w=62 l=6
+ ad=1171 pd=320 as=0 ps=0 
M2634 Vdd n_29 n_29 GND dfet w=9 l=14
+ ad=0 pd=0 as=456 ps=124 
M2635 n_819 pipephi2Reset0 GND GND efet w=67 l=7
+ ad=1260 pd=254 as=0 ps=0 
M2636 GND pipeUNK23 n_819 GND efet w=80 l=7
+ ad=0 pd=0 as=0 ps=0 
M2637 n_334 brk_done GND GND efet w=45 l=6
+ ad=2314 pd=662 as=0 ps=0 
M2638 n_533 pipeUNK22 GND GND efet w=44 l=7
+ ad=808 pd=238 as=0 ps=0 
M2639 pipeUNK22 cclk n_29 GND efet w=13 l=8
+ ad=231 pd=80 as=0 ps=0 
M2640 n_1347 nnT2BR GND GND efet w=31 l=7
+ ad=0 pd=0 as=0 ps=0 
M2641 GND n_223 n_1357 GND efet w=136 l=7
+ ad=0 pd=0 as=1803 ps=390 
M2642 n_223 cp1 n_1215 GND efet w=12 l=8
+ ad=174 pd=74 as=3489 ps=816 
M2643 n_1357 n_1357 Vdd GND dfet w=10 l=8
+ ad=6107 pd=2008 as=0 ps=0 
M2644 n_104 nnT2BR GND GND efet w=49 l=6
+ ad=0 pd=0 as=0 ps=0 
M2645 pipephi2Reset0 cclk Reset0 GND efet w=12 l=8
+ ad=140 pd=58 as=0 ps=0 
M2646 Vdd n_819 n_819 GND dfet w=9 l=10
+ ad=0 pd=0 as=4692 ps=1604 
M2647 n_533 n_533 Vdd GND dfet w=9 l=19
+ ad=1662 pd=530 as=0 ps=0 
M2648 pipeUNK23 cclk n_1085 GND efet w=13 l=9
+ ad=144 pd=66 as=0 ps=0 
M2649 n_590 cp1 n_1178 GND efet w=12 l=7
+ ad=192 pd=80 as=0 ps=0 
M2650 GND op_ANDS op_SUMS GND efet w=28 l=7
+ ad=0 pd=0 as=1421 ps=364 
M2651 op_SUMS op_EORS GND GND efet w=29 l=7
+ ad=0 pd=0 as=0 ps=0 
M2652 GND op_ORS op_SUMS GND efet w=45 l=6
+ ad=0 pd=0 as=0 ps=0 
M2653 op_SUMS op_SUMS Vdd GND dfet w=9 l=15
+ ad=304 pd=82 as=0 ps=0 
M2654 op_ANDS cclk n_1574 GND efet w=12 l=8
+ ad=0 pd=0 as=164 ps=78 
M2655 n_796 cclk n_396 GND efet w=12 l=9
+ ad=126 pd=68 as=0 ps=0 
M2656 GND n_590 alucin GND efet w=68 l=6
+ ad=0 pd=0 as=685 ps=220 
M2657 op_SUMS op_SRS GND GND efet w=33 l=6
+ ad=0 pd=0 as=0 ps=0 
M2658 notRdy0 cp1 n_1679 GND efet w=12 l=7
+ ad=0 pd=0 as=198 ps=78 
M2659 n_1262 n_1679 GND GND efet w=44 l=7
+ ad=786 pd=204 as=0 ps=0 
M2660 GND n_236 n_506 GND efet w=38 l=6
+ ad=0 pd=0 as=0 ps=0 
M2661 GND n_46 n_1508 GND efet w=96 l=6
+ ad=0 pd=0 as=0 ps=0 
M2662 GND op_T2_pha n_1037 GND efet w=35 l=6
+ ad=0 pd=0 as=1905 ps=506 
M2663 n_824 n_824 Vdd GND dfet w=10 l=15
+ ad=8959 pd=2948 as=0 ps=0 
M2664 Vdd op_SRS op_SRS GND dfet w=9 l=11
+ ad=0 pd=0 as=11360 ps=4024 
M2665 op_SRS n_366 GND GND efet w=33 l=6
+ ad=0 pd=0 as=0 ps=0 
M2666 n_1280 op_sta_cmp n_1037 GND efet w=54 l=6
+ ad=395 pd=126 as=0 ps=0 
M2667 GND n_335 n_1280 GND efet w=56 l=6
+ ad=0 pd=0 as=0 ps=0 
M2668 n_1225 op_T2_ind GND GND efet w=45 l=6
+ ad=1699 pd=598 as=0 ps=0 
M2669 n_272 op_T2_abs_access GND GND efet w=54 l=7
+ ad=2232 pd=742 as=0 ps=0 
M2670 GND op_T5_rts n_272 GND efet w=36 l=7
+ ad=0 pd=0 as=0 ps=0 
M2671 n_256 op_T4 GND GND efet w=45 l=6
+ ad=0 pd=0 as=0 ps=0 
M2672 GND op_T3 n_256 GND efet w=41 l=7
+ ad=0 pd=0 as=0 ps=0 
M2673 n_726 op_T5_ind_x GND GND efet w=42 l=6
+ ad=1572 pd=502 as=0 ps=0 
M2674 n_256 op_T0_brk_rti GND GND efet w=43 l=7
+ ad=0 pd=0 as=0 ps=0 
M2675 n_1225 n_1225 Vdd GND dfet w=10 l=9
+ ad=12615 pd=4282 as=0 ps=0 
M2676 n_272 n_272 Vdd GND dfet w=9 l=13
+ ad=7941 pd=2612 as=0 ps=0 
M2677 GND op_T2_zp_zp_idx n_1225 GND efet w=64 l=7
+ ad=0 pd=0 as=0 ps=0 
M2678 n_636 op_T2_branch GND GND efet w=25 l=7
+ ad=516 pd=156 as=0 ps=0 
M2679 n_256 op_T5_rts GND GND efet w=35 l=7
+ ad=0 pd=0 as=0 ps=0 
M2680 GND op_T0_jmp n_256 GND efet w=42 l=6
+ ad=0 pd=0 as=0 ps=0 
M2681 GND op_T3_abs_idx_ind n_726 GND efet w=38 l=6
+ ad=0 pd=0 as=0 ps=0 
M2682 n_256 op_T5_ind_x GND GND efet w=38 l=6
+ ad=0 pd=0 as=0 ps=0 
M2683 n_726 n_726 Vdd GND dfet w=9 l=13
+ ad=1344 pd=460 as=0 ps=0 
M2684 n_256 n_256 Vdd GND dfet w=10 l=15
+ ad=4505 pd=1638 as=0 ps=0 
M2685 GND Reset0 n_501 GND efet w=55 l=6
+ ad=0 pd=0 as=1915 ps=526 
M2686 pipeUNK34 cclk n_824 GND efet w=11 l=8
+ ad=162 pd=76 as=0 ps=0 
M2687 n_1215 brk_done GND GND efet w=160 l=6
+ ad=0 pd=0 as=0 ps=0 
M2688 n_272 n_236 GND GND efet w=31 l=7
+ ad=0 pd=0 as=0 ps=0 
M2689 n_720 pipeUNK34 GND GND efet w=69 l=6
+ ad=1722 pd=446 as=0 ps=0 
M2690 n_636 n_636 Vdd GND dfet w=10 l=16
+ ad=1250 pd=396 as=0 ps=0 
M2691 GND pipeUNK35 n_238 GND efet w=59 l=6
+ ad=0 pd=0 as=972 ps=284 
M2692 n_261 x_op_T4_ind_y GND GND efet w=36 l=6
+ ad=644 pd=246 as=0 ps=0 
M2693 GND x_op_T3_abs_idx n_261 GND efet w=38 l=7
+ ad=0 pd=0 as=0 ps=0 
M2694 n_726 x_op_T4_ind_y GND GND efet w=37 l=6
+ ad=0 pd=0 as=0 ps=0 
M2695 n_134 op_brk_rti GND GND efet w=38 l=7
+ ad=1124 pd=256 as=0 ps=0 
M2696 GND op_jsr n_134 GND efet w=27 l=6
+ ad=0 pd=0 as=0 ps=0 
M2697 n_261 n_261 Vdd GND dfet w=10 l=14
+ ad=1342 pd=464 as=0 ps=0 
M2698 n_501 cclk pipeUNK35 GND efet w=11 l=7
+ ad=0 pd=0 as=138 ps=58 
M2699 n_726 op_T5_rts GND GND efet w=33 l=7
+ ad=0 pd=0 as=0 ps=0 
M2700 n_238 n_238 Vdd GND dfet w=10 l=16
+ ad=1834 pd=570 as=0 ps=0 
M2701 Vdd nnT2BR nnT2BR GND dfet w=10 l=10
+ ad=0 pd=0 as=8649 ps=2854 
M2702 n_720 notRdy0 GND GND efet w=37 l=7
+ ad=0 pd=0 as=0 ps=0 
M2703 n_272 n_862 GND GND efet w=24 l=7
+ ad=0 pd=0 as=0 ps=0 
M2704 GND nnT2BR n_272 GND efet w=23 l=6
+ ad=0 pd=0 as=0 ps=0 
M2705 nnT2BR n_636 GND GND efet w=38 l=7
+ ad=1354 pd=392 as=0 ps=0 
M2706 n_720 n_720 Vdd GND dfet w=9 l=13
+ ad=1639 pd=572 as=0 ps=0 
M2707 n_680 cclk n_1688 GND efet w=12 l=9
+ ad=285 pd=112 as=0 ps=0 
M2708 op_EORS cclk n_982 GND efet w=11 l=7
+ ad=0 pd=0 as=148 ps=72 
M2709 op_ORS cclk n_88 GND efet w=12 l=7
+ ad=0 pd=0 as=164 ps=78 
M2710 Vdd n_1089 n_1089 GND dfet w=9 l=17
+ ad=0 pd=0 as=902 ps=258 
M2711 n_1089 n_1574 GND GND efet w=59 l=7
+ ad=731 pd=236 as=0 ps=0 
M2712 Vdd n_1141 n_1141 GND dfet w=9 l=15
+ ad=0 pd=0 as=434 ps=120 
M2713 alucin alucin Vdd GND dfet w=9 l=12
+ ad=1293 pd=422 as=0 ps=0 
M2714 Vdd n_1262 n_1262 GND dfet w=9 l=17
+ ad=0 pd=0 as=1925 ps=574 
M2715 n_1225 cclk pipedpc28 GND efet w=12 l=8
+ ad=0 pd=0 as=159 ps=70 
M2716 n_1407 n_1262 n_933 GND efet w=62 l=7
+ ad=470 pd=144 as=868 ps=238 
M2717 GND n_572 n_1407 GND efet w=65 l=7
+ ad=0 pd=0 as=0 ps=0 
M2718 Vdd n_10 n_10 GND dfet w=9 l=12
+ ad=0 pd=0 as=2446 ps=874 
M2719 n_1215 n_1215 Vdd GND dfet w=15 l=7
+ ad=2365 pd=860 as=0 ps=0 
M2720 GND x_op_jmp n_134 GND efet w=34 l=7
+ ad=0 pd=0 as=0 ps=0 
M2721 n_510 x_op_jmp GND GND efet w=37 l=6
+ ad=1639 pd=402 as=0 ps=0 
M2722 GND op_store nop_store GND efet w=49 l=7
+ ad=0 pd=0 as=754 ps=198 
M2723 n_1391 op_T4_brk GND GND efet w=39 l=7
+ ad=1223 pd=362 as=0 ps=0 
M2724 GND op_T2_php n_1391 GND efet w=38 l=7
+ ad=0 pd=0 as=0 ps=0 
M2725 n_368 op_T2_php_pha GND GND efet w=28 l=6
+ ad=2039 pd=478 as=0 ps=0 
M2726 GND op_T4_jmp n_368 GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M2727 n_368 op_T5_rti_rts GND GND efet w=28 l=6
+ ad=0 pd=0 as=0 ps=0 
M2728 GND xx_op_T5_jsr n_368 GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M2729 n_368 op_T2_jmp_abs GND GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M2730 GND x_op_T3_plp_pla n_368 GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M2731 n_790 op_lsr_ror_dec_inc GND GND efet w=27 l=7
+ ad=835 pd=208 as=0 ps=0 
M2732 GND op_asl_rol n_790 GND efet w=27 l=6
+ ad=0 pd=0 as=0 ps=0 
M2733 n_1065 op_T0_cli_sei GND GND efet w=27 l=6
+ ad=672 pd=178 as=0 ps=0 
M2734 n_134 n_134 Vdd GND dfet w=9 l=16
+ ad=4342 pd=1596 as=0 ps=0 
M2735 Vdd nop_store nop_store GND dfet w=10 l=12
+ ad=0 pd=0 as=1791 ps=588 
M2736 GND n_726 n_630 GND efet w=60 l=7
+ ad=0 pd=0 as=924 ps=260 
M2737 Vdd short_circuit_idx_add short_circuit_idx_add GND dfet w=9 l=11
+ ad=0 pd=0 as=1382 ps=424 
M2738 GND n_238 n_1215 GND efet w=174 l=6
+ ad=0 pd=0 as=0 ps=0 
M2739 GND pipeUNK36 short_circuit_idx_add GND efet w=102 l=7
+ ad=0 pd=0 as=1472 ps=388 
M2740 short_circuit_idx_add n_1137 GND GND efet w=40 l=7
+ ad=0 pd=0 as=0 ps=0 
M2741 n_1215 short_circuit_idx_add GND GND efet w=121 l=6
+ ad=0 pd=0 as=0 ps=0 
M2742 n_335 n_335 Vdd GND dfet w=9 l=7
+ ad=6382 pd=2174 as=0 ps=0 
M2743 n_630 n_630 Vdd GND dfet w=10 l=10
+ ad=4203 pd=1488 as=0 ps=0 
M2744 n_261 cclk pipeUNK36 GND efet w=12 l=8
+ ad=0 pd=0 as=346 ps=80 
M2745 short_circuit_idx_add n_916 GND GND efet w=39 l=6
+ ad=0 pd=0 as=0 ps=0 
M2746 n_10 op_branch_done GND GND efet w=53 l=5
+ ad=2102 pd=606 as=0 ps=0 
M2747 Vdd n_1211 n_1211 GND dfet w=8 l=11
+ ad=0 pd=0 as=5898 ps=2076 
M2748 GND op_T2_abs_access n_1211 GND efet w=44 l=5
+ ad=0 pd=0 as=2767 ps=782 
M2749 n_1211 nnT2BR GND GND efet w=19 l=8
+ ad=0 pd=0 as=0 ps=0 
M2750 GND n_1211 n_10 GND efet w=53 l=6
+ ad=0 pd=0 as=0 ps=0 
M2751 n_1211 nnT2BR GND GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M2752 GND n_862 n_1211 GND efet w=35 l=6
+ ad=0 pd=0 as=0 ps=0 
M2753 GND notRdy0 short_circuit_idx_add GND efet w=39 l=8
+ ad=0 pd=0 as=0 ps=0 
M2754 GND n_1716 n_180 GND efet w=36 l=6
+ ad=0 pd=0 as=834 ps=278 
M2755 n_720 cp1 n_1338 GND efet w=12 l=8
+ ad=0 pd=0 as=136 ps=72 
M2756 n_462 n_1338 GND GND efet w=77 l=6
+ ad=972 pd=314 as=0 ps=0 
M2757 Vdd n_462 n_462 GND dfet w=9 l=12
+ ad=0 pd=0 as=4437 ps=1502 
M2758 Vdd n_933 n_933 GND dfet w=9 l=12
+ ad=0 pd=0 as=1405 ps=430 
M2759 n_533 cp1 n_599 GND efet w=12 l=9
+ ad=0 pd=0 as=261 ps=74 
M2760 op_SUMS cclk n_415 GND efet w=11 l=8
+ ad=0 pd=0 as=276 ps=96 
M2761 op_SRS cclk n_968 GND efet w=12 l=8
+ ad=0 pd=0 as=188 ps=78 
M2762 Vdd notalucin notalucin GND dfet w=9 l=8
+ ad=0 pd=0 as=4636 ps=1634 
M2763 Vdd n_1375 n_1375 GND dfet w=10 l=16
+ ad=0 pd=0 as=955 ps=272 
M2764 GND n_982 n_1141 GND efet w=63 l=6
+ ad=0 pd=0 as=1092 ps=248 
M2765 n_1375 n_88 GND GND efet w=46 l=6
+ ad=657 pd=222 as=0 ps=0 
M2766 notalucin alucin GND GND efet w=63 l=7
+ ad=610 pd=196 as=0 ps=0 
M2767 Vdd n_1093 n_1093 GND dfet w=9 l=17
+ ad=0 pd=0 as=447 ps=106 
M2768 n_1526 n_1526 Vdd GND dfet w=9 l=13
+ ad=465 pd=150 as=0 ps=0 
M2769 GND n_968 n_1093 GND efet w=66 l=6
+ ad=0 pd=0 as=1123 ps=308 
M2770 n_931 n_415 GND GND efet w=53 l=7
+ ad=891 pd=318 as=0 ps=0 
M2771 Vdd n_931 n_931 GND dfet w=10 l=14
+ ad=0 pd=0 as=748 ps=252 
M2772 GND n_680 n_1526 GND efet w=63 l=6
+ ad=0 pd=0 as=962 ps=318 
M2773 n_1089 cp1 n_1529 GND efet w=11 l=8
+ ad=0 pd=0 as=285 ps=102 
M2774 n_1141 cp1 n_101 GND efet w=12 l=8
+ ad=0 pd=0 as=303 ps=82 
M2775 n_1375 cp1 n_95 GND efet w=12 l=8
+ ad=0 pd=0 as=321 ps=84 
M2776 n_779 cclk n_805 GND efet w=12 l=9
+ ad=0 pd=0 as=137 ps=68 
M2777 n_1594 cclk n_688 GND efet w=12 l=9
+ ad=0 pd=0 as=135 ps=68 
M2778 n_1649 cclk n_1027 GND efet w=12 l=9
+ ad=0 pd=0 as=132 ps=72 
M2779 n_795 cclk n_360 GND efet w=12 l=9
+ ad=0 pd=0 as=141 ps=72 
M2780 n_604 cclk n_1477 GND efet w=12 l=9
+ ad=0 pd=0 as=162 ps=72 
M2781 n_692 n_460 GND GND efet w=53 l=6
+ ad=843 pd=228 as=0 ps=0 
M2782 Vdd n_692 n_692 GND dfet w=9 l=13
+ ad=0 pd=0 as=1088 ps=338 
M2783 n_625 n_459 GND GND efet w=53 l=6
+ ad=878 pd=230 as=0 ps=0 
M2784 Vdd n_625 n_625 GND dfet w=9 l=13
+ ad=0 pd=0 as=1118 ps=340 
M2785 Vdd n_355 n_355 GND dfet w=9 l=10
+ ad=0 pd=0 as=1142 ps=388 
M2786 GND n_621 n_355 GND efet w=72 l=6
+ ad=0 pd=0 as=872 ps=206 
M2787 GND n_43 n_692 GND efet w=24 l=7
+ ad=0 pd=0 as=0 ps=0 
M2788 n_441 n_692 GND GND efet w=24 l=6
+ ad=366 pd=110 as=0 ps=0 
M2789 GND n_43 n_625 GND efet w=24 l=6
+ ad=0 pd=0 as=0 ps=0 
M2790 Vdd n_543 n_543 GND dfet w=9 l=10
+ ad=0 pd=0 as=1175 ps=384 
M2791 GND n_339 n_543 GND efet w=72 l=6
+ ad=0 pd=0 as=886 ps=210 
M2792 n_662 n_625 GND GND efet w=25 l=6
+ ad=368 pd=106 as=0 ps=0 
M2793 n_6 n_521 GND GND efet w=53 l=6
+ ad=881 pd=236 as=0 ps=0 
M2794 Vdd n_6 n_6 GND dfet w=10 l=13
+ ad=0 pd=0 as=1112 ps=342 
M2795 n_35 n_796 GND GND efet w=53 l=6
+ ad=878 pd=228 as=0 ps=0 
M2796 Vdd n_35 n_35 GND dfet w=10 l=13
+ ad=0 pd=0 as=1099 ps=340 
M2797 n_1534 n_805 GND GND efet w=53 l=6
+ ad=911 pd=230 as=0 ps=0 
M2798 Vdd n_1534 n_1534 GND dfet w=9 l=13
+ ad=0 pd=0 as=1128 ps=342 
M2799 n_1223 n_688 GND GND efet w=52 l=5
+ ad=899 pd=234 as=0 ps=0 
M2800 Vdd n_1223 n_1223 GND dfet w=10 l=13
+ ad=0 pd=0 as=1101 ps=340 
M2801 n_476 n_1027 GND GND efet w=53 l=6
+ ad=881 pd=230 as=0 ps=0 
M2802 Vdd n_476 n_476 GND dfet w=9 l=13
+ ad=0 pd=0 as=1131 ps=342 
M2803 GND n_43 n_6 GND efet w=26 l=6
+ ad=0 pd=0 as=0 ps=0 
M2804 n_593 n_355 GND GND efet w=25 l=6
+ ad=348 pd=108 as=0 ps=0 
M2805 n_441 n_441 Vdd GND dfet w=10 l=14
+ ad=1160 pd=362 as=0 ps=0 
M2806 Vdd n_692 dpc1_SBY GND dfet w=10 l=10
+ ad=0 pd=0 as=1780 ps=334 
M2807 n_662 n_662 Vdd GND dfet w=10 l=13
+ ad=1133 pd=354 as=0 ps=0 
M2808 n_196 n_543 GND GND efet w=25 l=6
+ ad=360 pd=104 as=0 ps=0 
M2809 Vdd n_625 dpc3_SBX GND dfet w=9 l=10
+ ad=0 pd=0 as=1744 ps=340 
M2810 n_593 n_593 Vdd GND dfet w=9 l=13
+ ad=1134 pd=364 as=0 ps=0 
M2811 n_282 n_6 GND GND efet w=25 l=6
+ ad=368 pd=108 as=0 ps=0 
M2812 GND n_43 n_35 GND efet w=25 l=7
+ ad=0 pd=0 as=0 ps=0 
M2813 Vdd n_355 dpc4_SSB GND dfet w=10 l=9
+ ad=0 pd=0 as=1361 ps=316 
M2814 n_196 n_196 Vdd GND dfet w=9 l=14
+ ad=1171 pd=362 as=0 ps=0 
M2815 dpc1_SBY n_1247 GND GND efet w=74 l=6
+ ad=0 pd=0 as=0 ps=0 
M2816 GND n_441 dpc1_SBY GND efet w=77 l=6
+ ad=0 pd=0 as=0 ps=0 
M2817 dpc3_SBX n_1247 GND GND efet w=76 l=7
+ ad=0 pd=0 as=0 ps=0 
M2818 GND n_662 dpc3_SBX GND efet w=77 l=6
+ ad=0 pd=0 as=0 ps=0 
M2819 GND n_593 dpc4_SSB GND efet w=98 l=6
+ ad=0 pd=0 as=0 ps=0 
M2820 Vdd n_543 dpc5_SADL GND dfet w=10 l=8
+ ad=0 pd=0 as=1328 ps=314 
M2821 n_71 n_35 GND GND efet w=25 l=6
+ ad=391 pd=112 as=0 ps=0 
M2822 GND n_43 n_1534 GND efet w=25 l=6
+ ad=0 pd=0 as=0 ps=0 
M2823 n_1230 n_360 GND GND efet w=53 l=6
+ ad=879 pd=232 as=0 ps=0 
M2824 Vdd n_1230 n_1230 GND dfet w=11 l=13
+ ad=0 pd=0 as=1100 ps=338 
M2825 n_1541 n_1477 GND GND efet w=53 l=6
+ ad=882 pd=232 as=0 ps=0 
M2826 Vdd n_1541 n_1541 GND dfet w=10 l=13
+ ad=0 pd=0 as=1090 ps=338 
M2827 n_91 n_1529 GND GND efet w=76 l=6
+ ad=749 pd=218 as=0 ps=0 
M2828 Vdd n_91 n_91 GND dfet w=10 l=11
+ ad=0 pd=0 as=1436 ps=472 
M2829 n_282 n_282 Vdd GND dfet w=9 l=13
+ ad=1132 pd=356 as=0 ps=0 
M2830 GND n_196 dpc5_SADL GND efet w=97 l=6
+ ad=0 pd=0 as=0 ps=0 
M2831 Vdd n_6 dpc6_SBS GND dfet w=10 l=9
+ ad=0 pd=0 as=1931 ps=376 
M2832 n_763 n_1534 GND GND efet w=24 l=6
+ ad=373 pd=110 as=0 ps=0 
M2833 GND n_43 n_1223 GND efet w=24 l=6
+ ad=0 pd=0 as=0 ps=0 
M2834 n_71 n_71 Vdd GND dfet w=10 l=13
+ ad=1137 pd=356 as=0 ps=0 
M2835 Vdd n_35 dpc7_SS GND dfet w=10 l=10
+ ad=0 pd=0 as=2147 ps=426 
M2836 n_225 n_1223 GND GND efet w=25 l=6
+ ad=386 pd=110 as=0 ps=0 
M2837 GND n_43 n_476 GND efet w=24 l=6
+ ad=0 pd=0 as=0 ps=0 
M2838 n_763 n_763 Vdd GND dfet w=10 l=13
+ ad=1129 pd=356 as=0 ps=0 
M2839 Vdd n_1534 dpc8_nDBADD GND dfet w=10 l=10
+ ad=0 pd=0 as=1841 ps=342 
M2840 dpc6_SBS n_1247 GND GND efet w=76 l=6
+ ad=0 pd=0 as=0 ps=0 
M2841 GND n_282 dpc6_SBS GND efet w=78 l=6
+ ad=0 pd=0 as=0 ps=0 
M2842 n_956 n_476 GND GND efet w=25 l=6
+ ad=425 pd=112 as=0 ps=0 
M2843 GND n_43 n_1230 GND efet w=24 l=7
+ ad=0 pd=0 as=0 ps=0 
M2844 n_225 n_225 Vdd GND dfet w=9 l=13
+ ad=1229 pd=354 as=0 ps=0 
M2845 Vdd n_1223 dpc9_DBADD GND dfet w=10 l=9
+ ad=0 pd=0 as=1818 ps=344 
M2846 dpc7_SS n_1247 GND GND efet w=76 l=6
+ ad=0 pd=0 as=0 ps=0 
M2847 GND n_71 dpc7_SS GND efet w=77 l=6
+ ad=0 pd=0 as=0 ps=0 
M2848 n_708 n_1230 GND GND efet w=25 l=6
+ ad=406 pd=110 as=0 ps=0 
M2849 GND n_43 n_1541 GND efet w=25 l=6
+ ad=0 pd=0 as=0 ps=0 
M2850 Vdd n_1364 n_1364 GND dfet w=9 l=11
+ ad=0 pd=0 as=1347 ps=448 
M2851 n_956 n_956 Vdd GND dfet w=10 l=13
+ ad=1127 pd=352 as=0 ps=0 
M2852 Vdd n_476 dpc12_0ADD GND dfet w=9 l=10
+ ad=0 pd=0 as=1943 ps=386 
M2853 dpc8_nDBADD n_1247 GND GND efet w=76 l=7
+ ad=0 pd=0 as=0 ps=0 
M2854 GND n_763 dpc8_nDBADD GND efet w=78 l=6
+ ad=0 pd=0 as=0 ps=0 
M2855 n_491 n_1541 GND GND efet w=25 l=6
+ ad=380 pd=108 as=0 ps=0 
M2856 GND n_91 n_1256 GND efet w=25 l=6
+ ad=0 pd=0 as=409 ps=132 
M2857 n_708 n_708 Vdd GND dfet w=9 l=13
+ ad=1133 pd=354 as=0 ps=0 
M2858 Vdd n_1230 dpc11_SBADD GND dfet w=10 l=10
+ ad=0 pd=0 as=2268 ps=424 
M2859 dpc9_DBADD n_1247 GND GND efet w=76 l=6
+ ad=0 pd=0 as=0 ps=0 
M2860 GND n_225 dpc9_DBADD GND efet w=77 l=6
+ ad=0 pd=0 as=0 ps=0 
M2861 n_491 n_491 Vdd GND dfet w=10 l=13
+ ad=1139 pd=356 as=0 ps=0 
M2862 Vdd n_1541 dpc10_ADLADD GND dfet w=9 l=10
+ ad=0 pd=0 as=1889 ps=322 
M2863 dpc12_0ADD n_1247 GND GND efet w=76 l=6
+ ad=0 pd=0 as=0 ps=0 
M2864 GND n_956 dpc12_0ADD GND efet w=77 l=6
+ ad=0 pd=0 as=0 ps=0 
M2865 dpc11_SBADD n_1247 GND GND efet w=76 l=7
+ ad=0 pd=0 as=0 ps=0 
M2866 GND n_708 dpc11_SBADD GND efet w=77 l=6
+ ad=0 pd=0 as=0 ps=0 
M2867 n_1256 n_1256 Vdd GND dfet w=10 l=14
+ ad=1525 pd=406 as=0 ps=0 
M2868 dpc10_ADLADD n_1247 GND GND efet w=74 l=6
+ ad=0 pd=0 as=0 ps=0 
M2869 GND n_491 dpc10_ADLADD GND efet w=76 l=6
+ ad=0 pd=0 as=0 ps=0 
M2870 dpc15_ANDS n_1256 GND GND efet w=126 l=7
+ ad=1088 pd=288 as=0 ps=0 
M2871 Vdd n_91 dpc15_ANDS GND dfet w=9 l=8
+ ad=0 pd=0 as=0 ps=0 
M2872 GND n_101 n_1364 GND efet w=75 l=6
+ ad=0 pd=0 as=737 ps=208 
M2873 n_531 n_95 GND GND efet w=75 l=6
+ ad=730 pd=206 as=0 ps=0 
M2874 Vdd n_531 n_531 GND dfet w=9 l=10
+ ad=0 pd=0 as=1439 ps=452 
M2875 GND n_1364 n_108 GND efet w=24 l=6
+ ad=0 pd=0 as=359 ps=108 
M2876 GND n_531 n_1255 GND efet w=24 l=6
+ ad=0 pd=0 as=362 ps=108 
M2877 n_108 n_108 Vdd GND dfet w=10 l=14
+ ad=1169 pd=384 as=0 ps=0 
M2878 Vdd n_1364 dpc16_EORS GND dfet w=9 l=9
+ ad=0 pd=0 as=965 ps=282 
M2879 n_1255 n_1255 Vdd GND dfet w=9 l=14
+ ad=1358 pd=382 as=0 ps=0 
M2880 adl0 n_0_ADL0 GND GND efet w=15 l=7
+ ad=2953 pd=756 as=0 ps=0 
M2881 nABL0 cclk n_1100 GND efet w=12 l=8
+ ad=288 pd=90 as=0 ps=0 
M2882 n_246 ADL_ABL nABL0 GND efet w=12 l=6
+ ad=96 pd=40 as=0 ps=0 
M2883 n_123 cp1 n_246 GND efet w=12 l=7
+ ad=909 pd=256 as=0 ps=0 
M2884 abl0 nABL0 GND GND efet w=94 l=7
+ ad=839 pd=248 as=0 ps=0 
M2885 abl0 abl0 Vdd GND dfet w=9 l=14
+ ad=2842 pd=836 as=0 ps=0 
M2886 ab0 n_855 Vdd GND efet w=110 l=7
+ ad=0 pd=0 as=0 ps=0 
M2887 GND n_66 ab1 GND efet w=126 l=6
+ ad=0 pd=0 as=16284 ps=2466 
M2888 ab1 n_66 GND GND efet w=302 l=7
+ ad=0 pd=0 as=0 ps=0 
M2889 ab1 n_66 GND GND efet w=355 l=6
+ ad=0 pd=0 as=0 ps=0 
M2890 ab1 n_66 GND GND efet w=171 l=7
+ ad=0 pd=0 as=0 ps=0 
M2891 GND n_842 n_1479 GND efet w=127 l=7
+ ad=0 pd=0 as=1560 ps=374 
M2892 Vdd n_1479 ab1 GND efet w=68 l=6
+ ad=0 pd=0 as=0 ps=0 
M2893 Vdd n_1479 ab1 GND efet w=240 l=7
+ ad=0 pd=0 as=0 ps=0 
M2894 n_842 abl1 GND GND efet w=36 l=7
+ ad=453 pd=134 as=0 ps=0 
M2895 Vdd n_1479 ab1 GND efet w=240 l=7
+ ad=0 pd=0 as=0 ps=0 
M2896 n_842 n_842 Vdd GND dfet w=10 l=11
+ ad=1708 pd=542 as=0 ps=0 
M2897 GND abl1 n_66 GND efet w=154 l=7
+ ad=0 pd=0 as=1492 ps=404 
M2898 n_1479 abl1 Vdd GND dfet w=17 l=6
+ ad=0 pd=0 as=0 ps=0 
M2899 Vdd n_1479 ab1 GND efet w=239 l=6
+ ad=0 pd=0 as=0 ps=0 
M2900 n_66 n_842 Vdd GND dfet w=20 l=7
+ ad=0 pd=0 as=0 ps=0 
M2901 GND adl0 n_123 GND efet w=83 l=7
+ ad=0 pd=0 as=0 ps=0 
M2902 n_123 n_123 Vdd GND dfet w=10 l=12
+ ad=309 pd=82 as=0 ps=0 
M2903 GND n_0_ADL1 adl1 GND efet w=16 l=8
+ ad=0 pd=0 as=2847 ps=720 
M2904 nABL1 cclk n_66 GND efet w=11 l=7
+ ad=272 pd=90 as=0 ps=0 
M2905 n_416 ADL_ABL nABL1 GND efet w=11 l=6
+ ad=88 pd=38 as=0 ps=0 
M2906 n_1016 cp1 n_416 GND efet w=11 l=9
+ ad=924 pd=262 as=0 ps=0 
M2907 abl1 nABL1 GND GND efet w=96 l=6
+ ad=938 pd=254 as=0 ps=0 
M2908 abl1 abl1 Vdd GND dfet w=10 l=13
+ ad=2819 pd=840 as=0 ps=0 
M2909 ab1 n_1479 Vdd GND efet w=111 l=7
+ ad=0 pd=0 as=0 ps=0 
M2910 GND n_642 ab2 GND efet w=127 l=7
+ ad=0 pd=0 as=16693 ps=2482 
M2911 GND n_951 n_1152 GND efet w=126 l=7
+ ad=0 pd=0 as=1698 ps=378 
M2912 ab2 n_642 GND GND efet w=302 l=6
+ ad=0 pd=0 as=0 ps=0 
M2913 ab2 n_642 GND GND efet w=355 l=7
+ ad=0 pd=0 as=0 ps=0 
M2914 ab2 n_642 GND GND efet w=171 l=7
+ ad=0 pd=0 as=0 ps=0 
M2915 n_951 abl2 GND GND efet w=36 l=7
+ ad=427 pd=134 as=0 ps=0 
M2916 Vdd n_1152 ab2 GND efet w=68 l=6
+ ad=0 pd=0 as=0 ps=0 
M2917 Vdd n_1152 ab2 GND efet w=240 l=6
+ ad=0 pd=0 as=0 ps=0 
M2918 n_951 n_951 Vdd GND dfet w=10 l=11
+ ad=1839 pd=540 as=0 ps=0 
M2919 GND abl2 n_642 GND efet w=155 l=7
+ ad=0 pd=0 as=1576 ps=418 
M2920 n_1152 abl2 Vdd GND dfet w=17 l=6
+ ad=0 pd=0 as=0 ps=0 
M2921 n_642 n_951 Vdd GND dfet w=21 l=7
+ ad=0 pd=0 as=0 ps=0 
M2922 GND adl1 n_1016 GND efet w=82 l=7
+ ad=0 pd=0 as=0 ps=0 
M2923 n_1016 n_1016 Vdd GND dfet w=10 l=10
+ ad=249 pd=74 as=0 ps=0 
M2924 Vdd n_564 n_564 GND dfet w=10 l=17
+ ad=0 pd=0 as=377 ps=104 
M2925 GND noty0 n_564 GND efet w=55 l=6
+ ad=0 pd=0 as=1479 ps=318 
M2926 Vdd noty0 noty0 GND dfet w=10 l=21
+ ad=0 pd=0 as=858 ps=248 
M2927 noty0 y0 GND GND efet w=36 l=7
+ ad=547 pd=166 as=0 ps=0 
M2928 y0 cclk n_564 GND efet w=12 l=9
+ ad=250 pd=86 as=0 ps=0 
M2929 n_564 dpc0_YSB sb0 GND efet w=14 l=7
+ ad=0 pd=0 as=4619 ps=1126 
M2930 y0 dpc1_SBY sb0 GND efet w=12 l=7
+ ad=0 pd=0 as=0 ps=0 
M2931 GND n_0_ADL2 adl2 GND efet w=16 l=7
+ ad=0 pd=0 as=2803 ps=710 
M2932 Vdd n_767 n_767 GND dfet w=10 l=17
+ ad=0 pd=0 as=309 ps=82 
M2933 GND noty1 n_767 GND efet w=55 l=7
+ ad=0 pd=0 as=1546 ps=354 
M2934 Vdd noty1 noty1 GND dfet w=10 l=21
+ ad=0 pd=0 as=967 ps=256 
M2935 noty1 y1 GND GND efet w=35 l=6
+ ad=569 pd=170 as=0 ps=0 
M2936 y1 cclk n_767 GND efet w=12 l=8
+ ad=278 pd=98 as=0 ps=0 
M2937 n_767 dpc0_YSB sb1 GND efet w=14 l=7
+ ad=0 pd=0 as=4095 ps=982 
M2938 nABL2 cclk n_642 GND efet w=12 l=8
+ ad=300 pd=92 as=0 ps=0 
M2939 n_1636 ADL_ABL nABL2 GND efet w=12 l=6
+ ad=96 pd=40 as=0 ps=0 
M2940 n_935 cp1 n_1636 GND efet w=12 l=8
+ ad=864 pd=262 as=0 ps=0 
M2941 abl2 nABL2 GND GND efet w=94 l=6
+ ad=890 pd=252 as=0 ps=0 
M2942 abl2 abl2 Vdd GND dfet w=9 l=13
+ ad=2840 pd=840 as=0 ps=0 
M2943 Vdd n_1152 ab2 GND efet w=241 l=6
+ ad=0 pd=0 as=0 ps=0 
M2944 Vdd n_1152 ab2 GND efet w=241 l=6
+ ad=0 pd=0 as=0 ps=0 
M2945 ab2 n_1152 Vdd GND efet w=112 l=7
+ ad=0 pd=0 as=0 ps=0 
M2946 GND n_990 n_1041 GND efet w=126 l=7
+ ad=0 pd=0 as=1920 ps=438 
M2947 n_990 abl3 GND GND efet w=35 l=8
+ ad=410 pd=132 as=0 ps=0 
M2948 GND n_138 ab3 GND efet w=127 l=7
+ ad=0 pd=0 as=16511 ps=2472 
M2949 n_990 n_990 Vdd GND dfet w=10 l=10
+ ad=1851 pd=540 as=0 ps=0 
M2950 GND abl3 n_138 GND efet w=155 l=7
+ ad=0 pd=0 as=1599 ps=418 
M2951 n_1041 abl3 Vdd GND dfet w=18 l=6
+ ad=0 pd=0 as=0 ps=0 
M2952 ab3 n_138 GND GND efet w=302 l=7
+ ad=0 pd=0 as=0 ps=0 
M2953 ab3 n_138 GND GND efet w=355 l=7
+ ad=0 pd=0 as=0 ps=0 
M2954 ab3 n_138 GND GND efet w=171 l=7
+ ad=0 pd=0 as=0 ps=0 
M2955 n_138 n_990 Vdd GND dfet w=22 l=8
+ ad=0 pd=0 as=0 ps=0 
M2956 GND adl2 n_935 GND efet w=83 l=6
+ ad=0 pd=0 as=0 ps=0 
M2957 y1 dpc1_SBY sb1 GND efet w=11 l=8
+ ad=0 pd=0 as=0 ps=0 
M2958 Vdd n_1491 n_1491 GND dfet w=10 l=17
+ ad=0 pd=0 as=309 ps=82 
M2959 Vdd n_1169 n_1169 GND dfet w=10 l=16
+ ad=0 pd=0 as=294 ps=80 
M2960 GND notx0 n_1169 GND efet w=55 l=7
+ ad=0 pd=0 as=1511 ps=352 
M2961 Vdd notx0 notx0 GND dfet w=9 l=21
+ ad=0 pd=0 as=969 ps=256 
M2962 notx0 x0 GND GND efet w=35 l=6
+ ad=481 pd=164 as=0 ps=0 
M2963 x0 cclk n_1169 GND efet w=12 l=8
+ ad=266 pd=92 as=0 ps=0 
M2964 n_1169 dpc2_XSB sb0 GND efet w=13 l=8
+ ad=0 pd=0 as=0 ps=0 
M2965 Vdd n_332 n_332 GND dfet w=10 l=17
+ ad=0 pd=0 as=370 ps=102 
M2966 n_332 dpc5_SADL adl0 GND efet w=16 l=7
+ ad=1966 pd=458 as=0 ps=0 
M2967 Vdd n_983 n_983 GND dfet w=9 l=20
+ ad=0 pd=0 as=488 ps=132 
M2968 x0 dpc3_SBX sb0 GND efet w=11 l=8
+ ad=0 pd=0 as=0 ps=0 
M2969 Vdd n_1709 n_1709 GND dfet w=10 l=16
+ ad=0 pd=0 as=294 ps=80 
M2970 GND notx1 n_1709 GND efet w=55 l=6
+ ad=0 pd=0 as=1463 ps=354 
M2971 Vdd notx1 notx1 GND dfet w=10 l=21
+ ad=0 pd=0 as=953 ps=258 
M2972 notx1 x1 GND GND efet w=35 l=7
+ ad=532 pd=168 as=0 ps=0 
M2973 x1 cclk n_1709 GND efet w=11 l=7
+ ad=251 pd=94 as=0 ps=0 
M2974 n_332 dpc4_SSB sb0 GND efet w=17 l=8
+ ad=0 pd=0 as=0 ps=0 
M2975 GND nots0 n_332 GND efet w=45 l=7
+ ad=0 pd=0 as=0 ps=0 
M2976 n_983 s0 GND GND efet w=32 l=7
+ ad=849 pd=230 as=0 ps=0 
M2977 n_983 cclk nots0 GND efet w=12 l=7
+ ad=0 pd=0 as=324 ps=104 
M2978 n_332 dpc7_SS s0 GND efet w=12 l=8
+ ad=0 pd=0 as=333 ps=76 
M2979 s0 dpc6_SBS sb0 GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M2980 sb0 cclk Vdd GND efet w=24 l=7
+ ad=0 pd=0 as=0 ps=0 
M2981 Vdd n_694 n_694 GND dfet w=10 l=17
+ ad=0 pd=0 as=378 ps=102 
M2982 n_694 dpc5_SADL adl1 GND efet w=15 l=8
+ ad=1897 pd=454 as=0 ps=0 
M2983 Vdd n_1711 n_1711 GND dfet w=9 l=20
+ ad=0 pd=0 as=488 ps=132 
M2984 n_1709 dpc2_XSB sb1 GND efet w=13 l=8
+ ad=0 pd=0 as=0 ps=0 
M2985 x1 dpc3_SBX sb1 GND efet w=11 l=8
+ ad=0 pd=0 as=0 ps=0 
M2986 GND noty2 n_1491 GND efet w=56 l=6
+ ad=0 pd=0 as=1549 ps=356 
M2987 Vdd noty2 noty2 GND dfet w=9 l=21
+ ad=0 pd=0 as=964 ps=258 
M2988 noty2 y2 GND GND efet w=37 l=7
+ ad=529 pd=164 as=0 ps=0 
M2989 y2 cclk n_1491 GND efet w=12 l=8
+ ad=281 pd=96 as=0 ps=0 
M2990 n_935 n_935 Vdd GND dfet w=9 l=11
+ ad=250 pd=74 as=0 ps=0 
M2991 n_1491 dpc0_YSB sb2 GND efet w=13 l=7
+ ad=0 pd=0 as=3995 ps=980 
M2992 nABL3 cclk n_138 GND efet w=12 l=8
+ ad=282 pd=92 as=0 ps=0 
M2993 n_864 ADL_ABL nABL3 GND efet w=12 l=7
+ ad=84 pd=38 as=0 ps=0 
M2994 n_1507 cp1 n_864 GND efet w=12 l=8
+ ad=1104 pd=288 as=0 ps=0 
M2995 abl3 nABL3 GND GND efet w=94 l=7
+ ad=879 pd=250 as=0 ps=0 
M2996 abl3 abl3 Vdd GND dfet w=10 l=14
+ ad=2730 pd=824 as=0 ps=0 
M2997 Vdd n_1041 ab3 GND efet w=69 l=6
+ ad=0 pd=0 as=0 ps=0 
M2998 GND adl3 n_1507 GND efet w=87 l=7
+ ad=0 pd=0 as=0 ps=0 
M2999 n_1507 n_1507 Vdd GND dfet w=9 l=10
+ ad=220 pd=70 as=0 ps=0 
M3000 y2 dpc1_SBY sb2 GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M3001 Vdd n_1531 n_1531 GND dfet w=10 l=16
+ ad=0 pd=0 as=304 ps=80 
M3002 GND noty3 n_1531 GND efet w=56 l=6
+ ad=0 pd=0 as=1486 ps=358 
M3003 Vdd noty3 noty3 GND dfet w=9 l=21
+ ad=0 pd=0 as=964 ps=258 
M3004 noty3 y3 GND GND efet w=37 l=6
+ ad=512 pd=164 as=0 ps=0 
M3005 y3 cclk n_1531 GND efet w=11 l=9
+ ad=265 pd=96 as=0 ps=0 
M3006 n_1531 dpc0_YSB sb3 GND efet w=13 l=8
+ ad=0 pd=0 as=4031 ps=980 
M3007 Vdd n_1041 ab3 GND efet w=241 l=7
+ ad=0 pd=0 as=0 ps=0 
M3008 Vdd n_1041 ab3 GND efet w=241 l=7
+ ad=0 pd=0 as=0 ps=0 
M3009 Vdd n_1041 ab3 GND efet w=240 l=6
+ ad=0 pd=0 as=0 ps=0 
M3010 ab3 n_1041 Vdd GND efet w=111 l=7
+ ad=0 pd=0 as=0 ps=0 
M3011 GND n_1676 n_634 GND efet w=126 l=7
+ ad=0 pd=0 as=1583 ps=376 
M3012 n_1676 abl4 GND GND efet w=36 l=7
+ ad=481 pd=134 as=0 ps=0 
M3013 n_1676 n_1676 Vdd GND dfet w=10 l=10
+ ad=1792 pd=542 as=0 ps=0 
M3014 GND abl4 n_86 GND efet w=155 l=7
+ ad=0 pd=0 as=1595 ps=422 
M3015 n_634 abl4 Vdd GND dfet w=18 l=6
+ ad=0 pd=0 as=0 ps=0 
M3016 n_86 n_1676 Vdd GND dfet w=22 l=7
+ ad=0 pd=0 as=0 ps=0 
M3017 y3 dpc1_SBY sb3 GND efet w=11 l=8
+ ad=0 pd=0 as=0 ps=0 
M3018 nABL4 cclk n_86 GND efet w=12 l=8
+ ad=282 pd=92 as=0 ps=0 
M3019 n_738 ADL_ABL nABL4 GND efet w=12 l=7
+ ad=84 pd=38 as=0 ps=0 
M3020 n_1519 cp1 n_738 GND efet w=12 l=8
+ ad=903 pd=266 as=0 ps=0 
M3021 abl4 nABL4 GND GND efet w=95 l=6
+ ad=889 pd=254 as=0 ps=0 
M3022 abl4 abl4 Vdd GND dfet w=9 l=14
+ ad=2720 pd=836 as=0 ps=0 
M3023 GND n_86 ab4 GND efet w=126 l=7
+ ad=0 pd=0 as=16302 ps=2466 
M3024 ab4 n_86 GND GND efet w=301 l=7
+ ad=0 pd=0 as=0 ps=0 
M3025 ab4 n_86 GND GND efet w=356 l=7
+ ad=0 pd=0 as=0 ps=0 
M3026 ab4 n_86 GND GND efet w=172 l=7
+ ad=0 pd=0 as=0 ps=0 
M3027 Vdd n_634 ab4 GND efet w=68 l=6
+ ad=0 pd=0 as=0 ps=0 
M3028 Vdd n_634 ab4 GND efet w=238 l=7
+ ad=0 pd=0 as=0 ps=0 
M3029 Vdd n_634 ab4 GND efet w=239 l=6
+ ad=0 pd=0 as=0 ps=0 
M3030 Vdd n_634 ab4 GND efet w=239 l=6
+ ad=0 pd=0 as=0 ps=0 
M3031 ab4 n_634 Vdd GND efet w=111 l=7
+ ad=0 pd=0 as=0 ps=0 
M3032 GND n_172 n_1633 GND efet w=126 l=7
+ ad=0 pd=0 as=1594 ps=376 
M3033 n_172 abl5 GND GND efet w=36 l=8
+ ad=410 pd=134 as=0 ps=0 
M3034 GND n_210 ab5 GND efet w=126 l=7
+ ad=0 pd=0 as=16631 ps=2472 
M3035 ab5 n_210 GND GND efet w=302 l=7
+ ad=0 pd=0 as=0 ps=0 
M3036 ab5 n_210 GND GND efet w=358 l=7
+ ad=0 pd=0 as=0 ps=0 
M3037 ab5 n_210 GND GND efet w=171 l=6
+ ad=0 pd=0 as=0 ps=0 
M3038 n_172 n_172 Vdd GND dfet w=11 l=10
+ ad=1719 pd=540 as=0 ps=0 
M3039 GND abl5 n_210 GND efet w=154 l=7
+ ad=0 pd=0 as=1607 ps=400 
M3040 n_1633 abl5 Vdd GND dfet w=19 l=6
+ ad=0 pd=0 as=0 ps=0 
M3041 n_210 n_172 Vdd GND dfet w=21 l=7
+ ad=0 pd=0 as=0 ps=0 
M3042 GND adl4 n_1519 GND efet w=83 l=6
+ ad=0 pd=0 as=0 ps=0 
M3043 Vdd n_658 n_658 GND dfet w=10 l=16
+ ad=0 pd=0 as=304 ps=80 
M3044 GND noty4 n_658 GND efet w=56 l=7
+ ad=0 pd=0 as=1430 ps=348 
M3045 Vdd noty4 noty4 GND dfet w=10 l=21
+ ad=0 pd=0 as=975 ps=258 
M3046 noty4 y4 GND GND efet w=35 l=7
+ ad=522 pd=166 as=0 ps=0 
M3047 y4 cclk n_658 GND efet w=11 l=8
+ ad=262 pd=90 as=0 ps=0 
M3048 n_1519 n_1519 Vdd GND dfet w=9 l=10
+ ad=224 pd=72 as=0 ps=0 
M3049 n_658 dpc0_YSB sb4 GND efet w=13 l=8
+ ad=0 pd=0 as=4148 ps=1052 
M3050 y4 dpc1_SBY sb4 GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M3051 nABL5 cclk n_210 GND efet w=11 l=7
+ ad=272 pd=90 as=0 ps=0 
M3052 n_463 ADL_ABL nABL5 GND efet w=11 l=7
+ ad=77 pd=36 as=0 ps=0 
M3053 n_1094 cp1 n_463 GND efet w=11 l=8
+ ad=933 pd=268 as=0 ps=0 
M3054 abl5 nABL5 GND GND efet w=97 l=6
+ ad=942 pd=254 as=0 ps=0 
M3055 abl5 abl5 Vdd GND dfet w=10 l=14
+ ad=2812 pd=836 as=0 ps=0 
M3056 Vdd n_1633 ab5 GND efet w=69 l=6
+ ad=0 pd=0 as=0 ps=0 
M3057 Vdd n_1633 ab5 GND efet w=241 l=7
+ ad=0 pd=0 as=0 ps=0 
M3058 Vdd n_1633 ab5 GND efet w=240 l=7
+ ad=0 pd=0 as=0 ps=0 
M3059 Vdd n_1633 ab5 GND efet w=239 l=6
+ ad=0 pd=0 as=0 ps=0 
M3060 ab5 n_1633 Vdd GND efet w=111 l=7
+ ad=0 pd=0 as=0 ps=0 
M3061 GND n_1195 n_1191 GND efet w=127 l=7
+ ad=0 pd=0 as=1584 ps=374 
M3062 n_1195 abl6 GND GND efet w=36 l=7
+ ad=428 pd=134 as=0 ps=0 
M3063 n_1195 n_1195 Vdd GND dfet w=10 l=11
+ ad=1708 pd=542 as=0 ps=0 
M3064 GND abl6 n_1254 GND efet w=156 l=7
+ ad=0 pd=0 as=1510 ps=408 
M3065 n_1191 abl6 Vdd GND dfet w=19 l=7
+ ad=0 pd=0 as=0 ps=0 
M3066 n_1254 n_1195 Vdd GND dfet w=20 l=7
+ ad=0 pd=0 as=0 ps=0 
M3067 GND adl5 n_1094 GND efet w=84 l=7
+ ad=0 pd=0 as=0 ps=0 
M3068 Vdd n_733 n_733 GND dfet w=9 l=17
+ ad=0 pd=0 as=320 ps=82 
M3069 GND noty5 n_733 GND efet w=57 l=7
+ ad=0 pd=0 as=1467 ps=352 
M3070 Vdd noty5 noty5 GND dfet w=9 l=20
+ ad=0 pd=0 as=957 ps=256 
M3071 noty5 y5 GND GND efet w=35 l=7
+ ad=491 pd=162 as=0 ps=0 
M3072 y5 cclk n_733 GND efet w=11 l=8
+ ad=264 pd=90 as=0 ps=0 
M3073 n_1094 n_1094 Vdd GND dfet w=9 l=11
+ ad=267 pd=76 as=0 ps=0 
M3074 n_733 dpc0_YSB sb5 GND efet w=13 l=8
+ ad=0 pd=0 as=4004 ps=980 
M3075 y5 dpc1_SBY sb5 GND efet w=11 l=7
+ ad=0 pd=0 as=0 ps=0 
M3076 nABL6 cclk n_1254 GND efet w=12 l=7
+ ad=294 pd=94 as=0 ps=0 
M3077 n_524 ADL_ABL nABL6 GND efet w=12 l=7
+ ad=84 pd=38 as=0 ps=0 
M3078 n_1548 cp1 n_524 GND efet w=12 l=8
+ ad=953 pd=264 as=0 ps=0 
M3079 abl6 nABL6 GND GND efet w=97 l=6
+ ad=915 pd=250 as=0 ps=0 
M3080 abl6 abl6 Vdd GND dfet w=10 l=14
+ ad=2853 pd=838 as=0 ps=0 
M3081 GND n_1254 ab6 GND efet w=139 l=7
+ ad=0 pd=0 as=16917 ps=2466 
M3082 ab6 n_1254 GND GND efet w=325 l=7
+ ad=0 pd=0 as=0 ps=0 
M3083 ab6 n_1254 GND GND efet w=359 l=7
+ ad=0 pd=0 as=0 ps=0 
M3084 GND n_1026 n_322 GND efet w=125 l=6
+ ad=0 pd=0 as=1761 ps=390 
M3085 n_1026 abl7 GND GND efet w=36 l=7
+ ad=435 pd=134 as=0 ps=0 
M3086 Vdd n_1191 ab6 GND efet w=124 l=7
+ ad=0 pd=0 as=0 ps=0 
M3087 ab6 n_1254 GND GND efet w=210 l=6
+ ad=0 pd=0 as=0 ps=0 
M3088 Vdd n_1191 ab6 GND efet w=239 l=7
+ ad=0 pd=0 as=0 ps=0 
M3089 Vdd n_1191 ab6 GND efet w=239 l=6
+ ad=0 pd=0 as=0 ps=0 
M3090 Vdd n_1191 ab6 GND efet w=250 l=7
+ ad=0 pd=0 as=0 ps=0 
M3091 n_1026 n_1026 Vdd GND dfet w=11 l=10
+ ad=1692 pd=536 as=0 ps=0 
M3092 GND abl7 n_171 GND efet w=155 l=7
+ ad=0 pd=0 as=1569 ps=414 
M3093 n_322 abl7 Vdd GND dfet w=18 l=7
+ ad=0 pd=0 as=0 ps=0 
M3094 n_171 n_1026 Vdd GND dfet w=20 l=7
+ ad=0 pd=0 as=0 ps=0 
M3095 GND adl6 n_1548 GND efet w=83 l=6
+ ad=0 pd=0 as=0 ps=0 
M3096 Vdd n_518 n_518 GND dfet w=10 l=16
+ ad=0 pd=0 as=304 ps=80 
M3097 Vdd n_1694 n_1694 GND dfet w=10 l=17
+ ad=0 pd=0 as=309 ps=82 
M3098 GND notx2 n_1694 GND efet w=56 l=6
+ ad=0 pd=0 as=1485 ps=356 
M3099 Vdd notx2 notx2 GND dfet w=10 l=21
+ ad=0 pd=0 as=947 ps=256 
M3100 n_694 dpc4_SSB sb1 GND efet w=17 l=7
+ ad=0 pd=0 as=0 ps=0 
M3101 notx2 x2 GND GND efet w=36 l=7
+ ad=537 pd=166 as=0 ps=0 
M3102 x2 cclk n_1694 GND efet w=12 l=9
+ ad=266 pd=96 as=0 ps=0 
M3103 GND nots1 n_694 GND efet w=43 l=6
+ ad=0 pd=0 as=0 ps=0 
M3104 n_1711 s1 GND GND efet w=32 l=7
+ ad=875 pd=232 as=0 ps=0 
M3105 n_1711 cclk nots1 GND efet w=12 l=8
+ ad=0 pd=0 as=279 ps=100 
M3106 n_694 dpc7_SS s1 GND efet w=12 l=9
+ ad=0 pd=0 as=342 ps=76 
M3107 s1 dpc6_SBS sb1 GND efet w=13 l=8
+ ad=0 pd=0 as=0 ps=0 
M3108 sb1 cclk Vdd GND efet w=24 l=7
+ ad=0 pd=0 as=0 ps=0 
M3109 Vdd n_1389 n_1389 GND dfet w=10 l=17
+ ad=0 pd=0 as=372 ps=102 
M3110 n_1389 dpc5_SADL adl2 GND efet w=16 l=5
+ ad=1915 pd=462 as=0 ps=0 
M3111 Vdd n_1190 n_1190 GND dfet w=9 l=20
+ ad=0 pd=0 as=482 ps=130 
M3112 n_1694 dpc2_XSB sb2 GND efet w=13 l=8
+ ad=0 pd=0 as=0 ps=0 
M3113 x2 dpc3_SBX sb2 GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M3114 Vdd n_242 n_242 GND dfet w=10 l=16
+ ad=0 pd=0 as=294 ps=80 
M3115 GND notx3 n_242 GND efet w=55 l=6
+ ad=0 pd=0 as=1587 ps=354 
M3116 Vdd notx3 notx3 GND dfet w=9 l=21
+ ad=0 pd=0 as=947 ps=256 
M3117 notx3 x3 GND GND efet w=36 l=6
+ ad=557 pd=168 as=0 ps=0 
M3118 x3 cclk n_242 GND efet w=12 l=8
+ ad=289 pd=96 as=0 ps=0 
M3119 n_242 dpc2_XSB sb3 GND efet w=13 l=8
+ ad=0 pd=0 as=0 ps=0 
M3120 n_1389 dpc4_SSB sb2 GND efet w=17 l=8
+ ad=0 pd=0 as=0 ps=0 
M3121 GND nots2 n_1389 GND efet w=44 l=7
+ ad=0 pd=0 as=0 ps=0 
M3122 n_1190 s2 GND GND efet w=33 l=7
+ ad=874 pd=230 as=0 ps=0 
M3123 n_1190 cclk nots2 GND efet w=12 l=8
+ ad=0 pd=0 as=272 ps=100 
M3124 GND n_108 dpc16_EORS GND efet w=111 l=5
+ ad=0 pd=0 as=0 ps=0 
M3125 dpc13_ORS n_1255 GND GND efet w=111 l=7
+ ad=955 pd=260 as=0 ps=0 
M3126 Vdd n_531 dpc13_ORS GND dfet w=9 l=9
+ ad=0 pd=0 as=0 ps=0 
M3127 GND pipedpc28 dpc28_0ADH0 GND efet w=94 l=6
+ ad=0 pd=0 as=1028 ps=276 
M3128 n_877 n_506 GND GND efet w=56 l=6
+ ad=1112 pd=332 as=0 ps=0 
M3129 Vdd dpc28_0ADH0 dpc28_0ADH0 GND dfet w=9 l=16
+ ad=0 pd=0 as=4160 ps=1520 
M3130 n_674 n_674 Vdd GND dfet w=9 l=11
+ ad=671 pd=240 as=0 ps=0 
M3131 Vdd dpc22_nDSA dpc22_nDSA GND dfet w=9 l=12
+ ad=0 pd=0 as=6783 ps=2702 
M3132 n_674 n_25 GND GND efet w=50 l=6
+ ad=936 pd=322 as=0 ps=0 
M3133 n_80 n_267 GND GND efet w=38 l=7
+ ad=927 pd=250 as=0 ps=0 
M3134 GND n_1130 n_80 GND efet w=46 l=5
+ ad=0 pd=0 as=0 ps=0 
M3135 GND n_599 dpc22_nDSA GND efet w=79 l=6
+ ad=0 pd=0 as=668 ps=210 
M3136 Vdd n_80 n_80 GND dfet w=8 l=10
+ ad=0 pd=0 as=230 ps=72 
M3137 n_1245 n_1245 Vdd GND dfet w=10 l=8
+ ad=3156 pd=1042 as=0 ps=0 
M3138 n_1245 aluvout GND GND efet w=74 l=6
+ ad=909 pd=250 as=0 ps=0 
M3139 GND n_933 n_877 GND efet w=49 l=7
+ ad=0 pd=0 as=0 ps=0 
M3140 n_1211 n_1002 GND GND efet w=36 l=6
+ ad=0 pd=0 as=0 ps=0 
M3141 n_182 n_182 Vdd GND dfet w=10 l=12
+ ad=3753 pd=1308 as=0 ps=0 
M3142 GND op_T5_rts n_182 GND efet w=29 l=6
+ ad=0 pd=0 as=2882 ps=798 
M3143 n_1151 n_1262 GND GND efet w=68 l=6
+ ad=414 pd=150 as=0 ps=0 
M3144 GND n_467 n_10 GND efet w=28 l=6
+ ad=0 pd=0 as=0 ps=0 
M3145 n_182 n_236 n_1151 GND efet w=68 l=6
+ ad=0 pd=0 as=0 ps=0 
M3146 GND n_1286 n_1211 GND efet w=45 l=7
+ ad=0 pd=0 as=0 ps=0 
M3147 Vdd n_467 n_467 GND dfet w=9 l=14
+ ad=0 pd=0 as=1216 ps=386 
M3148 GND nnT2BR n_1427 GND efet w=46 l=7
+ ad=0 pd=0 as=1281 ps=400 
M3149 n_1427 n_1427 Vdd GND dfet w=9 l=17
+ ad=1924 pd=652 as=0 ps=0 
M3150 n_930 n_930 Vdd GND dfet w=9 l=17
+ ad=1403 pd=434 as=0 ps=0 
M3151 n_930 n_134 GND GND efet w=34 l=6
+ ad=1190 pd=360 as=0 ps=0 
M3152 n_1705 n_467 GND GND efet w=32 l=6
+ ad=1337 pd=378 as=0 ps=0 
M3153 n_877 n_877 Vdd GND dfet w=9 l=10
+ ad=950 pd=310 as=0 ps=0 
M3154 n_1093 cp1 n_226 GND efet w=12 l=8
+ ad=0 pd=0 as=280 ps=80 
M3155 n_931 cp1 n_1674 GND efet w=12 l=8
+ ad=0 pd=0 as=294 ps=82 
M3156 n_1526 cp1 n_1450 GND efet w=12 l=8
+ ad=0 pd=0 as=316 ps=112 
M3157 n_80 cclk n_1333 GND efet w=12 l=9
+ ad=0 pd=0 as=189 ps=78 
M3158 n_1130 cclk n_512 GND efet w=12 l=9
+ ad=0 pd=0 as=213 ps=82 
M3159 n_674 cclk n_745 GND efet w=12 l=9
+ ad=0 pd=0 as=183 ps=62 
M3160 Vdd n_1593 n_1593 GND dfet w=9 l=12
+ ad=0 pd=0 as=1492 ps=462 
M3161 GND n_226 n_1593 GND efet w=74 l=7
+ ad=0 pd=0 as=714 ps=204 
M3162 n_772 n_1674 GND GND efet w=73 l=6
+ ad=634 pd=220 as=0 ps=0 
M3163 Vdd n_772 n_772 GND dfet w=9 l=11
+ ad=0 pd=0 as=1304 ps=452 
M3164 GND n_1593 n_1552 GND efet w=24 l=6
+ ad=0 pd=0 as=345 ps=106 
M3165 GND n_772 n_1305 GND efet w=24 l=6
+ ad=0 pd=0 as=377 ps=110 
M3166 n_1552 n_1552 Vdd GND dfet w=8 l=14
+ ad=1393 pd=396 as=0 ps=0 
M3167 Vdd n_1593 dpc14_SRS GND dfet w=8 l=9
+ ad=0 pd=0 as=864 ps=232 
M3168 n_1305 n_1305 Vdd GND dfet w=10 l=14
+ ad=1378 pd=402 as=0 ps=0 
M3169 dpc14_SRS n_1552 GND GND efet w=120 l=6
+ ad=0 pd=0 as=0 ps=0 
M3170 dpc17_SUMS n_1305 GND GND efet w=122 l=7
+ ad=1093 pd=322 as=0 ps=0 
M3171 Vdd n_772 dpc17_SUMS GND dfet w=11 l=9
+ ad=0 pd=0 as=0 ps=0 
M3172 Vdd n_1499 n_1499 GND dfet w=9 l=12
+ ad=0 pd=0 as=1310 ps=450 
M3173 GND n_1450 n_1499 GND efet w=76 l=6
+ ad=0 pd=0 as=818 ps=222 
M3174 n_906 n_1333 GND GND efet w=76 l=6
+ ad=823 pd=226 as=0 ps=0 
M3175 Vdd n_906 n_906 GND dfet w=9 l=10
+ ad=0 pd=0 as=1950 ps=632 
M3176 Vdd n_154 n_154 GND dfet w=9 l=12
+ ad=0 pd=0 as=1289 ps=446 
M3177 n_714 n_906 GND GND efet w=43 l=5
+ ad=492 pd=142 as=0 ps=0 
M3178 GND n_1499 n_709 GND efet w=24 l=6
+ ad=0 pd=0 as=352 ps=108 
M3179 GND n_512 n_154 GND efet w=74 l=7
+ ad=0 pd=0 as=663 ps=218 
M3180 n_241 n_745 GND GND efet w=73 l=6
+ ad=682 pd=204 as=0 ps=0 
M3181 Vdd n_241 n_241 GND dfet w=8 l=10
+ ad=0 pd=0 as=1418 ps=450 
M3182 GND n_154 n_75 GND efet w=25 l=6
+ ad=0 pd=0 as=376 ps=112 
M3183 GND n_241 n_1033 GND efet w=24 l=6
+ ad=0 pd=0 as=336 ps=104 
M3184 n_709 n_709 Vdd GND dfet w=9 l=14
+ ad=1314 pd=404 as=0 ps=0 
M3185 Vdd n_1499 dpc18_nDAA GND dfet w=9 l=9
+ ad=0 pd=0 as=1263 ps=352 
M3186 n_714 n_714 Vdd GND dfet w=9 l=15
+ ad=705 pd=190 as=0 ps=0 
M3187 adl0 dpc10_ADLADD alub0 GND efet w=11 l=7
+ ad=0 pd=0 as=562 ps=144 
M3188 alub0 dpc8_nDBADD n_624 GND efet w=11 l=7
+ ad=0 pd=0 as=884 ps=274 
M3189 alub0 dpc9_DBADD idb0 GND efet w=11 l=7
+ ad=0 pd=0 as=2127 ps=558 
M3190 GND idb0 n_624 GND efet w=60 l=7
+ ad=0 pd=0 as=0 ps=0 
M3191 n_624 n_624 Vdd GND dfet w=10 l=18
+ ad=358 pd=88 as=0 ps=0 
M3192 n_316 alua0 GND GND efet w=61 l=6
+ ad=305 pd=132 as=0 ps=0 
M3193 nA_B0 alub0 n_316 GND efet w=61 l=7
+ ad=1049 pd=290 as=0 ps=0 
M3194 Vdd nA_B0 nA_B0 GND dfet w=10 l=22
+ ad=0 pd=0 as=2507 ps=772 
M3195 naluresult0 dpc13_ORS n_A_B_0 GND efet w=13 l=8
+ ad=1631 pd=444 as=1074 ps=288 
M3196 GND dpc12_0ADD alua0 GND efet w=13 l=6
+ ad=0 pd=0 as=555 ps=144 
M3197 alua0 dpc11_SBADD sb0 GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M3198 adl1 dpc10_ADLADD alub1 GND efet w=11 l=7
+ ad=0 pd=0 as=579 ps=144 
M3199 alub1 dpc8_nDBADD n_583 GND efet w=12 l=8
+ ad=0 pd=0 as=981 ps=278 
M3200 alub1 dpc9_DBADD idb1 GND efet w=12 l=7
+ ad=0 pd=0 as=2139 ps=552 
M3201 GND idb1 n_583 GND efet w=61 l=7
+ ad=0 pd=0 as=0 ps=0 
M3202 n_583 n_583 Vdd GND dfet w=8 l=17
+ ad=332 pd=86 as=0 ps=0 
M3203 n_A_B_0 alua0 GND GND efet w=32 l=6
+ ad=0 pd=0 as=0 ps=0 
M3204 GND alub0 n_A_B_0 GND efet w=32 l=7
+ ad=0 pd=0 as=0 ps=0 
M3205 Vdd n_A_B_0 n_A_B_0 GND dfet w=10 l=23
+ ad=0 pd=0 as=2377 ps=764 
M3206 n_189 alua1 GND GND efet w=61 l=6
+ ad=366 pd=134 as=0 ps=0 
M3207 nA_B1 alub1 n_189 GND efet w=61 l=6
+ ad=1110 pd=296 as=0 ps=0 
M3208 Vdd nA_B1 nA_B1 GND dfet w=9 l=22
+ ad=0 pd=0 as=932 ps=242 
M3209 A_B0 A_B0 Vdd GND dfet w=10 l=15
+ ad=887 pd=262 as=0 ps=0 
M3210 GND n_709 dpc18_nDAA GND efet w=122 l=6
+ ad=0 pd=0 as=0 ps=0 
M3211 dpc19_ADDSB7 n_906 GND GND efet w=114 l=6
+ ad=1025 pd=310 as=0 ps=0 
M3212 Vdd n_714 dpc19_ADDSB7 GND dfet w=10 l=9
+ ad=0 pd=0 as=0 ps=0 
M3213 n_75 n_75 Vdd GND dfet w=9 l=14
+ ad=1295 pd=392 as=0 ps=0 
M3214 Vdd n_154 dpc20_ADDSB06 GND dfet w=9 l=9
+ ad=0 pd=0 as=1108 ps=322 
M3215 n_1033 n_1033 Vdd GND dfet w=9 l=15
+ ad=1333 pd=378 as=0 ps=0 
M3216 GND n_75 dpc20_ADDSB06 GND efet w=118 l=6
+ ad=0 pd=0 as=0 ps=0 
M3217 dpc21_ADDADL n_1033 GND GND efet w=111 l=6
+ ad=1007 pd=302 as=0 ps=0 
M3218 Vdd n_241 dpc21_ADDADL GND dfet w=9 l=8
+ ad=0 pd=0 as=0 ps=0 
M3219 Vdd n_105 n_105 GND dfet w=10 l=16
+ ad=0 pd=0 as=1218 ps=344 
M3220 n_105 notalucin GND GND efet w=18 l=6
+ ad=318 pd=98 as=0 ps=0 
M3221 A_B0 n_A_B_0 GND GND efet w=18 l=6
+ ad=336 pd=92 as=0 ps=0 
M3222 n_1348 A_B0 n_AxB_0 GND efet w=36 l=6
+ ad=189 pd=82 as=769 ps=236 
M3223 naluresult0 dpc15_ANDS nA_B0 GND efet w=11 l=8
+ ad=0 pd=0 as=0 ps=0 
M3224 n_AxB_0 dpc16_EORS naluresult0 GND efet w=11 l=8
+ ad=0 pd=0 as=0 ps=0 
M3225 nA_B1 dpc14_SRS naluresult0 GND efet w=11 l=8
+ ad=0 pd=0 as=0 ps=0 
M3226 naluresult1 dpc13_ORS n_A_B_1 GND efet w=12 l=8
+ ad=1883 pd=500 as=1061 ps=282 
M3227 GND dpc12_0ADD alua1 GND efet w=12 l=6
+ ad=0 pd=0 as=563 ps=140 
M3228 alua1 dpc11_SBADD sb1 GND efet w=12 l=9
+ ad=0 pd=0 as=0 ps=0 
M3229 n_1389 dpc7_SS s2 GND efet w=12 l=7
+ ad=0 pd=0 as=345 ps=78 
M3230 s2 dpc6_SBS sb2 GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M3231 sb2 cclk Vdd GND efet w=23 l=7
+ ad=0 pd=0 as=0 ps=0 
M3232 Vdd n_998 n_998 GND dfet w=9 l=16
+ ad=0 pd=0 as=363 ps=102 
M3233 n_998 dpc5_SADL adl3 GND efet w=15 l=6
+ ad=1989 pd=464 as=2512 ps=628 
M3234 Vdd n_34 n_34 GND dfet w=9 l=20
+ ad=0 pd=0 as=482 ps=130 
M3235 x3 dpc3_SBX sb3 GND efet w=12 l=7
+ ad=0 pd=0 as=0 ps=0 
M3236 Vdd n_436 n_436 GND dfet w=10 l=16
+ ad=0 pd=0 as=304 ps=80 
M3237 n_998 dpc4_SSB sb3 GND efet w=16 l=7
+ ad=0 pd=0 as=0 ps=0 
M3238 GND notx4 n_436 GND efet w=56 l=7
+ ad=0 pd=0 as=1454 ps=352 
M3239 Vdd notx4 notx4 GND dfet w=10 l=21
+ ad=0 pd=0 as=975 ps=258 
M3240 notx4 x4 GND GND efet w=35 l=6
+ ad=524 pd=166 as=0 ps=0 
M3241 x4 cclk n_436 GND efet w=11 l=8
+ ad=262 pd=92 as=0 ps=0 
M3242 GND nots3 n_998 GND efet w=44 l=6
+ ad=0 pd=0 as=0 ps=0 
M3243 n_34 s3 GND GND efet w=34 l=6
+ ad=919 pd=228 as=0 ps=0 
M3244 n_34 cclk nots3 GND efet w=11 l=8
+ ad=0 pd=0 as=289 ps=100 
M3245 n_998 dpc7_SS s3 GND efet w=11 l=8
+ ad=0 pd=0 as=334 ps=76 
M3246 s3 dpc6_SBS sb3 GND efet w=12 l=7
+ ad=0 pd=0 as=0 ps=0 
M3247 sb3 cclk Vdd GND efet w=22 l=6
+ ad=0 pd=0 as=0 ps=0 
M3248 Vdd n_3 n_3 GND dfet w=9 l=17
+ ad=0 pd=0 as=358 ps=100 
M3249 n_3 dpc5_SADL adl4 GND efet w=14 l=7
+ ad=1943 pd=454 as=2433 ps=608 
M3250 Vdd n_973 n_973 GND dfet w=9 l=21
+ ad=0 pd=0 as=500 ps=132 
M3251 n_436 dpc2_XSB sb4 GND efet w=13 l=7
+ ad=0 pd=0 as=0 ps=0 
M3252 x4 dpc3_SBX sb4 GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M3253 Vdd n_578 n_578 GND dfet w=9 l=16
+ ad=0 pd=0 as=294 ps=80 
M3254 GND notx5 n_578 GND efet w=56 l=7
+ ad=0 pd=0 as=1571 ps=356 
M3255 Vdd notx5 notx5 GND dfet w=9 l=21
+ ad=0 pd=0 as=965 ps=256 
M3256 notx5 x5 GND GND efet w=36 l=7
+ ad=521 pd=168 as=0 ps=0 
M3257 x5 cclk n_578 GND efet w=11 l=8
+ ad=264 pd=92 as=0 ps=0 
M3258 n_3 dpc4_SSB sb4 GND efet w=16 l=9
+ ad=0 pd=0 as=0 ps=0 
M3259 GND nots4 n_3 GND efet w=44 l=6
+ ad=0 pd=0 as=0 ps=0 
M3260 n_973 s4 GND GND efet w=34 l=6
+ ad=886 pd=230 as=0 ps=0 
M3261 n_973 cclk nots4 GND efet w=12 l=8
+ ad=0 pd=0 as=283 ps=98 
M3262 n_3 dpc7_SS s4 GND efet w=11 l=8
+ ad=0 pd=0 as=322 ps=74 
M3263 s4 dpc6_SBS sb4 GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M3264 sb4 cclk Vdd GND efet w=23 l=7
+ ad=0 pd=0 as=0 ps=0 
M3265 Vdd n_280 n_280 GND dfet w=9 l=16
+ ad=0 pd=0 as=359 ps=102 
M3266 n_280 dpc5_SADL adl5 GND efet w=15 l=6
+ ad=1941 pd=454 as=2491 ps=618 
M3267 Vdd n_496 n_496 GND dfet w=9 l=20
+ ad=0 pd=0 as=468 ps=128 
M3268 n_578 dpc2_XSB sb5 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M3269 x5 dpc3_SBX sb5 GND efet w=11 l=8
+ ad=0 pd=0 as=0 ps=0 
M3270 GND noty6 n_518 GND efet w=57 l=7
+ ad=0 pd=0 as=1474 ps=356 
M3271 Vdd noty6 noty6 GND dfet w=10 l=20
+ ad=0 pd=0 as=957 ps=256 
M3272 noty6 y6 GND GND efet w=35 l=6
+ ad=541 pd=168 as=0 ps=0 
M3273 y6 cclk n_518 GND efet w=11 l=8
+ ad=260 pd=92 as=0 ps=0 
M3274 n_1548 n_1548 Vdd GND dfet w=9 l=10
+ ad=240 pd=74 as=0 ps=0 
M3275 n_518 dpc0_YSB sb6 GND efet w=13 l=8
+ ad=0 pd=0 as=4155 ps=988 
M3276 y6 dpc1_SBY sb6 GND efet w=11 l=7
+ ad=0 pd=0 as=0 ps=0 
M3277 nABL7 cclk n_171 GND efet w=12 l=8
+ ad=294 pd=94 as=0 ps=0 
M3278 n_577 ADL_ABL nABL7 GND efet w=12 l=7
+ ad=84 pd=38 as=0 ps=0 
M3279 n_1046 cp1 n_577 GND efet w=12 l=7
+ ad=1036 pd=260 as=0 ps=0 
M3280 abl7 nABL7 GND GND efet w=95 l=6
+ ad=964 pd=256 as=0 ps=0 
M3281 abl7 abl7 Vdd GND dfet w=9 l=14
+ ad=2772 pd=836 as=0 ps=0 
M3282 Vdd n_1668 n_1668 GND dfet w=9 l=10
+ ad=0 pd=0 as=327 ps=104 
M3283 GND adh0 n_1668 GND efet w=77 l=7
+ ad=0 pd=0 as=1123 ps=270 
M3284 abh0 nABH0 GND GND efet w=66 l=7
+ ad=515 pd=196 as=0 ps=0 
M3285 GND adl7 n_1046 GND efet w=81 l=6
+ ad=0 pd=0 as=0 ps=0 
M3286 Vdd n_1251 n_1251 GND dfet w=10 l=16
+ ad=0 pd=0 as=294 ps=80 
M3287 GND noty7 n_1251 GND efet w=56 l=7
+ ad=0 pd=0 as=1557 ps=350 
M3288 Vdd noty7 noty7 GND dfet w=9 l=20
+ ad=0 pd=0 as=957 ps=256 
M3289 noty7 y7 GND GND efet w=35 l=7
+ ad=531 pd=168 as=0 ps=0 
M3290 y7 cclk n_1251 GND efet w=11 l=8
+ ad=260 pd=90 as=0 ps=0 
M3291 n_1046 n_1046 Vdd GND dfet w=10 l=11
+ ad=237 pd=72 as=0 ps=0 
M3292 n_1251 dpc0_YSB sb7 GND efet w=14 l=8
+ ad=0 pd=0 as=4081 ps=1000 
M3293 y7 dpc1_SBY sb7 GND efet w=11 l=8
+ ad=0 pd=0 as=0 ps=0 
M3294 Vdd n_1724 n_1724 GND dfet w=10 l=16
+ ad=0 pd=0 as=304 ps=80 
M3295 GND notx6 n_1724 GND efet w=56 l=7
+ ad=0 pd=0 as=1563 ps=352 
M3296 Vdd notx6 notx6 GND dfet w=9 l=20
+ ad=0 pd=0 as=945 ps=256 
M3297 n_280 dpc4_SSB sb5 GND efet w=16 l=8
+ ad=0 pd=0 as=0 ps=0 
M3298 notx6 x6 GND GND efet w=36 l=6
+ ad=573 pd=170 as=0 ps=0 
M3299 x6 cclk n_1724 GND efet w=12 l=8
+ ad=270 pd=90 as=0 ps=0 
M3300 GND nots5 n_280 GND efet w=44 l=6
+ ad=0 pd=0 as=0 ps=0 
M3301 n_496 s5 GND GND efet w=33 l=6
+ ad=900 pd=228 as=0 ps=0 
M3302 n_496 cclk nots5 GND efet w=12 l=8
+ ad=0 pd=0 as=283 ps=98 
M3303 n_280 dpc7_SS s5 GND efet w=11 l=8
+ ad=0 pd=0 as=328 ps=76 
M3304 s5 dpc6_SBS sb5 GND efet w=12 l=7
+ ad=0 pd=0 as=0 ps=0 
M3305 sb5 cclk Vdd GND efet w=23 l=7
+ ad=0 pd=0 as=0 ps=0 
M3306 Vdd n_618 n_618 GND dfet w=9 l=17
+ ad=0 pd=0 as=358 ps=100 
M3307 n_618 dpc5_SADL adl6 GND efet w=15 l=5
+ ad=1885 pd=454 as=2476 ps=616 
M3308 Vdd n_1187 n_1187 GND dfet w=10 l=20
+ ad=0 pd=0 as=457 ps=130 
M3309 n_1724 dpc2_XSB sb6 GND efet w=13 l=7
+ ad=0 pd=0 as=0 ps=0 
M3310 x6 dpc3_SBX sb6 GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M3311 Vdd n_871 n_871 GND dfet w=10 l=16
+ ad=0 pd=0 as=294 ps=80 
M3312 GND notx7 n_871 GND efet w=57 l=7
+ ad=0 pd=0 as=1449 ps=354 
M3313 Vdd notx7 notx7 GND dfet w=10 l=20
+ ad=0 pd=0 as=957 ps=256 
M3314 notx7 x7 GND GND efet w=34 l=6
+ ad=538 pd=168 as=0 ps=0 
M3315 x7 cclk n_871 GND efet w=11 l=8
+ ad=264 pd=90 as=0 ps=0 
M3316 n_871 dpc2_XSB sb7 GND efet w=13 l=8
+ ad=0 pd=0 as=0 ps=0 
M3317 n_618 dpc4_SSB sb6 GND efet w=17 l=9
+ ad=0 pd=0 as=0 ps=0 
M3318 GND nots6 n_618 GND efet w=45 l=7
+ ad=0 pd=0 as=0 ps=0 
M3319 n_1187 s6 GND GND efet w=33 l=6
+ ad=849 pd=230 as=0 ps=0 
M3320 n_1187 cclk nots6 GND efet w=11 l=8
+ ad=0 pd=0 as=273 ps=94 
M3321 adl2 dpc10_ADLADD alub2 GND efet w=12 l=8
+ ad=0 pd=0 as=593 ps=148 
M3322 alub2 dpc8_nDBADD n_458 GND efet w=12 l=7
+ ad=0 pd=0 as=965 ps=276 
M3323 alub2 dpc9_DBADD idb2 GND efet w=12 l=7
+ ad=0 pd=0 as=2131 ps=558 
M3324 GND idb2 n_458 GND efet w=60 l=7
+ ad=0 pd=0 as=0 ps=0 
M3325 n_458 n_458 Vdd GND dfet w=9 l=17
+ ad=332 pd=86 as=0 ps=0 
M3326 n_A_B_1 alua1 GND GND efet w=31 l=6
+ ad=0 pd=0 as=0 ps=0 
M3327 GND alub1 n_A_B_1 GND efet w=31 l=7
+ ad=0 pd=0 as=0 ps=0 
M3328 Vdd n_A_B_1 n_A_B_1 GND dfet w=9 l=23
+ ad=0 pd=0 as=1402 ps=412 
M3329 naluresult1 dpc15_ANDS nA_B1 GND efet w=11 l=8
+ ad=0 pd=0 as=0 ps=0 
M3330 n_452 alua2 GND GND efet w=61 l=7
+ ad=305 pd=132 as=0 ps=0 
M3331 nA_B2 alub2 n_452 GND efet w=61 l=7
+ ad=1140 pd=302 as=0 ps=0 
M3332 Vdd nA_B2 nA_B2 GND dfet w=10 l=21
+ ad=0 pd=0 as=2310 ps=710 
M3333 GND nA_B0 n_1348 GND efet w=34 l=7
+ ad=0 pd=0 as=0 ps=0 
M3334 C01 n_A_B_0 GND GND efet w=28 l=6
+ ad=1033 pd=264 as=0 ps=0 
M3335 n_942 nA_B0 C01 GND efet w=56 l=6
+ ad=479 pd=162 as=0 ps=0 
M3336 GND notalucin n_942 GND efet w=73 l=6
+ ad=0 pd=0 as=0 ps=0 
M3337 n_406 n_AxB_0 GND GND efet w=35 l=7
+ ad=175 pd=80 as=0 ps=0 
M3338 n_AxBxC_0 n_105 n_406 GND efet w=35 l=7
+ ad=837 pd=218 as=0 ps=0 
M3339 Vdd n_AxBxC_0 n_AxBxC_0 GND dfet w=9 l=18
+ ad=0 pd=0 as=456 ps=104 
M3340 GND n_134 n_467 GND efet w=26 l=6
+ ad=0 pd=0 as=917 ps=212 
M3341 GND n_236 n_1427 GND efet w=39 l=6
+ ad=0 pd=0 as=0 ps=0 
M3342 GND n_470 n_467 GND efet w=29 l=5
+ ad=0 pd=0 as=0 ps=0 
M3343 n_930 n_1276 GND GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M3344 n_180 n_180 Vdd GND dfet w=10 l=12
+ ad=971 pd=292 as=0 ps=0 
M3345 n_501 n_501 Vdd GND dfet w=9 l=12
+ ad=1783 pd=640 as=0 ps=0 
M3346 n_501 n_180 GND GND efet w=38 l=6
+ ad=0 pd=0 as=0 ps=0 
M3347 n_180 notRdy0 GND GND efet w=41 l=7
+ ad=0 pd=0 as=0 ps=0 
M3348 GND op_T3_branch n_1708 GND efet w=38 l=7
+ ad=0 pd=0 as=651 ps=186 
M3349 n_1716 op_T3_branch GND GND efet w=30 l=6
+ ad=1725 pd=408 as=0 ps=0 
M3350 GND n_510 n_1716 GND efet w=31 l=6
+ ad=0 pd=0 as=0 ps=0 
M3351 n_510 n_347 GND GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M3352 GND op_rmw n_510 GND efet w=33 l=7
+ ad=0 pd=0 as=0 ps=0 
M3353 Vdd op_rmw op_rmw GND dfet w=8 l=13
+ ad=0 pd=0 as=641 ps=178 
M3354 n_510 n_510 Vdd GND dfet w=10 l=16
+ ad=801 pd=248 as=0 ps=0 
M3355 op_rmw n_790 GND GND efet w=37 l=7
+ ad=404 pd=124 as=0 ps=0 
M3356 n_335 nop_store GND GND efet w=88 l=6
+ ad=1094 pd=326 as=0 ps=0 
M3357 GND n_368 n_218 GND efet w=38 l=7
+ ad=0 pd=0 as=819 ps=232 
M3358 n_368 n_368 Vdd GND dfet w=11 l=16
+ ad=813 pd=244 as=0 ps=0 
M3359 n_790 n_790 Vdd GND dfet w=9 l=16
+ ad=2930 pd=964 as=0 ps=0 
M3360 Vdd n_218 n_218 GND dfet w=10 l=10
+ ad=0 pd=0 as=745 ps=262 
M3361 GND n_347 n_335 GND efet w=87 l=7
+ ad=0 pd=0 as=0 ps=0 
M3362 n_1708 n_1708 Vdd GND dfet w=10 l=13
+ ad=4739 pd=1630 as=0 ps=0 
M3363 n_1716 n_1716 Vdd GND dfet w=10 l=13
+ ad=2265 pd=758 as=0 ps=0 
M3364 Vdd n_944 n_944 GND dfet w=10 l=12
+ ad=0 pd=0 as=327 ps=94 
M3365 GND n_1449 n_944 GND efet w=50 l=7
+ ad=0 pd=0 as=1416 ps=358 
M3366 GND n_1708 n_236 GND efet w=65 l=6
+ ad=0 pd=0 as=717 ps=174 
M3367 n_944 cclk pipeUNK37 GND efet w=14 l=7
+ ad=0 pd=0 as=156 ps=76 
M3368 GND pipeUNK37 n_198 GND efet w=93 l=6
+ ad=0 pd=0 as=1043 ps=274 
M3369 n_198 pipeUNK37 GND GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M3370 GND n_759 n_944 GND efet w=78 l=6
+ ad=0 pd=0 as=0 ps=0 
M3371 n_236 n_236 Vdd GND dfet w=9 l=8
+ ad=7578 pd=2500 as=0 ps=0 
M3372 n_501 n_819 GND GND efet w=42 l=6
+ ad=0 pd=0 as=0 ps=0 
M3373 GND op_T2_abs_access n_773 GND efet w=32 l=6
+ ad=0 pd=0 as=776 ps=208 
M3374 n_1272 cp1 notRdy0 GND efet w=11 l=8
+ ad=385 pd=140 as=0 ps=0 
M3375 n_773 n_646 GND GND efet w=44 l=7
+ ad=0 pd=0 as=0 ps=0 
M3376 n_773 n_773 Vdd GND dfet w=9 l=13
+ ad=1131 pd=342 as=0 ps=0 
M3377 Vdd n_275 n_275 GND dfet w=9 l=11
+ ad=0 pd=0 as=762 ps=212 
M3378 n_275 n_1697 GND GND efet w=50 l=9
+ ad=744 pd=204 as=0 ps=0 
M3379 notRdy0 cp1 n_1276 GND efet w=12 l=8
+ ad=0 pd=0 as=264 ps=66 
M3380 GND n_630 n_1705 GND efet w=28 l=7
+ ad=0 pd=0 as=0 ps=0 
M3381 n_930 n_1276 GND GND efet w=17 l=7
+ ad=0 pd=0 as=0 ps=0 
M3382 Vdd n_1655 n_1655 GND dfet w=9 l=10
+ ad=0 pd=0 as=825 ps=264 
M3383 n_1655 n_1211 GND GND efet w=37 l=6
+ ad=331 pd=104 as=0 ps=0 
M3384 GND n_236 n_176 GND efet w=41 l=6
+ ad=0 pd=0 as=987 ps=300 
M3385 n_176 n_10 GND GND efet w=44 l=6
+ ad=0 pd=0 as=0 ps=0 
M3386 GND n_646 n_272 GND efet w=31 l=6
+ ad=0 pd=0 as=0 ps=0 
M3387 n_1278 n_824 n_1642 GND efet w=84 l=6
+ ad=472 pd=178 as=760 ps=204 
M3388 GND n_462 n_1278 GND efet w=83 l=7
+ ad=0 pd=0 as=0 ps=0 
M3389 n_1642 n_1642 Vdd GND dfet w=10 l=10
+ ad=4432 pd=1610 as=0 ps=0 
M3390 n_182 n_1655 GND GND efet w=27 l=6
+ ad=0 pd=0 as=0 ps=0 
M3391 n_176 n_176 Vdd GND dfet w=10 l=11
+ ad=2638 pd=944 as=0 ps=0 
M3392 Vdd n_952 n_952 GND dfet w=10 l=9
+ ad=0 pd=0 as=3796 ps=1322 
M3393 n_952 n_272 GND GND efet w=56 l=7
+ ad=812 pd=254 as=0 ps=0 
M3394 n_182 n_646 GND GND efet w=44 l=6
+ ad=0 pd=0 as=0 ps=0 
M3395 GND n_930 n_1286 GND efet w=66 l=6
+ ad=0 pd=0 as=1050 ps=238 
M3396 GND n_773 n_275 GND efet w=43 l=6
+ ad=0 pd=0 as=0 ps=0 
M3397 GND n_1272 n_608 GND efet w=52 l=7
+ ad=0 pd=0 as=697 ps=214 
M3398 Vdd n_608 n_608 GND dfet w=9 l=17
+ ad=0 pd=0 as=361 ps=90 
M3399 n_559 cclk n_608 GND efet w=12 l=9
+ ad=214 pd=92 as=0 ps=0 
M3400 Vdd n_916 n_916 GND dfet w=9 l=9
+ ad=0 pd=0 as=2489 ps=838 
M3401 GND n_275 n_104 GND efet w=39 l=8
+ ad=0 pd=0 as=0 ps=0 
M3402 n_916 n_1517 GND GND efet w=63 l=6
+ ad=1575 pd=378 as=0 ps=0 
M3403 n_387 n_206 n_916 GND efet w=120 l=6
+ ad=653 pd=252 as=0 ps=0 
M3404 GND n_853 n_387 GND efet w=120 l=6
+ ad=0 pd=0 as=0 ps=0 
M3405 notRdy0 n_198 GND GND efet w=136 l=7
+ ad=0 pd=0 as=0 ps=0 
M3406 nWR op_T4_brk GND GND efet w=35 l=6
+ ad=3126 pd=730 as=0 ps=0 
M3407 GND op_T2_php_pha nWR GND efet w=35 l=7
+ ad=0 pd=0 as=0 ps=0 
M3408 n_191 n_790 GND GND efet w=39 l=7
+ ad=1078 pd=312 as=0 ps=0 
M3409 n_1065 n_1065 Vdd GND dfet w=10 l=16
+ ad=863 pd=258 as=0 ps=0 
M3410 n_591 n_1258 GND GND efet w=84 l=7
+ ad=507 pd=196 as=0 ps=0 
M3411 nop_set_C op_asl_rol n_591 GND efet w=68 l=6
+ ad=3038 pd=732 as=0 ps=0 
M3412 GND op_T3_mem_zp_idx n_347 GND efet w=37 l=7
+ ad=0 pd=0 as=1693 ps=452 
M3413 nop_set_C x_op_T__adc_sbc GND GND efet w=30 l=6
+ ad=0 pd=0 as=0 ps=0 
M3414 n_327 op_T0_plp GND GND efet w=31 l=7
+ ad=944 pd=258 as=0 ps=0 
M3415 GND x_op_T4_rti n_327 GND efet w=38 l=7
+ ad=0 pd=0 as=0 ps=0 
M3416 nop_set_C op_T__cmp GND GND efet w=26 l=6
+ ad=0 pd=0 as=0 ps=0 
M3417 GND op_T__cpx_cpy_abs nop_set_C GND efet w=25 l=6
+ ad=0 pd=0 as=0 ps=0 
M3418 nop_set_C op_T__asl_rol_a GND GND efet w=34 l=6
+ ad=0 pd=0 as=0 ps=0 
M3419 nop_set_C nop_set_C Vdd GND dfet w=10 l=17
+ ad=948 pd=278 as=0 ps=0 
M3420 GND op_T__cpx_cpy_imm_zp nop_set_C GND efet w=37 l=6
+ ad=0 pd=0 as=0 ps=0 
M3421 n_327 n_327 Vdd GND dfet w=11 l=18
+ ad=895 pd=266 as=0 ps=0 
M3422 GND op_T0_cld_sed n_774 GND efet w=28 l=7
+ ad=0 pd=0 as=1241 ps=314 
M3423 n_347 op_T3_mem_abs GND GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M3424 GND op_T2_mem_zp n_347 GND efet w=33 l=6
+ ad=0 pd=0 as=0 ps=0 
M3425 n_347 op_T5_mem_ind_idx GND GND efet w=40 l=6
+ ad=0 pd=0 as=0 ps=0 
M3426 GND op_T4_mem_abs_idx n_347 GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M3427 Vdd n_1137 n_1137 GND dfet w=9 l=13
+ ad=0 pd=0 as=763 ps=216 
M3428 Vdd nWR nWR GND dfet w=9 l=11
+ ad=0 pd=0 as=263 ps=72 
M3429 GND n_218 n_1716 GND efet w=36 l=5
+ ad=0 pd=0 as=0 ps=0 
M3430 GND n_347 n_191 GND efet w=32 l=6
+ ad=0 pd=0 as=0 ps=0 
M3431 Vdd n_1258 n_1258 GND dfet w=10 l=6
+ ad=0 pd=0 as=4400 ps=1430 
M3432 n_1391 n_1391 Vdd GND dfet w=11 l=15
+ ad=6832 pd=2480 as=0 ps=0 
M3433 n_816 n_790 n_1137 GND efet w=46 l=7
+ ad=432 pd=158 as=725 ps=178 
M3434 GND nop_store n_816 GND efet w=56 l=6
+ ad=0 pd=0 as=0 ps=0 
M3435 n_198 n_198 Vdd GND dfet w=10 l=11
+ ad=1854 pd=558 as=0 ps=0 
M3436 notRnWprepad cp1 n_759 GND efet w=11 l=9
+ ad=0 pd=0 as=153 ps=76 
M3437 Vdd n_424 notRdy0 GND dfet w=18 l=6
+ ad=0 pd=0 as=0 ps=0 
M3438 notRnWprepad notRnWprepad Vdd GND dfet w=9 l=9
+ ad=6826 pd=2258 as=0 ps=0 
M3439 GND n_1258 nWR GND efet w=37 l=6
+ ad=0 pd=0 as=0 ps=0 
M3440 nWR n_335 GND GND efet w=64 l=5
+ ad=0 pd=0 as=0 ps=0 
M3441 GND n_440 nWR GND efet w=54 l=6
+ ad=0 pd=0 as=0 ps=0 
M3442 GND n_1642 nWR GND efet w=36 l=6
+ ad=0 pd=0 as=0 ps=0 
M3443 GND n_1258 n_1716 GND efet w=38 l=6
+ ad=0 pd=0 as=0 ps=0 
M3444 n_191 n_191 Vdd GND dfet w=11 l=11
+ ad=594 pd=222 as=0 ps=0 
M3445 GND notRdy0 n_191 GND efet w=28 l=6
+ ad=0 pd=0 as=0 ps=0 
M3446 Vdd n_1120 n_1120 GND dfet w=10 l=11
+ ad=0 pd=0 as=626 ps=216 
M3447 n_1258 n_390 GND GND efet w=72 l=6
+ ad=789 pd=204 as=0 ps=0 
M3448 n_889 op_T0_clc_sec GND GND efet w=27 l=7
+ ad=885 pd=278 as=0 ps=0 
M3449 n_347 n_347 Vdd GND dfet w=9 l=16
+ ad=4296 pd=1396 as=0 ps=0 
M3450 GND n_1533 clock2 GND efet w=130 l=6
+ ad=0 pd=0 as=2105 ps=460 
M3451 Vdd clock2 clock2 GND dfet w=9 l=6
+ ad=0 pd=0 as=20352 ps=6126 
M3452 n_664 n_664 Vdd GND dfet w=10 l=16
+ ad=727 pd=202 as=0 ps=0 
M3453 GND op_implied n_664 GND efet w=40 l=6
+ ad=0 pd=0 as=598 ps=164 
M3454 GND pd6_clearIR n_1309 GND efet w=72 l=7
+ ad=0 pd=0 as=0 ps=0 
M3455 n_1309 n_1309 Vdd GND dfet w=11 l=7
+ ad=712 pd=260 as=0 ps=0 
M3456 GND notRdy0 n_1180 GND efet w=43 l=7
+ ad=0 pd=0 as=1106 ps=262 
M3457 n_1533 cp1 n_1180 GND efet w=16 l=8
+ ad=164 pd=86 as=0 ps=0 
M3458 n_1180 pipenT0 GND GND efet w=46 l=6
+ ad=0 pd=0 as=0 ps=0 
M3459 n_390 n_653 GND GND efet w=48 l=6
+ ad=537 pd=130 as=0 ps=0 
M3460 Vdd n_390 n_390 GND dfet w=9 l=21
+ ad=0 pd=0 as=1553 ps=444 
M3461 n_889 n_889 Vdd GND dfet w=12 l=20
+ ad=468 pd=126 as=0 ps=0 
M3462 Vdd n_1180 n_1180 GND dfet w=9 l=17
+ ad=0 pd=0 as=435 ps=102 
M3463 n_653 cp1 n_1497 GND efet w=13 l=8
+ ad=168 pd=72 as=916 ps=272 
M3464 GND n_1533 n_964 GND efet w=55 l=7
+ ad=0 pd=0 as=974 ps=222 
M3465 n_1497 pipeUNK41 GND GND efet w=51 l=6
+ ad=0 pd=0 as=0 ps=0 
M3466 n_191 cclk pipeUNK40 GND efet w=13 l=9
+ ad=0 pd=0 as=153 ps=64 
M3467 nWR cclk pipenWR_phi2 GND efet w=12 l=8
+ ad=0 pd=0 as=281 ps=92 
M3468 GND C1x5Reset notRnWprepad GND efet w=70 l=6
+ ad=0 pd=0 as=0 ps=0 
M3469 Vdd n_424 n_424 GND dfet w=10 l=7
+ ad=0 pd=0 as=679 ps=252 
M3470 n_424 n_198 GND GND efet w=60 l=6
+ ad=956 pd=228 as=0 ps=0 
M3471 GND Reset0 n_14 GND efet w=20 l=7
+ ad=0 pd=0 as=1796 ps=432 
M3472 GND n_666 n_862 GND efet w=151 l=6
+ ad=0 pd=0 as=0 ps=0 
M3473 notRnWprepad notRdy0 GND GND efet w=55 l=6
+ ad=0 pd=0 as=0 ps=0 
M3474 n_14 n_14 Vdd GND dfet w=10 l=19
+ ad=1974 pd=694 as=0 ps=0 
M3475 n_862 n_862 Vdd GND dfet w=9 l=8
+ ad=14778 pd=4932 as=0 ps=0 
M3476 n_109 n_1380 GND GND efet w=91 l=6
+ ad=1150 pd=348 as=0 ps=0 
M3477 notRnWprepad pipenWR_phi2 GND GND efet w=87 l=6
+ ad=0 pd=0 as=0 ps=0 
M3478 n_104 op_T4_jmp GND GND efet w=42 l=6
+ ad=0 pd=0 as=0 ps=0 
M3479 n_964 pipenT0 GND GND efet w=46 l=6
+ ad=0 pd=0 as=0 ps=0 
M3480 GND n_664 n_1697 GND efet w=32 l=7
+ ad=0 pd=0 as=780 ps=204 
M3481 Vdd n_409 n_409 GND dfet w=12 l=6
+ ad=0 pd=0 as=1821 ps=598 
M3482 Vdd n_1497 n_1497 GND dfet w=10 l=16
+ ad=0 pd=0 as=627 ps=170 
M3483 n_889 cclk pipeUNK42 GND efet w=12 l=8
+ ad=0 pd=0 as=278 ps=68 
M3484 pipenT0 cclk n_17 GND efet w=12 l=8
+ ad=453 pd=130 as=985 ps=200 
M3485 pipeUNK41 cclk n_504 GND efet w=12 l=8
+ ad=230 pd=82 as=1249 ps=310 
M3486 Vdd n_964 n_964 GND dfet w=10 l=16
+ ad=0 pd=0 as=1493 ps=444 
M3487 n_1697 n_1697 Vdd GND dfet w=10 l=11
+ ad=1464 pd=440 as=0 ps=0 
M3488 nTWOCYCLE PD_xxx010x1 GND GND efet w=48 l=6
+ ad=2074 pd=532 as=0 ps=0 
M3489 Vdd n_1641 n_1641 GND dfet w=12 l=7
+ ad=0 pd=0 as=1531 ps=512 
M3490 GND pd0_clearIR n_409 GND efet w=76 l=6
+ ad=0 pd=0 as=0 ps=0 
M3491 n_1641 pd1_clearIR GND GND efet w=75 l=6
+ ad=0 pd=0 as=0 ps=0 
M3492 Vdd n_1605 n_1605 GND dfet w=12 l=6
+ ad=0 pd=0 as=2192 ps=736 
M3493 Vdd n_227 n_227 GND dfet w=12 l=6
+ ad=0 pd=0 as=976 ps=326 
M3494 GND pd7_clearIR n_1605 GND efet w=74 l=6
+ ad=0 pd=0 as=0 ps=0 
M3495 n_227 pd4_clearIR GND GND efet w=72 l=6
+ ad=0 pd=0 as=0 ps=0 
M3496 clock1 n_964 GND GND efet w=84 l=6
+ ad=1387 pd=224 as=0 ps=0 
M3497 GND n_964 n_17 GND efet w=37 l=7
+ ad=0 pd=0 as=0 ps=0 
M3498 GND n_440 n_812 GND efet w=62 l=7
+ ad=0 pd=0 as=775 ps=222 
M3499 n_104 n_440 GND GND efet w=40 l=6
+ ad=0 pd=0 as=0 ps=0 
M3500 n_812 n_646 GND GND efet w=61 l=6
+ ad=0 pd=0 as=0 ps=0 
M3501 Vdd n_109 n_109 GND dfet w=9 l=6
+ ad=0 pd=0 as=3185 ps=1092 
M3502 n_770 n_559 GND GND efet w=54 l=7
+ ad=529 pd=170 as=0 ps=0 
M3503 n_666 cp1 n_1380 GND efet w=12 l=8
+ ad=147 pd=68 as=1202 ps=320 
M3504 GND notRdy0 n_1718 GND efet w=40 l=6
+ ad=0 pd=0 as=680 ps=196 
M3505 GND notRdy0 n_1120 GND efet w=35 l=6
+ ad=0 pd=0 as=727 ps=204 
M3506 n_137 n_1120 GND GND efet w=34 l=6
+ ad=204 pd=80 as=0 ps=0 
M3507 n_504 n_440 n_137 GND efet w=34 l=6
+ ad=0 pd=0 as=0 ps=0 
M3508 Vdd n_504 n_504 GND dfet w=10 l=15
+ ad=0 pd=0 as=426 ps=116 
M3509 n_17 n_17 Vdd GND dfet w=9 l=9
+ ad=1605 pd=524 as=0 ps=0 
M3510 n_1065 cclk n_1124 GND efet w=15 l=8
+ ad=0 pd=0 as=285 ps=68 
M3511 n_17 n_732 GND GND efet w=37 l=7
+ ad=0 pd=0 as=0 ps=0 
M3512 clock1 n_732 GND GND efet w=75 l=7
+ ad=0 pd=0 as=0 ps=0 
M3513 Vdd n_17 clock1 GND dfet w=11 l=7
+ ad=0 pd=0 as=0 ps=0 
M3514 GND PD_1xx000x0 nTWOCYCLE GND efet w=45 l=6
+ ad=0 pd=0 as=0 ps=0 
M3515 PD_xxx010x1 PD_xxx010x1 Vdd GND dfet w=10 l=10
+ ad=1023 pd=348 as=0 ps=0 
M3516 n_928 n_928 Vdd GND dfet w=12 l=6
+ ad=870 pd=294 as=0 ps=0 
M3517 Vdd n_1083 n_1083 GND dfet w=12 l=7
+ ad=0 pd=0 as=1714 ps=608 
M3518 Vdd n_571 n_571 GND dfet w=13 l=6
+ ad=0 pd=0 as=986 ps=358 
M3519 GND pd3_clearIR n_1083 GND efet w=75 l=7
+ ad=0 pd=0 as=0 ps=0 
M3520 n_571 pd2_clearIR GND GND efet w=72 l=6
+ ad=0 pd=0 as=0 ps=0 
M3521 GND pd5_clearIR n_928 GND efet w=89 l=7
+ ad=0 pd=0 as=0 ps=0 
M3522 nTWOCYCLE PD_xxxx10x0 n_1515 GND efet w=101 l=5
+ ad=0 pd=0 as=755 ps=216 
M3523 Vdd nTWOCYCLE nTWOCYCLE GND dfet w=9 l=10
+ ad=0 pd=0 as=933 ps=304 
M3524 n_646 n_17 GND GND efet w=65 l=6
+ ad=999 pd=212 as=0 ps=0 
M3525 nTWOCYCLE cp1 nTWOCYCLE_phi1 GND efet w=14 l=7
+ ad=0 pd=0 as=167 ps=84 
M3526 n_1039 pipeUNK40 GND GND efet w=60 l=7
+ ad=1132 pd=308 as=0 ps=0 
M3527 n_2 notRdy0 n_1039 GND efet w=53 l=6
+ ad=814 pd=242 as=0 ps=0 
M3528 GND pipeUNK39 n_2 GND efet w=85 l=7
+ ad=0 pd=0 as=0 ps=0 
M3529 n_440 cclk pipeUNK39 GND efet w=12 l=8
+ ad=1270 pd=382 as=183 ps=76 
M3530 n_253 pipeUNK42 GND GND efet w=45 l=7
+ ad=809 pd=198 as=0 ps=0 
M3531 n_1718 n_1718 Vdd GND dfet w=9 l=17
+ ad=1146 pd=372 as=0 ps=0 
M3532 n_770 n_770 Vdd GND dfet w=9 l=17
+ ad=1668 pd=540 as=0 ps=0 
M3533 Vdd n_586 n_586 GND dfet w=8 l=10
+ ad=0 pd=0 as=1328 ps=466 
M3534 n_1330 BRtaken n_586 GND efet w=49 l=7
+ ad=655 pd=178 as=2141 ps=678 
M3535 n_1286 n_470 GND GND efet w=40 l=7
+ ad=0 pd=0 as=0 ps=0 
M3536 n_470 n_646 GND GND efet w=52 l=7
+ ad=600 pd=186 as=0 ps=0 
M3537 n_1286 n_1286 Vdd GND dfet w=10 l=10
+ ad=2206 pd=734 as=0 ps=0 
M3538 n_1448 n_1427 GND GND efet w=35 l=7
+ ad=450 pd=146 as=0 ps=0 
M3539 n_1330 BRtaken n_586 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M3540 GND nnT2BR n_1330 GND efet w=72 l=6
+ ad=0 pd=0 as=0 ps=0 
M3541 n_853 n_770 GND GND efet w=22 l=7
+ ad=300 pd=98 as=0 ps=0 
M3542 n_1409 cp1 n_916 GND efet w=12 l=8
+ ad=245 pd=90 as=0 ps=0 
M3543 n_853 n_853 Vdd GND dfet w=10 l=16
+ ad=2239 pd=668 as=0 ps=0 
M3544 n_1380 n_1154 GND GND efet w=65 l=7
+ ad=0 pd=0 as=0 ps=0 
M3545 GND n_819 n_1380 GND efet w=52 l=7
+ ad=0 pd=0 as=0 ps=0 
M3546 n_781 notRdy0 GND GND efet w=15 l=7
+ ad=1598 pd=418 as=0 ps=0 
M3547 n_781 notRdy0 GND GND efet w=17 l=7
+ ad=0 pd=0 as=0 ps=0 
M3548 n_1055 n_1708 GND GND efet w=42 l=6
+ ad=1040 pd=334 as=0 ps=0 
M3549 n_1380 n_1380 Vdd GND dfet w=10 l=7
+ ad=1067 pd=354 as=0 ps=0 
M3550 n_1154 notRdy0 GND GND efet w=61 l=6
+ ad=1121 pd=344 as=0 ps=0 
M3551 n_1517 n_572 GND GND efet w=37 l=6
+ ad=1085 pd=292 as=0 ps=0 
M3552 Vdd n_1517 n_1517 GND dfet w=10 l=9
+ ad=0 pd=0 as=1033 ps=336 
M3553 Vdd n_1231 n_1231 GND dfet w=9 l=20
+ ad=0 pd=0 as=448 ps=110 
M3554 n_470 n_470 Vdd GND dfet w=10 l=10
+ ad=1641 pd=574 as=0 ps=0 
M3555 n_1448 n_1448 Vdd GND dfet w=10 l=12
+ ad=1011 pd=322 as=0 ps=0 
M3556 Vdd n_572 n_572 GND dfet w=10 l=13
+ ad=0 pd=0 as=2325 ps=752 
M3557 n_586 n_1619 GND GND efet w=43 l=6
+ ad=0 pd=0 as=0 ps=0 
M3558 Vdd n_442 n_442 GND dfet w=9 l=13
+ ad=0 pd=0 as=1665 ps=570 
M3559 GND n_182 n_442 GND efet w=50 l=6
+ ad=0 pd=0 as=1061 ps=334 
M3560 n_1347 cclk n_1527 GND efet w=12 l=9
+ ad=0 pd=0 as=151 ps=60 
M3561 n_1455 cclk n_1505 GND efet w=13 l=9
+ ad=0 pd=0 as=152 ps=74 
M3562 GND pipeUNK21 n_572 GND efet w=77 l=6
+ ad=0 pd=0 as=921 ps=220 
M3563 n_1231 n_1409 GND GND efet w=36 l=7
+ ad=873 pd=248 as=0 ps=0 
M3564 Vdd n_19 n_19 GND dfet w=10 l=16
+ ad=0 pd=0 as=361 ps=98 
M3565 Vdd n_1154 n_1154 GND dfet w=8 l=7
+ ad=0 pd=0 as=711 ps=236 
M3566 n_1718 cp1 n_671 GND efet w=12 l=8
+ ad=0 pd=0 as=136 ps=72 
M3567 n_812 n_812 Vdd GND dfet w=10 l=10
+ ad=755 pd=244 as=0 ps=0 
M3568 n_104 n_104 Vdd GND dfet w=10 l=11
+ ad=4812 pd=1628 as=0 ps=0 
M3569 n_1044 n_812 GND GND efet w=43 l=6
+ ad=1583 pd=420 as=0 ps=0 
M3570 Vdd n_1044 n_1044 GND dfet w=10 l=12
+ ad=0 pd=0 as=2740 ps=998 
M3571 n_1039 n_1039 Vdd GND dfet w=9 l=21
+ ad=453 pd=100 as=0 ps=0 
M3572 n_1161 cp1 n_109 GND efet w=14 l=9
+ ad=294 pd=92 as=0 ps=0 
M3573 Vdd n_253 n_253 GND dfet w=10 l=19
+ ad=0 pd=0 as=4197 ps=1372 
M3574 GND x_op_T0_bit n_1379 GND efet w=30 l=6
+ ad=0 pd=0 as=1443 ps=340 
M3575 Vdd n_646 n_646 GND dfet w=10 l=7
+ ad=0 pd=0 as=12020 ps=4204 
M3576 GND n_1161 n_732 GND efet w=78 l=6
+ ad=0 pd=0 as=1832 ps=458 
M3577 Vdd n_732 n_732 GND dfet w=11 l=10
+ ad=0 pd=0 as=1206 ps=364 
M3578 PD_xxxx10x0 PD_xxxx10x0 Vdd GND dfet w=10 l=9
+ ad=2138 pd=760 as=0 ps=0 
M3579 n_1515 PD_n_0xx0xx0x GND GND efet w=100 l=6
+ ad=0 pd=0 as=0 ps=0 
M3580 GND n_409 PD_xxx010x1 GND efet w=32 l=7
+ ad=0 pd=0 as=1658 ps=424 
M3581 PD_xxxx10x0 pd0_clearIR GND GND efet w=38 l=6
+ ad=1792 pd=434 as=0 ps=0 
M3582 GND PD_0xx0xx0x PD_n_0xx0xx0x GND efet w=65 l=7
+ ad=0 pd=0 as=976 ps=260 
M3583 PD_0xx0xx0x PD_0xx0xx0x Vdd GND dfet w=9 l=11
+ ad=1105 pd=354 as=0 ps=0 
M3584 PD_n_0xx0xx0x PD_n_0xx0xx0x Vdd GND dfet w=9 l=7
+ ad=1140 pd=398 as=0 ps=0 
M3585 PD_1xx000x0 PD_1xx000x0 Vdd GND dfet w=10 l=10
+ ad=1790 pd=646 as=0 ps=0 
M3586 GND pd1_clearIR PD_0xx0xx0x GND efet w=31 l=6
+ ad=0 pd=0 as=1605 ps=408 
M3587 PD_xxx010x1 pd4_clearIR GND GND efet w=48 l=6
+ ad=0 pd=0 as=0 ps=0 
M3588 GND n_1083 PD_xxx010x1 GND efet w=46 l=6
+ ad=0 pd=0 as=0 ps=0 
M3589 PD_1xx000x0 pd0_clearIR GND GND efet w=31 l=6
+ ad=2006 pd=504 as=0 ps=0 
M3590 GND PD_xxxx10x0 n_231 GND efet w=87 l=6
+ ad=0 pd=0 as=1413 ps=332 
M3591 Vdd n_231 n_231 GND dfet w=9 l=7
+ ad=0 pd=0 as=1060 ps=376 
M3592 n_106 nTWOCYCLE_phi1 n_732 GND efet w=150 l=6
+ ad=1007 pd=314 as=0 ps=0 
M3593 n_1528 cp1 n_1215 GND efet w=14 l=9
+ ad=207 pd=82 as=0 ps=0 
M3594 n_106 n_1528 GND GND efet w=150 l=6
+ ad=0 pd=0 as=0 ps=0 
M3595 GND pd7_clearIR PD_0xx0xx0x GND efet w=45 l=6
+ ad=0 pd=0 as=0 ps=0 
M3596 PD_1xx000x0 n_1605 GND GND efet w=33 l=6
+ ad=0 pd=0 as=0 ps=0 
M3597 ONEBYTE n_231 GND GND efet w=74 l=6
+ ad=783 pd=254 as=0 ps=0 
M3598 GND D1x1 n_380 GND efet w=56 l=6
+ ad=0 pd=0 as=336 ps=124 
M3599 n_1039 cp1 n_24 GND efet w=13 l=8
+ ad=0 pd=0 as=198 ps=78 
M3600 n_440 n_24 GND GND efet w=149 l=7
+ ad=0 pd=0 as=0 ps=0 
M3601 Vdd n_440 n_440 GND dfet w=11 l=9
+ ad=0 pd=0 as=7163 ps=2416 
M3602 GND n_31 n_1044 GND efet w=42 l=7
+ ad=0 pd=0 as=0 ps=0 
M3603 p2 cp1 n_845 GND efet w=12 l=8
+ ad=155 pd=58 as=1663 ps=480 
M3604 GND p2 n_334 GND efet w=77 l=8
+ ad=0 pd=0 as=0 ps=0 
M3605 Vdd n_334 n_334 GND dfet w=9 l=9
+ ad=0 pd=0 as=4511 ps=1544 
M3606 Vdd n_845 n_845 GND dfet w=10 l=19
+ ad=0 pd=0 as=854 ps=270 
M3607 Vdd n_553 n_553 GND dfet w=10 l=16
+ ad=0 pd=0 as=856 ps=262 
M3608 ONEBYTE ONEBYTE Vdd GND dfet w=10 l=7
+ ad=6889 pd=2364 as=0 ps=0 
M3609 n_380 fetch clearIR GND efet w=56 l=7
+ ad=0 pd=0 as=778 ps=190 
M3610 Vdd clearIR clearIR GND dfet w=10 l=12
+ ad=0 pd=0 as=3607 ps=1108 
M3611 PD_0xx0xx0x pd4_clearIR GND GND efet w=31 l=6
+ ad=0 pd=0 as=0 ps=0 
M3612 GND n_1083 PD_xxxx10x0 GND efet w=40 l=6
+ ad=0 pd=0 as=0 ps=0 
M3613 GND pd2_clearIR PD_xxx010x1 GND efet w=32 l=6
+ ad=0 pd=0 as=0 ps=0 
M3614 GND pd2_clearIR PD_xxxx10x0 GND efet w=39 l=6
+ ad=0 pd=0 as=0 ps=0 
M3615 PD_1xx000x0 pd3_clearIR GND GND efet w=41 l=7
+ ad=0 pd=0 as=0 ps=0 
M3616 PD_1xx000x0 pd4_clearIR GND GND efet w=32 l=6
+ ad=0 pd=0 as=0 ps=0 
M3617 GND pd2_clearIR PD_1xx000x0 GND efet w=32 l=6
+ ad=0 pd=0 as=0 ps=0 
M3618 GND pd3 pd3_clearIR GND efet w=84 l=6
+ ad=0 pd=0 as=1162 ps=306 
M3619 pd5_clearIR pd5 GND GND efet w=85 l=7
+ ad=1073 pd=284 as=0 ps=0 
M3620 GND pd0 pd0_clearIR GND efet w=84 l=7
+ ad=0 pd=0 as=1021 ps=300 
M3621 pd1_clearIR pd1 GND GND efet w=85 l=7
+ ad=1019 pd=298 as=0 ps=0 
M3622 n_1662 n_1124 GND GND efet w=49 l=7
+ ad=708 pd=198 as=0 ps=0 
M3623 GND clearIR pd4_clearIR GND efet w=32 l=6
+ ad=0 pd=0 as=983 ps=296 
M3624 GND notRdy0 fetch GND efet w=38 l=6
+ ad=0 pd=0 as=879 ps=200 
M3625 n_1662 n_1662 Vdd GND dfet w=9 l=23
+ ad=1631 pd=474 as=0 ps=0 
M3626 GND op_T__bit n_513 GND efet w=48 l=7
+ ad=0 pd=0 as=1233 ps=322 
M3627 n_1426 n_270 GND GND efet w=38 l=7
+ ad=645 pd=162 as=0 ps=0 
M3628 n_845 n_1662 n_1426 GND efet w=40 l=6
+ ad=0 pd=0 as=0 ps=0 
M3629 n_511 n_553 n_845 GND efet w=56 l=6
+ ad=512 pd=146 as=0 ps=0 
M3630 Vdd n_1055 n_1055 GND dfet w=10 l=13
+ ad=0 pd=0 as=4878 ps=1728 
M3631 n_1154 n_959 GND GND efet w=50 l=6
+ ad=0 pd=0 as=0 ps=0 
M3632 n_19 n_770 GND GND efet w=35 l=7
+ ad=786 pd=182 as=0 ps=0 
M3633 GND n_1708 n_19 GND efet w=40 l=6
+ ad=0 pd=0 as=0 ps=0 
M3634 GND n_853 n_1517 GND efet w=46 l=6
+ ad=0 pd=0 as=0 ps=0 
M3635 n_1055 n_771 GND GND efet w=26 l=7
+ ad=0 pd=0 as=0 ps=0 
M3636 n_19 cclk pipeUNK18 GND efet w=12 l=9
+ ad=0 pd=0 as=175 ps=70 
M3637 n_1231 cclk pipeUNK21 GND efet w=11 l=8
+ ad=0 pd=0 as=411 ps=126 
M3638 n_14 n_671 GND GND efet w=37 l=7
+ ad=0 pd=0 as=0 ps=0 
M3639 n_1550 n_781 GND GND efet w=40 l=7
+ ad=340 pd=112 as=0 ps=0 
M3640 n_845 n_1573 n_1550 GND efet w=50 l=6
+ ad=0 pd=0 as=0 ps=0 
M3641 GND pipeUNK17 n_511 GND efet w=64 l=7
+ ad=0 pd=0 as=0 ps=0 
M3642 n_14 n_323 GND GND efet w=47 l=6
+ ad=0 pd=0 as=0 ps=0 
M3643 n_959 short_circuit_branch_add GND GND efet w=160 l=7
+ ad=1738 pd=490 as=0 ps=0 
M3644 n_323 cp1 n_959 GND efet w=12 l=8
+ ad=156 pd=68 as=0 ps=0 
M3645 GND pipeUNK18 n_850 GND efet w=77 l=6
+ ad=0 pd=0 as=774 ps=198 
M3646 Vdd n_1619 n_1619 GND dfet w=10 l=17
+ ad=0 pd=0 as=974 ps=314 
M3647 n_1619 n_1448 GND GND efet w=30 l=7
+ ad=1199 pd=344 as=0 ps=0 
M3648 n_1619 n_182 GND GND efet w=30 l=7
+ ad=0 pd=0 as=0 ps=0 
M3649 n_465 n_465 Vdd GND dfet w=9 l=7
+ ad=235 pd=90 as=0 ps=0 
M3650 Vdd n_1446 n_1446 GND dfet w=10 l=13
+ ad=0 pd=0 as=541 ps=162 
M3651 n_850 n_850 Vdd GND dfet w=10 l=16
+ ad=1382 pd=404 as=0 ps=0 
M3652 GND pipeUNK20 n_959 GND efet w=163 l=6
+ ad=0 pd=0 as=0 ps=0 
M3653 n_14 cclk pipeUNK20 GND efet w=12 l=8
+ ad=0 pd=0 as=203 ps=78 
M3654 pipeBRtaken cclk n_586 GND efet w=14 l=7
+ ad=353 pd=96 as=0 ps=0 
M3655 Vdd n_959 n_959 GND dfet w=8 l=8
+ ad=0 pd=0 as=659 ps=226 
M3656 GND n_206 n_465 GND efet w=75 l=6
+ ad=0 pd=0 as=1149 ps=302 
M3657 n_1446 n_771 GND GND efet w=53 l=6
+ ad=941 pd=268 as=0 ps=0 
M3658 GND n_850 n_1446 GND efet w=45 l=7
+ ad=0 pd=0 as=0 ps=0 
M3659 short_circuit_branch_add cp1 n_1570 GND efet w=13 l=8
+ ad=1990 pd=526 as=170 ps=70 
M3660 short_circuit_branch_add n_771 n_465 GND efet w=18 l=8
+ ad=0 pd=0 as=0 ps=0 
M3661 n_206 n_1446 short_circuit_branch_add GND efet w=18 l=7
+ ad=1879 pd=466 as=0 ps=0 
M3662 short_circuit_branch_add n_850 GND GND efet w=76 l=6
+ ad=0 pd=0 as=0 ps=0 
M3663 n_1472 cp1 D1x1 GND efet w=14 l=7
+ ad=284 pd=108 as=0 ps=0 
M3664 n_1275 pipeBRtaken GND GND efet w=97 l=6
+ ad=1633 pd=410 as=0 ps=0 
M3665 Vdd n_1275 n_1275 GND dfet w=10 l=11
+ ad=0 pd=0 as=266 ps=88 
M3666 Vdd dpc36_nIPC dpc36_nIPC GND dfet w=10 l=13
+ ad=0 pd=0 as=2720 ps=832 
M3667 n_1480 n_1472 GND GND efet w=161 l=6
+ ad=3122 pd=672 as=0 ps=0 
M3668 dpc36_nIPC n_1570 n_1480 GND efet w=157 l=5
+ ad=1910 pd=486 as=0 ps=0 
M3669 GND notRdy0 n_1275 GND efet w=49 l=6
+ ad=0 pd=0 as=0 ps=0 
M3670 n_1705 n_1705 Vdd GND dfet w=10 l=11
+ ad=2616 pd=834 as=0 ps=0 
M3671 GND ONEBYTE n_1275 GND efet w=45 l=6
+ ad=0 pd=0 as=0 ps=0 
M3672 n_1275 cp1 n_1581 GND efet w=13 l=7
+ ad=0 pd=0 as=154 ps=72 
M3673 n_506 cclk n_1602 GND efet w=12 l=8
+ ad=0 pd=0 as=160 ps=78 
M3674 n_1683 cclk n_1090 GND efet w=12 l=8
+ ad=167 pd=60 as=0 ps=0 
M3675 n_11 cclk n_55 GND efet w=12 l=9
+ ad=0 pd=0 as=160 ps=74 
M3676 n_1037 cclk n_266 GND efet w=11 l=9
+ ad=0 pd=0 as=148 ps=62 
M3677 n_272 cclk n_1162 GND efet w=13 l=9
+ ad=0 pd=0 as=149 ps=74 
M3678 n_952 cclk n_1509 GND efet w=12 l=8
+ ad=0 pd=0 as=149 ps=76 
M3679 n_824 cclk n_398 GND efet w=12 l=8
+ ad=0 pd=0 as=179 ps=62 
M3680 Vdd n_1295 n_1295 GND dfet w=9 l=10
+ ad=0 pd=0 as=1322 ps=394 
M3681 GND n_1527 n_1295 GND efet w=72 l=7
+ ad=0 pd=0 as=807 ps=210 
M3682 n_830 n_1505 GND GND efet w=52 l=7
+ ad=877 pd=224 as=0 ps=0 
M3683 Vdd n_830 n_830 GND dfet w=9 l=15
+ ad=0 pd=0 as=1257 ps=336 
M3684 Vdd n_1596 n_1596 GND dfet w=9 l=11
+ ad=0 pd=0 as=1269 ps=398 
M3685 GND n_1602 n_1596 GND efet w=72 l=6
+ ad=0 pd=0 as=829 ps=204 
M3686 GND n_43 n_830 GND efet w=26 l=6
+ ad=0 pd=0 as=0 ps=0 
M3687 Vdd n_966 n_966 GND dfet w=8 l=10
+ ad=0 pd=0 as=1190 ps=390 
M3688 GND n_1683 n_966 GND efet w=72 l=6
+ ad=0 pd=0 as=832 ps=208 
M3689 n_1238 n_1295 GND GND efet w=24 l=7
+ ad=335 pd=106 as=0 ps=0 
M3690 n_1047 n_830 GND GND efet w=23 l=8
+ ad=334 pd=100 as=0 ps=0 
M3691 n_628 n_55 GND GND efet w=59 l=5
+ ad=861 pd=222 as=0 ps=0 
M3692 Vdd n_628 n_628 GND dfet w=10 l=13
+ ad=0 pd=0 as=946 ps=322 
M3693 n_1238 n_1238 Vdd GND dfet w=9 l=14
+ ad=1331 pd=356 as=0 ps=0 
M3694 n_1271 n_1596 GND GND efet w=25 l=7
+ ad=369 pd=104 as=0 ps=0 
M3695 n_462 cclk n_878 GND efet w=13 l=9
+ ad=0 pd=0 as=169 ps=62 
M3696 n_598 cclk n_176 GND efet w=12 l=9
+ ad=152 pd=60 as=0 ps=0 
M3697 n_442 cclk n_509 GND efet w=12 l=9
+ ad=0 pd=0 as=144 ps=74 
M3698 n_1211 cclk n_897 GND efet w=12 l=10
+ ad=0 pd=0 as=150 ps=58 
M3699 n_182 cclk n_265 GND efet w=12 l=10
+ ad=0 pd=0 as=155 ps=72 
M3700 Vdd n_525 n_525 GND dfet w=10 l=12
+ ad=0 pd=0 as=1038 ps=322 
M3701 GND n_266 n_525 GND efet w=57 l=5
+ ad=0 pd=0 as=946 ps=226 
M3702 n_21 n_1162 GND GND efet w=54 l=6
+ ad=872 pd=222 as=0 ps=0 
M3703 Vdd n_21 n_21 GND dfet w=9 l=13
+ ad=0 pd=0 as=1259 ps=340 
M3704 GND cclk n_628 GND efet w=25 l=5
+ ad=0 pd=0 as=0 ps=0 
M3705 n_525 cclk GND GND efet w=25 l=6
+ ad=0 pd=0 as=0 ps=0 
M3706 n_611 n_1509 GND GND efet w=54 l=6
+ ad=834 pd=226 as=0 ps=0 
M3707 Vdd n_611 n_611 GND dfet w=9 l=14
+ ad=0 pd=0 as=1270 ps=338 
M3708 n_1047 n_1047 Vdd GND dfet w=10 l=15
+ ad=1218 pd=360 as=0 ps=0 
M3709 n_1635 n_966 GND GND efet w=24 l=6
+ ad=337 pd=104 as=0 ps=0 
M3710 Vdd n_1295 dpc25_SBDB GND dfet w=11 l=10
+ ad=0 pd=0 as=1353 ps=316 
M3711 GND n_1238 dpc25_SBDB GND efet w=94 l=8
+ ad=0 pd=0 as=0 ps=0 
M3712 Vdd n_830 dpc23_SBAC GND dfet w=10 l=10
+ ad=0 pd=0 as=1997 ps=402 
M3713 n_1271 n_1271 Vdd GND dfet w=9 l=15
+ ad=1249 pd=358 as=0 ps=0 
M3714 n_1335 n_628 GND GND efet w=25 l=5
+ ad=367 pd=108 as=0 ps=0 
M3715 GND n_43 n_21 GND efet w=25 l=7
+ ad=0 pd=0 as=0 ps=0 
M3716 Vdd n_321 n_321 GND dfet w=10 l=10
+ ad=0 pd=0 as=1199 ps=392 
M3717 GND n_398 n_321 GND efet w=73 l=7
+ ad=0 pd=0 as=793 ps=216 
M3718 n_1635 n_1635 Vdd GND dfet w=9 l=14
+ ad=1229 pd=360 as=0 ps=0 
M3719 Vdd n_1596 dpc27_SBADH GND dfet w=9 l=9
+ ad=0 pd=0 as=1290 ps=282 
M3720 dpc23_SBAC n_1247 GND GND efet w=76 l=6
+ ad=0 pd=0 as=0 ps=0 
M3721 GND n_1047 dpc23_SBAC GND efet w=77 l=7
+ ad=0 pd=0 as=0 ps=0 
M3722 GND n_1271 dpc27_SBADH GND efet w=96 l=7
+ ad=0 pd=0 as=0 ps=0 
M3723 Vdd n_966 dpc29_0ADH17 GND dfet w=10 l=9
+ ad=0 pd=0 as=1217 ps=262 
M3724 n_1335 n_1335 Vdd GND dfet w=9 l=12
+ ad=1063 pd=356 as=0 ps=0 
M3725 GND n_1635 dpc29_0ADH17 GND efet w=96 l=6
+ ad=0 pd=0 as=0 ps=0 
M3726 Vdd n_628 dpc24_ACSB GND dfet w=10 l=8
+ ad=0 pd=0 as=1779 ps=384 
M3727 GND n_525 n_800 GND efet w=26 l=6
+ ad=0 pd=0 as=390 ps=108 
M3728 n_228 n_21 GND GND efet w=26 l=8
+ ad=336 pd=106 as=0 ps=0 
M3729 GND n_43 n_611 GND efet w=24 l=6
+ ad=0 pd=0 as=0 ps=0 
M3730 Vdd n_631 n_631 GND dfet w=9 l=10
+ ad=0 pd=0 as=1231 ps=396 
M3731 GND n_878 n_631 GND efet w=73 l=7
+ ad=0 pd=0 as=824 ps=214 
M3732 n_800 n_800 Vdd GND dfet w=10 l=12
+ ad=1099 pd=362 as=0 ps=0 
M3733 Vdd n_525 dpc26_ACDB GND dfet w=9 l=9
+ ad=0 pd=0 as=1902 ps=428 
M3734 n_255 n_611 GND GND efet w=24 l=8
+ ad=316 pd=102 as=0 ps=0 
M3735 Vdd n_1260 n_1260 GND dfet w=9 l=10
+ ad=0 pd=0 as=1200 ps=398 
M3736 GND n_598 n_1260 GND efet w=73 l=7
+ ad=0 pd=0 as=760 ps=210 
M3737 n_1270 n_509 GND GND efet w=53 l=5
+ ad=925 pd=222 as=0 ps=0 
M3738 Vdd n_1270 n_1270 GND dfet w=10 l=15
+ ad=0 pd=0 as=1151 ps=336 
M3739 Vdd n_1369 n_1369 GND dfet w=9 l=10
+ ad=0 pd=0 as=1276 ps=400 
M3740 GND n_897 n_1369 GND efet w=74 l=7
+ ad=0 pd=0 as=806 ps=216 
M3741 GND n_43 n_1270 GND efet w=27 l=8
+ ad=0 pd=0 as=0 ps=0 
M3742 n_228 n_228 Vdd GND dfet w=10 l=15
+ ad=1297 pd=358 as=0 ps=0 
M3743 Vdd n_21 dpc30_ADHPCH GND dfet w=10 l=11
+ ad=0 pd=0 as=1887 ps=446 
M3744 DA_C01 DA_C01 Vdd GND dfet w=10 l=16
+ ad=1643 pd=502 as=0 ps=0 
M3745 naluresult0 dpc17_SUMS n_AxBxC_0 GND efet w=10 l=7
+ ad=0 pd=0 as=0 ps=0 
M3746 n_AxBxC_0 _AxB_0_nC0in GND GND efet w=24 l=6
+ ad=0 pd=0 as=0 ps=0 
M3747 _AxB_0_nC0in n_AxB_0 GND GND efet w=18 l=7
+ ad=654 pd=222 as=0 ps=0 
M3748 n_AxB_0 n_AxB_0 Vdd GND dfet w=9 l=17
+ ad=1298 pd=384 as=0 ps=0 
M3749 GND n_105 _AxB_0_nC0in GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M3750 C01 C01 Vdd GND dfet w=10 l=10
+ ad=1119 pd=384 as=0 ps=0 
M3751 Vdd n_936 n_936 GND dfet w=9 l=17
+ ad=0 pd=0 as=2425 ps=804 
M3752 Vdd A_B1 A_B1 GND dfet w=9 l=16
+ ad=0 pd=0 as=865 ps=252 
M3753 Vdd _AxB_0_nC0in _AxB_0_nC0in GND dfet w=10 l=16
+ ad=0 pd=0 as=954 ps=294 
M3754 Vdd nC01 nC01 GND dfet w=9 l=16
+ ad=0 pd=0 as=1133 ps=336 
M3755 n_936 nA_B1 GND GND efet w=18 l=6
+ ad=703 pd=188 as=0 ps=0 
M3756 nC01 C01 GND GND efet w=18 l=6
+ ad=284 pd=96 as=0 ps=0 
M3757 DA_C01 n_A_B_0 GND GND efet w=25 l=6
+ ad=861 pd=214 as=0 ps=0 
M3758 n_1707 n_936 GND GND efet w=54 l=6
+ ad=324 pd=120 as=0 ps=0 
M3759 n_319 DA_C01 n_1707 GND efet w=54 l=6
+ ad=666 pd=192 as=0 ps=0 
M3760 n_1354 nA_B0 DA_C01 GND efet w=53 l=6
+ ad=265 pd=116 as=0 ps=0 
M3761 GND notalucin n_1354 GND efet w=53 l=7
+ ad=0 pd=0 as=0 ps=0 
M3762 GND n_A_B_1 A_B1 GND efet w=24 l=7
+ ad=0 pd=0 as=574 ps=170 
M3763 n_1510 A_B1 GND GND efet w=54 l=6
+ ad=316 pd=120 as=0 ps=0 
M3764 nC12 C01 n_1510 GND efet w=54 l=6
+ ad=820 pd=230 as=0 ps=0 
M3765 n_AxB_1 dpc16_EORS naluresult1 GND efet w=11 l=8
+ ad=455 pd=136 as=0 ps=0 
M3766 GND AxB1 n_AxB_1 GND efet w=29 l=6
+ ad=0 pd=0 as=0 ps=0 
M3767 AxB1 n_936 GND GND efet w=18 l=6
+ ad=552 pd=164 as=0 ps=0 
M3768 GND n_A_B_1 AxB1 GND efet w=18 l=7
+ ad=0 pd=0 as=0 ps=0 
M3769 GND n_936 nC12 GND efet w=26 l=6
+ ad=0 pd=0 as=0 ps=0 
M3770 n_1388 AxB1 GND GND efet w=35 l=6
+ ad=210 pd=82 as=0 ps=0 
M3771 n_AxBxC_1 nC01 n_1388 GND efet w=35 l=6
+ ad=845 pd=216 as=0 ps=0 
M3772 Vdd n_AxBxC_1 n_AxBxC_1 GND dfet w=10 l=17
+ ad=0 pd=0 as=472 ps=106 
M3773 n_319 n_319 Vdd GND dfet w=9 l=16
+ ad=3363 pd=1088 as=0 ps=0 
M3774 n_388 n_388 Vdd GND dfet w=10 l=13
+ ad=3118 pd=1108 as=0 ps=0 
M3775 n_388 DA_C01 GND GND efet w=33 l=6
+ ad=1493 pd=378 as=0 ps=0 
M3776 n_388 DA_AxB2 GND GND efet w=34 l=6
+ ad=0 pd=0 as=0 ps=0 
M3777 n_AxBxC_1 n_AxB1__C01 GND GND efet w=27 l=6
+ ad=0 pd=0 as=0 ps=0 
M3778 naluresult1 dpc17_SUMS n_AxBxC_1 GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M3779 n_388 n_936 GND GND efet w=27 l=6
+ ad=0 pd=0 as=0 ps=0 
M3780 GND AxB1 n_388 GND efet w=30 l=6
+ ad=0 pd=0 as=0 ps=0 
M3781 n_AxB1__C01 AxB1 GND GND efet w=18 l=6
+ ad=523 pd=166 as=0 ps=0 
M3782 n_AxB_1 n_AxB_1 Vdd GND dfet w=9 l=16
+ ad=427 pd=120 as=0 ps=0 
M3783 AxB1 AxB1 Vdd GND dfet w=9 l=16
+ ad=2426 pd=804 as=0 ps=0 
M3784 GND nC01 n_AxB1__C01 GND efet w=35 l=7
+ ad=0 pd=0 as=0 ps=0 
M3785 Vdd nC12 nC12 GND dfet w=9 l=9
+ ad=0 pd=0 as=1458 ps=460 
M3786 n_AxB1__C01 n_AxB1__C01 Vdd GND dfet w=10 l=17
+ ad=771 pd=228 as=0 ps=0 
M3787 A_B2 A_B2 Vdd GND dfet w=9 l=16
+ ad=889 pd=266 as=0 ps=0 
M3788 Vdd C12 C12 GND dfet w=9 l=16
+ ad=0 pd=0 as=1053 ps=344 
M3789 nA_B2 dpc14_SRS naluresult1 GND efet w=11 l=7
+ ad=0 pd=0 as=0 ps=0 
M3790 naluresult2 dpc13_ORS n_A_B_2 GND efet w=12 l=7
+ ad=1656 pd=438 as=1013 ps=278 
M3791 GND dpc12_0ADD alua2 GND efet w=12 l=6
+ ad=0 pd=0 as=573 ps=142 
M3792 alua2 dpc11_SBADD sb2 GND efet w=12 l=7
+ ad=0 pd=0 as=0 ps=0 
M3793 n_A_B_2 alua2 GND GND efet w=31 l=7
+ ad=0 pd=0 as=0 ps=0 
M3794 GND alub2 n_A_B_2 GND efet w=32 l=6
+ ad=0 pd=0 as=0 ps=0 
M3795 Vdd n_A_B_2 n_A_B_2 GND dfet w=9 l=21
+ ad=0 pd=0 as=3438 ps=1062 
M3796 adl3 dpc10_ADLADD alub3 GND efet w=11 l=7
+ ad=0 pd=0 as=575 ps=144 
M3797 alub3 dpc8_nDBADD n_1621 GND efet w=11 l=8
+ ad=0 pd=0 as=924 ps=278 
M3798 alub3 dpc9_DBADD idb3 GND efet w=12 l=6
+ ad=0 pd=0 as=2106 ps=550 
M3799 GND idb3 n_1621 GND efet w=62 l=7
+ ad=0 pd=0 as=0 ps=0 
M3800 n_1621 n_1621 Vdd GND dfet w=9 l=17
+ ad=343 pd=86 as=0 ps=0 
M3801 n_313 alua3 GND GND efet w=61 l=6
+ ad=366 pd=134 as=0 ps=0 
M3802 nA_B3 alub3 n_313 GND efet w=61 l=6
+ ad=1193 pd=306 as=0 ps=0 
M3803 Vdd nA_B3 nA_B3 GND dfet w=10 l=21
+ ad=0 pd=0 as=986 ps=248 
M3804 C12 nC12 GND GND efet w=17 l=6
+ ad=270 pd=96 as=0 ps=0 
M3805 A_B2 n_A_B_2 GND GND efet w=18 l=8
+ ad=306 pd=88 as=0 ps=0 
M3806 n_716 A_B2 n_AxB_2 GND efet w=36 l=6
+ ad=197 pd=84 as=807 ps=236 
M3807 naluresult2 dpc15_ANDS nA_B2 GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M3808 n_AxB_2 dpc16_EORS naluresult2 GND efet w=12 l=7
+ ad=0 pd=0 as=0 ps=0 
M3809 GND nA_B2 n_716 GND efet w=34 l=6
+ ad=0 pd=0 as=0 ps=0 
M3810 C23 n_A_B_2 GND GND efet w=28 l=6
+ ad=997 pd=262 as=0 ps=0 
M3811 n_433 nA_B2 C23 GND efet w=55 l=6
+ ad=500 pd=162 as=0 ps=0 
M3812 GND nC12 n_433 GND efet w=72 l=6
+ ad=0 pd=0 as=0 ps=0 
M3813 n_1572 n_AxB_2 GND GND efet w=36 l=7
+ ad=216 pd=84 as=0 ps=0 
M3814 n_AxBxC_2 C12 n_1572 GND efet w=36 l=5
+ ad=966 pd=238 as=0 ps=0 
M3815 Vdd n_AxBxC_2 n_AxBxC_2 GND dfet w=9 l=17
+ ad=0 pd=0 as=452 ps=104 
M3816 DA_AxB2 DA_AB2 GND GND efet w=33 l=5
+ ad=1284 pd=314 as=0 ps=0 
M3817 n_1610 AxB3 GND GND efet w=41 l=7
+ ad=604 pd=184 as=0 ps=0 
M3818 GND DA_AB2 n_1610 GND efet w=27 l=6
+ ad=0 pd=0 as=0 ps=0 
M3819 n_1610 n_1610 Vdd GND dfet w=10 l=16
+ ad=2349 pd=730 as=0 ps=0 
M3820 naluresult2 dpc17_SUMS n_AxBxC_2 GND efet w=11 l=7
+ ad=0 pd=0 as=0 ps=0 
M3821 n_AxBxC_2 _AxB_2_nC12 GND GND efet w=27 l=6
+ ad=0 pd=0 as=0 ps=0 
M3822 _AxB_2_nC12 n_AxB_2 GND GND efet w=18 l=5
+ ad=646 pd=210 as=0 ps=0 
M3823 nA_B3 dpc14_SRS naluresult2 GND efet w=11 l=7
+ ad=0 pd=0 as=0 ps=0 
M3824 naluresult3 dpc13_ORS n_A_B_3 GND efet w=13 l=7
+ ad=1864 pd=500 as=1054 ps=282 
M3825 GND dpc12_0ADD alua3 GND efet w=13 l=7
+ ad=0 pd=0 as=552 ps=144 
M3826 alua3 dpc11_SBADD sb3 GND efet w=12 l=7
+ ad=0 pd=0 as=0 ps=0 
M3827 adl4 dpc10_ADLADD alub4 GND efet w=11 l=6
+ ad=0 pd=0 as=565 ps=144 
M3828 alub4 dpc8_nDBADD n_478 GND efet w=12 l=9
+ ad=0 pd=0 as=921 ps=276 
M3829 alub4 dpc9_DBADD idb4 GND efet w=12 l=8
+ ad=0 pd=0 as=2179 ps=562 
M3830 GND idb4 n_478 GND efet w=62 l=7
+ ad=0 pd=0 as=0 ps=0 
M3831 n_478 n_478 Vdd GND dfet w=9 l=17
+ ad=332 pd=86 as=0 ps=0 
M3832 n_A_B_3 alua3 GND GND efet w=32 l=6
+ ad=0 pd=0 as=0 ps=0 
M3833 GND alub3 n_A_B_3 GND efet w=31 l=7
+ ad=0 pd=0 as=0 ps=0 
M3834 Vdd n_A_B_3 n_A_B_3 GND dfet w=10 l=22
+ ad=0 pd=0 as=1370 ps=416 
M3835 n_185 alua4 GND GND efet w=61 l=6
+ ad=366 pd=134 as=0 ps=0 
M3836 nA_B4 alub4 n_185 GND efet w=61 l=7
+ ad=1110 pd=296 as=0 ps=0 
M3837 Vdd nA_B4 nA_B4 GND dfet w=9 l=21
+ ad=0 pd=0 as=1613 ps=434 
M3838 naluresult3 dpc15_ANDS nA_B3 GND efet w=12 l=7
+ ad=0 pd=0 as=0 ps=0 
M3839 n_AxB_2 n_AxB_2 Vdd GND dfet w=9 l=16
+ ad=1197 pd=382 as=0 ps=0 
M3840 GND C12 _AxB_2_nC12 GND efet w=26 l=7
+ ad=0 pd=0 as=0 ps=0 
M3841 DA_AB2 nA_B2 GND GND efet w=27 l=6
+ ad=969 pd=304 as=0 ps=0 
M3842 C23 C23 Vdd GND dfet w=10 l=9
+ ad=1120 pd=382 as=0 ps=0 
M3843 Vdd n_988 n_988 GND dfet w=10 l=17
+ ad=0 pd=0 as=940 ps=304 
M3844 Vdd A_B3 A_B3 GND dfet w=10 l=17
+ ad=0 pd=0 as=824 ps=250 
M3845 n_988 nA_B3 GND GND efet w=17 l=7
+ ad=722 pd=196 as=0 ps=0 
M3846 Vdd _AxB_2_nC12 _AxB_2_nC12 GND dfet w=8 l=17
+ ad=0 pd=0 as=964 ps=292 
M3847 Vdd nC23 nC23 GND dfet w=10 l=16
+ ad=0 pd=0 as=1142 ps=340 
M3848 DA_AB2 DA_AB2 Vdd GND dfet w=9 l=16
+ ad=1719 pd=590 as=0 ps=0 
M3849 DA_AxB2 DA_AxB2 Vdd GND dfet w=10 l=17
+ ad=859 pd=268 as=0 ps=0 
M3850 DA_AxB2 n_A_B_2 GND GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M3851 nC23 C23 GND GND efet w=18 l=6
+ ad=340 pd=94 as=0 ps=0 
M3852 n_AxB_3 dpc16_EORS naluresult3 GND efet w=12 l=7
+ ad=475 pd=140 as=0 ps=0 
M3853 GND AxB3 n_AxB_3 GND efet w=29 l=6
+ ad=0 pd=0 as=0 ps=0 
M3854 GND n_A_B_3 A_B3 GND efet w=24 l=7
+ ad=0 pd=0 as=593 ps=196 
M3855 AxB3 n_988 GND GND efet w=18 l=6
+ ad=592 pd=184 as=0 ps=0 
M3856 GND n_A_B_3 AxB3 GND efet w=18 l=7
+ ad=0 pd=0 as=0 ps=0 
M3857 n_924 A_B3 GND GND efet w=53 l=6
+ ad=318 pd=118 as=0 ps=0 
M3858 nC34 C23 n_924 GND efet w=53 l=6
+ ad=1030 pd=268 as=0 ps=0 
M3859 GND n_988 nC34 GND efet w=26 l=6
+ ad=0 pd=0 as=0 ps=0 
M3860 n_136 AxB3 GND GND efet w=35 l=6
+ ad=210 pd=82 as=0 ps=0 
M3861 n_AxBxC_3 nC23 n_136 GND efet w=35 l=6
+ ad=828 pd=210 as=0 ps=0 
M3862 Vdd n_AxBxC_3 n_AxBxC_3 GND dfet w=10 l=17
+ ad=0 pd=0 as=482 ps=106 
M3863 n_AxBxC_3 n_AxB3__C23 GND GND efet w=26 l=6
+ ad=0 pd=0 as=0 ps=0 
M3864 naluresult3 dpc17_SUMS n_AxBxC_3 GND efet w=11 l=8
+ ad=0 pd=0 as=0 ps=0 
M3865 GND DC34 nC34 GND efet w=27 l=6
+ ad=0 pd=0 as=0 ps=0 
M3866 n_AxB3__C23 AxB3 GND GND efet w=18 l=6
+ ad=550 pd=168 as=0 ps=0 
M3867 GND nC23 n_AxB3__C23 GND efet w=34 l=6
+ ad=0 pd=0 as=0 ps=0 
M3868 n_AxB_3 n_AxB_3 Vdd GND dfet w=8 l=17
+ ad=445 pd=122 as=0 ps=0 
M3869 AxB3 AxB3 Vdd GND dfet w=9 l=16
+ ad=3793 pd=1274 as=0 ps=0 
M3870 nC34 nC34 Vdd GND dfet w=9 l=10
+ ad=1355 pd=442 as=0 ps=0 
M3871 A_B4 A_B4 Vdd GND dfet w=10 l=15
+ ad=791 pd=246 as=0 ps=0 
M3872 nA_B4 dpc14_SRS naluresult3 GND efet w=11 l=8
+ ad=0 pd=0 as=0 ps=0 
M3873 naluresult4 dpc13_ORS n_A_B_4 GND efet w=12 l=7
+ ad=1635 pd=448 as=988 ps=276 
M3874 GND dpc12_0ADD alua4 GND efet w=12 l=7
+ ad=0 pd=0 as=489 ps=134 
M3875 alua4 dpc11_SBADD sb4 GND efet w=11 l=8
+ ad=0 pd=0 as=0 ps=0 
M3876 adl5 dpc10_ADLADD alub5 GND efet w=10 l=8
+ ad=0 pd=0 as=568 ps=144 
M3877 alub5 dpc8_nDBADD n_1383 GND efet w=12 l=7
+ ad=0 pd=0 as=969 ps=276 
M3878 alub5 dpc9_DBADD idb5 GND efet w=12 l=8
+ ad=0 pd=0 as=1738 ps=448 
M3879 GND idb5 n_1383 GND efet w=61 l=7
+ ad=0 pd=0 as=0 ps=0 
M3880 n_1383 n_1383 Vdd GND dfet w=8 l=17
+ ad=332 pd=86 as=0 ps=0 
M3881 n_A_B_4 alua4 GND GND efet w=31 l=6
+ ad=0 pd=0 as=0 ps=0 
M3882 GND alub4 n_A_B_4 GND efet w=32 l=6
+ ad=0 pd=0 as=0 ps=0 
M3883 Vdd n_A_B_4 n_A_B_4 GND dfet w=10 l=22
+ ad=0 pd=0 as=1646 ps=524 
M3884 A_B4 n_A_B_4 GND GND efet w=18 l=6
+ ad=558 pd=158 as=0 ps=0 
M3885 n_AxB3__C23 n_AxB3__C23 Vdd GND dfet w=9 l=17
+ ad=764 pd=230 as=0 ps=0 
M3886 n_972 n_A_B_2 GND GND efet w=56 l=7
+ ad=1691 pd=430 as=0 ps=0 
M3887 GND n_319 n_972 GND efet w=67 l=6
+ ad=0 pd=0 as=0 ps=0 
M3888 adl0 dpc21_ADDADL alu0 GND efet w=16 l=8
+ ad=0 pd=0 as=1615 ps=422 
M3889 naluresult0 cclk notalu0 GND efet w=11 l=8
+ ad=0 pd=0 as=184 ps=76 
M3890 GND notalu0 alu0 GND efet w=100 l=6
+ ad=0 pd=0 as=0 ps=0 
M3891 alu0 dpc20_ADDSB06 sb0 GND efet w=21 l=8
+ ad=0 pd=0 as=0 ps=0 
M3892 alu0 alu0 Vdd GND dfet w=10 l=13
+ ad=355 pd=104 as=0 ps=0 
M3893 adl1 dpc21_ADDADL alu1 GND efet w=16 l=8
+ ad=0 pd=0 as=1537 ps=422 
M3894 naluresult1 cclk notalu1 GND efet w=11 l=9
+ ad=0 pd=0 as=164 ps=72 
M3895 GND notalu1 alu1 GND efet w=102 l=7
+ ad=0 pd=0 as=0 ps=0 
M3896 alu1 dpc20_ADDSB06 sb1 GND efet w=21 l=8
+ ad=0 pd=0 as=0 ps=0 
M3897 n_700 dpc18_nDAA GND GND efet w=27 l=6
+ ad=850 pd=254 as=0 ps=0 
M3898 n_972 n_1610 DC34 GND efet w=59 l=7
+ ad=0 pd=0 as=1126 ps=348 
M3899 n_972 n_388 DC34 GND efet w=59 l=6
+ ad=0 pd=0 as=0 ps=0 
M3900 n_700 n_700 Vdd GND dfet w=9 l=15
+ ad=1667 pd=526 as=0 ps=0 
M3901 n_700 cclk n_1565 GND efet w=12 l=8
+ ad=0 pd=0 as=140 ps=68 
M3902 GND dpc18_nDAA DC34 GND efet w=34 l=6
+ ad=0 pd=0 as=0 ps=0 
M3903 Vdd C34 C34 GND dfet w=10 l=15
+ ad=0 pd=0 as=2619 ps=840 
M3904 DC34 DC34 Vdd GND dfet w=10 l=10
+ ad=1083 pd=356 as=0 ps=0 
M3905 n_1218 n_1565 GND GND efet w=26 l=7
+ ad=730 pd=206 as=0 ps=0 
M3906 GND n_1565 n_1218 GND efet w=23 l=6
+ ad=0 pd=0 as=0 ps=0 
M3907 C34 nC34 GND GND efet w=18 l=7
+ ad=332 pd=120 as=0 ps=0 
M3908 naluresult4 dpc15_ANDS nA_B4 GND efet w=11 l=7
+ ad=0 pd=0 as=0 ps=0 
M3909 n_AxB_4 dpc16_EORS naluresult4 GND efet w=11 l=7
+ ad=874 pd=256 as=0 ps=0 
M3910 n_1559 alua5 GND GND efet w=61 l=7
+ ad=305 pd=132 as=0 ps=0 
M3911 nA_B5 alub5 n_1559 GND efet w=61 l=6
+ ad=1170 pd=300 as=0 ps=0 
M3912 Vdd nA_B5 nA_B5 GND dfet w=9 l=21
+ ad=0 pd=0 as=969 ps=244 
M3913 nA_B5 dpc14_SRS naluresult4 GND efet w=11 l=7
+ ad=0 pd=0 as=0 ps=0 
M3914 naluresult5 dpc13_ORS n_A_B_5 GND efet w=12 l=8
+ ad=1862 pd=504 as=927 ps=274 
M3915 GND dpc12_0ADD alua5 GND efet w=12 l=7
+ ad=0 pd=0 as=519 ps=138 
M3916 alua5 dpc11_SBADD sb5 GND efet w=11 l=8
+ ad=0 pd=0 as=0 ps=0 
M3917 n_618 dpc7_SS s6 GND efet w=12 l=8
+ ad=0 pd=0 as=312 ps=74 
M3918 s6 dpc6_SBS sb6 GND efet w=12 l=7
+ ad=0 pd=0 as=0 ps=0 
M3919 sb6 cclk Vdd GND efet w=22 l=6
+ ad=0 pd=0 as=0 ps=0 
M3920 Vdd n_721 n_721 GND dfet w=10 l=17
+ ad=0 pd=0 as=355 ps=100 
M3921 n_721 dpc5_SADL adl7 GND efet w=15 l=7
+ ad=1947 pd=452 as=2485 ps=626 
M3922 Vdd n_548 n_548 GND dfet w=9 l=20
+ ad=0 pd=0 as=480 ps=130 
M3923 x7 dpc3_SBX sb7 GND efet w=11 l=8
+ ad=0 pd=0 as=0 ps=0 
M3924 n_721 dpc4_SSB sb7 GND efet w=16 l=8
+ ad=0 pd=0 as=0 ps=0 
M3925 GND nots7 n_721 GND efet w=44 l=6
+ ad=0 pd=0 as=0 ps=0 
M3926 n_548 s7 GND GND efet w=33 l=6
+ ad=879 pd=232 as=0 ps=0 
M3927 n_548 cclk nots7 GND efet w=12 l=8
+ ad=0 pd=0 as=283 ps=98 
M3928 n_721 dpc7_SS s7 GND efet w=12 l=8
+ ad=0 pd=0 as=352 ps=78 
M3929 s7 dpc6_SBS sb7 GND efet w=12 l=7
+ ad=0 pd=0 as=0 ps=0 
M3930 sb7 cclk Vdd GND efet w=22 l=7
+ ad=0 pd=0 as=0 ps=0 
M3931 adl6 dpc10_ADLADD alub6 GND efet w=12 l=7
+ ad=0 pd=0 as=596 ps=150 
M3932 alub6 dpc8_nDBADD n_351 GND efet w=12 l=7
+ ad=0 pd=0 as=973 ps=280 
M3933 alub6 dpc9_DBADD idb6 GND efet w=11 l=7
+ ad=0 pd=0 as=1974 ps=542 
M3934 GND idb6 n_351 GND efet w=60 l=7
+ ad=0 pd=0 as=0 ps=0 
M3935 n_351 n_351 Vdd GND dfet w=9 l=17
+ ad=343 pd=86 as=0 ps=0 
M3936 n_A_B_5 alua5 GND GND efet w=32 l=7
+ ad=0 pd=0 as=0 ps=0 
M3937 GND alub5 n_A_B_5 GND efet w=32 l=7
+ ad=0 pd=0 as=0 ps=0 
M3938 naluresult5 dpc15_ANDS nA_B5 GND efet w=11 l=8
+ ad=0 pd=0 as=0 ps=0 
M3939 Vdd n_A_B_5 n_A_B_5 GND dfet w=9 l=22
+ ad=0 pd=0 as=1428 ps=414 
M3940 n_1483 alua6 GND GND efet w=61 l=6
+ ad=366 pd=134 as=0 ps=0 
M3941 nA_B6 alub6 n_1483 GND efet w=61 l=6
+ ad=1089 pd=300 as=0 ps=0 
M3942 Vdd nA_B6 nA_B6 GND dfet w=10 l=22
+ ad=0 pd=0 as=2389 ps=732 
M3943 n_1583 nA_B4 n_AxB_4 GND efet w=33 l=7
+ ad=198 pd=78 as=0 ps=0 
M3944 GND A_B4 n_1583 GND efet w=33 l=6
+ ad=0 pd=0 as=0 ps=0 
M3945 C45 n_A_B_4 GND GND efet w=29 l=6
+ ad=854 pd=222 as=0 ps=0 
M3946 n_1310 nC34 C45 GND efet w=54 l=6
+ ad=277 pd=118 as=0 ps=0 
M3947 GND nA_B4 n_1310 GND efet w=52 l=7
+ ad=0 pd=0 as=0 ps=0 
M3948 n_375 n_AxB_4 GND GND efet w=35 l=7
+ ad=210 pd=82 as=0 ps=0 
M3949 n_AxBxC_4 C34 n_375 GND efet w=35 l=5
+ ad=911 pd=222 as=0 ps=0 
M3950 Vdd n_AxBxC_4 n_AxBxC_4 GND dfet w=9 l=18
+ ad=0 pd=0 as=487 ps=106 
M3951 naluresult4 dpc17_SUMS n_AxBxC_4 GND efet w=11 l=7
+ ad=0 pd=0 as=0 ps=0 
M3952 Vdd DA_C45 DA_C45 GND dfet w=9 l=17
+ ad=0 pd=0 as=1799 ps=574 
M3953 n_AxBxC_4 _AxB_4_nC34 GND GND efet w=30 l=6
+ ad=0 pd=0 as=0 ps=0 
M3954 _AxB_4_nC34 n_AxB_4 GND GND efet w=18 l=7
+ ad=531 pd=178 as=0 ps=0 
M3955 DA_C45 nC45 GND GND efet w=27 l=6
+ ad=296 pd=110 as=0 ps=0 
M3956 n_AxB_4 n_AxB_4 Vdd GND dfet w=9 l=17
+ ad=1195 pd=342 as=0 ps=0 
M3957 GND C34 _AxB_4_nC34 GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M3958 C45 C45 Vdd GND dfet w=9 l=9
+ ad=1183 pd=406 as=0 ps=0 
M3959 Vdd n_647 n_647 GND dfet w=8 l=17
+ ad=0 pd=0 as=2179 ps=700 
M3960 Vdd A_B5 A_B5 GND dfet w=9 l=16
+ ad=0 pd=0 as=890 ps=254 
M3961 n_647 nA_B5 GND GND efet w=18 l=7
+ ad=748 pd=196 as=0 ps=0 
M3962 Vdd _AxB_4_nC34 _AxB_4_nC34 GND dfet w=9 l=16
+ ad=0 pd=0 as=912 ps=280 
M3963 Vdd nC45 nC45 GND dfet w=10 l=17
+ ad=0 pd=0 as=2281 ps=708 
M3964 n_1218 n_1218 Vdd GND dfet w=9 l=17
+ ad=1174 pd=344 as=0 ps=0 
M3965 Vdd alucout alucout GND dfet w=11 l=7
+ ad=0 pd=0 as=7047 ps=2420 
M3966 Vdd n_757 n_757 GND dfet w=9 l=16
+ ad=0 pd=0 as=2795 ps=986 
M3967 n_939 n_647 GND GND efet w=53 l=6
+ ad=371 pd=120 as=0 ps=0 
M3968 n_757 DA_C45 n_939 GND efet w=53 l=6
+ ad=675 pd=176 as=0 ps=0 
M3969 nC45 C45 GND GND efet w=18 l=6
+ ad=299 pd=98 as=0 ps=0 
M3970 GND n_A_B_5 A_B5 GND efet w=23 l=7
+ ad=0 pd=0 as=565 ps=170 
M3971 n_165 A_B5 GND GND efet w=55 l=6
+ ad=327 pd=122 as=0 ps=0 
M3972 nC56 C45 n_165 GND efet w=55 l=6
+ ad=782 pd=226 as=0 ps=0 
M3973 n_AxB_5 dpc16_EORS naluresult5 GND efet w=11 l=7
+ ad=456 pd=140 as=0 ps=0 
M3974 GND AxB5 n_AxB_5 GND efet w=29 l=7
+ ad=0 pd=0 as=0 ps=0 
M3975 AxB5 n_647 GND GND efet w=18 l=6
+ ad=579 pd=164 as=0 ps=0 
M3976 GND n_A_B_5 AxB5 GND efet w=18 l=8
+ ad=0 pd=0 as=0 ps=0 
M3977 GND n_647 nC56 GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M3978 n_547 AxB5 GND GND efet w=35 l=6
+ ad=210 pd=82 as=0 ps=0 
M3979 n_AxBxC_5 nC45 n_547 GND efet w=35 l=6
+ ad=876 pd=210 as=0 ps=0 
M3980 Vdd n_AxBxC_5 n_AxBxC_5 GND dfet w=9 l=18
+ ad=0 pd=0 as=478 ps=112 
M3981 n_1257 n_1218 GND GND efet w=35 l=7
+ ad=1122 pd=268 as=0 ps=0 
M3982 alucout notalucout GND GND efet w=76 l=6
+ ad=969 pd=262 as=0 ps=0 
M3983 n_1257 notalucout GND GND efet w=38 l=7
+ ad=0 pd=0 as=0 ps=0 
M3984 n_1257 n_1257 Vdd GND dfet w=10 l=10
+ ad=3784 pd=1410 as=0 ps=0 
M3985 n_AxBxC_5 n_AxB5__C45 GND GND efet w=26 l=6
+ ad=0 pd=0 as=0 ps=0 
M3986 naluresult5 dpc17_SUMS n_AxBxC_5 GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M3987 n_AxB5__C45 AxB5 GND GND efet w=18 l=6
+ ad=531 pd=164 as=0 ps=0 
M3988 n_AxB_5 n_AxB_5 Vdd GND dfet w=9 l=17
+ ad=435 pd=122 as=0 ps=0 
M3989 AxB5 AxB5 Vdd GND dfet w=10 l=16
+ ad=2291 pd=712 as=0 ps=0 
M3990 GND nC45 n_AxB5__C45 GND efet w=36 l=7
+ ad=0 pd=0 as=0 ps=0 
M3991 Vdd nC56 nC56 GND dfet w=9 l=10
+ ad=0 pd=0 as=1479 ps=480 
M3992 n_570 AxB5 GND GND efet w=26 l=6
+ ad=1103 pd=306 as=0 ps=0 
M3993 GND n_647 n_570 GND efet w=26 l=6
+ ad=0 pd=0 as=0 ps=0 
M3994 n_570 DA_C45 GND GND efet w=26 l=7
+ ad=0 pd=0 as=0 ps=0 
M3995 GND n_122 n_570 GND efet w=26 l=6
+ ad=0 pd=0 as=0 ps=0 
M3996 A_B6 A_B6 Vdd GND dfet w=9 l=16
+ ad=880 pd=246 as=0 ps=0 
M3997 nA_B6 dpc14_SRS naluresult5 GND efet w=11 l=7
+ ad=0 pd=0 as=0 ps=0 
M3998 naluresult6 dpc13_ORS n_A_B_6 GND efet w=12 l=7
+ ad=1717 pd=450 as=962 ps=278 
M3999 GND dpc12_0ADD alua6 GND efet w=13 l=7
+ ad=0 pd=0 as=539 ps=136 
M4000 alua6 dpc11_SBADD sb6 GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M4001 adl7 dpc10_ADLADD alub7 GND efet w=10 l=8
+ ad=0 pd=0 as=610 ps=148 
M4002 alub7 dpc8_nDBADD n_423 GND efet w=12 l=8
+ ad=0 pd=0 as=981 ps=274 
M4003 alub7 dpc9_DBADD idb7 GND efet w=12 l=7
+ ad=0 pd=0 as=2101 ps=560 
M4004 GND idb7 n_423 GND efet w=60 l=7
+ ad=0 pd=0 as=0 ps=0 
M4005 n_423 n_423 Vdd GND dfet w=8 l=17
+ ad=352 pd=86 as=0 ps=0 
M4006 n_A_B_6 alua6 GND GND efet w=30 l=6
+ ad=0 pd=0 as=0 ps=0 
M4007 GND alub6 n_A_B_6 GND efet w=30 l=7
+ ad=0 pd=0 as=0 ps=0 
M4008 Vdd n_A_B_6 n_A_B_6 GND dfet w=10 l=22
+ ad=0 pd=0 as=1643 ps=516 
M4009 n_1695 alua7 GND GND efet w=61 l=6
+ ad=366 pd=134 as=0 ps=0 
M4010 nA_B7 alub7 n_1695 GND efet w=61 l=7
+ ad=1431 pd=394 as=0 ps=0 
M4011 Vdd nA_B7 nA_B7 GND dfet w=10 l=21
+ ad=0 pd=0 as=1708 ps=526 
M4012 A_B6 n_A_B_6 GND GND efet w=18 l=6
+ ad=514 pd=162 as=0 ps=0 
M4013 n_AxB5__C45 n_AxB5__C45 Vdd GND dfet w=10 l=18
+ ad=781 pd=228 as=0 ps=0 
M4014 n_570 n_570 Vdd GND dfet w=10 l=13
+ ad=2490 pd=806 as=0 ps=0 
M4015 GND nA_B6 n_1038 GND efet w=36 l=6
+ ad=0 pd=0 as=392 ps=130 
M4016 Vdd C56 C56 GND dfet w=9 l=16
+ ad=0 pd=0 as=1145 ps=330 
M4017 C56 nC56 GND GND efet w=18 l=6
+ ad=386 pd=126 as=0 ps=0 
M4018 naluresult6 dpc15_ANDS nA_B6 GND efet w=12 l=7
+ ad=0 pd=0 as=0 ps=0 
M4019 n_AxB_6 dpc16_EORS naluresult6 GND efet w=12 l=7
+ ad=828 pd=252 as=0 ps=0 
M4020 n_482 nA_B6 n_AxB_6 GND efet w=34 l=6
+ ad=204 pd=80 as=0 ps=0 
M4021 GND A_B6 n_482 GND efet w=34 l=7
+ ad=0 pd=0 as=0 ps=0 
M4022 C67 n_A_B_6 GND GND efet w=28 l=6
+ ad=838 pd=220 as=0 ps=0 
M4023 n_112 nC56 C67 GND efet w=54 l=6
+ ad=328 pd=120 as=0 ps=0 
M4024 GND nA_B6 n_112 GND efet w=53 l=6
+ ad=0 pd=0 as=0 ps=0 
M4025 n_1390 n_AxB_6 GND GND efet w=35 l=7
+ ad=175 pd=80 as=0 ps=0 
M4026 n_AxBxC_6 C56 n_1390 GND efet w=35 l=7
+ ad=841 pd=218 as=0 ps=0 
M4027 Vdd n_AxBxC_6 n_AxBxC_6 GND dfet w=10 l=17
+ ad=0 pd=0 as=458 ps=106 
M4028 n_1038 n_1038 Vdd GND dfet w=10 l=15
+ ad=821 pd=312 as=0 ps=0 
M4029 naluresult6 dpc17_SUMS n_AxBxC_6 GND efet w=11 l=7
+ ad=0 pd=0 as=0 ps=0 
M4030 n_AxBxC_6 _AxB_6_nC56 GND GND efet w=29 l=6
+ ad=0 pd=0 as=0 ps=0 
M4031 _AxB_6_nC56 n_AxB_6 GND GND efet w=17 l=7
+ ad=540 pd=178 as=0 ps=0 
M4032 nA_B7 dpc14_SRS naluresult6 GND efet w=11 l=7
+ ad=0 pd=0 as=0 ps=0 
M4033 naluresult7 dpc13_ORS n_A_B_7 GND efet w=12 l=7
+ ad=1297 pd=326 as=986 ps=280 
M4034 GND dpc12_0ADD alua7 GND efet w=12 l=7
+ ad=0 pd=0 as=535 ps=140 
M4035 alua7 dpc11_SBADD sb7 GND efet w=11 l=9
+ ad=0 pd=0 as=0 ps=0 
M4036 n_A_B_7 alua7 GND GND efet w=31 l=6
+ ad=0 pd=0 as=0 ps=0 
M4037 GND alub7 n_A_B_7 GND efet w=31 l=6
+ ad=0 pd=0 as=0 ps=0 
M4038 naluresult7 dpc14_SRS Vdd GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M4039 naluresult7 dpc15_ANDS nA_B7 GND efet w=10 l=7
+ ad=0 pd=0 as=0 ps=0 
M4040 n_AxB_6 n_AxB_6 Vdd GND dfet w=9 l=10
+ ad=1889 pd=598 as=0 ps=0 
M4041 C67 C67 Vdd GND dfet w=10 l=10
+ ad=3132 pd=1004 as=0 ps=0 
M4042 GND C56 _AxB_6_nC56 GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M4043 Vdd n_748 n_748 GND dfet w=9 l=17
+ ad=0 pd=0 as=996 ps=312 
M4044 Vdd A_B7 A_B7 GND dfet w=9 l=17
+ ad=0 pd=0 as=896 ps=264 
M4045 n_748 nA_B7 GND GND efet w=19 l=6
+ ad=706 pd=192 as=0 ps=0 
M4046 Vdd n_122 n_122 GND dfet w=9 l=16
+ ad=0 pd=0 as=1223 ps=390 
M4047 n_122 n_AxB_6 GND GND efet w=35 l=6
+ ad=569 pd=182 as=0 ps=0 
M4048 n_269 AxB7 GND GND efet w=26 l=7
+ ad=582 pd=156 as=0 ps=0 
M4049 GND n_1038 n_269 GND efet w=26 l=6
+ ad=0 pd=0 as=0 ps=0 
M4050 Vdd _AxB_6_nC56 _AxB_6_nC56 GND dfet w=9 l=16
+ ad=0 pd=0 as=892 ps=276 
M4051 Vdd nC67 nC67 GND dfet w=9 l=17
+ ad=0 pd=0 as=1139 ps=336 
M4052 nC67 C67 GND GND efet w=18 l=6
+ ad=280 pd=96 as=0 ps=0 
M4053 n_1030 n_757 GND GND efet w=51 l=6
+ ad=1839 pd=420 as=0 ps=0 
M4054 n_269 n_269 Vdd GND dfet w=10 l=17
+ ad=1188 pd=368 as=0 ps=0 
M4055 GND n_AxB_6 n_1030 GND efet w=52 l=6
+ ad=0 pd=0 as=0 ps=0 
M4056 GND n_A_B_7 A_B7 GND efet w=23 l=7
+ ad=0 pd=0 as=606 ps=196 
M4057 n_1617 A_B7 GND GND efet w=55 l=6
+ ad=295 pd=122 as=0 ps=0 
M4058 nC78 C67 n_1617 GND efet w=55 l=6
+ ad=799 pd=226 as=0 ps=0 
M4059 n_AxB_7 dpc16_EORS naluresult7 GND efet w=11 l=7
+ ad=469 pd=134 as=0 ps=0 
M4060 Vdd n_A_B_7 n_A_B_7 GND dfet w=9 l=22
+ ad=0 pd=0 as=2858 ps=830 
M4061 dpc0_YSB cclk GND GND efet w=27 l=8
+ ad=0 pd=0 as=0 ps=0 
M4062 dpc1_SBY cclk GND GND efet w=28 l=8
+ ad=0 pd=0 as=0 ps=0 
M4063 dpc2_XSB cclk GND GND efet w=25 l=8
+ ad=0 pd=0 as=0 ps=0 
M4064 dpc3_SBX cclk GND GND efet w=27 l=8
+ ad=0 pd=0 as=0 ps=0 
M4065 GND AxB7 n_AxB_7 GND efet w=29 l=7
+ ad=0 pd=0 as=0 ps=0 
M4066 AxB7 n_748 GND GND efet w=24 l=7
+ ad=563 pd=170 as=0 ps=0 
M4067 GND n_A_B_7 AxB7 GND efet w=17 l=7
+ ad=0 pd=0 as=0 ps=0 
M4068 GND n_748 nC78 GND efet w=26 l=6
+ ad=0 pd=0 as=0 ps=0 
M4069 n_1013 AxB7 GND GND efet w=35 l=7
+ ad=175 pd=80 as=0 ps=0 
M4070 n_AxBxC_7 nC67 n_1013 GND efet w=35 l=7
+ ad=866 pd=218 as=0 ps=0 
M4071 Vdd n_AxBxC_7 n_AxBxC_7 GND dfet w=9 l=16
+ ad=0 pd=0 as=436 ps=104 
M4072 n_1030 n_269 DC78 GND efet w=60 l=6
+ ad=0 pd=0 as=1343 ps=412 
M4073 n_1030 n_570 DC78 GND efet w=59 l=7
+ ad=0 pd=0 as=0 ps=0 
M4074 n_AxBxC_7 n_AxB7__C67 GND GND efet w=30 l=6
+ ad=0 pd=0 as=0 ps=0 
M4075 naluresult7 dpc17_SUMS n_AxBxC_7 GND efet w=11 l=8
+ ad=0 pd=0 as=0 ps=0 
M4076 n_AxB_7 n_AxB_7 Vdd GND dfet w=10 l=17
+ ad=443 pd=120 as=0 ps=0 
M4077 AxB7 AxB7 Vdd GND dfet w=9 l=16
+ ad=3048 pd=980 as=0 ps=0 
M4078 n_AxB7__C67 AxB7 GND GND efet w=18 l=7
+ ad=495 pd=162 as=0 ps=0 
M4079 GND nC67 n_AxB7__C67 GND efet w=34 l=7
+ ad=0 pd=0 as=0 ps=0 
M4080 alu1 alu1 Vdd GND dfet w=9 l=12
+ ad=893 pd=272 as=0 ps=0 
M4081 dpc24_ACSB n_1247 GND GND efet w=73 l=5
+ ad=0 pd=0 as=0 ps=0 
M4082 GND n_1335 dpc24_ACSB GND efet w=76 l=6
+ ad=0 pd=0 as=0 ps=0 
M4083 dpc26_ACDB n_800 GND GND efet w=76 l=6
+ ad=0 pd=0 as=0 ps=0 
M4084 n_849 n_321 GND GND efet w=25 l=7
+ ad=363 pd=106 as=0 ps=0 
M4085 Vdd n_255 n_255 GND dfet w=9 l=15
+ ad=0 pd=0 as=1203 ps=354 
M4086 n_1323 n_631 GND GND efet w=25 l=6
+ ad=348 pd=106 as=0 ps=0 
M4087 Vdd n_611 dpc31_PCHPCH GND dfet w=10 l=11
+ ad=0 pd=0 as=1890 ps=396 
M4088 n_849 n_849 Vdd GND dfet w=9 l=15
+ ad=1253 pd=358 as=0 ps=0 
M4089 n_1413 n_1260 GND GND efet w=24 l=7
+ ad=354 pd=106 as=0 ps=0 
M4090 n_1518 n_1270 GND GND efet w=25 l=6
+ ad=355 pd=104 as=0 ps=0 
M4091 n_818 n_265 GND GND efet w=54 l=6
+ ad=876 pd=220 as=0 ps=0 
M4092 Vdd n_818 n_818 GND dfet w=10 l=14
+ ad=0 pd=0 as=1153 ps=344 
M4093 n_1480 n_1581 dpc36_nIPC GND efet w=154 l=6
+ ad=0 pd=0 as=0 ps=0 
M4094 pipeUNK17 cclk n_334 GND efet w=12 l=9
+ ad=233 pd=78 as=0 ps=0 
M4095 nop_set_C cclk pipeUNK08 GND efet w=12 l=9
+ ad=0 pd=0 as=170 ps=76 
M4096 n_513 n_885 GND GND efet w=52 l=6
+ ad=0 pd=0 as=0 ps=0 
M4097 Vdd n_513 n_513 GND dfet w=10 l=8
+ ad=0 pd=0 as=203 ps=72 
M4098 n_553 n_1662 GND GND efet w=30 l=7
+ ad=1155 pd=302 as=0 ps=0 
M4099 n_553 n_781 GND GND efet w=41 l=7
+ ad=0 pd=0 as=0 ps=0 
M4100 n_954 n_954 Vdd GND dfet w=11 l=12
+ ad=4193 pd=1400 as=0 ps=0 
M4101 GND n_954 n_513 GND efet w=41 l=7
+ ad=0 pd=0 as=0 ps=0 
M4102 GND pipeUNK08 n_954 GND efet w=83 l=6
+ ad=0 pd=0 as=1076 ps=270 
M4103 n_1379 cclk pipeUNK07 GND efet w=11 l=9
+ ad=0 pd=0 as=119 ps=60 
M4104 Vdd n_1379 n_1379 GND dfet w=10 l=18
+ ad=0 pd=0 as=450 ps=102 
M4105 n_327 cclk pipeUNK09 GND efet w=15 l=8
+ ad=0 pd=0 as=160 ps=78 
M4106 GND pipeUNK09 n_941 GND efet w=62 l=6
+ ad=0 pd=0 as=488 ps=172 
M4107 pipeUNK11 cclk n_862 GND efet w=12 l=7
+ ad=163 pd=76 as=0 ps=0 
M4108 Vdd fetch fetch GND dfet w=9 l=10
+ ad=0 pd=0 as=9410 ps=2802 
M4109 n_941 pipeUNK07 n_1111 GND efet w=76 l=6
+ ad=0 pd=0 as=1087 ps=250 
M4110 Vdd n_774 n_774 GND dfet w=10 l=18
+ ad=0 pd=0 as=1876 ps=618 
M4111 n_513 cclk pipeUNK06 GND efet w=12 l=8
+ ad=0 pd=0 as=189 ps=82 
M4112 n_754 n_754 Vdd GND dfet w=10 l=19
+ ad=4647 pd=1464 as=0 ps=0 
M4113 n_1225 cclk n_1121 GND efet w=12 l=10
+ ad=0 pd=0 as=144 ps=66 
M4114 n_1705 cclk n_1020 GND efet w=12 l=10
+ ad=0 pd=0 as=226 ps=80 
M4115 n_104 cclk n_1221 GND efet w=12 l=9
+ ad=0 pd=0 as=226 ps=80 
M4116 n_754 n_1673 GND GND efet w=40 l=7
+ ad=1270 pd=272 as=0 ps=0 
M4117 n_1422 pipeUNK06 n_754 GND efet w=77 l=5
+ ad=519 pd=190 as=0 ps=0 
M4118 GND pipeUNK09 n_1422 GND efet w=90 l=7
+ ad=0 pd=0 as=0 ps=0 
M4119 n_781 pipeUNK09 GND GND efet w=77 l=6
+ ad=0 pd=0 as=0 ps=0 
M4120 Vdd n_781 n_781 GND dfet w=10 l=10
+ ad=0 pd=0 as=6320 ps=2092 
M4121 n_1111 n_1111 Vdd GND dfet w=10 l=23
+ ad=3848 pd=1116 as=0 ps=0 
M4122 nnT2BR cclk n_1269 GND efet w=13 l=8
+ ad=0 pd=0 as=179 ps=74 
M4123 Vdd n_1401 n_1401 GND dfet w=10 l=18
+ ad=0 pd=0 as=836 ps=264 
M4124 fetch n_1214 GND GND efet w=38 l=7
+ ad=0 pd=0 as=0 ps=0 
M4125 GND pipeUNK11 n_1214 GND efet w=44 l=7
+ ad=0 pd=0 as=580 ps=150 
M4126 Vdd n_1214 n_1214 GND dfet w=11 l=15
+ ad=0 pd=0 as=912 ps=284 
M4127 pd3_clearIR clearIR GND GND efet w=30 l=7
+ ad=0 pd=0 as=0 ps=0 
M4128 pd4_clearIR pd4 GND GND efet w=75 l=7
+ ad=0 pd=0 as=0 ps=0 
M4129 GND clearIR pd5_clearIR GND efet w=30 l=7
+ ad=0 pd=0 as=0 ps=0 
M4130 pd0_clearIR clearIR GND GND efet w=30 l=6
+ ad=0 pd=0 as=0 ps=0 
M4131 GND clearIR pd1_clearIR GND efet w=31 l=7
+ ad=0 pd=0 as=0 ps=0 
M4132 pd7_clearIR clearIR GND GND efet w=41 l=6
+ ad=1057 pd=300 as=0 ps=0 
M4133 pd3_clearIR pd3_clearIR Vdd GND dfet w=10 l=10
+ ad=2003 pd=648 as=0 ps=0 
M4134 Vdd pd4_clearIR pd4_clearIR GND dfet w=10 l=11
+ ad=0 pd=0 as=2353 ps=764 
M4135 GND pd7 pd7_clearIR GND efet w=90 l=7
+ ad=0 pd=0 as=0 ps=0 
M4136 pd2_clearIR pd2 GND GND efet w=101 l=7
+ ad=1018 pd=296 as=0 ps=0 
M4137 GND clearIR pd2_clearIR GND efet w=31 l=6
+ ad=0 pd=0 as=0 ps=0 
M4138 pd6_clearIR clearIR GND GND efet w=31 l=7
+ ad=1009 pd=292 as=0 ps=0 
M4139 GND pd6 pd6_clearIR GND efet w=88 l=7
+ ad=0 pd=0 as=0 ps=0 
M4140 pd5_clearIR pd5_clearIR Vdd GND dfet w=10 l=11
+ ad=2520 pd=738 as=0 ps=0 
M4141 pd0_clearIR pd0_clearIR Vdd GND dfet w=11 l=9
+ ad=2205 pd=752 as=0 ps=0 
M4142 pd1_clearIR pd1_clearIR Vdd GND dfet w=10 l=10
+ ad=2321 pd=770 as=0 ps=0 
M4143 pd7_clearIR pd7_clearIR Vdd GND dfet w=10 l=10
+ ad=2335 pd=754 as=0 ps=0 
M4144 pd2_clearIR pd2_clearIR Vdd GND dfet w=10 l=10
+ ad=2237 pd=748 as=0 ps=0 
M4145 pd6_clearIR pd6_clearIR Vdd GND dfet w=11 l=10
+ ad=3257 pd=1066 as=0 ps=0 
M4146 pd4 cclk n_1075 GND efet w=15 l=7
+ ad=226 pd=88 as=1446 ps=356 
M4147 pd3 cclk n_1281 GND efet w=16 l=9
+ ad=178 pd=76 as=1451 ps=348 
M4148 pd5 cclk n_1588 GND efet w=15 l=9
+ ad=154 pd=62 as=1560 ps=364 
M4149 pd0 cclk n_93 GND efet w=16 l=9
+ ad=175 pd=78 as=1557 ps=360 
M4150 pd1 cclk n_1319 GND efet w=14 l=9
+ ad=144 pd=60 as=1476 ps=346 
M4151 pd7 cclk n_62 GND efet w=15 l=9
+ ad=164 pd=74 as=1414 ps=356 
M4152 pd2 cclk n_111 GND efet w=15 l=9
+ ad=152 pd=62 as=1457 ps=340 
M4153 pd6 cclk n_374 GND efet w=15 l=9
+ ad=219 pd=78 as=1439 ps=378 
M4154 GND op_clv n_340 GND efet w=45 l=6
+ ad=0 pd=0 as=574 ps=150 
M4155 n_503 notir5 GND GND efet w=36 l=6
+ ad=475 pd=120 as=0 ps=0 
M4156 n_340 n_340 Vdd GND dfet w=10 l=16
+ ad=447 pd=116 as=0 ps=0 
M4157 Vdd n_587 n_587 GND dfet w=10 l=18
+ ad=0 pd=0 as=3507 ps=1190 
M4158 n_340 cclk pipeUNK12 GND efet w=12 l=8
+ ad=0 pd=0 as=142 ps=62 
M4159 n_1673 cclk op_T__bit GND efet w=12 l=8
+ ad=149 pd=60 as=0 ps=0 
M4160 n_160 op_SRS GND GND efet w=33 l=6
+ ad=1054 pd=282 as=0 ps=0 
M4161 GND n_781 n_160 GND efet w=30 l=7
+ ad=0 pd=0 as=0 ps=0 
M4162 n_1049 cclk n_160 GND efet w=13 l=8
+ ad=149 pd=68 as=0 ps=0 
M4163 GND n_1049 n_507 GND efet w=58 l=6
+ ad=0 pd=0 as=689 ps=188 
M4164 n_160 n_160 Vdd GND dfet w=10 l=13
+ ad=325 pd=94 as=0 ps=0 
M4165 n_507 n_507 Vdd GND dfet w=10 l=15
+ ad=1101 pd=340 as=0 ps=0 
M4166 Vdd n_279 n_279 GND dfet w=9 l=15
+ ad=0 pd=0 as=1123 ps=352 
M4167 n_279 n_253 GND GND efet w=33 l=7
+ ad=1081 pd=252 as=0 ps=0 
M4168 n_279 n_954 GND GND efet w=23 l=6
+ ad=0 pd=0 as=0 ps=0 
M4169 GND n_507 n_279 GND efet w=24 l=6
+ ad=0 pd=0 as=0 ps=0 
M4170 n_1692 n_270 n_1082 GND efet w=35 l=6
+ ad=193 pd=82 as=2477 ps=578 
M4171 GND n_253 n_1692 GND efet w=35 l=6
+ ad=0 pd=0 as=0 ps=0 
M4172 GND pipeUNK06 n_755 GND efet w=61 l=7
+ ad=0 pd=0 as=787 ps=204 
M4173 n_1401 n_1269 GND GND efet w=56 l=6
+ ad=749 pd=206 as=0 ps=0 
M4174 n_1249 n_1269 GND GND efet w=90 l=7
+ ad=747 pd=168 as=0 ps=0 
M4175 n_755 n_755 Vdd GND dfet w=10 l=18
+ ad=4389 pd=1488 as=0 ps=0 
M4176 Vdd n_771 n_771 GND dfet w=10 l=14
+ ad=0 pd=0 as=2531 ps=798 
M4177 GND pipeUNK01 n_1198 GND efet w=62 l=6
+ ad=0 pd=0 as=601 ps=166 
M4178 Vdd n_503 n_503 GND dfet w=10 l=16
+ ad=0 pd=0 as=752 ps=204 
M4179 GND pipeUNK12 n_587 GND efet w=53 l=6
+ ad=0 pd=0 as=775 ps=204 
M4180 n_1198 n_1401 n_626 GND efet w=36 l=6
+ ad=0 pd=0 as=1063 ps=250 
M4181 n_626 DBNeg n_1249 GND efet w=45 l=7
+ ad=0 pd=0 as=0 ps=0 
M4182 Vdd n_1110 n_1110 GND dfet w=10 l=10
+ ad=0 pd=0 as=1199 ps=388 
M4183 n_626 n_626 Vdd GND dfet w=9 l=19
+ ad=438 pd=114 as=0 ps=0 
M4184 pipeUNK01 cclk n_1110 GND efet w=12 l=9
+ ad=144 pd=56 as=1660 ps=398 
M4185 GND n_756 n_1110 GND efet w=134 l=7
+ ad=0 pd=0 as=0 ps=0 
M4186 n_626 cp1 n_756 GND efet w=11 l=8
+ ad=0 pd=0 as=220 ps=86 
M4187 GND n_1110 n_771 GND efet w=35 l=8
+ ad=0 pd=0 as=724 ps=198 
M4188 n_367 n_954 GND GND efet w=35 l=6
+ ad=335 pd=114 as=0 ps=0 
M4189 n_1082 n_206 n_367 GND efet w=37 l=6
+ ad=0 pd=0 as=0 ps=0 
M4190 n_186 n_507 n_1082 GND efet w=31 l=7
+ ad=155 pd=72 as=0 ps=0 
M4191 GND n_1224 n_186 GND efet w=31 l=7
+ ad=0 pd=0 as=0 ps=0 
M4192 Vdd n_132 n_132 GND dfet w=9 l=9
+ ad=0 pd=0 as=6213 ps=2188 
M4193 GND n_31 n_132 GND efet w=46 l=6
+ ad=0 pd=0 as=0 ps=0 
M4194 GND n_43 n_818 GND efet w=24 l=6
+ ad=0 pd=0 as=0 ps=0 
M4195 Vdd n_291 n_291 GND dfet w=9 l=11
+ ad=0 pd=0 as=1314 ps=392 
M4196 GND n_1121 n_291 GND efet w=78 l=6
+ ad=0 pd=0 as=844 ps=200 
M4197 n_1277 n_1020 GND GND efet w=72 l=6
+ ad=784 pd=206 as=0 ps=0 
M4198 Vdd n_1277 n_1277 GND dfet w=10 l=11
+ ad=0 pd=0 as=1159 ps=382 
M4199 Vdd n_321 dpc33_PCHDB GND dfet w=8 l=9
+ ad=0 pd=0 as=1187 ps=278 
M4200 n_1323 n_1323 Vdd GND dfet w=9 l=14
+ ad=1179 pd=362 as=0 ps=0 
M4201 GND n_1247 dpc26_ACDB GND efet w=75 l=6
+ ad=0 pd=0 as=0 ps=0 
M4202 dpc30_ADHPCH n_1247 GND GND efet w=77 l=8
+ ad=0 pd=0 as=0 ps=0 
M4203 GND n_228 dpc30_ADHPCH GND efet w=78 l=7
+ ad=0 pd=0 as=0 ps=0 
M4204 dpc31_PCHPCH n_1247 GND GND efet w=76 l=8
+ ad=0 pd=0 as=0 ps=0 
M4205 GND n_255 dpc31_PCHPCH GND efet w=75 l=6
+ ad=0 pd=0 as=0 ps=0 
M4206 GND n_849 dpc33_PCHDB GND efet w=97 l=7
+ ad=0 pd=0 as=0 ps=0 
M4207 Vdd n_631 dpc37_PCLDB GND dfet w=8 l=9
+ ad=0 pd=0 as=1232 ps=274 
M4208 n_1413 n_1413 Vdd GND dfet w=10 l=15
+ ad=1277 pd=360 as=0 ps=0 
M4209 n_1462 n_1369 GND GND efet w=25 l=6
+ ad=364 pd=106 as=0 ps=0 
M4210 n_1518 n_1518 Vdd GND dfet w=10 l=14
+ ad=1324 pd=396 as=0 ps=0 
M4211 n_1043 n_818 GND GND efet w=26 l=6
+ ad=424 pd=110 as=0 ps=0 
M4212 GND dpc34_PCLC n_1007 GND efet w=22 l=6
+ ad=0 pd=0 as=358 ps=114 
M4213 adl2 dpc21_ADDADL alu2 GND efet w=15 l=8
+ ad=0 pd=0 as=1563 ps=422 
M4214 naluresult2 cclk notalu2 GND efet w=11 l=8
+ ad=0 pd=0 as=186 ps=74 
M4215 GND notalu2 alu2 GND efet w=101 l=6
+ ad=0 pd=0 as=0 ps=0 
M4216 alu2 dpc20_ADDSB06 sb2 GND efet w=21 l=8
+ ad=0 pd=0 as=0 ps=0 
M4217 alu2 alu2 Vdd GND dfet w=9 l=12
+ ad=1287 pd=400 as=0 ps=0 
M4218 adl3 dpc21_ADDADL alu3 GND efet w=16 l=8
+ ad=0 pd=0 as=1527 ps=422 
M4219 naluresult3 cclk notalu3 GND efet w=11 l=8
+ ad=0 pd=0 as=190 ps=74 
M4220 GND notalu3 alu3 GND efet w=100 l=6
+ ad=0 pd=0 as=0 ps=0 
M4221 alu3 dpc20_ADDSB06 sb3 GND efet w=21 l=8
+ ad=0 pd=0 as=0 ps=0 
M4222 alu3 alu3 Vdd GND dfet w=10 l=12
+ ad=358 pd=104 as=0 ps=0 
M4223 adl4 dpc21_ADDADL alu4 GND efet w=16 l=7
+ ad=0 pd=0 as=1598 ps=420 
M4224 naluresult4 cclk notalu4 GND efet w=12 l=9
+ ad=0 pd=0 as=174 ps=74 
M4225 GND notalu4 alu4 GND efet w=98 l=6
+ ad=0 pd=0 as=0 ps=0 
M4226 alu4 dpc20_ADDSB06 sb4 GND efet w=21 l=8
+ ad=0 pd=0 as=0 ps=0 
M4227 alu4 alu4 Vdd GND dfet w=9 l=12
+ ad=358 pd=104 as=0 ps=0 
M4228 adl5 dpc21_ADDADL alu5 GND efet w=16 l=8
+ ad=0 pd=0 as=1589 ps=422 
M4229 naluresult5 cclk notalu5 GND efet w=12 l=9
+ ad=0 pd=0 as=174 ps=74 
M4230 GND notalu5 alu5 GND efet w=99 l=7
+ ad=0 pd=0 as=0 ps=0 
M4231 Vdd notalucout notalucout GND dfet w=9 l=16
+ ad=0 pd=0 as=3974 ps=1284 
M4232 DC78 dpc18_nDAA GND GND efet w=27 l=6
+ ad=0 pd=0 as=0 ps=0 
M4233 Vdd nC78 nC78 GND dfet w=10 l=9
+ ad=0 pd=0 as=1420 ps=514 
M4234 n_1489 n_A_B_7 GND GND efet w=55 l=7
+ ad=555 pd=172 as=0 ps=0 
M4235 dpc6_SBS cclk GND GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M4236 dpc7_SS cclk GND GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M4237 dpc8_nDBADD cclk GND GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M4238 dpc9_DBADD cclk GND GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M4239 dpc10_ADLADD cclk GND GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M4240 dpc11_SBADD cclk GND GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M4241 dpc12_0ADD cclk GND GND efet w=26 l=8
+ ad=0 pd=0 as=0 ps=0 
M4242 n_637 nA_B7 GND GND efet w=24 l=6
+ ad=518 pd=166 as=0 ps=0 
M4243 GND C67 n_637 GND efet w=30 l=6
+ ad=0 pd=0 as=0 ps=0 
M4244 notaluvout C67 n_1489 GND efet w=52 l=7
+ ad=1059 pd=330 as=0 ps=0 
M4245 DC78 DC78 Vdd GND dfet w=9 l=11
+ ad=621 pd=194 as=0 ps=0 
M4246 n_AxB7__C67 n_AxB7__C67 Vdd GND dfet w=10 l=16
+ ad=751 pd=228 as=0 ps=0 
M4247 Vdd C78 C78 GND dfet w=9 l=8
+ ad=0 pd=0 as=304 ps=104 
M4248 notalucout DC78_phi2 GND GND efet w=42 l=6
+ ad=1073 pd=246 as=0 ps=0 
M4249 GND C78_phi2 notalucout GND efet w=42 l=6
+ ad=0 pd=0 as=0 ps=0 
M4250 alu5 dpc20_ADDSB06 sb5 GND efet w=21 l=7
+ ad=0 pd=0 as=0 ps=0 
M4251 alu5 alu5 Vdd GND dfet w=9 l=13
+ ad=867 pd=242 as=0 ps=0 
M4252 adl6 dpc21_ADDADL alu6 GND efet w=15 l=9
+ ad=0 pd=0 as=1563 ps=418 
M4253 naluresult6 cclk notalu6 GND efet w=11 l=9
+ ad=0 pd=0 as=178 ps=76 
M4254 GND notalu6 alu6 GND efet w=99 l=6
+ ad=0 pd=0 as=0 ps=0 
M4255 alu6 dpc20_ADDSB06 sb6 GND efet w=21 l=7
+ ad=0 pd=0 as=0 ps=0 
M4256 alu6 alu6 Vdd GND dfet w=9 l=12
+ ad=854 pd=262 as=0 ps=0 
M4257 notalu7 cclk naluresult7 GND efet w=11 l=8
+ ad=216 pd=78 as=0 ps=0 
M4258 n_1556 nDA_ADD1 GND GND efet w=34 l=7
+ ad=225 pd=86 as=0 ps=0 
M4259 n_986 nDA_ADD2 n_1556 GND efet w=37 l=7
+ ad=479 pd=132 as=0 ps=0 
M4260 Vdd n_986 n_986 GND dfet w=9 l=17
+ ad=0 pd=0 as=3627 ps=1274 
M4261 Vdd n_1682 n_1682 GND dfet w=9 l=17
+ ad=0 pd=0 as=798 ps=226 
M4262 n_36 n_36 Vdd GND dfet w=9 l=17
+ ad=1925 pd=654 as=0 ps=0 
M4263 n_36 n_8 GND GND efet w=19 l=7
+ ad=862 pd=252 as=0 ps=0 
M4264 n_867 nDA_ADD1 GND GND efet w=27 l=7
+ ad=746 pd=170 as=0 ps=0 
M4265 GND nDA_ADD2 n_867 GND efet w=34 l=7
+ ad=0 pd=0 as=0 ps=0 
M4266 n_867 n_867 Vdd GND dfet w=10 l=17
+ ad=1587 pd=480 as=0 ps=0 
M4267 Vdd nDA_ADD1 nDA_ADD1 GND dfet w=11 l=16
+ ad=0 pd=0 as=2021 ps=614 
M4268 n_1682 nDA_ADD1 GND GND efet w=18 l=7
+ ad=349 pd=120 as=0 ps=0 
M4269 n_150 n_1682 n_613 GND efet w=37 l=6
+ ad=389 pd=94 as=1311 ps=372 
M4270 GND n_8 n_150 GND efet w=35 l=7
+ ad=0 pd=0 as=0 ps=0 
M4271 n_36 n_600 GND GND efet w=21 l=7
+ ad=0 pd=0 as=0 ps=0 
M4272 n_1362 nDA_ADD1 GND GND efet w=53 l=6
+ ad=475 pd=142 as=0 ps=0 
M4273 n_613 n_600 n_1362 GND efet w=78 l=6
+ ad=0 pd=0 as=0 ps=0 
M4274 nDA_ADD1 alu1 GND GND efet w=46 l=7
+ ad=565 pd=158 as=0 ps=0 
M4275 nDA_ADD2 alu2 GND GND efet w=44 l=6
+ ad=448 pd=146 as=0 ps=0 
M4276 GND n_867 n_876 GND efet w=18 l=6
+ ad=0 pd=0 as=447 ps=138 
M4277 nDA_ADD2 nDA_ADD2 Vdd GND dfet w=10 l=17
+ ad=2225 pd=672 as=0 ps=0 
M4278 n_876 n_876 Vdd GND dfet w=9 l=16
+ ad=2057 pd=682 as=0 ps=0 
M4279 Vdd n_600 n_600 GND dfet w=9 l=10
+ ad=0 pd=0 as=3914 ps=1374 
M4280 n_600 n_1341 GND GND efet w=79 l=7
+ ad=930 pd=228 as=0 ps=0 
M4281 Vdd n_146 n_146 GND dfet w=10 l=12
+ ad=0 pd=0 as=354 ps=108 
M4282 GND n_1323 dpc37_PCLDB GND efet w=95 l=6
+ ad=0 pd=0 as=0 ps=0 
M4283 Vdd n_1260 dpc32_PCHADH GND dfet w=10 l=9
+ ad=0 pd=0 as=1256 ps=304 
M4284 GND n_1413 dpc32_PCHADH GND efet w=98 l=7
+ ad=0 pd=0 as=0 ps=0 
M4285 Vdd n_1270 dpc39_PCLPCL GND dfet w=9 l=10
+ ad=0 pd=0 as=1915 ps=346 
M4286 n_1462 n_1462 Vdd GND dfet w=10 l=14
+ ad=1264 pd=368 as=0 ps=0 
M4287 n_1043 n_1043 Vdd GND dfet w=10 l=14
+ ad=1228 pd=352 as=0 ps=0 
M4288 Vdd n_1369 dpc38_PCLADL GND dfet w=10 l=10
+ ad=0 pd=0 as=1190 ps=256 
M4289 GND n_1462 dpc38_PCLADL GND efet w=99 l=7
+ ad=0 pd=0 as=0 ps=0 
M4290 dpc39_PCLPCL n_1247 GND GND efet w=84 l=6
+ ad=0 pd=0 as=0 ps=0 
M4291 GND n_1518 dpc39_PCLPCL GND efet w=91 l=6
+ ad=0 pd=0 as=0 ps=0 
M4292 Vdd n_818 dpc40_ADLPCL GND dfet w=9 l=11
+ ad=0 pd=0 as=1718 ps=312 
M4293 n_1566 n_1221 GND GND efet w=70 l=6
+ ad=801 pd=202 as=0 ps=0 
M4294 Vdd n_1566 n_1566 GND dfet w=10 l=11
+ ad=0 pd=0 as=1129 ps=398 
M4295 GND n_334 Pout2 GND efet w=67 l=7
+ ad=0 pd=0 as=1198 ps=310 
M4296 p7 n_1045 GND GND efet w=67 l=7
+ ad=1171 pd=300 as=0 ps=0 
M4297 Vdd Pout2 Pout2 GND dfet w=10 l=10
+ ad=0 pd=0 as=278 ps=86 
M4298 p7 p7 Vdd GND dfet w=10 l=9
+ ad=264 pd=86 as=0 ps=0 
M4299 Pout2 H1x1 idb2 GND efet w=25 l=8
+ ad=0 pd=0 as=0 ps=0 
M4300 p7 H1x1 idb7 GND efet w=24 l=8
+ ad=0 pd=0 as=0 ps=0 
M4301 n_1007 n_1007 Vdd GND dfet w=10 l=17
+ ad=1101 pd=324 as=0 ps=0 
M4302 dpc40_ADLPCL n_1247 GND GND efet w=75 l=7
+ ad=0 pd=0 as=0 ps=0 
M4303 GND n_1043 dpc40_ADLPCL GND efet w=77 l=7
+ ad=0 pd=0 as=0 ps=0 
M4304 dpc35_PCHC n_1007 GND GND efet w=55 l=6
+ ad=2900 pd=802 as=0 ps=0 
M4305 n_1157 n_291 GND GND efet w=25 l=6
+ ad=352 pd=102 as=0 ps=0 
M4306 n_1157 n_1157 Vdd GND dfet w=10 l=14
+ ad=1270 pd=372 as=0 ps=0 
M4307 n_1441 n_1441 Vdd GND dfet w=10 l=14
+ ad=1354 pd=396 as=0 ps=0 
M4308 GND n_1277 n_1441 GND efet w=25 l=6
+ ad=0 pd=0 as=460 ps=116 
M4309 GND n_1566 n_1240 GND efet w=25 l=6
+ ad=0 pd=0 as=358 ps=102 
M4310 GND idb2 n_1573 GND efet w=72 l=6
+ ad=0 pd=0 as=816 ps=220 
M4311 DBNeg idb7 GND GND efet w=84 l=6
+ ad=747 pd=194 as=0 ps=0 
M4312 Vdd n_291 dpc41_DL_ADL GND dfet w=9 l=9
+ ad=0 pd=0 as=1203 ps=252 
M4313 Vdd n_1277 dpc42_DL_ADH GND dfet w=10 l=9
+ ad=0 pd=0 as=1118 ps=262 
M4314 n_1240 n_1240 Vdd GND dfet w=9 l=14
+ ad=1328 pd=388 as=0 ps=0 
M4315 n_1573 n_1573 Vdd GND dfet w=9 l=12
+ ad=3500 pd=1226 as=0 ps=0 
M4316 DBNeg DBNeg Vdd GND dfet w=10 l=8
+ ad=6758 pd=2352 as=0 ps=0 
M4317 GND n_90 p6 GND efet w=66 l=6
+ ad=0 pd=0 as=1165 ps=300 
M4318 Pout3 n_1194 GND GND efet w=99 l=6
+ ad=1543 pd=364 as=0 ps=0 
M4319 Vdd p6 p6 GND dfet w=10 l=11
+ ad=0 pd=0 as=291 ps=84 
M4320 Pout3 Pout3 Vdd GND dfet w=10 l=10
+ ad=4962 pd=1668 as=0 ps=0 
M4321 p6 H1x1 idb6 GND efet w=25 l=8
+ ad=0 pd=0 as=0 ps=0 
M4322 Pout3 H1x1 idb3 GND efet w=25 l=8
+ ad=0 pd=0 as=0 ps=0 
M4323 GND idb6 n_1416 GND efet w=73 l=6
+ ad=0 pd=0 as=800 ps=224 
M4324 n_1600 idb3 GND GND efet w=73 l=6
+ ad=800 pd=226 as=0 ps=0 
M4325 n_455 n_279 GND GND efet w=61 l=6
+ ad=366 pd=134 as=0 ps=0 
M4326 n_1082 pipeUNK16 n_455 GND efet w=61 l=6
+ ad=0 pd=0 as=0 ps=0 
M4327 n_31 p0 GND GND efet w=65 l=6
+ ad=1273 pd=308 as=0 ps=0 
M4328 Vdd n_1471 n_1471 GND dfet w=10 l=17
+ ad=0 pd=0 as=1451 ps=424 
M4329 p0 cp1 n_1082 GND efet w=13 l=8
+ ad=193 pd=70 as=0 ps=0 
M4330 n_31 n_31 Vdd GND dfet w=10 l=12
+ ad=8672 pd=2864 as=0 ps=0 
M4331 n_1471 D1x1 GND GND efet w=40 l=6
+ ad=434 pd=142 as=0 ps=0 
M4332 n_1082 n_1082 Vdd GND dfet w=10 l=21
+ ad=457 pd=110 as=0 ps=0 
M4333 n_31 cclk pipeUNK16 GND efet w=12 l=7
+ ad=0 pd=0 as=163 ps=64 
M4334 p4 n_1471 GND GND efet w=89 l=7
+ ad=1588 pd=386 as=0 ps=0 
M4335 p4 p4 Vdd GND dfet w=11 l=10
+ ad=282 pd=86 as=0 ps=0 
M4336 n_270 n_503 GND GND efet w=32 l=7
+ ad=486 pd=146 as=0 ps=0 
M4337 Vdd n_270 n_270 GND dfet w=10 l=13
+ ad=0 pd=0 as=11979 ps=4098 
M4338 pipeUNK02 cclk n_774 GND efet w=10 l=8
+ ad=146 pd=68 as=0 ps=0 
M4339 GND pipeUNK02 n_1492 GND efet w=41 l=6
+ ad=0 pd=0 as=517 ps=142 
M4340 GND db4 n_1075 GND efet w=135 l=7
+ ad=0 pd=0 as=0 ps=0 
M4341 n_1281 db3 GND GND efet w=138 l=6
+ ad=0 pd=0 as=0 ps=0 
M4342 n_1075 n_1075 Vdd GND dfet w=10 l=7
+ ad=175 pd=64 as=0 ps=0 
M4343 GND db5 n_1588 GND efet w=138 l=5
+ ad=0 pd=0 as=0 ps=0 
M4344 n_93 db0 GND GND efet w=143 l=11
+ ad=0 pd=0 as=0 ps=0 
M4345 Vdd n_1281 n_1281 GND dfet w=10 l=7
+ ad=0 pd=0 as=182 ps=66 
M4346 n_1588 n_1588 Vdd GND dfet w=10 l=7
+ ad=175 pd=64 as=0 ps=0 
M4347 Vdd n_1492 n_1492 GND dfet w=9 l=18
+ ad=0 pd=0 as=2536 ps=786 
M4348 GND db1 n_1319 GND efet w=138 l=7
+ ad=0 pd=0 as=0 ps=0 
M4349 n_62 db7 GND GND efet w=139 l=6
+ ad=0 pd=0 as=0 ps=0 
M4350 Vdd n_93 n_93 GND dfet w=10 l=8
+ ad=0 pd=0 as=200 ps=66 
M4351 n_1319 n_1319 Vdd GND dfet w=10 l=7
+ ad=175 pd=64 as=0 ps=0 
M4352 Vdd n_62 n_62 GND dfet w=10 l=6
+ ad=0 pd=0 as=150 ps=62 
M4353 n_111 n_111 Vdd GND dfet w=10 l=7
+ ad=175 pd=64 as=0 ps=0 
M4354 GND db2 n_111 GND efet w=123 l=7
+ ad=0 pd=0 as=0 ps=0 
M4355 GND db6 n_374 GND efet w=123 l=7
+ ad=0 pd=0 as=0 ps=0 
M4356 n_374 n_374 Vdd GND dfet w=9 l=8
+ ad=200 pd=66 as=0 ps=0 
M4357 pipeUNK04 cclk n_1194 GND efet w=12 l=8
+ ad=308 pd=84 as=1052 ps=290 
M4358 GND p3 n_1194 GND efet w=60 l=7
+ ad=0 pd=0 as=0 ps=0 
M4359 n_1495 cp1 p3 GND efet w=12 l=8
+ ad=1311 pd=284 as=184 ps=80 
M4360 n_1194 n_1194 Vdd GND dfet w=10 l=14
+ ad=2585 pd=806 as=0 ps=0 
M4361 n_1495 n_1495 Vdd GND dfet w=11 l=20
+ ad=380 pd=92 as=0 ps=0 
M4362 n_1644 n_1457 n_1495 GND efet w=33 l=6
+ ad=684 pd=160 as=0 ps=0 
M4363 GND pipeUNK04 n_1644 GND efet w=66 l=7
+ ad=0 pd=0 as=0 ps=0 
M4364 GND DBNeg n_648 GND efet w=47 l=6
+ ad=0 pd=0 as=273 ps=106 
M4365 n_648 n_754 n_1181 GND efet w=47 l=6
+ ad=0 pd=0 as=1245 ps=326 
M4366 n_1069 cclk n_1177 GND efet w=11 l=7
+ ad=0 pd=0 as=342 ps=112 
M4367 GND n_587 n_299 GND efet w=21 l=7
+ ad=0 pd=0 as=1373 ps=346 
M4368 x_op_T__adc_sbc cclk pipeUNK03 GND efet w=12 l=9
+ ad=0 pd=0 as=356 ps=108 
M4369 n_299 n_1245 n_1723 GND efet w=32 l=7
+ ad=0 pd=0 as=565 ps=154 
M4370 Vdd n_299 n_299 GND dfet w=10 l=20
+ ad=0 pd=0 as=715 ps=200 
M4371 n_1723 pipeUNK03 GND GND efet w=67 l=6
+ ad=0 pd=0 as=0 ps=0 
M4372 Vdd n_1614 n_1614 GND dfet w=10 l=18
+ ad=0 pd=0 as=1116 ps=304 
M4373 n_1614 n_1177 GND GND efet w=44 l=6
+ ad=1626 pd=438 as=0 ps=0 
M4374 n_1595 n_754 GND GND efet w=28 l=7
+ ad=312 pd=118 as=0 ps=0 
M4375 n_1181 n_1181 Vdd GND dfet w=10 l=20
+ ad=1179 pd=324 as=0 ps=0 
M4376 Vdd n_1595 n_1595 GND dfet w=10 l=16
+ ad=0 pd=0 as=1148 ps=334 
M4377 n_1181 n_1595 n_793 GND efet w=31 l=6
+ ad=0 pd=0 as=548 ps=150 
M4378 n_793 pipeUNK13 GND GND efet w=65 l=6
+ ad=0 pd=0 as=0 ps=0 
M4379 n_1614 pipeUNK03 GND GND efet w=42 l=6
+ ad=0 pd=0 as=0 ps=0 
M4380 GND n_1111 n_1470 GND efet w=32 l=7
+ ad=0 pd=0 as=192 ps=76 
M4381 n_1546 n_781 GND GND efet w=32 l=7
+ ad=192 pd=76 as=0 ps=0 
M4382 n_1495 n_1600 n_1546 GND efet w=32 l=6
+ ad=0 pd=0 as=0 ps=0 
M4383 n_1445 n_270 n_1495 GND efet w=32 l=7
+ ad=160 pd=74 as=0 ps=0 
M4384 GND n_1492 n_1445 GND efet w=32 l=6
+ ad=0 pd=0 as=0 ps=0 
M4385 n_1470 n_1416 n_299 GND efet w=32 l=7
+ ad=0 pd=0 as=0 ps=0 
M4386 GND n_1111 n_1614 GND efet w=20 l=7
+ ad=0 pd=0 as=0 ps=0 
M4387 pipeUNK13 cclk n_1045 GND efet w=12 l=10
+ ad=135 pd=70 as=814 ps=250 
M4388 n_1181 cp1 n_69 GND efet w=13 l=9
+ ad=0 pd=0 as=156 ps=80 
M4389 n_1045 n_1045 Vdd GND dfet w=11 l=12
+ ad=5012 pd=1594 as=0 ps=0 
M4390 GND n_69 n_1045 GND efet w=80 l=6
+ ad=0 pd=0 as=0 ps=0 
M4391 n_299 n_1614 n_1616 GND efet w=32 l=8
+ ad=0 pd=0 as=517 ps=152 
M4392 n_1457 n_1457 Vdd GND dfet w=11 l=14
+ ad=858 pd=264 as=0 ps=0 
M4393 n_1457 n_781 GND GND efet w=25 l=7
+ ad=880 pd=172 as=0 ps=0 
M4394 GND n_1492 n_1457 GND efet w=25 l=7
+ ad=0 pd=0 as=0 ps=0 
M4395 n_1616 pipeUNK05 GND GND efet w=68 l=6
+ ad=0 pd=0 as=0 ps=0 
M4396 n_307 n_31 GND GND efet w=38 l=7
+ ad=1428 pd=380 as=0 ps=0 
M4397 n_299 cp1 n_1625 GND efet w=13 l=8
+ ad=0 pd=0 as=191 ps=80 
M4398 GND nop_branch_bit7 n_307 GND efet w=40 l=6
+ ad=0 pd=0 as=0 ps=0 
M4399 GND n_1625 n_90 GND efet w=69 l=6
+ ad=0 pd=0 as=900 ps=242 
M4400 pipeUNK05 cclk n_90 GND efet w=13 l=8
+ ad=210 pd=72 as=0 ps=0 
M4401 n_307 n_846 GND GND efet w=41 l=6
+ ad=0 pd=0 as=0 ps=0 
M4402 GND n_31 Pout0 GND efet w=67 l=7
+ ad=0 pd=0 as=1099 ps=310 
M4403 Pout1 n_318 GND GND efet w=84 l=6
+ ad=1243 pd=324 as=0 ps=0 
M4404 n_1416 n_1416 Vdd GND dfet w=10 l=12
+ ad=3292 pd=1104 as=0 ps=0 
M4405 n_1600 n_1600 Vdd GND dfet w=10 l=11
+ ad=2259 pd=832 as=0 ps=0 
M4406 GND alucout n_206 GND efet w=126 l=6
+ ad=0 pd=0 as=0 ps=0 
M4407 p4 H1x1 idb4 GND efet w=25 l=7
+ ad=0 pd=0 as=0 ps=0 
M4408 GND dpc36_nIPC dpc34_PCLC GND efet w=56 l=8
+ ad=0 pd=0 as=4543 ps=1300 
M4409 n_146 cclk a0 GND efet w=12 l=7
+ ad=1655 pd=400 as=437 ps=136 
M4410 a0 dpc23_SBAC sb0 GND efet w=11 l=7
+ ad=0 pd=0 as=0 ps=0 
M4411 n_146 n_5 GND GND efet w=80 l=6
+ ad=0 pd=0 as=0 ps=0 
M4412 n_613 n_613 Vdd GND dfet w=10 l=16
+ ad=2232 pd=752 as=0 ps=0 
M4413 Vdd dasb1 dasb1 GND dfet w=9 l=17
+ ad=0 pd=0 as=390 ps=102 
M4414 GND a0 n_5 GND efet w=44 l=6
+ ad=0 pd=0 as=784 ps=192 
M4415 n_146 dpc26_ACDB idb0 GND efet w=13 l=8
+ ad=0 pd=0 as=0 ps=0 
M4416 idb0 dpc25_SBDB sb0 GND efet w=23 l=7
+ ad=0 pd=0 as=0 ps=0 
M4417 sb0 dpc24_ACSB n_146 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M4418 Vdd n_5 n_5 GND dfet w=10 l=16
+ ad=0 pd=0 as=1009 ps=290 
M4419 n_1322 n_320 GND GND efet w=35 l=6
+ ad=210 pd=82 as=0 ps=0 
M4420 dasb1 n_36 n_1322 GND efet w=35 l=6
+ ad=738 pd=182 as=0 ps=0 
M4421 a1 dpc23_SBAC dasb1 GND efet w=11 l=7
+ ad=453 pd=140 as=0 ps=0 
M4422 GND n_735 dasb1 GND efet w=18 l=6
+ ad=0 pd=0 as=0 ps=0 
M4423 n_735 n_320 GND GND efet w=23 l=6
+ ad=570 pd=158 as=0 ps=0 
M4424 GND n_36 n_735 GND efet w=25 l=6
+ ad=0 pd=0 as=0 ps=0 
M4425 n_1341 cclk n_695 GND efet w=11 l=8
+ ad=129 pd=56 as=747 ps=230 
M4426 Vdd n_695 n_695 GND dfet w=9 l=15
+ ad=0 pd=0 as=571 ps=170 
M4427 n_619 n_700 GND GND efet w=47 l=6
+ ad=280 pd=106 as=0 ps=0 
M4428 n_695 C34 n_619 GND efet w=47 l=6
+ ad=0 pd=0 as=0 ps=0 
M4429 n_320 sb1 GND GND efet w=54 l=7
+ ad=465 pd=146 as=0 ps=0 
M4430 n_735 n_735 Vdd GND dfet w=9 l=17
+ ad=892 pd=266 as=0 ps=0 
M4431 Vdd n_929 n_929 GND dfet w=10 l=12
+ ad=0 pd=0 as=327 ps=96 
M4432 n_929 cclk a1 GND efet w=12 l=8
+ ad=1586 pd=380 as=0 ps=0 
M4433 n_929 n_1549 GND GND efet w=80 l=7
+ ad=0 pd=0 as=0 ps=0 
M4434 GND a1 n_1549 GND efet w=46 l=6
+ ad=0 pd=0 as=670 ps=200 
M4435 Vdd n_320 n_320 GND dfet w=9 l=17
+ ad=0 pd=0 as=1020 ps=318 
M4436 Vdd dasb2 dasb2 GND dfet w=9 l=17
+ ad=0 pd=0 as=390 ps=102 
M4437 n_1656 n_1580 GND GND efet w=39 l=6
+ ad=209 pd=90 as=0 ps=0 
M4438 dasb2 n_613 n_1656 GND efet w=37 l=6
+ ad=786 pd=188 as=0 ps=0 
M4439 adh0 dpc27_SBADH sb0 GND efet w=21 l=7
+ ad=1645 pd=438 as=0 ps=0 
M4440 GND dpc28_0ADH0 adh0 GND efet w=21 l=8
+ ad=0 pd=0 as=0 ps=0 
M4441 n_929 dpc26_ACDB idb1 GND efet w=15 l=8
+ ad=0 pd=0 as=0 ps=0 
M4442 idb1 dpc25_SBDB sb1 GND efet w=22 l=7
+ ad=0 pd=0 as=0 ps=0 
M4443 sb1 dpc24_ACSB n_929 GND efet w=13 l=8
+ ad=0 pd=0 as=0 ps=0 
M4444 Vdd n_1549 n_1549 GND dfet w=9 l=16
+ ad=0 pd=0 as=1055 ps=284 
M4445 a2 dpc23_SBAC dasb2 GND efet w=11 l=7
+ ad=433 pd=138 as=0 ps=0 
M4446 Vdd n_1618 n_1618 GND dfet w=10 l=13
+ ad=0 pd=0 as=318 ps=98 
M4447 GND n_1159 dasb2 GND efet w=18 l=6
+ ad=0 pd=0 as=0 ps=0 
M4448 n_1159 n_1580 GND GND efet w=20 l=6
+ ad=520 pd=142 as=0 ps=0 
M4449 GND n_613 n_1159 GND efet w=24 l=6
+ ad=0 pd=0 as=0 ps=0 
M4450 n_1580 sb2 GND GND efet w=15 l=5
+ ad=634 pd=184 as=0 ps=0 
M4451 Vdd n_1580 n_1580 GND dfet w=8 l=14
+ ad=0 pd=0 as=905 ps=282 
M4452 n_1159 n_1159 Vdd GND dfet w=9 l=17
+ ad=885 pd=252 as=0 ps=0 
M4453 n_1580 sb2 GND GND efet w=46 l=6
+ ad=0 pd=0 as=0 ps=0 
M4454 Vdd dasb3 dasb3 GND dfet w=10 l=17
+ ad=0 pd=0 as=390 ps=102 
M4455 n_1179 C34 GND GND efet w=24 l=6
+ ad=1185 pd=346 as=0 ps=0 
M4456 GND dpc22_nDSA n_1179 GND efet w=21 l=7
+ ad=0 pd=0 as=0 ps=0 
M4457 n_1584 n_876 GND GND efet w=51 l=6
+ ad=275 pd=112 as=0 ps=0 
M4458 n_345 n_8 n_1584 GND efet w=50 l=7
+ ad=992 pd=228 as=0 ps=0 
M4459 n_1686 n_432 GND GND efet w=34 l=7
+ ad=170 pd=78 as=0 ps=0 
M4460 dasb3 n_345 n_1686 GND efet w=34 l=6
+ ad=735 pd=172 as=0 ps=0 
M4461 n_1618 cclk a2 GND efet w=11 l=8
+ ad=1613 pd=388 as=0 ps=0 
M4462 n_1618 n_419 GND GND efet w=81 l=6
+ ad=0 pd=0 as=0 ps=0 
M4463 GND a2 n_419 GND efet w=44 l=6
+ ad=0 pd=0 as=739 ps=204 
M4464 Vdd cclk adh0 GND efet w=23 l=7
+ ad=0 pd=0 as=0 ps=0 
M4465 GND dpc29_0ADH17 adh1 GND efet w=23 l=8
+ ad=0 pd=0 as=1644 ps=408 
M4466 adh1 dpc27_SBADH sb1 GND efet w=23 l=7
+ ad=0 pd=0 as=0 ps=0 
M4467 Vdd cclk adh1 GND efet w=24 l=6
+ ad=0 pd=0 as=0 ps=0 
M4468 dpc35_PCHC dpc35_PCHC Vdd GND dfet w=13 l=7
+ ad=5733 pd=2144 as=0 ps=0 
M4469 n_311 n_311 Vdd GND dfet w=9 l=16
+ ad=1361 pd=420 as=0 ps=0 
M4470 Vdd cclk adl0 GND efet w=22 l=7
+ ad=0 pd=0 as=0 ps=0 
M4471 Vdd n_919 n_919 GND dfet w=9 l=15
+ ad=0 pd=0 as=2179 ps=696 
M4472 n_1229 cclk npchp0 GND efet w=12 l=8
+ ad=931 pd=234 as=222 ps=80 
M4473 pchp0 dpc31_PCHPCH pch0 GND efet w=14 l=9
+ ad=1504 pd=376 as=590 ps=156 
M4474 pch0 dpc30_ADHPCH adh0 GND efet w=14 l=8
+ ad=0 pd=0 as=0 ps=0 
M4475 GND npchp0 pchp0 GND efet w=42 l=7
+ ad=0 pd=0 as=0 ps=0 
M4476 n_856 dpc34_PCLC n_919 GND efet w=45 l=7
+ ad=473 pd=122 as=521 ps=146 
M4477 GND n_311 n_856 GND efet w=44 l=6
+ ad=0 pd=0 as=0 ps=0 
M4478 n_1010 pch0 GND GND efet w=39 l=6
+ ad=417 pd=118 as=0 ps=0 
M4479 Vdd n_1010 n_1010 GND dfet w=10 l=20
+ ad=0 pd=0 as=1107 ps=344 
M4480 pchp0 dpc33_PCHDB idb0 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M4481 adh0 dpc32_PCHADH pchp0 GND efet w=14 l=8
+ ad=0 pd=0 as=0 ps=0 
M4482 adl1 cclk Vdd GND efet w=22 l=7
+ ad=0 pd=0 as=0 ps=0 
M4483 pchp1 dpc31_PCHPCH pch1 GND efet w=14 l=8
+ ad=1705 pd=426 as=592 ps=158 
M4484 pch1 dpc30_ADHPCH adh1 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M4485 n_1618 dpc26_ACDB idb2 GND efet w=14 l=8
+ ad=0 pd=0 as=0 ps=0 
M4486 idb2 dpc25_SBDB sb2 GND efet w=22 l=5
+ ad=0 pd=0 as=0 ps=0 
M4487 sb2 dpc24_ACSB n_1618 GND efet w=15 l=8
+ ad=0 pd=0 as=0 ps=0 
M4488 Vdd n_419 n_419 GND dfet w=10 l=16
+ ad=0 pd=0 as=1003 ps=282 
M4489 a3 dpc23_SBAC dasb3 GND efet w=11 l=7
+ ad=457 pd=136 as=0 ps=0 
M4490 Vdd n_1654 n_1654 GND dfet w=10 l=13
+ ad=0 pd=0 as=318 ps=98 
M4491 GND n_1097 dasb3 GND efet w=25 l=6
+ ad=0 pd=0 as=0 ps=0 
M4492 n_1279 n_986 n_345 GND efet w=39 l=6
+ ad=234 pd=90 as=0 ps=0 
M4493 GND n_600 n_1279 GND efet w=39 l=6
+ ad=0 pd=0 as=0 ps=0 
M4494 n_1097 n_432 GND GND efet w=31 l=6
+ ad=559 pd=180 as=0 ps=0 
M4495 n_1179 n_1179 Vdd GND dfet w=9 l=15
+ ad=714 pd=202 as=0 ps=0 
M4496 n_8 n_551 GND GND efet w=37 l=6
+ ad=448 pd=124 as=0 ps=0 
M4497 GND n_345 n_1097 GND efet w=32 l=6
+ ad=0 pd=0 as=0 ps=0 
M4498 n_345 n_345 Vdd GND dfet w=10 l=16
+ ad=942 pd=290 as=0 ps=0 
M4499 n_432 sb3 GND GND efet w=13 l=7
+ ad=858 pd=242 as=0 ps=0 
M4500 n_8 n_8 Vdd GND dfet w=10 l=10
+ ad=4195 pd=1410 as=0 ps=0 
M4501 n_1097 n_1097 Vdd GND dfet w=9 l=16
+ ad=1021 pd=306 as=0 ps=0 
M4502 n_1179 cclk n_393 GND efet w=11 l=8
+ ad=0 pd=0 as=115 ps=54 
M4503 Vdd n_306 n_306 GND dfet w=10 l=16
+ ad=0 pd=0 as=476 ps=124 
M4504 n_306 cclk n_581 GND efet w=12 l=8
+ ad=745 pd=232 as=177 ps=70 
M4505 GND dpc22_nDSA n_306 GND efet w=36 l=6
+ ad=0 pd=0 as=0 ps=0 
M4506 n_432 sb3 GND GND efet w=34 l=7
+ ad=0 pd=0 as=0 ps=0 
M4507 Vdd n_432 n_432 GND dfet w=9 l=16
+ ad=0 pd=0 as=1180 ps=360 
M4508 n_1654 cclk a3 GND efet w=12 l=7
+ ad=1661 pd=384 as=0 ps=0 
M4509 n_1654 n_947 GND GND efet w=81 l=6
+ ad=0 pd=0 as=0 ps=0 
M4510 GND a3 n_947 GND efet w=44 l=7
+ ad=0 pd=0 as=767 ps=204 
M4511 adh2 dpc27_SBADH sb2 GND efet w=22 l=8
+ ad=1772 pd=456 as=0 ps=0 
M4512 GND dpc29_0ADH17 adh2 GND efet w=22 l=7
+ ad=0 pd=0 as=0 ps=0 
M4513 n_1654 dpc26_ACDB idb3 GND efet w=14 l=8
+ ad=0 pd=0 as=0 ps=0 
M4514 idb3 dpc25_SBDB sb3 GND efet w=22 l=6
+ ad=0 pd=0 as=0 ps=0 
M4515 sb3 dpc24_ACSB n_1654 GND efet w=14 l=9
+ ad=0 pd=0 as=0 ps=0 
M4516 Vdd n_947 n_947 GND dfet w=10 l=16
+ ad=0 pd=0 as=971 ps=282 
M4517 GND alucout n_811 GND efet w=41 l=6
+ ad=0 pd=0 as=929 ps=222 
M4518 n_753 n_811 GND GND efet w=12 l=6
+ ad=1080 pd=282 as=0 ps=0 
M4519 a4 dpc23_SBAC sb4 GND efet w=12 l=7
+ ad=423 pd=134 as=0 ps=0 
M4520 n_551 n_393 GND GND efet w=44 l=7
+ ad=577 pd=182 as=0 ps=0 
M4521 GND n_581 n_838 GND efet w=45 l=6
+ ad=0 pd=0 as=671 ps=178 
M4522 n_811 n_838 GND GND efet w=49 l=7
+ ad=0 pd=0 as=0 ps=0 
M4523 n_753 n_811 GND GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M4524 n_753 n_1257 GND GND efet w=31 l=6
+ ad=0 pd=0 as=0 ps=0 
M4525 n_551 n_551 Vdd GND dfet w=9 l=15
+ ad=1586 pd=526 as=0 ps=0 
M4526 n_838 n_838 Vdd GND dfet w=10 l=17
+ ad=873 pd=242 as=0 ps=0 
M4527 n_811 n_811 Vdd GND dfet w=9 l=9
+ ad=3739 pd=1334 as=0 ps=0 
M4528 Vdd n_761 n_761 GND dfet w=8 l=16
+ ad=0 pd=0 as=3156 ps=1014 
M4529 GND alu5 n_761 GND efet w=37 l=8
+ ad=0 pd=0 as=669 ps=184 
M4530 Vdd n_233 n_233 GND dfet w=9 l=16
+ ad=0 pd=0 as=3064 ps=1048 
M4531 n_233 n_761 n_970 GND efet w=45 l=6
+ ad=730 pd=214 as=405 ps=114 
M4532 n_970 n_149 GND GND efet w=38 l=6
+ ad=0 pd=0 as=0 ps=0 
M4533 n_753 n_753 Vdd GND dfet w=9 l=16
+ ad=1219 pd=370 as=0 ps=0 
M4534 n_762 n_149 GND GND efet w=36 l=6
+ ad=664 pd=190 as=0 ps=0 
M4535 GND n_761 n_762 GND efet w=36 l=7
+ ad=0 pd=0 as=0 ps=0 
M4536 adl7 dpc21_ADDADL alu7 GND efet w=16 l=8
+ ad=0 pd=0 as=1243 ps=346 
M4537 GND notalu7 alu7 GND efet w=101 l=7
+ ad=0 pd=0 as=0 ps=0 
M4538 Vdd notaluvout notaluvout GND dfet w=10 l=16
+ ad=0 pd=0 as=667 ps=226 
M4539 GND n_1315 n_826 GND efet w=114 l=8
+ ad=0 pd=0 as=1817 ps=394 
M4540 GND n_617 n_1140 GND efet w=114 l=6
+ ad=0 pd=0 as=1870 ps=400 
M4541 Vdd abh0 abh0 GND dfet w=9 l=15
+ ad=0 pd=0 as=2571 ps=784 
M4542 GND n_171 ab7 GND efet w=116 l=36
+ ad=0 pd=0 as=19404 ps=2768 
M4543 n_1668 cp1 n_705 GND efet w=11 l=9
+ ad=0 pd=0 as=66 ps=34 
M4544 n_705 ADH_ABH nABH0 GND efet w=11 l=8
+ ad=0 pd=0 as=380 ps=120 
M4545 GND n_171 ab7 GND efet w=212 l=6
+ ad=0 pd=0 as=0 ps=0 
M4546 ab7 n_171 GND GND efet w=212 l=6
+ ad=0 pd=0 as=0 ps=0 
M4547 ab7 n_171 GND GND efet w=437 l=6
+ ad=0 pd=0 as=0 ps=0 
M4548 n_826 abh0 Vdd GND dfet w=18 l=7
+ ad=0 pd=0 as=0 ps=0 
M4549 Vdd n_1315 n_1315 GND dfet w=9 l=10
+ ad=0 pd=0 as=2052 ps=612 
M4550 Vdd n_322 ab7 GND efet w=256 l=6
+ ad=0 pd=0 as=0 ps=0 
M4551 nABH0 cclk n_381 GND efet w=11 l=7
+ ad=0 pd=0 as=1283 ps=378 
M4552 Vdd n_1315 n_381 GND dfet w=21 l=8
+ ad=0 pd=0 as=0 ps=0 
M4553 GND abh0 n_1315 GND efet w=36 l=7
+ ad=0 pd=0 as=459 ps=130 
M4554 GND abh0 n_381 GND efet w=155 l=7
+ ad=0 pd=0 as=0 ps=0 
M4555 GND n_381 ab8 GND efet w=14 l=6
+ ad=0 pd=0 as=18277 ps=2308 
M4556 GND n_381 ab8 GND efet w=42 l=6
+ ad=0 pd=0 as=0 ps=0 
M4557 Vdd n_322 ab7 GND efet w=264 l=7
+ ad=0 pd=0 as=0 ps=0 
M4558 Vdd n_322 ab7 GND efet w=235 l=7
+ ad=0 pd=0 as=0 ps=0 
M4559 Vdd n_322 ab7 GND efet w=233 l=6
+ ad=0 pd=0 as=0 ps=0 
M4560 ab8 n_381 GND GND efet w=163 l=6
+ ad=0 pd=0 as=0 ps=0 
M4561 GND n_381 ab8 GND efet w=163 l=7
+ ad=0 pd=0 as=0 ps=0 
M4562 ab8 n_381 GND GND efet w=163 l=7
+ ad=0 pd=0 as=0 ps=0 
M4563 GND n_381 ab8 GND efet w=163 l=7
+ ad=0 pd=0 as=0 ps=0 
M4564 ab8 n_381 GND GND efet w=163 l=6
+ ad=0 pd=0 as=0 ps=0 
M4565 Vdd n_826 ab8 GND efet w=414 l=6
+ ad=0 pd=0 as=0 ps=0 
M4566 Vdd n_826 ab8 GND efet w=317 l=6
+ ad=0 pd=0 as=0 ps=0 
M4567 Vdd n_826 ab8 GND efet w=159 l=7
+ ad=0 pd=0 as=0 ps=0 
M4568 ab9 n_1140 Vdd GND efet w=159 l=6
+ ad=18412 pd=2314 as=0 ps=0 
M4569 Vdd n_1140 ab9 GND efet w=317 l=7
+ ad=0 pd=0 as=0 ps=0 
M4570 Vdd n_1140 ab9 GND efet w=416 l=6
+ ad=0 pd=0 as=0 ps=0 
M4571 Vdd abh1 n_1140 GND dfet w=18 l=8
+ ad=0 pd=0 as=0 ps=0 
M4572 n_617 abh1 GND GND efet w=45 l=7
+ ad=445 pd=144 as=0 ps=0 
M4573 Vdd n_617 n_617 GND dfet w=10 l=10
+ ad=0 pd=0 as=2008 ps=680 
M4574 abh1 abh1 Vdd GND dfet w=9 l=14
+ ad=2441 pd=662 as=0 ps=0 
M4575 GND nABH1 abh1 GND efet w=65 l=7
+ ad=0 pd=0 as=602 ps=186 
M4576 n_637 n_637 Vdd GND dfet w=9 l=15
+ ad=1300 pd=448 as=0 ps=0 
M4577 GND n_637 notaluvout GND efet w=30 l=6
+ ad=0 pd=0 as=0 ps=0 
M4578 alu7 dpc19_ADDSB7 sb7 GND efet w=20 l=7
+ ad=0 pd=0 as=0 ps=0 
M4579 DC78_phi2 cclk DC78 GND efet w=12 l=8
+ ad=162 pd=72 as=0 ps=0 
M4580 C78_phi2 cclk C78 GND efet w=11 l=8
+ ad=145 pd=70 as=1078 ps=296 
M4581 alu7 alu7 Vdd GND dfet w=10 l=13
+ ad=355 pd=104 as=0 ps=0 
M4582 n_762 n_762 Vdd GND dfet w=9 l=16
+ ad=2300 pd=738 as=0 ps=0 
M4583 Vdd n_149 n_149 GND dfet w=9 l=17
+ ad=0 pd=0 as=1009 ps=310 
M4584 GND alu6 n_149 GND efet w=49 l=6
+ ad=0 pd=0 as=837 ps=234 
M4585 C78 nC78 GND GND efet w=59 l=6
+ ad=0 pd=0 as=0 ps=0 
M4586 n_408 cclk notaluvout GND efet w=11 l=7
+ ad=211 pd=86 as=0 ps=0 
M4587 GND n_408 aluvout GND efet w=130 l=7
+ ad=0 pd=0 as=1644 ps=394 
M4588 n_1203 n_1135 GND GND efet w=46 l=6
+ ad=286 pd=104 as=0 ps=0 
M4589 Vdd dasb5 dasb5 GND dfet w=9 l=17
+ ad=0 pd=0 as=393 ps=102 
M4590 Vdd n_1344 n_1344 GND dfet w=10 l=13
+ ad=0 pd=0 as=346 ps=100 
M4591 n_1344 cclk a4 GND efet w=11 l=8
+ ad=1499 pd=386 as=0 ps=0 
M4592 n_1344 n_556 GND GND efet w=82 l=7
+ ad=0 pd=0 as=0 ps=0 
M4593 GND a4 n_556 GND efet w=43 l=6
+ ad=0 pd=0 as=755 ps=204 
M4594 Vdd cclk adh2 GND efet w=22 l=7
+ ad=0 pd=0 as=0 ps=0 
M4595 adh3 dpc27_SBADH sb3 GND efet w=21 l=7
+ ad=1987 pd=498 as=0 ps=0 
M4596 GND dpc29_0ADH17 adh3 GND efet w=21 l=8
+ ad=0 pd=0 as=0 ps=0 
M4597 n_1344 dpc26_ACDB idb4 GND efet w=14 l=8
+ ad=0 pd=0 as=0 ps=0 
M4598 idb4 dpc25_SBDB sb4 GND efet w=22 l=5
+ ad=0 pd=0 as=0 ps=0 
M4599 sb4 dpc24_ACSB n_1344 GND efet w=14 l=8
+ ad=0 pd=0 as=0 ps=0 
M4600 Vdd n_556 n_556 GND dfet w=9 l=16
+ ad=0 pd=0 as=1032 ps=284 
M4601 dasb5 n_753 n_1203 GND efet w=34 l=6
+ ad=659 pd=184 as=0 ps=0 
M4602 a5 dpc23_SBAC dasb5 GND efet w=11 l=7
+ ad=475 pd=140 as=0 ps=0 
M4603 Vdd n_831 n_831 GND dfet w=9 l=13
+ ad=0 pd=0 as=318 ps=98 
M4604 GND n_1629 dasb5 GND efet w=18 l=7
+ ad=0 pd=0 as=0 ps=0 
M4605 GND sb5 n_1135 GND efet w=62 l=7
+ ad=0 pd=0 as=1308 ps=360 
M4606 n_1629 n_1135 GND GND efet w=18 l=6
+ ad=587 pd=164 as=0 ps=0 
M4607 GND n_753 n_1629 GND efet w=26 l=7
+ ad=0 pd=0 as=0 ps=0 
M4608 Vdd n_1056 n_1056 GND dfet w=10 l=16
+ ad=0 pd=0 as=972 ps=298 
M4609 GND n_761 n_1056 GND efet w=29 l=7
+ ad=0 pd=0 as=379 ps=124 
M4610 n_1629 n_1629 Vdd GND dfet w=10 l=17
+ ad=958 pd=270 as=0 ps=0 
M4611 Vdd n_1135 n_1135 GND dfet w=9 l=14
+ ad=0 pd=0 as=1127 ps=340 
M4612 Vdd dasb6 dasb6 GND dfet w=9 l=17
+ ad=0 pd=0 as=358 ps=104 
M4613 n_1554 n_61 GND GND efet w=36 l=6
+ ad=216 pd=84 as=0 ps=0 
M4614 dasb6 n_739 n_1554 GND efet w=36 l=7
+ ad=673 pd=190 as=0 ps=0 
M4615 n_831 cclk a5 GND efet w=12 l=8
+ ad=1536 pd=384 as=0 ps=0 
M4616 n_831 n_1719 GND GND efet w=80 l=6
+ ad=0 pd=0 as=0 ps=0 
M4617 GND a5 n_1719 GND efet w=44 l=7
+ ad=0 pd=0 as=679 ps=202 
M4618 adh4 dpc27_SBADH sb4 GND efet w=22 l=7
+ ad=1644 pd=404 as=0 ps=0 
M4619 GND dpc29_0ADH17 adh4 GND efet w=22 l=8
+ ad=0 pd=0 as=0 ps=0 
M4620 n_831 dpc26_ACDB idb5 GND efet w=14 l=8
+ ad=0 pd=0 as=0 ps=0 
M4621 idb5 dpc25_SBDB sb5 GND efet w=21 l=7
+ ad=0 pd=0 as=0 ps=0 
M4622 sb5 dpc24_ACSB n_831 GND efet w=14 l=8
+ ad=0 pd=0 as=0 ps=0 
M4623 Vdd n_1719 n_1719 GND dfet w=9 l=16
+ ad=0 pd=0 as=1042 ps=284 
M4624 a6 dpc23_SBAC dasb6 GND efet w=12 l=7
+ ad=462 pd=140 as=0 ps=0 
M4625 Vdd n_326 n_326 GND dfet w=10 l=13
+ ad=0 pd=0 as=331 ps=100 
M4626 n_1080 n_811 GND GND efet w=35 l=7
+ ad=175 pd=80 as=0 ps=0 
M4627 n_739 n_1056 n_1080 GND efet w=35 l=6
+ ad=918 pd=236 as=0 ps=0 
M4628 GND n_479 dasb6 GND efet w=18 l=7
+ ad=0 pd=0 as=0 ps=0 
M4629 n_479 n_61 GND GND efet w=20 l=6
+ ad=636 pd=170 as=0 ps=0 
M4630 GND n_739 n_479 GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M4631 n_711 n_761 n_739 GND efet w=34 l=6
+ ad=204 pd=80 as=0 ps=0 
M4632 GND n_1257 n_711 GND efet w=34 l=6
+ ad=0 pd=0 as=0 ps=0 
M4633 Vdd n_61 n_61 GND dfet w=10 l=17
+ ad=0 pd=0 as=867 ps=270 
M4634 n_739 n_739 Vdd GND dfet w=9 l=17
+ ad=1054 pd=314 as=0 ps=0 
M4635 n_61 sb6 GND GND efet w=50 l=6
+ ad=583 pd=174 as=0 ps=0 
M4636 n_479 n_479 Vdd GND dfet w=10 l=17
+ ad=980 pd=276 as=0 ps=0 
M4637 Vdd dasb7 dasb7 GND dfet w=10 l=16
+ ad=0 pd=0 as=355 ps=104 
M4638 GND n_762 n_1018 GND efet w=42 l=7
+ ad=0 pd=0 as=588 ps=168 
M4639 n_100 n_1018 GND GND efet w=47 l=6
+ ad=290 pd=108 as=0 ps=0 
M4640 n_1205 n_811 n_100 GND efet w=48 l=6
+ ad=868 pd=236 as=0 ps=0 
M4641 n_1454 n_852 GND GND efet w=36 l=7
+ ad=216 pd=84 as=0 ps=0 
M4642 dasb7 n_1205 n_1454 GND efet w=36 l=7
+ ad=701 pd=180 as=0 ps=0 
M4643 n_326 cclk a6 GND efet w=12 l=8
+ ad=1516 pd=388 as=0 ps=0 
M4644 n_326 n_1356 GND GND efet w=82 l=6
+ ad=0 pd=0 as=0 ps=0 
M4645 GND a6 n_1356 GND efet w=44 l=7
+ ad=0 pd=0 as=721 ps=198 
M4646 adh5 dpc27_SBADH sb5 GND efet w=22 l=7
+ ad=1667 pd=430 as=0 ps=0 
M4647 GND dpc29_0ADH17 adh5 GND efet w=22 l=8
+ ad=0 pd=0 as=0 ps=0 
M4648 n_326 dpc26_ACDB idb6 GND efet w=14 l=8
+ ad=0 pd=0 as=0 ps=0 
M4649 idb6 dpc25_SBDB sb6 GND efet w=22 l=7
+ ad=0 pd=0 as=0 ps=0 
M4650 sb6 dpc24_ACSB n_326 GND efet w=13 l=8
+ ad=0 pd=0 as=0 ps=0 
M4651 Vdd n_1356 n_1356 GND dfet w=8 l=17
+ ad=0 pd=0 as=1016 ps=284 
M4652 a7 dpc23_SBAC dasb7 GND efet w=12 l=8
+ ad=433 pd=136 as=0 ps=0 
M4653 GND n_260 dasb7 GND efet w=18 l=6
+ ad=0 pd=0 as=0 ps=0 
M4654 n_260 n_852 GND GND efet w=19 l=7
+ ad=612 pd=170 as=0 ps=0 
M4655 GND n_1205 n_260 GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M4656 n_1018 n_1018 Vdd GND dfet w=9 l=10
+ ad=756 pd=238 as=0 ps=0 
M4657 n_569 n_233 n_1205 GND efet w=36 l=7
+ ad=180 pd=82 as=0 ps=0 
M4658 GND n_1257 n_569 GND efet w=36 l=6
+ ad=0 pd=0 as=0 ps=0 
M4659 n_852 sb7 GND GND efet w=28 l=6
+ ad=525 pd=152 as=0 ps=0 
M4660 Vdd n_852 n_852 GND dfet w=10 l=16
+ ad=0 pd=0 as=962 ps=276 
M4661 n_1205 n_1205 Vdd GND dfet w=9 l=17
+ ad=1050 pd=294 as=0 ps=0 
M4662 n_852 sb7 GND GND efet w=19 l=6
+ ad=0 pd=0 as=0 ps=0 
M4663 n_260 n_260 Vdd GND dfet w=9 l=17
+ ad=1047 pd=278 as=0 ps=0 
M4664 Vdd n_1592 n_1592 GND dfet w=10 l=14
+ ad=0 pd=0 as=364 ps=100 
M4665 n_1592 cclk a7 GND efet w=11 l=7
+ ad=1433 pd=372 as=0 ps=0 
M4666 n_1592 n_128 GND GND efet w=77 l=6
+ ad=0 pd=0 as=0 ps=0 
M4667 GND a7 n_128 GND efet w=45 l=6
+ ad=0 pd=0 as=736 ps=204 
M4668 adh6 dpc27_SBADH sb6 GND efet w=22 l=8
+ ad=1781 pd=428 as=0 ps=0 
M4669 GND dpc29_0ADH17 adh6 GND efet w=22 l=9
+ ad=0 pd=0 as=0 ps=0 
M4670 pchp0 pchp0 Vdd GND dfet w=10 l=18
+ ad=479 pd=126 as=0 ps=0 
M4671 n_835 n_919 n_1229 GND efet w=58 l=6
+ ad=1312 pd=346 as=0 ps=0 
M4672 n_311 n_1010 GND GND efet w=22 l=6
+ ad=1156 pd=270 as=0 ps=0 
M4673 n_835 dpc34_PCLC GND GND efet w=55 l=6
+ ad=0 pd=0 as=0 ps=0 
M4674 n_1229 n_1229 Vdd GND dfet w=10 l=17
+ ad=394 pd=112 as=0 ps=0 
M4675 GND n_311 n_835 GND efet w=54 l=6
+ ad=0 pd=0 as=0 ps=0 
M4676 dpc35_PCHC n_1010 GND GND efet w=56 l=6
+ ad=0 pd=0 as=0 ps=0 
M4677 Vdd pchp1 pchp1 GND dfet w=9 l=16
+ ad=0 pd=0 as=435 ps=126 
M4678 Vdd npchp1 npchp1 GND dfet w=10 l=16
+ ad=0 pd=0 as=1052 ps=326 
M4679 Vdd n_1486 n_1486 GND dfet w=9 l=17
+ ad=0 pd=0 as=332 ps=86 
M4680 n_1486 cclk n_126 GND efet w=11 l=7
+ ad=874 pd=228 as=166 ps=62 
M4681 GND npchp1 pchp1 GND efet w=61 l=6
+ ad=0 pd=0 as=0 ps=0 
M4682 pchp1 dpc33_PCHDB idb1 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M4683 n_1070 pch1 GND GND efet w=34 l=6
+ ad=750 pd=198 as=0 ps=0 
M4684 GND n_126 npchp1 GND efet w=42 l=6
+ ad=0 pd=0 as=849 ps=246 
M4685 n_1486 n_200 GND GND efet w=33 l=6
+ ad=0 pd=0 as=0 ps=0 
M4686 n_1538 n_919 n_1486 GND efet w=43 l=6
+ ad=258 pd=98 as=0 ps=0 
M4687 GND n_1070 n_1538 GND efet w=43 l=6
+ ad=0 pd=0 as=0 ps=0 
M4688 dpc35_PCHC n_1070 GND GND efet w=57 l=7
+ ad=0 pd=0 as=0 ps=0 
M4689 n_200 n_1070 GND GND efet w=24 l=7
+ ad=1128 pd=294 as=0 ps=0 
M4690 GND n_919 n_200 GND efet w=22 l=6
+ ad=0 pd=0 as=0 ps=0 
M4691 adh1 dpc32_PCHADH pchp1 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M4692 n_1070 n_1070 Vdd GND dfet w=10 l=21
+ ad=1643 pd=480 as=0 ps=0 
M4693 n_200 n_200 Vdd GND dfet w=9 l=14
+ ad=2067 pd=638 as=0 ps=0 
M4694 n_1202 n_1202 Vdd GND dfet w=10 l=17
+ ad=1271 pd=408 as=0 ps=0 
M4695 GND n_1157 dpc41_DL_ADL GND efet w=96 l=7
+ ad=0 pd=0 as=0 ps=0 
M4696 dpc42_DL_ADH n_1441 GND GND efet w=98 l=6
+ ad=0 pd=0 as=0 ps=0 
M4697 dpc43_DL_DB n_1240 GND GND efet w=103 l=6
+ ad=958 pd=244 as=0 ps=0 
M4698 Vdd n_1566 dpc43_DL_DB GND dfet w=9 l=9
+ ad=0 pd=0 as=0 ps=0 
M4699 DBZ idb2 GND GND efet w=54 l=6
+ ad=2373 pd=588 as=0 ps=0 
M4700 GND idb7 DBZ GND efet w=68 l=6
+ ad=0 pd=0 as=0 ps=0 
M4701 DBZ idb6 GND GND efet w=51 l=6
+ ad=0 pd=0 as=0 ps=0 
M4702 GND idb3 DBZ GND efet w=38 l=5
+ ad=0 pd=0 as=0 ps=0 
M4703 Vdd n_206 n_206 GND dfet w=14 l=7
+ ad=0 pd=0 as=5645 ps=1900 
M4704 Pout0 Pout0 Vdd GND dfet w=9 l=10
+ ad=615 pd=218 as=0 ps=0 
M4705 Pout1 Pout1 Vdd GND dfet w=10 l=10
+ ad=265 pd=86 as=0 ps=0 
M4706 Pout0 H1x1 idb0 GND efet w=24 l=8
+ ad=0 pd=0 as=0 ps=0 
M4707 Pout1 H1x1 idb1 GND efet w=25 l=8
+ ad=0 pd=0 as=0 ps=0 
M4708 GND idb0 n_1224 GND efet w=71 l=6
+ ad=0 pd=0 as=827 ps=216 
M4709 n_243 idb1 GND GND efet w=71 l=6
+ ad=760 pd=224 as=0 ps=0 
M4710 n_1391 cclk pipeUNK15 GND efet w=12 l=9
+ ad=0 pd=0 as=159 ps=66 
M4711 GND pipeUNK15 H1x1 GND efet w=83 l=5
+ ad=0 pd=0 as=1174 ps=256 
M4712 Vdd n_307 n_307 GND dfet w=9 l=11
+ ad=0 pd=0 as=1254 ps=438 
M4713 n_90 n_90 Vdd GND dfet w=10 l=11
+ ad=2476 pd=844 as=0 ps=0 
M4714 GND n_90 n_1433 GND efet w=41 l=6
+ ad=0 pd=0 as=1123 ps=340 
M4715 GND n_620 n_922 GND efet w=81 l=7
+ ad=0 pd=0 as=405 ps=172 
M4716 n_922 n_270 BRtaken GND efet w=81 l=6
+ ad=0 pd=0 as=1068 ps=260 
M4717 BRtaken BRtaken Vdd GND dfet w=9 l=9
+ ad=4602 pd=1580 as=0 ps=0 
M4718 GND n_1115 BRtaken GND efet w=51 l=7
+ ad=0 pd=0 as=0 ps=0 
M4719 n_1433 nop_branch_bit6 GND GND efet w=41 l=7
+ ad=0 pd=0 as=0 ps=0 
M4720 n_1170 n_755 GND GND efet w=25 l=7
+ ad=713 pd=176 as=0 ps=0 
M4721 GND n_781 n_1170 GND efet w=26 l=7
+ ad=0 pd=0 as=0 ps=0 
M4722 n_1170 n_1170 Vdd GND dfet w=10 l=15
+ ad=780 pd=236 as=0 ps=0 
M4723 n_580 nDBZ GND GND efet w=49 l=6
+ ad=405 pd=136 as=0 ps=0 
M4724 n_1224 n_1224 Vdd GND dfet w=10 l=12
+ ad=2917 pd=928 as=0 ps=0 
M4725 GND n_937 dpc34_PCLC GND efet w=48 l=6
+ ad=0 pd=0 as=0 ps=0 
M4726 n_1706 n_937 GND GND efet w=40 l=7
+ ad=200 pd=90 as=0 ps=0 
M4727 n_1500 dpc36_nIPC n_1706 GND efet w=40 l=6
+ ad=916 pd=220 as=0 ps=0 
M4728 Vdd n_1500 n_1500 GND dfet w=10 l=16
+ ad=0 pd=0 as=319 ps=82 
M4729 Vdd npclp0 npclp0 GND dfet w=10 l=21
+ ad=0 pd=0 as=1132 ps=344 
M4730 n_526 cclk n_1500 GND efet w=12 l=9
+ ad=167 pd=74 as=0 ps=0 
M4731 GND n_937 n_1345 GND efet w=24 l=6
+ ad=0 pd=0 as=1155 ps=318 
M4732 GND n_1345 n_1500 GND efet w=33 l=6
+ ad=0 pd=0 as=0 ps=0 
M4733 Vdd pclp0 pclp0 GND dfet w=10 l=15
+ ad=0 pd=0 as=418 ps=124 
M4734 n_1345 dpc36_nIPC GND GND efet w=22 l=6
+ ad=0 pd=0 as=0 ps=0 
M4735 npclp0 n_526 GND GND efet w=35 l=7
+ ad=745 pd=228 as=0 ps=0 
M4736 GND pcl0 n_937 GND efet w=34 l=7
+ ad=0 pd=0 as=730 ps=186 
M4737 pclp0 npclp0 GND GND efet w=61 l=6
+ ad=1631 pd=392 as=0 ps=0 
M4738 Vdd cclk adl2 GND efet w=22 l=6
+ ad=0 pd=0 as=0 ps=0 
M4739 Vdd n_293 n_293 GND dfet w=11 l=15
+ ad=0 pd=0 as=2168 ps=692 
M4740 n_1402 cclk npchp2 GND efet w=11 l=8
+ ad=806 pd=232 as=217 ps=80 
M4741 pchp2 dpc31_PCHPCH pch2 GND efet w=15 l=7
+ ad=1589 pd=390 as=611 ps=158 
M4742 pch2 dpc30_ADHPCH adh2 GND efet w=14 l=8
+ ad=0 pd=0 as=0 ps=0 
M4743 n_1592 dpc26_ACDB idb7 GND efet w=14 l=8
+ ad=0 pd=0 as=0 ps=0 
M4744 idb7 dpc25_SBDB sb7 GND efet w=21 l=7
+ ad=0 pd=0 as=0 ps=0 
M4745 sb7 dpc24_ACSB n_1592 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M4746 Vdd n_128 n_128 GND dfet w=10 l=16
+ ad=0 pd=0 as=1062 ps=284 
M4747 adh7 dpc27_SBADH sb7 GND efet w=22 l=8
+ ad=1928 pd=478 as=0 ps=0 
M4748 GND dpc29_0ADH17 adh7 GND efet w=22 l=8
+ ad=0 pd=0 as=0 ps=0 
M4749 GND npchp2 pchp2 GND efet w=43 l=6
+ ad=0 pd=0 as=0 ps=0 
M4750 n_1367 n_200 n_293 GND efet w=43 l=7
+ ad=431 pd=120 as=501 ps=144 
M4751 GND n_1202 n_1367 GND efet w=45 l=6
+ ad=0 pd=0 as=0 ps=0 
M4752 n_1265 pch2 GND GND efet w=44 l=7
+ ad=462 pd=126 as=0 ps=0 
M4753 Vdd n_1265 n_1265 GND dfet w=9 l=20
+ ad=0 pd=0 as=1099 ps=342 
M4754 pchp2 dpc33_PCHDB idb2 GND efet w=15 l=7
+ ad=0 pd=0 as=0 ps=0 
M4755 n_57 n_293 n_1402 GND efet w=57 l=6
+ ad=1242 pd=338 as=0 ps=0 
M4756 n_1202 n_1265 GND GND efet w=23 l=6
+ ad=1206 pd=272 as=0 ps=0 
M4757 Vdd n_1166 n_1166 GND dfet w=10 l=16
+ ad=0 pd=0 as=1363 ps=414 
M4758 n_1345 n_1345 Vdd GND dfet w=10 l=14
+ ad=1974 pd=630 as=0 ps=0 
M4759 n_937 n_937 Vdd GND dfet w=10 l=20
+ ad=1493 pd=434 as=0 ps=0 
M4760 adl0 dpc38_PCLADL pclp0 GND efet w=14 l=8
+ ad=0 pd=0 as=0 ps=0 
M4761 adl0 dpc40_ADLPCL pcl0 GND efet w=14 l=8
+ ad=0 pd=0 as=476 ps=96 
M4762 pcl0 dpc39_PCLPCL pclp0 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M4763 idb0 dpc37_PCLDB pclp0 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M4764 Vdd n_329 n_329 GND dfet w=10 l=20
+ ad=0 pd=0 as=1280 ps=344 
M4765 GND pcl1 n_329 GND efet w=41 l=6
+ ad=0 pd=0 as=401 ps=122 
M4766 GND n_329 n_1166 GND efet w=23 l=7
+ ad=0 pd=0 as=1137 ps=270 
M4767 n_1685 n_1166 GND GND efet w=43 l=7
+ ad=464 pd=120 as=0 ps=0 
M4768 Vdd n_1542 n_1542 GND dfet w=10 l=13
+ ad=0 pd=0 as=2181 ps=694 
M4769 n_1542 n_1345 n_1685 GND efet w=45 l=6
+ ad=603 pd=146 as=0 ps=0 
M4770 npclp1 cclk n_1099 GND efet w=11 l=8
+ ad=227 pd=92 as=1133 ps=292 
M4771 adl1 dpc38_PCLADL pclp1 GND efet w=14 l=7
+ ad=0 pd=0 as=1536 ps=352 
M4772 GND n_329 dpc34_PCLC GND efet w=55 l=7
+ ad=0 pd=0 as=0 ps=0 
M4773 n_1568 n_1166 GND GND efet w=56 l=7
+ ad=1215 pd=334 as=0 ps=0 
M4774 GND n_1345 n_1568 GND efet w=53 l=7
+ ad=0 pd=0 as=0 ps=0 
M4775 n_1099 n_1542 n_1568 GND efet w=58 l=6
+ ad=0 pd=0 as=0 ps=0 
M4776 pclp1 npclp1 GND GND efet w=57 l=6
+ ad=0 pd=0 as=0 ps=0 
M4777 adl1 dpc40_ADLPCL pcl1 GND efet w=14 l=9
+ ad=0 pd=0 as=462 ps=94 
M4778 pcl1 dpc39_PCLPCL pclp1 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M4779 n_1099 n_1099 Vdd GND dfet w=10 l=16
+ ad=394 pd=112 as=0 ps=0 
M4780 idb1 dpc37_PCLDB pclp1 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M4781 adh2 dpc32_PCHADH pchp2 GND efet w=14 l=8
+ ad=0 pd=0 as=0 ps=0 
M4782 adl3 cclk Vdd GND efet w=23 l=7
+ ad=0 pd=0 as=0 ps=0 
M4783 pchp3 dpc31_PCHPCH pch3 GND efet w=14 l=8
+ ad=1661 pd=418 as=596 ps=156 
M4784 pch3 dpc30_ADHPCH adh3 GND efet w=14 l=8
+ ad=0 pd=0 as=0 ps=0 
M4785 dpc23_SBAC cclk GND GND efet w=26 l=7
+ ad=0 pd=0 as=0 ps=0 
M4786 dpc24_ACSB cclk GND GND efet w=26 l=7
+ ad=0 pd=0 as=0 ps=0 
M4787 dpc26_ACDB cclk GND GND efet w=27 l=7
+ ad=0 pd=0 as=0 ps=0 
M4788 pchp2 pchp2 Vdd GND dfet w=9 l=19
+ ad=476 pd=124 as=0 ps=0 
M4789 n_57 n_200 GND GND efet w=54 l=6
+ ad=0 pd=0 as=0 ps=0 
M4790 n_1402 n_1402 Vdd GND dfet w=10 l=17
+ ad=383 pd=112 as=0 ps=0 
M4791 GND n_1202 n_57 GND efet w=55 l=6
+ ad=0 pd=0 as=0 ps=0 
M4792 dpc35_PCHC n_1265 GND GND efet w=54 l=6
+ ad=0 pd=0 as=0 ps=0 
M4793 Vdd pchp3 pchp3 GND dfet w=10 l=16
+ ad=0 pd=0 as=446 ps=124 
M4794 Vdd npchp3 npchp3 GND dfet w=10 l=16
+ ad=0 pd=0 as=1102 ps=326 
M4795 Vdd n_207 n_207 GND dfet w=9 l=16
+ ad=0 pd=0 as=306 ps=84 
M4796 n_207 cclk n_1061 GND efet w=11 l=8
+ ad=922 pd=242 as=142 ps=74 
M4797 GND npchp3 pchp3 GND efet w=59 l=6
+ ad=0 pd=0 as=0 ps=0 
M4798 pchp3 dpc33_PCHDB idb3 GND efet w=13 l=8
+ ad=0 pd=0 as=0 ps=0 
M4799 n_923 pch3 GND GND efet w=33 l=6
+ ad=715 pd=200 as=0 ps=0 
M4800 GND n_1061 npchp3 GND efet w=45 l=7
+ ad=0 pd=0 as=882 ps=250 
M4801 n_207 n_810 GND GND efet w=33 l=6
+ ad=0 pd=0 as=0 ps=0 
M4802 n_356 n_293 n_207 GND efet w=44 l=6
+ ad=308 pd=102 as=0 ps=0 
M4803 GND n_923 n_356 GND efet w=44 l=5
+ ad=0 pd=0 as=0 ps=0 
M4804 dpc35_PCHC n_923 GND GND efet w=58 l=6
+ ad=0 pd=0 as=0 ps=0 
M4805 GND n_293 n_810 GND efet w=21 l=6
+ ad=0 pd=0 as=1074 ps=312 
M4806 n_810 n_923 GND GND efet w=25 l=6
+ ad=0 pd=0 as=0 ps=0 
M4807 adh3 dpc32_PCHADH pchp3 GND efet w=14 l=8
+ ad=0 pd=0 as=0 ps=0 
M4808 pchp4 dpc31_PCHPCH pch4 GND efet w=14 l=7
+ ad=1593 pd=394 as=626 ps=158 
M4809 pch4 dpc30_ADHPCH adh4 GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M4810 n_923 n_923 Vdd GND dfet w=9 l=20
+ ad=1509 pd=478 as=0 ps=0 
M4811 n_810 n_810 Vdd GND dfet w=10 l=15
+ ad=812 pd=252 as=0 ps=0 
M4812 n_83 n_83 Vdd GND dfet w=8 l=16
+ ad=1341 pd=394 as=0 ps=0 
M4813 n_1657 cclk npchp4 GND efet w=11 l=8
+ ad=1122 pd=292 as=192 ps=82 
M4814 Vdd n_523 n_523 GND dfet w=10 l=15
+ ad=0 pd=0 as=2251 ps=688 
M4815 GND npchp4 pchp4 GND efet w=57 l=6
+ ad=0 pd=0 as=0 ps=0 
M4816 n_949 n_83 n_523 GND efet w=43 l=7
+ ad=455 pd=116 as=420 ps=138 
M4817 GND dpc35_PCHC n_949 GND efet w=44 l=6
+ ad=0 pd=0 as=0 ps=0 
M4818 n_1400 pch4 GND GND efet w=43 l=7
+ ad=400 pd=118 as=0 ps=0 
M4819 Vdd n_1400 n_1400 GND dfet w=9 l=21
+ ad=0 pd=0 as=794 ps=222 
M4820 pchp4 dpc33_PCHDB idb4 GND efet w=14 l=8
+ ad=0 pd=0 as=0 ps=0 
M4821 n_1406 n_523 n_1657 GND efet w=57 l=7
+ ad=1191 pd=338 as=0 ps=0 
M4822 n_83 n_1400 GND GND efet w=22 l=6
+ ad=1169 pd=266 as=0 ps=0 
M4823 adh4 dpc32_PCHADH pchp4 GND efet w=14 l=8
+ ad=0 pd=0 as=0 ps=0 
M4824 pchp5 dpc31_PCHPCH pch5 GND efet w=14 l=7
+ ad=1613 pd=418 as=618 ps=156 
M4825 pch5 dpc30_ADHPCH adh5 GND efet w=13 l=7
+ ad=0 pd=0 as=0 ps=0 
M4826 pchp4 pchp4 Vdd GND dfet w=10 l=18
+ ad=486 pd=126 as=0 ps=0 
M4827 n_1406 n_83 GND GND efet w=55 l=7
+ ad=0 pd=0 as=0 ps=0 
M4828 n_1657 n_1657 Vdd GND dfet w=10 l=16
+ ad=373 pd=110 as=0 ps=0 
M4829 GND dpc35_PCHC n_1406 GND efet w=56 l=6
+ ad=0 pd=0 as=0 ps=0 
M4830 GND n_783 dpc34_PCLC GND efet w=56 l=6
+ ad=0 pd=0 as=0 ps=0 
M4831 pclp1 pclp1 Vdd GND dfet w=10 l=18
+ ad=489 pd=128 as=0 ps=0 
M4832 n_1158 n_783 GND GND efet w=39 l=6
+ ad=195 pd=88 as=0 ps=0 
M4833 n_515 n_1542 n_1158 GND efet w=39 l=7
+ ad=933 pd=240 as=0 ps=0 
M4834 Vdd n_515 n_515 GND dfet w=9 l=17
+ ad=0 pd=0 as=338 ps=84 
M4835 Vdd npclp2 npclp2 GND dfet w=11 l=21
+ ad=0 pd=0 as=1129 ps=342 
M4836 GND n_783 n_1253 GND efet w=24 l=6
+ ad=0 pd=0 as=1107 ps=314 
M4837 GND n_1253 n_515 GND efet w=34 l=6
+ ad=0 pd=0 as=0 ps=0 
M4838 n_515 cclk n_1411 GND efet w=12 l=8
+ ad=0 pd=0 as=160 ps=76 
M4839 Vdd pclp2 pclp2 GND dfet w=10 l=16
+ ad=0 pd=0 as=458 ps=122 
M4840 n_1253 n_1542 GND GND efet w=22 l=7
+ ad=0 pd=0 as=0 ps=0 
M4841 npclp2 n_1411 GND GND efet w=33 l=7
+ ad=857 pd=234 as=0 ps=0 
M4842 GND pcl2 n_783 GND efet w=33 l=7
+ ad=0 pd=0 as=720 ps=176 
M4843 pclp2 npclp2 GND GND efet w=61 l=6
+ ad=1678 pd=392 as=0 ps=0 
M4844 Vdd n_163 n_163 GND dfet w=9 l=16
+ ad=0 pd=0 as=1423 ps=416 
M4845 n_1253 n_1253 Vdd GND dfet w=9 l=13
+ ad=1893 pd=626 as=0 ps=0 
M4846 n_783 n_783 Vdd GND dfet w=10 l=20
+ ad=1550 pd=472 as=0 ps=0 
M4847 adl2 dpc38_PCLADL pclp2 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M4848 DBZ idb4 GND GND efet w=38 l=6
+ ad=0 pd=0 as=0 ps=0 
M4849 GND idb5 DBZ GND efet w=50 l=5
+ ad=0 pd=0 as=0 ps=0 
M4850 H1x1 H1x1 Vdd GND dfet w=11 l=16
+ ad=2685 pd=734 as=0 ps=0 
M4851 n_243 n_243 Vdd GND dfet w=10 l=12
+ ad=2207 pd=794 as=0 ps=0 
M4852 DBZ idb0 GND GND efet w=50 l=5
+ ad=0 pd=0 as=0 ps=0 
M4853 GND idb1 DBZ GND efet w=38 l=4
+ ad=0 pd=0 as=0 ps=0 
M4854 Vdd DBZ DBZ GND dfet w=10 l=10
+ ad=0 pd=0 as=882 ps=248 
M4855 n_566 n_755 n_580 GND efet w=39 l=5
+ ad=1342 pd=356 as=0 ps=0 
M4856 n_661 n_1170 n_566 GND efet w=58 l=6
+ ad=829 pd=182 as=0 ps=0 
M4857 n_318 cclk pipeUNK14 GND efet w=13 l=8
+ ad=1605 pd=364 as=150 ps=80 
M4858 GND pipeUNK14 n_661 GND efet w=81 l=5
+ ad=0 pd=0 as=0 ps=0 
M4859 GND p1 n_318 GND efet w=86 l=6
+ ad=0 pd=0 as=0 ps=0 
M4860 n_1115 n_1115 Vdd GND dfet w=10 l=12
+ ad=782 pd=226 as=0 ps=0 
M4861 n_1115 n_270 GND GND efet w=32 l=7
+ ad=641 pd=182 as=0 ps=0 
M4862 GND n_201 n_1433 GND efet w=41 l=7
+ ad=0 pd=0 as=0 ps=0 
M4863 Vdd n_1433 n_1433 GND dfet w=9 l=11
+ ad=0 pd=0 as=1414 ps=434 
M4864 n_1371 n_1045 GND GND efet w=40 l=6
+ ad=1047 pd=342 as=0 ps=0 
M4865 n_318 n_318 Vdd GND dfet w=9 l=12
+ ad=3100 pd=1018 as=0 ps=0 
M4866 Vdd n_1371 n_1371 GND dfet w=10 l=12
+ ad=0 pd=0 as=1327 ps=408 
M4867 n_1115 n_620 GND GND efet w=35 l=6
+ ad=0 pd=0 as=0 ps=0 
M4868 GND n_307 n_620 GND efet w=40 l=6
+ ad=0 pd=0 as=2023 ps=506 
M4869 GND n_201 n_1371 GND efet w=41 l=7
+ ad=0 pd=0 as=0 ps=0 
M4870 n_620 n_1433 GND GND efet w=41 l=7
+ ad=0 pd=0 as=0 ps=0 
M4871 n_1371 n_846 GND GND efet w=41 l=6
+ ad=0 pd=0 as=0 ps=0 
M4872 n_802 n_781 GND GND efet w=39 l=6
+ ad=273 pd=92 as=0 ps=0 
M4873 n_566 n_243 n_802 GND efet w=39 l=5
+ ad=0 pd=0 as=0 ps=0 
M4874 Vdd n_566 n_566 GND dfet w=9 l=13
+ ad=0 pd=0 as=341 ps=92 
M4875 p1 cp1 n_566 GND efet w=11 l=9
+ ad=153 pd=58 as=0 ps=0 
M4876 GND n_1371 n_620 GND efet w=41 l=7
+ ad=0 pd=0 as=0 ps=0 
M4877 n_620 n_620 Vdd GND dfet w=9 l=10
+ ad=1994 pd=624 as=0 ps=0 
M4878 GND n_1293 n_620 GND efet w=55 l=7
+ ad=0 pd=0 as=0 ps=0 
M4879 GND n_318 n_1293 GND efet w=41 l=7
+ ad=0 pd=0 as=1223 ps=336 
M4880 n_1579 cp1 notRnWprepad GND efet w=12 l=8
+ ad=174 pd=80 as=0 ps=0 
M4881 nDBE cclk GND GND efet w=123 l=6
+ ad=1525 pd=434 as=0 ps=0 
M4882 GND n_251 n_1028 GND efet w=90 l=6
+ ad=0 pd=0 as=785 ps=222 
M4883 n_1028 n_1028 Vdd GND dfet w=9 l=7
+ ad=704 pd=234 as=0 ps=0 
M4884 RnWstretched n_1028 Vdd GND dfet w=21 l=5
+ ad=4882 pd=920 as=0 ps=0 
M4885 GND n_251 RnWstretched GND efet w=164 l=6
+ ad=0 pd=0 as=0 ps=0 
M4886 n_251 n_221 GND GND efet w=103 l=6
+ ad=1659 pd=470 as=0 ps=0 
M4887 GND nDBE n_251 GND efet w=134 l=6
+ ad=0 pd=0 as=0 ps=0 
M4888 nDBZ DBZ GND GND efet w=63 l=7
+ ad=919 pd=282 as=0 ps=0 
M4889 RnWstretched n_251 GND GND efet w=161 l=8
+ ad=0 pd=0 as=0 ps=0 
M4890 GND n_251 RnWstretched GND efet w=157 l=7
+ ad=0 pd=0 as=0 ps=0 
M4891 GND n_962 nDBE GND efet w=118 l=6
+ ad=0 pd=0 as=0 ps=0 
M4892 n_1585 cclk GND GND efet w=35 l=7
+ ad=446 pd=152 as=0 ps=0 
M4893 n_1585 n_1585 Vdd GND dfet w=9 l=20
+ ad=844 pd=242 as=0 ps=0 
M4894 GND n_1579 n_221 GND efet w=75 l=6
+ ad=0 pd=0 as=910 ps=222 
M4895 n_962 n_1585 GND GND efet w=36 l=5
+ ad=640 pd=176 as=0 ps=0 
M4896 n_1293 nop_branch_bit6 GND GND efet w=40 l=6
+ ad=0 pd=0 as=0 ps=0 
M4897 Vdd n_1293 n_1293 GND dfet w=9 l=11
+ ad=0 pd=0 as=1264 ps=424 
M4898 GND nop_branch_bit6 n_846 GND efet w=27 l=7
+ ad=0 pd=0 as=964 ps=220 
M4899 GND nop_branch_bit7 n_1293 GND efet w=38 l=6
+ ad=0 pd=0 as=0 ps=0 
M4900 n_201 nop_branch_bit7 GND GND efet w=27 l=6
+ ad=666 pd=186 as=0 ps=0 
M4901 n_846 n_846 Vdd GND dfet w=10 l=17
+ ad=1856 pd=560 as=0 ps=0 
M4902 n_201 n_201 Vdd GND dfet w=9 l=16
+ ad=2964 pd=958 as=0 ps=0 
M4903 n_221 n_221 Vdd GND dfet w=10 l=12
+ ad=1720 pd=522 as=0 ps=0 
M4904 nDBZ nDBZ Vdd GND dfet w=11 l=11
+ ad=1668 pd=614 as=0 ps=0 
M4905 n_719 dpc41_DL_ADL adl0 GND efet w=63 l=7
+ ad=1959 pd=500 as=0 ps=0 
M4906 adl2 dpc40_ADLPCL pcl2 GND efet w=14 l=7
+ ad=0 pd=0 as=490 ps=98 
M4907 pcl2 dpc39_PCLPCL pclp2 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M4908 idb2 dpc37_PCLDB pclp2 GND efet w=13 l=8
+ ad=0 pd=0 as=0 ps=0 
M4909 Vdd n_249 n_249 GND dfet w=10 l=21
+ ad=0 pd=0 as=1268 ps=340 
M4910 GND pcl3 n_249 GND efet w=42 l=6
+ ad=0 pd=0 as=493 ps=122 
M4911 GND n_249 n_163 GND efet w=22 l=7
+ ad=0 pd=0 as=1178 ps=268 
M4912 n_1498 n_163 GND GND efet w=43 l=7
+ ad=465 pd=120 as=0 ps=0 
M4913 Vdd n_1184 n_1184 GND dfet w=10 l=14
+ ad=0 pd=0 as=2135 ps=720 
M4914 n_1184 n_1253 n_1498 GND efet w=43 l=6
+ ad=564 pd=138 as=0 ps=0 
M4915 npclp3 cclk n_1631 GND efet w=12 l=7
+ ad=216 pd=90 as=1186 ps=296 
M4916 GND n_249 dpc34_PCLC GND efet w=55 l=7
+ ad=0 pd=0 as=0 ps=0 
M4917 n_903 n_163 GND GND efet w=56 l=7
+ ad=1300 pd=340 as=0 ps=0 
M4918 GND n_1253 n_903 GND efet w=54 l=5
+ ad=0 pd=0 as=0 ps=0 
M4919 n_1631 n_1184 n_903 GND efet w=57 l=6
+ ad=0 pd=0 as=0 ps=0 
M4920 pclp3 npclp3 GND GND efet w=57 l=6
+ ad=1605 pd=364 as=0 ps=0 
M4921 adl3 dpc38_PCLADL pclp3 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M4922 adl3 dpc40_ADLPCL pcl3 GND efet w=14 l=8
+ ad=0 pd=0 as=469 ps=96 
M4923 pcl3 dpc39_PCLPCL pclp3 GND efet w=13 l=7
+ ad=0 pd=0 as=0 ps=0 
M4924 n_1631 n_1631 Vdd GND dfet w=10 l=16
+ ad=403 pd=110 as=0 ps=0 
M4925 idb3 dpc37_PCLDB pclp3 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M4926 pclp3 pclp3 Vdd GND dfet w=10 l=19
+ ad=476 pd=128 as=0 ps=0 
M4927 GND n_1643 dpc34_PCLC GND efet w=57 l=6
+ ad=0 pd=0 as=0 ps=0 
M4928 n_766 n_1643 GND GND efet w=39 l=6
+ ad=234 pd=90 as=0 ps=0 
M4929 n_474 n_1184 n_766 GND efet w=39 l=6
+ ad=947 pd=240 as=0 ps=0 
M4930 Vdd n_474 n_474 GND dfet w=9 l=15
+ ad=0 pd=0 as=284 ps=80 
M4931 Vdd npclp4 npclp4 GND dfet w=9 l=20
+ ad=0 pd=0 as=1149 ps=340 
M4932 GND n_1643 n_410 GND efet w=25 l=6
+ ad=0 pd=0 as=1130 ps=320 
M4933 GND n_410 n_474 GND efet w=34 l=6
+ ad=0 pd=0 as=0 ps=0 
M4934 n_474 cclk n_15 GND efet w=12 l=8
+ ad=0 pd=0 as=174 ps=74 
M4935 Vdd pclp4 pclp4 GND dfet w=9 l=16
+ ad=0 pd=0 as=390 ps=114 
M4936 n_410 n_1184 GND GND efet w=21 l=6
+ ad=0 pd=0 as=0 ps=0 
M4937 npclp4 n_15 GND GND efet w=33 l=6
+ ad=769 pd=230 as=0 ps=0 
M4938 GND pcl4 n_1643 GND efet w=33 l=7
+ ad=0 pd=0 as=744 ps=180 
M4939 pclp4 npclp4 GND GND efet w=60 l=6
+ ad=1633 pd=392 as=0 ps=0 
M4940 Vdd n_392 n_392 GND dfet w=9 l=16
+ ad=0 pd=0 as=1341 ps=412 
M4941 Vdd pchp5 pchp5 GND dfet w=10 l=15
+ ad=0 pd=0 as=429 ps=122 
M4942 Vdd npchp5 npchp5 GND dfet w=10 l=16
+ ad=0 pd=0 as=1114 ps=330 
M4943 Vdd n_875 n_875 GND dfet w=9 l=17
+ ad=0 pd=0 as=326 ps=84 
M4944 n_875 cclk n_469 GND efet w=12 l=8
+ ad=907 pd=238 as=162 ps=70 
M4945 GND npchp5 pchp5 GND efet w=61 l=6
+ ad=0 pd=0 as=0 ps=0 
M4946 pchp5 dpc33_PCHDB idb5 GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M4947 n_499 pch5 GND GND efet w=34 l=7
+ ad=704 pd=200 as=0 ps=0 
M4948 GND n_469 npchp5 GND efet w=42 l=7
+ ad=0 pd=0 as=812 ps=246 
M4949 n_875 n_743 GND GND efet w=33 l=6
+ ad=0 pd=0 as=0 ps=0 
M4950 n_1659 n_523 n_875 GND efet w=44 l=6
+ ad=264 pd=100 as=0 ps=0 
M4951 GND n_499 n_1659 GND efet w=44 l=6
+ ad=0 pd=0 as=0 ps=0 
M4952 GND n_523 n_743 GND efet w=22 l=6
+ ad=0 pd=0 as=1100 ps=298 
M4953 GND n_499 n_743 GND efet w=29 l=6
+ ad=0 pd=0 as=0 ps=0 
M4954 adh5 dpc32_PCHADH pchp5 GND efet w=13 l=7
+ ad=0 pd=0 as=0 ps=0 
M4955 pchp6 dpc31_PCHPCH pch6 GND efet w=14 l=7
+ ad=1596 pd=402 as=578 ps=156 
M4956 pch6 dpc30_ADHPCH adh6 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M4957 n_499 n_499 Vdd GND dfet w=9 l=20
+ ad=1682 pd=534 as=0 ps=0 
M4958 n_410 n_410 Vdd GND dfet w=9 l=13
+ ad=2045 pd=628 as=0 ps=0 
M4959 n_1643 n_1643 Vdd GND dfet w=10 l=21
+ ad=1548 pd=480 as=0 ps=0 
M4960 adl4 dpc38_PCLADL pclp4 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M4961 adl4 dpc40_ADLPCL pcl4 GND efet w=14 l=7
+ ad=0 pd=0 as=490 ps=98 
M4962 pcl4 dpc39_PCLPCL pclp4 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M4963 idb4 dpc37_PCLDB pclp4 GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M4964 Vdd n_386 n_386 GND dfet w=11 l=21
+ ad=0 pd=0 as=1148 ps=342 
M4965 GND pcl5 n_386 GND efet w=42 l=7
+ ad=0 pd=0 as=420 ps=126 
M4966 GND n_386 n_392 GND efet w=23 l=6
+ ad=0 pd=0 as=1155 ps=270 
M4967 n_814 n_392 GND GND efet w=43 l=7
+ ad=426 pd=118 as=0 ps=0 
M4968 Vdd n_344 n_344 GND dfet w=10 l=13
+ ad=0 pd=0 as=2033 ps=690 
M4969 n_344 n_410 n_814 GND efet w=45 l=7
+ ad=591 pd=146 as=0 ps=0 
M4970 npclp5 cclk n_1073 GND efet w=12 l=8
+ ad=204 pd=88 as=1175 ps=294 
M4971 n_743 n_743 Vdd GND dfet w=10 l=14
+ ad=2075 pd=634 as=0 ps=0 
M4972 n_1488 n_1488 Vdd GND dfet w=9 l=16
+ ad=1321 pd=404 as=0 ps=0 
M4973 n_1192 cclk npchp6 GND efet w=12 l=7
+ ad=1092 pd=288 as=193 ps=84 
M4974 Vdd n_609 n_609 GND dfet w=9 l=14
+ ad=0 pd=0 as=2141 ps=688 
M4975 GND npchp6 pchp6 GND efet w=57 l=6
+ ad=0 pd=0 as=0 ps=0 
M4976 n_545 n_743 n_609 GND efet w=44 l=7
+ ad=424 pd=120 as=472 ps=144 
M4977 GND n_1488 n_545 GND efet w=44 l=6
+ ad=0 pd=0 as=0 ps=0 
M4978 n_278 pch6 GND GND efet w=42 l=7
+ ad=408 pd=118 as=0 ps=0 
M4979 Vdd n_278 n_278 GND dfet w=10 l=20
+ ad=0 pd=0 as=782 ps=222 
M4980 pchp6 dpc33_PCHDB idb6 GND efet w=13 l=7
+ ad=0 pd=0 as=0 ps=0 
M4981 n_1547 n_609 n_1192 GND efet w=56 l=6
+ ad=1210 pd=342 as=0 ps=0 
M4982 n_1488 n_278 GND GND efet w=23 l=6
+ ad=1110 pd=270 as=0 ps=0 
M4983 GND n_386 dpc34_PCLC GND efet w=55 l=6
+ ad=0 pd=0 as=0 ps=0 
M4984 n_557 n_392 GND GND efet w=56 l=6
+ ad=1215 pd=336 as=0 ps=0 
M4985 GND n_410 n_557 GND efet w=52 l=7
+ ad=0 pd=0 as=0 ps=0 
M4986 n_1073 n_344 n_557 GND efet w=58 l=6
+ ad=0 pd=0 as=0 ps=0 
M4987 pclp5 npclp5 GND GND efet w=58 l=6
+ ad=1550 pd=352 as=0 ps=0 
M4988 adl5 dpc38_PCLADL pclp5 GND efet w=14 l=8
+ ad=0 pd=0 as=0 ps=0 
M4989 adl5 dpc40_ADLPCL pcl5 GND efet w=14 l=8
+ ad=0 pd=0 as=462 ps=94 
M4990 pcl5 dpc39_PCLPCL pclp5 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M4991 GND n_232 dpc34_PCLC GND efet w=56 l=7
+ ad=0 pd=0 as=0 ps=0 
M4992 n_1073 n_1073 Vdd GND dfet w=9 l=16
+ ad=394 pd=112 as=0 ps=0 
M4993 idb5 dpc37_PCLDB pclp5 GND efet w=14 l=6
+ ad=0 pd=0 as=0 ps=0 
M4994 pclp5 pclp5 Vdd GND dfet w=9 l=18
+ ad=485 pd=128 as=0 ps=0 
M4995 n_585 n_232 GND GND efet w=39 l=7
+ ad=195 pd=88 as=0 ps=0 
M4996 n_20 n_344 n_585 GND efet w=39 l=6
+ ad=976 pd=240 as=0 ps=0 
M4997 Vdd n_20 n_20 GND dfet w=10 l=17
+ ad=0 pd=0 as=337 ps=84 
M4998 Vdd npclp6 npclp6 GND dfet w=10 l=20
+ ad=0 pd=0 as=1100 ps=336 
M4999 adh6 dpc32_PCHADH pchp6 GND efet w=13 l=7
+ ad=0 pd=0 as=0 ps=0 
M5000 pchp7 dpc31_PCHPCH pch7 GND efet w=14 l=8
+ ad=1670 pd=424 as=599 ps=154 
M5001 pch7 dpc30_ADHPCH adh7 GND efet w=13 l=7
+ ad=0 pd=0 as=0 ps=0 
M5002 pchp6 pchp6 Vdd GND dfet w=11 l=18
+ ad=454 pd=120 as=0 ps=0 
M5003 n_1547 n_743 GND GND efet w=55 l=6
+ ad=0 pd=0 as=0 ps=0 
M5004 n_1192 n_1192 Vdd GND dfet w=10 l=16
+ ad=394 pd=112 as=0 ps=0 
M5005 GND n_1488 n_1547 GND efet w=54 l=6
+ ad=0 pd=0 as=0 ps=0 
M5006 Vdd pchp7 pchp7 GND dfet w=10 l=15
+ ad=0 pd=0 as=427 ps=122 
M5007 Vdd npchp7 npchp7 GND dfet w=10 l=16
+ ad=0 pd=0 as=1094 ps=328 
M5008 Vdd n_1209 n_1209 GND dfet w=9 l=17
+ ad=0 pd=0 as=326 ps=84 
M5009 n_1209 cclk n_663 GND efet w=11 l=8
+ ad=897 pd=234 as=155 ps=78 
M5010 GND npchp7 pchp7 GND efet w=60 l=6
+ ad=0 pd=0 as=0 ps=0 
M5011 pchp7 dpc33_PCHDB idb7 GND efet w=15 l=8
+ ad=0 pd=0 as=0 ps=0 
M5012 n_453 pch7 GND GND efet w=32 l=6
+ ad=688 pd=198 as=0 ps=0 
M5013 GND n_663 npchp7 GND efet w=42 l=6
+ ad=0 pd=0 as=898 ps=248 
M5014 n_1209 n_1213 GND GND efet w=33 l=7
+ ad=0 pd=0 as=0 ps=0 
M5015 n_1264 n_609 n_1209 GND efet w=44 l=6
+ ad=264 pd=100 as=0 ps=0 
M5016 GND n_453 n_1264 GND efet w=44 l=6
+ ad=0 pd=0 as=0 ps=0 
M5017 GND n_609 n_1213 GND efet w=23 l=6
+ ad=0 pd=0 as=1169 ps=312 
M5018 n_1213 n_453 GND GND efet w=22 l=6
+ ad=0 pd=0 as=0 ps=0 
M5019 GND n_232 n_1316 GND efet w=24 l=7
+ ad=0 pd=0 as=1181 ps=292 
M5020 GND n_1316 n_20 GND efet w=34 l=6
+ ad=0 pd=0 as=0 ps=0 
M5021 n_20 cclk n_993 GND efet w=13 l=9
+ ad=0 pd=0 as=172 ps=74 
M5022 Vdd pclp6 pclp6 GND dfet w=10 l=16
+ ad=0 pd=0 as=422 ps=116 
M5023 n_1316 n_344 GND GND efet w=21 l=6
+ ad=0 pd=0 as=0 ps=0 
M5024 npclp6 n_993 GND GND efet w=34 l=7
+ ad=788 pd=228 as=0 ps=0 
M5025 GND pcl6 n_232 GND efet w=33 l=7
+ ad=0 pd=0 as=720 ps=176 
M5026 pclp6 npclp6 GND GND efet w=61 l=6
+ ad=1713 pd=394 as=0 ps=0 
M5027 Vdd n_715 n_715 GND dfet w=10 l=16
+ ad=0 pd=0 as=1377 ps=414 
M5028 n_1316 n_1316 Vdd GND dfet w=9 l=13
+ ad=2039 pd=630 as=0 ps=0 
M5029 n_232 n_232 Vdd GND dfet w=10 l=21
+ ad=1632 pd=466 as=0 ps=0 
M5030 adl6 dpc38_PCLADL pclp6 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M5031 nDBE nDBE Vdd GND dfet w=9 l=8
+ ad=1521 pd=480 as=0 ps=0 
M5032 RnWstretched n_251 GND GND efet w=174 l=7
+ ad=0 pd=0 as=0 ps=0 
M5033 n_251 n_221 GND GND efet w=32 l=7
+ ad=0 pd=0 as=0 ps=0 
M5034 n_962 n_962 Vdd GND dfet w=9 l=13
+ ad=1247 pd=382 as=0 ps=0 
M5035 Vdd n_251 n_251 GND dfet w=18 l=7
+ ad=0 pd=0 as=6031 ps=1834 
M5036 Vdd n_1687 n_1687 GND dfet w=9 l=16
+ ad=0 pd=0 as=322 ps=84 
M5037 idl0 idl0 Vdd GND dfet w=10 l=17
+ ad=337 pd=84 as=0 ps=0 
M5038 n_1687 cp1 notdor0 GND efet w=12 l=8
+ ad=901 pd=270 as=215 ps=84 
M5039 idl0 cp1 n_719 GND efet w=61 l=7
+ ad=1393 pd=334 as=0 ps=0 
M5040 n_719 dpc42_DL_ADH adh0 GND efet w=43 l=7
+ ad=0 pd=0 as=0 ps=0 
M5041 GND idb0 n_1687 GND efet w=46 l=6
+ ad=0 pd=0 as=0 ps=0 
M5042 dor0 notdor0 GND GND efet w=69 l=6
+ ad=854 pd=252 as=0 ps=0 
M5043 GND notidl0 idl0 GND efet w=38 l=6
+ ad=0 pd=0 as=0 ps=0 
M5044 Vdd n_718 n_718 GND dfet w=10 l=7
+ ad=0 pd=0 as=256 ps=98 
M5045 db0 GND GND GND efet w=54 l=7
+ ad=26200 pd=4358 as=0 ps=0 
M5046 n_718 cclk notidl0 GND efet w=14 l=8
+ ad=1723 pd=380 as=234 ps=82 
M5047 GND db0 n_718 GND efet w=134 l=6
+ ad=0 pd=0 as=0 ps=0 
M5048 n_87 dpc41_DL_ADL adl1 GND efet w=62 l=7
+ ad=1952 pd=502 as=0 ps=0 
M5049 idb0 dpc43_DL_DB n_719 GND efet w=43 l=7
+ ad=0 pd=0 as=0 ps=0 
M5050 GND notidl0 idl0 GND efet w=33 l=5
+ ad=0 pd=0 as=0 ps=0 
M5051 db0 n_1325 Vdd GND efet w=637 l=7
+ ad=0 pd=0 as=0 ps=0 
M5052 n_1325 RnWstretched GND GND efet w=151 l=6
+ ad=2345 pd=548 as=0 ps=0 
M5053 GND RnWstretched n_1325 GND efet w=155 l=6
+ ad=0 pd=0 as=0 ps=0 
M5054 idl0 notidl0 GND GND efet w=49 l=6
+ ad=0 pd=0 as=0 ps=0 
M5055 GND RnWstretched n_769 GND efet w=72 l=6
+ ad=0 pd=0 as=799 ps=214 
M5056 GND n_769 n_1325 GND efet w=138 l=6
+ ad=0 pd=0 as=0 ps=0 
M5057 Vdd cclk idb0 GND efet w=22 l=8
+ ad=0 pd=0 as=0 ps=0 
M5058 n_1325 dor0 Vdd GND dfet w=16 l=7
+ ad=0 pd=0 as=0 ps=0 
M5059 Vdd n_769 n_769 GND dfet w=10 l=8
+ ad=0 pd=0 as=1463 ps=492 
M5060 n_1072 n_769 Vdd GND dfet w=17 l=6
+ ad=2457 pd=552 as=0 ps=0 
M5061 GND RnWstretched n_1072 GND efet w=94 l=6
+ ad=0 pd=0 as=0 ps=0 
M5062 GND RnWstretched n_1072 GND efet w=201 l=6
+ ad=0 pd=0 as=0 ps=0 
M5063 n_1072 dor0 GND GND efet w=148 l=6
+ ad=0 pd=0 as=0 ps=0 
M5064 n_769 dor0 GND GND efet w=59 l=6
+ ad=0 pd=0 as=0 ps=0 
M5065 db0 n_1072 GND GND efet w=111 l=6
+ ad=0 pd=0 as=0 ps=0 
M5066 GND n_1072 db0 GND efet w=216 l=6
+ ad=0 pd=0 as=0 ps=0 
M5067 db0 n_1072 GND GND efet w=213 l=6
+ ad=0 pd=0 as=0 ps=0 
M5068 db0 n_1325 Vdd GND efet w=634 l=7
+ ad=0 pd=0 as=0 ps=0 
M5069 GND n_1072 db0 GND efet w=11 l=6
+ ad=0 pd=0 as=0 ps=0 
M5070 dor0 dor0 Vdd GND dfet w=10 l=11
+ ad=2138 pd=672 as=0 ps=0 
M5071 Vdd n_1474 n_1474 GND dfet w=9 l=16
+ ad=0 pd=0 as=316 ps=82 
M5072 idl1 idl1 Vdd GND dfet w=9 l=17
+ ad=317 pd=84 as=0 ps=0 
M5073 n_1474 cp1 notdor1 GND efet w=11 l=9
+ ad=857 pd=262 as=216 ps=82 
M5074 idl1 cp1 n_87 GND efet w=63 l=7
+ ad=1347 pd=338 as=0 ps=0 
M5075 Vdd cclk adh3 GND efet w=22 l=6
+ ad=0 pd=0 as=0 ps=0 
M5076 adl4 cclk Vdd GND efet w=22 l=7
+ ad=0 pd=0 as=0 ps=0 
M5077 adl6 dpc40_ADLPCL pcl6 GND efet w=14 l=8
+ ad=0 pd=0 as=482 ps=96 
M5078 pcl6 dpc39_PCLPCL pclp6 GND efet w=15 l=8
+ ad=0 pd=0 as=0 ps=0 
M5079 idb6 dpc37_PCLDB pclp6 GND efet w=13 l=7
+ ad=0 pd=0 as=0 ps=0 
M5080 Vdd n_641 n_641 GND dfet w=10 l=21
+ ad=0 pd=0 as=1213 ps=322 
M5081 GND pcl7 n_641 GND efet w=43 l=6
+ ad=0 pd=0 as=474 ps=120 
M5082 GND n_641 n_715 GND efet w=23 l=7
+ ad=0 pd=0 as=1184 ps=276 
M5083 n_426 n_715 GND GND efet w=44 l=7
+ ad=481 pd=122 as=0 ps=0 
M5084 Vdd n_1386 n_1386 GND dfet w=10 l=15
+ ad=0 pd=0 as=1120 ps=322 
M5085 n_1386 n_1316 n_426 GND efet w=46 l=6
+ ad=501 pd=144 as=0 ps=0 
M5086 npclp7 cclk n_484 GND efet w=11 l=8
+ ad=217 pd=90 as=1075 ps=292 
M5087 adh7 dpc32_PCHADH pchp7 GND efet w=14 l=8
+ ad=0 pd=0 as=0 ps=0 
M5088 n_453 n_453 Vdd GND dfet w=9 l=21
+ ad=1116 pd=334 as=0 ps=0 
M5089 n_1213 n_1213 Vdd GND dfet w=10 l=14
+ ad=825 pd=254 as=0 ps=0 
M5090 dpc34_PCLC dpc34_PCLC Vdd GND dfet w=11 l=6
+ ad=9843 pd=3498 as=0 ps=0 
M5091 GND n_641 dpc34_PCLC GND efet w=47 l=7
+ ad=0 pd=0 as=0 ps=0 
M5092 n_914 n_715 GND GND efet w=56 l=6
+ ad=1196 pd=332 as=0 ps=0 
M5093 GND n_1316 n_914 GND efet w=52 l=6
+ ad=0 pd=0 as=0 ps=0 
M5094 n_484 n_1386 n_914 GND efet w=57 l=6
+ ad=0 pd=0 as=0 ps=0 
M5095 pclp7 npclp7 GND GND efet w=58 l=7
+ ad=1543 pd=384 as=0 ps=0 
M5096 adl7 dpc38_PCLADL pclp7 GND efet w=14 l=8
+ ad=0 pd=0 as=0 ps=0 
M5097 adl7 dpc40_ADLPCL pcl7 GND efet w=14 l=8
+ ad=0 pd=0 as=454 ps=92 
M5098 pcl7 dpc39_PCLPCL pclp7 GND efet w=14 l=8
+ ad=0 pd=0 as=0 ps=0 
M5099 n_484 n_484 Vdd GND dfet w=10 l=16
+ ad=394 pd=112 as=0 ps=0 
M5100 idb7 dpc37_PCLDB pclp7 GND efet w=14 l=7
+ ad=0 pd=0 as=0 ps=0 
M5101 pclp7 pclp7 Vdd GND dfet w=10 l=18
+ ad=474 pd=126 as=0 ps=0 
M5102 GND cclk dpc30_ADHPCH GND efet w=26 l=8
+ ad=0 pd=0 as=0 ps=0 
M5103 n_87 dpc42_DL_ADH adh1 GND efet w=43 l=7
+ ad=0 pd=0 as=0 ps=0 
M5104 GND idb1 n_1474 GND efet w=45 l=6
+ ad=0 pd=0 as=0 ps=0 
M5105 dor1 notdor1 GND GND efet w=69 l=6
+ ad=845 pd=250 as=0 ps=0 
M5106 GND notidl1 idl1 GND efet w=37 l=7
+ ad=0 pd=0 as=0 ps=0 
M5107 Vdd n_213 n_213 GND dfet w=10 l=7
+ ad=0 pd=0 as=246 ps=100 
M5108 db0 n_1072 GND GND efet w=211 l=6
+ ad=0 pd=0 as=0 ps=0 
M5109 GND n_1072 db0 GND efet w=11 l=6
+ ad=0 pd=0 as=0 ps=0 
M5110 n_213 cclk notidl1 GND efet w=14 l=8
+ ad=1840 pd=390 as=236 ps=78 
M5111 GND db1 n_213 GND efet w=135 l=6
+ ad=0 pd=0 as=0 ps=0 
M5112 n_1424 dpc41_DL_ADL adl2 GND efet w=62 l=6
+ ad=2072 pd=506 as=0 ps=0 
M5113 idb1 dpc43_DL_DB n_87 GND efet w=43 l=7
+ ad=0 pd=0 as=0 ps=0 
M5114 GND notidl1 idl1 GND efet w=33 l=6
+ ad=0 pd=0 as=0 ps=0 
M5115 n_798 RnWstretched GND GND efet w=151 l=6
+ ad=2291 pd=546 as=0 ps=0 
M5116 n_798 RnWstretched GND GND efet w=153 l=6
+ ad=0 pd=0 as=0 ps=0 
M5117 idl1 notidl1 GND GND efet w=49 l=6
+ ad=0 pd=0 as=0 ps=0 
M5118 GND n_288 n_798 GND efet w=139 l=6
+ ad=0 pd=0 as=0 ps=0 
M5119 GND RnWstretched n_288 GND efet w=73 l=7
+ ad=0 pd=0 as=770 ps=208 
M5120 Vdd cclk idb1 GND efet w=21 l=9
+ ad=0 pd=0 as=0 ps=0 
M5121 n_798 dor1 Vdd GND dfet w=17 l=7
+ ad=0 pd=0 as=0 ps=0 
M5122 Vdd n_288 n_288 GND dfet w=10 l=8
+ ad=0 pd=0 as=1507 ps=490 
M5123 n_794 n_288 Vdd GND dfet w=17 l=6
+ ad=2509 pd=558 as=0 ps=0 
M5124 GND RnWstretched n_794 GND efet w=95 l=6
+ ad=0 pd=0 as=0 ps=0 
M5125 db0 n_1072 GND GND efet w=157 l=6
+ ad=0 pd=0 as=0 ps=0 
M5126 db0 n_1072 GND GND efet w=130 l=7
+ ad=0 pd=0 as=0 ps=0 
M5127 GND n_794 db1 GND efet w=157 l=7
+ ad=0 pd=0 as=26638 ps=4386 
M5128 GND n_794 db1 GND efet w=130 l=7
+ ad=0 pd=0 as=0 ps=0 
M5129 db1 n_798 Vdd GND efet w=638 l=6
+ ad=0 pd=0 as=0 ps=0 
M5130 db1 n_794 GND GND efet w=281 l=6
+ ad=0 pd=0 as=0 ps=0 
M5131 GND RnWstretched n_794 GND efet w=200 l=6
+ ad=0 pd=0 as=0 ps=0 
M5132 n_794 dor1 GND GND efet w=149 l=6
+ ad=0 pd=0 as=0 ps=0 
M5133 n_288 dor1 GND GND efet w=58 l=6
+ ad=0 pd=0 as=0 ps=0 
M5134 GND n_794 db1 GND efet w=12 l=6
+ ad=0 pd=0 as=0 ps=0 
M5135 dor1 dor1 Vdd GND dfet w=9 l=12
+ ad=2173 pd=678 as=0 ps=0 
M5136 Vdd n_1376 n_1376 GND dfet w=10 l=16
+ ad=0 pd=0 as=326 ps=84 
M5137 idl2 idl2 Vdd GND dfet w=9 l=16
+ ad=301 pd=82 as=0 ps=0 
M5138 n_1376 cp1 notdor2 GND efet w=11 l=8
+ ad=903 pd=266 as=223 ps=82 
M5139 idl2 cp1 n_1424 GND efet w=60 l=7
+ ad=1368 pd=338 as=0 ps=0 
M5140 n_1424 dpc42_DL_ADH adh2 GND efet w=44 l=8
+ ad=0 pd=0 as=0 ps=0 
M5141 GND idb2 n_1376 GND efet w=46 l=6
+ ad=0 pd=0 as=0 ps=0 
M5142 dor2 notdor2 GND GND efet w=70 l=6
+ ad=855 pd=254 as=0 ps=0 
M5143 GND notidl2 idl2 GND efet w=38 l=6
+ ad=0 pd=0 as=0 ps=0 
M5144 Vdd n_1199 n_1199 GND dfet w=9 l=7
+ ad=0 pd=0 as=251 ps=96 
M5145 db1 n_794 GND GND efet w=223 l=5
+ ad=0 pd=0 as=0 ps=0 
M5146 db1 n_798 Vdd GND efet w=639 l=6
+ ad=0 pd=0 as=0 ps=0 
M5147 GND n_794 db1 GND efet w=11 l=6
+ ad=0 pd=0 as=0 ps=0 
M5148 n_1661 dpc41_DL_ADL adl3 GND efet w=60 l=7
+ ad=1972 pd=500 as=0 ps=0 
M5149 adh4 cclk Vdd GND efet w=22 l=6
+ ad=0 pd=0 as=0 ps=0 
M5150 adl5 cclk Vdd GND efet w=23 l=6
+ ad=0 pd=0 as=0 ps=0 
M5151 adh5 cclk Vdd GND efet w=25 l=7
+ ad=0 pd=0 as=0 ps=0 
M5152 idb2 dpc43_DL_DB n_1424 GND efet w=44 l=7
+ ad=0 pd=0 as=0 ps=0 
M5153 GND notidl2 idl2 GND efet w=33 l=5
+ ad=0 pd=0 as=0 ps=0 
M5154 n_1199 cclk notidl2 GND efet w=14 l=7
+ ad=1730 pd=384 as=219 ps=72 
M5155 GND db2 n_1199 GND efet w=132 l=6
+ ad=0 pd=0 as=0 ps=0 
M5156 idl2 notidl2 GND GND efet w=49 l=7
+ ad=0 pd=0 as=0 ps=0 
M5157 n_520 RnWstretched GND GND efet w=153 l=6
+ ad=2224 pd=550 as=0 ps=0 
M5158 n_520 RnWstretched GND GND efet w=154 l=5
+ ad=0 pd=0 as=0 ps=0 
M5159 GND n_224 n_520 GND efet w=140 l=6
+ ad=0 pd=0 as=0 ps=0 
M5160 GND RnWstretched n_224 GND efet w=74 l=6
+ ad=0 pd=0 as=756 ps=212 
M5161 Vdd cclk idb2 GND efet w=22 l=8
+ ad=0 pd=0 as=0 ps=0 
M5162 n_520 dor2 Vdd GND dfet w=16 l=7
+ ad=0 pd=0 as=0 ps=0 
M5163 Vdd n_224 n_224 GND dfet w=9 l=8
+ ad=0 pd=0 as=1623 ps=492 
M5164 n_37 n_224 Vdd GND dfet w=17 l=7
+ ad=2514 pd=558 as=0 ps=0 
M5165 GND RnWstretched n_37 GND efet w=95 l=6
+ ad=0 pd=0 as=0 ps=0 
M5166 GND RnWstretched n_37 GND efet w=201 l=6
+ ad=0 pd=0 as=0 ps=0 
M5167 n_37 dor2 GND GND efet w=148 l=6
+ ad=0 pd=0 as=0 ps=0 
M5168 n_224 dor2 GND GND efet w=60 l=7
+ ad=0 pd=0 as=0 ps=0 
M5169 GND n_794 db1 GND efet w=245 l=6
+ ad=0 pd=0 as=0 ps=0 
M5170 GND GND db1 GND efet w=57 l=8
+ ad=0 pd=0 as=0 ps=0 
M5171 GND GND db2 GND efet w=55 l=6
+ ad=0 pd=0 as=24805 ps=4260 
M5172 db2 n_520 Vdd GND efet w=639 l=7
+ ad=0 pd=0 as=0 ps=0 
M5173 dor2 dor2 Vdd GND dfet w=10 l=12
+ ad=2317 pd=676 as=0 ps=0 
M5174 Vdd n_457 n_457 GND dfet w=9 l=17
+ ad=0 pd=0 as=338 ps=86 
M5175 idl3 idl3 Vdd GND dfet w=9 l=17
+ ad=317 pd=84 as=0 ps=0 
M5176 n_457 cp1 notdor3 GND efet w=12 l=8
+ ad=955 pd=274 as=203 ps=80 
M5177 idl3 cp1 n_1661 GND efet w=60 l=7
+ ad=1315 pd=330 as=0 ps=0 
M5178 n_1661 dpc42_DL_ADH adh3 GND efet w=44 l=8
+ ad=0 pd=0 as=0 ps=0 
M5179 GND idb3 n_457 GND efet w=46 l=6
+ ad=0 pd=0 as=0 ps=0 
M5180 dor3 notdor3 GND GND efet w=68 l=6
+ ad=874 pd=248 as=0 ps=0 
M5181 GND notidl3 idl3 GND efet w=37 l=7
+ ad=0 pd=0 as=0 ps=0 
M5182 Vdd n_896 n_896 GND dfet w=10 l=7
+ ad=0 pd=0 as=256 ps=98 
M5183 db2 n_37 db2 GND efet w=8 l=6
+ ad=0 pd=0 as=0 ps=0 
M5184 n_896 cclk notidl3 GND efet w=14 l=8
+ ad=1754 pd=384 as=226 ps=74 
M5185 db2 n_37 GND GND efet w=225 l=6
+ ad=0 pd=0 as=0 ps=0 
M5186 GND n_37 db2 GND efet w=8 l=6
+ ad=0 pd=0 as=0 ps=0 
M5187 GND db3 n_896 GND efet w=134 l=7
+ ad=0 pd=0 as=0 ps=0 
M5188 n_1095 dpc41_DL_ADL adl4 GND efet w=61 l=7
+ ad=2025 pd=504 as=0 ps=0 
M5189 idb3 dpc43_DL_DB n_1661 GND efet w=43 l=6
+ ad=0 pd=0 as=0 ps=0 
M5190 GND notidl3 idl3 GND efet w=34 l=6
+ ad=0 pd=0 as=0 ps=0 
M5191 n_42 RnWstretched GND GND efet w=152 l=6
+ ad=2217 pd=550 as=0 ps=0 
M5192 n_42 RnWstretched GND GND efet w=153 l=5
+ ad=0 pd=0 as=0 ps=0 
M5193 idl3 notidl3 GND GND efet w=48 l=6
+ ad=0 pd=0 as=0 ps=0 
M5194 GND n_1613 n_42 GND efet w=141 l=6
+ ad=0 pd=0 as=0 ps=0 
M5195 GND RnWstretched n_1613 GND efet w=74 l=7
+ ad=0 pd=0 as=750 ps=210 
M5196 Vdd cclk idb3 GND efet w=23 l=8
+ ad=0 pd=0 as=0 ps=0 
M5197 n_42 dor3 Vdd GND dfet w=16 l=7
+ ad=0 pd=0 as=0 ps=0 
M5198 db2 n_37 GND GND efet w=225 l=6
+ ad=0 pd=0 as=0 ps=0 
M5199 db2 n_520 Vdd GND efet w=638 l=6
+ ad=0 pd=0 as=0 ps=0 
M5200 GND n_37 db2 GND efet w=11 l=6
+ ad=0 pd=0 as=0 ps=0 
M5201 Vdd n_1613 n_1613 GND dfet w=10 l=8
+ ad=0 pd=0 as=1542 ps=490 
M5202 n_643 n_1613 Vdd GND dfet w=17 l=6
+ ad=2544 pd=556 as=0 ps=0 
M5203 GND RnWstretched n_643 GND efet w=94 l=6
+ ad=0 pd=0 as=0 ps=0 
M5204 GND RnWstretched n_643 GND efet w=200 l=6
+ ad=0 pd=0 as=0 ps=0 
M5205 n_643 dor3 GND GND efet w=148 l=6
+ ad=0 pd=0 as=0 ps=0 
M5206 n_1613 dor3 GND GND efet w=59 l=7
+ ad=0 pd=0 as=0 ps=0 
M5207 dor3 dor3 Vdd GND dfet w=10 l=12
+ ad=2316 pd=674 as=0 ps=0 
M5208 Vdd n_797 n_797 GND dfet w=9 l=17
+ ad=0 pd=0 as=348 ps=86 
M5209 idl4 idl4 Vdd GND dfet w=10 l=17
+ ad=343 pd=86 as=0 ps=0 
M5210 n_797 cp1 notdor4 GND efet w=11 l=8
+ ad=844 pd=268 as=194 ps=78 
M5211 idl4 cp1 n_1095 GND efet w=62 l=7
+ ad=1291 pd=334 as=0 ps=0 
M5212 n_1095 dpc42_DL_ADH adh4 GND efet w=43 l=8
+ ad=0 pd=0 as=0 ps=0 
M5213 GND idb4 n_797 GND efet w=46 l=6
+ ad=0 pd=0 as=0 ps=0 
M5214 dor4 notdor4 GND GND efet w=69 l=6
+ ad=878 pd=250 as=0 ps=0 
M5215 GND notidl4 idl4 GND efet w=38 l=7
+ ad=0 pd=0 as=0 ps=0 
M5216 db2 n_37 GND GND efet w=242 l=6
+ ad=0 pd=0 as=0 ps=0 
M5217 GND n_37 db2 GND efet w=11 l=6
+ ad=0 pd=0 as=0 ps=0 
M5218 db2 n_37 GND GND efet w=182 l=6
+ ad=0 pd=0 as=0 ps=0 
M5219 db2 n_37 GND GND efet w=156 l=6
+ ad=0 pd=0 as=0 ps=0 
M5220 GND n_643 db3 GND efet w=156 l=7
+ ad=0 pd=0 as=25724 ps=4350 
M5221 GND n_643 db3 GND efet w=236 l=7
+ ad=0 pd=0 as=0 ps=0 
M5222 Vdd n_490 n_490 GND dfet w=10 l=8
+ ad=0 pd=0 as=279 ps=100 
M5223 db3 n_42 Vdd GND efet w=636 l=6
+ ad=0 pd=0 as=0 ps=0 
M5224 db3 n_643 GND GND efet w=212 l=6
+ ad=0 pd=0 as=0 ps=0 
M5225 n_490 cclk notidl4 GND efet w=13 l=8
+ ad=1750 pd=378 as=214 ps=76 
M5226 GND db4 n_490 GND efet w=132 l=6
+ ad=0 pd=0 as=0 ps=0 
M5227 n_1387 dpc41_DL_ADL adl5 GND efet w=61 l=6
+ ad=2026 pd=506 as=0 ps=0 
M5228 adl6 cclk Vdd GND efet w=23 l=7
+ ad=0 pd=0 as=0 ps=0 
M5229 Vdd cclk adh6 GND efet w=25 l=7
+ ad=0 pd=0 as=0 ps=0 
M5230 Vdd cclk adl7 GND efet w=23 l=7
+ ad=0 pd=0 as=0 ps=0 
M5231 dpc31_PCHPCH cclk GND GND efet w=26 l=7
+ ad=0 pd=0 as=0 ps=0 
M5232 aluvout aluvout Vdd GND dfet w=10 l=7
+ ad=10389 pd=3534 as=0 ps=0 
M5233 n_1267 n_1267 Vdd GND dfet w=9 l=10
+ ad=232 pd=74 as=0 ps=0 
M5234 n_676 abh1 GND GND efet w=147 l=7
+ ad=1092 pd=352 as=0 ps=0 
M5235 Vdd n_617 n_676 GND dfet w=19 l=7
+ ad=0 pd=0 as=0 ps=0 
M5236 nABH1 cclk n_676 GND efet w=12 l=8
+ ad=408 pd=118 as=0 ps=0 
M5237 n_1298 ADH_ABH nABH1 GND efet w=12 l=8
+ ad=72 pd=36 as=0 ps=0 
M5238 n_1267 cp1 n_1298 GND efet w=12 l=7
+ ad=922 pd=242 as=0 ps=0 
M5239 GND adh1 n_1267 GND efet w=75 l=7
+ ad=0 pd=0 as=0 ps=0 
M5240 n_168 adh2 GND GND efet w=75 l=7
+ ad=871 pd=244 as=0 ps=0 
M5241 Vdd n_168 n_168 GND dfet w=10 l=9
+ ad=0 pd=0 as=203 ps=72 
M5242 abh2 nABH2 GND GND efet w=66 l=7
+ ad=522 pd=190 as=0 ps=0 
M5243 Vdd abh2 abh2 GND dfet w=9 l=15
+ ad=0 pd=0 as=2166 ps=662 
M5244 GND n_1034 n_1545 GND efet w=113 l=5
+ ad=0 pd=0 as=1934 ps=404 
M5245 GND n_1346 n_1296 GND efet w=113 l=5
+ ad=0 pd=0 as=1922 ps=404 
M5246 n_1545 abh2 Vdd GND dfet w=17 l=6
+ ad=0 pd=0 as=0 ps=0 
M5247 Vdd n_1034 n_1034 GND dfet w=9 l=10
+ ad=0 pd=0 as=1974 ps=680 
M5248 GND abh2 n_1034 GND efet w=44 l=7
+ ad=0 pd=0 as=471 ps=146 
M5249 n_836 cp1 n_168 GND efet w=12 l=8
+ ad=60 pd=34 as=0 ps=0 
M5250 nABH2 ADH_ABH n_836 GND efet w=12 l=8
+ ad=397 pd=114 as=0 ps=0 
M5251 nABH2 cclk n_994 GND efet w=12 l=8
+ ad=0 pd=0 as=1180 ps=356 
M5252 Vdd n_1034 n_994 GND dfet w=18 l=8
+ ad=0 pd=0 as=0 ps=0 
M5253 GND abh2 n_994 GND efet w=148 l=7
+ ad=0 pd=0 as=0 ps=0 
M5254 GND n_676 ab9 GND efet w=41 l=5
+ ad=0 pd=0 as=0 ps=0 
M5255 GND n_676 ab9 GND efet w=12 l=5
+ ad=0 pd=0 as=0 ps=0 
M5256 GND n_676 ab9 GND efet w=163 l=7
+ ad=0 pd=0 as=0 ps=0 
M5257 ab9 n_676 GND GND efet w=163 l=7
+ ad=0 pd=0 as=0 ps=0 
M5258 GND n_676 ab9 GND efet w=163 l=6
+ ad=0 pd=0 as=0 ps=0 
M5259 ab9 n_676 GND GND efet w=163 l=7
+ ad=0 pd=0 as=0 ps=0 
M5260 GND n_676 ab9 GND efet w=163 l=7
+ ad=0 pd=0 as=0 ps=0 
M5261 GND n_994 ab10 GND efet w=13 l=6
+ ad=0 pd=0 as=18798 ps=2312 
M5262 GND n_994 ab10 GND efet w=41 l=6
+ ad=0 pd=0 as=0 ps=0 
M5263 ab10 n_994 GND GND efet w=163 l=6
+ ad=0 pd=0 as=0 ps=0 
M5264 GND n_994 ab10 GND efet w=163 l=6
+ ad=0 pd=0 as=0 ps=0 
M5265 ab10 n_994 GND GND efet w=163 l=6
+ ad=0 pd=0 as=0 ps=0 
M5266 GND n_994 ab10 GND efet w=163 l=7
+ ad=0 pd=0 as=0 ps=0 
M5267 ab10 n_994 GND GND efet w=163 l=7
+ ad=0 pd=0 as=0 ps=0 
M5268 Vdd n_1545 ab10 GND efet w=416 l=6
+ ad=0 pd=0 as=0 ps=0 
M5269 Vdd n_1545 ab10 GND efet w=316 l=6
+ ad=0 pd=0 as=0 ps=0 
M5270 Vdd n_1545 ab10 GND efet w=159 l=7
+ ad=0 pd=0 as=0 ps=0 
M5271 ab11 n_1296 Vdd GND efet w=159 l=7
+ ad=18508 pd=2312 as=0 ps=0 
M5272 Vdd n_1296 ab11 GND efet w=318 l=6
+ ad=0 pd=0 as=0 ps=0 
M5273 Vdd n_1296 ab11 GND efet w=418 l=7
+ ad=0 pd=0 as=0 ps=0 
M5274 Vdd abh3 n_1296 GND dfet w=17 l=7
+ ad=0 pd=0 as=0 ps=0 
M5275 n_1346 abh3 GND GND efet w=46 l=7
+ ad=463 pd=134 as=0 ps=0 
M5276 Vdd n_1346 n_1346 GND dfet w=9 l=10
+ ad=0 pd=0 as=1873 ps=680 
M5277 abh3 abh3 Vdd GND dfet w=8 l=13
+ ad=2305 pd=660 as=0 ps=0 
M5278 GND nABH3 abh3 GND efet w=65 l=6
+ ad=0 pd=0 as=622 ps=188 
M5279 n_883 n_883 Vdd GND dfet w=9 l=9
+ ad=213 pd=72 as=0 ps=0 
M5280 n_359 abh3 GND GND efet w=149 l=7
+ ad=1045 pd=346 as=0 ps=0 
M5281 Vdd n_1346 n_359 GND dfet w=19 l=6
+ ad=0 pd=0 as=0 ps=0 
M5282 nABH3 cclk n_359 GND efet w=11 l=7
+ ad=392 pd=118 as=0 ps=0 
M5283 n_1667 ADH_ABH nABH3 GND efet w=11 l=8
+ ad=55 pd=32 as=0 ps=0 
M5284 n_883 cp1 n_1667 GND efet w=11 l=7
+ ad=957 pd=240 as=0 ps=0 
M5285 GND adh3 n_883 GND efet w=75 l=6
+ ad=0 pd=0 as=0 ps=0 
M5286 n_212 adh4 GND GND efet w=75 l=6
+ ad=802 pd=244 as=0 ps=0 
M5287 Vdd n_212 n_212 GND dfet w=9 l=10
+ ad=0 pd=0 as=242 ps=76 
M5288 abh4 nABH4 GND GND efet w=65 l=7
+ ad=503 pd=184 as=0 ps=0 
M5289 Vdd abh4 abh4 GND dfet w=9 l=14
+ ad=0 pd=0 as=2256 ps=660 
M5290 GND n_1677 n_475 GND efet w=112 l=7
+ ad=0 pd=0 as=1681 ps=386 
M5291 GND n_1423 n_1608 GND efet w=113 l=7
+ ad=0 pd=0 as=1723 ps=388 
M5292 n_475 abh4 Vdd GND dfet w=17 l=7
+ ad=0 pd=0 as=0 ps=0 
M5293 Vdd n_1677 n_1677 GND dfet w=10 l=9
+ ad=0 pd=0 as=2162 ps=676 
M5294 GND abh4 n_1677 GND efet w=45 l=6
+ ad=0 pd=0 as=552 ps=154 
M5295 n_1451 cp1 n_212 GND efet w=12 l=8
+ ad=48 pd=32 as=0 ps=0 
M5296 nABH4 ADH_ABH n_1451 GND efet w=12 l=8
+ ad=385 pd=112 as=0 ps=0 
M5297 nABH4 cclk n_999 GND efet w=11 l=8
+ ad=0 pd=0 as=1216 ps=356 
M5298 Vdd n_1677 n_999 GND dfet w=20 l=7
+ ad=0 pd=0 as=0 ps=0 
M5299 GND abh4 n_999 GND efet w=147 l=6
+ ad=0 pd=0 as=0 ps=0 
M5300 GND n_359 ab11 GND efet w=41 l=6
+ ad=0 pd=0 as=0 ps=0 
M5301 GND n_359 ab11 GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M5302 GND n_359 ab11 GND efet w=163 l=6
+ ad=0 pd=0 as=0 ps=0 
M5303 ab11 n_359 GND GND efet w=163 l=6
+ ad=0 pd=0 as=0 ps=0 
M5304 GND n_359 ab11 GND efet w=163 l=6
+ ad=0 pd=0 as=0 ps=0 
M5305 ab11 n_359 GND GND efet w=163 l=8
+ ad=0 pd=0 as=0 ps=0 
M5306 GND n_359 ab11 GND efet w=163 l=7
+ ad=0 pd=0 as=0 ps=0 
M5307 GND n_999 ab12 GND efet w=13 l=5
+ ad=0 pd=0 as=18767 ps=2320 
M5308 GND n_999 ab12 GND efet w=41 l=5
+ ad=0 pd=0 as=0 ps=0 
M5309 ab12 n_999 GND GND efet w=164 l=7
+ ad=0 pd=0 as=0 ps=0 
M5310 GND n_999 ab12 GND efet w=164 l=6
+ ad=0 pd=0 as=0 ps=0 
M5311 ab12 n_999 GND GND efet w=164 l=6
+ ad=0 pd=0 as=0 ps=0 
M5312 GND n_999 ab12 GND efet w=163 l=6
+ ad=0 pd=0 as=0 ps=0 
M5313 ab12 n_999 GND GND efet w=163 l=6
+ ad=0 pd=0 as=0 ps=0 
M5314 Vdd n_475 ab12 GND efet w=416 l=7
+ ad=0 pd=0 as=0 ps=0 
M5315 Vdd n_475 ab12 GND efet w=315 l=6
+ ad=0 pd=0 as=0 ps=0 
M5316 Vdd n_475 ab12 GND efet w=160 l=7
+ ad=0 pd=0 as=0 ps=0 
M5317 ab13 n_1608 Vdd GND efet w=160 l=7
+ ad=18253 pd=2310 as=0 ps=0 
M5318 Vdd n_1608 ab13 GND efet w=316 l=6
+ ad=0 pd=0 as=0 ps=0 
M5319 Vdd n_1608 ab13 GND efet w=416 l=7
+ ad=0 pd=0 as=0 ps=0 
M5320 Vdd abh5 n_1608 GND dfet w=17 l=7
+ ad=0 pd=0 as=0 ps=0 
M5321 n_1423 abh5 GND GND efet w=44 l=7
+ ad=443 pd=134 as=0 ps=0 
M5322 Vdd n_1423 n_1423 GND dfet w=9 l=11
+ ad=0 pd=0 as=2215 ps=682 
M5323 abh5 abh5 Vdd GND dfet w=10 l=13
+ ad=2150 pd=660 as=0 ps=0 
M5324 GND nABH5 abh5 GND efet w=66 l=7
+ ad=0 pd=0 as=659 ps=192 
M5325 Vdd cclk adh7 GND efet w=23 l=7
+ ad=0 pd=0 as=0 ps=0 
M5326 dpc39_PCLPCL cclk GND GND efet w=27 l=9
+ ad=0 pd=0 as=0 ps=0 
M5327 dpc40_ADLPCL cclk GND GND efet w=26 l=9
+ ad=0 pd=0 as=0 ps=0 
M5328 idb4 dpc43_DL_DB n_1095 GND efet w=44 l=7
+ ad=0 pd=0 as=0 ps=0 
M5329 GND notidl4 idl4 GND efet w=33 l=6
+ ad=0 pd=0 as=0 ps=0 
M5330 n_1076 RnWstretched GND GND efet w=152 l=6
+ ad=2321 pd=550 as=0 ps=0 
M5331 GND RnWstretched n_1076 GND efet w=156 l=6
+ ad=0 pd=0 as=0 ps=0 
M5332 idl4 notidl4 GND GND efet w=48 l=7
+ ad=0 pd=0 as=0 ps=0 
M5333 GND RnWstretched n_1463 GND efet w=73 l=6
+ ad=0 pd=0 as=765 ps=208 
M5334 GND n_1463 n_1076 GND efet w=137 l=6
+ ad=0 pd=0 as=0 ps=0 
M5335 Vdd cclk idb4 GND efet w=22 l=8
+ ad=0 pd=0 as=0 ps=0 
M5336 n_1076 dor4 Vdd GND dfet w=16 l=7
+ ad=0 pd=0 as=0 ps=0 
M5337 GND n_643 db3 GND efet w=12 l=6
+ ad=0 pd=0 as=0 ps=0 
M5338 Vdd n_1463 n_1463 GND dfet w=9 l=8
+ ad=0 pd=0 as=1554 ps=492 
M5339 n_147 n_1463 Vdd GND dfet w=17 l=7
+ ad=2471 pd=548 as=0 ps=0 
M5340 GND RnWstretched n_147 GND efet w=95 l=6
+ ad=0 pd=0 as=0 ps=0 
M5341 GND RnWstretched n_147 GND efet w=201 l=6
+ ad=0 pd=0 as=0 ps=0 
M5342 n_147 dor4 GND GND efet w=147 l=6
+ ad=0 pd=0 as=0 ps=0 
M5343 n_1463 dor4 GND GND efet w=58 l=6
+ ad=0 pd=0 as=0 ps=0 
M5344 dor4 dor4 Vdd GND dfet w=9 l=11
+ ad=2156 pd=674 as=0 ps=0 
M5345 Vdd n_961 n_961 GND dfet w=10 l=17
+ ad=0 pd=0 as=332 ps=84 
M5346 idl5 idl5 Vdd GND dfet w=9 l=17
+ ad=317 pd=84 as=0 ps=0 
M5347 n_961 cp1 notdor5 GND efet w=11 l=8
+ ad=863 pd=270 as=215 ps=78 
M5348 idl5 cp1 n_1387 GND efet w=63 l=7
+ ad=1369 pd=336 as=0 ps=0 
M5349 n_1387 dpc42_DL_ADH adh5 GND efet w=43 l=8
+ ad=0 pd=0 as=0 ps=0 
M5350 GND idb5 n_961 GND efet w=46 l=6
+ ad=0 pd=0 as=0 ps=0 
M5351 dor5 notdor5 GND GND efet w=69 l=6
+ ad=920 pd=254 as=0 ps=0 
M5352 GND notidl5 idl5 GND efet w=38 l=7
+ ad=0 pd=0 as=0 ps=0 
M5353 Vdd n_568 n_568 GND dfet w=10 l=7
+ ad=0 pd=0 as=262 ps=98 
M5354 n_568 cclk notidl5 GND efet w=14 l=8
+ ad=1845 pd=382 as=217 ps=76 
M5355 GND db5 n_568 GND efet w=133 l=6
+ ad=0 pd=0 as=0 ps=0 
M5356 n_1014 dpc41_DL_ADL adl6 GND efet w=64 l=7
+ ad=2002 pd=506 as=0 ps=0 
M5357 idb5 dpc43_DL_DB n_1387 GND efet w=43 l=7
+ ad=0 pd=0 as=0 ps=0 
M5358 GND notidl5 idl5 GND efet w=33 l=6
+ ad=0 pd=0 as=0 ps=0 
M5359 db3 n_643 GND GND efet w=212 l=6
+ ad=0 pd=0 as=0 ps=0 
M5360 GND n_643 db3 GND efet w=11 l=6
+ ad=0 pd=0 as=0 ps=0 
M5361 db3 n_42 Vdd GND efet w=640 l=6
+ ad=0 pd=0 as=0 ps=0 
M5362 GND n_643 db3 GND efet w=234 l=6
+ ad=0 pd=0 as=0 ps=0 
M5363 GND GND db3 GND efet w=54 l=7
+ ad=0 pd=0 as=0 ps=0 
M5364 GND GND db4 GND efet w=55 l=7
+ ad=0 pd=0 as=27574 ps=4708 
M5365 n_373 RnWstretched GND GND efet w=152 l=6
+ ad=2299 pd=548 as=0 ps=0 
M5366 n_373 RnWstretched GND GND efet w=155 l=6
+ ad=0 pd=0 as=0 ps=0 
M5367 idl5 notidl5 GND GND efet w=48 l=7
+ ad=0 pd=0 as=0 ps=0 
M5368 GND n_1720 n_373 GND efet w=139 l=6
+ ad=0 pd=0 as=0 ps=0 
M5369 GND RnWstretched n_1720 GND efet w=74 l=7
+ ad=0 pd=0 as=746 ps=212 
M5370 Vdd cclk idb5 GND efet w=21 l=8
+ ad=0 pd=0 as=0 ps=0 
M5371 n_373 dor5 Vdd GND dfet w=17 l=7
+ ad=0 pd=0 as=0 ps=0 
M5372 db4 n_1076 Vdd GND efet w=639 l=7
+ ad=0 pd=0 as=0 ps=0 
M5373 db4 n_147 db4 GND efet w=9 l=5
+ ad=0 pd=0 as=0 ps=0 
M5374 Vdd n_1720 n_1720 GND dfet w=10 l=8
+ ad=0 pd=0 as=1505 ps=490 
M5375 n_612 n_1720 Vdd GND dfet w=17 l=6
+ ad=2345 pd=552 as=0 ps=0 
M5376 GND RnWstretched n_612 GND efet w=95 l=7
+ ad=0 pd=0 as=0 ps=0 
M5377 GND RnWstretched n_612 GND efet w=201 l=7
+ ad=0 pd=0 as=0 ps=0 
M5378 n_612 dor5 GND GND efet w=147 l=6
+ ad=0 pd=0 as=0 ps=0 
M5379 n_1720 dor5 GND GND efet w=59 l=7
+ ad=0 pd=0 as=0 ps=0 
M5380 db4 n_147 GND GND efet w=216 l=6
+ ad=0 pd=0 as=0 ps=0 
M5381 GND n_147 db4 GND efet w=9 l=5
+ ad=0 pd=0 as=0 ps=0 
M5382 dor5 dor5 Vdd GND dfet w=9 l=12
+ ad=2316 pd=674 as=0 ps=0 
M5383 Vdd n_1684 n_1684 GND dfet w=9 l=17
+ ad=0 pd=0 as=343 ps=86 
M5384 idl6 idl6 Vdd GND dfet w=9 l=16
+ ad=317 pd=84 as=0 ps=0 
M5385 n_1684 cp1 notdor6 GND efet w=12 l=8
+ ad=852 pd=272 as=190 ps=78 
M5386 idl6 cp1 n_1014 GND efet w=65 l=7
+ ad=1398 pd=342 as=0 ps=0 
M5387 n_1014 dpc42_DL_ADH adh6 GND efet w=43 l=8
+ ad=0 pd=0 as=0 ps=0 
M5388 GND idb6 n_1684 GND efet w=46 l=6
+ ad=0 pd=0 as=0 ps=0 
M5389 dor6 notdor6 GND GND efet w=70 l=6
+ ad=889 pd=252 as=0 ps=0 
M5390 GND notidl6 idl6 GND efet w=37 l=6
+ ad=0 pd=0 as=0 ps=0 
M5391 Vdd n_1638 n_1638 GND dfet w=8 l=7
+ ad=0 pd=0 as=256 ps=98 
M5392 n_1638 cclk notidl6 GND efet w=14 l=8
+ ad=1846 pd=382 as=219 ps=74 
M5393 GND db6 n_1638 GND efet w=133 l=6
+ ad=0 pd=0 as=0 ps=0 
M5394 n_1147 dpc41_DL_ADL adl7 GND efet w=62 l=7
+ ad=2058 pd=510 as=0 ps=0 
M5395 idb6 dpc43_DL_DB n_1014 GND efet w=43 l=7
+ ad=0 pd=0 as=0 ps=0 
M5396 GND notidl6 idl6 GND efet w=34 l=6
+ ad=0 pd=0 as=0 ps=0 
M5397 n_7 RnWstretched GND GND efet w=152 l=6
+ ad=2284 pd=548 as=0 ps=0 
M5398 n_7 RnWstretched GND GND efet w=154 l=6
+ ad=0 pd=0 as=0 ps=0 
M5399 idl6 notidl6 GND GND efet w=50 l=6
+ ad=0 pd=0 as=0 ps=0 
M5400 GND n_466 n_7 GND efet w=138 l=6
+ ad=0 pd=0 as=0 ps=0 
M5401 GND RnWstretched n_466 GND efet w=75 l=7
+ ad=0 pd=0 as=804 ps=214 
M5402 Vdd cclk idb6 GND efet w=22 l=7
+ ad=0 pd=0 as=0 ps=0 
M5403 n_7 dor6 Vdd GND dfet w=17 l=7
+ ad=0 pd=0 as=0 ps=0 
M5404 Vdd n_466 n_466 GND dfet w=8 l=8
+ ad=0 pd=0 as=1550 ps=492 
M5405 n_471 n_466 Vdd GND dfet w=17 l=7
+ ad=2636 pd=552 as=0 ps=0 
M5406 GND RnWstretched n_471 GND efet w=95 l=6
+ ad=0 pd=0 as=0 ps=0 
M5407 db4 n_147 GND GND efet w=214 l=6
+ ad=0 pd=0 as=0 ps=0 
M5408 db4 n_1076 Vdd GND efet w=634 l=7
+ ad=0 pd=0 as=0 ps=0 
M5409 GND n_147 db4 GND efet w=11 l=5
+ ad=0 pd=0 as=0 ps=0 
M5410 db4 n_147 GND GND efet w=215 l=6
+ ad=0 pd=0 as=0 ps=0 
M5411 GND n_147 db4 GND efet w=11 l=5
+ ad=0 pd=0 as=0 ps=0 
M5412 db4 n_147 GND GND efet w=156 l=7
+ ad=0 pd=0 as=0 ps=0 
M5413 db4 n_147 GND GND efet w=228 l=6
+ ad=0 pd=0 as=0 ps=0 
M5414 GND n_612 db5 GND efet w=155 l=7
+ ad=0 pd=0 as=29707 ps=5060 
M5415 GND n_612 db5 GND efet w=228 l=7
+ ad=0 pd=0 as=0 ps=0 
M5416 GND RnWstretched n_471 GND efet w=201 l=6
+ ad=0 pd=0 as=0 ps=0 
M5417 n_471 dor6 GND GND efet w=148 l=6
+ ad=0 pd=0 as=0 ps=0 
M5418 n_466 dor6 GND GND efet w=60 l=6
+ ad=0 pd=0 as=0 ps=0 
M5419 db5 n_373 Vdd GND efet w=637 l=6
+ ad=0 pd=0 as=0 ps=0 
M5420 dor6 dor6 Vdd GND dfet w=10 l=12
+ ad=2151 pd=678 as=0 ps=0 
M5421 db5 n_612 GND GND efet w=213 l=6
+ ad=0 pd=0 as=0 ps=0 
M5422 Vdd n_789 n_789 GND dfet w=9 l=17
+ ad=0 pd=0 as=343 ps=86 
M5423 idl7 idl7 Vdd GND dfet w=9 l=17
+ ad=334 pd=86 as=0 ps=0 
M5424 n_789 cp1 notdor7 GND efet w=12 l=8
+ ad=953 pd=268 as=228 ps=86 
M5425 idl7 cp1 n_1147 GND efet w=65 l=7
+ ad=1351 pd=340 as=0 ps=0 
M5426 n_1147 dpc42_DL_ADH adh7 GND efet w=43 l=7
+ ad=0 pd=0 as=0 ps=0 
M5427 GND idb7 n_789 GND efet w=44 l=6
+ ad=0 pd=0 as=0 ps=0 
M5428 dor7 notdor7 GND GND efet w=69 l=6
+ ad=884 pd=250 as=0 ps=0 
M5429 GND notidl7 idl7 GND efet w=36 l=6
+ ad=0 pd=0 as=0 ps=0 
M5430 Vdd n_588 n_588 GND dfet w=10 l=7
+ ad=0 pd=0 as=256 ps=98 
M5431 GND n_612 db5 GND efet w=13 l=7
+ ad=0 pd=0 as=0 ps=0 
M5432 idb7 dpc43_DL_DB n_1147 GND efet w=44 l=7
+ ad=0 pd=0 as=0 ps=0 
M5433 GND notidl7 idl7 GND efet w=35 l=6
+ ad=0 pd=0 as=0 ps=0 
M5434 n_588 cclk notidl7 GND efet w=14 l=8
+ ad=1760 pd=382 as=211 ps=72 
M5435 GND db7 n_588 GND efet w=134 l=7
+ ad=0 pd=0 as=0 ps=0 
M5436 GND notidl7 idl7 GND efet w=48 l=7
+ ad=0 pd=0 as=0 ps=0 
M5437 n_298 RnWstretched GND GND efet w=152 l=6
+ ad=2245 pd=552 as=0 ps=0 
M5438 n_298 RnWstretched GND GND efet w=157 l=6
+ ad=0 pd=0 as=0 ps=0 
M5439 GND n_23 n_298 GND efet w=138 l=6
+ ad=0 pd=0 as=0 ps=0 
M5440 GND RnWstretched n_23 GND efet w=74 l=6
+ ad=0 pd=0 as=788 ps=214 
M5441 Vdd cclk idb7 GND efet w=23 l=7
+ ad=0 pd=0 as=0 ps=0 
M5442 n_298 dor7 Vdd GND dfet w=16 l=7
+ ad=0 pd=0 as=0 ps=0 
M5443 Vdd n_23 n_23 GND dfet w=9 l=8
+ ad=0 pd=0 as=1602 ps=496 
M5444 n_1501 n_23 Vdd GND dfet w=17 l=7
+ ad=2493 pd=548 as=0 ps=0 
M5445 GND RnWstretched n_1501 GND efet w=95 l=6
+ ad=0 pd=0 as=0 ps=0 
M5446 GND RnWstretched n_1501 GND efet w=199 l=6
+ ad=0 pd=0 as=0 ps=0 
M5447 n_1501 dor7 GND GND efet w=148 l=6
+ ad=0 pd=0 as=0 ps=0 
M5448 n_23 dor7 GND GND efet w=60 l=7
+ ad=0 pd=0 as=0 ps=0 
M5449 dor7 dor7 Vdd GND dfet w=10 l=12
+ ad=2308 pd=674 as=0 ps=0 
M5450 db5 n_612 GND GND efet w=212 l=6
+ ad=0 pd=0 as=0 ps=0 
M5451 db5 n_373 Vdd GND efet w=639 l=6
+ ad=0 pd=0 as=0 ps=0 
M5452 GND n_612 db5 GND efet w=11 l=7
+ ad=0 pd=0 as=0 ps=0 
M5453 GND n_612 db5 GND efet w=232 l=6
+ ad=0 pd=0 as=0 ps=0 
M5454 GND GND db5 GND efet w=54 l=7
+ ad=0 pd=0 as=0 ps=0 
M5455 GND GND db6 GND efet w=56 l=7
+ ad=0 pd=0 as=25581 ps=4358 
M5456 db6 n_7 Vdd GND efet w=146 l=7
+ ad=0 pd=0 as=0 ps=0 
M5457 n_254 n_254 Vdd GND dfet w=10 l=10
+ ad=212 pd=72 as=0 ps=0 
M5458 n_869 abh5 GND GND efet w=148 l=6
+ ad=1167 pd=354 as=0 ps=0 
M5459 Vdd n_1423 n_869 GND dfet w=20 l=7
+ ad=0 pd=0 as=0 ps=0 
M5460 nABH5 cclk n_869 GND efet w=12 l=8
+ ad=405 pd=118 as=0 ps=0 
M5461 n_1353 ADH_ABH nABH5 GND efet w=11 l=8
+ ad=55 pd=32 as=0 ps=0 
M5462 n_254 cp1 n_1353 GND efet w=11 l=7
+ ad=978 pd=240 as=0 ps=0 
M5463 GND adh5 n_254 GND efet w=76 l=6
+ ad=0 pd=0 as=0 ps=0 
M5464 n_880 adh6 GND GND efet w=76 l=7
+ ad=799 pd=246 as=0 ps=0 
M5465 Vdd n_880 n_880 GND dfet w=9 l=9
+ ad=0 pd=0 as=206 ps=70 
M5466 abh6 nABH6 GND GND efet w=66 l=7
+ ad=584 pd=192 as=0 ps=0 
M5467 Vdd abh6 abh6 GND dfet w=9 l=14
+ ad=0 pd=0 as=2126 ps=662 
M5468 GND n_1523 n_963 GND efet w=113 l=6
+ ad=0 pd=0 as=1900 ps=398 
M5469 n_963 abh6 Vdd GND dfet w=17 l=7
+ ad=0 pd=0 as=0 ps=0 
M5470 Vdd n_1523 n_1523 GND dfet w=9 l=10
+ ad=0 pd=0 as=1959 ps=670 
M5471 GND abh6 n_1523 GND efet w=45 l=6
+ ad=0 pd=0 as=509 ps=144 
M5472 n_1514 cp1 n_880 GND efet w=12 l=7
+ ad=60 pd=34 as=0 ps=0 
M5473 nABH6 ADH_ABH n_1514 GND efet w=12 l=8
+ ad=402 pd=110 as=0 ps=0 
M5474 n_635 cclk nABH6 GND efet w=14 l=9
+ ad=1186 pd=358 as=0 ps=0 
M5475 Vdd n_1523 n_635 GND dfet w=20 l=6
+ ad=0 pd=0 as=0 ps=0 
M5476 GND abh6 n_635 GND efet w=147 l=6
+ ad=0 pd=0 as=0 ps=0 
M5477 GND n_869 ab13 GND efet w=41 l=6
+ ad=0 pd=0 as=0 ps=0 
M5478 GND n_869 ab13 GND efet w=13 l=6
+ ad=0 pd=0 as=0 ps=0 
M5479 GND n_869 ab13 GND efet w=163 l=6
+ ad=0 pd=0 as=0 ps=0 
M5480 ab13 n_869 GND GND efet w=163 l=6
+ ad=0 pd=0 as=0 ps=0 
M5481 GND n_869 ab13 GND efet w=164 l=6
+ ad=0 pd=0 as=0 ps=0 
M5482 ab13 n_869 GND GND efet w=164 l=8
+ ad=0 pd=0 as=0 ps=0 
M5483 GND n_869 ab13 GND efet w=164 l=7
+ ad=0 pd=0 as=0 ps=0 
M5484 GND n_635 ab14 GND efet w=13 l=5
+ ad=0 pd=0 as=18651 ps=2324 
M5485 GND n_635 ab14 GND efet w=42 l=5
+ ad=0 pd=0 as=0 ps=0 
M5486 ab14 n_635 GND GND efet w=164 l=6
+ ad=0 pd=0 as=0 ps=0 
M5487 GND n_635 ab14 GND efet w=164 l=7
+ ad=0 pd=0 as=0 ps=0 
M5488 ab14 n_635 GND GND efet w=164 l=6
+ ad=0 pd=0 as=0 ps=0 
M5489 GND n_635 ab14 GND efet w=164 l=6
+ ad=0 pd=0 as=0 ps=0 
M5490 ab14 n_635 GND GND efet w=164 l=6
+ ad=0 pd=0 as=0 ps=0 
M5491 Vdd n_963 ab14 GND efet w=419 l=7
+ ad=0 pd=0 as=0 ps=0 
M5492 Vdd n_963 ab14 GND efet w=317 l=6
+ ad=0 pd=0 as=0 ps=0 
M5493 Vdd n_963 ab14 GND efet w=160 l=7
+ ad=0 pd=0 as=0 ps=0 
M5494 GND n_1153 n_1639 GND efet w=131 l=6
+ ad=0 pd=0 as=2134 ps=430 
M5495 n_494 adh7 GND GND efet w=76 l=7
+ ad=747 pd=234 as=0 ps=0 
M5496 Vdd n_494 n_494 GND dfet w=10 l=10
+ ad=0 pd=0 as=232 ps=74 
M5497 abh7 nABH7 GND GND efet w=67 l=7
+ ad=521 pd=178 as=0 ps=0 
M5498 Vdd abh7 abh7 GND dfet w=10 l=12
+ ad=0 pd=0 as=2007 ps=658 
M5499 n_1639 abh7 Vdd GND dfet w=17 l=6
+ ad=0 pd=0 as=0 ps=0 
M5500 Vdd n_1153 n_1153 GND dfet w=9 l=9
+ ad=0 pd=0 as=1961 ps=666 
M5501 GND abh7 n_1153 GND efet w=47 l=6
+ ad=0 pd=0 as=525 ps=144 
M5502 n_514 cp1 n_494 GND efet w=12 l=7
+ ad=72 pd=36 as=0 ps=0 
M5503 nABH7 ADH_ABH n_514 GND efet w=12 l=7
+ ad=388 pd=120 as=0 ps=0 
M5504 n_659 cclk nABH7 GND efet w=11 l=8
+ ad=1137 pd=368 as=0 ps=0 
M5505 Vdd n_1153 n_659 GND dfet w=19 l=7
+ ad=0 pd=0 as=0 ps=0 
M5506 GND abh7 n_659 GND efet w=148 l=6
+ ad=0 pd=0 as=0 ps=0 
M5507 ab15 n_659 GND GND efet w=178 l=6
+ ad=19416 pd=2334 as=0 ps=0 
M5508 GND n_659 ab15 GND efet w=51 l=6
+ ad=0 pd=0 as=0 ps=0 
M5509 GND n_659 ab15 GND efet w=162 l=6
+ ad=0 pd=0 as=0 ps=0 
M5510 ab15 n_659 GND GND efet w=162 l=6
+ ad=0 pd=0 as=0 ps=0 
M5511 GND n_659 ab15 GND efet w=162 l=6
+ ad=0 pd=0 as=0 ps=0 
M5512 ab15 n_659 GND GND efet w=162 l=7
+ ad=0 pd=0 as=0 ps=0 
M5513 Vdd n_1639 ab15 GND efet w=411 l=6
+ ad=0 pd=0 as=0 ps=0 
M5514 Vdd n_1639 ab15 GND efet w=315 l=6
+ ad=0 pd=0 as=0 ps=0 
M5515 Vdd n_1639 ab15 GND efet w=163 l=6
+ ad=0 pd=0 as=0 ps=0 
M5516 db6 n_471 db6 GND efet w=8 l=6
+ ad=0 pd=0 as=0 ps=0 
M5517 db6 n_7 Vdd GND efet w=470 l=6
+ ad=0 pd=0 as=0 ps=0 
M5518 db6 n_471 GND GND efet w=213 l=6
+ ad=0 pd=0 as=0 ps=0 
M5519 GND n_471 db6 GND efet w=9 l=6
+ ad=0 pd=0 as=0 ps=0 
M5520 db6 n_471 GND GND efet w=211 l=6
+ ad=0 pd=0 as=0 ps=0 
M5521 db6 n_7 Vdd GND efet w=626 l=6
+ ad=0 pd=0 as=0 ps=0 
M5522 GND n_471 db6 GND efet w=11 l=6
+ ad=0 pd=0 as=0 ps=0 
M5523 db6 n_471 GND GND efet w=215 l=6
+ ad=0 pd=0 as=0 ps=0 
M5524 GND n_471 db6 GND efet w=11 l=6
+ ad=0 pd=0 as=0 ps=0 
M5525 db6 n_471 GND GND efet w=150 l=6
+ ad=0 pd=0 as=0 ps=0 
M5526 db6 n_471 GND GND efet w=229 l=6
+ ad=0 pd=0 as=0 ps=0 
M5527 GND GND db7 GND efet w=46 l=7
+ ad=0 pd=0 as=28444 ps=4486 
M5528 Vdd n_298 db7 GND efet w=297 l=6
+ ad=0 pd=0 as=0 ps=0 
M5529 db7 n_1501 GND GND efet w=261 l=6
+ ad=0 pd=0 as=0 ps=0 
M5530 Vdd n_298 db7 GND efet w=293 l=6
+ ad=0 pd=0 as=0 ps=0 
M5531 Vdd n_298 db7 GND efet w=293 l=7
+ ad=0 pd=0 as=0 ps=0 
M5532 Vdd n_298 db7 GND efet w=291 l=7
+ ad=0 pd=0 as=0 ps=0 
M5533 GND n_1501 db7 GND efet w=261 l=5
+ ad=0 pd=0 as=0 ps=0 
M5534 db7 n_1501 GND GND efet w=262 l=6
+ ad=0 pd=0 as=0 ps=0 
M5535 db7 n_1501 GND GND efet w=261 l=6
+ ad=0 pd=0 as=0 ps=0 
C0 metal_3743_71# gnd! 14.4fF ;**FLOATING
C1 metal_3722_71# gnd! 14.4fF ;**FLOATING
C2 metal_3645_77# gnd! 75.6fF ;**FLOATING
C3 metal_3743_108# gnd! 14.4fF ;**FLOATING
C4 metal_3722_96# gnd! 14.4fF ;**FLOATING
C5 metal_252_84# gnd! 85.6fF ;**FLOATING
C6 testpad_8 gnd! 459.4fF ;**FLOATING
C7 metal_1733_2073# gnd! 568.8fF ;**FLOATING
C8 metal_772_2304# gnd! 69.6fF ;**FLOATING
C9 metal_1625_2379# gnd! 453.6fF ;**FLOATING
C10 metal_790_2348# gnd! 31.2fF ;**FLOATING
C11 metal_772_2348# gnd! 34.3fF ;**FLOATING
C12 metal_853_2540# gnd! 99.6fF ;**FLOATING
C13 metal_2585_3058# gnd! 547.2fF ;**FLOATING
C14 pad_nc1 gnd! 1494.7fF ;**FLOATING
C15 diff_3703_71# gnd! 18.8fF ;**FLOATING
C16 diff_3681_71# gnd! 19.8fF ;**FLOATING
C17 n_915 gnd! 81.2fF ;**FLOATING
C18 n_749 gnd! 78.4fF ;**FLOATING
C19 diff_3703_109# gnd! 14.6fF ;**FLOATING
C20 diff_3681_97# gnd! 18.4fF ;**FLOATING
C21 n_1208 gnd! 86.8fF ;**FLOATING
C22 n_908 gnd! 86.8fF ;**FLOATING
C23 n_144 gnd! 303.6fF ;**FLOATING
C24 ab15 gnd! 11093.3fF
C25 n_659 gnd! 1828.6fF
C26 n_514 gnd! 36.0fF
C27 n_1639 gnd! 2254.2fF
C28 abh7 gnd! 735.6fF
C29 n_494 gnd! 412.0fF
C30 n_1153 gnd! 648.2fF
C31 nABH7 gnd! 329.0fF
C32 ab14 gnd! 10567.1fF
C33 n_635 gnd! 1795.2fF
C34 n_1514 gnd! 30.8fF
C35 n_963 gnd! 2193.4fF
C36 n_1523 gnd! 649.8fF
C37 abh6 gnd! 785.6fF
C38 n_1353 gnd! 28.4fF
C39 n_869 gnd! 1883.8fF
C40 n_880 gnd! 424.8fF
C41 nABH6 gnd! 327.4fF
C42 n_1501 gnd! 3203.1fF
C43 n_23 gnd! 690.2fF
C44 n_298 gnd! 3286.8fF
C45 n_588 gnd! 840.4fF
C46 dor7 gnd! 969.4fF
C47 notdor7 gnd! 224.4fF
C48 n_789 gnd! 517.8fF
C49 notidl7 gnd! 363.6fF
C50 idl7 gnd! 683.6fF
C51 n_471 gnd! 3199.9fF
C52 n_466 gnd! 690.6fF
C53 n_7 gnd! 3429.9fF
C54 n_1147 gnd! 1112.4fF
C55 n_1638 gnd! 876.4fF
C56 dor6 gnd! 925.6fF
C57 notdor6 gnd! 206.8fF
C58 n_1684 gnd! 478.2fF
C59 notidl6 gnd! 369.2fF
C60 idl6 gnd! 701.0fF
C61 n_612 gnd! 2847.4fF
C62 n_1720 gnd! 652.8fF
C63 n_373 gnd! 3295.0fF
C64 n_542 gnd! 2666.7fF ;**FLOATING
C65 n_1014 gnd! 1090.2fF
C66 n_568 gnd! 879.6fF
C67 dor5 gnd! 978.2fF
C68 notdor5 gnd! 221.2fF
C69 n_961 gnd! 478.2fF
C70 notidl5 gnd! 389.6fF
C71 idl5 gnd! 688.4fF
C72 n_147 gnd! 3008.8fF
C73 n_1463 gnd! 669.6fF
C74 n_1076 gnd! 3257.8fF
C75 n_254 gnd! 494.8fF
C76 ab13 gnd! 10399.4fF
C77 ab12 gnd! 10603.2fF
C78 n_999 gnd! 1809.8fF
C79 n_1451 gnd! 25.6fF
C80 n_1608 gnd! 2100.4fF
C81 n_475 gnd! 2105.8fF
C82 abh5 gnd! 809.4fF
C83 nABH5 gnd! 334.2fF
C84 n_1423 gnd! 668.6fF
C85 n_1677 gnd! 704.4fF
C86 abh4 gnd! 767.2fF
C87 n_212 gnd! 432.6fF
C88 nABH4 gnd! 327.0fF
C89 n_1667 gnd! 28.4fF
C90 n_359 gnd! 1842.6fF
C91 n_883 gnd! 488.0fF
C92 nABH3 gnd! 311.6fF
C93 ab11 gnd! 10480.6fF
C94 ab10 gnd! 10617.8fF
C95 n_994 gnd! 1870.2fF
C96 n_836 gnd! 30.8fF
C97 n_1296 gnd! 2192.0fF
C98 n_1545 gnd! 2179.8fF
C99 abh3 gnd! 826.6fF
C100 n_1346 gnd! 609.0fF
C101 n_1034 gnd! 632.6fF
C102 abh2 gnd! 760.2fF
C103 n_1298 gnd! 36.0fF
C104 n_676 gnd! 1860.6fF
C105 n_168 gnd! 449.6fF
C106 nABH2 gnd! 326.6fF
C107 n_1387 gnd! 1101.0fF
C108 n_490 gnd! 840.2fF
C109 dor4 gnd! 923.6fF
C110 notdor4 gnd! 207.4fF
C111 n_797 gnd! 475.8fF
C112 notidl4 gnd! 381.0fF
C113 idl4 gnd! 662.6fF
C114 n_643 gnd! 2831.3fF
C115 n_1613 gnd! 658.4fF
C116 n_42 gnd! 3270.1fF
C117 n_1095 gnd! 1098.0fF
C118 n_896 gnd! 839.8fF
C119 dor3 gnd! 959.2fF
C120 notdor3 gnd! 221.2fF
C121 n_457 gnd! 516.8fF
C122 notidl3 gnd! 366.6fF
C123 idl3 gnd! 664.0fF
C124 n_37 gnd! 2990.2fF
C125 n_224 gnd! 682.2fF
C126 n_520 gnd! 3093.2fF
C127 n_1661 gnd! 1073.4fF
C128 n_1199 gnd! 829.6fF
C129 dor2 gnd! 949.8fF
C130 notdor2 gnd! 219.4fF
C131 n_1376 gnd! 492.0fF
C132 notidl2 gnd! 355.4fF
C133 idl2 gnd! 685.2fF
C134 n_794 gnd! 2947.2fF
C135 n_288 gnd! 663.8fF
C136 n_798 gnd! 3086.7fF
C137 n_1424 gnd! 1115.3fF
C138 n_213 gnd! 874.0fF
C139 dor1 gnd! 915.8fF
C140 pclp7 gnd! 876.2fF
C141 n_914 gnd! 544.8fF
C142 n_484 gnd! 586.4fF
C143 npclp7 gnd! 255.4fF
C144 n_1386 gnd! 468.6fF
C145 n_426 gnd! 216.8fF
C146 pcl7 gnd! 527.8fF
C147 n_641 gnd! 477.2fF
C148 notdor1 gnd! 228.2fF
C149 notidl1 gnd! 385.4fF
C150 idl1 gnd! 680.0fF
C151 n_1474 gnd! 471.0fF
C152 n_769 gnd! 669.0fF
C153 n_87 gnd! 1065.8fF
C154 n_1325 gnd! 3070.4fF
C155 n_1072 gnd! 2839.4fF
C156 n_718 gnd! 830.0fF
C157 dor0 gnd! 911.6fF
C158 notdor0 gnd! 219.8fF
C159 n_1687 gnd! 493.2fF
C160 notidl0 gnd! 364.4fF
C161 idl0 gnd! 702.2fF
C162 n_715 gnd! 888.6fF
C163 pcl6 gnd! 464.2fF
C164 n_993 gnd! 169.0fF
C165 n_1264 gnd! 125.6fF
C166 n_663 gnd! 166.4fF
C167 n_1213 gnd! 712.6fF
C168 n_453 gnd! 672.2fF
C169 n_1209 gnd! 483.6fF
C170 npchp7 gnd! 643.0fF
C171 pchp7 gnd! 939.0fF
C172 n_1316 gnd! 969.4fF
C173 pclp6 gnd! 944.9fF
C174 npclp6 gnd! 601.2fF
C175 n_585 gnd! 95.6fF
C176 n_20 gnd! 516.6fF
C177 n_232 gnd! 785.6fF
C178 pclp5 gnd! 887.9fF
C179 n_557 gnd! 553.2fF
C180 n_1547 gnd! 552.4fF
C181 n_278 gnd! 358.4fF
C182 n_545 gnd! 193.6fF
C183 n_1192 gnd! 589.6fF
C184 npchp6 gnd! 239.4fF
C185 n_609 gnd! 667.2fF
C186 n_1488 gnd! 851.2fF
C187 n_1073 gnd! 626.8fF
C188 npclp5 gnd! 241.2fF
C189 n_344 gnd! 694.0fF
C190 n_814 gnd! 194.0fF
C191 pcl5 gnd! 543.9fF
C192 n_386 gnd! 436.2fF
C193 pch7 gnd! 542.2fF
C194 pchp6 gnd! 901.4fF
C195 pch6 gnd! 617.8fF
C196 n_1659 gnd! 125.6fF
C197 n_469 gnd! 171.6fF
C198 n_743 gnd! 934.6fF
C199 n_499 gnd! 787.0fF
C200 n_875 gnd! 486.2fF
C201 npchp5 gnd! 614.8fF
C202 n_392 gnd! 894.9fF
C203 pcl4 gnd! 459.2fF
C204 n_15 gnd! 158.4fF
C205 n_410 gnd! 942.6fF
C206 pclp4 gnd! 900.2fF
C207 npclp4 gnd! 602.4fF
C208 n_766 gnd! 111.6fF
C209 n_474 gnd! 492.2fF
C210 n_1643 gnd! 771.6fF
C211 pclp3 gnd! 882.2fF
C212 n_903 gnd! 588.0fF
C213 n_1631 gnd! 634.8fF
C214 npclp3 gnd! 244.0fF
C215 n_1184 gnd! 698.2fF
C216 n_1498 gnd! 210.0fF
C217 pcl3 gnd! 540.2fF
C218 n_249 gnd! 502.0fF
C219 n_719 gnd! 1087.7fF
C220 n_1585 gnd! 390.4fF
C221 RnWstretched gnd! 11409.0fF
C222 n_221 gnd! 925.3fF
C223 n_1028 gnd! 523.0fF
C224 n_251 gnd! 1997.0fF
C225 n_962 gnd! 560.2fF
C226 n_1579 gnd! 225.4fF
C227 nDBE gnd! 1032.0fF
C228 n_1293 gnd! 824.2fF
C229 n_802 gnd! 127.6fF
C230 n_1371 gnd! 765.4fF
C231 n_201 gnd! 1031.4fF
C232 p1 gnd! 232.8fF
C233 n_661 gnd! 368.0fF
C234 n_163 gnd! 898.5fF
C235 pcl2 gnd! 466.6fF
C236 n_1411 gnd! 169.8fF
C237 n_1253 gnd! 910.6fF
C238 pclp2 gnd! 934.2fF
C239 npclp2 gnd! 639.0fF
C240 n_1158 gnd! 95.6fF
C241 n_515 gnd! 503.8fF
C242 pchp5 gnd! 903.3fF
C243 n_1406 gnd! 544.0fF
C244 n_1400 gnd! 354.8fF
C245 n_949 gnd! 205.2fF
C246 n_1657 gnd! 601.6fF
C247 npchp4 gnd! 225.0fF
C248 n_523 gnd! 669.2fF
C249 n_83 gnd! 910.4fF
C250 pch5 gnd! 552.4fF
C251 pchp4 gnd! 902.4fF
C252 n_356 gnd! 143.6fF
C253 n_1061 gnd! 173.4fF
C254 n_810 gnd! 674.4fF
C255 n_923 gnd! 757.4fF
C256 n_207 gnd! 490.0fF
C257 npchp3 gnd! 641.2fF
C258 pch4 gnd! 637.5fF
C259 pchp3 gnd! 930.1fF
C260 pch3 gnd! 533.9fF
C261 n_783 gnd! 770.6fF
C262 pclp1 gnd! 877.2fF
C263 n_1568 gnd! 552.8fF
C264 n_1099 gnd! 609.6fF
C265 npclp1 gnd! 250.4fF
C266 n_1542 gnd! 725.6fF
C267 n_1685 gnd! 209.6fF
C268 pcl1 gnd! 540.2fF
C269 n_329 gnd! 456.2fF
C270 n_57 gnd! 564.4fF
C271 n_1265 gnd! 438.4fF
C272 adh7 gnd! 2142.8fF
C273 pchp2 gnd! 880.3fF
C274 n_1402 gnd! 470.4fF
C275 npchp2 gnd! 184.4fF
C276 n_1367 gnd! 196.4fF
C277 n_293 gnd! 679.6fF
C278 n_1166 gnd! 905.8fF
C279 pcl0 gnd! 488.5fF
C280 n_526 gnd! 168.4fF
C281 n_1345 gnd! 936.4fF
C282 pclp0 gnd! 909.3fF
C283 npclp0 gnd! 580.8fF
C284 n_1706 gnd! 98.0fF
C285 n_1500 gnd! 491.4fF
C286 n_937 gnd! 768.4fF
C287 n_580 gnd! 189.2fF
C288 n_566 gnd! 895.8fF
C289 pipeUNK14 gnd! 225.2fF
C290 n_1170 gnd! 490.2fF
C291 nDBZ gnd! 785.2fF
C292 n_1115 gnd! 457.8fF
C293 n_922 gnd! 196.4fF
C294 n_620 gnd! 1338.0fF
C295 n_1433 gnd! 810.8fF
C296 pipeUNK15 gnd! 213.8fF
C297 n_243 gnd! 1092.0fF
C298 DBZ gnd! 1742.7fF
C299 dpc43_DL_DB gnd! 2350.4fF
C300 n_1202 gnd! 900.0fF
C301 pch2 gnd! 675.0fF
C302 n_1538 gnd! 122.8fF
C303 n_126 gnd! 168.8fF
C304 n_200 gnd! 944.6fF
C305 n_1070 gnd! 800.0fF
C306 n_1486 gnd! 474.4fF
C307 npchp1 gnd! 614.6fF
C308 n_835 gnd! 594.0fF
C309 adh6 gnd! 2462.2fF
C310 n_128 gnd! 565.8fF
C311 n_1592 gnd! 820.6fF
C312 n_569 gnd! 88.4fF
C313 n_260 gnd! 504.6fF
C314 a7 gnd! 300.8fF
C315 adh5 gnd! 2608.2fF
C316 n_1356 gnd! 555.8fF
C317 n_1454 gnd! 103.2fF
C318 n_100 gnd! 137.6fF
C319 n_1205 gnd! 793.8fF
C320 n_852 gnd! 454.4fF
C321 dasb7 gnd! 400.6fF
C322 n_1018 gnd! 443.6fF
C323 n_711 gnd! 97.6fF
C324 n_1080 gnd! 86.0fF
C325 n_479 gnd! 503.6fF
C326 n_326 gnd! 868.7fF
C327 a6 gnd! 327.4fF
C328 adh4 gnd! 3889.8fF
C329 n_1719 gnd! 540.2fF
C330 n_1554 gnd! 103.2fF
C331 n_739 gnd! 783.3fF
C332 n_61 gnd! 455.8fF
C333 dasb6 gnd! 388.8fF
C334 n_1056 gnd! 388.0fF
C335 n_1629 gnd! 483.4fF
C336 n_831 gnd! 875.9fF
C337 a5 gnd! 327.2fF
C338 adh3 gnd! 3615.8fF
C339 n_556 gnd! 568.2fF
C340 n_1344 gnd! 851.9fF
C341 n_1203 gnd! 135.2fF
C342 n_408 gnd! 439.4fF
C343 n_1267 gnd! 478.4fF
C344 ab9 gnd! 10415.9fF
C345 diff_272_79# gnd! 79.6fF ;**FLOATING
C346 diff_247_79# gnd! 74.0fF ;**FLOATING
C347 diff_272_107# gnd! 64.4fF ;**FLOATING
C348 n_290 gnd! 59.6fF ;**FLOATING
C349 n_1461 gnd! 69.6fF ;**FLOATING
C350 diff_247_120# gnd! 66.8fF ;**FLOATING
C351 diff_272_148# gnd! 67.6fF ;**FLOATING
C352 diff_247_140# gnd! 65.2fF ;**FLOATING
C353 diff_272_161# gnd! 67.6fF ;**FLOATING
C354 diff_247_161# gnd! 65.2fF ;**FLOATING
C355 diff_272_189# gnd! 67.6fF ;**FLOATING
C356 n_30 gnd! 65.2fF ;**FLOATING
C357 ab8 gnd! 10314.2fF
C358 n_381 gnd! 1948.4fF
C359 ab7 gnd! 11349.6fF
C360 n_705 gnd! 33.2fF
C361 n_826 gnd! 2150.8fF
C362 n_1140 gnd! 2161.4fF
C363 abh1 gnd! 846.4fF
C364 nABH1 gnd! 335.2fF
C365 n_617 gnd! 630.4fF
C366 n_1315 gnd! 718.6fF
C367 alu7 gnd! 655.4fF
C368 notalu7 gnd! 281.2fF
C369 n_762 gnd! 785.0fF
C370 n_1135 gnd! 852.8fF
C371 dasb5 gnd! 391.8fF
C372 n_970 gnd! 184.8fF
C373 n_149 gnd! 601.4fF
C374 n_233 gnd! 1063.6fF
C375 n_761 gnd! 1039.1fF
C376 n_838 gnd! 500.6fF
C377 a4 gnd! 295.2fF
C378 n_753 gnd! 750.8fF
C379 n_811 gnd! 1243.4fF
C380 n_947 gnd! 557.8fF
C381 n_581 gnd! 183.4fF
C382 n_306 gnd! 454.4fF
C383 n_393 gnd! 161.4fF
C384 n_551 gnd! 595.2fF
C385 n_1279 gnd! 111.6fF
C386 n_1097 gnd! 476.0fF
C387 n_1654 gnd! 923.1fF
C388 a3 gnd! 316.8fF
C389 pchp1 gnd! 942.9fF
C390 pch1 gnd! 528.4fF
C391 n_1010 gnd! 422.0fF
C392 pchp0 gnd! 854.0fF
C393 n_1229 gnd! 519.0fF
C394 npchp0 gnd! 200.4fF
C395 n_856 gnd! 213.6fF
C396 n_919 gnd! 686.6fF
C397 pch0 gnd! 614.6fF
C398 n_311 gnd! 890.8fF
C399 adh1 gnd! 4233.2fF
C400 n_419 gnd! 554.4fF
C401 n_1686 gnd! 83.6fF
C402 n_1584 gnd! 132.4fF
C403 n_1179 gnd! 716.6fF
C404 n_345 gnd! 759.3fF
C405 n_432 gnd! 650.2fF
C406 dasb3 gnd! 417.0fF
C407 n_1159 gnd! 435.0fF
C408 n_1618 gnd! 904.7fF
C409 a2 gnd! 301.2fF
C410 n_1656 gnd! 101.6fF
C411 n_1580 gnd! 491.4fF
C412 dasb2 gnd! 442.6fF
C413 n_1549 gnd! 541.0fF
C414 n_929 gnd! 871.4fF
C415 n_619 gnd! 133.2fF
C416 n_695 gnd! 495.8fF
C417 n_735 gnd! 456.2fF
C418 a1 gnd! 303.4fF
C419 n_1322 gnd! 100.4fF
C420 n_320 gnd! 443.0fF
C421 dasb1 gnd! 420.2fF
C422 n_5 gnd! 565.4fF
C423 a0 gnd! 280.8fF
C424 dpc41_DL_ADL gnd! 2700.9fF
C425 dpc42_DL_ADH gnd! 2581.2fF
C426 Pout1 gnd! 625.2fF
C427 Pout0 gnd! 643.4fF
C428 n_318 gnd! 1704.0fF
C429 n_846 gnd! 1018.3fF
C430 n_1625 gnd! 226.6fF
C431 n_307 gnd! 910.8fF
C432 pipeUNK05 gnd! 282.0fF
C433 n_1616 gnd! 237.2fF
C434 n_69 gnd! 216.6fF
C435 n_1445 gnd! 78.8fF
C436 n_1546 gnd! 92.0fF
C437 n_1470 gnd! 92.0fF
C438 pipeUNK13 gnd! 205.6fF
C439 n_793 gnd! 249.0fF
C440 n_1595 gnd! 400.6fF
C441 n_1181 gnd! 842.8fF
C442 n_1614 gnd! 994.2fF
C443 pipeUNK03 gnd! 366.4fF
C444 n_1723 gnd! 256.8fF
C445 n_1177 gnd! 257.4fF
C446 n_299 gnd! 999.2fF
C447 n_648 gnd! 130.4fF
C448 n_1644 gnd! 305.4fF
C449 n_1457 gnd! 656.4fF
C450 n_1495 gnd! 819.1fF
C451 p3 gnd! 213.8fF
C452 pipeUNK04 gnd! 280.0fF
C453 db6 gnd! 17512.5fF
C454 db2 gnd! 15679.1fF
C455 n_1492 gnd! 884.0fF
C456 db0 gnd! 20891.1fF
C457 db5 gnd! 18618.8fF
C458 pipeUNK02 gnd! 148.8fF
C459 p4 gnd! 777.6fF
C460 n_1471 gnd! 514.2fF
C461 p0 gnd! 212.4fF
C462 n_455 gnd! 173.2fF
C463 p6 gnd! 606.4fF
C464 n_1240 gnd! 440.0fF
C465 n_1441 gnd! 489.8fF
C466 n_1157 gnd! 426.0fF
C467 dpc35_PCHC gnd! 2545.6fF
C468 H1x1 gnd! 1589.9fF
C469 n_1416 gnd! 1605.7fF
C470 n_1600 gnd! 1267.8fF
C471 n_90 gnd! 1519.6fF
C472 p7 gnd! 596.0fF
C473 Pout2 gnd! 605.6fF
C474 n_1566 gnd! 601.2fF
C475 dpc40_ADLPCL gnd! 2790.4fF
C476 dpc38_PCLADL gnd! 2513.2fF
C477 dpc39_PCLPCL gnd! 2627.7fF
C478 dpc32_PCHADH gnd! 2302.6fF
C479 n_146 gnd! 913.0fF
C480 n_1341 gnd! 213.2fF
C481 n_876 gnd! 634.4fF
C482 n_1362 gnd! 218.4fF
C483 n_600 gnd! 1427.1fF
C484 n_150 gnd! 174.4fF
C485 n_613 gnd! 1148.8fF
C486 n_867 gnd! 718.3fF
C487 n_8 gnd! 1152.0fF
C488 n_1682 gnd! 336.0fF
C489 n_986 gnd! 958.6fF
C490 n_1556 gnd! 107.2fF
C491 nDA_ADD2 gnd! 676.4fF
C492 nDA_ADD1 gnd! 775.9fF
C493 notalu6 gnd! 256.2fF
C494 alu6 gnd! 970.8fF
C495 C78 gnd! 562.0fF
C496 C78_phi2 gnd! 155.6fF
C497 DC78_phi2 gnd! 162.8fF
C498 notaluvout gnd! 650.8fF
C499 adh2 gnd! 4487.3fF
C500 n_637 gnd! 520.0fF
C501 n_1489 gnd! 256.4fF
C502 notalu5 gnd! 266.0fF
C503 alu5 gnd! 989.0fF
C504 notalu4 gnd! 260.6fF
C505 alu4 gnd! 810.2fF
C506 notalu3 gnd! 256.8fF
C507 alu3 gnd! 782.0fF
C508 notalu2 gnd! 252.4fF
C509 alu2 gnd! 1067.8fF
C510 dpc37_PCLDB gnd! 2233.7fF
C511 n_1007 gnd! 399.0fF
C512 dpc34_PCLC gnd! 4407.3fF
C513 n_1043 gnd! 455.2fF
C514 n_1462 gnd! 430.4fF
C515 dpc33_PCHDB gnd! 2164.9fF
C516 n_36 gnd! 799.6fF
C517 n_1277 gnd! 603.0fF
C518 n_291 gnd! 667.2fF
C519 n_1221 gnd! 223.8fF
C520 n_1020 gnd! 222.2fF
C521 n_1121 gnd! 217.4fF
C522 n_1045 gnd! 2216.3fF
C523 n_186 gnd! 76.4fF
C524 n_367 gnd! 156.8fF
C525 n_1224 gnd! 968.2fF
C526 pipeUNK16 gnd! 303.2fF
C527 n_756 gnd! 350.2fF
C528 n_1110 gnd! 1157.0fF
C529 n_626 gnd! 575.4fF
C530 pipeUNK12 gnd! 178.2fF
C531 n_1198 gnd! 273.6fF
C532 n_1249 gnd! 332.4fF
C533 pipeUNK01 gnd! 201.2fF
C534 n_755 gnd! 1304.3fF
C535 n_1692 gnd! 93.6fF
C536 n_1082 gnd! 1394.6fF
C537 n_279 gnd! 804.2fF
C538 n_507 gnd! 542.0fF
C539 n_1049 gnd! 198.0fF
C540 n_1194 gnd! 1496.7fF
C541 n_160 gnd! 553.8fF
C542 db4 gnd! 17619.4fF
C543 n_374 gnd! 714.8fF
C544 n_111 gnd! 703.4fF
C545 n_62 gnd! 681.6fF
C546 db7 gnd! 19610.5fF
C547 db1 gnd! 21502.0fF
C548 n_1319 gnd! 711.4fF
C549 n_93 gnd! 754.8fF
C550 n_1588 gnd! 748.6fF
C551 n_1281 gnd! 703.4fF
C552 db3 gnd! 17055.4fF
C553 n_1075 gnd! 702.4fF
C554 n_587 gnd! 1060.8fF
C555 n_503 gnd! 380.0fF
C556 n_340 gnd! 371.6fF
C557 pd4 gnd! 252.6fF
C558 n_1214 gnd! 462.6fF
C559 n_1401 gnd! 540.4fF
C560 n_1269 gnd! 325.4fF
C561 DBNeg gnd! 2209.8fF
C562 n_1673 gnd! 174.4fF
C563 n_754 gnd! 1846.0fF
C564 n_1422 gnd! 245.6fF
C565 pipeUNK06 gnd! 357.4fF
C566 n_1111 gnd! 1459.0fF
C567 pipeUNK11 gnd! 221.8fF
C568 pipeUNK07 gnd! 199.4fF
C569 n_941 gnd! 229.6fF
C570 pipeUNK09 gnd! 786.9fF
C571 n_954 gnd! 1498.7fF
C572 pipeUNK08 gnd! 246.4fF
C573 n_818 gnd! 651.4fF
C574 n_1518 gnd! 436.2fF
C575 n_1413 gnd! 431.6fF
C576 dpc31_PCHPCH gnd! 2516.0fF
C577 n_1323 gnd! 409.4fF
C578 n_849 gnd! 431.4fF
C579 dpc30_ADHPCH gnd! 2594.2fF
C580 n_AxB7__C67 gnd! 389.2fF
C581 DC78 gnd! 767.8fF
C582 n_AxBxC_7 gnd! 487.8fF
C583 n_1013 gnd! 86.0fF
C584 n_AxB_7 gnd! 316.4fF
C585 nC78 gnd! 662.6fF
C586 n_1617 gnd! 142.4fF
C587 n_1030 gnd! 819.6fF
C588 nC67 gnd! 383.0fF
C589 n_269 gnd! 510.2fF
C590 AxB7 gnd! 1046.9fF
C591 A_B7 gnd! 484.8fF
C592 n_748 gnd! 660.0fF
C593 n_A_B_7 gnd! 1215.8fF
C594 naluresult7 gnd! 1141.0fF
C595 _AxB_6_nC56 gnd! 445.4fF
C596 n_1038 gnd! 359.8fF
C597 n_AxBxC_6 gnd! 482.4fF
C598 n_1390 gnd! 86.0fF
C599 n_112 gnd! 155.2fF
C600 C67 gnd! 1015.8fF
C601 n_482 gnd! 97.6fF
C602 n_AxB_6 gnd! 1079.2fF
C603 C56 gnd! 421.4fF
C604 nA_B7 gnd! 1153.4fF
C605 n_1695 gnd! 173.2fF
C606 alua7 gnd! 456.0fF
C607 n_423 gnd! 530.6fF
C608 idb7 gnd! 4875.8fF
C609 alub7 gnd! 696.9fF
C610 n_A_B_6 gnd! 946.7fF
C611 naluresult6 gnd! 1424.3fF
C612 A_B6 gnd! 426.8fF
C613 n_570 gnd! 1102.7fF
C614 n_AxB5__C45 gnd! 412.2fF
C615 n_122 gnd! 518.8fF
C616 n_1257 gnd! 1617.6fF
C617 n_AxBxC_5 gnd! 498.8fF
C618 n_547 gnd! 100.4fF
C619 n_AxB_5 gnd! 315.2fF
C620 nC56 gnd! 672.6fF
C621 n_165 gnd! 155.2fF
C622 AxB5 gnd! 899.0fF
C623 n_939 gnd! 172.4fF
C624 n_757 gnd! 987.0fF
C625 notalucout gnd! 1286.0fF
C626 alucout gnd! 3193.0fF
C627 A_B5 gnd! 460.8fF
C628 n_647 gnd! 1031.2fF
C629 nC45 gnd! 671.8fF
C630 _AxB_4_nC34 gnd! 441.2fF
C631 DA_C45 gnd! 520.2fF
C632 n_AxBxC_4 gnd! 516.8fF
C633 n_375 gnd! 100.4fF
C634 n_1310 gnd! 134.4fF
C635 C45 gnd! 635.4fF
C636 n_1583 gnd! 94.8fF
C637 nA_B6 gnd! 1347.4fF
C638 n_1483 gnd! 173.2fF
C639 alua6 gnd! 448.6fF
C640 n_351 gnd! 524.6fF
C641 idb6 gnd! 4804.6fF
C642 alub6 gnd! 687.9fF
C643 s7 gnd! 285.0fF
C644 nots7 gnd! 214.4fF
C645 n_548 gnd! 506.8fF
C646 n_721 gnd! 1090.8fF
C647 n_A_B_5 gnd! 923.4fF
C648 naluresult5 gnd! 1514.7fF
C649 nA_B5 gnd! 870.2fF
C650 n_1559 gnd! 148.4fF
C651 alua5 gnd! 465.8fF
C652 n_AxB_4 gnd! 750.2fF
C653 n_1218 gnd! 579.8fF
C654 C34 gnd! 1083.4fF
C655 n_1565 gnd! 219.2fF
C656 n_700 gnd! 920.3fF
C657 notalu1 gnd! 266.0fF
C658 alu1 gnd! 1007.4fF
C659 notalu0 gnd! 262.2fF
C660 alu0 gnd! 819.0fF
C661 n_972 gnd! 762.4fF
C662 n_1383 gnd! 521.8fF
C663 idb5 gnd! 4500.4fF
C664 alub5 gnd! 669.6fF
C665 n_A_B_4 gnd! 939.5fF
C666 naluresult4 gnd! 1392.6fF
C667 A_B4 gnd! 425.4fF
C668 DC34 gnd! 875.4fF
C669 n_AxB3__C23 gnd! 417.2fF
C670 n_AxBxC_3 gnd! 482.6fF
C671 n_136 gnd! 100.4fF
C672 nC34 gnd! 746.2fF
C673 n_924 gnd! 150.8fF
C674 n_AxB_3 gnd! 323.6fF
C675 nC23 gnd! 398.2fF
C676 A_B3 gnd! 459.2fF
C677 n_988 gnd! 657.4fF
C678 nA_B4 gnd! 1063.0fF
C679 n_185 gnd! 173.2fF
C680 alua4 gnd! 429.4fF
C681 n_478 gnd! 500.6fF
C682 idb4 gnd! 4430.1fF
C683 alub4 gnd! 666.6fF
C684 n_A_B_3 gnd! 963.3fF
C685 naluresult3 gnd! 1547.7fF
C686 _AxB_2_nC12 gnd! 503.8fF
C687 n_1610 gnd! 763.0fF
C688 AxB3 gnd! 1217.0fF
C689 DA_AB2 gnd! 826.4fF
C690 n_AxBxC_2 gnd! 535.2fF
C691 n_1572 gnd! 103.2fF
C692 n_433 gnd! 232.4fF
C693 C23 gnd! 691.2fF
C694 n_716 gnd! 95.6fF
C695 n_AxB_2 gnd! 702.6fF
C696 nA_B3 gnd! 884.0fF
C697 n_313 gnd! 173.2fF
C698 alua3 gnd! 451.2fF
C699 n_1621 gnd! 506.6fF
C700 idb3 gnd! 4368.3fF
C701 alub3 gnd! 661.8fF
C702 n_A_B_2 gnd! 1520.7fF
C703 naluresult2 gnd! 1415.6fF
C704 C12 gnd! 354.4fF
C705 A_B2 gnd! 328.6fF
C706 n_AxB1__C01 gnd! 407.4fF
C707 DA_AxB2 gnd! 780.2fF
C708 n_388 gnd! 1309.0fF
C709 n_AxBxC_1 gnd! 491.0fF
C710 n_1388 gnd! 100.4fF
C711 n_AxB_1 gnd! 313.6fF
C712 nC12 gnd! 686.0fF
C713 n_1510 gnd! 150.4fF
C714 n_1354 gnd! 129.2fF
C715 n_319 gnd! 1066.1fF
C716 n_1707 gnd! 153.6fF
C717 AxB1 gnd! 916.4fF
C718 nC01 gnd! 377.4fF
C719 n_936 gnd! 1036.4fF
C720 A_B1 gnd! 456.6fF
C721 _AxB_0_nC0in gnd! 512.2fF
C722 DA_C01 gnd! 723.8fF
C723 dpc26_ACDB gnd! 2650.2fF
C724 n_1369 gnd! 641.8fF
C725 n_1270 gnd! 671.8fF
C726 n_1260 gnd! 612.0fF
C727 n_255 gnd! 404.8fF
C728 n_631 gnd! 638.0fF
C729 n_228 gnd! 431.4fF
C730 dpc24_ACSB gnd! 2289.2fF
C731 dpc29_0ADH17 gnd! 2517.6fF
C732 dpc27_SBADH gnd! 2132.6fF
C733 n_800 gnd! 415.2fF
C734 n_321 gnd! 615.8fF
C735 n_1335 gnd! 395.6fF
C736 dpc23_SBAC gnd! 2323.2fF
C737 dpc25_SBDB gnd! 2380.1fF
C738 n_1635 gnd! 414.6fF
C739 n_265 gnd! 181.6fF
C740 n_897 gnd! 215.6fF
C741 n_611 gnd! 663.2fF
C742 n_21 gnd! 683.2fF
C743 n_525 gnd! 676.8fF
C744 n_598 gnd! 222.6fF
C745 n_878 gnd! 231.8fF
C746 n_509 gnd! 163.6fF
C747 n_398 gnd! 227.2fF
C748 n_1509 gnd! 172.4fF
C749 n_1162 gnd! 168.8fF
C750 n_266 gnd! 170.8fF
C751 n_1271 gnd! 428.2fF
C752 n_628 gnd! 617.2fF
C753 n_1047 gnd! 414.2fF
C754 n_1238 gnd! 435.8fF
C755 n_966 gnd! 630.8fF
C756 n_1596 gnd! 647.4fF
C757 n_830 gnd! 675.0fF
C758 n_1295 gnd! 653.0fF
C759 n_55 gnd! 183.2fF
C760 n_1683 gnd! 215.6fF
C761 n_1602 gnd! 206.8fF
C762 n_1505 gnd! 181.4fF
C763 n_1527 gnd! 222.2fF
C764 n_1581 gnd! 318.4fF
C765 n_1480 gnd! 1485.4fF
C766 dpc36_nIPC gnd! 1439.6fF
C767 n_1275 gnd! 796.6fF
C768 n_1570 gnd! 307.8fF
C769 n_1472 gnd! 367.2fF
C770 pipeBRtaken gnd! 374.8fF
C771 n_1446 gnd! 575.4fF
C772 n_465 gnd! 576.4fF
C773 pipeUNK20 gnd! 324.4fF
C774 n_850 gnd! 635.8fF
C775 short_circuit_branch_add gnd! 1166.4fF
C776 n_323 gnd! 172.8fF
C777 n_1550 gnd! 158.4fF
C778 pipeUNK18 gnd! 252.0fF
C779 n_771 gnd! 1536.8fF
C780 n_959 gnd! 968.0fF
C781 n_671 gnd! 180.0fF
C782 n_1573 gnd! 1094.4fF
C783 n_511 gnd! 234.0fF
C784 pipeUNK17 gnd! 240.4fF
C785 n_270 gnd! 3283.9fF
C786 n_1426 gnd! 290.4fF
C787 n_513 gnd! 623.8fF
C788 pd6 gnd! 350.0fF
C789 pd2 gnd! 300.0fF
C790 pd7 gnd! 285.2fF
C791 pd1 gnd! 264.4fF
C792 pd0 gnd! 299.0fF
C793 pd5 gnd! 274.6fF
C794 pd3 gnd! 273.8fF
C795 clearIR gnd! 1491.2fF
C796 n_380 gnd! 159.2fF
C797 n_1662 gnd! 842.2fF
C798 n_553 gnd! 839.6fF
C799 n_845 gnd! 980.2fF
C800 p2 gnd! 235.4fF
C801 n_31 gnd! 3174.0fF
C802 n_24 gnd! 335.6fF
C803 n_1528 gnd! 341.8fF
C804 n_106 gnd! 465.6fF
C805 n_231 gnd! 868.4fF
C806 PD_0xx0xx0x gnd! 1163.1fF
C807 PD_n_0xx0xx0x gnd! 701.0fF
C808 n_1515 gnd! 345.2fF
C809 nTWOCYCLE_phi1 gnd! 376.4fF
C810 n_1379 gnd! 965.6fF
C811 n_1161 gnd! 338.2fF
C812 n_253 gnd! 1337.6fF
C813 n_19 gnd! 431.8fF
C814 n_442 gnd! 875.4fF
C815 n_1619 gnd! 774.8fF
C816 pipeUNK21 gnd! 329.6fF
C817 n_1231 gnd! 506.6fF
C818 n_781 gnd! 2688.7fF
C819 n_1154 gnd! 679.4fF
C820 n_1409 gnd! 271.0fF
C821 n_1448 gnd! 429.4fF
C822 n_1330 gnd! 297.6fF
C823 n_2 gnd! 374.0fF
C824 n_1039 gnd! 628.6fF
C825 n_1124 gnd! 489.4fF
C826 pipeUNK39 gnd! 245.6fF
C827 PD_xxxx10x0 gnd! 1575.1fF
C828 pd2_clearIR gnd! 959.8fF
C829 pd3_clearIR gnd! 1222.4fF
C830 pd5_clearIR gnd! 1220.1fF
C831 PD_1xx000x0 gnd! 1566.1fF
C832 n_732 gnd! 1189.6fF
C833 n_137 gnd! 97.6fF
C834 n_1718 gnd! 582.8fF
C835 n_770 gnd! 606.2fF
C836 n_812 gnd! 518.2fF
C837 pd4_clearIR gnd! 1272.2fF
C838 pd7_clearIR gnd! 984.0fF
C839 pd1_clearIR gnd! 964.8fF
C840 pd0_clearIR gnd! 934.2fF
C841 PD_xxx010x1 gnd! 1211.5fF
C842 n_17 gnd! 774.4fF
C843 n_504 gnd! 666.6fF
C844 pipeUNK42 gnd! 421.0fF
C845 nTWOCYCLE gnd! 1162.8fF
C846 pipeUNK40 gnd! 246.8fF
C847 n_1380 gnd! 787.8fF
C848 n_14 gnd! 1426.9fF
C849 n_666 gnd! 297.0fF
C850 ONEBYTE gnd! 2057.0fF
C851 pipenWR_phi2 gnd! 271.8fF
C852 pipeUNK41 gnd! 222.8fF
C853 n_1497 gnd! 571.2fF
C854 n_964 gnd! 743.4fF
C855 n_653 gnd! 230.4fF
C856 pipenT0 gnd! 489.6fF
C857 n_1180 gnd! 594.6fF
C858 n_1533 gnd! 524.4fF
C859 n_664 gnd! 428.2fF
C860 n_889 gnd! 531.4fF
C861 n_390 gnd! 572.0fF
C862 n_1120 gnd! 468.6fF
C863 n_424 gnd! 576.6fF
C864 n_109 gnd! 1644.7fF
C865 n_816 gnd! 204.4fF
C866 n_774 gnd! 1528.9fF
C867 n_327 gnd! 1032.2fF
C868 n_591 gnd! 242.0fF
C869 nop_set_C gnd! 2191.1fF
C870 n_191 gnd! 642.0fF
C871 nWR gnd! 1532.5fF
C872 n_387 gnd! 311.6fF
C873 n_586 gnd! 1590.1fF
C874 n_1517 gnd! 828.6fF
C875 n_853 gnd! 595.0fF
C876 n_206 gnd! 2633.4fF
C877 n_559 gnd! 231.4fF
C878 n_608 gnd! 412.6fF
C879 n_1278 gnd! 224.4fF
C880 n_1642 gnd! 2087.5fF
C881 n_176 gnd! 1006.4fF
C882 n_1655 gnd! 343.0fF
C883 n_1697 gnd! 2248.4fF
C884 n_275 gnd! 542.0fF
C885 n_1272 gnd! 298.2fF
C886 n_773 gnd! 591.2fF
C887 n_759 gnd! 219.4fF
C888 n_198 gnd! 874.4fF
C889 pipeUNK37 gnd! 303.2fF
C890 n_944 gnd! 713.6fF
C891 n_218 gnd! 533.6fF
C892 n_470 gnd! 631.2fF
C893 n_1276 gnd! 291.0fF
C894 n_AxBxC_0 gnd! 478.4fF
C895 n_406 gnd! 86.0fF
C896 n_942 gnd! 224.0fF
C897 C01 gnd! 709.8fF
C898 nA_B2 gnd! 1312.8fF
C899 n_452 gnd! 148.4fF
C900 alua2 gnd! 484.2fF
C901 n_458 gnd! 518.2fF
C902 idb2 gnd! 4120.2fF
C903 alub2 gnd! 679.4fF
C904 s6 gnd! 269.9fF
C905 nots6 gnd! 219.8fF
C906 x7 gnd! 203.0fF
C907 notx7 gnd! 450.2fF
C908 n_871 gnd! 720.0fF
C909 n_1187 gnd! 487.2fF
C910 n_618 gnd! 1067.0fF
C911 s5 gnd! 279.6fF
C912 nots5 gnd! 213.2fF
C913 x6 gnd! 205.0fF
C914 notx6 gnd! 462.2fF
C915 sb7 gnd! 3483.2fF
C916 y7 gnd! 210.4fF
C917 noty7 gnd! 447.4fF
C918 n_1251 gnd! 760.4fF
C919 abh0 gnd! 777.2fF
C920 nABH0 gnd! 378.2fF
C921 n_1668 gnd! 588.6fF
C922 adh0 gnd! 5243.6fF
C923 n_577 gnd! 41.2fF
C924 nABL7 gnd! 296.6fF
C925 n_1046 gnd! 528.0fF
C926 adl7 gnd! 3591.6fF
C927 sb6 gnd! 3523.2fF
C928 y6 gnd! 201.6fF
C929 noty6 gnd! 451.4fF
C930 n_1724 gnd! 765.2fF
C931 n_496 gnd! 507.8fF
C932 n_280 gnd! 1091.2fF
C933 s4 gnd! 275.8fF
C934 nots4 gnd! 214.4fF
C935 x5 gnd! 216.6fF
C936 notx5 gnd! 447.6fF
C937 n_578 gnd! 771.2fF
C938 n_973 gnd! 513.2fF
C939 n_3 gnd! 1090.6fF
C940 s3 gnd! 276.3fF
C941 nots3 gnd! 219.2fF
C942 x4 gnd! 202.4fF
C943 notx4 gnd! 450.4fF
C944 n_436 gnd! 721.6fF
C945 n_34 gnd! 520.4fF
C946 n_998 gnd! 1104.7fF
C947 n_A_B_1 gnd! 974.0fF
C948 naluresult1 gnd! 1563.3fF
C949 n_1348 gnd! 92.0fF
C950 n_AxB_0 gnd! 714.3fF
C951 dpc21_ADDADL gnd! 2090.8fF
C952 dpc20_ADDSB06 gnd! 1842.2fF
C953 n_1033 gnd! 434.8fF
C954 n_75 gnd! 444.6fF
C955 dpc19_ADDSB7 gnd! 1781.6fF
C956 A_B0 gnd! 341.0fF
C957 n_105 gnd! 411.0fF
C958 nA_B1 gnd! 837.0fF
C959 n_189 gnd! 173.2fF
C960 alua1 gnd! 460.6fF
C961 n_583 gnd! 527.0fF
C962 idb1 gnd! 4026.4fF
C963 alub1 gnd! 667.2fF
C964 n_A_B_0 gnd! 1378.2fF
C965 naluresult0 gnd! 1452.8fF
C966 nA_B0 gnd! 1574.8fF
C967 n_316 gnd! 148.4fF
C968 alua0 gnd! 458.0fF
C969 n_624 gnd! 495.4fF
C970 idb0 gnd! 3953.4fF
C971 dpc18_nDAA gnd! 2219.6fF
C972 n_241 gnd! 625.0fF
C973 n_714 gnd! 374.8fF
C974 n_709 gnd! 437.8fF
C975 n_154 gnd! 581.6fF
C976 n_906 gnd! 782.0fF
C977 n_1499 gnd! 652.6fF
C978 dpc17_SUMS gnd! 1964.2fF
C979 n_1305 gnd! 459.2fF
C980 n_1552 gnd! 448.6fF
C981 n_772 gnd! 577.0fF
C982 n_1593 gnd! 643.0fF
C983 n_745 gnd! 225.6fF
C984 n_512 gnd! 248.0fF
C985 n_1333 gnd! 216.2fF
C986 n_1450 gnd! 285.4fF
C987 n_1674 gnd! 274.2fF
C988 n_226 gnd! 277.8fF
C989 n_1705 gnd! 1819.0fF
C990 n_930 gnd! 859.4fF
C991 n_1427 gnd! 1024.6fF
C992 n_1151 gnd! 195.6fF
C993 n_467 gnd! 848.9fF
C994 n_1286 gnd! 1004.6fF
C995 aluvout gnd! 2899.8fF
C996 n_1245 gnd! 2869.0fF
C997 n_80 gnd! 479.4fF
C998 dpc22_nDSA gnd! 1810.8fF
C999 n_674 gnd! 611.2fF
C1000 dpc14_SRS gnd! 2037.1fF
C1001 dpc13_ORS gnd! 2108.0fF
C1002 dpc16_EORS gnd! 1919.8fF
C1003 alub0 gnd! 689.3fF
C1004 s2 gnd! 290.0fF
C1005 nots2 gnd! 226.8fF
C1006 x3 gnd! 215.4fF
C1007 notx3 gnd! 456.4fF
C1008 n_242 gnd! 775.2fF
C1009 n_1190 gnd! 504.8fF
C1010 n_1389 gnd! 1085.0fF
C1011 s1 gnd! 294.0fF
C1012 nots1 gnd! 215.2fF
C1013 x2 gnd! 222.4fF
C1014 notx2 gnd! 448.0fF
C1015 n_1694 gnd! 739.8fF
C1016 n_518 gnd! 732.4fF
C1017 abl7 gnd! 1003.0fF
C1018 n_1026 gnd! 551.4fF
C1019 n_322 gnd! 2648.6fF
C1020 ab6 gnd! 10469.3fF
C1021 n_171 gnd! 2545.4fF
C1022 n_524 gnd! 41.2fF
C1023 nABL6 gnd! 302.2fF
C1024 n_1548 gnd! 500.8fF
C1025 adl6 gnd! 3731.4fF
C1026 sb5 gnd! 3457.6fF
C1027 y5 gnd! 210.2fF
C1028 noty5 gnd! 428.0fF
C1029 n_733 gnd! 732.0fF
C1030 abl6 gnd! 1001.4fF
C1031 n_1195 gnd! 551.4fF
C1032 n_1191 gnd! 2312.6fF
C1033 n_1254 gnd! 2877.0fF
C1034 n_463 gnd! 38.0fF
C1035 nABL5 gnd! 290.6fF
C1036 n_1094 gnd! 503.6fF
C1037 adl5 gnd! 3701.7fF
C1038 sb4 gnd! 3511.6fF
C1039 y4 gnd! 211.2fF
C1040 noty4 gnd! 449.6fF
C1041 ab5 gnd! 10332.1fF
C1042 abl5 gnd! 1002.8fF
C1043 n_172 gnd! 546.8fF
C1044 n_1633 gnd! 2357.6fF
C1045 n_210 gnd! 2796.6fF
C1046 ab4 gnd! 10233.7fF
C1047 n_738 gnd! 41.2fF
C1048 nABL4 gnd! 291.4fF
C1049 n_1519 gnd! 473.8fF
C1050 adl4 gnd! 3784.1fF
C1051 n_658 gnd! 711.2fF
C1052 abl4 gnd! 960.6fF
C1053 n_1676 gnd! 589.8fF
C1054 n_634 gnd! 2328.4fF
C1055 n_86 gnd! 2722.4fF
C1056 sb3 gnd! 3487.7fF
C1057 y3 gnd! 207.8fF
C1058 noty3 gnd! 441.0fF
C1059 n_1531 gnd! 739.6fF
C1060 n_864 gnd! 41.2fF
C1061 nABL3 gnd! 301.6fF
C1062 n_1507 gnd! 558.6fF
C1063 adl3 gnd! 3738.0fF
C1064 sb2 gnd! 3511.7fF
C1065 y2 gnd! 224.4fF
C1066 noty2 gnd! 447.4fF
C1067 n_1711 gnd! 506.8fF
C1068 n_694 gnd! 1080.2fF
C1069 s0 gnd! 290.2fF
C1070 nots0 gnd! 247.0fF
C1071 x1 gnd! 213.8fF
C1072 notx1 gnd! 449.6fF
C1073 n_1709 gnd! 725.6fF
C1074 n_983 gnd! 495.8fF
C1075 n_332 gnd! 1105.0fF
C1076 x0 gnd! 211.0fF
C1077 notx0 gnd! 429.6fF
C1078 n_1169 gnd! 744.4fF
C1079 n_1491 gnd! 765.4fF
C1080 ab3 gnd! 10296.1fF
C1081 abl3 gnd! 962.4fF
C1082 n_990 gnd! 572.8fF
C1083 n_1041 gnd! 2356.4fF
C1084 n_138 gnd! 2698.2fF
C1085 n_1636 gnd! 46.4fF
C1086 nABL2 gnd! 298.0fF
C1087 n_935 gnd! 465.6fF
C1088 adl2 gnd! 3845.4fF
C1089 sb1 gnd! 3480.7fF
C1090 y1 gnd! 213.2fF
C1091 noty1 gnd! 465.2fF
C1092 n_767 gnd! 763.8fF
C1093 sb0 gnd! 3696.3fF
C1094 y0 gnd! 198.4fF
C1095 noty0 gnd! 437.2fF
C1096 abl2 gnd! 989.2fF
C1097 n_951 gnd! 577.6fF
C1098 ab2 gnd! 10429.3fF
C1099 n_1152 gnd! 2198.2fF
C1100 n_642 gnd! 2500.0fF
C1101 n_416 gnd! 42.8fF
C1102 nABL1 gnd! 285.8fF
C1103 n_1016 gnd! 492.6fF
C1104 adl1 gnd! 3855.3fF
C1105 n_564 gnd! 753.6fF
C1106 abl1 gnd! 1004.6fF
C1107 n_842 gnd! 561.4fF
C1108 ab1 gnd! 10245.0fF
C1109 n_1479 gnd! 2167.4fF
C1110 n_66 gnd! 2454.8fF
C1111 n_246 gnd! 46.4fF
C1112 nABL0 gnd! 302.0fF
C1113 n_123 gnd! 510.4fF
C1114 adl0 gnd! 4018.2fF
C1115 n_1255 gnd! 450.8fF
C1116 n_108 gnd! 411.6fF
C1117 n_531 gnd! 645.2fF
C1118 dpc15_ANDS gnd! 2057.7fF
C1119 dpc10_ADLADD gnd! 3055.4fF
C1120 n_1256 gnd! 512.8fF
C1121 dpc11_SBADD gnd! 2742.9fF
C1122 n_491 gnd! 412.6fF
C1123 dpc12_0ADD gnd! 2388.4fF
C1124 n_1364 gnd! 621.2fF
C1125 n_708 gnd! 426.4fF
C1126 dpc9_DBADD gnd! 2576.8fF
C1127 n_956 gnd! 434.0fF
C1128 dpc8_nDBADD gnd! 2434.2fF
C1129 n_225 gnd! 443.2fF
C1130 dpc7_SS gnd! 2743.4fF
C1131 n_763 gnd! 418.0fF
C1132 dpc6_SBS gnd! 2403.2fF
C1133 dpc5_SADL gnd! 2036.6fF
C1134 n_95 gnd! 283.0fF
C1135 n_91 gnd! 654.4fF
C1136 n_1541 gnd! 650.0fF
C1137 n_1230 gnd! 650.2fF
C1138 n_71 gnd! 423.8fF
C1139 dpc4_SSB gnd! 2456.6fF
C1140 n_282 gnd! 411.6fF
C1141 dpc3_SBX gnd! 2501.0fF
C1142 n_196 gnd! 408.2fF
C1143 dpc1_SBY gnd! 2319.4fF
C1144 n_593 gnd! 397.8fF
C1145 n_476 gnd! 659.6fF
C1146 n_1223 gnd! 659.4fF
C1147 n_1534 gnd! 669.2fF
C1148 n_35 gnd! 649.6fF
C1149 n_6 gnd! 658.4fF
C1150 n_662 gnd! 411.2fF
C1151 n_543 gnd! 654.0fF
C1152 n_101 gnd! 275.4fF
C1153 n_1529 gnd! 271.0fF
C1154 n_1477 gnd! 175.4fF
C1155 n_360 gnd! 167.6fF
C1156 n_1027 gnd! 164.6fF
C1157 n_688 gnd! 151.2fF
C1158 n_805 gnd! 163.8fF
C1159 n_441 gnd! 415.8fF
C1160 n_355 gnd! 639.6fF
C1161 n_625 gnd! 658.8fF
C1162 n_692 gnd! 631.6fF
C1163 n_931 gnd! 612.0fF
C1164 n_1526 gnd! 596.4fF
C1165 n_968 gnd! 199.2fF
C1166 n_1093 gnd! 617.0fF
C1167 n_1375 gnd! 535.2fF
C1168 notalucin gnd! 1412.7fF
C1169 n_415 gnd! 250.0fF
C1170 n_599 gnd! 330.2fF
C1171 dpc28_0ADH0 gnd! 1751.4fF
C1172 n_182 gnd! 2285.3fF
C1173 n_462 gnd! 1386.4fF
C1174 n_1338 gnd! 235.6fF
C1175 n_180 gnd! 631.6fF
C1176 n_1716 gnd! 1706.1fF
C1177 n_1211 gnd! 2506.6fF
C1178 n_916 gnd! 1227.4fF
C1179 n_1708 gnd! 1262.2fF
C1180 op_rmw gnd! 330.2fF
C1181 n_1137 gnd! 891.6fF
C1182 pipeUNK36 gnd! 500.4fF
C1183 short_circuit_idx_add gnd! 965.4fF
C1184 n_347 gnd! 2327.2fF
C1185 n_1065 gnd! 691.5fF
C1186 n_790 gnd! 1219.8fF
C1187 n_368 gnd! 1181.0fF
C1188 n_1391 gnd! 2352.8fF
C1189 nop_store gnd! 727.2fF
C1190 n_510 gnd! 908.2fF
C1191 n_10 gnd! 1505.6fF
C1192 n_1407 gnd! 216.8fF
C1193 n_933 gnd! 690.6fF
C1194 pipedpc28 gnd! 263.0fF
C1195 n_1141 gnd! 586.0fF
C1196 n_1089 gnd! 554.4fF
C1197 n_88 gnd! 193.8fF
C1198 n_982 gnd! 194.0fF
C1199 n_680 gnd! 358.6fF
C1200 n_572 gnd! 1434.5fF
C1201 n_261 gnd! 605.0fF
C1202 pipeUNK35 gnd! 187.4fF
C1203 n_720 gnd! 1138.2fF
C1204 pipeUNK34 gnd! 209.4fF
C1205 n_238 gnd! 822.6fF
C1206 n_501 gnd! 1248.2fF
C1207 n_636 gnd! 500.0fF
C1208 n_726 gnd! 1046.0fF
C1209 n_1280 gnd! 183.2fF
C1210 n_1262 gnd! 1063.2fF
C1211 n_1679 gnd! 225.4fF
C1212 n_1574 gnd! 230.8fF
C1213 n_796 gnd! 158.8fF
C1214 op_SUMS gnd! 983.6fF
C1215 alucin gnd! 585.4fF
C1216 n_590 gnd! 212.0fF
C1217 n_1215 gnd! 3390.6fF
C1218 n_223 gnd! 346.0fF
C1219 n_533 gnd! 724.8fF
C1220 pipeUNK22 gnd! 201.8fF
C1221 pipeUNK23 gnd! 228.2fF
C1222 n_819 gnd! 2639.2fF
C1223 pipephi2Reset0 gnd! 207.0fF
C1224 n_29 gnd! 640.4fF
C1225 n_51 gnd! 150.8fF
C1226 n_1688 gnd! 1089.0fF
C1227 n_334 gnd! 3253.2fF
C1228 n_1508 gnd! 374.0fF
C1229 n_46 gnd! 682.6fF
C1230 n_272 gnd! 3004.2fF
C1231 n_239 gnd! 119.6fF
C1232 n_992 gnd! 432.8fF
C1233 n_813 gnd! 659.2fF
C1234 n_25 gnd! 1253.0fF
C1235 n_1053 gnd! 223.6fF
C1236 n_1440 gnd! 356.6fF
C1237 Pout3 gnd! 3269.2fF
C1238 n_506 gnd! 1795.4fF
C1239 n_550 gnd! 683.0fF
C1240 n_885 gnd! 2469.4fF
C1241 n_1219 gnd! 364.8fF
C1242 n_1004 gnd! 186.4fF
C1243 n_979 gnd! 375.2fF
C1244 n_1347 gnd! 2822.5fF
C1245 n_134 gnd! 1851.0fF
C1246 n_1037 gnd! 2447.8fF
C1247 n_824 gnd! 2427.0fF
C1248 n_1012 gnd! 172.2fF
C1249 n_366 gnd! 583.4fF
C1250 nop_branch_done gnd! 422.0fF
C1251 n_595 gnd! 636.0fF
C1252 n_669 gnd! 441.0fF
C1253 n_1225 gnd! 4309.4fF
C1254 n_1412 gnd! 404.2fF
C1255 n_1222 gnd! 535.0fF
C1256 n_384 gnd! 1391.6fF
C1257 n_1681 gnd! 132.0fF
C1258 n_905 gnd! 406.6fF
C1259 n_1090 gnd! 2086.9fF
C1260 n_1563 gnd! 123.6fF
C1261 n_397 gnd! 468.2fF
C1262 n_11 gnd! 2472.5fF
C1263 n_1455 gnd! 2876.9fF
C1264 n_928 gnd! 1003.4fF
C1265 n_1378 gnd! 57.2fF
C1266 n_605 gnd! 811.6fF
C1267 n_673 gnd! 494.8fF
C1268 n_1304 gnd! 768.4fF
C1269 n_521 gnd! 167.4fF
C1270 n_339 gnd! 198.4fF
C1271 n_621 gnd! 200.4fF
C1272 n_459 gnd! 174.2fF
C1273 n_460 gnd! 174.8fF
C1274 n_795 gnd! 422.8fF
C1275 n_656 gnd! 131.6fF
C1276 n_396 gnd! 385.4fF
C1277 n_1594 gnd! 582.4fF
C1278 D1x1 gnd! 4848.8fF
C1279 n_760 gnd! 267.6fF
C1280 n_236 gnd! 3463.8fF
C1281 n_405 gnd! 245.0fF
C1282 n_1343 gnd! 527.4fF
C1283 n_877 gnd! 1512.7fF
C1284 n_779 gnd! 1670.0fF
C1285 n_1172 gnd! 549.2fF
C1286 BRtaken gnd! 4036.6fF
C1287 n_1085 gnd! 1154.7fF
C1288 n_1365 gnd! 114.4fF
C1289 n_104 gnd! 4161.6fF
C1290 n_1408 gnd! 585.8fF
C1291 n_1044 gnd! 2513.2fF
C1292 INTG gnd! 1121.0fF
C1293 n_372 gnd! 371.2fF
C1294 op_EORS gnd! 954.0fF
C1295 n_630 gnd! 2774.8fF
C1296 n_256 gnd! 3483.3fF
C1297 n_847 gnd! 503.2fF
C1298 n_1258 gnd! 2903.2fF
C1299 n_1130 gnd! 2216.4fF
C1300 n_192 gnd! 1893.6fF
C1301 n_1081 gnd! 1233.9fF
C1302 pipeUNK32 gnd! 285.5fF
C1303 pipeUNK33 gnd! 234.8fF
C1304 n_152 gnd! 906.2fF
C1305 abl0 gnd! 968.4fF
C1306 n_1660 gnd! 585.6fF
C1307 n_855 gnd! 2162.2fF
C1308 ab0 gnd! 9352.2fF
C1309 dpc2_XSB gnd! 2468.5fF
C1310 dpc0_YSB gnd! 2544.7fF
C1311 n_1100 gnd! 2444.8fF
C1312 n_1701 gnd! 1105.5fF
C1313 diff_237_1656# gnd! 337.2fF
C1314 testpad_6 gnd! 796.3fF
C1315 ADL_ABL gnd! 1777.0fF
C1316 ADH_ABH gnd! 5620.7fF
C1317 n_602 gnd! 409.8fF
C1318 n_969 gnd! 414.2fF
C1319 n_130 gnd! 419.8fF
C1320 n_1067 gnd! 463.4fF
C1321 n_38 gnd! 494.0fF
C1322 testpad_4 gnd! 551.3fF
C1323 testpad_2 gnd! 3869.8fF
C1324 n_1127 gnd! 924.8fF
C1325 testpad_5 gnd! 2739.1fF
C1326 testpad_1 gnd! 1656.8fF
C1327 n_1247 gnd! 6019.8fF
C1328 n_133 gnd! 636.6fF
C1329 n_1404 gnd! 170.0fF
C1330 n_161 gnd! 617.6fF
C1331 n_220 gnd! 644.8fF
C1332 n_839 gnd! 489.2fF
C1333 n_43 gnd! 4654.0fF
C1334 n_582 gnd! 671.0fF
C1335 n_1113 gnd! 192.0fF
C1336 n_190 gnd! 214.4fF
C1337 n_610 gnd! 231.8fF
C1338 n_0_ADL2 gnd! 1257.2fF
C1339 n_0_ADL1 gnd! 1214.2fF
C1340 pipeVectorA1 gnd! 246.2fF
C1341 n_1117 gnd! 475.2fF
C1342 n_815 gnd! 569.2fF
C1343 n_952 gnd! 2585.6fF
C1344 n_50 gnd! 182.0fF
C1345 pipeUNK31 gnd! 233.0fF
C1346 n_1178 gnd! 1569.8fF
C1347 pipeUNK30 gnd! 252.8fF
C1348 n_473 gnd! 1167.0fF
C1349 n_1002 gnd! 2128.3fF
C1350 n_629 gnd! 1226.8fF
C1351 n_646 gnd! 5419.1fF
C1352 n_202 gnd! 422.4fF
C1353 op_ORS gnd! 1288.1fF
C1354 n_385 gnd! 489.2fF
C1355 n_782 gnd! 1300.6fF
C1356 n_1040 gnd! 498.4fF
C1357 n_1377 gnd! 446.8fF
C1358 nnT2BR gnd! 5072.3fF
C1359 n_1092 gnd! 848.1fF
C1360 n_118 gnd! 1142.0fF
C1361 n_480 gnd! 819.8fF
C1362 op_ANDS gnd! 2789.4fF
C1363 n_837 gnd! 1100.6fF
C1364 n_1145 gnd! 650.6fF
C1365 n_980 gnd! 771.2fF
C1366 n_389 gnd! 956.3fF
C1367 n_1055 gnd! 2751.9fF
C1368 n_1560 gnd! 626.8fF
C1369 n_1000 gnd! 526.8fF
C1370 n_300 gnd! 1709.0fF
C1371 n_1555 gnd! 129.2fF
C1372 n_1118 gnd! 156.4fF
C1373 n_1649 gnd! 3040.6fF
C1374 n_1107 gnd! 960.2fF
C1375 n_440 gnd! 3709.7fF
C1376 n_638 gnd! 431.4fF
C1377 n_604 gnd! 3022.8fF
C1378 pipeVectorA2 gnd! 206.0fF
C1379 n_70 gnd! 617.6fF
C1380 n_1054 gnd! 468.6fF
C1381 pipeVectorA0 gnd! 350.6fF
C1382 n_911 gnd! 1706.7fF
C1383 n_0_ADL0 gnd! 1666.9fF
C1384 n_696 gnd! 1177.4fF
C1385 n_1361 gnd! 272.8fF ;**FLOATING
C1386 n_79 gnd! 1494.4fF
C1387 diff_713_2318# gnd! 73.4fF ;**FLOATING
C1388 diff_726_2349# gnd! 43.2fF ;**FLOATING
C1389 diff_713_2349# gnd! 43.2fF ;**FLOATING
C1390 n_1132 gnd! 213.8fF
C1391 pipephi2Reset0x gnd! 175.8fF
C1392 n_1087 gnd! 665.8fF
C1393 n_717 gnd! 717.0fF
C1394 n_1712 gnd! 1224.9fF
C1395 n_1317 gnd! 335.2fF ;**FLOATING
C1396 n_1261 gnd! 127.2fF ;**FLOATING
C1397 n_1207 gnd! 127.2fF ;**FLOATING
C1398 n_728 gnd! 917.2fF
C1399 n_411 gnd! 39.6fF ;**FLOATING
C1400 n_1663 gnd! 394.8fF ;**FLOATING
C1401 diff_822_2540# gnd! 160.6fF ;**FLOATING
C1402 n_497 gnd! 358.8fF ;**FLOATING
C1403 n_563 gnd! 384.8fF ;**FLOATING
C1404 op_SRS gnd! 4814.2fF
C1405 n_902 gnd! 341.0fF
C1406 n_920 gnd! 397.0fF
C1407 pipeUNK27 gnd! 167.8fF
C1408 n_1598 gnd! 234.4fF
C1409 n_1511 gnd! 418.6fF
C1410 n_785 gnd! 167.8fF
C1411 pipeUNK28 gnd! 197.6fF
C1412 n_1189 gnd! 357.2fF
C1413 n_1624 gnd! 277.0fF
C1414 n_139 gnd! 821.8fF
C1415 n_267 gnd! 2761.2fF
C1416 n_383 gnd! 1113.0fF
C1417 n_917 gnd! 529.4fF
C1418 n_1058 gnd! 145.2fF
C1419 n_262 gnd! 799.8fF
C1420 pipeUNK29 gnd! 486.0fF
C1421 n_169 gnd! 513.4fF
C1422 n_1175 gnd! 605.6fF
C1423 n_1447 gnd! 268.0fF
C1424 sync gnd! 10766.4fF
C1425 n_417 gnd! 2295.2fF
C1426 n_1101 gnd! 3418.2fF
C1427 n_132 gnd! 4034.6fF
C1428 pipeUNK26 gnd! 176.6fF
C1429 n_317 gnd! 533.2fF
C1430 n_1714 gnd! 893.8fF
C1431 C1x5Reset gnd! 4819.8fF
C1432 n_1289 gnd! 723.6fF
C1433 n_1358 gnd! 1956.4fF
C1434 n_632 gnd! 1711.8fF
C1435 n_1109 gnd! 2010.8fF
C1436 n_544 gnd! 1081.4fF
C1437 n_454 gnd! 182.4fF
C1438 n_689 gnd! 956.2fF
C1439 n_1586 gnd! 1807.6fF
C1440 n_946 gnd! 1941.2fF
C1441 n_734 gnd! 287.6fF
C1442 n_1103 gnd! 117.6fF
C1443 n_445 gnd! 2263.8fF
C1444 n_1464 gnd! 1137.6fF
C1445 n_616 gnd! 2466.3fF
C1446 n_844 gnd! 2181.6fF
C1447 n_1351 gnd! 226.8fF
C1448 n_1244 gnd! 435.2fF
C1449 n_1106 gnd! 2931.1fF
C1450 n_1604 gnd! 143.6fF
C1451 n_1397 gnd! 143.6fF
C1452 n_698 gnd! 276.0fF
C1453 VEC0 gnd! 2595.0fF
C1454 n_508 gnd! 275.2fF
C1455 n_335 gnd! 4511.8fF
C1456 n_1303 gnd! 2171.0fF
C1457 n_1717 gnd! 2883.4fF
C1458 n_1126 gnd! 195.0fF
C1459 n_1290 gnd! 832.0fF
C1460 n_912 gnd! 201.2fF
C1461 VEC1 gnd! 1056.8fF
C1462 n_1452 gnd! 262.6fF
C1463 n_861 gnd! 909.6fF
C1464 brk_done gnd! 6060.2fF
C1465 n_1291 gnd! 238.6fF
C1466 clock2 gnd! 5079.3fF
C1467 n_1312 gnd! 610.6fF
C1468 n_1609 gnd! 399.2fF
C1469 pd6_clearIR gnd! 1142.8fF
C1470 n_1309 gnd! 759.0fF
C1471 n_74 gnd! 57.2fF
C1472 clock1 gnd! 4729.0fF
C1473 notir5 gnd! 5653.2fF
C1474 n_1693 gnd! 258.0fF
C1475 nNMIG gnd! 3105.0fF
C1476 n_799 gnd! 263.2fF
C1477 n_1675 gnd! 411.8fF
C1478 n_1149 gnd! 273.2fF
C1479 n_1339 gnd! 431.2fF
C1480 nVEC gnd! 2809.8fF
C1481 ir5 gnd! 4602.6fF
C1482 notir6 gnd! 4627.6fF
C1483 n_571 gnd! 1044.2fF
C1484 n_343 gnd! 57.2fF
C1485 n_1300 gnd! 416.8fF
C1486 ir6 gnd! 4539.6fF
C1487 notir2 gnd! 4693.4fF
C1488 diff_3658_3262# gnd! 235.6fF ;**FLOATING
C1489 n_1083 gnd! 1158.3fF
C1490 n_1590 gnd! 59.6fF
C1491 n_597 gnd! 203.8fF
C1492 ir2 gnd! 4569.6fF
C1493 diff_3658_3288# gnd! 213.2fF ;**FLOATING
C1494 n_1620 gnd! 429.6fF
C1495 notir3 gnd! 4570.6fF
C1496 diff_3658_3314# gnd! 202.2fF ;**FLOATING
C1497 ir3 gnd! 4582.2fF
C1498 n_1252 gnd! 289.8fF
C1499 pipenVEC gnd! 263.4fF
C1500 n_1578 gnd! 404.0fF
C1501 n_882 gnd! 671.8fF
C1502 n_562 gnd! 369.4fF
C1503 NMIL gnd! 866.4fF
C1504 n_227 gnd! 1223.2fF
C1505 n_703 gnd! 59.6fF
C1506 notir4 gnd! 4694.8fF
C1507 n_927 gnd! 413.4fF
C1508 n_1368 gnd! 1468.6fF
C1509 n_862 gnd! 7487.1fF
C1510 pipeT_SYNC gnd! 326.6fF
C1511 ir4 gnd! 4567.6fF
C1512 diff_3659_3362# gnd! 642.6fF ;**FLOATING
C1513 diff_3704_3419# gnd! 209.8fF ;**FLOATING
C1514 diff_3681_3419# gnd! 220.8fF ;**FLOATING
C1515 n_1183 gnd! 54.8fF
C1516 n_1605 gnd! 1532.9fF
C1517 n_541 gnd! 390.4fF
C1518 diff_3658_3431# gnd! 205.2fF ;**FLOATING
C1519 n_363 gnd! 446.8fF
C1520 notir7 gnd! 4676.4fF
C1521 n_1091 gnd! 566.2fF
C1522 n_1360 gnd! 220.2fF
C1523 ir7 gnd! 4568.6fF
C1524 notir0 gnd! 4460.4fF
C1525 n_409 gnd! 1598.5fF
C1526 n_724 gnd! 57.2fF
C1527 n_310 gnd! 392.4fF
C1528 n_1641 gnd! 1474.4fF
C1529 n_237 gnd! 54.8fF
C1530 fetch gnd! 3027.4fF
C1531 irline3 gnd! 4175.4fF
C1532 n_12 gnd! 278.8fF
C1533 n_1575 gnd! 746.6fF
C1534 n_644 gnd! 234.4fF
C1535 _t2 gnd! 4149.6fF
C1536 pipeT2out gnd! 528.8fF
C1537 n_1558 gnd! 452.0fF
C1538 n_428 gnd! 639.0fF
C1539 n_119 gnd! 424.6fF
C1540 n_1133 gnd! 780.4fF
C1541 ir1 gnd! 705.8fF
C1542 _t3 gnd! 4217.2fF
C1543 n_678 gnd! 1002.2fF
C1544 notir1 gnd! 4482.8fF
C1545 notRnWprepad gnd! 4978.8fF
C1546 ir0 gnd! 1275.4fF
C1547 op_clv gnd! 2556.7fF
C1548 op_T4_mem_abs_idx gnd! 1323.6fF
C1549 op_implied gnd! 1463.4fF
C1550 nop_branch_bit7 gnd! 3285.9fF
C1551 op_T2_mem_zp gnd! 1410.8fF
C1552 nop_branch_bit6 gnd! 3180.8fF
C1553 x_op_push_pull gnd! 1549.6fF
C1554 op_T__asl_rol_a gnd! 1615.3fF
C1555 op_T5_mem_ind_idx gnd! 1422.8fF
C1556 op_T3_mem_abs gnd! 1417.5fF
C1557 op_T0_cld_sed gnd! 1581.1fF
C1558 op_T__cpx_cpy_imm_zp gnd! 1526.3fF
C1559 op_T__cmp gnd! 1414.8fF
C1560 op_T__cpx_cpy_abs gnd! 1593.3fF
C1561 op_T0_plp gnd! 1636.5fF
C1562 x_op_T4_rti gnd! 1680.3fF
C1563 x_op_T__adc_sbc gnd! 3214.0fF
C1564 op_T0_clc_sec gnd! 1826.1fF
C1565 n_1363 gnd! 866.0fF
C1566 op_asl_rol gnd! 1400.3fF
C1567 x_op_T3_plp_pla gnd! 1630.0fF
C1568 x_op_T0_bit gnd! 1980.7fF
C1569 op_T3_mem_zp_idx gnd! 1282.0fF
C1570 op_T__bit gnd! 2618.2fF
C1571 op_T0_cli_sei gnd! 1554.6fF
C1572 op_lsr_ror_dec_inc gnd! 1127.1fF
C1573 op_T5_rti_rts gnd! 1716.5fF
C1574 op_T4_jmp gnd! 2180.4fF
C1575 op_T2_php gnd! 1839.3fF
C1576 op_store gnd! 1293.4fF
C1577 op_T2_jmp_abs gnd! 1745.7fF
C1578 xx_op_T5_jsr gnd! 1794.9fF
C1579 n_173 gnd! 838.1fF
C1580 op_T2_php_pha gnd! 1757.4fF
C1581 op_T4_brk gnd! 2008.7fF
C1582 op_push_pull gnd! 1778.3fF
C1583 op_jsr gnd! 1760.0fF
C1584 op_T3_branch gnd! 1650.2fF
C1585 x_op_T4_ind_y gnd! 1463.6fF
C1586 op_T3_abs_idx_ind gnd! 1260.8fF
C1587 n_9 gnd! 116.4fF
C1588 diff_2598_3600# gnd! 73.8fF
C1589 x_op_jmp gnd! 1698.2fF
C1590 op_brk_rti gnd! 1582.2fF
C1591 op_T0_jmp gnd! 1818.8fF
C1592 x_op_T3_abs_idx gnd! 1304.8fF
C1593 op_T3 gnd! 1122.0fF
C1594 op_T5_ind_x gnd! 1543.6fF
C1595 op_T0_brk_rti gnd! 1712.3fF
C1596 op_T5_rts gnd! 3343.6fF
C1597 op_T4 gnd! 1063.2fF
C1598 op_T2_ind gnd! 1403.1fF
C1599 op_T2_branch gnd! 1559.6fF
C1600 op_T2_abs_access gnd! 2382.0fF
C1601 n_402 gnd! 250.8fF
C1602 n_400 gnd! 553.6fF
C1603 n_1059 gnd! 496.4fF
C1604 n_834 gnd! 856.3fF
C1605 rw gnd! 10912.8fF
C1606 n_633 gnd! 185.2fF
C1607 n_102 gnd! 2422.7fF
C1608 n_1129 gnd! 2108.2fF
C1609 n_1399 gnd! 1920.6fF
C1610 op_T2_zp_zp_idx gnd! 1444.7fF
C1611 op_T3_jsr gnd! 1885.2fF
C1612 op_sta_cmp gnd! 1838.9fF
C1613 op_shift_right gnd! 1390.2fF
C1614 op_T2_brk gnd! 1798.9fF
C1615 op_T2_pha gnd! 1878.4fF
C1616 op_T0_shift_right_a gnd! 1649.9fF
C1617 op_T4_abs_idx gnd! 1342.2fF
C1618 op_T0_bit gnd! 1645.2fF
C1619 op_branch_done gnd! 2400.2fF
C1620 op_T5_ind_y gnd! 1433.4fF
C1621 op_T0_and gnd! 1344.6fF
C1622 op_T0_shift_a gnd! 1896.0fF
C1623 op_T0_tax gnd! 1530.0fF
C1624 op_T0_acc gnd! 1243.5fF
C1625 op_T0_tay gnd! 1541.0fF
C1626 op_T0_pla gnd! 1692.5fF
C1627 op_T0_lda gnd! 1471.9fF
C1628 op_T__shift_a gnd! 1600.2fF
C1629 op_T0_txa gnd! 1673.4fF
C1630 op_T__ora_and_eor_adc gnd! 1397.2fF
C1631 n_1456 gnd! 362.4fF
C1632 op_T__adc_sbc gnd! 1481.0fF
C1633 op_T2_stack_access gnd! 1765.2fF
C1634 op_T0_tya gnd! 1775.5fF
C1635 op_shift gnd! 1523.4fF
C1636 op_T5_jsr gnd! 2323.1fF
C1637 op_rol_ror gnd! 1463.4fF
C1638 op_T0_sbc gnd! 2285.0fF
C1639 op_T3_jmp gnd! 1764.4fF
C1640 op_T0_adc_sbc gnd! 1862.0fF
C1641 op_T0_cpx_cpy_inx_iny gnd! 1468.0fF
C1642 op_T0_cmp gnd! 1410.3fF
C1643 op_rti_rts gnd! 2259.2fF
C1644 op_T2_jsr gnd! 2332.8fF
C1645 op_T4_ind_x gnd! 1726.0fF
C1646 x_op_T3_ind_y gnd! 1442.7fF
C1647 op_plp_pla gnd! 1538.3fF
C1648 op_inc_nop gnd! 1484.5fF
C1649 op_T2_ind_y gnd! 1475.0fF
C1650 op_T3_abs_idx gnd! 1295.1fF
C1651 op_T3_ind_x gnd! 1616.4fF
C1652 op_T4_ind_y gnd! 1405.8fF
C1653 op_T4_brk_jsr gnd! 1764.2fF
C1654 op_T4_rti gnd! 1719.6fF
C1655 op_T2_stack gnd! 2194.0fF
C1656 op_T3_stack_bit_jmp gnd! 1385.0fF
C1657 op_T2_ADL_ADD gnd! 1421.2fF
C1658 op_T0 gnd! 1108.6fF
C1659 op_T2_abs gnd! 1679.6fF
C1660 op_T0_ora gnd! 1698.6fF
C1661 op_T0_eor gnd! 1732.6fF
C1662 op_jmp gnd! 1862.2fF
C1663 op_ror gnd! 1689.1fF
C1664 op_T2 gnd! 2016.3fF
C1665 op_T3_plp_pla gnd! 1676.4fF
C1666 op_T0_php_pha gnd! 1669.3fF
C1667 op_T5_rti gnd! 2807.4fF
C1668 op_T4_rts gnd! 1879.8fF
C1669 op_T0_jsr gnd! 2064.6fF
C1670 op_T5_brk gnd! 2103.6fF
C1671 op_T0_tay_ldy_not_idx gnd! 1421.3fF
C1672 op_T__iny_dey gnd! 1606.3fF
C1673 op_T__inx gnd! 1699.1fF
C1674 op_T0_ldy_mem gnd! 1461.3fF
C1675 op_T0_tsx gnd! 1824.4fF
C1676 op_T0_ldx_tax_tsx gnd! 1389.6fF
C1677 op_T__dex gnd! 1509.8fF
C1678 op_from_x gnd! 2064.0fF
C1679 op_T0_txs gnd! 2432.5fF
C1680 op_T0_dex gnd! 1522.3fF
C1681 op_T2_ind_x gnd! 1543.8fF
C1682 op_T0_cpx_inx gnd! 1462.1fF
C1683 x_op_T0_txa gnd! 1678.9fF
C1684 op_T2_idx_x_xy gnd! 1719.7fF
C1685 op_T0_cpy_iny gnd! 1437.3fF
C1686 op_xy gnd! 1549.7fF
C1687 op_T0_iny_dey gnd! 1535.6fF
C1688 x_op_T0_tya gnd! 1787.7fF
C1689 op_T3_ind_y gnd! 1475.3fF
C1690 op_T2_abs_y gnd! 1427.7fF
C1691 n_1606 gnd! 227.2fF
C1692 _t4 gnd! 4005.8fF
C1693 op_sty_cpy_mem gnd! 1777.9fF
C1694 n_913 gnd! 486.8fF
C1695 n_1699 gnd! 174.2fF
C1696 n_1069 gnd! 4145.8fF
C1697 n_1274 gnd! 237.2fF
C1698 n_1024 gnd! 920.4fF
C1699 n_94 gnd! 215.0fF
C1700 n_1650 gnd! 730.6fF
C1701 n_1105 gnd! 2889.2fF
C1702 n_1715 gnd! 2108.2fF
C1703 n_1467 gnd! 2618.8fF
C1704 n_358 gnd! 2308.7fF
C1705 n_1696 gnd! 2046.4fF
C1706 so gnd! 4874.6fF
C1707 n_127 gnd! 2180.5fF
C1708 n_1395 gnd! 371.6fF
C1709 n_742 gnd! 114.8fF
C1710 n_975 gnd! 495.6fF
C1711 n_886 gnd! 114.8fF
C1712 n_995 gnd! 524.8fF
C1713 n_854 gnd! 796.4fF
C1714 n_312 gnd! 792.4fF
C1715 Reset0 gnd! 6836.8fF
C1716 clk2out gnd! 6771.0fF
C1717 n_603 gnd! 1371.4fF
C1718 n_47 gnd! 205.8fF
C1719 n_865 gnd! 201.8fF
C1720 n_420 gnd! 528.2fF
C1721 n_1449 gnd! 3413.0fF
C1722 n_958 gnd! 1048.0fF
C1723 clk0 gnd! 7799.9fF
C1724 res gnd! 4096.7fF
C1725 n_519 gnd! 2691.0fF
C1726 n_135 gnd! 2919.7fF
C1727 n_670 gnd! 2516.0fF
C1728 n_747 gnd! 2777.0fF
C1729 nIRQP gnd! 2631.4fF
C1730 IRQP gnd! 332.8fF
C1731 n_806 gnd! 1446.4fF
C1732 n_431 gnd! 294.4fF
C1733 n_330 gnd! 767.4fF
C1734 n_881 gnd! 357.6fF
C1735 n_538 gnd! 428.2fF
C1736 n_807 gnd! 620.0fF
C1737 n_1599 gnd! 840.0fF
C1738 n_346 gnd! 114.8fF
C1739 nNMIP gnd! 512.2fF
C1740 pipeT3out gnd! 487.6fF
C1741 n_1366 gnd! 498.2fF
C1742 n_188 gnd! 1098.0fF
C1743 n_1357 gnd! 4410.1fF
C1744 n_891 gnd! 214.4fF
C1745 n_284 gnd! 446.6fF
C1746 NMIP gnd! 747.8fF
C1747 _t5 gnd! 4572.8fF
C1748 cclk gnd! 100774.0fF
C1749 n_472 gnd! 576.6fF
C1750 cp1 gnd! 58835.8fF
C1751 n_378 gnd! 793.6fF
C1752 n_18 gnd! 263.4fF
C1753 pipeT5out gnd! 315.2fF
C1754 n_468 gnd! 522.6fF
C1755 n_395 gnd! 376.8fF
C1756 n_16 gnd! 1524.1fF
C1757 pipeT4out gnd! 488.4fF
C1758 n_1703 gnd! 610.8fF
C1759 notRdy0 gnd! 12415.5fF
C1760 n_1615 gnd! 510.4fF
C1761 n_645 gnd! 1638.4fF
C1762 Vdd gnd! 399097.0fF
C1763 n_1392 gnd! 813.2fF
C1764 clk1out gnd! 8088.6fF
C1765 n_1417 gnd! 3277.2fF
C1766 irq gnd! 3731.8fF
C1767 rdy gnd! 4320.9fF
C1768 nmi gnd! 3889.9fF
