`include "common.h"

module chip_6502(
  input eclk, ereset,
  output ab0,
  output ab1,
  output ab2,
  output ab3,
  output ab4,
  output ab5,
  output ab6,
  output ab7,
  output ab8,
  output ab9,
  output ab10,
  output ab11,
  output ab12,
  output ab13,
  output ab14,
  output ab15,
  input db0_i,
  output db0_o,
  output db0_t,
  input db1_i,
  output db1_o,
  output db1_t,
  input db2_i,
  output db2_o,
  output db2_t,
  input db3_i,
  output db3_o,
  output db3_t,
  input db4_i,
  output db4_o,
  output db4_t,
  input db5_i,
  output db5_o,
  output db5_t,
  input db6_i,
  output db6_o,
  output db6_t,
  input db7_i,
  output db7_o,
  output db7_t,
  input res,
  output rw,
  output sync,
  input so,
  input clk0,
  output clk1out,
  output clk2out,
  input rdy,
  input nmi,
  input irq
);

  wire signed [`W-1:0] dor5_port_3, dor5_port_4, dor5_v;
  wire signed [`W-1:0] dor4_port_3, dor4_port_4, dor4_v;
  wire signed [`W-1:0] dor7_port_0, dor7_port_4, dor7_v;
  wire signed [`W-1:0] dor6_port_2, dor6_port_4, dor6_v;
  wire signed [`W-1:0] dor1_port_0, dor1_port_4, dor1_v;
  wire signed [`W-1:0] dor0_port_0, dor0_port_4, dor0_v;
  wire signed [`W-1:0] dor3_port_3, dor3_port_4, dor3_v;
  wire signed [`W-1:0] dor2_port_3, dor2_port_4, dor2_v;
  wire signed [`W-1:0] _DBZ_port_2, _DBZ_port_0, _DBZ_v;
  wire signed [`W-1:0] _DBE_port_3, _DBE_port_5, _DBE_v;
  wire signed [`W-1:0] n_1714_port_2, n_1714_port_1, n_1714_v;
  wire signed [`W-1:0] n_1715_port_2, n_1715_port_3, n_1715_v;
  wire signed [`W-1:0] n_1716_port_6, n_1716_port_5, n_1716_v;
  wire signed [`W-1:0] n_1717_port_8, n_1717_port_12, n_1717_v;
  wire signed [`W-1:0] n_1247_port_13, n_1247_port_0, n_1247_v;
  wire signed [`W-1:0] n_1244_port_2, n_1244_port_1, n_1244_v;
  wire signed [`W-1:0] n_1245_port_2, n_1245_port_1, n_1245_v;
  wire signed [`W-1:0] n_1718_port_2, n_1718_port_1, n_1718_v;
  wire signed [`W-1:0] n_1719_port_2, n_1719_port_0, n_1719_v;
  wire signed [`W-1:0] _ABL7_port_3, _ABL7_port_1, _ABL7_v;
  wire signed [`W-1:0] _ABL6_port_3, _ABL6_port_1, _ABL6_v;
  wire signed [`W-1:0] _ABL5_port_3, _ABL5_port_0, _ABL5_v;
  wire signed [`W-1:0] _ABL3_port_3, _ABL3_port_0, _ABL3_v;
  wire signed [`W-1:0] _ABL2_port_2, _ABL2_port_3, _ABL2_v;
  wire signed [`W-1:0] _ABL1_port_2, _ABL1_port_3, _ABL1_v;
  wire signed [`W-1:0] _ABL0_port_2, _ABL0_port_3, _ABL0_v;
  wire signed [`W-1:0] dpc5_SADL_port_0, dpc5_SADL_port_7, dpc5_SADL_v;
  wire signed [`W-1:0] n_604_port_10, n_604_port_15, n_604_v;
  wire signed [`W-1:0] n_600_port_1, n_600_port_4, n_600_v;
  wire signed [`W-1:0] n_602_port_2, n_602_port_0, n_602_v;
  wire signed [`W-1:0] n_603_port_2, n_603_port_1, n_603_v;
  wire signed [`W-1:0] n_608_port_2, n_608_port_0, n_608_v;
  wire signed [`W-1:0] n_609_port_6, n_609_port_4, n_609_v;
  wire signed [`W-1:0] pd6_clearIR_port_3, pd6_clearIR_port_4, pd6_clearIR_v;
  wire signed [`W-1:0] n_462_port_2, n_462_port_3, n_462_v;
  wire signed [`W-1:0] n_465_port_2, n_465_port_0, n_465_port_1, n_465_v;
  wire signed [`W-1:0] n_466_port_6, n_466_port_4, n_466_v;
  wire signed [`W-1:0] n_467_port_6, n_467_port_4, n_467_v;
  wire signed [`W-1:0] n_468_port_3, n_468_port_6, n_468_v;
  wire signed [`W-1:0] op_T4_brk_port_10, op_T4_brk_port_12, op_T4_brk_v;
  wire signed [`W-1:0] rw_port_0, rw_port_1, rw_v;
  wire signed [`W-1:0] x_op_T3_plp_pla_port_8, x_op_T3_plp_pla_port_10, x_op_T3_plp_pla_v;
  wire signed [`W-1:0] idl7_port_2, idl7_port_0, idl7_port_1, idl7_v;
  wire signed [`W-1:0] idl6_port_2, idl6_port_0, idl6_port_1, idl6_v;
  wire signed [`W-1:0] idl5_port_2, idl5_port_0, idl5_port_1, idl5_v;
  wire signed [`W-1:0] idl4_port_2, idl4_port_0, idl4_port_1, idl4_v;
  wire signed [`W-1:0] idl3_port_2, idl3_port_0, idl3_port_1, idl3_v;
  wire signed [`W-1:0] idl2_port_2, idl2_port_0, idl2_port_1, idl2_v;
  wire signed [`W-1:0] idl1_port_2, idl1_port_0, idl1_port_1, idl1_v;
  wire signed [`W-1:0] idl0_port_2, idl0_port_0, idl0_port_1, idl0_v;
  wire signed [`W-1:0] n_1523_port_2, n_1523_port_3, n_1523_v;
  wire signed [`W-1:0] n_1521_port_2, n_1521_port_1, n_1521_v;
  wire signed [`W-1:0] n_1526_port_2, n_1526_port_1, n_1526_v;
  wire signed [`W-1:0] n_733_port_2, n_733_port_3, n_733_port_0, n_733_port_1, n_733_v;
  wire signed [`W-1:0] dpc20_ADDSB06_port_0, dpc20_ADDSB06_port_5, dpc20_ADDSB06_v;
  wire signed [`W-1:0] n_1389_port_2, n_1389_port_3, n_1389_port_0, n_1389_port_1, n_1389_port_4, n_1389_v;
  wire signed [`W-1:0] n_1387_port_2, n_1387_port_3, n_1387_port_0, n_1387_port_1, n_1387_v;
  wire signed [`W-1:0] n_1386_port_2, n_1386_port_3, n_1386_v;
  wire signed [`W-1:0] n_1383_port_2, n_1383_port_0, n_1383_port_1, n_1383_v;
  wire signed [`W-1:0] n_1380_port_4, n_1380_port_5, n_1380_v;
  wire signed [`W-1:0] n_917_port_3, n_917_port_5, n_917_v;
  wire signed [`W-1:0] x6_port_0, x6_port_1, x6_v;
  wire signed [`W-1:0] n_819_port_6, n_819_port_4, n_819_v;
  wire signed [`W-1:0] n_818_port_4, n_818_port_5, n_818_v;
  wire signed [`W-1:0] n_811_port_7, n_811_port_5, n_811_v;
  wire signed [`W-1:0] n_810_port_3, n_810_port_4, n_810_v;
  wire signed [`W-1:0] n_813_port_3, n_813_port_4, n_813_v;
  wire signed [`W-1:0] n_812_port_3, n_812_port_4, n_812_v;
  wire signed [`W-1:0] n_815_port_2, n_815_port_0, n_815_v;
  wire signed [`W-1:0] irq_port_2, irq_v;
  wire signed [`W-1:0] ir0_port_3, ir0_port_4, ir0_v;
  wire signed [`W-1:0] ir1_port_2, ir1_port_3, ir1_v;
  wire signed [`W-1:0] ir2_port_72, ir2_port_0, ir2_v;
  wire signed [`W-1:0] ir3_port_1, ir3_port_41, ir3_v;
  wire signed [`W-1:0] ir4_port_70, ir4_port_68, ir4_v;
  wire signed [`W-1:0] ir5_port_0, ir5_port_33, ir5_v;
  wire signed [`W-1:0] ir6_port_42, ir6_port_43, ir6_v;
  wire signed [`W-1:0] ir7_port_59, ir7_port_60, ir7_v;
  wire signed [`W-1:0] n_1267_port_2, n_1267_port_3, n_1267_port_0, n_1267_v;
  wire signed [`W-1:0] n_1260_port_2, n_1260_port_3, n_1260_v;
  wire signed [`W-1:0] op_T__inx_port_9, op_T__inx_port_11, op_T__inx_v;
  wire signed [`W-1:0] n_5_port_2, n_5_port_0, n_5_v;
  wire signed [`W-1:0] n_6_port_4, n_6_port_5, n_6_v;
  wire signed [`W-1:0] n_7_port_2, n_7_port_4, n_7_v;
  wire signed [`W-1:0] n_3_port_2, n_3_port_3, n_3_port_0, n_3_port_1, n_3_port_4, n_3_v;
  wire signed [`W-1:0] aluanandb0_port_9, aluanandb0_port_3, aluanandb0_port_5, aluanandb0_v;
  wire signed [`W-1:0] aluanandb1_port_0, aluanandb1_port_1, aluanandb1_port_4, aluanandb1_port_5, aluanandb1_v;
  wire signed [`W-1:0] n_1240_port_2, n_1240_port_1, n_1240_v;
  wire signed [`W-1:0] n_1711_port_2, n_1711_port_1, n_1711_v;
  wire signed [`W-1:0] n_1712_port_4, n_1712_port_5, n_1712_v;
  wire signed [`W-1:0] op_T0_php_pha_port_8, op_T0_php_pha_port_10, op_T0_php_pha_v;
  wire signed [`W-1:0] dasb6_port_3, dasb6_port_0, dasb6_port_5, dasb6_v;
  wire signed [`W-1:0] dasb5_port_3, dasb5_port_1, dasb5_port_5, dasb5_v;
  wire signed [`W-1:0] dasb3_port_3, dasb3_port_1, dasb3_port_5, dasb3_v;
  wire signed [`W-1:0] dasb2_port_3, dasb2_port_1, dasb2_port_5, dasb2_v;
  wire signed [`W-1:0] dasb1_port_3, dasb1_port_0, dasb1_port_5, dasb1_v;
  wire signed [`W-1:0] n_662_port_2, n_662_port_0, n_662_v;
  wire signed [`W-1:0] n_664_port_2, n_664_port_1, n_664_v;
  wire signed [`W-1:0] alu4_port_2, alu4_port_3, alu4_port_0, alu4_port_1, alu4_v;
  wire signed [`W-1:0] alu5_port_3, alu5_port_0, alu5_port_1, alu5_port_4, alu5_v;
  wire signed [`W-1:0] alu6_port_2, alu6_port_0, alu6_port_1, alu6_port_4, alu6_v;
  wire signed [`W-1:0] alu7_port_2, alu7_port_3, alu7_port_0, alu7_port_1, alu7_v;
  wire signed [`W-1:0] alu0_port_2, alu0_port_3, alu0_port_0, alu0_port_1, alu0_v;
  wire signed [`W-1:0] alu1_port_3, alu1_port_0, alu1_port_1, alu1_port_4, alu1_v;
  wire signed [`W-1:0] alu2_port_3, alu2_port_0, alu2_port_1, alu2_port_4, alu2_v;
  wire signed [`W-1:0] alu3_port_2, alu3_port_3, alu3_port_0, alu3_port_1, alu3_v;
  wire signed [`W-1:0] _ABL4_port_3, _ABL4_port_1, _ABL4_v;
  wire signed [`W-1:0] n_488_port_2, n_488_port_3, n_488_port_0, n_488_port_1, n_488_port_4, n_488_v;
  wire signed [`W-1:0] n_484_port_2, n_484_port_3, n_484_v;
  wire signed [`W-1:0] n_485_port_2, n_485_port_1, n_485_v;
  wire signed [`W-1:0] n_480_port_2, n_480_port_4, n_480_v;
  wire signed [`W-1:0] n_481_port_2, n_481_port_3, n_481_port_0, n_481_port_1, n_481_port_4, n_481_v;
  wire signed [`W-1:0] PD_xxx010x1_port_6, PD_xxx010x1_port_5, PD_xxx010x1_v;
  wire signed [`W-1:0] op_shift_port_4, op_shift_port_5, op_shift_v;
  wire signed [`W-1:0] op_xy_port_6, op_xy_port_5, op_xy_v;
  wire signed [`W-1:0] op_T0_cld_sed_port_8, op_T0_cld_sed_port_9, op_T0_cld_sed_v;
  wire signed [`W-1:0] n_327_port_3, n_327_port_4, n_327_v;
  wire signed [`W-1:0] n_326_port_2, n_326_port_3, n_326_port_0, n_326_port_1, n_326_port_4, n_326_v;
  wire signed [`W-1:0] _AxB_0__C0in_port_3, _AxB_0__C0in_port_4, _AxB_0__C0in_v;
  wire signed [`W-1:0] n_321_port_2, n_321_port_3, n_321_v;
  wire signed [`W-1:0] n_320_port_3, n_320_port_0, n_320_v;
  wire signed [`W-1:0] n_1105_port_2, n_1105_port_0, n_1105_v;
  wire signed [`W-1:0] n_1107_port_7, n_1107_port_10, n_1107_v;
  wire signed [`W-1:0] n_1106_port_8, n_1106_port_12, n_1106_v;
  wire signed [`W-1:0] n_1101_port_2, n_1101_port_3, n_1101_v;
  wire signed [`W-1:0] n_1100_port_2, n_1100_port_3, n_1100_port_0, n_1100_v;
  wire signed [`W-1:0] n_1109_port_9, n_1109_port_5, n_1109_v;
  wire signed [`W-1:0] pd4_clearIR_port_8, pd4_clearIR_port_6, pd4_clearIR_v;
  wire signed [`W-1:0] op_ror_port_6, op_ror_port_5, op_ror_v;
  wire signed [`W-1:0] dpc6_SBS_port_11, dpc6_SBS_port_12, dpc6_SBS_v;
  wire signed [`W-1:0] n_345_port_4, n_345_port_10, n_345_v;
  wire signed [`W-1:0] n_347_port_8, n_347_port_9, n_347_v;
  wire signed [`W-1:0] n_340_port_2, n_340_port_0, n_340_v;
  wire signed [`W-1:0] n_831_port_2, n_831_port_3, n_831_port_0, n_831_port_1, n_831_port_4, n_831_v;
  wire signed [`W-1:0] n_830_port_4, n_830_port_5, n_830_v;
  wire signed [`W-1:0] n_839_port_2, n_839_port_1, n_839_v;
  wire signed [`W-1:0] n_838_port_2, n_838_port_0, n_838_v;
  wire signed [`W-1:0] op_T0_ldy_mem_port_8, op_T0_ldy_mem_port_7, op_T0_ldy_mem_v;
  wire signed [`W-1:0] D1x1_port_6, D1x1_port_5, D1x1_v;
  wire signed [`W-1:0] s3_port_0, s3_port_1, s3_v;
  wire signed [`W-1:0] s2_port_0, s2_port_1, s2_v;
  wire signed [`W-1:0] s1_port_0, s1_port_1, s1_v;
  wire signed [`W-1:0] s0_port_0, s0_port_1, s0_v;
  wire signed [`W-1:0] s7_port_2, s7_port_0, s7_v;
  wire signed [`W-1:0] s6_port_0, s6_port_1, s6_v;
  wire signed [`W-1:0] s5_port_0, s5_port_1, s5_v;
  wire signed [`W-1:0] s4_port_0, s4_port_1, s4_v;
  wire signed [`W-1:0] so_port_2, so_port_3, so_v;
  wire signed [`W-1:0] dpc15_ANDS_port_9, dpc15_ANDS_port_0, dpc15_ANDS_v;
  wire signed [`W-1:0] n_1585_port_2, n_1585_port_1, n_1585_v;
  wire signed [`W-1:0] n_1586_port_2, n_1586_port_1, n_1586_v;
  wire signed [`W-1:0] _TWOCYCLE_port_7, _TWOCYCLE_port_4, _TWOCYCLE_v;
  wire signed [`W-1:0] dpc27_SBADH_port_9, dpc27_SBADH_port_0, dpc27_SBADH_v;
  wire signed [`W-1:0] pd3_clearIR_port_6, pd3_clearIR_port_4, pd3_clearIR_v;
  wire signed [`W-1:0] n_649_port_0, n_649_port_7, n_649_port_5, n_649_v;
  wire signed [`W-1:0] n_138_port_2, n_138_port_0, n_138_port_1, n_138_v;
  wire signed [`W-1:0] n_139_port_2, n_139_port_1, n_139_v;
  wire signed [`W-1:0] n_641_port_3, n_641_port_0, n_641_v;
  wire signed [`W-1:0] n_642_port_3, n_642_port_0, n_642_port_1, n_642_v;
  wire signed [`W-1:0] n_643_port_3, n_643_port_4, n_643_v;
  wire signed [`W-1:0] n_132_port_2, n_132_port_1, n_132_v;
  wire signed [`W-1:0] n_645_port_2, n_645_port_3, n_645_v;
  wire signed [`W-1:0] n_646_port_8, n_646_port_2, n_646_v;
  wire signed [`W-1:0] n_647_port_3, n_647_port_5, n_647_v;
  wire signed [`W-1:0] n_1632_port_7, n_1632_port_4, n_1632_port_5, n_1632_v;
  wire signed [`W-1:0] n_1635_port_2, n_1635_port_1, n_1635_v;
  wire signed [`W-1:0] _AxB_6__C56_port_3, _AxB_6__C56_port_4, _AxB_6__C56_v;
  wire signed [`W-1:0] pd0_clearIR_port_8, pd0_clearIR_port_5, pd0_clearIR_v;
  wire signed [`W-1:0] op_T0_shift_a_port_8, op_T0_shift_a_port_11, op_T0_shift_a_v;
  wire signed [`W-1:0] __AxB7__C67_port_3, __AxB7__C67_port_4, __AxB7__C67_v;
  wire signed [`W-1:0] n_1439_port_2, n_1439_port_1, n_1439_v;
  wire signed [`W-1:0] _VEC_port_8, _VEC_port_5, _VEC_v;
  wire signed [`W-1:0] n_1129_port_4, n_1129_port_5, n_1129_v;
  wire signed [`W-1:0] n_1120_port_2, n_1120_port_1, n_1120_v;
  wire signed [`W-1:0] n_587_port_2, n_587_port_1, n_587_v;
  wire signed [`W-1:0] n_586_port_3, n_586_port_5, n_586_v;
  wire signed [`W-1:0] n_583_port_2, n_583_port_0, n_583_port_1, n_583_v;
  wire signed [`W-1:0] n_582_port_2, n_582_port_3, n_582_v;
  wire signed [`W-1:0] n_588_port_2, n_588_port_0, n_588_v;
  wire signed [`W-1:0] op_rmw_port_2, op_rmw_port_0, op_rmw_v;
  wire signed [`W-1:0] n_366_port_3, n_366_port_5, n_366_v;
  wire signed [`W-1:0] n_368_port_8, n_368_port_7, n_368_v;
  wire signed [`W-1:0] op_jmp_port_8, op_jmp_port_7, op_jmp_v;
  wire signed [`W-1:0] C12_port_2, C12_port_3, C12_v;
  wire signed [`W-1:0] n_1433_port_6, n_1433_port_4, n_1433_v;
  wire signed [`W-1:0] op_shift_right_port_4, op_shift_right_port_5, op_shift_right_v;
  wire signed [`W-1:0] op_EORS_port_2, op_EORS_port_3, op_EORS_v;
  wire signed [`W-1:0] x_op_T__adc_sbc_port_8, x_op_T__adc_sbc_port_6, x_op_T__adc_sbc_v;
  wire signed [`W-1:0] n_1631_port_2, n_1631_port_3, n_1631_v;
  wire signed [`W-1:0] notir0_port_0, notir0_port_1, notir0_port_28, notir0_v;
  wire signed [`W-1:0] notir1_port_21, notir1_port_23, notir1_port_22, notir1_v;
  wire signed [`W-1:0] notir2_port_19, notir2_port_0, notir2_port_20, notir2_v;
  wire signed [`W-1:0] notir3_port_51, notir3_port_0, notir3_port_1, notir3_v;
  wire signed [`W-1:0] notir4_port_25, notir4_port_24, notir4_port_26, notir4_v;
  wire signed [`W-1:0] notir5_port_36, notir5_port_37, notir5_port_0, notir5_v;
  wire signed [`W-1:0] notir6_port_0, notir6_port_1, notir6_port_39, notir6_v;
  wire signed [`W-1:0] notir7_port_34, notir7_port_35, notir7_port_33, notir7_v;
  wire signed [`W-1:0] n_93_port_2, n_93_port_0, n_93_v;
  wire signed [`W-1:0] n_90_port_3, n_90_port_4, n_90_v;
  wire signed [`W-1:0] n_91_port_3, n_91_port_0, n_91_v;
  wire signed [`W-1:0] op_lsr_ror_dec_inc_port_3, op_lsr_ror_dec_inc_port_4, op_lsr_ror_dec_inc_v;
  wire signed [`W-1:0] n_110_port_2, n_110_port_1, n_110_v;
  wire signed [`W-1:0] n_111_port_2, n_111_port_1, n_111_v;
  wire signed [`W-1:0] n_118_port_2, n_118_port_1, n_118_v;
  wire signed [`W-1:0] n_119_port_3, n_119_port_0, n_119_v;
  wire signed [`W-1:0] cp1_port_75, cp1_port_50, cp1_v;
  wire signed [`W-1:0] a3_port_0, a3_port_1, a3_v;
  wire signed [`W-1:0] a6_port_2, a6_port_0, a6_v;
  wire signed [`W-1:0] n_696_port_3, n_696_port_5, n_696_v;
  wire signed [`W-1:0] n_1199_port_2, n_1199_port_0, n_1199_v;
  wire signed [`W-1:0] n_930_port_3, n_930_port_4, n_930_v;
  wire signed [`W-1:0] DA_AxB2_port_3, DA_AxB2_port_5, DA_AxB2_v;
  wire signed [`W-1:0] n_1479_port_0, n_1479_port_1, n_1479_v;
  wire signed [`W-1:0] sync_port_0, sync_port_1, sync_v;
  wire signed [`W-1:0] n_1499_port_3, n_1499_port_0, n_1499_v;
  wire signed [`W-1:0] n_1325_port_2, n_1325_port_4, n_1325_v;
  wire signed [`W-1:0] n_1496_port_2, n_1496_port_3, n_1496_port_0, n_1496_port_1, n_1496_port_4, n_1496_v;
  wire signed [`W-1:0] n_1495_port_8, n_1495_port_4, n_1495_v;
  wire signed [`W-1:0] n_1492_port_3, n_1492_port_0, n_1492_v;
  wire signed [`W-1:0] n_1323_port_2, n_1323_port_0, n_1323_v;
  wire signed [`W-1:0] n_1141_port_2, n_1141_port_1, n_1141_v;
  wire signed [`W-1:0] n_568_port_2, n_568_port_1, n_568_v;
  wire signed [`W-1:0] n_565_port_2, n_565_port_0, n_565_v;
  wire signed [`W-1:0] n_564_port_2, n_564_port_3, n_564_port_0, n_564_port_1, n_564_v;
  wire signed [`W-1:0] n_567_port_0, n_567_port_4, n_567_v;
  wire signed [`W-1:0] n_566_port_8, n_566_port_4, n_566_v;
  wire signed [`W-1:0] __AxBxC_6_port_3, __AxBxC_6_port_1, __AxBxC_6_port_5, __AxBxC_6_v;
  wire signed [`W-1:0] __AxBxC_7_port_3, __AxBxC_7_port_0, __AxBxC_7_port_5, __AxBxC_7_v;
  wire signed [`W-1:0] __AxBxC_4_port_2, __AxBxC_4_port_3, __AxBxC_4_port_5, __AxBxC_4_v;
  wire signed [`W-1:0] __AxBxC_5_port_3, __AxBxC_5_port_1, __AxBxC_5_port_5, __AxBxC_5_v;
  wire signed [`W-1:0] __AxBxC_2_port_3, __AxBxC_2_port_1, __AxBxC_2_port_5, __AxBxC_2_v;
  wire signed [`W-1:0] __AxBxC_3_port_3, __AxBxC_3_port_1, __AxBxC_3_port_5, __AxBxC_3_v;
  wire signed [`W-1:0] __AxBxC_0_port_2, __AxBxC_0_port_3, __AxBxC_0_port_5, __AxBxC_0_v;
  wire signed [`W-1:0] __AxBxC_1_port_3, __AxBxC_1_port_1, __AxBxC_1_port_5, __AxBxC_1_v;
  wire signed [`W-1:0] n_300_port_8, n_300_port_7, n_300_v;
  wire signed [`W-1:0] n_304_port_2, n_304_port_3, n_304_port_0, n_304_port_1, n_304_port_4, n_304_v;
  wire signed [`W-1:0] n_307_port_6, n_307_port_4, n_307_v;
  wire signed [`W-1:0] n_306_port_2, n_306_port_0, n_306_v;
  wire signed [`W-1:0] aluaorb0_port_2, aluaorb0_port_1, aluaorb0_v;
  wire signed [`W-1:0] x_op_T0_tya_port_9, x_op_T0_tya_port_10, x_op_T0_tya_v;
  wire signed [`W-1:0] x_op_T4_ind_y_port_7, x_op_T4_ind_y_port_10, x_op_T4_ind_y_v;
  wire signed [`W-1:0] pclp0_port_2, pclp0_port_1, pclp0_v;
  wire signed [`W-1:0] pclp2_port_2, pclp2_port_1, pclp2_v;
  wire signed [`W-1:0] pclp4_port_2, pclp4_port_0, pclp4_v;
  wire signed [`W-1:0] pclp6_port_2, pclp6_port_0, pclp6_v;
  wire signed [`W-1:0] op_T3_branch_port_8, op_T3_branch_port_7, op_T3_branch_v;
  wire signed [`W-1:0] ab12_port_0, ab12_port_1, ab12_v;
  wire signed [`W-1:0] ab13_port_0, ab13_port_1, ab13_v;
  wire signed [`W-1:0] ab10_port_0, ab10_port_1, ab10_v;
  wire signed [`W-1:0] ab11_port_0, ab11_port_1, ab11_v;
  wire signed [`W-1:0] n_79_port_2, n_79_port_1, n_79_v;
  wire signed [`W-1:0] ab14_port_0, ab14_port_1, ab14_v;
  wire signed [`W-1:0] ab15_port_0, ab15_port_1, ab15_v;
  wire signed [`W-1:0] n_75_port_2, n_75_port_0, n_75_v;
  wire signed [`W-1:0] n_70_port_3, n_70_port_4, n_70_v;
  wire signed [`W-1:0] n_71_port_2, n_71_port_0, n_71_v;
  wire signed [`W-1:0] n_72_port_2, n_72_port_3, n_72_port_0, n_72_port_1, n_72_port_4, n_72_v;
  wire signed [`W-1:0] n_1705_port_3, n_1705_port_4, n_1705_v;
  wire signed [`W-1:0] n_1256_port_2, n_1256_port_0, n_1256_v;
  wire signed [`W-1:0] op_T0_tya_port_9, op_T0_tya_port_11, op_T0_tya_v;
  wire signed [`W-1:0] n_172_port_2, n_172_port_3, n_172_v;
  wire signed [`W-1:0] n_176_port_3, n_176_port_4, n_176_v;
  wire signed [`W-1:0] n_177_port_2, n_177_port_0, n_177_port_1, n_177_v;
  wire signed [`W-1:0] n_797_port_2, n_797_port_1, n_797_v;
  wire signed [`W-1:0] n_794_port_1, n_794_port_4, n_794_v;
  wire signed [`W-1:0] n_795_port_2, n_795_port_0, n_795_v;
  wire signed [`W-1:0] n_790_port_7, n_790_port_5, n_790_v;
  wire signed [`W-1:0] n_798_port_1, n_798_port_4, n_798_v;
  wire signed [`W-1:0] n_1305_port_2, n_1305_port_1, n_1305_v;
  wire signed [`W-1:0] n_1304_port_3, n_1304_port_4, n_1304_v;
  wire signed [`W-1:0] n_1303_port_3, n_1303_port_7, n_1303_v;
  wire signed [`W-1:0] n_1301_port_2, n_1301_port_3, n_1301_port_0, n_1301_port_1, n_1301_port_4, n_1301_v;
  wire signed [`W-1:0] n_1300_port_2, n_1300_port_3, n_1300_v;
  wire signed [`W-1:0] n_1309_port_2, n_1309_port_3, n_1309_port_1, n_1309_v;
  wire signed [`W-1:0] n_330_port_7, n_330_port_4, n_330_v;
  wire signed [`W-1:0] n_332_port_2, n_332_port_3, n_332_port_0, n_332_port_1, n_332_port_4, n_332_v;
  wire signed [`W-1:0] n_1166_port_2, n_1166_port_3, n_1166_v;
  wire signed [`W-1:0] n_1169_port_2, n_1169_port_3, n_1169_port_0, n_1169_port_1, n_1169_v;
  wire signed [`W-1:0] PD_1xx000x0_port_6, PD_1xx000x0_port_7, PD_1xx000x0_v;
  wire signed [`W-1:0] n_548_port_2, n_548_port_0, n_548_v;
  wire signed [`W-1:0] op_T2_brk_port_9, op_T2_brk_port_10, op_T2_brk_v;
  wire signed [`W-1:0] n_543_port_3, n_543_port_0, n_543_v;
  wire signed [`W-1:0] n_541_port_3, n_541_port_1, n_541_v;
  wire signed [`W-1:0] n_544_port_2, n_544_port_1, n_544_v;
  wire signed [`W-1:0] C56_port_3, C56_port_0, C56_v;
  wire signed [`W-1:0] n_890_port_2, n_890_port_1, n_890_v;
  wire signed [`W-1:0] n_322_port_2, n_322_port_1, n_322_v;
  wire signed [`W-1:0] n_896_port_2, n_896_port_1, n_896_v;
  wire signed [`W-1:0] n_329_port_3, n_329_port_0, n_329_v;
  wire signed [`W-1:0] xx_op_T5_jsr_port_9, xx_op_T5_jsr_port_11, xx_op_T5_jsr_v;
  wire signed [`W-1:0] PD_xxxx10x0_port_6, PD_xxxx10x0_port_5, PD_xxxx10x0_v;
  wire signed [`W-1:0] n_1028_port_2, n_1028_port_0, n_1028_v;
  wire signed [`W-1:0] dpc24_ACSB_port_1, dpc24_ACSB_port_12, dpc24_ACSB_v;
  wire signed [`W-1:0] n_152_port_6, n_152_port_5, n_152_v;
  wire signed [`W-1:0] n_154_port_2, n_154_port_3, n_154_v;
  wire signed [`W-1:0] rdy_port_2, rdy_port_3, rdy_v;
  wire signed [`W-1:0] n_1347_port_8, n_1347_port_7, n_1347_v;
  wire signed [`W-1:0] op_ORS_port_2, op_ORS_port_3, op_ORS_v;
  wire signed [`W-1:0] n_1346_port_3, n_1346_port_0, n_1346_v;
  wire signed [`W-1:0] _AxB_2__C12_port_3, _AxB_2__C12_port_4, _AxB_2__C12_v;
  wire signed [`W-1:0] n_1364_port_3, n_1364_port_0, n_1364_v;
  wire signed [`W-1:0] n_1369_port_2, n_1369_port_3, n_1369_v;
  wire signed [`W-1:0] n_1368_port_4, n_1368_port_5, n_1368_v;
  wire signed [`W-1:0] clearIR_port_9, clearIR_port_18, clearIR_v;
  wire signed [`W-1:0] op_T__cpx_cpy_imm_zp_port_8, op_T__cpx_cpy_imm_zp_port_7, op_T__cpx_cpy_imm_zp_v;
  wire signed [`W-1:0] n_1187_port_2, n_1187_port_0, n_1187_v;
  wire signed [`W-1:0] n_1181_port_3, n_1181_port_6, n_1181_v;
  wire signed [`W-1:0] n_1180_port_3, n_1180_port_4, n_1180_v;
  wire signed [`W-1:0] op_T5_mem_ind_idx_port_7, op_T5_mem_ind_idx_port_5, op_T5_mem_ind_idx_v;
  wire signed [`W-1:0] n_520_port_0, n_520_port_4, n_520_v;
  wire signed [`W-1:0] n_523_port_6, n_523_port_4, n_523_v;
  wire signed [`W-1:0] n_525_port_4, n_525_port_5, n_525_v;
  wire signed [`W-1:0] C78_port_2, C78_port_1, C78_v;
  wire signed [`W-1:0] dpc21_ADDADL_port_9, dpc21_ADDADL_port_0, dpc21_ADDADL_v;
  wire signed [`W-1:0] n_1592_port_2, n_1592_port_3, n_1592_port_0, n_1592_port_1, n_1592_port_4, n_1592_v;
  wire signed [`W-1:0] n_31_port_0, n_31_port_6, n_31_v;
  wire signed [`W-1:0] n_34_port_2, n_34_port_1, n_34_v;
  wire signed [`W-1:0] n_35_port_4, n_35_port_5, n_35_v;
  wire signed [`W-1:0] n_36_port_6, n_36_port_4, n_36_v;
  wire signed [`W-1:0] n_37_port_3, n_37_port_4, n_37_v;
  wire signed [`W-1:0] db1_port_1, db1_port_4, db1_port_5, db1_v;
  wire signed [`W-1:0] db0_port_1, db0_port_4, db0_port_5, db0_v;
  wire signed [`W-1:0] db3_port_2, db3_port_3, db3_port_5, db3_v;
  wire signed [`W-1:0] db2_port_2, db2_port_3, db2_port_5, db2_v;
  wire signed [`W-1:0] db5_port_0, db5_port_4, db5_port_5, db5_v;
  wire signed [`W-1:0] db4_port_3, db4_port_0, db4_port_5, db4_v;
  wire signed [`W-1:0] db7_port_3, db7_port_1, db7_port_5, db7_v;
  wire signed [`W-1:0] db6_port_0, db6_port_4, db6_port_5, db6_v;
  wire signed [`W-1:0] pchp5_port_2, pchp5_port_1, pchp5_v;
  wire signed [`W-1:0] pchp7_port_2, pchp7_port_0, pchp7_v;
  wire signed [`W-1:0] pchp1_port_2, pchp1_port_0, pchp1_v;
  wire signed [`W-1:0] pchp3_port_2, pchp3_port_0, pchp3_v;
  wire signed [`W-1:0] clk1out_port_0, clk1out_port_1, clk1out_v;
  wire signed [`W-1:0] _WR_port_8, _WR_port_7, _WR_v;
  wire signed [`W-1:0] n_1647_port_2, n_1647_port_3, n_1647_port_0, n_1647_port_1, n_1647_port_4, n_1647_v;
  wire signed [`W-1:0] n_1642_port_2, n_1642_port_4, n_1642_v;
  wire signed [`W-1:0] n_1643_port_3, n_1643_port_4, n_1643_v;
  wire signed [`W-1:0] n_1640_port_2, n_1640_port_0, n_1640_v;
  wire signed [`W-1:0] n_1641_port_2, n_1641_port_3, n_1641_port_1, n_1641_v;
  wire signed [`W-1:0] n_1649_port_11, n_1649_port_12, n_1649_v;
  wire signed [`W-1:0] _op_branch_bit6_port_0, _op_branch_bit6_port_4, _op_branch_bit6_v;
  wire signed [`W-1:0] _op_branch_bit7_port_1, _op_branch_bit7_port_4, _op_branch_bit7_v;
  wire signed [`W-1:0] n_1184_port_8, n_1184_port_4, n_1184_v;
  wire signed [`W-1:0] op_rol_ror_port_7, op_rol_ror_port_5, op_rol_ror_v;
  wire signed [`W-1:0] n_1491_port_2, n_1491_port_3, n_1491_port_0, n_1491_port_1, n_1491_v;
  wire signed [`W-1:0] n_201_port_3, n_201_port_1, n_201_v;
  wire signed [`W-1:0] n_206_port_3, n_206_port_0, n_206_port_5, n_206_v;
  wire signed [`W-1:0] clock1_port_68, clock1_port_40, clock1_v;
  wire signed [`W-1:0] clock2_port_12, clock2_port_13, clock2_v;
  wire signed [`W-1:0] n_1434_port_2, n_1434_port_0, n_1434_v;
  wire signed [`W-1:0] n_1344_port_2, n_1344_port_3, n_1344_port_0, n_1344_port_1, n_1344_port_4, n_1344_v;
  wire signed [`W-1:0] op_asl_rol_port_7, op_asl_rol_port_5, op_asl_rol_v;
  wire signed [`W-1:0] short_circuit_idx_add_port_7, short_circuit_idx_add_port_5, short_circuit_idx_add_v;
  wire signed [`W-1:0] n_507_port_2, n_507_port_3, n_507_v;
  wire signed [`W-1:0] n_506_port_4, n_506_port_5, n_506_v;
  wire signed [`W-1:0] n_504_port_2, n_504_port_3, n_504_v;
  wire signed [`W-1:0] n_503_port_2, n_503_port_0, n_503_v;
  wire signed [`W-1:0] n_501_port_4, n_501_port_5, n_501_v;
  wire signed [`W-1:0] x_op_T0_bit_port_8, x_op_T0_bit_port_9, x_op_T0_bit_v;
  wire signed [`W-1:0] n_16_port_0, n_16_port_5, n_16_v;
  wire signed [`W-1:0] n_17_port_6, n_17_port_5, n_17_v;
  wire signed [`W-1:0] n_14_port_4, n_14_port_5, n_14_v;
  wire signed [`W-1:0] n_10_port_6, n_10_port_4, n_10_v;
  wire signed [`W-1:0] n_11_port_9, n_11_port_6, n_11_v;
  wire signed [`W-1:0] n_1084_port_0, n_1084_port_6, n_1084_port_5, n_1084_v;
  wire signed [`W-1:0] n_1085_port_3, n_1085_port_6, n_1085_v;
  wire signed [`W-1:0] n_1087_port_3, n_1087_port_4, n_1087_v;
  wire signed [`W-1:0] n_1081_port_2, n_1081_port_3, n_1081_v;
  wire signed [`W-1:0] n_1082_port_5, n_1082_port_10, n_1082_v;
  wire signed [`W-1:0] n_1083_port_1, n_1083_port_7, n_1083_port_4, n_1083_v;
  wire signed [`W-1:0] n_1089_port_2, n_1089_port_1, n_1089_v;
  wire signed [`W-1:0] dpc35_PCHC_port_8, dpc35_PCHC_port_7, dpc35_PCHC_v;
  wire signed [`W-1:0] n_1265_port_2, n_1265_port_3, n_1265_v;
  wire signed [`W-1:0] n_1661_port_2, n_1661_port_3, n_1661_port_0, n_1661_port_1, n_1661_v;
  wire signed [`W-1:0] n_1662_port_3, n_1662_port_1, n_1662_v;
  wire signed [`W-1:0] n_1262_port_2, n_1262_port_3, n_1262_v;
  wire signed [`W-1:0] n_1668_port_2, n_1668_port_3, n_1668_port_0, n_1668_v;
  wire signed [`W-1:0] op_T2_abs_y_port_6, op_T2_abs_y_port_7, op_T2_abs_y_v;
  wire signed [`W-1:0] n_267_port_4, n_267_port_5, n_267_v;
  wire signed [`W-1:0] n_264_port_8, n_264_port_6, n_264_v;
  wire signed [`W-1:0] n_262_port_3, n_262_port_6, n_262_v;
  wire signed [`W-1:0] n_260_port_3, n_260_port_4, n_260_v;
  wire signed [`W-1:0] n_261_port_3, n_261_port_4, n_261_v;
  wire signed [`W-1:0] n_269_port_3, n_269_port_4, n_269_v;
  wire signed [`W-1:0] dpc32_PCHADH_port_0, dpc32_PCHADH_port_1, dpc32_PCHADH_v;
  wire signed [`W-1:0] idb1_port_8, idb1_port_9, idb1_port_3, idb1_port_0, idb1_port_7, idb1_port_4, idb1_port_5, idb1_port_10, idb1_v;
  wire signed [`W-1:0] idb0_port_8, idb0_port_2, idb0_port_1, idb0_port_6, idb0_port_7, idb0_port_4, idb0_port_5, idb0_port_10, idb0_v;
  wire signed [`W-1:0] idb3_port_8, idb3_port_9, idb3_port_3, idb3_port_0, idb3_port_1, idb3_port_6, idb3_port_5, idb3_port_10, idb3_v;
  wire signed [`W-1:0] idb2_port_9, idb2_port_3, idb2_port_0, idb2_port_1, idb2_port_6, idb2_port_4, idb2_port_5, idb2_port_10, idb2_v;
  wire signed [`W-1:0] idb5_port_8, idb5_port_9, idb5_port_2, idb5_port_6, idb5_port_7, idb5_port_4, idb5_port_5, idb5_v;
  wire signed [`W-1:0] idb4_port_8, idb4_port_9, idb4_port_0, idb4_port_6, idb4_port_7, idb4_port_4, idb4_port_5, idb4_port_10, idb4_v;
  wire signed [`W-1:0] idb7_port_8, idb7_port_9, idb7_port_2, idb7_port_3, idb7_port_0, idb7_port_7, idb7_port_4, idb7_port_10, idb7_v;
  wire signed [`W-1:0] idb6_port_9, idb6_port_3, idb6_port_0, idb6_port_6, idb6_port_7, idb6_port_5, idb6_port_10, idb6_port_11, idb6_v;
  wire signed [`W-1:0] n_8_port_1, n_8_port_4, n_8_v;
  wire signed [`W-1:0] op_T3_mem_abs_port_7, op_T3_mem_abs_port_5, op_T3_mem_abs_v;
  wire signed [`W-1:0] op_T2_ADL_ADD_port_3, op_T2_ADL_ADD_port_4, op_T2_ADL_ADD_v;
  wire signed [`W-1:0] n_1417_port_2, n_1417_port_0, n_1417_v;
  wire signed [`W-1:0] n_1416_port_2, n_1416_port_0, n_1416_v;
  wire signed [`W-1:0] n_1413_port_2, n_1413_port_1, n_1413_v;
  wire signed [`W-1:0] n_1412_port_2, n_1412_port_0, n_1412_v;
  wire signed [`W-1:0] n_381_port_2, n_381_port_3, n_381_port_1, n_381_v;
  wire signed [`W-1:0] n_383_port_3, n_383_port_0, n_383_v;
  wire signed [`W-1:0] n_385_port_3, n_385_port_4, n_385_v;
  wire signed [`W-1:0] n_384_port_8, n_384_port_6, n_384_v;
  wire signed [`W-1:0] n_386_port_3, n_386_port_0, n_386_v;
  wire signed [`W-1:0] n_389_port_1, n_389_port_4, n_389_v;
  wire signed [`W-1:0] n_388_port_6, n_388_port_5, n_388_v;
  wire signed [`W-1:0] op_T__shift_a_port_9, op_T__shift_a_port_7, op_T__shift_a_v;
  wire signed [`W-1:0] n_927_port_3, n_927_port_1, n_927_v;
  wire signed [`W-1:0] n_920_port_2, n_920_port_1, n_920_v;
  wire signed [`W-1:0] n_923_port_0, n_923_port_4, n_923_v;
  wire signed [`W-1:0] n_928_port_2, n_928_port_3, n_928_port_1, n_928_v;
  wire signed [`W-1:0] n_1039_port_3, n_1039_port_5, n_1039_v;
  wire signed [`W-1:0] alub2_port_0, alub2_port_1, alub2_port_4, alub2_v;
  wire signed [`W-1:0] pch7_port_2, pch7_port_1, pch7_v;
  wire signed [`W-1:0] pch6_port_2, pch6_port_0, pch6_v;
  wire signed [`W-1:0] pch5_port_2, pch5_port_0, pch5_v;
  wire signed [`W-1:0] pch4_port_2, pch4_port_1, pch4_v;
  wire signed [`W-1:0] pch3_port_2, pch3_port_1, pch3_v;
  wire signed [`W-1:0] pch2_port_0, pch2_port_1, pch2_v;
  wire signed [`W-1:0] pch1_port_2, pch1_port_1, pch1_v;
  wire signed [`W-1:0] pch0_port_2, pch0_port_1, pch0_v;
  wire signed [`W-1:0] op_T3_mem_zp_idx_port_7, op_T3_mem_zp_idx_port_5, op_T3_mem_zp_idx_v;
  wire signed [`W-1:0] notalucin_port_2, notalucin_port_4, notalucin_v;
  wire signed [`W-1:0] dpc13_ORS_port_8, dpc13_ORS_port_5, dpc13_ORS_v;
  wire signed [`W-1:0] n_1069_port_3, n_1069_port_4, n_1069_v;
  wire signed [`W-1:0] n_1067_port_2, n_1067_port_0, n_1067_v;
  wire signed [`W-1:0] n_1065_port_2, n_1065_port_1, n_1065_v;
  wire signed [`W-1:0] n_1063_port_2, n_1063_port_7, n_1063_port_4, n_1063_port_5, n_1063_v;
  wire signed [`W-1:0] op_T0_tay_port_9, op_T0_tay_port_11, op_T0_tay_v;
  wire signed [`W-1:0] op_T0_tax_port_9, op_T0_tax_port_10, op_T0_tax_v;
  wire signed [`W-1:0] n_1608_port_2, n_1608_port_1, n_1608_v;
  wire signed [`W-1:0] n_1609_port_3, n_1609_port_0, n_1609_v;
  wire signed [`W-1:0] n_1605_port_3, n_1605_port_0, n_1605_port_5, n_1605_v;
  wire signed [`W-1:0] op_T0_brk_rti_port_8, op_T0_brk_rti_port_9, op_T0_brk_rti_v;
  wire signed [`W-1:0] n_249_port_3, n_249_port_0, n_249_v;
  wire signed [`W-1:0] n_718_port_2, n_718_port_1, n_718_v;
  wire signed [`W-1:0] n_719_port_2, n_719_port_3, n_719_port_0, n_719_port_1, n_719_v;
  wire signed [`W-1:0] n_717_port_4, n_717_port_5, n_717_v;
  wire signed [`W-1:0] n_715_port_2, n_715_port_3, n_715_v;
  wire signed [`W-1:0] n_241_port_2, n_241_port_3, n_241_v;
  wire signed [`W-1:0] n_242_port_2, n_242_port_3, n_242_port_0, n_242_port_1, n_242_v;
  wire signed [`W-1:0] n_243_port_2, n_243_port_1, n_243_v;
  wire signed [`W-1:0] dasb7_port_3, dasb7_port_1, dasb7_port_5, dasb7_v;
  wire signed [`W-1:0] op_T5_rti_rts_port_8, op_T5_rti_rts_port_10, op_T5_rti_rts_v;
  wire signed [`W-1:0] n_669_port_3, n_669_port_4, n_669_v;
  wire signed [`W-1:0] _C23_port_2, _C23_port_3, _C23_v;
  wire signed [`W-1:0] nnT2BR_port_5, nnT2BR_port_10, nnT2BR_v;
  wire signed [`W-1:0] n_1474_port_2, n_1474_port_0, n_1474_v;
  wire signed [`W-1:0] op_T4_ind_x_port_9, op_T4_ind_x_port_7, op_T4_ind_x_v;
  wire signed [`W-1:0] op_T4_ind_y_port_8, op_T4_ind_y_port_6, op_T4_ind_y_v;
  wire signed [`W-1:0] n_1295_port_2, n_1295_port_3, n_1295_v;
  wire signed [`W-1:0] n_1296_port_2, n_1296_port_0, n_1296_v;
  wire signed [`W-1:0] n_1290_port_3, n_1290_port_5, n_1290_v;
  wire signed [`W-1:0] n_1293_port_6, n_1293_port_4, n_1293_v;
  wire signed [`W-1:0] dpc7_SS_port_7, dpc7_SS_port_12, dpc7_SS_v;
  wire signed [`W-1:0] op_T__iny_dey_port_8, op_T__iny_dey_port_9, op_T__iny_dey_v;
  wire signed [`W-1:0] n_906_port_3, n_906_port_0, n_906_v;
  wire signed [`W-1:0] n_905_port_2, n_905_port_3, n_905_v;
  wire signed [`W-1:0] n_1356_port_2, n_1356_port_0, n_1356_v;
  wire signed [`W-1:0] n_1423_port_3, n_1423_port_0, n_1423_v;
  wire signed [`W-1:0] n_38_port_2, n_38_port_1, n_38_v;
  wire signed [`W-1:0] n_1599_port_2, n_1599_port_3, n_1599_v;
  wire signed [`W-1:0] n_1041_port_0, n_1041_port_1, n_1041_v;
  wire signed [`W-1:0] n_1043_port_2, n_1043_port_0, n_1043_v;
  wire signed [`W-1:0] n_1596_port_3, n_1596_port_0, n_1596_v;
  wire signed [`W-1:0] n_1045_port_3, n_1045_port_4, n_1045_v;
  wire signed [`W-1:0] n_1046_port_2, n_1046_port_3, n_1046_port_0, n_1046_v;
  wire signed [`W-1:0] n_1595_port_2, n_1595_port_1, n_1595_v;
  wire signed [`W-1:0] n_1620_port_3, n_1620_port_0, n_1620_v;
  wire signed [`W-1:0] n_1621_port_2, n_1621_port_0, n_1621_port_1, n_1621_v;
  wire signed [`W-1:0] n_1629_port_3, n_1629_port_4, n_1629_v;
  wire signed [`W-1:0] n_228_port_2, n_228_port_0, n_228_v;
  wire signed [`W-1:0] n_220_port_3, n_220_port_0, n_220_v;
  wire signed [`W-1:0] n_221_port_2, n_221_port_1, n_221_v;
  wire signed [`W-1:0] n_227_port_2, n_227_port_3, n_227_port_0, n_227_v;
  wire signed [`W-1:0] n_224_port_4, n_224_port_5, n_224_v;
  wire signed [`W-1:0] n_225_port_2, n_225_port_0, n_225_v;
  wire signed [`W-1:0] op_T4_abs_idx_port_6, op_T4_abs_idx_port_4, op_T4_abs_idx_v;
  wire signed [`W-1:0] op_implied_port_6, op_implied_port_5, op_implied_v;
  wire signed [`W-1:0] n_735_port_3, n_735_port_4, n_735_v;
  wire signed [`W-1:0] n_730_port_2, n_730_port_1, n_730_v;
  wire signed [`W-1:0] n_732_port_8, n_732_port_4, n_732_v;
  wire signed [`W-1:0] dpc22__DSA_port_3, dpc22__DSA_port_0, dpc22__DSA_v;
  wire signed [`W-1:0] n_739_port_9, n_739_port_4, n_739_v;
  wire signed [`W-1:0] x2_port_0, x2_port_1, x2_v;
  wire signed [`W-1:0] x3_port_0, x3_port_1, x3_v;
  wire signed [`W-1:0] x0_port_0, x0_port_1, x0_v;
  wire signed [`W-1:0] x1_port_0, x1_port_1, x1_v;
  wire signed [`W-1:0] op_T__dex_port_9, op_T__dex_port_10, op_T__dex_v;
  wire signed [`W-1:0] x7_port_2, x7_port_1, x7_v;
  wire signed [`W-1:0] x4_port_0, x4_port_1, x4_v;
  wire signed [`W-1:0] x5_port_2, x5_port_1, x5_v;
  wire signed [`W-1:0] _C01_port_2, _C01_port_3, _C01_v;
  wire signed [`W-1:0] op_T0_sbc_port_8, op_T0_sbc_port_9, op_T0_sbc_v;
  wire signed [`W-1:0] n_410_port_6, n_410_port_5, n_410_v;
  wire signed [`W-1:0] n_1458_port_2, n_1458_port_3, n_1458_port_0, n_1458_port_1, n_1458_port_4, n_1458_v;
  wire signed [`W-1:0] n_1457_port_3, n_1457_port_4, n_1457_v;
  wire signed [`W-1:0] n_1455_port_9, n_1455_port_10, n_1455_v;
  wire signed [`W-1:0] DA_AB2_port_2, DA_AB2_port_3, DA_AB2_v;
  wire signed [`W-1:0] n_692_port_4, n_692_port_5, n_692_v;
  wire signed [`W-1:0] n_695_port_2, n_695_port_3, n_695_v;
  wire signed [`W-1:0] n_694_port_2, n_694_port_3, n_694_port_0, n_694_port_1, n_694_port_4, n_694_v;
  wire signed [`W-1:0] n_969_port_2, n_969_port_0, n_969_v;
  wire signed [`W-1:0] n_961_port_2, n_961_port_0, n_961_v;
  wire signed [`W-1:0] n_963_port_2, n_963_port_1, n_963_v;
  wire signed [`W-1:0] n_962_port_2, n_962_port_1, n_962_v;
  wire signed [`W-1:0] n_964_port_7, n_964_port_4, n_964_v;
  wire signed [`W-1:0] n_966_port_3, n_966_port_0, n_966_v;
  wire signed [`W-1:0] irline3_port_0, irline3_port_64, irline3_v;
  wire signed [`W-1:0] pcl3_port_2, pcl3_port_1, pcl3_v;
  wire signed [`W-1:0] pcl2_port_2, pcl2_port_1, pcl2_v;
  wire signed [`W-1:0] pcl1_port_2, pcl1_port_1, pcl1_v;
  wire signed [`W-1:0] pcl0_port_2, pcl0_port_1, pcl0_v;
  wire signed [`W-1:0] pcl7_port_2, pcl7_port_1, pcl7_v;
  wire signed [`W-1:0] pcl6_port_2, pcl6_port_1, pcl6_v;
  wire signed [`W-1:0] pcl5_port_2, pcl5_port_1, pcl5_v;
  wire signed [`W-1:0] pcl4_port_2, pcl4_port_1, pcl4_v;
  wire signed [`W-1:0] dpc0_YSB_port_3, dpc0_YSB_port_12, dpc0_YSB_v;
  wire signed [`W-1:0] n_1026_port_3, n_1026_port_0, n_1026_v;
  wire signed [`W-1:0] n_1024_port_3, n_1024_port_0, n_1024_v;
  wire signed [`W-1:0] n_1025_port_2, n_1025_port_1, n_1025_v;
  wire signed [`W-1:0] alua6_port_0, alua6_port_1, alua6_v;
  wire signed [`W-1:0] alua7_port_3, alua7_port_0, alua7_v;
  wire signed [`W-1:0] alua4_port_0, alua4_port_1, alua4_v;
  wire signed [`W-1:0] alua5_port_0, alua5_port_1, alua5_v;
  wire signed [`W-1:0] alua2_port_0, alua2_port_1, alua2_v;
  wire signed [`W-1:0] alua3_port_0, alua3_port_1, alua3_v;
  wire signed [`W-1:0] alua0_port_0, alua0_port_1, alua0_v;
  wire signed [`W-1:0] alua1_port_2, alua1_port_3, alua1_v;
  wire signed [`W-1:0] n_1271_port_2, n_1271_port_0, n_1271_v;
  wire signed [`W-1:0] nmi_port_2, nmi_v;
  wire signed [`W-1:0] op_T2_branch_port_6, op_T2_branch_port_7, op_T2_branch_v;
  wire signed [`W-1:0] dpc41_DL_ADL_port_9, dpc41_DL_ADL_port_0, dpc41_DL_ADL_v;
  wire signed [`W-1:0] n_200_port_7, n_200_port_5, n_200_v;
  wire signed [`W-1:0] n_753_port_4, n_753_port_5, n_753_v;
  wire signed [`W-1:0] n_757_port_2, n_757_port_5, n_757_v;
  wire signed [`W-1:0] n_754_port_8, n_754_port_4, n_754_v;
  wire signed [`W-1:0] n_207_port_3, n_207_port_5, n_207_v;
  wire signed [`W-1:0] n_208_port_2, n_208_port_3, n_208_port_0, n_208_port_1, n_208_port_4, n_208_v;
  wire signed [`W-1:0] n_209_port_2, n_209_port_3, n_209_port_0, n_209_port_1, n_209_port_4, n_209_v;
  wire signed [`W-1:0] _C67_port_3, _C67_port_0, _C67_v;
  wire signed [`W-1:0] dpc37_PCLDB_port_0, dpc37_PCLDB_port_4, dpc37_PCLDB_v;
  wire signed [`W-1:0] __AxB3__C23_port_3, __AxB3__C23_port_4, __AxB3__C23_v;
  wire signed [`W-1:0] pd5_clearIR_port_3, pd5_clearIR_port_4, pd5_clearIR_v;
  wire signed [`W-1:0] dpc12_0ADD_port_9, dpc12_0ADD_port_12, dpc12_0ADD_v;
  wire signed [`W-1:0] dpc4_SSB_port_9, dpc4_SSB_port_0, dpc4_SSB_v;
  wire signed [`W-1:0] n_134_port_7, n_134_port_5, n_134_v;
  wire signed [`W-1:0] n_947_port_2, n_947_port_1, n_947_v;
  wire signed [`W-1:0] n_946_port_2, n_946_port_4, n_946_v;
  wire signed [`W-1:0] n_417_port_0, n_417_port_1, n_417_v;
  wire signed [`W-1:0] n_944_port_3, n_944_port_4, n_944_v;
  wire signed [`W-1:0] op_T0_cpy_iny_port_9, op_T0_cpy_iny_port_7, op_T0_cpy_iny_v;
  wire signed [`W-1:0] n_419_port_2, n_419_port_0, n_419_v;
  wire signed [`W-1:0] y1_port_2, y1_port_0, y1_v;
  wire signed [`W-1:0] y0_port_2, y0_port_0, y0_v;
  wire signed [`W-1:0] y3_port_2, y3_port_0, y3_v;
  wire signed [`W-1:0] y2_port_2, y2_port_0, y2_v;
  wire signed [`W-1:0] y5_port_0, y5_port_1, y5_v;
  wire signed [`W-1:0] y4_port_2, y4_port_0, y4_v;
  wire signed [`W-1:0] y7_port_0, y7_port_1, y7_v;
  wire signed [`W-1:0] y6_port_0, y6_port_1, y6_v;
  wire signed [`W-1:0] n_1007_port_2, n_1007_port_1, n_1007_v;
  wire signed [`W-1:0] n_1002_port_1, n_1002_port_5, n_1002_v;
  wire signed [`W-1:0] abh5_port_3, abh5_port_4, abh5_v;
  wire signed [`W-1:0] abh4_port_0, abh4_port_4, abh4_v;
  wire signed [`W-1:0] abh7_port_0, abh7_port_4, abh7_v;
  wire signed [`W-1:0] abh6_port_3, abh6_port_4, abh6_v;
  wire signed [`W-1:0] abh1_port_3, abh1_port_4, abh1_v;
  wire signed [`W-1:0] abh0_port_3, abh0_port_4, abh0_v;
  wire signed [`W-1:0] abh3_port_3, abh3_port_4, abh3_v;
  wire signed [`W-1:0] abh2_port_0, abh2_port_4, abh2_v;
  wire signed [`W-1:0] n_1552_port_2, n_1552_port_0, n_1552_v;
  wire signed [`W-1:0] alucin_port_2, alucin_port_1, alucin_v;
  wire signed [`W-1:0] x_op_push_pull_port_8, x_op_push_pull_port_6, x_op_push_pull_v;
  wire signed [`W-1:0] dpc11_SBADD_port_9, dpc11_SBADD_port_12, dpc11_SBADD_v;
  wire signed [`W-1:0] dpc10_ADLADD_port_5, dpc10_ADLADD_port_12, dpc10_ADLADD_v;
  wire signed [`W-1:0] n_779_port_3, n_779_port_5, n_779_v;
  wire signed [`W-1:0] n_770_port_3, n_770_port_1, n_770_v;
  wire signed [`W-1:0] n_771_port_1, n_771_port_4, n_771_v;
  wire signed [`W-1:0] n_772_port_2, n_772_port_3, n_772_v;
  wire signed [`W-1:0] n_773_port_3, n_773_port_5, n_773_v;
  wire signed [`W-1:0] n_774_port_2, n_774_port_0, n_774_v;
  wire signed [`W-1:0] n_837_port_2, n_837_port_0, n_837_v;
  wire signed [`W-1:0] op_T0_bit_port_8, op_T0_bit_port_10, op_T0_bit_v;
  wire signed [`W-1:0] n_344_port_8, n_344_port_4, n_344_v;
  wire signed [`W-1:0] n_834_port_2, n_834_port_4, n_834_v;
  wire signed [`W-1:0] dpc29_0ADH17_port_2, dpc29_0ADH17_port_1, dpc29_0ADH17_v;
  wire signed [`W-1:0] dpc26_ACDB_port_0, dpc26_ACDB_port_12, dpc26_ACDB_v;
  wire signed [`W-1:0] _C45_port_1, _C45_port_4, _C45_v;
  wire signed [`W-1:0] VEC0_port_6, VEC0_port_5, VEC0_v;
  wire signed [`W-1:0] VEC1_port_3, VEC1_port_4, VEC1_v;
  wire signed [`W-1:0] op_T4_rts_port_9, op_T4_rts_port_11, op_T4_rts_v;
  wire signed [`W-1:0] n_430_port_2, n_430_port_3, n_430_port_1, n_430_v;
  wire signed [`W-1:0] n_436_port_2, n_436_port_3, n_436_port_0, n_436_port_1, n_436_v;
  wire signed [`W-1:0] op_T4_rti_port_9, op_T4_rti_port_10, op_T4_rti_v;
  wire signed [`W-1:0] op_SRS_port_2, op_SRS_port_6, op_SRS_v;
  wire signed [`W-1:0] n_1343_port_3, n_1343_port_5, n_1343_v;
  wire signed [`W-1:0] n_1345_port_7, n_1345_port_5, n_1345_v;
  wire signed [`W-1:0] n_1578_port_2, n_1578_port_1, n_1578_v;
  wire signed [`W-1:0] n_1573_port_2, n_1573_port_0, n_1573_v;
  wire signed [`W-1:0] DC78_port_7, DC78_port_4, DC78_v;
  wire signed [`W-1:0] op_sta_cmp_port_6, op_sta_cmp_port_5, op_sta_cmp_v;
  wire signed [`W-1:0] op_SUMS_port_6, op_SUMS_port_5, op_SUMS_v;
  wire signed [`W-1:0] n_1688_port_2, n_1688_port_0, n_1688_v;
  wire signed [`W-1:0] n_404_port_2, n_404_port_6, n_404_port_5, n_404_v;
  wire signed [`W-1:0] n_954_port_3, n_954_port_4, n_954_v;
  wire signed [`W-1:0] n_400_port_2, n_400_port_3, n_400_v;
  wire signed [`W-1:0] op_T4_brk_jsr_port_8, op_T4_brk_jsr_port_9, op_T4_brk_jsr_v;
  wire signed [`W-1:0] n_1219_port_2, n_1219_port_1, n_1219_v;
  wire signed [`W-1:0] n_1215_port_6, n_1215_port_5, n_1215_v;
  wire signed [`W-1:0] n_1214_port_2, n_1214_port_0, n_1214_v;
  wire signed [`W-1:0] n_1211_port_8, n_1211_port_9, n_1211_v;
  wire signed [`W-1:0] n_1213_port_3, n_1213_port_4, n_1213_v;
  wire signed [`W-1:0] n_1655_port_2, n_1655_port_1, n_1655_v;
  wire signed [`W-1:0] pd2_clearIR_port_6, pd2_clearIR_port_7, pd2_clearIR_v;
  wire signed [`W-1:0] n_1654_port_2, n_1654_port_3, n_1654_port_0, n_1654_port_1, n_1654_port_4, n_1654_v;
  wire signed [`W-1:0] n_1657_port_2, n_1657_port_3, n_1657_v;
  wire signed [`W-1:0] n_1650_port_2, n_1650_port_0, n_1650_v;
  wire signed [`W-1:0] n_182_port_7, n_182_port_11, n_182_v;
  wire signed [`W-1:0] n_180_port_3, n_180_port_5, n_180_v;
  wire signed [`W-1:0] n_184_port_2, n_184_port_0, n_184_v;
  wire signed [`W-1:0] n_635_port_3, n_635_port_0, n_635_port_1, n_635_v;
  wire signed [`W-1:0] n_634_port_0, n_634_port_1, n_634_v;
  wire signed [`W-1:0] n_637_port_3, n_637_port_4, n_637_v;
  wire signed [`W-1:0] n_636_port_2, n_636_port_0, n_636_v;
  wire signed [`W-1:0] n_631_port_2, n_631_port_3, n_631_v;
  wire signed [`W-1:0] n_630_port_3, n_630_port_0, n_630_v;
  wire signed [`W-1:0] n_633_port_0, n_633_v;
  wire signed [`W-1:0] n_632_port_3, n_632_port_5, n_632_v;
  wire signed [`W-1:0] n_458_port_2, n_458_port_0, n_458_port_1, n_458_v;
  wire signed [`W-1:0] n_988_port_3, n_988_port_1, n_988_v;
  wire signed [`W-1:0] n_983_port_2, n_983_port_1, n_983_v;
  wire signed [`W-1:0] n_981_port_2, n_981_port_1, n_981_v;
  wire signed [`W-1:0] n_987_port_2, n_987_port_1, n_987_v;
  wire signed [`W-1:0] n_986_port_2, n_986_port_3, n_986_v;
  wire signed [`W-1:0] n_457_port_2, n_457_port_1, n_457_v;
  wire signed [`W-1:0] op_T0_lda_port_9, op_T0_lda_port_7, op_T0_lda_v;
  wire signed [`W-1:0] abl1_port_3, abl1_port_4, abl1_v;
  wire signed [`W-1:0] abl0_port_3, abl0_port_4, abl0_v;
  wire signed [`W-1:0] abl4_port_0, abl4_port_4, abl4_v;
  wire signed [`W-1:0] op_T3_plp_pla_port_8, op_T3_plp_pla_port_10, op_T3_plp_pla_v;
  wire signed [`W-1:0] n_1517_port_3, n_1517_port_4, n_1517_v;
  wire signed [`W-1:0] n_1518_port_2, n_1518_port_1, n_1518_v;
  wire signed [`W-1:0] n_1519_port_2, n_1519_port_3, n_1519_port_0, n_1519_v;
  wire signed [`W-1:0] n_279_port_4, n_279_port_5, n_279_v;
  wire signed [`W-1:0] n_846_port_3, n_846_port_1, n_846_v;
  wire signed [`W-1:0] n_847_port_2, n_847_port_1, n_847_v;
  wire signed [`W-1:0] n_844_port_6, n_844_port_5, n_844_v;
  wire signed [`W-1:0] n_845_port_8, n_845_port_4, n_845_v;
  wire signed [`W-1:0] n_842_port_3, n_842_port_0, n_842_v;
  wire signed [`W-1:0] op_T3_jmp_port_8, op_T3_jmp_port_9, op_T3_jmp_v;
  wire signed [`W-1:0] n_849_port_2, n_849_port_0, n_849_v;
  wire signed [`W-1:0] __AxB5__C45_port_3, __AxB5__C45_port_4, __AxB5__C45_v;
  wire signed [`W-1:0] dpc16_EORS_port_8, dpc16_EORS_port_9, dpc16_EORS_v;
  wire signed [`W-1:0] n_1231_port_2, n_1231_port_1, n_1231_v;
  wire signed [`W-1:0] n_1230_port_4, n_1230_port_5, n_1230_v;
  wire signed [`W-1:0] n_1238_port_2, n_1238_port_1, n_1238_v;
  wire signed [`W-1:0] n_1722_port_2, n_1722_port_3, n_1722_port_0, n_1722_port_1, n_1722_port_4, n_1722_v;
  wire signed [`W-1:0] op_branch_done_port_8, op_branch_done_port_9, op_branch_done_v;
  wire signed [`W-1:0] aluvout_port_2, aluvout_port_0, aluvout_v;
  wire signed [`W-1:0] n_618_port_2, n_618_port_3, n_618_port_0, n_618_port_1, n_618_port_4, n_618_v;
  wire signed [`W-1:0] n_613_port_4, n_613_port_10, n_613_v;
  wire signed [`W-1:0] n_612_port_0, n_612_port_4, n_612_v;
  wire signed [`W-1:0] n_611_port_4, n_611_port_5, n_611_v;
  wire signed [`W-1:0] n_617_port_3, n_617_port_0, n_617_v;
  wire signed [`W-1:0] n_616_port_6, n_616_port_5, n_616_v;
  wire signed [`W-1:0] n_1137_port_2, n_1137_port_4, n_1137_v;
  wire signed [`W-1:0] n_620_port_6, n_620_port_7, n_620_v;
  wire signed [`W-1:0] n_884_port_2, n_884_port_0, n_884_port_1, n_884_v;
  wire signed [`W-1:0] Pout0_port_2, Pout0_port_0, Pout0_port_1, Pout0_v;
  wire signed [`W-1:0] n_1545_port_2, n_1545_port_1, n_1545_v;
  wire signed [`W-1:0] n_1010_port_3, n_1010_port_0, n_1010_v;
  wire signed [`W-1:0] n_1017_port_2, n_1017_port_0, n_1017_v;
  wire signed [`W-1:0] n_1542_port_6, n_1542_port_4, n_1542_v;
  wire signed [`W-1:0] dpc19_ADDSB7_port_2, dpc19_ADDSB7_port_0, dpc19_ADDSB7_v;
  wire signed [`W-1:0] n_477_port_3, n_477_port_1, n_477_port_4, n_477_port_5, n_477_v;
  wire signed [`W-1:0] n_476_port_4, n_476_port_5, n_476_v;
  wire signed [`W-1:0] n_475_port_2, n_475_port_0, n_475_v;
  wire signed [`W-1:0] n_474_port_3, n_474_port_5, n_474_v;
  wire signed [`W-1:0] n_473_port_2, n_473_port_3, n_473_v;
  wire signed [`W-1:0] n_472_port_3, n_472_port_6, n_472_v;
  wire signed [`W-1:0] n_471_port_3, n_471_port_4, n_471_v;
  wire signed [`W-1:0] n_470_port_2, n_470_port_3, n_470_v;
  wire signed [`W-1:0] n_479_port_3, n_479_port_4, n_479_v;
  wire signed [`W-1:0] n_478_port_2, n_478_port_0, n_478_port_1, n_478_v;
  wire signed [`W-1:0] brk_done_port_9, brk_done_port_12, brk_done_v;
  wire signed [`W-1:0] op_T0_txa_port_9, op_T0_txa_port_11, op_T0_txa_v;
  wire signed [`W-1:0] p6_port_2, p6_port_0, p6_port_1, p6_v;
  wire signed [`W-1:0] p7_port_2, p7_port_0, p7_port_1, p7_v;
  wire signed [`W-1:0] DC34_port_9, DC34_port_4, DC34_v;
  wire signed [`W-1:0] op_T2_stack_port_8, op_T2_stack_port_7, op_T2_stack_v;
  wire signed [`W-1:0] n_1534_port_4, n_1534_port_5, n_1534_v;
  wire signed [`W-1:0] n_1531_port_2, n_1531_port_3, n_1531_port_0, n_1531_port_1, n_1531_v;
  wire signed [`W-1:0] n_1391_port_3, n_1391_port_4, n_1391_v;
  wire signed [`W-1:0] n_1392_port_2, n_1392_port_3, n_1392_v;
  wire signed [`W-1:0] n_1398_port_8, n_1398_port_1, n_1398_port_6, n_1398_v;
  wire signed [`W-1:0] n_1399_port_3, n_1399_port_0, n_1399_v;
  wire signed [`W-1:0] n_288_port_6, n_288_port_4, n_288_v;
  wire signed [`W-1:0] n_280_port_2, n_280_port_3, n_280_port_0, n_280_port_1, n_280_port_4, n_280_v;
  wire signed [`W-1:0] n_282_port_2, n_282_port_1, n_282_v;
  wire signed [`W-1:0] n_284_port_2, n_284_port_0, n_284_v;
  wire signed [`W-1:0] n_135_port_2, n_135_port_1, n_135_v;
  wire signed [`W-1:0] n_133_port_4, n_133_port_5, n_133_v;
  wire signed [`W-1:0] n_130_port_2, n_130_port_0, n_130_v;
  wire signed [`W-1:0] n_869_port_2, n_869_port_3, n_869_port_1, n_869_v;
  wire signed [`W-1:0] n_866_v;
  wire signed [`W-1:0] n_867_port_3, n_867_port_4, n_867_v;
  wire signed [`W-1:0] n_861_port_2, n_861_port_0, n_861_v;
  wire signed [`W-1:0] n_862_port_9, n_862_port_4, n_862_v;
  wire signed [`W-1:0] n_350_port_3, n_350_port_1, n_350_port_4, n_350_port_5, n_350_v;
  wire signed [`W-1:0] dpc17_SUMS_port_0, dpc17_SUMS_port_1, dpc17_SUMS_v;
  wire signed [`W-1:0] _op_branch_done_port_2, _op_branch_done_port_0, _op_branch_done_v;
  wire signed [`W-1:0] op_T0_acc_port_3, op_T0_acc_port_4, op_T0_acc_v;
  wire signed [`W-1:0] BRtaken_port_4, BRtaken_port_10, BRtaken_v;
  wire signed [`W-1:0] n_1251_port_2, n_1251_port_3, n_1251_port_0, n_1251_port_1, n_1251_v;
  wire signed [`W-1:0] n_1253_port_7, n_1253_port_5, n_1253_v;
  wire signed [`W-1:0] n_1257_port_7, n_1257_port_5, n_1257_v;
  wire signed [`W-1:0] n_1258_port_7, n_1258_port_4, n_1258_v;
  wire signed [`W-1:0] n_1709_port_2, n_1709_port_3, n_1709_port_0, n_1709_port_1, n_1709_v;
  wire signed [`W-1:0] n_1708_port_3, n_1708_port_4, n_1708_v;
  wire signed [`W-1:0] dpc3_SBX_port_9, dpc3_SBX_port_12, dpc3_SBX_v;
  wire signed [`W-1:0] op_T2_php_port_9, op_T2_php_port_10, op_T2_php_v;
  wire signed [`W-1:0] op_T2_pha_port_9, op_T2_pha_port_10, op_T2_pha_v;
  wire signed [`W-1:0] dpc31_PCHPCH_port_11, dpc31_PCHPCH_port_12, dpc31_PCHPCH_v;
  wire signed [`W-1:0] n_670_port_2, n_670_port_3, n_670_v;
  wire signed [`W-1:0] n_673_port_2, n_673_port_4, n_673_v;
  wire signed [`W-1:0] n_674_port_2, n_674_port_0, n_674_v;
  wire signed [`W-1:0] n_676_port_2, n_676_port_3, n_676_port_0, n_676_v;
  wire signed [`W-1:0] n_678_port_4, n_678_port_5, n_678_v;
  wire signed [`W-1:0] Pout1_port_2, Pout1_port_0, Pout1_port_1, Pout1_v;
  wire signed [`W-1:0] Pout3_port_2, Pout3_port_3, Pout3_port_4, Pout3_v;
  wire signed [`W-1:0] Pout2_port_2, Pout2_port_0, Pout2_port_1, Pout2_v;
  wire signed [`W-1:0] n_499_port_3, n_499_port_0, n_499_v;
  wire signed [`W-1:0] n_494_port_2, n_494_port_3, n_494_port_1, n_494_v;
  wire signed [`W-1:0] n_496_port_2, n_496_port_1, n_496_v;
  wire signed [`W-1:0] n_491_port_2, n_491_port_1, n_491_v;
  wire signed [`W-1:0] n_490_port_2, n_490_port_1, n_490_v;
  wire signed [`W-1:0] pd7_clearIR_port_4, pd7_clearIR_port_5, pd7_clearIR_v;
  wire signed [`W-1:0] n_1401_port_2, n_1401_port_0, n_1401_v;
  wire signed [`W-1:0] op_T4_jmp_port_9, op_T4_jmp_port_11, op_T4_jmp_v;
  wire signed [`W-1:0] n_19_port_3, n_19_port_4, n_19_v;
  wire signed [`W-1:0] n_1117_port_2, n_1117_port_1, n_1117_v;
  wire signed [`W-1:0] n_1115_port_3, n_1115_port_4, n_1115_v;
  wire signed [`W-1:0] n_1110_port_3, n_1110_port_1, n_1110_v;
  wire signed [`W-1:0] n_1111_port_3, n_1111_port_6, n_1111_v;
  wire signed [`W-1:0] n_803_port_2, n_803_port_0, n_803_v;
  wire signed [`W-1:0] n_800_port_2, n_800_port_0, n_800_v;
  wire signed [`W-1:0] n_806_v;
  wire signed [`W-1:0] n_807_port_3, n_807_port_5, n_807_v;
  wire signed [`W-1:0] n_432_port_2, n_432_port_3, n_432_v;
  wire signed [`W-1:0] n_1277_port_3, n_1277_port_0, n_1277_v;
  wire signed [`W-1:0] n_1275_port_4, n_1275_port_5, n_1275_v;
  wire signed [`W-1:0] n_1660_port_3, n_1660_port_0, n_1660_v;
  wire signed [`W-1:0] op_inc_nop_port_6, op_inc_nop_port_5, op_inc_nop_v;
  wire signed [`W-1:0] n_128_port_2, n_128_port_0, n_128_v;
  wire signed [`W-1:0] n_659_port_2, n_659_port_3, n_659_port_1, n_659_v;
  wire signed [`W-1:0] n_658_port_2, n_658_port_3, n_658_port_0, n_658_port_1, n_658_v;
  wire signed [`W-1:0] n_127_port_4, n_127_port_5, n_127_v;
  wire signed [`W-1:0] n_652_port_2, n_652_port_3, n_652_port_0, n_652_port_1, n_652_port_4, n_652_v;
  wire signed [`W-1:0] n_123_port_2, n_123_port_3, n_123_port_0, n_123_v;
  wire signed [`W-1:0] n_122_port_2, n_122_port_0, n_122_v;
  wire signed [`W-1:0] op_T0_shift_right_a_port_8, op_T0_shift_right_a_port_9, op_T0_shift_right_a_v;
  wire signed [`W-1:0] op_T0_adc_sbc_port_8, op_T0_adc_sbc_port_6, op_T0_adc_sbc_v;
  wire signed [`W-1:0] op_push_pull_port_8, op_push_pull_port_7, op_push_pull_v;
  wire signed [`W-1:0] n_1130_port_8, n_1130_port_7, n_1130_v;
  wire signed [`W-1:0] n_1133_port_3, n_1133_port_4, n_1133_v;
  wire signed [`W-1:0] n_1135_port_2, n_1135_port_3, n_1135_v;
  wire signed [`W-1:0] n_1138_port_2, n_1138_port_0, n_1138_v;
  wire signed [`W-1:0] op_T2_mem_zp_port_7, op_T2_mem_zp_port_5, op_T2_mem_zp_v;
  wire signed [`W-1:0] n_355_port_3, n_355_port_0, n_355_v;
  wire signed [`W-1:0] n_824_port_6, n_824_port_5, n_824_v;
  wire signed [`W-1:0] n_826_port_2, n_826_port_1, n_826_v;
  wire signed [`W-1:0] n_351_port_2, n_351_port_0, n_351_port_1, n_351_v;
  wire signed [`W-1:0] dpc9_DBADD_port_1, dpc9_DBADD_port_12, dpc9_DBADD_v;
  wire signed [`W-1:0] n_358_port_2, n_358_port_4, n_358_v;
  wire signed [`W-1:0] n_359_port_2, n_359_port_0, n_359_port_1, n_359_v;
  wire signed [`W-1:0] dpc33_PCHDB_port_0, dpc33_PCHDB_port_1, dpc33_PCHDB_v;
  wire signed [`W-1:0] INTG_port_6, INTG_port_4, INTG_v;
  wire signed [`W-1:0] n_755_port_3, n_755_port_0, n_755_v;
  wire signed [`W-1:0] op_T2_ind_port_6, op_T2_ind_port_5, op_T2_ind_v;
  wire signed [`W-1:0] op_rti_rts_port_9, op_rti_rts_port_10, op_rti_rts_v;
  wire signed [`W-1:0] dpc8_nDBADD_port_6, dpc8_nDBADD_port_12, dpc8_nDBADD_v;
  wire signed [`W-1:0] n_109_port_2, n_109_port_0, n_109_v;
  wire signed [`W-1:0] n_108_port_2, n_108_port_1, n_108_v;
  wire signed [`W-1:0] n_102_port_2, n_102_port_0, n_102_v;
  wire signed [`W-1:0] n_105_port_2, n_105_port_3, n_105_v;
  wire signed [`W-1:0] n_104_port_6, n_104_port_7, n_104_v;
  wire signed [`W-1:0] n_1575_port_4, n_1575_port_5, n_1575_v;
  wire signed [`W-1:0] dpc39_PCLPCL_port_11, dpc39_PCLPCL_port_12, dpc39_PCLPCL_v;
  wire signed [`W-1:0] ADH_ABH_port_7, ADH_ABH_port_4, ADH_ABH_v;
  wire signed [`W-1:0] Reset0_port_4, Reset0_port_5, Reset0_v;
  wire signed [`W-1:0] dpc25_SBDB_port_9, dpc25_SBDB_port_0, dpc25_SBDB_v;
  wire signed [`W-1:0] n_1541_port_4, n_1541_port_5, n_1541_v;
  wire signed [`W-1:0] dpc23_SBAC_port_11, dpc23_SBAC_port_12, dpc23_SBAC_v;
  wire signed [`W-1:0] n_1484_port_2, n_1484_port_0, n_1484_v;
  wire signed [`W-1:0] x_op_jmp_port_8, x_op_jmp_port_9, x_op_jmp_v;
  wire signed [`W-1:0] n_1339_port_2, n_1339_port_1, n_1339_v;
  wire signed [`W-1:0] n_1488_port_3, n_1488_port_0, n_1488_v;
  wire signed [`W-1:0] n_1335_port_2, n_1335_port_0, n_1335_v;
  wire signed [`W-1:0] n_1159_port_3, n_1159_port_4, n_1159_v;
  wire signed [`W-1:0] n_1152_port_2, n_1152_port_0, n_1152_v;
  wire signed [`W-1:0] n_1157_port_2, n_1157_port_0, n_1157_v;
  wire signed [`W-1:0] n_1154_port_3, n_1154_port_5, n_1154_v;
  wire signed [`W-1:0] _t2_port_0, _t2_port_21, _t2_v;
  wire signed [`W-1:0] _t3_port_15, _t3_port_16, _t3_v;
  wire signed [`W-1:0] n_595_port_4, n_595_port_5, n_595_v;
  wire signed [`W-1:0] _t4_port_0, _t4_port_13, _t4_v;
  wire signed [`W-1:0] _t5_port_0, _t5_port_10, _t5_v;
  wire signed [`W-1:0] n_1682_port_2, n_1682_port_1, n_1682_v;
  wire signed [`W-1:0] n_378_port_4, n_378_port_5, n_378_v;
  wire signed [`W-1:0] n_374_port_2, n_374_port_1, n_374_v;
  wire signed [`W-1:0] n_372_port_2, n_372_port_0, n_372_v;
  wire signed [`W-1:0] n_373_port_0, n_373_port_4, n_373_v;
  wire signed [`W-1:0] x_op_T0_txa_port_9, x_op_T0_txa_port_11, x_op_T0_txa_v;
  wire signed [`W-1:0] C01_port_8, C01_port_4, C01_v;
  wire signed [`W-1:0] op_store_port_4, op_store_port_5, op_store_v;
  wire signed [`W-1:0] n_1687_port_2, n_1687_port_1, n_1687_v;
  wire signed [`W-1:0] ab0_port_0, ab0_port_1, ab0_v;
  wire signed [`W-1:0] ab1_port_0, ab1_port_1, ab1_v;
  wire signed [`W-1:0] ab2_port_0, ab2_port_1, ab2_v;
  wire signed [`W-1:0] ab3_port_0, ab3_port_1, ab3_v;
  wire signed [`W-1:0] ab4_port_0, ab4_port_1, ab4_v;
  wire signed [`W-1:0] ab5_port_0, ab5_port_1, ab5_v;
  wire signed [`W-1:0] ab6_port_0, ab6_port_1, ab6_v;
  wire signed [`W-1:0] ab7_port_0, ab7_port_1, ab7_v;
  wire signed [`W-1:0] ab8_port_0, ab8_port_1, ab8_v;
  wire signed [`W-1:0] ab9_port_0, ab9_port_1, ab9_v;
  wire signed [`W-1:0] n_80_port_3, n_80_port_4, n_80_v;
  wire signed [`W-1:0] n_83_port_3, n_83_port_0, n_83_v;
  wire signed [`W-1:0] n_87_port_2, n_87_port_3, n_87_port_0, n_87_port_1, n_87_v;
  wire signed [`W-1:0] n_86_port_2, n_86_port_3, n_86_port_0, n_86_v;
  wire signed [`W-1:0] n_1684_port_2, n_1684_port_1, n_1684_v;
  wire signed [`W-1:0] n_161_port_4, n_161_port_5, n_161_v;
  wire signed [`W-1:0] n_160_port_3, n_160_port_4, n_160_v;
  wire signed [`W-1:0] n_163_port_2, n_163_port_3, n_163_v;
  wire signed [`W-1:0] n_169_port_3, n_169_port_4, n_169_v;
  wire signed [`W-1:0] n_168_port_2, n_168_port_3, n_168_port_0, n_168_v;
  wire signed [`W-1:0] n_781_port_9, n_781_port_13, n_781_v;
  wire signed [`W-1:0] n_783_port_3, n_783_port_4, n_783_v;
  wire signed [`W-1:0] n_782_port_2, n_782_port_4, n_782_v;
  wire signed [`W-1:0] n_789_port_2, n_789_port_0, n_789_v;
  wire signed [`W-1:0] sb2_port_8, sb2_port_9, sb2_port_2, sb2_port_3, sb2_port_0, sb2_port_1, sb2_port_6, sb2_port_7, sb2_port_4, sb2_port_10, sb2_port_11, sb2_port_12, sb2_v;
  wire signed [`W-1:0] sb3_port_8, sb3_port_9, sb3_port_2, sb3_port_3, sb3_port_0, sb3_port_1, sb3_port_6, sb3_port_7, sb3_port_4, sb3_port_5, sb3_port_10, sb3_port_11, sb3_v;
  wire signed [`W-1:0] sb0_port_8, sb0_port_9, sb0_port_2, sb0_port_3, sb0_port_0, sb0_port_1, sb0_port_6, sb0_port_7, sb0_port_4, sb0_port_5, sb0_port_10, sb0_port_11, sb0_port_12, sb0_v;
  wire signed [`W-1:0] sb1_port_8, sb1_port_9, sb1_port_2, sb1_port_0, sb1_port_1, sb1_port_6, sb1_port_7, sb1_port_4, sb1_port_5, sb1_port_10, sb1_port_11, sb1_port_12, sb1_v;
  wire signed [`W-1:0] sb6_port_8, sb6_port_9, sb6_port_2, sb6_port_3, sb6_port_0, sb6_port_1, sb6_port_6, sb6_port_7, sb6_port_4, sb6_port_10, sb6_port_11, sb6_port_12, sb6_v;
  wire signed [`W-1:0] sb7_port_8, sb7_port_9, sb7_port_2, sb7_port_3, sb7_port_0, sb7_port_1, sb7_port_6, sb7_port_7, sb7_port_4, sb7_port_5, sb7_port_10, sb7_port_11, sb7_v;
  wire signed [`W-1:0] sb4_port_8, sb4_port_9, sb4_port_2, sb4_port_3, sb4_port_0, sb4_port_1, sb4_port_6, sb4_port_7, sb4_port_4, sb4_port_5, sb4_port_10, sb4_port_11, sb4_port_12, sb4_v;
  wire signed [`W-1:0] sb5_port_8, sb5_port_2, sb5_port_3, sb5_port_0, sb5_port_1, sb5_port_6, sb5_port_7, sb5_port_4, sb5_port_5, sb5_port_10, sb5_port_11, sb5_port_12, sb5_v;
  wire signed [`W-1:0] __AxB_6_port_2, __AxB_6_port_6, __AxB_6_port_11, __AxB_6_v;
  wire signed [`W-1:0] __AxB_4_port_0, __AxB_4_port_6, __AxB_4_port_4, __AxB_4_v;
  wire signed [`W-1:0] __AxB_2_port_0, __AxB_2_port_7, __AxB_2_port_4, __AxB_2_v;
  wire signed [`W-1:0] __AxB_0_port_2, __AxB_0_port_6, __AxB_0_port_4, __AxB_0_v;
  wire signed [`W-1:0] n_1318_port_2, n_1318_port_3, n_1318_port_7, n_1318_port_5, n_1318_v;
  wire signed [`W-1:0] n_1319_port_2, n_1319_port_0, n_1319_v;
  wire signed [`W-1:0] n_1312_port_3, n_1312_port_5, n_1312_v;
  wire signed [`W-1:0] n_1315_port_3, n_1315_port_0, n_1315_v;
  wire signed [`W-1:0] n_1316_port_7, n_1316_port_5, n_1316_v;
  wire signed [`W-1:0] dpc2_XSB_port_2, dpc2_XSB_port_12, dpc2_XSB_v;
  wire signed [`W-1:0] n_1175_port_3, n_1175_port_1, n_1175_v;
  wire signed [`W-1:0] n_1170_port_3, n_1170_port_4, n_1170_v;
  wire signed [`W-1:0] n_1178_port_6, n_1178_port_5, n_1178_v;
  wire signed [`W-1:0] n_1179_port_3, n_1179_port_4, n_1179_v;
  wire signed [`W-1:0] n_578_port_2, n_578_port_3, n_578_port_0, n_578_port_1, n_578_v;
  wire signed [`W-1:0] n_572_port_3, n_572_port_0, n_572_v;
  wire signed [`W-1:0] n_570_port_6, n_570_port_5, n_570_v;
  wire signed [`W-1:0] n_571_port_2, n_571_port_3, n_571_port_1, n_571_v;
  wire signed [`W-1:0] n_318_port_1, n_318_port_4, n_318_v;
  wire signed [`W-1:0] n_319_port_2, n_319_port_4, n_319_v;
  wire signed [`W-1:0] n_312_port_2, n_312_port_3, n_312_v;
  wire signed [`W-1:0] n_310_port_3, n_310_port_0, n_310_v;
  wire signed [`W-1:0] n_311_port_2, n_311_port_3, n_311_v;
  wire signed [`W-1:0] n_317_port_2, n_317_port_0, n_317_v;
  wire signed [`W-1:0] PD_n_0xx0xx0x_port_2, PD_n_0xx0xx0x_port_0, PD_n_0xx0xx0x_v;
  wire signed [`W-1:0] C23_port_7, C23_port_4, C23_v;
  wire signed [`W-1:0] PD_0xx0xx0x_port_4, PD_0xx0xx0x_port_5, PD_0xx0xx0x_v;
  wire signed [`W-1:0] op_T0_dex_port_9, op_T0_dex_port_11, op_T0_dex_v;
  wire signed [`W-1:0] op_T__ora_and_eor_adc_port_6, op_T__ora_and_eor_adc_port_4, op_T__ora_and_eor_adc_v;
  wire signed [`W-1:0] dpc14_SRS_port_2, dpc14_SRS_port_1, dpc14_SRS_v;
  wire signed [`W-1:0] op_T2_ind_x_port_8, op_T2_ind_x_port_6, op_T2_ind_x_v;
  wire signed [`W-1:0] op_T2_ind_y_port_8, op_T2_ind_y_port_6, op_T2_ind_y_v;
  wire signed [`W-1:0] op_plp_pla_port_9, op_plp_pla_port_7, op_plp_pla_v;
  wire signed [`W-1:0] op_T0_txs_port_10, op_T0_txs_port_12, op_T0_txs_v;
  wire signed [`W-1:0] n_66_port_2, n_66_port_3, n_66_port_1, n_66_v;
  wire signed [`W-1:0] n_62_port_2, n_62_port_1, n_62_v;
  wire signed [`W-1:0] n_61_port_3, n_61_port_0, n_61_v;
  wire signed [`W-1:0] n_149_port_3, n_149_port_0, n_149_v;
  wire signed [`W-1:0] n_147_port_3, n_147_port_4, n_147_v;
  wire signed [`W-1:0] n_146_port_2, n_146_port_3, n_146_port_0, n_146_port_1, n_146_port_4, n_146_v;
  wire signed [`W-1:0] n_141_port_2, n_141_port_3, n_141_port_0, n_141_port_1, n_141_port_4, n_141_v;
  wire signed [`W-1:0] _op_set_C_port_7, _op_set_C_port_10, _op_set_C_v;
  wire signed [`W-1:0] op_T5_rti_port_10, op_T5_rti_port_13, op_T5_rti_v;
  wire signed [`W-1:0] op_T5_ind_y_port_8, op_T5_ind_y_port_6, op_T5_ind_y_v;
  wire signed [`W-1:0] op_T5_ind_x_port_9, op_T5_ind_x_port_7, op_T5_ind_x_v;
  wire signed [`W-1:0] op_T3_jsr_port_9, op_T3_jsr_port_10, op_T3_jsr_v;
  wire signed [`W-1:0] op_T5_brk_port_10, op_T5_brk_port_12, op_T5_brk_v;
  wire signed [`W-1:0] ADL_ABL_port_0, ADL_ABL_port_5, ADL_ABL_v;
  wire signed [`W-1:0] n_1371_port_6, n_1371_port_4, n_1371_v;
  wire signed [`W-1:0] n_1376_port_2, n_1376_port_1, n_1376_v;
  wire signed [`W-1:0] n_1377_port_2, n_1377_port_1, n_1377_v;
  wire signed [`W-1:0] n_1374_port_4, n_1374_port_5, n_1374_v;
  wire signed [`W-1:0] n_1375_port_2, n_1375_port_0, n_1375_v;
  wire signed [`W-1:0] n_1379_port_2, n_1379_port_1, n_1379_v;
  wire signed [`W-1:0] n_1724_port_2, n_1724_port_3, n_1724_port_0, n_1724_port_1, n_1724_v;
  wire signed [`W-1:0] n_1194_port_2, n_1194_port_3, n_1194_v;
  wire signed [`W-1:0] n_1195_port_2, n_1195_port_3, n_1195_v;
  wire signed [`W-1:0] n_1192_port_2, n_1192_port_3, n_1192_v;
  wire signed [`W-1:0] n_1190_port_2, n_1190_port_0, n_1190_v;
  wire signed [`W-1:0] n_1191_port_2, n_1191_port_0, n_1191_v;
  wire signed [`W-1:0] n_708_port_2, n_708_port_1, n_708_v;
  wire signed [`W-1:0] n_556_port_2, n_556_port_0, n_556_v;
  wire signed [`W-1:0] n_550_port_3, n_550_port_5, n_550_v;
  wire signed [`W-1:0] n_551_port_2, n_551_port_1, n_551_v;
  wire signed [`W-1:0] n_553_port_3, n_553_port_4, n_553_v;
  wire signed [`W-1:0] C45_port_7, C45_port_4, C45_v;
  wire signed [`W-1:0] x_op_T3_ind_y_port_6, x_op_T3_ind_y_port_7, x_op_T3_ind_y_v;
  wire signed [`W-1:0] op_T__asl_rol_a_port_8, op_T__asl_rol_a_port_10, op_T__asl_rol_a_v;
  wire signed [`W-1:0] n_882_port_3, n_882_port_5, n_882_v;
  wire signed [`W-1:0] n_883_port_2, n_883_port_3, n_883_port_1, n_883_v;
  wire signed [`W-1:0] n_880_port_2, n_880_port_3, n_880_port_0, n_880_v;
  wire signed [`W-1:0] n_334_port_6, n_334_port_5, n_334_v;
  wire signed [`W-1:0] n_335_port_8, n_335_port_10, n_335_v;
  wire signed [`W-1:0] n_336_port_3, n_336_port_1, n_336_port_6, n_336_port_7, n_336_v;
  wire signed [`W-1:0] n_885_port_2, n_885_port_0, n_885_v;
  wire signed [`W-1:0] n_888_port_2, n_888_port_0, n_888_v;
  wire signed [`W-1:0] n_889_port_2, n_889_port_1, n_889_v;
  wire signed [`W-1:0] _AxB_4__C34_port_3, _AxB_4__C34_port_4, _AxB_4__C34_v;
  wire signed [`W-1:0] dpc28_0ADH0_port_2, dpc28_0ADH0_port_0, dpc28_0ADH0_v;
  wire signed [`W-1:0] fetch_port_11, fetch_port_12, fetch_v;
  wire signed [`W-1:0] op_ANDS_port_6, op_ANDS_port_5, op_ANDS_v;
  wire signed [`W-1:0] n_46_port_3, n_46_port_4, n_46_v;
  wire signed [`W-1:0] n_43_port_11, n_43_port_13, n_43_v;
  wire signed [`W-1:0] n_42_port_0, n_42_port_4, n_42_v;
  wire signed [`W-1:0] op_T__cpx_cpy_abs_port_8, op_T__cpx_cpy_abs_port_10, op_T__cpx_cpy_abs_v;
  wire signed [`W-1:0] n_1153_port_3, n_1153_port_0, n_1153_v;
  wire signed [`W-1:0] res_port_2, res_v;
  wire signed [`W-1:0] adl7_port_2, adl7_port_3, adl7_port_0, adl7_port_6, adl7_port_7, adl7_port_4, adl7_port_5, adl7_v;
  wire signed [`W-1:0] adl6_port_2, adl6_port_3, adl6_port_1, adl6_port_6, adl6_port_7, adl6_port_4, adl6_port_5, adl6_v;
  wire signed [`W-1:0] adl5_port_2, adl5_port_3, adl5_port_0, adl5_port_1, adl5_port_7, adl5_port_4, adl5_port_5, adl5_v;
  wire signed [`W-1:0] adl4_port_3, adl4_port_0, adl4_port_1, adl4_port_6, adl4_port_7, adl4_port_4, adl4_port_5, adl4_v;
  wire signed [`W-1:0] adl3_port_2, adl3_port_3, adl3_port_0, adl3_port_1, adl3_port_6, adl3_port_7, adl3_port_4, adl3_v;
  wire signed [`W-1:0] adl2_port_8, adl2_port_2, adl2_port_3, adl2_port_0, adl2_port_1, adl2_port_6, adl2_port_4, adl2_port_5, adl2_v;
  wire signed [`W-1:0] adl1_port_8, adl1_port_2, adl1_port_3, adl1_port_0, adl1_port_1, adl1_port_7, adl1_port_4, adl1_port_5, adl1_v;
  wire signed [`W-1:0] adl0_port_8, adl0_port_3, adl0_port_0, adl0_port_1, adl0_port_6, adl0_port_7, adl0_port_4, adl0_port_5, adl0_v;
  wire signed [`W-1:0] n_1014_port_2, n_1014_port_3, n_1014_port_0, n_1014_port_1, n_1014_v;
  wire signed [`W-1:0] n_0_ADL1_port_2, n_0_ADL1_port_0, n_0_ADL1_v;
  wire signed [`W-1:0] n_0_ADL0_port_3, n_0_ADL0_port_0, n_0_ADL0_v;
  wire signed [`W-1:0] n_0_ADL2_port_2, n_0_ADL2_port_0, n_0_ADL2_v;
  wire signed [`W-1:0] op_T3_abs_idx_port_6, op_T3_abs_idx_port_4, op_T3_abs_idx_v;
  wire signed [`W-1:0] op_jsr_port_8, op_jsr_port_9, op_jsr_v;
  wire signed [`W-1:0] dpc40_ADLPCL_port_0, dpc40_ADLPCL_port_12, dpc40_ADLPCL_v;
  wire signed [`W-1:0] n_593_port_2, n_593_port_1, n_593_v;
  wire signed [`W-1:0] n_929_port_2, n_929_port_3, n_929_port_0, n_929_port_1, n_929_port_4, n_929_v;
  wire signed [`W-1:0] n_1255_port_2, n_1255_port_1, n_1255_v;
  wire signed [`W-1:0] n_1358_port_6, n_1358_port_5, n_1358_v;
  wire signed [`W-1:0] n_1427_port_3, n_1427_port_4, n_1427_v;
  wire signed [`W-1:0] n_1424_port_2, n_1424_port_3, n_1424_port_0, n_1424_port_1, n_1424_v;
  wire signed [`W-1:0] n_1357_port_0, n_1357_port_5, n_1357_v;
  wire signed [`W-1:0] notaluoutmux0_port_2, notaluoutmux0_port_3, notaluoutmux0_port_0, notaluoutmux0_port_1, notaluoutmux0_port_5, notaluoutmux0_v;
  wire signed [`W-1:0] notaluoutmux1_port_2, notaluoutmux1_port_0, notaluoutmux1_port_1, notaluoutmux1_port_4, notaluoutmux1_port_5, notaluoutmux1_v;
  wire signed [`W-1:0] n_533_port_2, n_533_port_1, n_533_v;
  wire signed [`W-1:0] n_531_port_3, n_531_port_0, n_531_v;
  wire signed [`W-1:0] n_538_port_2, n_538_port_1, n_538_v;
  wire signed [`W-1:0] C67_port_6, C67_port_11, C67_v;
  wire signed [`W-1:0] C1x5Reset_port_2, C1x5Reset_port_5, C1x5Reset_v;
  wire signed [`W-1:0] op_T__adc_sbc_port_7, op_T__adc_sbc_port_5, op_T__adc_sbc_v;
  wire signed [`W-1:0] op_T0_cmp_port_6, op_T0_cmp_port_7, op_T0_cmp_v;
  wire signed [`W-1:0] n_1218_port_2, n_1218_port_1, n_1218_v;
  wire signed [`W-1:0] dpc30_ADHPCH_port_10, dpc30_ADHPCH_port_12, dpc30_ADHPCH_v;
  wire signed [`W-1:0] dpc43_DL_DB_port_9, dpc43_DL_DB_port_0, dpc43_DL_DB_v;
  wire signed [`W-1:0] n_23_port_4, n_23_port_5, n_23_v;
  wire signed [`W-1:0] n_21_port_4, n_21_port_5, n_21_v;
  wire signed [`W-1:0] n_20_port_3, n_20_port_5, n_20_v;
  wire signed [`W-1:0] n_27_port_2, n_27_port_3, n_27_port_0, n_27_port_1, n_27_port_4, n_27_v;
  wire signed [`W-1:0] aluanorb0_port_1, aluanorb0_port_6, aluanorb0_port_7, aluanorb0_v;
  wire signed [`W-1:0] n_25_port_3, n_25_port_4, n_25_v;
  wire signed [`W-1:0] n_29_port_2, n_29_port_3, n_29_v;
  wire signed [`W-1:0] n_1694_port_2, n_1694_port_3, n_1694_port_0, n_1694_port_1, n_1694_v;
  wire signed [`W-1:0] a1_port_0, a1_port_1, a1_v;
  wire signed [`W-1:0] a0_port_0, a0_port_1, a0_v;
  wire signed [`W-1:0] a2_port_2, a2_port_1, a2_v;
  wire signed [`W-1:0] a5_port_2, a5_port_0, a5_v;
  wire signed [`W-1:0] a4_port_2, a4_port_0, a4_v;
  wire signed [`W-1:0] a7_port_2, a7_port_1, a7_v;
  wire signed [`W-1:0] n_275_port_3, n_275_port_4, n_275_v;
  wire signed [`W-1:0] n_277_port_2, n_277_port_3, n_277_port_1, n_277_port_4, n_277_port_5, n_277_v;
  wire signed [`W-1:0] n_270_port_2, n_270_port_6, n_270_v;
  wire signed [`W-1:0] n_272_port_8, n_272_port_9, n_272_v;
  wire signed [`W-1:0] n_278_port_2, n_278_port_0, n_278_v;
  wire signed [`W-1:0] n_1486_port_3, n_1486_port_5, n_1486_v;
  wire signed [`W-1:0] n_638_port_2, n_638_port_0, n_638_v;
  wire signed [`W-1:0] n_1408_port_2, n_1408_port_3, n_1408_v;
  wire signed [`W-1:0] n_188_port_4, n_188_port_5, n_188_v;
  wire signed [`W-1:0] n_1400_port_2, n_1400_port_0, n_1400_v;
  wire signed [`W-1:0] n_1402_port_2, n_1402_port_3, n_1402_v;
  wire signed [`W-1:0] op_T0_ora_port_6, op_T0_ora_port_7, op_T0_ora_v;
  wire signed [`W-1:0] n_518_port_2, n_518_port_3, n_518_port_0, n_518_port_1, n_518_v;
  wire signed [`W-1:0] n_519_port_2, n_519_port_4, n_519_v;
  wire signed [`W-1:0] n_510_port_6, n_510_port_4, n_510_v;
  wire signed [`W-1:0] n_513_port_4, n_513_port_5, n_513_v;
  wire signed [`W-1:0] n_515_port_3, n_515_port_5, n_515_v;
  wire signed [`W-1:0] n_1463_port_4, n_1463_port_5, n_1463_v;
  wire signed [`W-1:0] n_453_port_3, n_453_port_1, n_453_v;
  wire signed [`W-1:0] n_1467_port_0, n_1467_port_1, n_1467_v;
  wire signed [`W-1:0] n_980_port_2, n_980_port_0, n_980_v;
  wire signed [`W-1:0] n_1464_port_8, n_1464_port_7, n_1464_v;
  wire signed [`W-1:0] alucout_port_3, alucout_port_0, alucout_v;
  wire signed [`W-1:0] op_brk_rti_port_8, op_brk_rti_port_7, op_brk_rti_v;
  wire signed [`W-1:0] DBZ_port_9, DBZ_port_10, DBZ_v;
  wire signed [`W-1:0] n_1600_port_2, n_1600_port_0, n_1600_v;
  wire signed [`W-1:0] n_1093_port_2, n_1093_port_1, n_1093_v;
  wire signed [`W-1:0] n_1091_port_3, n_1091_port_6, n_1091_v;
  wire signed [`W-1:0] n_1090_port_3, n_1090_port_4, n_1090_v;
  wire signed [`W-1:0] n_1097_port_3, n_1097_port_4, n_1097_v;
  wire signed [`W-1:0] n_1095_port_2, n_1095_port_3, n_1095_port_0, n_1095_port_1, n_1095_v;
  wire signed [`W-1:0] n_1094_port_2, n_1094_port_3, n_1094_port_1, n_1094_v;
  wire signed [`W-1:0] n_1099_port_2, n_1099_port_3, n_1099_v;
  wire signed [`W-1:0] n_1677_port_2, n_1677_port_3, n_1677_v;
  wire signed [`W-1:0] n_1676_port_2, n_1676_port_3, n_1676_v;
  wire signed [`W-1:0] n_1675_port_3, n_1675_port_0, n_1675_v;
  wire signed [`W-1:0] adh3_port_2, adh3_port_3, adh3_port_0, adh3_port_6, adh3_port_4, adh3_port_5, adh3_v;
  wire signed [`W-1:0] adh2_port_3, adh2_port_0, adh2_port_1, adh2_port_6, adh2_port_4, adh2_port_5, adh2_v;
  wire signed [`W-1:0] adh1_port_2, adh1_port_0, adh1_port_1, adh1_port_6, adh1_port_4, adh1_port_5, adh1_v;
  wire signed [`W-1:0] adh0_port_2, adh0_port_3, adh0_port_0, adh0_port_1, adh0_port_6, adh0_port_4, adh0_v;
  wire signed [`W-1:0] adh7_port_2, adh7_port_3, adh7_port_0, adh7_port_1, adh7_port_4, adh7_port_5, adh7_v;
  wire signed [`W-1:0] adh6_port_3, adh6_port_0, adh6_port_1, adh6_port_6, adh6_port_4, adh6_port_5, adh6_v;
  wire signed [`W-1:0] adh5_port_2, adh5_port_3, adh5_port_0, adh5_port_1, adh5_port_4, adh5_port_5, adh5_v;
  wire signed [`W-1:0] adh4_port_2, adh4_port_0, adh4_port_1, adh4_port_6, adh4_port_4, adh4_port_5, adh4_v;
  wire signed [`W-1:0] op_T5_rts_port_12, op_T5_rts_port_14, op_T5_rts_v;
  wire signed [`W-1:0] n_253_port_2, n_253_port_3, n_253_v;
  wire signed [`W-1:0] n_251_port_4, n_251_port_5, n_251_v;
  wire signed [`W-1:0] n_709_port_2, n_709_port_0, n_709_v;
  wire signed [`W-1:0] n_256_port_8, n_256_port_9, n_256_v;
  wire signed [`W-1:0] n_255_port_2, n_255_port_1, n_255_v;
  wire signed [`W-1:0] n_254_port_2, n_254_port_3, n_254_port_1, n_254_v;
  wire signed [`W-1:0] n_700_port_3, n_700_port_1, n_700_v;
  wire signed [`W-1:0] n_1462_port_2, n_1462_port_0, n_1462_v;
  wire signed [`W-1:0] n_1469_port_2, n_1469_port_0, n_1469_port_1, n_1469_v;
  wire signed [`W-1:0] n_714_port_2, n_714_port_1, n_714_v;
  wire signed [`W-1:0] n_1286_port_3, n_1286_port_5, n_1286_v;
  wire signed [`W-1:0] n_1281_port_2, n_1281_port_0, n_1281_v;
  wire signed [`W-1:0] n_1289_port_2, n_1289_port_1, n_1289_v;
  wire signed [`W-1:0] A_B7_port_2, A_B7_port_1, A_B7_v;
  wire signed [`W-1:0] A_B5_port_2, A_B5_port_1, A_B5_v;
  wire signed [`W-1:0] A_B3_port_2, A_B3_port_1, A_B3_v;
  wire signed [`W-1:0] A_B1_port_2, A_B1_port_0, A_B1_v;
  wire signed [`W-1:0] n_392_port_2, n_392_port_3, n_392_v;
  wire signed [`W-1:0] n_390_port_2, n_390_port_0, n_390_v;
  wire signed [`W-1:0] n_396_port_2, n_396_port_1, n_396_v;
  wire signed [`W-1:0] n_397_port_2, n_397_port_0, n_397_v;
  wire signed [`W-1:0] n_1497_port_2, n_1497_port_1, n_1497_v;
  wire signed [`W-1:0] n_936_port_4, n_936_port_5, n_936_v;
  wire signed [`W-1:0] n_937_port_0, n_937_port_4, n_937_v;
  wire signed [`W-1:0] n_935_port_2, n_935_port_3, n_935_port_1, n_935_v;
  wire signed [`W-1:0] n_933_port_2, n_933_port_4, n_933_v;
  wire signed [`W-1:0] n_931_port_2, n_931_port_1, n_931_v;
  wire signed [`W-1:0] op_T2_php_pha_port_9, op_T2_php_pha_port_12, op_T2_php_pha_v;
  wire signed [`W-1:0] ONEBYTE_port_2, ONEBYTE_port_1, ONEBYTE_v;
  wire signed [`W-1:0] NMIP_port_7, NMIP_port_4, NMIP_v;
  wire signed [`W-1:0] n_1075_port_2, n_1075_port_1, n_1075_v;
  wire signed [`W-1:0] n_1076_port_0, n_1076_port_4, n_1076_v;
  wire signed [`W-1:0] n_1071_port_2, n_1071_port_3, n_1071_port_0, n_1071_port_4, n_1071_port_5, n_1071_v;
  wire signed [`W-1:0] n_1070_port_3, n_1070_port_4, n_1070_v;
  wire signed [`W-1:0] n_1073_port_2, n_1073_port_3, n_1073_v;
  wire signed [`W-1:0] n_1072_port_2, n_1072_port_4, n_1072_v;
  wire signed [`W-1:0] abl2_port_3, abl2_port_4, abl2_v;
  wire signed [`W-1:0] abl5_port_0, abl5_port_4, abl5_v;
  wire signed [`W-1:0] abl6_port_0, abl6_port_4, abl6_v;
  wire signed [`W-1:0] n_1619_port_3, n_1619_port_4, n_1619_v;
  wire signed [`W-1:0] notaluvout_port_3, notaluvout_port_5, notaluvout_v;
  wire signed [`W-1:0] n_1140_port_2, n_1140_port_1, n_1140_v;
  wire signed [`W-1:0] n_1614_port_4, n_1614_port_5, n_1614_v;
  wire signed [`W-1:0] n_1145_port_3, n_1145_port_4, n_1145_v;
  wire signed [`W-1:0] n_1147_port_2, n_1147_port_3, n_1147_port_0, n_1147_port_1, n_1147_v;
  wire signed [`W-1:0] dpc34_PCLC_port_12, dpc34_PCLC_port_14, dpc34_PCLC_v;
  wire signed [`W-1:0] aluanorb1_port_7, aluanorb1_port_4, aluanorb1_port_5, aluanorb1_v;
  wire signed [`W-1:0] H1x1_port_8, H1x1_port_4, H1x1_v;
  wire signed [`W-1:0] n_238_port_2, n_238_port_1, n_238_v;
  wire signed [`W-1:0] n_728_port_2, n_728_port_0, n_728_v;
  wire signed [`W-1:0] n_723_port_2, n_723_port_3, n_723_port_0, n_723_port_1, n_723_port_4, n_723_v;
  wire signed [`W-1:0] n_722_port_2, n_722_port_0, n_722_port_1, n_722_port_4, n_722_port_5, n_722_v;
  wire signed [`W-1:0] n_721_port_2, n_721_port_3, n_721_port_0, n_721_port_1, n_721_port_4, n_721_v;
  wire signed [`W-1:0] n_720_port_3, n_720_port_4, n_720_v;
  wire signed [`W-1:0] n_726_port_6, n_726_port_5, n_726_v;
  wire signed [`W-1:0] dpc1_SBY_port_3, dpc1_SBY_port_12, dpc1_SBY_v;
  wire signed [`W-1:0] op_T2_abs_port_7, op_T2_abs_port_5, op_T2_abs_v;
  wire signed [`W-1:0] op_T0_plp_port_9, op_T0_plp_port_10, op_T0_plp_v;
  wire signed [`W-1:0] op_T0_pla_port_9, op_T0_pla_port_11, op_T0_pla_v;
  wire signed [`W-1:0] op_T2_jmp_abs_port_9, op_T2_jmp_abs_port_11, op_T2_jmp_abs_v;
  wire signed [`W-1:0] _C34_port_9, _C34_port_5, _C34_v;
  wire signed [`W-1:0] DA_C01_port_8, DA_C01_port_4, DA_C01_v;
  wire signed [`W-1:0] n_1448_port_2, n_1448_port_0, n_1448_v;
  wire signed [`W-1:0] n_1449_port_2, n_1449_port_1, n_1449_v;
  wire signed [`W-1:0] cclk_port_236, cclk_port_28, cclk_v;
  wire signed [`W-1:0] n_1446_port_3, n_1446_port_4, n_1446_v;
  wire signed [`W-1:0] n_1440_port_2, n_1440_port_1, n_1440_v;
  wire signed [`W-1:0] n_1441_port_2, n_1441_port_1, n_1441_v;
  wire signed [`W-1:0] notRnWprepad_port_6, notRnWprepad_port_7, notRnWprepad_v;
  wire signed [`W-1:0] n_1511_port_2, n_1511_port_1, n_1511_v;
  wire signed [`W-1:0] n_918_port_2, n_918_port_1, n_918_v;
  wire signed [`W-1:0] n_919_port_6, n_919_port_4, n_919_v;
  wire signed [`W-1:0] n_916_port_7, n_916_port_4, n_916_v;
  wire signed [`W-1:0] RnWstretched_port_23, RnWstretched_port_22, RnWstretched_v;
  wire signed [`W-1:0] n_913_port_2, n_913_port_0, n_913_v;
  wire signed [`W-1:0] op_T0_tay_ldy_not_idx_port_8, op_T0_tay_ldy_not_idx_port_7, op_T0_tay_ldy_not_idx_v;
  wire signed [`W-1:0] op_T0_port_2, op_T0_port_1, op_T0_v;
  wire signed [`W-1:0] op_T3_port_2, op_T3_port_0, op_T3_v;
  wire signed [`W-1:0] op_T2_port_2, op_T2_port_0, op_T2_v;
  wire signed [`W-1:0] op_T4_port_2, op_T4_port_1, op_T4_v;
  wire signed [`W-1:0] n_1224_port_2, n_1224_port_0, n_1224_v;
  wire signed [`W-1:0] op_T3_stack_bit_jmp_port_7, op_T3_stack_bit_jmp_port_5, op_T3_stack_bit_jmp_v;
  wire signed [`W-1:0] op_T5_jsr_port_9, op_T5_jsr_port_10, op_T5_jsr_v;
  wire signed [`W-1:0] op_T2_stack_access_port_6, op_T2_stack_access_port_7, op_T2_stack_access_v;
  wire signed [`W-1:0] n_1056_port_2, n_1056_port_0, n_1056_v;
  wire signed [`W-1:0] n_1055_port_3, n_1055_port_5, n_1055_v;
  wire signed [`W-1:0] n_1054_port_2, n_1054_port_0, n_1054_v;
  wire signed [`W-1:0] op_T4_mem_abs_idx_port_6, op_T4_mem_abs_idx_port_4, op_T4_mem_abs_idx_v;
  wire signed [`W-1:0] n_1059_port_0, n_1059_v;
  wire signed [`W-1:0] n_1588_port_2, n_1588_port_1, n_1588_v;
  wire signed [`W-1:0] n_1580_port_3, n_1580_port_0, n_1580_v;
  wire signed [`W-1:0] n_1633_port_2, n_1633_port_0, n_1633_v;
  wire signed [`W-1:0] n_1639_port_2, n_1639_port_0, n_1639_v;
  wire signed [`W-1:0] n_1638_port_2, n_1638_port_1, n_1638_v;
  wire signed [`W-1:0] C34_port_2, C34_port_5, C34_v;
  wire signed [`W-1:0] _DA_ADD2_port_2, _DA_ADD2_port_3, _DA_ADD2_v;
  wire signed [`W-1:0] _DA_ADD1_port_0, _DA_ADD1_port_5, _DA_ADD1_v;
  wire signed [`W-1:0] n_740_port_2, n_740_port_3, n_740_port_0, n_740_port_1, n_740_port_4, n_740_v;
  wire signed [`W-1:0] n_743_port_7, n_743_port_5, n_743_v;
  wire signed [`W-1:0] n_213_port_2, n_213_port_0, n_213_v;
  wire signed [`W-1:0] n_212_port_2, n_212_port_3, n_212_port_1, n_212_v;
  wire signed [`W-1:0] n_747_port_3, n_747_port_0, n_747_v;
  wire signed [`W-1:0] n_210_port_3, n_210_port_0, n_210_port_1, n_210_v;
  wire signed [`W-1:0] n_748_port_3, n_748_port_0, n_748_v;
  wire signed [`W-1:0] n_218_port_2, n_218_port_0, n_218_v;
  wire signed [`W-1:0] notRdy0_port_3, notRdy0_port_4, notRdy0_v;
  wire signed [`W-1:0] notalucout_port_4, notalucout_port_5, notalucout_v;
  wire signed [`W-1:0] dpc36_IPC_port_5, dpc36_IPC_port_10, dpc36_IPC_v;
  wire signed [`W-1:0] op_T0_cpx_cpy_inx_iny_port_6, op_T0_cpx_cpy_inx_iny_port_7, op_T0_cpx_cpy_inx_iny_v;
  wire signed [`W-1:0] n_624_port_2, n_624_port_0, n_624_port_1, n_624_v;
  wire signed [`W-1:0] op_T2_zp_zp_idx_port_4, op_T2_zp_zp_idx_port_5, op_T2_zp_zp_idx_v;
  wire signed [`W-1:0] _C12_port_7, _C12_port_4, _C12_v;
  wire signed [`W-1:0] clk2out_port_0, clk2out_port_1, clk2out_v;
  wire signed [`W-1:0] n_689_port_2, n_689_port_0, n_689_v;
  wire signed [`W-1:0] n_681_port_8, n_681_port_3, n_681_port_1, n_681_port_6, n_681_v;
  wire signed [`W-1:0] n_1471_port_2, n_1471_port_1, n_1471_v;
  wire signed [`W-1:0] n_979_port_2, n_979_port_1, n_979_v;
  wire signed [`W-1:0] n_973_port_2, n_973_port_1, n_973_v;
  wire signed [`W-1:0] n_976_port_2, n_976_port_3, n_976_port_0, n_976_port_1, n_976_port_4, n_976_v;
  wire signed [`W-1:0] n_975_port_3, n_975_port_6, n_975_v;
  wire signed [`W-1:0] op_T__bit_port_9, op_T__bit_port_10, op_T__bit_v;
  wire signed [`W-1:0] op_T0_iny_dey_port_8, op_T0_iny_dey_port_9, op_T0_iny_dey_v;
  wire signed [`W-1:0] n_1270_port_4, n_1270_port_5, n_1270_v;
  wire signed [`W-1:0] op_T__cmp_port_8, op_T__cmp_port_6, op_T__cmp_v;
  wire signed [`W-1:0] n_1618_port_2, n_1618_port_3, n_1618_port_0, n_1618_port_1, n_1618_port_4, n_1618_v;
  wire signed [`W-1:0] op_T0_jsr_port_10, op_T0_jsr_port_12, op_T0_jsr_v;
  wire signed [`W-1:0] n_1610_port_3, n_1610_port_5, n_1610_v;
  wire signed [`W-1:0] op_T2_abs_access_port_9, op_T2_abs_access_port_6, op_T2_abs_access_v;
  wire signed [`W-1:0] n_1613_port_4, n_1613_port_5, n_1613_v;
  wire signed [`W-1:0] n_1033_port_2, n_1033_port_0, n_1033_v;
  wire signed [`W-1:0] n_1034_port_3, n_1034_port_0, n_1034_v;
  wire signed [`W-1:0] n_1037_port_3, n_1037_port_5, n_1037_v;
  wire signed [`W-1:0] alub3_port_2, alub3_port_3, alub3_port_4, alub3_v;
  wire signed [`W-1:0] n_1038_port_2, n_1038_port_1, n_1038_v;
  wire signed [`W-1:0] alub1_port_0, alub1_port_1, alub1_port_4, alub1_v;
  wire signed [`W-1:0] alub0_port_2, alub0_port_3, alub0_port_4, alub0_v;
  wire signed [`W-1:0] alub7_port_3, alub7_port_0, alub7_port_4, alub7_v;
  wire signed [`W-1:0] alub6_port_2, alub6_port_3, alub6_port_4, alub6_v;
  wire signed [`W-1:0] alub5_port_2, alub5_port_3, alub5_port_4, alub5_v;
  wire signed [`W-1:0] alub4_port_3, alub4_port_0, alub4_port_4, alub4_v;
  wire signed [`W-1:0] x_op_T4_rti_port_9, x_op_T4_rti_port_10, x_op_T4_rti_v;
  wire signed [`W-1:0] dpc42_DL_ADH_port_8, dpc42_DL_ADH_port_9, dpc42_DL_ADH_v;
  wire signed [`W-1:0] n_769_port_6, n_769_port_4, n_769_v;
  wire signed [`W-1:0] n_767_port_2, n_767_port_3, n_767_port_0, n_767_port_1, n_767_v;
  wire signed [`W-1:0] n_763_port_2, n_763_port_1, n_763_v;
  wire signed [`W-1:0] n_762_port_3, n_762_port_4, n_762_v;
  wire signed [`W-1:0] n_761_port_4, n_761_port_5, n_761_v;
  wire signed [`W-1:0] op_T3_abs_idx_ind_port_6, op_T3_abs_idx_ind_port_4, op_T3_abs_idx_ind_v;
  wire signed [`W-1:0] op_T2_jsr_port_11, op_T2_jsr_port_13, op_T2_jsr_v;
  wire signed [`W-1:0] DA_C45_port_3, DA_C45_port_1, DA_C45_v;
  wire signed [`W-1:0] n_231_port_2, n_231_port_1, n_231_v;
  wire signed [`W-1:0] _C78_port_3, _C78_port_5, _C78_v;
  wire signed [`W-1:0] n_233_port_2, n_233_port_4, n_233_v;
  wire signed [`W-1:0] n_232_port_0, n_232_port_4, n_232_v;
  wire signed [`W-1:0] n_236_port_3, n_236_port_7, n_236_v;
  wire signed [`W-1:0] n_951_port_3, n_951_port_0, n_951_v;
  wire signed [`W-1:0] n_952_port_3, n_952_port_0, n_952_v;
  wire signed [`W-1:0] n_953_port_2, n_953_port_0, n_953_port_1, n_953_v;
  wire signed [`W-1:0] n_958_port_3, n_958_port_0, n_958_v;
  wire signed [`W-1:0] n_959_port_4, n_959_port_5, n_959_v;
  wire signed [`W-1:0] n_409_port_3, n_409_port_0, n_409_port_5, n_409_v;
  wire signed [`W-1:0] op_T0_eor_port_6, op_T0_eor_port_7, op_T0_eor_v;
  wire signed [`W-1:0] pd1_clearIR_port_6, pd1_clearIR_port_4, pd1_clearIR_v;
  wire signed [`W-1:0] abl3_port_3, abl3_port_4, abl3_v;
  wire signed [`W-1:0] op_T0_jmp_port_8, op_T0_jmp_port_9, op_T0_jmp_v;
  wire signed [`W-1:0] n_1018_port_2, n_1018_port_0, n_1018_v;
  wire signed [`W-1:0] n_1549_port_2, n_1549_port_1, n_1549_v;
  wire signed [`W-1:0] n_1548_port_2, n_1548_port_3, n_1548_port_1, n_1548_v;
  wire signed [`W-1:0] n_1016_port_2, n_1016_port_3, n_1016_port_1, n_1016_v;
  wire signed [`W-1:0] p4_port_2, p4_port_0, p4_port_1, p4_v;
  wire signed [`W-1:0] __AxB1__C01_port_3, __AxB1__C01_port_4, __AxB1__C01_v;
  wire signed [`W-1:0] op_T2_idx_x_xy_port_6, op_T2_idx_x_xy_port_5, op_T2_idx_x_xy_v;
  wire signed [`W-1:0] op_clv_port_8, op_clv_port_9, op_clv_v;
  wire signed [`W-1:0] op_T0_and_port_8, op_T0_and_port_6, op_T0_and_v;
  wire signed [`W-1:0] n_171_port_3, n_171_port_0, n_171_port_1, n_171_v;
  wire signed [`W-1:0] clk0_port_3, clk0_v;
  wire signed [`W-1:0] op_T0_clc_sec_port_8, op_T0_clc_sec_port_9, op_T0_clc_sec_v;
  wire signed [`W-1:0] _C56_port_8, _C56_port_4, _C56_v;
  wire signed [`W-1:0] n_1209_port_3, n_1209_port_5, n_1209_v;
  wire signed [`W-1:0] n_1206_port_2, n_1206_port_3, n_1206_port_0, n_1206_port_1, n_1206_port_4, n_1206_v;
  wire signed [`W-1:0] n_1205_port_4, n_1205_port_10, n_1205_v;
  wire signed [`W-1:0] n_1202_port_2, n_1202_port_3, n_1202_v;
  wire signed [`W-1:0] n_1500_port_3, n_1500_port_5, n_1500_v;
  wire signed [`W-1:0] _ABH3_port_3, _ABH3_port_1, _ABH3_v;
  wire signed [`W-1:0] _ABH2_port_2, _ABH2_port_3, _ABH2_v;
  wire signed [`W-1:0] _ABH1_port_3, _ABH1_port_0, _ABH1_v;
  wire signed [`W-1:0] _ABH0_port_2, _ABH0_port_3, _ABH0_v;
  wire signed [`W-1:0] _ABH7_port_2, _ABH7_port_3, _ABH7_v;
  wire signed [`W-1:0] _ABH6_port_2, _ABH6_port_3, _ABH6_v;
  wire signed [`W-1:0] _ABH5_port_2, _ABH5_port_3, _ABH5_v;
  wire signed [`W-1:0] _ABH4_port_2, _ABH4_port_3, _ABH4_v;
  wire signed [`W-1:0] n_1507_port_2, n_1507_port_3, n_1507_port_1, n_1507_v;
  wire signed [`W-1:0] n_428_port_3, n_428_port_6, n_428_v;
  wire signed [`W-1:0] n_424_port_2, n_424_port_1, n_424_v;
  wire signed [`W-1:0] n_420_port_2, n_420_port_1, n_420_v;
  wire signed [`W-1:0] n_423_port_2, n_423_port_0, n_423_port_1, n_423_v;
  wire signed [`W-1:0] op_sty_cpy_mem_port_8, op_sty_cpy_mem_port_7, op_sty_cpy_mem_v;
  wire signed [`W-1:0] n_1254_port_2, n_1254_port_0, n_1254_port_1, n_1254_v;
  wire signed [`W-1:0] dpc18__DAA_port_2, dpc18__DAA_port_1, dpc18__DAA_v;
  wire signed [`W-1:0] n_1720_port_4, n_1720_port_5, n_1720_v;
  wire signed [`W-1:0] AxB5_port_6, AxB5_port_7, AxB5_v;
  wire signed [`W-1:0] AxB7_port_8, AxB7_port_6, AxB7_v;
  wire signed [`W-1:0] AxB1_port_8, AxB1_port_6, AxB1_v;
  wire signed [`W-1:0] AxB3_port_8, AxB3_port_6, AxB3_v;
  wire signed [`W-1:0] op_T3_ind_y_port_6, op_T3_ind_y_port_7, op_T3_ind_y_v;
  wire signed [`W-1:0] op_T3_ind_x_port_7, op_T3_ind_x_port_10, op_T3_ind_x_v;
  wire signed [`W-1:0] n_1566_port_3, n_1566_port_0, n_1566_v;
  wire signed [`W-1:0] n_1561_port_2, n_1561_port_0, n_1561_v;
  wire signed [`W-1:0] n_1560_port_4, n_1560_port_5, n_1560_v;
  wire signed [`W-1:0] dpc38_PCLADL_port_9, dpc38_PCLADL_port_0, dpc38_PCLADL_v;
  wire signed [`W-1:0] n_1691_port_8, n_1691_port_1, n_1691_port_7, n_1691_v;
  wire signed [`W-1:0] n_1697_port_2, n_1697_port_0, n_1697_v;
  wire signed [`W-1:0] n_1696_port_0, n_1696_port_1, n_1696_v;
  wire signed [`W-1:0] x_op_T3_abs_idx_port_6, x_op_T3_abs_idx_port_4, x_op_T3_abs_idx_v;
  wire signed [`W-1:0] op_from_x_port_6, op_from_x_port_7, op_from_x_v;
  wire signed [`W-1:0] n_855_port_2, n_855_port_0, n_855_v;
  wire signed [`W-1:0] n_854_port_6, n_854_port_4, n_854_v;
  wire signed [`W-1:0] n_850_port_3, n_850_port_0, n_850_v;
  wire signed [`W-1:0] n_853_port_2, n_853_port_3, n_853_v;
  wire signed [`W-1:0] n_852_port_2, n_852_port_3, n_852_v;
  wire signed [`W-1:0] op_T0_cli_sei_port_8, op_T0_cli_sei_port_9, op_T0_cli_sei_v;
  wire signed [`W-1:0] op_T0_ldx_tax_tsx_port_8, op_T0_ldx_tax_tsx_port_6, op_T0_ldx_tax_tsx_v;
  wire signed [`W-1:0] n_1229_port_2, n_1229_port_3, n_1229_v;
  wire signed [`W-1:0] n_1593_port_2, n_1593_port_3, n_1593_v;
  wire signed [`W-1:0] n_1222_port_2, n_1222_port_0, n_1222_v;
  wire signed [`W-1:0] n_1223_port_4, n_1223_port_5, n_1223_v;
  wire signed [`W-1:0] n_1225_port_6, n_1225_port_5, n_1225_v;
  wire signed [`W-1:0] n_1044_port_3, n_1044_port_4, n_1044_v;
  wire signed [`W-1:0] n_1594_port_2, n_1594_port_3, n_1594_v;
  wire signed [`W-1:0] n_1047_port_2, n_1047_port_1, n_1047_v;
  wire signed [`W-1:0] n_198_port_2, n_198_port_3, n_198_v;
  wire signed [`W-1:0] n_628_port_4, n_628_port_5, n_628_v;
  wire signed [`W-1:0] n_629_port_3, n_629_port_5, n_629_v;
  wire signed [`W-1:0] n_626_port_3, n_626_port_6, n_626_v;
  wire signed [`W-1:0] n_196_port_2, n_196_port_0, n_196_v;
  wire signed [`W-1:0] n_625_port_4, n_625_port_5, n_625_v;
  wire signed [`W-1:0] n_191_port_4, n_191_port_5, n_191_v;
  wire signed [`W-1:0] n_192_port_8, n_192_port_4, n_192_v;
  wire signed [`W-1:0] n_442_port_2, n_442_port_0, n_442_v;
  wire signed [`W-1:0] n_440_port_7, n_440_port_10, n_440_v;
  wire signed [`W-1:0] n_441_port_2, n_441_port_0, n_441_v;
  wire signed [`W-1:0] n_445_port_3, n_445_port_4, n_445_v;
  wire signed [`W-1:0] DBNeg_port_3, DBNeg_port_1, DBNeg_v;
  wire signed [`W-1:0] op_T0_tsx_port_9, op_T0_tsx_port_10, op_T0_tsx_v;
  wire signed [`W-1:0] n_994_port_2, n_994_port_3, n_994_port_1, n_994_v;
  wire signed [`W-1:0] n_995_port_2, n_995_port_1, n_995_v;
  wire signed [`W-1:0] n_990_port_3, n_990_port_0, n_990_v;
  wire signed [`W-1:0] n_992_port_2, n_992_port_0, n_992_v;
  wire signed [`W-1:0] n_998_port_2, n_998_port_3, n_998_port_0, n_998_port_1, n_998_port_4, n_998_v;
  wire signed [`W-1:0] n_999_port_2, n_999_port_3, n_999_port_1, n_999_v;
  wire signed [`W-1:0] _op_store_port_2, _op_store_port_3, _op_store_v;
  wire signed [`W-1:0] n_1501_port_1, n_1501_port_4, n_1501_v;
  wire signed [`W-1:0] op_T0_cpx_inx_port_9, op_T0_cpx_inx_port_7, op_T0_cpx_inx_v;
  wire signed [`W-1:0] n_299_port_9, n_299_port_5, n_299_v;
  wire signed [`W-1:0] n_298_port_3, n_298_port_4, n_298_v;
  wire signed [`W-1:0] n_297_port_3, n_297_port_5, n_297_v;
  wire signed [`W-1:0] n_296_port_3, n_296_port_0, n_296_port_1, n_296_port_4, n_296_port_5, n_296_v;
  wire signed [`W-1:0] n_293_port_8, n_293_port_4, n_293_v;
  wire signed [`W-1:0] n_291_port_2, n_291_port_3, n_291_v;
  wire signed [`W-1:0] n_871_port_2, n_871_port_3, n_871_port_0, n_871_port_1, n_871_v;
  wire signed [`W-1:0] n_877_port_3, n_877_port_5, n_877_v;
  wire signed [`W-1:0] n_876_port_2, n_876_port_0, n_876_v;
  wire signed [`W-1:0] n_875_port_3, n_875_port_5, n_875_v;
  wire signed [`W-1:0] n_956_port_2, n_956_port_1, n_956_v;

  wire pipedpc28_v;
  wire n_460_v;
  wire n_469_v;
  wire n_1162_v;
  wire n_1161_v;
  wire n_1529_v;
  wire n_1528_v;
  wire n_1527_v;
  wire n_599_v;
  wire n_9_v;
  wire n_663_v;
  wire n_666_v;
  wire n_1450_v;
  wire n_1126_v;
  wire n_1124_v;
  wire n_1121_v;
  wire n_360_v;
  wire n_94_v;
  wire n_95_v;
  wire n_698_v;
  wire pipeVectorA2_v;
  wire n_745_v;
  wire n_562_v;
  wire pclp1_v;
  wire pclp3_v;
  wire pclp5_v;
  wire pclp7_v;
  wire n_1252_v;
  wire n_796_v;
  wire n_799_v;
  wire pd7_v;
  wire pd6_v;
  wire pd5_v;
  wire pd4_v;
  wire pd3_v;
  wire pd2_v;
  wire pd1_v;
  wire pd0_v;
  wire n_339_v;
  wire n_323_v;
  wire n_897_v;
  wire n_50_v;
  wire n_55_v;
  wire n_1360_v;
  wire n_521_v;
  wire n_526_v;
  wire pchp4_v;
  wire pchp6_v;
  wire pchp0_v;
  wire pchp2_v;
  wire n_1341_v;
  wire n_509_v;
  wire n_18_v;
  wire n_15_v;
  wire n_1269_v;
  wire n_265_v;
  wire n_1411_v;
  wire n_1061_v;
  wire n_1606_v;
  wire notidl0_v;
  wire pipeT3out_v;
  wire n_1472_v;
  wire n_1477_v;
  wire n_1291_v;
  wire n_902_v;
  wire pipeUNK18_v;
  wire pipeUNK16_v;
  wire pipeUNK17_v;
  wire pipeUNK14_v;
  wire pipeUNK15_v;
  wire pipeUNK12_v;
  wire pipeUNK13_v;
  wire pipeUNK11_v;
  wire n_1624_v;
  wire n_1625_v;
  wire n_223_v;
  wire n_226_v;
  wire n_415_v;
  wire n_1452_v;
  wire n_968_v;
  wire pipeUNK34_v;
  wire pipeUNK35_v;
  wire pipeUNK36_v;
  wire pipeUNK37_v;
  wire pipeUNK30_v;
  wire pipeUNK31_v;
  wire pipeUNK32_v;
  wire pipeUNK33_v;
  wire pipeUNK39_v;
  wire n_1020_v;
  wire n_1027_v;
  wire n_756_v;
  wire n_759_v;
  wire pipephi2Reset0_v;
  wire n_1579_v;
  wire n_1574_v;
  wire pipeT2out_v;
  wire n_459_v;
  wire n_982_v;
  wire pipe_WR_phi2_v;
  wire DC78_phi2_v;
  wire n_610_v;
  wire p2_v;
  wire p3_v;
  wire p0_v;
  wire n_1533_v;
  wire n_1395_v;
  wire n_644_v;
  wire n_865_v;
  wire pipeT4out_v;
  wire pipeT_SYNC_v;
  wire n_671_v;
  wire n_675_v;
  wire n_1404_v;
  wire n_1113_v;
  wire n_805_v;
  wire n_1272_v;
  wire n_1276_v;
  wire n_1274_v;
  wire n_126_v;
  wire n_653_v;
  wire pipe_VEC_v;
  wire n_266_v;
  wire n_1132_v;
  wire notdor1_v;
  wire notdor0_v;
  wire notdor3_v;
  wire notdor2_v;
  wire notdor5_v;
  wire notdor4_v;
  wire notdor7_v;
  wire notdor6_v;
  wire n_1570_v;
  wire n_101_v;
  wire n_581_v;
  wire n_1338_v;
  wire n_1333_v;
  wire n_597_v;
  wire nots3_v;
  wire nots2_v;
  wire nots1_v;
  wire nots0_v;
  wire nots7_v;
  wire nots6_v;
  wire nots5_v;
  wire nots4_v;
  wire n_1683_v;
  wire n_88_v;
  wire n_785_v;
  wire n_1177_v;
  wire C78_phi2_v;
  wire n_69_v;
  wire n_559_v;
  wire n_47_v;
  wire n_590_v;
  wire n_598_v;
  wire pipeBRtaken_v;
  wire pipeUNK41_v;
  wire pipeUNK40_v;
  wire pipeUNK42_v;
  wire n_24_v;
  wire n_1693_v;
  wire pipephi2Reset0x_v;
  wire n_1409_v;
  wire n_512_v;
  wire pipeVectorA0_v;
  wire pipeVectorA1_v;
  wire n_1602_v;
  wire pipeT5out_v;
  wire n_1679_v;
  wire n_1674_v;
  wire n_1673_v;
  wire n_393_v;
  wire n_398_v;
  wire pipeUNK09_v;
  wire pipeUNK08_v;
  wire pipeUNK05_v;
  wire pipeUNK04_v;
  wire pipeUNK07_v;
  wire pipeUNK06_v;
  wire pipeUNK01_v;
  wire pipeUNK03_v;
  wire pipeUNK02_v;
  wire n_1149_v;
  wire pipe_T0_v;
  wire n_1447_v;
  wire pipeUNK23_v;
  wire pipeUNK22_v;
  wire pipeUNK21_v;
  wire pipeUNK20_v;
  wire pipeUNK27_v;
  wire pipeUNK26_v;
  wire pipeUNK29_v;
  wire pipeUNK28_v;
  wire n_1581_v;
  wire n_688_v;
  wire n_680_v;
  wire notalu4_v;
  wire notalu5_v;
  wire notalu6_v;
  wire notalu7_v;
  wire notalu0_v;
  wire notalu1_v;
  wire notalu2_v;
  wire notalu3_v;
  wire notidl6_v;
  wire n_760_v;
  wire notidl4_v;
  wire notidl1_v;
  wire n_402_v;
  wire n_408_v;
  wire p1_v;
  wire _TWOCYCLE_phi1_v;
  wire notidl5_v;
  wire n_1565_v;
  wire n_1699_v;
  wire n_1049_v;
  wire n_1221_v;
  wire n_190_v;
  wire n_621_v;
  wire notidl7_v;
  wire notidl3_v;
  wire notidl2_v;
  wire n_993_v;
  wire n_1505_v;
  wire n_1509_v;
  wire n_878_v;

  spice_pin_input pin_4286(nmi, nmi_v, nmi_port_2);
  spice_pin_input pin_4287(irq, irq_v, irq_port_2);
  spice_pin_input pin_4285(rdy, rdy_v, rdy_port_3);
  spice_pin_input pin_4282(clk0, clk0_v, clk0_port_3);
  spice_pin_input pin_4281(so, so_v, so_port_3);
  spice_pin_input pin_4278(res, res_v, res_port_2);

  spice_pin_output pin_4284(clk2out, clk2out_v);
  spice_pin_output pin_4283(clk1out, clk1out_v);
  spice_pin_output pin_4280(sync, sync_v);
  spice_pin_output pin_4268(ab14, ab14_v);
  spice_pin_output pin_4264(ab10, ab10_v);
  spice_pin_output pin_4266(ab12, ab12_v);
  spice_pin_output pin_4260(ab6, ab6_v);
  spice_pin_output pin_4261(ab7, ab7_v);
  spice_pin_output pin_4262(ab8, ab8_v);
  spice_pin_output pin_4263(ab9, ab9_v);
  spice_pin_output pin_4269(ab15, ab15_v);
  spice_pin_output pin_4265(ab11, ab11_v);
  spice_pin_output pin_4267(ab13, ab13_v);
  spice_pin_output pin_4279(rw, rw_v);
  spice_pin_output pin_4255(ab1, ab1_v);
  spice_pin_output pin_4254(ab0, ab0_v);
  spice_pin_output pin_4257(ab3, ab3_v);
  spice_pin_output pin_4256(ab2, ab2_v);
  spice_pin_output pin_4259(ab5, ab5_v);
  spice_pin_output pin_4258(ab4, ab4_v);

  spice_pin_bidirectional pin_4277(db7_i, db7_o, db7_t, db7_v, db7_port_5);
  spice_pin_bidirectional pin_4276(db6_i, db6_o, db6_t, db6_v, db6_port_5);
  spice_pin_bidirectional pin_4275(db5_i, db5_o, db5_t, db5_v, db5_port_5);
  spice_pin_bidirectional pin_4274(db4_i, db4_o, db4_t, db4_v, db4_port_5);
  spice_pin_bidirectional pin_4273(db3_i, db3_o, db3_t, db3_v, db3_port_5);
  spice_pin_bidirectional pin_4272(db2_i, db2_o, db2_t, db2_v, db2_port_5);
  spice_pin_bidirectional pin_4271(db1_i, db1_o, db1_t, db1_v, db1_port_5);
  spice_pin_bidirectional pin_4270(db0_i, db0_o, db0_t, db0_v, db0_port_5);

  spice_transistor_nmos_gnd g_4389((~n_1662_v[`W-1]|~n_781_v[`W-1]), n_553_v, n_553_port_4);
  spice_transistor_nmos_gnd g_4388((~dor3_v[`W-1]|~RnWstretched_v[`W-1]), n_1613_v, n_1613_port_5);
  spice_transistor_nmos_gnd g_4383((~ir7_v[`W-1]|~irline3_v[`W-1]|~ir2_v[`W-1]|~notir3_v[`W-1]|~clock1_v[`W-1]|~notir4_v[`W-1]|~notir6_v[`W-1]), op_T0_cli_sei_v, op_T0_cli_sei_port_9);
  spice_transistor_nmos_gnd g_4382((~irline3_v[`W-1]|~notir5_v[`W-1]|~ir4_v[`W-1]|~notir3_v[`W-1]|~ir7_v[`W-1]|~_t3_v[`W-1]|~ir2_v[`W-1]), x_op_T3_plp_pla_v, x_op_T3_plp_pla_port_10);
  spice_transistor_nmos_gnd g_4381((~notir4_v[`W-1]|~irline3_v[`W-1]|~ir6_v[`W-1]|~notir7_v[`W-1]|~ir2_v[`W-1]|~notir3_v[`W-1]|~notir5_v[`W-1]), op_clv_v, op_clv_port_9);
  spice_transistor_nmos_gnd g_4380((~notir3_v[`W-1]|~x_op_push_pull_v[`W-1]|~ir0_v[`W-1]|~ir2_v[`W-1]), op_implied_v, op_implied_port_6);
  spice_transistor_nmos_gnd g_4387((~op_T5_ind_y_v[`W-1]|~op_T4_abs_idx_v[`W-1]), n_595_v, n_595_port_5);
  spice_transistor_nmos_gnd g_4386((~dor3_v[`W-1]|~RnWstretched_v[`W-1]), n_643_v, n_643_port_4);
  spice_transistor_nmos_gnd g_4385((~notir3_v[`W-1]|~ir2_v[`W-1]|~ir4_v[`W-1]|~clock1_v[`W-1]|~notir5_v[`W-1]|~notir7_v[`W-1]|~ir6_v[`W-1]|~notir1_v[`W-1]), op_T0_tax_v, op_T0_tax_port_10);
  spice_transistor_nmos_gnd g_4384((~_t4_v[`W-1]|~notir3_v[`W-1]|~notir4_v[`W-1]), op_T4_mem_abs_idx_v, op_T4_mem_abs_idx_port_6);
  spice_transistor_nmos t3178(~dpc39_PCLPCL_v[`W-1], pcl0_v, n_488_v, pcl0_port_1, n_488_port_3);
  spice_transistor_nmos t3179(~dpc39_PCLPCL_v[`W-1], pcl3_v, n_723_v, pcl3_port_1, n_723_port_3);
  spice_transistor_nmos t3174(~dpc39_PCLPCL_v[`W-1], pcl4_v, n_208_v, pcl4_port_1, n_208_port_3);
  spice_transistor_nmos t3175(~dpc39_PCLPCL_v[`W-1], pcl7_v, n_1647_v, pcl7_port_2, n_1647_port_3);
  spice_transistor_nmos t3176(~dpc39_PCLPCL_v[`W-1], pcl6_v, n_1458_v, pcl6_port_1, n_1458_port_3);
  spice_transistor_nmos t3177(~dpc39_PCLPCL_v[`W-1], pcl1_v, n_976_v, pcl1_port_1, n_976_port_2);
  spice_transistor_nmos_gnd t3172(~n_366_v[`W-1], op_SRS_v, op_SRS_port_2);
  spice_transistor_nmos t3173(~dpc39_PCLPCL_v[`W-1], pcl5_v, n_72_v, pcl5_port_1, n_72_port_3);
  spice_transistor_nmos_gnd t985(~n_790_v[`W-1], op_rmw_v, op_rmw_port_0);
  spice_transistor_nmos t989(~dpc37_PCLDB_v[`W-1], idb0_v, n_488_v, idb0_port_6, n_488_port_1);
  spice_transistor_nmos_gnd t988(~sb1_v[`W-1], n_320_v, n_320_port_0);
  spice_transistor_nmos_gnd t1538(pipeUNK42_v, n_253_v, n_253_port_2);
  spice_transistor_nmos_gnd t1539(~n_1552_v[`W-1], dpc14_SRS_v, dpc14_SRS_port_2);
  spice_transistor_nmos_gnd t1531(~_ABL2_v[`W-1], abl2_v, abl2_port_3);
  spice_transistor_nmos_gnd g_4608((n_1291_v|n_1693_v), n_1312_v, n_1312_port_5);
  spice_transistor_nmos_gnd g_4609((~n_36_v[`W-1]|~n_320_v[`W-1]), n_735_v, n_735_port_4);
  spice_transistor_nmos_gnd g_4606((~op_T__iny_dey_v[`W-1]|~op_T0_tay_ldy_not_idx_v[`W-1]|~op_T0_ldy_mem_v[`W-1]), n_616_v, n_616_port_6);
  spice_transistor_nmos_gnd g_4604((~n_602_v[`W-1]|~n_1247_v[`W-1]|~cclk_v[`W-1]), dpc2_XSB_v, dpc2_XSB_port_12);
  spice_transistor_nmos_gnd g_4602((~n_885_v[`W-1]|~n_954_v[`W-1]|~op_T__bit_v[`W-1]), n_513_v, n_513_port_5);
  spice_transistor_nmos_gnd g_4603((~notRdy0_v[`W-1]|~n_383_v[`W-1]), n_917_v, n_917_port_5);
  spice_transistor_nmos_gnd g_4600((~alub0_v[`W-1]|~alua0_v[`W-1]), aluanorb0_v, aluanorb0_port_7);
  spice_transistor_nmos_gnd g_4601((n_805_v|~n_43_v[`W-1]), n_1534_v, n_1534_port_5);
  spice_transistor_nmos_gnd t3365(~adl5_v[`W-1], n_1094_v, n_1094_port_1);
  spice_transistor_nmos_vdd t167(~dor5_v[`W-1], n_373_v, n_373_port_0);
  spice_transistor_nmos_vdd t166(~n_1296_v[`W-1], ab11_v, ab11_port_0);
  spice_transistor_nmos_gnd t162(~n_272_v[`W-1], n_952_v, n_952_port_0);
  spice_transistor_nmos t1571(~cclk_v[`W-1], n_658_v, y4_v, n_658_port_0, y4_port_2);
  spice_transistor_nmos_gnd t1762(~n_761_v[`W-1], n_1056_v, n_1056_port_0);
  spice_transistor_nmos t2363(~dpc24_ACSB_v[`W-1], sb0_v, n_146_v, sb0_port_10, n_146_port_2);
  spice_transistor_nmos t2366(~dpc24_ACSB_v[`W-1], sb3_v, n_1654_v, sb3_port_10, n_1654_port_3);
  spice_transistor_nmos t2367(~dpc24_ACSB_v[`W-1], sb4_v, n_1344_v, sb4_port_11, n_1344_port_1);
  spice_transistor_nmos t2364(~dpc24_ACSB_v[`W-1], sb1_v, n_929_v, sb1_port_9, n_929_port_3);
  spice_transistor_nmos t2365(~dpc24_ACSB_v[`W-1], n_1618_v, sb2_v, n_1618_port_1, sb2_port_9);
  spice_transistor_nmos t2368(~dpc24_ACSB_v[`W-1], sb5_v, n_831_v, sb5_port_8, n_831_port_2);
  spice_transistor_nmos t2369(~dpc24_ACSB_v[`W-1], n_326_v, sb6_v, n_326_port_3, sb6_port_11);
  spice_transistor_nmos_vdd t570(~n_772_v[`W-1], dpc17_SUMS_v, dpc17_SUMS_port_1);
  spice_transistor_nmos_gnd t571(~s5_v[`W-1], n_496_v, n_496_port_1);
  spice_transistor_nmos_gnd t572(~pclp2_v[`W-1], n_481_v, n_481_port_0);
  spice_transistor_nmos_vdd t578(~dor2_v[`W-1], n_520_v, n_520_port_0);
  spice_transistor_nmos_gnd t2189(~n_890_v[`W-1], n_1694_v, n_1694_port_1);
  spice_transistor_nmos_gnd t2184(p3_v, n_1194_v, n_1194_port_2);
  spice_transistor_nmos_gnd t2185(~n_350_v[`W-1], n_988_v, n_988_port_1);
  spice_transistor_nmos_gnd t2180(n_398_v, n_321_v, n_321_port_2);
  spice_transistor_nmos_gnd g_4598((~n_43_v[`W-1]|n_1509_v), n_611_v, n_611_port_5);
  spice_transistor_nmos_gnd g_4599((~n_1613_v[`W-1]|~RnWstretched_v[`W-1]), n_42_v, n_42_port_4);
  spice_transistor_nmos_gnd g_4597((~op_T0_plp_v[`W-1]|~x_op_T4_rti_v[`W-1]), n_327_v, n_327_port_4);
  spice_transistor_nmos_gnd g_4594((~n_467_v[`W-1]|~op_branch_done_v[`W-1]|~n_1211_v[`W-1]), n_10_v, n_10_port_6);
  spice_transistor_nmos_gnd g_4595((~brk_done_v[`W-1]|n_760_v), INTG_v, INTG_port_6);
  spice_transistor_nmos_gnd g_4592((~ir3_v[`W-1]|~_t2_v[`W-1]), op_T2_ADL_ADD_v, op_T2_ADL_ADD_port_4);
  spice_transistor_nmos_gnd g_4593((~op_T2_ind_v[`W-1]|~op_T2_zp_zp_idx_v[`W-1]), n_1225_v, n_1225_port_6);
  spice_transistor_nmos_gnd g_4590((~ir1_v[`W-1]|~ir0_v[`W-1]), n_1133_v, n_1133_port_4);
  spice_transistor_nmos_gnd g_4591((~Reset0_v[`W-1]|n_323_v|n_671_v), n_14_v, n_14_port_5);
  spice_transistor_nmos_gnd t1983(~n_1033_v[`W-1], dpc21_ADDADL_v, dpc21_ADDADL_port_9);
  spice_transistor_nmos_gnd t1982(~idb3_v[`W-1], n_457_v, n_457_port_1);
  spice_transistor_nmos_gnd t1329(~dpc22__DSA_v[`W-1], n_306_v, n_306_port_0);
  spice_transistor_nmos_gnd t1189(n_526_v, pclp0_v, pclp0_port_1);
  spice_transistor_nmos_gnd t1188(~n_1392_v[`W-1], n_284_v, n_284_port_0);
  spice_transistor_nmos t1183(~cclk_v[`W-1], x1_v, n_1709_v, x1_port_0, n_1709_port_0);
  spice_transistor_nmos_gnd t1181(~abl1_v[`W-1], n_842_v, n_842_port_0);
  spice_transistor_nmos_gnd t1180(~abl1_v[`W-1], n_66_v, n_66_port_1);
  spice_transistor_nmos_gnd t1184(~n_0_ADL1_v[`W-1], adl1_v, adl1_port_1);
  spice_transistor_nmos_gnd t711(n_1529_v, n_91_v, n_91_port_0);
  spice_transistor_nmos t2197(~dpc27_SBADH_v[`W-1], adh4_v, sb4_v, adh4_port_4, sb4_port_9);
  spice_transistor_nmos t372(~dpc10_ADLADD_v[`W-1], adl0_v, alub0_v, adl0_port_1, alub0_port_2);
  spice_transistor_nmos_gnd t373(~C1x5Reset_v[`W-1], n_1054_v, n_1054_port_0);
  spice_transistor_nmos_gnd t370(~n_198_v[`W-1], n_424_v, n_424_port_1);
  spice_transistor_nmos_gnd t2522(~op_T0_eor_v[`W-1], n_837_v, n_837_port_0);
  spice_transistor_nmos t374(~dpc4_SSB_v[`W-1], n_694_v, sb1_v, n_694_port_1, sb1_port_2);
  spice_transistor_nmos_gnd t375(~n_869_v[`W-1], ab13_v, ab13_port_1);
  spice_transistor_nmos t2526(~dpc38_PCLADL_v[`W-1], n_72_v, adl5_v, n_72_port_2, adl5_port_4);
  spice_transistor_nmos t2527(~dpc38_PCLADL_v[`W-1], adl6_v, n_1458_v, adl6_port_4, n_1458_port_1);
  spice_transistor_nmos_gnd g_4837(((~n_888_v[`W-1]|~n_118_v[`W-1])&~n_264_v[`W-1]), n_480_v, n_480_port_4);
  spice_transistor_nmos_gnd g_4836((~n_790_v[`W-1]&~_op_store_v[`W-1]), n_1137_v, n_1137_port_4);
  spice_transistor_nmos_gnd g_4831((~n_761_v[`W-1]&~n_149_v[`W-1]), n_233_v, n_233_port_4);
  spice_transistor_nmos_gnd g_4832((~alua5_v[`W-1]&~alub5_v[`W-1]), n_477_v, n_477_port_5);
  spice_transistor_nmos g_4839((~cp1_v[`W-1]&~fetch_v[`W-1]), n_1641_v, n_119_v, n_1641_port_3, n_119_port_3);
  spice_transistor_nmos t3118(~dpc2_XSB_v[`W-1], n_1694_v, sb2_v, n_1694_port_2, sb2_port_10);
  spice_transistor_nmos t3119(~dpc2_XSB_v[`W-1], n_242_v, sb3_v, n_242_port_2, sb3_port_11);
  spice_transistor_nmos t3116(~dpc2_XSB_v[`W-1], n_1724_v, sb6_v, n_1724_port_2, sb6_port_12);
  spice_transistor_nmos_gnd t3117(~n_1256_v[`W-1], dpc15_ANDS_v, dpc15_ANDS_port_9);
  spice_transistor_nmos t3115(~dpc2_XSB_v[`W-1], n_578_v, sb5_v, n_578_port_1, sb5_port_10);
  spice_transistor_nmos_gnd t2645(notidl3_v, idl3_v, idl3_port_0);
  spice_transistor_nmos_gnd t2641(~idb2_v[`W-1], n_1573_v, n_1573_port_0);
  spice_transistor_nmos_gnd t2640(notalu5_v, alu5_v, alu5_port_3);
  spice_transistor_nmos_vdd t2643(~n_625_v[`W-1], dpc3_SBX_v, dpc3_SBX_port_9);
  spice_transistor_nmos_gnd t967(~n_368_v[`W-1], n_218_v, n_218_port_0);
  spice_transistor_nmos t963(~dpc6_SBS_v[`W-1], sb0_v, s0_v, sb0_port_3, s0_port_1);
  spice_transistor_nmos t962(~cclk_v[`W-1], n_1694_v, x2_v, n_1694_port_0, x2_port_0);
  spice_transistor_nmos_vdd t961(~cclk_v[`W-1], idb3_v, idb3_port_1);
  spice_transistor_nmos_gnd t1046(pchp2_v, n_1496_v, n_1496_port_0);
  spice_transistor_nmos t1047(~cclk_v[`W-1], n_1251_v, y7_v, n_1251_port_0, y7_port_0);
  spice_transistor_nmos_gnd t1040(~adh1_v[`W-1], n_1267_v, n_1267_port_0);
  spice_transistor_nmos_gnd t1518(~s3_v[`W-1], n_34_v, n_34_port_1);
  spice_transistor_nmos_gnd t1519(pchp6_v, n_652_v, n_652_port_0);
  spice_transistor_nmos_gnd t1048(~adl4_v[`W-1], n_1519_v, n_1519_port_0);
  spice_transistor_nmos_gnd g_4309((~notir4_v[`W-1]|~_t3_v[`W-1]|~irline3_v[`W-1]|~ir2_v[`W-1]|~ir3_v[`W-1]), op_T3_branch_v, op_T3_branch_port_8);
  spice_transistor_nmos_gnd g_4628((~n_43_v[`W-1]|n_265_v), n_818_v, n_818_port_5);
  spice_transistor_nmos_gnd g_4629((~dpc36_IPC_v[`W-1]|~n_937_v[`W-1]), n_1345_v, n_1345_port_7);
  spice_transistor_nmos_gnd g_4620((~n_1464_v[`W-1]|n_902_v), n_1109_v, n_1109_port_9);
  spice_transistor_nmos_gnd g_4621((~notir6_v[`W-1]|~notir1_v[`W-1]), op_lsr_ror_dec_inc_v, op_lsr_ror_dec_inc_port_4);
  spice_transistor_nmos_gnd g_4622((~notir7_v[`W-1]|~notir0_v[`W-1]|~ir5_v[`W-1]|~clock2_v[`W-1]|~notir6_v[`W-1]), op_T__cmp_v, op_T__cmp_port_8);
  spice_transistor_nmos_gnd g_4623((~n_43_v[`W-1]|n_688_v), n_1223_v, n_1223_port_5);
  spice_transistor_nmos_gnd g_4624((~n_689_v[`W-1]|~notRdy0_v[`W-1]), VEC0_v, VEC0_port_6);
  spice_transistor_nmos_gnd g_4625((~RnWstretched_v[`W-1]|~n_1463_v[`W-1]), n_1076_v, n_1076_port_4);
  spice_transistor_nmos_gnd g_4626((~n_1247_v[`W-1]|~n_228_v[`W-1]|~cclk_v[`W-1]), dpc30_ADHPCH_v, dpc30_ADHPCH_port_12);
  spice_transistor_nmos_gnd g_4627((~n_1154_v[`W-1]|~n_819_v[`W-1]), n_1380_v, n_1380_port_5);
  spice_transistor_nmos_gnd t3438(~n_906_v[`W-1], dpc19_ADDSB7_v, dpc19_ADDSB7_port_2);
  spice_transistor_nmos_gnd t3349(n_598_v, n_1260_v, n_1260_port_2);
  spice_transistor_nmos t1533(~dpc3_SBX_v[`W-1], x7_v, sb7_v, x7_port_1, sb7_port_2);
  spice_transistor_nmos t3347(~dpc11_SBADD_v[`W-1], sb7_v, alua7_v, sb7_port_10, alua7_port_3);
  spice_transistor_nmos_gnd t3346(pipeUNK08_v, n_954_v, n_954_port_3);
  spice_transistor_nmos_gnd t3345(n_1049_v, n_507_v, n_507_port_2);
  spice_transistor_nmos_gnd t3344(~cp1_v[`W-1], n_839_v, n_839_port_1);
  spice_transistor_nmos_vdd t3340(~cclk_v[`W-1], sb5_v, sb5_port_12);
  spice_transistor_nmos_vdd t1536(~n_520_v[`W-1], db2_v, db2_port_3);
  spice_transistor_nmos_gnd t1534(~a5_v[`W-1], n_1719_v, n_1719_port_0);
  spice_transistor_nmos_vdd t149(~n_154_v[`W-1], dpc20_ADDSB06_v, dpc20_ADDSB06_port_0);
  spice_transistor_nmos_gnd t148(~n_154_v[`W-1], n_75_v, n_75_port_0);
  spice_transistor_nmos_gnd t145(~idb7_v[`W-1], n_789_v, n_789_port_0);
  spice_transistor_nmos_gnd t144(~op_T0_lda_v[`W-1], n_397_v, n_397_port_0);
  spice_transistor_nmos_gnd t147(~idb0_v[`W-1], n_624_v, n_624_port_0);
  spice_transistor_nmos_gnd t146(~AxB3_v[`W-1], n_884_v, n_884_port_0);
  spice_transistor_nmos_gnd t141(~x5_v[`W-1], n_1017_v, n_1017_port_0);
  spice_transistor_nmos t142(~cp1_v[`W-1], n_1424_v, idl2_v, n_1424_port_0, idl2_port_1);
  spice_transistor_nmos_gnd t2346(~y0_v[`W-1], n_1025_v, n_1025_port_1);
  spice_transistor_nmos_gnd t2252(~abh2_v[`W-1], n_994_v, n_994_port_1);
  spice_transistor_nmos_vdd t2250(~abh2_v[`W-1], n_1545_v, n_1545_port_1);
  spice_transistor_nmos_gnd t2251(~abh2_v[`W-1], n_1034_v, n_1034_port_0);
  spice_transistor_nmos_gnd t551(~n_1417_v[`W-1], clk1out_v, clk1out_port_0);
  spice_transistor_nmos t2254(~dpc27_SBADH_v[`W-1], sb1_v, adh1_v, sb1_port_8, adh1_port_4);
  spice_transistor_nmos_gnd t2255(~dpc12_0ADD_v[`W-1], alua2_v, alua2_port_1);
  spice_transistor_nmos_gnd g_4314((~ir4_v[`W-1]|~notir5_v[`W-1]|~irline3_v[`W-1]|~ir2_v[`W-1]|~notir6_v[`W-1]|~ir7_v[`W-1]|~ir3_v[`W-1]|~_t5_v[`W-1]), op_T5_rts_v, op_T5_rts_port_14);
  spice_transistor_nmos_gnd g_4315((~ir4_v[`W-1]|~irline3_v[`W-1]|~ir2_v[`W-1]|~ir6_v[`W-1]|~ir3_v[`W-1]|~ir5_v[`W-1]|~_t2_v[`W-1]|~ir7_v[`W-1]), op_T2_brk_v, op_T2_brk_port_10);
  spice_transistor_nmos_gnd g_4316((~ir7_v[`W-1]|~irline3_v[`W-1]|~ir6_v[`W-1]|~_t3_v[`W-1]|~ir2_v[`W-1]|~ir4_v[`W-1]|~notir5_v[`W-1]|~ir3_v[`W-1]), op_T3_jsr_v, op_T3_jsr_port_10);
  spice_transistor_nmos_gnd g_4317((~notir5_v[`W-1]|~ir4_v[`W-1]|~ir3_v[`W-1]|~irline3_v[`W-1]|~ir7_v[`W-1]|~ir2_v[`W-1]|~ir6_v[`W-1]), op_jsr_v, op_jsr_port_9);
  spice_transistor_nmos_gnd g_4305((~n_964_v[`W-1]|~n_732_v[`W-1]), n_17_v, n_17_port_6);
  spice_transistor_nmos_gnd g_4310((~ir3_v[`W-1]|~ir5_v[`W-1]|~irline3_v[`W-1]|~ir2_v[`W-1]|~ir4_v[`W-1]|~ir7_v[`W-1]), op_brk_rti_v, op_brk_rti_port_8);
  spice_transistor_nmos_gnd g_4311((~ir7_v[`W-1]|~ir3_v[`W-1]|~irline3_v[`W-1]|~ir5_v[`W-1]|~ir2_v[`W-1]|~ir4_v[`W-1]|~clock1_v[`W-1]), op_T0_brk_rti_v, op_T0_brk_rti_port_9);
  spice_transistor_nmos_gnd t312(~n_445_v[`W-1], sync_v, sync_port_0);
  spice_transistor_nmos_gnd g_4312((~ir4_v[`W-1]|~ir7_v[`W-1]|~notir6_v[`W-1]|~notir3_v[`W-1]|~notir2_v[`W-1]|~irline3_v[`W-1]|~clock1_v[`W-1]), op_T0_jmp_v, op_T0_jmp_port_9);
  spice_transistor_nmos_gnd t317(~_ABH2_v[`W-1], abh2_v, abh2_port_0);
  spice_transistor_nmos_gnd g_4313((~_t2_v[`W-1]|~ir3_v[`W-1]|~irline3_v[`W-1]|~notir4_v[`W-1]|~ir2_v[`W-1]), op_T2_branch_v, op_T2_branch_port_7);
  spice_transistor_nmos_gnd g_4817((~alub1_v[`W-1]&~alua1_v[`W-1]), aluanandb1_v, aluanandb1_port_5);
  spice_transistor_nmos_gnd g_4816((~DA_C45_v[`W-1]&~n_647_v[`W-1]), n_757_v, n_757_port_5);
  spice_transistor_nmos_gnd g_4814(((~n_311_v[`W-1]|~dpc34_PCLC_v[`W-1])&~n_919_v[`W-1]), n_1229_v, n_1229_port_3);
  spice_transistor_nmos_gnd t3131(~n_531_v[`W-1], n_1255_v, n_1255_port_1);
  spice_transistor_nmos_vdd t3132(~n_531_v[`W-1], dpc13_ORS_v, dpc13_ORS_port_8);
  spice_transistor_nmos_vdd t3133(~dor7_v[`W-1], n_298_v, n_298_port_3);
  spice_transistor_nmos t3134(~cclk_v[`W-1], _ABH4_v, n_999_v, _ABH4_port_2, n_999_port_3);
  spice_transistor_nmos_gnd t3137(notidl5_v, idl5_v, idl5_port_1);
  spice_transistor_nmos_gnd t2086(~a4_v[`W-1], n_556_v, n_556_port_0);
  spice_transistor_nmos_gnd t2084(~n_646_v[`W-1], n_470_v, n_470_port_2);
  spice_transistor_nmos_gnd t2089(n_1121_v, n_291_v, n_291_port_2);
  spice_transistor_nmos_gnd t1280(~pd5_clearIR_v[`W-1], n_928_v, n_928_port_1);
  spice_transistor_nmos_gnd t1282(~pch1_v[`W-1], n_1070_v, n_1070_port_3);
  spice_transistor_nmos t941(~dpc16_EORS_v[`W-1], n_1469_v, n_277_v, n_1469_port_0, n_277_port_1);
  spice_transistor_nmos t940(~dpc16_EORS_v[`W-1], __AxB_4_v, n_296_v, __AxB_4_port_0, n_296_port_0);
  spice_transistor_nmos t943(~dpc16_EORS_v[`W-1], n_304_v, n_177_v, n_304_port_1, n_177_port_1);
  spice_transistor_nmos t942(~dpc16_EORS_v[`W-1], __AxB_6_v, n_722_v, __AxB_6_port_2, n_722_port_1);
  spice_transistor_nmos_gnd t2889(~ir4_v[`W-1], notir4_v, notir4_port_25);
  spice_transistor_nmos t2883(~n_771_v[`W-1], n_430_v, n_465_v, n_430_port_3, n_465_port_1);
  spice_transistor_nmos_gnd t2881(n_745_v, n_241_v, n_241_port_2);
  spice_transistor_nmos_gnd g_4642((~VEC1_v[`W-1]|~VEC0_v[`W-1]), _VEC_v, _VEC_port_8);
  spice_transistor_nmos_gnd g_4643((~op_T2_stack_access_v[`W-1]|~n_1222_v[`W-1]), n_1090_v, n_1090_port_4);
  spice_transistor_nmos_gnd g_4640((~n_441_v[`W-1]|~n_1247_v[`W-1]|~cclk_v[`W-1]), dpc1_SBY_v, dpc1_SBY_port_12);
  spice_transistor_nmos_gnd g_4641((n_55_v|~cclk_v[`W-1]), n_628_v, n_628_port_5);
  spice_transistor_nmos_gnd g_4646((~notir3_v[`W-1]|~notir4_v[`W-1]|~_t3_v[`W-1]), op_T3_abs_idx_v, op_T3_abs_idx_port_6);
  spice_transistor_nmos_gnd g_4647((~_t3_v[`W-1]|~notir3_v[`W-1]|~notir4_v[`W-1]), x_op_T3_abs_idx_v, x_op_T3_abs_idx_port_6);
  spice_transistor_nmos_gnd g_4644((~n_1448_v[`W-1]|~n_182_v[`W-1]), n_1619_v, n_1619_port_4);
  spice_transistor_nmos_gnd g_4648((~notRdy0_v[`W-1]|~n_1716_v[`W-1]), n_180_v, n_180_port_5);
  spice_transistor_nmos_gnd g_4649((~n_959_v[`W-1]|~notRdy0_v[`W-1]), n_1154_v, n_1154_port_5);
  spice_transistor_nmos t1476(~cclk_v[`W-1], n_676_v, _ABH1_v, n_676_port_0, _ABH1_port_0);
  spice_transistor_nmos_gnd t1472(n_339_v, n_543_v, n_543_port_0);
  spice_transistor_nmos_vdd t1471(~n_91_v[`W-1], dpc15_ANDS_v, dpc15_ANDS_port_0);
  spice_transistor_nmos_gnd t1126(~n_1025_v[`W-1], n_564_v, n_564_port_1);
  spice_transistor_nmos_gnd t1122(n_402_v, n_834_v, n_834_port_2);
  spice_transistor_nmos_gnd t129(~n_1369_v[`W-1], n_1462_v, n_1462_port_0);
  spice_transistor_nmos t128(~dpc4_SSB_v[`W-1], n_1389_v, sb2_v, n_1389_port_0, sb2_port_1);
  spice_transistor_nmos_gnd t121(pclp7_v, n_1647_v, n_1647_port_0);
  spice_transistor_nmos t127(~dpc4_SSB_v[`W-1], n_998_v, sb3_v, n_998_port_0, sb3_port_1);
  spice_transistor_nmos_gnd t124(~DBZ_v[`W-1], _DBZ_v, _DBZ_port_0);
  spice_transistor_nmos_gnd t1496(~n_1105_v[`W-1], cp1_v, cp1_port_50);
  spice_transistor_nmos t1723(~dpc5_SADL_v[`W-1], adl3_v, n_998_v, adl3_port_3, n_998_port_3);
  spice_transistor_nmos t1722(~dpc5_SADL_v[`W-1], adl4_v, n_3_v, adl4_port_4, n_3_port_3);
  spice_transistor_nmos t1721(~dpc5_SADL_v[`W-1], adl5_v, n_280_v, adl5_port_3, n_280_port_3);
  spice_transistor_nmos_gnd t1720(~notir5_v[`W-1], n_503_v, n_503_port_0);
  spice_transistor_nmos t1727(~dpc5_SADL_v[`W-1], n_721_v, adl7_v, n_721_port_3, adl7_port_2);
  spice_transistor_nmos t1724(~dpc5_SADL_v[`W-1], adl2_v, n_1389_v, adl2_port_3, n_1389_port_2);
  spice_transistor_nmos_gnd t1729(~_ABL1_v[`W-1], abl1_v, abl1_port_3);
  spice_transistor_nmos_gnd t338(~pclp0_v[`W-1], n_488_v, n_488_port_0);
  spice_transistor_nmos_gnd t332(~n_182_v[`W-1], n_442_v, n_442_port_0);
  spice_transistor_nmos_vdd t333(~dor1_v[`W-1], n_798_v, n_798_port_1);
  spice_transistor_nmos_gnd g_4789((~n_1440_v[`W-1]&(~n_1002_v[`W-1]|~n_1081_v[`W-1]|~op_T0_sbc_v[`W-1])), n_779_v, n_779_port_5);
  spice_transistor_nmos_gnd g_4788((~aluaorb0_v[`W-1]&~aluanandb0_v[`W-1]), __AxB_0_v, __AxB_0_port_6);
  spice_transistor_nmos_gnd g_4787(((~n_1316_v[`W-1]|~n_715_v[`W-1])&~n_1386_v[`W-1]), n_484_v, n_484_port_3);
  spice_transistor_nmos g_4784((~cp1_v[`W-1]&~ADL_ABL_v[`W-1]), n_1016_v, _ABL1_v, n_1016_port_3, _ABL1_port_3);
  spice_transistor_nmos g_4782((~ADL_ABL_v[`W-1]&~cp1_v[`W-1]), _ABL3_v, n_1507_v, _ABL3_port_3, n_1507_port_3);
  spice_transistor_nmos_gnd g_4879((~n_735_v[`W-1]|(~n_36_v[`W-1]&~n_320_v[`W-1])), dasb1_v, dasb1_port_5);
  spice_transistor_nmos_gnd g_4878(((~notRdy0_v[`W-1]&pipeT5out_v)|(~n_16_v[`W-1]&pipeT4out_v)), n_468_v, n_468_port_6);
  spice_transistor_nmos_gnd g_4871(((pipeUNK01_v&~n_1401_v[`W-1])|(~DBNeg_v[`W-1]&n_1269_v)), n_626_v, n_626_port_6);
  spice_transistor_nmos_gnd g_4870(((~n_253_v[`W-1]&~n_270_v[`W-1])|(~n_507_v[`W-1]&~n_1224_v[`W-1])|(~n_954_v[`W-1]&~n_206_v[`W-1])|(pipeUNK16_v&~n_279_v[`W-1])), n_1082_v, n_1082_port_10);
  spice_transistor_nmos_gnd g_4873(((~n_270_v[`W-1]&~n_1662_v[`W-1])|(pipeUNK17_v&~n_553_v[`W-1])|(~n_1573_v[`W-1]&~n_781_v[`W-1])), n_845_v, n_845_port_8);
  spice_transistor_nmos_gnd g_4872(((~n_1492_v[`W-1]&~n_270_v[`W-1])|(~n_781_v[`W-1]&~n_1600_v[`W-1])|(~n_1457_v[`W-1]&pipeUNK04_v)), n_1495_v, n_1495_port_8);
  spice_transistor_nmos_gnd g_4875((~n_1629_v[`W-1]|(~n_753_v[`W-1]&~n_1135_v[`W-1])), dasb5_v, dasb5_port_5);
  spice_transistor_nmos_gnd g_4877(((~n_16_v[`W-1]&pipeT_SYNC_v)|(~notRdy0_v[`W-1]&pipeT2out_v)), n_1091_v, n_1091_port_6);
  spice_transistor_nmos_gnd g_4876(((~op_sta_cmp_v[`W-1]&~n_335_v[`W-1])|~op_T2_pha_v[`W-1]), n_1037_v, n_1037_port_5);
  spice_transistor_nmos_gnd t1222(~n_1675_v[`W-1], ir6_v, ir6_port_42);
  spice_transistor_nmos_gnd t2068(pipe_VEC_v, n_1578_v, n_1578_port_1);
  spice_transistor_nmos_vdd t2066(~n_1028_v[`W-1], RnWstretched_v, RnWstretched_port_23);
  spice_transistor_nmos_gnd t1267(pipeUNK26_v, n_1714_v, n_1714_port_1);
  spice_transistor_nmos_gnd t1262(~n_1620_v[`W-1], ir3_v, ir3_port_1);
  spice_transistor_nmos t1228(~cclk_v[`W-1], n_1592_v, a7_v, n_1592_port_0, a7_port_1);
  spice_transistor_nmos_gnd t691(~pch6_v[`W-1], n_278_v, n_278_port_0);
  spice_transistor_nmos_gnd t922(~notRdy0_v[`W-1], n_372_v, n_372_port_0);
  spice_transistor_nmos_gnd t693(~n_567_v[`W-1], n_1026_v, n_1026_port_0);
  spice_transistor_nmos_gnd t692(~n_567_v[`W-1], n_171_v, n_171_port_0);
  spice_transistor_nmos_gnd t695(~n_551_v[`W-1], n_8_v, n_8_port_1);
  spice_transistor_nmos_vdd t694(~n_567_v[`W-1], n_322_v, n_322_port_1);
  spice_transistor_nmos t696(~cclk_v[`W-1], n_1620_v, notir3_v, n_1620_port_0, notir3_port_1);
  spice_transistor_nmos_gnd t929(notdor2_v, dor2_v, dor2_port_3);
  spice_transistor_nmos_gnd t2605(~n_1660_v[`W-1], n_855_v, n_855_port_2);
  spice_transistor_nmos_vdd t2606(~n_1660_v[`W-1], n_1100_v, n_1100_port_3);
  spice_transistor_nmos_gnd t1009(~ir2_v[`W-1], notir2_v, notir2_port_0);
  spice_transistor_nmos_gnd t1000(~n_1110_v[`W-1], n_771_v, n_771_port_1);
  spice_transistor_nmos_gnd t1006(pipeUNK27_v, n_920_v, n_920_port_1);
  spice_transistor_nmos_gnd g_4668((~dor6_v[`W-1]|~RnWstretched_v[`W-1]), n_471_v, n_471_port_4);
  spice_transistor_nmos_gnd g_4669((~n_916_v[`W-1]|pipeUNK36_v|~n_1137_v[`W-1]|~notRdy0_v[`W-1]), short_circuit_idx_add_v, short_circuit_idx_add_port_7);
  spice_transistor_nmos_gnd g_4664((~cclk_v[`W-1]|~n_255_v[`W-1]|~n_1247_v[`W-1]), dpc31_PCHPCH_v, dpc31_PCHPCH_port_12);
  spice_transistor_nmos_gnd g_4665((~n_134_v[`W-1]|n_1276_v), n_930_v, n_930_port_4);
  spice_transistor_nmos_gnd g_4666((~op_T2_abs_access_v[`W-1]|~n_646_v[`W-1]), n_773_v, n_773_port_5);
  spice_transistor_nmos_gnd g_4667((~n_930_v[`W-1]|~n_470_v[`W-1]), n_1286_v, n_1286_port_5);
  spice_transistor_nmos_gnd g_4660((~n_1542_v[`W-1]|~n_783_v[`W-1]), n_1253_v, n_1253_port_7);
  spice_transistor_nmos_gnd g_4661((~C34_v[`W-1]|~__AxB_4_v[`W-1]), _AxB_4__C34_v, _AxB_4__C34_port_4);
  spice_transistor_nmos_gnd g_4662((~dor5_v[`W-1]|~RnWstretched_v[`W-1]), n_1720_v, n_1720_port_5);
  spice_transistor_nmos_gnd g_4663((~n_1720_v[`W-1]|~RnWstretched_v[`W-1]), n_373_v, n_373_port_4);
  spice_transistor_nmos_vdd t104(~n_963_v[`W-1], ab14_v, ab14_port_0);
  spice_transistor_nmos_vdd t109(~abh3_v[`W-1], n_1296_v, n_1296_port_0);
  spice_transistor_nmos_gnd t2472(~db4_v[`W-1], n_1075_v, n_1075_port_1);
  spice_transistor_nmos_gnd t2473(~dpc34_PCLC_v[`W-1], n_1007_v, n_1007_port_1);
  spice_transistor_nmos_gnd t2470(~x0_v[`W-1], n_987_v, n_987_port_1);
  spice_transistor_nmos t2476(~dpc31_PCHPCH_v[`W-1], pch7_v, n_1206_v, pch7_port_2, n_1206_port_1);
  spice_transistor_nmos t2477(~dpc31_PCHPCH_v[`W-1], pch4_v, n_27_v, pch4_port_2, n_27_port_1);
  spice_transistor_nmos t2475(~dpc31_PCHPCH_v[`W-1], pch6_v, n_652_v, pch6_port_2, n_652_port_1);
  spice_transistor_nmos t2478(~dpc31_PCHPCH_v[`W-1], pch5_v, n_1301_v, pch5_port_2, n_1301_port_1);
  spice_transistor_nmos t2479(~dpc31_PCHPCH_v[`W-1], pch2_v, n_1496_v, pch2_port_1, n_1496_port_1);
  spice_transistor_nmos_vdd t1(~n_1608_v[`W-1], ab13_v, ab13_port_0);
  spice_transistor_nmos_gnd t1929(n_1450_v, n_1499_v, n_1499_port_0);
  spice_transistor_nmos_gnd t1928(~n_1609_v[`W-1], ir5_v, ir5_port_0);
  spice_transistor_nmos_gnd t1927(~n_1560_v[`W-1], n_1081_v, n_1081_port_2);
  spice_transistor_nmos_gnd t1920(~alu1_v[`W-1], _DA_ADD1_v, _DA_ADD1_port_0);
  spice_transistor_nmos_vdd t1922(~n_1152_v[`W-1], ab2_v, ab2_port_0);
  spice_transistor_nmos_vdd t481(~n_670_v[`W-1], n_1417_v, n_1417_port_0);
  spice_transistor_nmos_gnd t482(~n_994_v[`W-1], ab10_v, ab10_port_1);
  spice_transistor_nmos_gnd t489(~n_1439_v[`W-1], n_518_v, n_518_port_1);
  spice_transistor_nmos_vdd t1749(~n_1596_v[`W-1], dpc27_SBADH_v, dpc27_SBADH_port_0);
  spice_transistor_nmos_gnd t1748(~n_1596_v[`W-1], n_1271_v, n_1271_port_0);
  spice_transistor_nmos_gnd t1745(~n_966_v[`W-1], n_1635_v, n_1635_port_1);
  spice_transistor_nmos_gnd t1747(n_559_v, n_770_v, n_770_port_1);
  spice_transistor_nmos_vdd t1746(~n_966_v[`W-1], dpc29_0ADH17_v, dpc29_0ADH17_port_2);
  spice_transistor_nmos_gnd g_4343((~n_519_v[`W-1]|~cp1_v[`W-1]), n_127_v, n_127_port_5);
  spice_transistor_nmos g_4857((~ADH_ABH_v[`W-1]&~cp1_v[`W-1]), _ABH6_v, n_880_v, _ABH6_port_3, n_880_port_3);
  spice_transistor_nmos g_4858((~ADH_ABH_v[`W-1]&~cp1_v[`W-1]), _ABH3_v, n_883_v, _ABH3_port_3, n_883_port_3);
  spice_transistor_nmos_gnd g_4342((~C1x5Reset_v[`W-1]|~INTG_v[`W-1]), D1x1_v, D1x1_port_6);
  spice_transistor_nmos t83(~H1x1_v[`W-1], idb2_v, Pout2_v, idb2_port_0, Pout2_port_0);
  spice_transistor_nmos_gnd t2256(n_610_v, n_582_v, n_582_port_2);
  spice_transistor_nmos t2257(~dpc0_YSB_v[`W-1], n_1251_v, sb7_v, n_1251_port_1, sb7_port_8);
  spice_transistor_nmos t2745(~dpc37_PCLDB_v[`W-1], n_723_v, idb3_v, n_723_port_2, idb3_port_9);
  spice_transistor_nmos t2746(~dpc37_PCLDB_v[`W-1], n_976_v, idb1_v, n_976_port_1, idb1_port_8);
  spice_transistor_nmos_vdd t2598(~cclk_v[`W-1], idb6_v, idb6_port_9);
  spice_transistor_nmos_gnd t2049(~n_1455_v[`W-1], n_1412_v, n_1412_port_0);
  spice_transistor_nmos t2592(~dpc13_ORS_v[`W-1], n_404_v, n_296_v, n_404_port_2, n_296_port_5);
  spice_transistor_nmos_gnd t2044(~op_rti_rts_v[`W-1], n_1377_v, n_1377_port_1);
  spice_transistor_nmos_gnd t2623(~alu5_v[`W-1], n_761_v, n_761_port_4);
  spice_transistor_nmos_vdd t2622(~n_1153_v[`W-1], n_659_v, n_659_port_2);
  spice_transistor_nmos_gnd t2621(~n_1153_v[`W-1], n_1639_v, n_1639_port_2);
  spice_transistor_nmos_gnd t900(~aluanorb1_v[`W-1], A_B1_v, A_B1_port_0);
  spice_transistor_nmos_gnd t905(~n_635_v[`W-1], ab14_v, ab14_port_1);
  spice_transistor_nmos t1985(~dpc1_SBY_v[`W-1], y3_v, sb3_v, y3_port_2, sb3_port_8);
  spice_transistor_nmos t1984(~dpc40_ADLPCL_v[`W-1], pcl7_v, adl7_v, pcl7_port_1, adl7_port_4);
  spice_transistor_nmos_gnd t1327(~n_1484_v[`W-1], n_1491_v, n_1491_port_1);
  spice_transistor_nmos_gnd t1024(~n_471_v[`W-1], db6_v, db6_port_0);
  spice_transistor_nmos t1505(~dpc0_YSB_v[`W-1], n_1491_v, sb2_v, n_1491_port_2, sb2_port_3);
  spice_transistor_nmos_gnd t3420(~notRdy0_v[`W-1], n_1440_v, n_1440_port_1);
  spice_transistor_nmos_gnd t2458(~abh7_v[`W-1], n_1153_v, n_1153_port_0);
  spice_transistor_nmos_gnd t2459(~abh7_v[`W-1], n_659_v, n_659_port_1);
  spice_transistor_nmos t2450(~dpc30_ADHPCH_v[`W-1], pch1_v, adh1_v, pch1_port_1, adh1_port_5);
  spice_transistor_nmos_gnd t2452(~_ABH5_v[`W-1], abh5_v, abh5_port_3);
  spice_transistor_nmos t2453(~dpc30_ADHPCH_v[`W-1], pch0_v, adh0_v, pch0_port_1, adh0_port_4);
  spice_transistor_nmos_gnd t2454(~abh1_v[`W-1], n_617_v, n_617_port_0);
  spice_transistor_nmos_gnd t2455(~abh1_v[`W-1], n_676_v, n_676_port_2);
  spice_transistor_nmos_vdd t2457(~abh7_v[`W-1], n_1639_v, n_1639_port_0);
  spice_transistor_nmos_vdd t1182(~abl1_v[`W-1], n_1479_v, n_1479_port_0);
  spice_transistor_nmos_gnd t3057(~n_1467_v[`W-1], cclk_v, cclk_port_236);
  spice_transistor_nmos_vdd t3055(~n_1364_v[`W-1], dpc16_EORS_v, dpc16_EORS_port_9);
  spice_transistor_nmos_gnd t3054(~n_1364_v[`W-1], n_108_v, n_108_port_1);
  spice_transistor_nmos_vdd t3504(~cclk_v[`W-1], idb4_v, idb4_port_10);
  spice_transistor_nmos_vdd t3501(~n_951_v[`W-1], n_642_v, n_642_port_3);
  spice_transistor_nmos_gnd t3500(~n_951_v[`W-1], n_1152_v, n_1152_port_2);
  spice_transistor_nmos_vdd t3502(~cclk_v[`W-1], sb2_v, sb2_port_12);
  spice_transistor_nmos_vdd t2902(~n_830_v[`W-1], dpc23_SBAC_v, dpc23_SBAC_port_11);
  spice_transistor_nmos_gnd t2900(n_902_v, n_1289_v, n_1289_port_1);
  spice_transistor_nmos_gnd t2901(~n_830_v[`W-1], n_1047_v, n_1047_port_1);
  spice_transistor_nmos_gnd t1901(~C67_v[`W-1], _C67_v, _C67_port_0);
  spice_transistor_nmos_gnd t1907(n_1020_v, n_1277_v, n_1277_port_0);
  spice_transistor_nmos_gnd t1906(~s7_v[`W-1], n_548_v, n_548_port_0);
  spice_transistor_nmos_vdd t1760(~cclk_v[`W-1], idb2_v, idb2_port_4);
  spice_transistor_nmos_gnd g_4302((~n_1047_v[`W-1]|~n_1247_v[`W-1]|~cclk_v[`W-1]), dpc23_SBAC_v, dpc23_SBAC_port_12);
  spice_transistor_nmos_gnd g_4301((~n_1312_v[`W-1]|n_1149_v), n_264_v, n_264_port_8);
  spice_transistor_nmos_gnd g_4300((~n_646_v[`W-1]|~n_440_v[`W-1]), n_812_v, n_812_port_4);
  spice_transistor_nmos_gnd g_4307((~n_1371_v[`W-1]|~n_307_v[`W-1]|~n_1433_v[`W-1]|~n_1293_v[`W-1]), n_620_v, n_620_port_7);
  spice_transistor_nmos_gnd g_4304((~n_43_v[`W-1]|n_1505_v), n_830_v, n_830_port_5);
  spice_transistor_nmos_gnd g_4308((~n_43_v[`W-1]|n_460_v), n_692_v, n_692_port_5);
  spice_transistor_nmos_gnd t3193(~n_837_v[`W-1], op_EORS_v, op_EORS_port_2);
  spice_transistor_nmos_gnd t3196(~idb7_v[`W-1], n_423_v, n_423_port_1);
  spice_transistor_nmos_gnd t3194(n_590_v, alucin_v, alucin_port_1);
  spice_transistor_nmos t3195(~dpc4_SSB_v[`W-1], n_332_v, sb0_v, n_332_port_3, sb0_port_12);
  spice_transistor_nmos_gnd t2029(n_878_v, n_631_v, n_631_port_2);
  spice_transistor_nmos_vdd t2028(~cclk_v[`W-1], adh7_v, adh7_port_2);
  spice_transistor_nmos t521(~dpc21_ADDADL_v[`W-1], adl3_v, alu3_v, adl3_port_0, alu3_port_0);
  spice_transistor_nmos t520(~cp1_v[`W-1], n_87_v, idl1_v, n_87_port_1, idl1_port_0);
  spice_transistor_nmos t1599(~dpc1_SBY_v[`W-1], y2_v, sb2_v, y2_port_2, sb2_port_6);
  spice_transistor_nmos t1590(~dpc14_SRS_v[`W-1], aluanandb1_v, notaluoutmux0_v, aluanandb1_port_0, notaluoutmux0_port_2);
  spice_transistor_nmos t1591(~dpc14_SRS_v[`W-1], notaluoutmux1_v, n_681_v, notaluoutmux1_port_2, n_681_port_1);
  spice_transistor_nmos t1592(~dpc14_SRS_v[`W-1], n_350_v, n_740_v, n_350_port_1, n_740_port_3);
  spice_transistor_nmos t1593(~dpc14_SRS_v[`W-1], n_1071_v, n_1063_v, n_1071_port_4, n_1063_port_2);
  spice_transistor_nmos t1594(~dpc14_SRS_v[`W-1], n_296_v, n_477_v, n_296_port_3, n_477_port_1);
  spice_transistor_nmos t1595(~dpc14_SRS_v[`W-1], n_277_v, n_336_v, n_277_port_3, n_336_port_1);
  spice_transistor_nmos t1596(~dpc14_SRS_v[`W-1], n_722_v, n_1318_v, n_722_port_4, n_1318_port_2);
  spice_transistor_nmos_gnd t1980(~adh4_v[`W-1], n_212_v, n_212_port_1);
  spice_transistor_nmos t588(~dpc43_DL_DB_v[`W-1], idb3_v, n_1661_v, idb3_port_0, n_1661_port_1);
  spice_transistor_nmos_gnd t2112(~x1_v[`W-1], n_1434_v, n_1434_port_0);
  spice_transistor_nmos t585(~dpc43_DL_DB_v[`W-1], idb0_v, n_719_v, idb0_port_5, n_719_port_2);
  spice_transistor_nmos_gnd t855(~_op_branch_bit6_v[`W-1], n_846_v, n_846_port_1);
  spice_transistor_nmos_gnd t1640(~n_1521_v[`W-1], n_242_v, n_242_port_1);
  spice_transistor_nmos t1641(~dpc1_SBY_v[`W-1], y1_v, sb1_v, y1_port_2, sb1_port_5);
  spice_transistor_nmos_gnd t2648(~_C12_v[`W-1], C12_v, C12_port_2);
  spice_transistor_nmos_gnd t1960(~pcl6_v[`W-1], n_232_v, n_232_port_0);
  spice_transistor_nmos_gnd t3038(~n_147_v[`W-1], db4_v, db4_port_3);
  spice_transistor_nmos_gnd t3030(~n_90_v[`W-1], p6_v, p6_port_1);
  spice_transistor_nmos_vdd t3035(~n_769_v[`W-1], n_1072_v, n_1072_port_2);
  spice_transistor_nmos_gnd t3036(~pcl4_v[`W-1], n_1643_v, n_1643_port_3);
  spice_transistor_nmos t1961(~dpc5_SADL_v[`W-1], adl0_v, n_332_v, adl0_port_4, n_332_port_1);
  spice_transistor_nmos_gnd t1963(~s2_v[`W-1], n_1190_v, n_1190_port_0);
  spice_transistor_nmos t1964(~cclk_v[`W-1], n_1300_v, notir2_v, n_1300_port_2, notir2_port_19);
  spice_transistor_nmos_gnd t1967(~n_1691_v[`W-1], n_110_v, n_110_port_1);
  spice_transistor_nmos_gnd t1969(pclp3_v, n_723_v, n_723_port_0);
  spice_transistor_nmos_gnd t3372(~_ABH1_v[`W-1], abh1_v, abh1_port_3);
  spice_transistor_nmos t3373(~dpc40_ADLPCL_v[`W-1], pcl1_v, adl1_v, pcl1_port_2, adl1_port_8);
  spice_transistor_nmos_gnd t3370(pipeUNK35_v, n_238_v, n_238_port_1);
  spice_transistor_nmos_gnd t2920(n_1674_v, n_772_v, n_772_port_2);
  spice_transistor_nmos t3375(~dpc40_ADLPCL_v[`W-1], pcl3_v, adl3_v, pcl3_port_2, adl3_port_7);
  spice_transistor_nmos_gnd t1785(~db4_v[`W-1], n_490_v, n_490_port_1);
  spice_transistor_nmos t1782(~dpc1_SBY_v[`W-1], y7_v, sb7_v, y7_port_1, sb7_port_4);
  spice_transistor_nmos g_4728((~cp1_v[`W-1]&~fetch_v[`W-1]), n_1605_v, n_541_v, n_1605_port_5, n_541_port_3);
  spice_transistor_nmos_gnd g_4725((~n_595_v[`W-1]&~_op_branch_done_v[`W-1]), n_192_v, n_192_port_8);
  spice_transistor_nmos g_4726((~ADH_ABH_v[`W-1]&~cp1_v[`W-1]), _ABH7_v, n_494_v, _ABH7_port_3, n_494_port_3);
  spice_transistor_nmos_gnd g_4722((~Pout3_v[`W-1]&~op_T0_adc_sbc_v[`W-1]), n_673_v, n_673_port_4);
  spice_transistor_nmos_gnd g_4897(((~_C12_v[`W-1]&~n_681_v[`W-1])|~n_1691_v[`W-1]), C23_v, C23_port_7);
  spice_transistor_nmos_gnd g_4896((~n_748_v[`W-1]|(~C67_v[`W-1]&~A_B7_v[`W-1])), _C78_v, _C78_port_5);
  spice_transistor_nmos_gnd g_4895((~n_1253_v[`W-1]|(~n_783_v[`W-1]&~n_1542_v[`W-1])), n_515_v, n_515_port_5);
  spice_transistor_nmos_gnd g_4894((n_1126_v|(~VEC1_v[`W-1]&~notRdy0_v[`W-1])), n_1290_v, n_1290_port_5);
  spice_transistor_nmos_gnd g_4893(((~op_T2_ADL_ADD_v[`W-1]&~n_638_v[`W-1])|(~op_T2_stack_v[`W-1]|~notRdy0_v[`W-1]|~op_T3_stack_bit_jmp_v[`W-1]|~op_T4_rti_v[`W-1]|~op_T4_brk_jsr_v[`W-1]|~op_T3_ind_x_v[`W-1])), n_604_v, n_604_port_15);
  spice_transistor_nmos_gnd g_4892(((~_DA_ADD1_v[`W-1]&~n_600_v[`W-1])|(~n_8_v[`W-1]&~n_1682_v[`W-1])), n_613_v, n_613_port_10);
  spice_transistor_nmos_gnd g_4891((~__AxB7__C67_v[`W-1]|(~_C67_v[`W-1]&~AxB7_v[`W-1])), __AxBxC_7_v, __AxBxC_7_port_5);
  spice_transistor_nmos_gnd g_4890((~_AxB_0__C0in_v[`W-1]|(~n_105_v[`W-1]&~__AxB_0_v[`W-1])), __AxBxC_0_v, __AxBxC_0_port_5);
  spice_transistor_nmos_gnd g_4899((~__AxB1__C01_v[`W-1]|(~AxB1_v[`W-1]&~_C01_v[`W-1])), __AxBxC_1_v, __AxBxC_1_port_5);
  spice_transistor_nmos_gnd g_4898(((~n_1595_v[`W-1]&pipeUNK13_v)|(~DBNeg_v[`W-1]&~n_754_v[`W-1])), n_1181_v, n_1181_port_6);
  spice_transistor_nmos t49(~dpc11_SBADD_v[`W-1], alua4_v, sb4_v, alua4_port_0, sb4_port_1);
  spice_transistor_nmos t48(~dpc11_SBADD_v[`W-1], alua3_v, sb3_v, alua3_port_0, sb3_port_0);
  spice_transistor_nmos_gnd t42(~pd0_clearIR_v[`W-1], n_409_v, n_409_port_0);
  spice_transistor_nmos t47(~dpc11_SBADD_v[`W-1], sb2_v, alua2_v, sb2_port_0, alua2_port_0);
  spice_transistor_nmos t46(~dpc11_SBADD_v[`W-1], sb1_v, alua1_v, sb1_port_0, alua1_port_2);
  spice_transistor_nmos t45(~cclk_v[`W-1], y1_v, n_767_v, y1_port_0, n_767_port_0);
  spice_transistor_nmos_gnd t44(notalu4_v, alu4_v, alu4_port_0);
  spice_transistor_nmos t3203(~dpc10_ADLADD_v[`W-1], adl6_v, alub6_v, adl6_port_6, alub6_port_4);
  spice_transistor_nmos t3206(~dpc10_ADLADD_v[`W-1], adl1_v, alub1_v, adl1_port_7, alub1_port_4);
  spice_transistor_nmos t3207(~dpc10_ADLADD_v[`W-1], adl4_v, alub4_v, adl4_port_6, alub4_port_4);
  spice_transistor_nmos t3204(~dpc10_ADLADD_v[`W-1], adl7_v, alub7_v, adl7_port_6, alub7_port_4);
  spice_transistor_nmos t3208(~dpc10_ADLADD_v[`W-1], alub5_v, adl5_v, alub5_port_4, adl5_port_5);
  spice_transistor_nmos t283(~dpc7_SS_v[`W-1], n_618_v, s6_v, n_618_port_1, s6_port_1);
  spice_transistor_nmos_gnd t280(n_101_v, n_1364_v, n_1364_port_0);
  spice_transistor_nmos t286(~dpc7_SS_v[`W-1], n_998_v, s3_v, n_998_port_1, s3_port_1);
  spice_transistor_nmos t287(~dpc7_SS_v[`W-1], n_1389_v, s2_v, n_1389_port_1, s2_port_1);
  spice_transistor_nmos t284(~dpc7_SS_v[`W-1], n_280_v, s5_v, n_280_port_0, s5_port_1);
  spice_transistor_nmos t285(~dpc7_SS_v[`W-1], n_3_v, s4_v, n_3_port_1, s4_port_1);
  spice_transistor_nmos t288(~dpc7_SS_v[`W-1], n_694_v, s1_v, n_694_port_0, s1_port_1);
  spice_transistor_nmos_gnd t289(~adh3_v[`W-1], n_883_v, n_883_port_1);
  spice_transistor_nmos t2009(~cclk_v[`W-1], n_541_v, notir7_v, n_541_port_1, notir7_port_34);
  spice_transistor_nmos_gnd t2008(~n_1067_v[`W-1], ADH_ABH_v, ADH_ABH_port_7);
  spice_transistor_nmos_gnd t2556(~dpc18__DAA_v[`W-1], n_700_v, n_700_port_1);
  spice_transistor_nmos t2551(~dpc32_PCHADH_v[`W-1], adh3_v, n_141_v, adh3_port_6, n_141_port_2);
  spice_transistor_nmos t2550(~dpc32_PCHADH_v[`W-1], adh4_v, n_27_v, adh4_port_6, n_27_port_2);
  spice_transistor_nmos t2553(~dpc32_PCHADH_v[`W-1], adh1_v, n_209_v, adh1_port_6, n_209_port_1);
  spice_transistor_nmos t2552(~dpc32_PCHADH_v[`W-1], adh2_v, n_1496_v, adh2_port_6, n_1496_port_2);
  spice_transistor_nmos_gnd t1217(~adl0_v[`W-1], n_123_v, n_123_port_0);
  spice_transistor_nmos t637(~cclk_v[`W-1], y2_v, n_1491_v, y2_port_0, n_1491_port_0);
  spice_transistor_nmos_gnd t1216(n_1272_v, n_608_v, n_608_port_0);
  spice_transistor_nmos t1208(~dpc20_ADDSB06_v[`W-1], alu6_v, sb6_v, alu6_port_2, sb6_port_6);
  spice_transistor_nmos t1209(~dpc20_ADDSB06_v[`W-1], alu5_v, sb5_v, alu5_port_1, sb5_port_3);
  spice_transistor_nmos_gnd t1201(n_1221_v, n_1566_v, n_1566_port_0);
  spice_transistor_nmos_gnd t2357(~n_659_v[`W-1], ab15_v, ab15_port_0);
  spice_transistor_nmos_vdd t2353(~n_298_v[`W-1], db7_v, db7_port_3);
  spice_transistor_nmos_gnd t1780(pipeUNK15_v, H1x1_v, H1x1_port_4);
  spice_transistor_nmos_vdd t3016(~n_1034_v[`W-1], n_994_v, n_994_port_3);
  spice_transistor_nmos_gnd t3015(~n_1034_v[`W-1], n_1545_v, n_1545_port_2);
  spice_transistor_nmos_gnd t3013(~n_717_v[`W-1], C1x5Reset_v, C1x5Reset_port_2);
  spice_transistor_nmos_gnd t1949(n_94_v, n_1024_v, n_1024_port_0);
  spice_transistor_nmos_gnd t1947(~n_849_v[`W-1], dpc33_PCHDB_v, dpc33_PCHDB_port_1);
  spice_transistor_nmos_gnd t1946(n_1411_v, pclp2_v, pclp2_port_1);
  spice_transistor_nmos_gnd t1945(~y3_v[`W-1], n_184_v, n_184_port_0);
  spice_transistor_nmos_gnd t1944(~op_T5_jsr_v[`W-1], n_1219_v, n_1219_port_1);
  spice_transistor_nmos_gnd t1943(n_1574_v, n_1089_v, n_1089_port_1);
  spice_transistor_nmos_gnd t1942(~clk0_v[`W-1], n_519_v, n_519_port_2);
  spice_transistor_nmos_gnd g_4685((~n_105_v[`W-1]|~__AxB_0_v[`W-1]), _AxB_0__C0in_v, _AxB_0__C0in_port_4);
  spice_transistor_nmos_vdd t2942(~n_617_v[`W-1], n_676_v, n_676_port_3);
  spice_transistor_nmos t2762(~cp1_v[`W-1], n_1661_v, idl3_v, n_1661_port_3, idl3_port_1);
  spice_transistor_nmos_vdd t2768(~n_1026_v[`W-1], n_171_v, n_171_port_3);
  spice_transistor_nmos_vdd t1410(~n_321_v[`W-1], dpc33_PCHDB_v, dpc33_PCHDB_port_0);
  spice_transistor_nmos_gnd g_4376((~notir2_v[`W-1]|~ir6_v[`W-1]|~irline3_v[`W-1]|~notir7_v[`W-1]|~ir5_v[`W-1]), op_sty_cpy_mem_v, op_sty_cpy_mem_port_8);
  spice_transistor_nmos_gnd g_4377((~op_T0_txs_v[`W-1]|~n_917_v[`W-1]|~n_1109_v[`W-1]), n_1358_v, n_1358_port_6);
  spice_transistor_nmos_gnd g_4374((~ir4_v[`W-1]|~notir6_v[`W-1]|~ir3_v[`W-1]|~ir7_v[`W-1]|~ir2_v[`W-1]|~notir5_v[`W-1]|~_t4_v[`W-1]|~irline3_v[`W-1]), op_T4_rts_v, op_T4_rts_port_11);
  spice_transistor_nmos_gnd g_4375((~notir3_v[`W-1]|~notir5_v[`W-1]|~irline3_v[`W-1]|~ir4_v[`W-1]|~ir2_v[`W-1]|~_t3_v[`W-1]|~ir7_v[`W-1]), op_T3_plp_pla_v, op_T3_plp_pla_port_10);
  spice_transistor_nmos_gnd g_4372((~ir2_v[`W-1]|~ir3_v[`W-1]|~ir4_v[`W-1]|~notir6_v[`W-1]|~_t5_v[`W-1]|~ir7_v[`W-1]|~irline3_v[`W-1]|~ir5_v[`W-1]), op_T5_rti_v, op_T5_rti_port_13);
  spice_transistor_nmos_gnd g_4373((~notir6_v[`W-1]|~notir2_v[`W-1]|~notir3_v[`W-1]|~ir7_v[`W-1]|~irline3_v[`W-1]|~ir4_v[`W-1]), op_jmp_v, op_jmp_port_8);
  spice_transistor_nmos_gnd g_4370((~irline3_v[`W-1]|~notir3_v[`W-1]|~ir7_v[`W-1]|~notir2_v[`W-1]|~notir6_v[`W-1]|~ir4_v[`W-1]|~_t4_v[`W-1]), op_T4_jmp_v, op_T4_jmp_port_11);
  spice_transistor_nmos_gnd g_4371((~n_572_v[`W-1]|~n_853_v[`W-1]), n_1517_v, n_1517_port_4);
  spice_transistor_nmos_gnd g_4378((~notir4_v[`W-1]|~ir2_v[`W-1]|~notir3_v[`W-1]|~clock1_v[`W-1]|~ir7_v[`W-1]|~ir6_v[`W-1]|~irline3_v[`W-1]), op_T0_clc_sec_v, op_T0_clc_sec_port_9);
  spice_transistor_nmos_gnd g_4379((~ir4_v[`W-1]|~notir5_v[`W-1]|~ir2_v[`W-1]|~ir7_v[`W-1]|~clock1_v[`W-1]|~irline3_v[`W-1]|~notir3_v[`W-1]|~ir6_v[`W-1]), op_T0_plp_v, op_T0_plp_port_10);
  spice_transistor_nmos_gnd g_4707((~DA_C01_v[`W-1]&~n_936_v[`W-1]), n_319_v, n_319_port_4);
  spice_transistor_nmos_gnd g_4701(((~n_1202_v[`W-1]|~n_200_v[`W-1])&~n_293_v[`W-1]), n_1402_v, n_1402_port_3);
  spice_transistor_nmos_gnd g_4700((~n_743_v[`W-1]&~n_1488_v[`W-1]), n_609_v, n_609_port_6);
  spice_transistor_nmos_gnd g_4709((~alub3_v[`W-1]&~alua3_v[`W-1]), n_350_v, n_350_port_5);
  spice_transistor_nmos_gnd g_4708((~n_1120_v[`W-1]&~n_440_v[`W-1]), n_504_v, n_504_port_3);
  spice_transistor_nmos_gnd t64(notalu6_v, alu6_v, alu6_port_0);
  spice_transistor_nmos_gnd t67(notidl2_v, idl2_v, idl2_port_0);
  spice_transistor_nmos_gnd t60(~pch3_v[`W-1], n_923_v, n_923_port_0);
  spice_transistor_nmos t3225(~dpc2_XSB_v[`W-1], n_1709_v, sb1_v, n_1709_port_2, sb1_port_12);
  spice_transistor_nmos_gnd t3226(~n_669_v[`W-1], op_ANDS_v, op_ANDS_port_5);
  spice_transistor_nmos t3489(~dpc13_ORS_v[`W-1], aluanorb1_v, notaluoutmux1_v, aluanorb1_port_4, notaluoutmux1_port_5);
  spice_transistor_nmos_gnd t3486(n_1395_v, Reset0_v, Reset0_port_4);
  spice_transistor_nmos_vdd t2572(~n_1639_v[`W-1], ab15_v, ab15_port_1);
  spice_transistor_nmos_vdd t2570(~n_1541_v[`W-1], dpc10_ADLADD_v, dpc10_ADLADD_port_5);
  spice_transistor_nmos_gnd t2577(pipeUNK29_v, n_1511_v, n_1511_port_1);
  spice_transistor_nmos t2683(~dpc9_DBADD_v[`W-1], alub7_v, idb7_v, alub7_port_0, idb7_port_8);
  spice_transistor_nmos_gnd t2682(~idb1_v[`W-1], n_243_v, n_243_port_1);
  spice_transistor_nmos t2684(~dpc9_DBADD_v[`W-1], alub6_v, idb6_v, alub6_port_2, idb6_port_10);
  spice_transistor_nmos_gnd t613(~clock1_v[`W-1], op_T0_v, op_T0_port_1);
  spice_transistor_nmos t1883(~cclk_v[`W-1], _ABL7_v, n_171_v, _ABL7_port_1, n_171_port_1);
  spice_transistor_nmos_vdd t1880(~n_1295_v[`W-1], dpc25_SBDB_v, dpc25_SBDB_port_9);
  spice_transistor_nmos_gnd t1886(n_799_v, n_1339_v, n_1339_port_1);
  spice_transistor_nmos_gnd t1887(~n_643_v[`W-1], db3_v, db3_port_3);
  spice_transistor_nmos_gnd t2642(~n_625_v[`W-1], n_662_v, n_662_port_0);
  spice_transistor_nmos_gnd t1082(~dpc12_0ADD_v[`W-1], alua6_v, alua6_port_1);
  spice_transistor_nmos_gnd t1083(~dpc12_0ADD_v[`W-1], alua5_v, alua5_port_1);
  spice_transistor_nmos_gnd t1080(~dpc12_0ADD_v[`W-1], alua1_v, alua1_port_3);
  spice_transistor_nmos_gnd t1081(~dpc12_0ADD_v[`W-1], alua4_v, alua4_port_1);
  spice_transistor_nmos_gnd t1086(~notalucin_v[`W-1], n_105_v, n_105_port_2);
  spice_transistor_nmos_gnd t1089(~n_37_v[`W-1], db2_v, db2_port_2);
  spice_transistor_nmos_vdd t1991(~n_23_v[`W-1], n_1501_v, n_1501_port_1);
  spice_transistor_nmos_gnd t1992(n_968_v, n_1093_v, n_1093_port_1);
  spice_transistor_nmos_gnd t1337(~idb3_v[`W-1], n_1600_v, n_1600_port_0);
  spice_transistor_nmos_vdd t1516(~abh0_v[`W-1], n_826_v, n_826_port_1);
  spice_transistor_nmos_gnd t1626(~db5_v[`W-1], n_1588_v, n_1588_port_1);
  spice_transistor_nmos_gnd t1628(~pd6_clearIR_v[`W-1], n_1309_v, n_1309_port_1);
  spice_transistor_nmos_gnd t1629(~_op_branch_bit7_v[`W-1], n_201_v, n_201_port_1);
  spice_transistor_nmos_gnd t189(n_408_v, aluvout_v, aluvout_port_0);
  spice_transistor_nmos_gnd t185(notidl6_v, idl6_v, idl6_port_0);
  spice_transistor_nmos_gnd g_4918(((pipeT4out_v&~notRdy0_v[`W-1])|(pipeT3out_v&~n_16_v[`W-1])), n_472_v, n_472_port_6);
  spice_transistor_nmos_gnd g_4919(((~__AxB_6_v[`W-1]&~C56_v[`W-1])|~_AxB_6__C56_v[`W-1]), __AxBxC_6_v, __AxBxC_6_port_5);
  spice_transistor_nmos_gnd g_4912(((n_1528_v&_TWOCYCLE_phi1_v)|n_1161_v), n_732_v, n_732_port_8);
  spice_transistor_nmos_gnd g_4913(((~n_1262_v[`W-1]&~n_236_v[`W-1])|(~n_646_v[`W-1]|~n_1655_v[`W-1]|~op_T5_rts_v[`W-1])), n_182_v, n_182_port_11);
  spice_transistor_nmos_gnd g_4910((~n_260_v[`W-1]|(~n_852_v[`W-1]&~n_1205_v[`W-1])), dasb7_v, dasb7_port_5);
  spice_transistor_nmos_gnd g_4911((~n_1316_v[`W-1]|(~n_344_v[`W-1]&~n_232_v[`W-1])), n_20_v, n_20_port_5);
  spice_transistor_nmos_gnd g_4916((~__AxB5__C45_v[`W-1]|(~AxB5_v[`W-1]&~_C45_v[`W-1])), __AxBxC_5_v, __AxBxC_5_port_5);
  spice_transistor_nmos_gnd g_4917((n_1673_v|(pipeUNK09_v&pipeUNK06_v)), n_754_v, n_754_port_8);
  spice_transistor_nmos_gnd g_4914((~n_975_v[`W-1]|(~n_312_v[`W-1]&~cclk_v[`W-1])), n_854_v, n_854_port_6);
  spice_transistor_nmos_gnd g_4915(((~op_from_x_v[`W-1]&~n_335_v[`W-1])|(~op_T0_cpx_inx_v[`W-1]|~op_T0_dex_v[`W-1]|~op_T0_txs_v[`W-1]|~x_op_T0_txa_v[`W-1]|~op_T2_ind_x_v[`W-1])|(~op_T2_idx_x_xy_v[`W-1]&~n_1244_v[`W-1])), n_1106_v, n_1106_port_12);
  spice_transistor_nmos_gnd t2748(n_698_v, VEC1_v, VEC1_port_3);
  spice_transistor_nmos t2218(~dpc15_ANDS_v[`W-1], n_336_v, n_722_v, n_336_port_3, n_722_port_5);
  spice_transistor_nmos t2219(~dpc15_ANDS_v[`W-1], n_304_v, n_1318_v, n_304_port_4, n_1318_port_3);
  spice_transistor_nmos t2216(~dpc15_ANDS_v[`W-1], n_1063_v, n_296_v, n_1063_port_4, n_296_port_4);
  spice_transistor_nmos t2217(~dpc15_ANDS_v[`W-1], n_277_v, n_477_v, n_277_port_4, n_477_port_3);
  spice_transistor_nmos t2214(~dpc15_ANDS_v[`W-1], n_681_v, n_740_v, n_681_port_3, n_740_port_4);
  spice_transistor_nmos t2747(~dpc37_PCLDB_v[`W-1], idb7_v, n_1647_v, idb7_port_9, n_1647_port_2);
  spice_transistor_nmos t2212(~dpc15_ANDS_v[`W-1], aluanandb0_v, notaluoutmux0_v, aluanandb0_port_3, notaluoutmux0_port_5);
  spice_transistor_nmos t2213(~dpc15_ANDS_v[`W-1], aluanandb1_v, notaluoutmux1_v, aluanandb1_port_1, notaluoutmux1_port_4);
  spice_transistor_nmos_gnd t2210(~C45_v[`W-1], _C45_v, _C45_port_1);
  spice_transistor_nmos_gnd g_4350((~n_1642_v[`W-1]|~n_440_v[`W-1]|~op_T2_php_pha_v[`W-1]|~op_T4_brk_v[`W-1]|~n_1258_v[`W-1]|~n_335_v[`W-1]), _WR_v, _WR_port_8);
  spice_transistor_nmos_gnd g_4351((~_t3_v[`W-1]|~notir4_v[`W-1]|~notir0_v[`W-1]|~ir3_v[`W-1]|~ir2_v[`W-1]), op_T3_ind_y_v, op_T3_ind_y_port_7);
  spice_transistor_nmos_gnd g_4352((~_t2_v[`W-1]|~notir3_v[`W-1]|~ir2_v[`W-1]|~notir0_v[`W-1]|~notir4_v[`W-1]), op_T2_abs_y_v, op_T2_abs_y_port_7);
  spice_transistor_nmos_gnd g_4353((~clock1_v[`W-1]|~notir4_v[`W-1]|~ir5_v[`W-1]|~ir2_v[`W-1]|~irline3_v[`W-1]|~ir6_v[`W-1]|~notir3_v[`W-1]|~notir7_v[`W-1]), x_op_T0_tya_v, x_op_T0_tya_port_10);
  spice_transistor_nmos_gnd g_4356((~notir1_v[`W-1]|~clock1_v[`W-1]|~ir2_v[`W-1]|~notir3_v[`W-1]|~notir4_v[`W-1]|~notir7_v[`W-1]|~ir6_v[`W-1]|~notir5_v[`W-1]), op_T0_tsx_v, op_T0_tsx_port_10);
  spice_transistor_nmos_gnd g_4357((~_t4_v[`W-1]|~ir3_v[`W-1]|~ir2_v[`W-1]|~notir4_v[`W-1]|~notir0_v[`W-1]), op_T4_ind_y_v, op_T4_ind_y_port_8);
  spice_transistor_nmos_gnd t404(~db3_v[`W-1], n_1281_v, n_1281_port_0);
  spice_transistor_nmos_gnd t405(~_C56_v[`W-1], C56_v, C56_port_0);
  spice_transistor_nmos_gnd g_4942((~dpc18__DAA_v[`W-1]|((~n_269_v[`W-1]|~n_570_v[`W-1])&(~n_757_v[`W-1]|~__AxB_6_v[`W-1]))), DC78_v, DC78_port_7);
  spice_transistor_nmos_gnd g_4763((~n_344_v[`W-1]&(~n_392_v[`W-1]|~n_410_v[`W-1])), n_1073_v, n_1073_port_3);
  spice_transistor_nmos_gnd g_4767((~n_844_v[`W-1]&~n_616_v[`W-1]), n_946_v, n_946_port_4);
  spice_transistor_nmos_gnd t2511(~idb3_v[`W-1], n_1621_v, n_1621_port_1);
  spice_transistor_nmos_gnd g_4291((~clearIR_v[`W-1]|pd2_v), pd2_clearIR_v, pd2_clearIR_port_7);
  spice_transistor_nmos_gnd g_4290((~notir1_v[`W-1]|~notir6_v[`W-1]|~notir5_v[`W-1]|~ir7_v[`W-1]), op_ror_v, op_ror_port_6);
  spice_transistor_nmos_gnd g_4292((~op_T4_rts_v[`W-1]|~op_T0_php_pha_v[`W-1]|~op_T5_rti_v[`W-1]|~op_T0_jsr_v[`W-1]|~op_T5_brk_v[`W-1]|~op_T3_plp_pla_v[`W-1]), n_1464_v, n_1464_port_8);
  spice_transistor_nmos_gnd g_4295((~n_1054_v[`W-1]|~_VEC_v[`W-1]), n_70_v, n_70_port_4);
  spice_transistor_nmos_gnd g_4297((~C1x5Reset_v[`W-1]|~_VEC_v[`W-1]|~n_264_v[`W-1]), n_1712_v, n_1712_port_5);
  spice_transistor_nmos_gnd g_4296((~x_op_T4_ind_y_v[`W-1]|~x_op_T3_abs_idx_v[`W-1]), n_261_v, n_261_port_4);
  spice_transistor_nmos_gnd g_4298((~op_T5_rts_v[`W-1]|~op_T5_ind_x_v[`W-1]|~op_T3_abs_idx_ind_v[`W-1]|~x_op_T4_ind_y_v[`W-1]), n_726_v, n_726_port_6);
  spice_transistor_nmos_gnd t896(~abh6_v[`W-1], n_635_v, n_635_port_1);
  spice_transistor_nmos_gnd t895(~abh6_v[`W-1], n_1523_v, n_1523_port_2);
  spice_transistor_nmos_vdd t894(~abh6_v[`W-1], n_963_v, n_963_port_2);
  spice_transistor_nmos_gnd t1608(~n_334_v[`W-1], Pout2_v, Pout2_port_1);
  spice_transistor_nmos t2554(~dpc32_PCHADH_v[`W-1], adh0_v, n_1722_v, adh0_port_6, n_1722_port_2);
  spice_transistor_nmos t2557(~cclk_v[`W-1], _ABH0_v, n_381_v, _ABH0_port_2, n_381_port_2);
  spice_transistor_nmos_vdd t2000(~n_1633_v[`W-1], ab5_v, ab5_port_1);
  spice_transistor_nmos_gnd g_4934((~dpc18__DAA_v[`W-1]|((~n_319_v[`W-1]|~n_1691_v[`W-1])&(~n_388_v[`W-1]|~n_1610_v[`W-1]))), DC34_v, DC34_port_9);
  spice_transistor_nmos_gnd g_4935(((~n_1257_v[`W-1]&~n_233_v[`W-1])|(~n_1018_v[`W-1]&~n_811_v[`W-1])), n_1205_v, n_1205_port_10);
  spice_transistor_nmos_gnd g_4936(((~n_986_v[`W-1]&~n_600_v[`W-1])|(~n_8_v[`W-1]&~n_876_v[`W-1])), n_345_v, n_345_port_10);
  spice_transistor_nmos_gnd g_4937(((~n_284_v[`W-1]&~cclk_v[`W-1])|~n_297_v[`W-1]), NMIP_v, NMIP_port_7);
  spice_transistor_nmos_gnd g_4930((~n_1213_v[`W-1]|(~n_609_v[`W-1]&~n_453_v[`W-1])), n_1209_v, n_1209_port_5);
  spice_transistor_nmos_gnd g_4931((pipeUNK40_v|(pipeUNK39_v&~notRdy0_v[`W-1])), n_1039_v, n_1039_port_5);
  spice_transistor_nmos_gnd g_4932((~_AxB_2__C12_v[`W-1]|(~__AxB_2_v[`W-1]&~C12_v[`W-1])), __AxBxC_2_v, __AxBxC_2_port_5);
  spice_transistor_nmos_gnd g_4933(((~op_T0_jsr_v[`W-1]&~n_1289_v[`W-1])|~op_T2_stack_v[`W-1]), n_632_v, n_632_port_5);
  spice_transistor_nmos_gnd g_4938(((~op_T0_shift_a_v[`W-1]|~op_T0_tax_v[`W-1]|~op_T0_tay_v[`W-1]|~op_ANDS_v[`W-1])|(~op_T0_acc_v[`W-1]&~n_397_v[`W-1])), n_11_v, n_11_port_9);
  spice_transistor_nmos_gnd g_4939((~n_404_v[`W-1]|(~n_1063_v[`W-1]&~_C34_v[`W-1])), C45_v, C45_port_7);
  spice_transistor_nmos_gnd t2234(n_756_v, n_1110_v, n_1110_port_1);
  spice_transistor_nmos t2235(~dpc26_ACDB_v[`W-1], n_146_v, idb0_v, n_146_port_1, idb0_port_8);
  spice_transistor_nmos t2236(~dpc26_ACDB_v[`W-1], n_929_v, idb1_v, n_929_port_2, idb1_port_5);
  spice_transistor_nmos t2237(~dpc26_ACDB_v[`W-1], n_1618_v, idb2_v, n_1618_port_0, idb2_port_6);
  spice_transistor_nmos_gnd t2231(~n_31_v[`W-1], n_132_v, n_132_port_1);
  spice_transistor_nmos t2238(~dpc26_ACDB_v[`W-1], n_1654_v, idb3_v, n_1654_port_2, idb3_port_6);
  spice_transistor_nmos t2239(~dpc26_ACDB_v[`W-1], idb4_v, n_1344_v, idb4_port_6, n_1344_port_0);
  spice_transistor_nmos t2728(~dpc9_DBADD_v[`W-1], alub5_v, idb5_v, alub5_port_2, idb5_port_8);
  spice_transistor_nmos t2729(~dpc9_DBADD_v[`W-1], alub4_v, idb4_v, alub4_port_3, idb4_port_8);
  spice_transistor_nmos t2726(~dpc9_DBADD_v[`W-1], alub3_v, idb3_v, alub3_port_3, idb3_port_8);
  spice_transistor_nmos t2727(~dpc9_DBADD_v[`W-1], idb2_v, alub2_v, idb2_port_9, alub2_port_4);
  spice_transistor_nmos t2724(~cp1_v[`W-1], n_1147_v, idl7_v, n_1147_port_3, idl7_port_1);
  spice_transistor_nmos t2725(~dpc9_DBADD_v[`W-1], alub1_v, idb1_v, alub1_port_1, idb1_port_7);
  spice_transistor_nmos_gnd t3348(~y5_v[`W-1], n_981_v, n_981_port_1);
  spice_transistor_nmos_gnd t429(~_ABH4_v[`W-1], abh4_v, abh4_port_0);
  spice_transistor_nmos_gnd t422(~n_135_v[`W-1], clk2out_v, clk2out_port_1);
  spice_transistor_nmos_gnd t421(~n_762_v[`W-1], n_1018_v, n_1018_port_0);
  spice_transistor_nmos_vdd t426(~cclk_v[`W-1], adh4_v, adh4_port_2);
  spice_transistor_nmos_vdd t427(~cclk_v[`W-1], adl5_v, adl5_port_0);
  spice_transistor_nmos_gnd g_4334((~n_71_v[`W-1]|~n_1247_v[`W-1]|~cclk_v[`W-1]), dpc7_SS_v, dpc7_SS_port_12);
  spice_transistor_nmos t3342(~cp1_v[`W-1], n_1095_v, idl4_v, n_1095_port_3, idl4_port_1);
  spice_transistor_nmos_gnd g_4741((~n_440_v[`W-1]&~op_shift_v[`W-1]), n_905_v, n_905_port_3);
  spice_transistor_nmos_gnd g_4747((~n_572_v[`W-1]&~n_1262_v[`W-1]), n_933_v, n_933_port_4);
  spice_transistor_nmos g_4746((~ADL_ABL_v[`W-1]&~cp1_v[`W-1]), _ABL0_v, n_123_v, _ABL0_port_3, n_123_port_3);
  spice_transistor_nmos_gnd g_4478((~_t4_v[`W-1]|~ir7_v[`W-1]|~ir6_v[`W-1]|~ir2_v[`W-1]|~ir4_v[`W-1]|~irline3_v[`W-1]|~ir3_v[`W-1]), op_T4_brk_jsr_v, op_T4_brk_jsr_port_9);
  spice_transistor_nmos_gnd g_4476((~notir2_v[`W-1]|~_t2_v[`W-1]|~ir4_v[`W-1]|~notir3_v[`W-1]), op_T2_abs_v, op_T2_abs_port_7);
  spice_transistor_nmos_gnd t228(n_621_v, n_355_v, n_355_port_0);
  spice_transistor_nmos_gnd t225(n_1061_v, pchp3_v, pchp3_port_0);
  spice_transistor_nmos t226(~dpc7_SS_v[`W-1], n_332_v, s0_v, n_332_port_0, s0_port_0);
  spice_transistor_nmos_vdd t227(~cclk_v[`W-1], idb0_v, idb0_port_1);
  spice_transistor_nmos_gnd t25(~abl0_v[`W-1], n_1100_v, n_1100_port_0);
  spice_transistor_nmos_vdd t27(~abl0_v[`W-1], n_855_v, n_855_port_0);
  spice_transistor_nmos_gnd t26(~abl0_v[`W-1], n_1660_v, n_1660_port_0);
  spice_transistor_nmos_gnd t2538(~idb6_v[`W-1], n_1416_v, n_1416_port_0);
  spice_transistor_nmos_gnd t2537(~n_0_ADL2_v[`W-1], adl2_v, adl2_port_6);
  spice_transistor_nmos t2535(~cclk_v[`W-1], n_635_v, _ABH6_v, n_635_port_3, _ABH6_port_2);
  spice_transistor_nmos t2532(~dpc38_PCLADL_v[`W-1], n_723_v, adl3_v, n_723_port_1, adl3_port_4);
  spice_transistor_nmos t2531(~dpc38_PCLADL_v[`W-1], adl2_v, n_481_v, adl2_port_5, n_481_port_2);
  spice_transistor_nmos t2530(~dpc38_PCLADL_v[`W-1], n_976_v, adl1_v, n_976_port_0, adl1_port_5);
  spice_transistor_nmos_gnd t2777(~n_842_v[`W-1], n_1479_v, n_1479_port_1);
  spice_transistor_nmos_gnd t2773(~n_404_v[`W-1], n_918_v, n_918_port_1);
  spice_transistor_nmos t1848(~dpc23_SBAC_v[`W-1], dasb7_v, a7_v, dasb7_port_1, a7_port_2);
  spice_transistor_nmos_gnd t1849(~n_251_v[`W-1], n_1028_v, n_1028_port_0);
  spice_transistor_nmos t1846(~dpc23_SBAC_v[`W-1], dasb5_v, a5_v, dasb5_port_1, a5_port_2);
  spice_transistor_nmos t1847(~dpc23_SBAC_v[`W-1], dasb6_v, a6_v, dasb6_port_0, a6_port_2);
  spice_transistor_nmos t1844(~dpc23_SBAC_v[`W-1], dasb3_v, a3_v, dasb3_port_1, a3_port_1);
  spice_transistor_nmos t1845(~dpc23_SBAC_v[`W-1], sb4_v, a4_v, sb4_port_7, a4_port_0);
  spice_transistor_nmos t1842(~dpc23_SBAC_v[`W-1], dasb1_v, a1_v, dasb1_port_0, a1_port_1);
  spice_transistor_nmos t1843(~dpc23_SBAC_v[`W-1], a2_v, dasb2_v, a2_port_1, dasb2_port_1);
  spice_transistor_nmos t1841(~dpc23_SBAC_v[`W-1], sb0_v, a0_v, sb0_port_5, a0_port_1);
  spice_transistor_nmos_gnd g_4484((~clock2_v[`W-1]|~ir7_v[`W-1]|~notir3_v[`W-1]|~ir6_v[`W-1]|~notir1_v[`W-1]|~ir2_v[`W-1]|~ir4_v[`W-1]), op_T__asl_rol_a_v, op_T__asl_rol_a_port_10);
  spice_transistor_nmos_gnd g_4485((~op_rti_rts_v[`W-1]|~brk_done_v[`W-1]|~x_op_T3_ind_y_v[`W-1]|~op_T2_jsr_v[`W-1]|~op_T4_ind_x_v[`W-1]|~n_389_v[`W-1]), n_300_v, n_300_port_8);
  spice_transistor_nmos_gnd g_4486((~n_201_v[`W-1]|~_op_branch_bit6_v[`W-1]|~n_90_v[`W-1]), n_1433_v, n_1433_port_6);
  spice_transistor_nmos_gnd g_4480((~op_ANDS_v[`W-1]|~n_384_v[`W-1]), n_550_v, n_550_port_5);
  spice_transistor_nmos_gnd g_4482((pd5_v|~clearIR_v[`W-1]), pd5_clearIR_v, pd5_clearIR_port_4);
  spice_transistor_nmos_gnd g_4483((~n_964_v[`W-1]|~n_732_v[`W-1]), clock1_v, clock1_port_68);
  spice_transistor_nmos_gnd g_4488((~n_1205_v[`W-1]|~n_852_v[`W-1]), n_260_v, n_260_port_4);
  spice_transistor_nmos_gnd g_4489((~n_769_v[`W-1]|~RnWstretched_v[`W-1]), n_1325_v, n_1325_port_4);
  spice_transistor_nmos_gnd t2437(~n_1696_v[`W-1], rw_v, rw_port_1);
  spice_transistor_nmos_gnd t2345(n_24_v, n_440_v, n_440_port_7);
  spice_transistor_nmos_gnd t326(n_1699_v, n_913_v, n_913_port_0);
  spice_transistor_nmos_gnd t2258(~pcl0_v[`W-1], n_937_v, n_937_port_0);
  spice_transistor_nmos_gnd t440(~n_400_v[`W-1], n_102_v, n_102_port_0);
  spice_transistor_nmos_vdd t441(~n_400_v[`W-1], n_1696_v, n_1696_port_0);
  spice_transistor_nmos_gnd t442(~n_834_v[`W-1], n_1696_v, n_1696_port_1);
  spice_transistor_nmos_gnd t443(~n_834_v[`W-1], n_400_v, n_400_port_2);
  spice_transistor_nmos_gnd t444(~x7_v[`W-1], n_1561_v, n_1561_port_0);
  spice_transistor_nmos_vdd t446(~n_1545_v[`W-1], ab10_v, ab10_port_0);
  spice_transistor_nmos_gnd g_4318((~notir3_v[`W-1]|~notir2_v[`W-1]|~notir6_v[`W-1]|~ir4_v[`W-1]|~irline3_v[`W-1]|~ir7_v[`W-1]), x_op_jmp_v, x_op_jmp_port_9);
  spice_transistor_nmos_gnd g_4319((~n_1024_v[`W-1]|n_1274_v), n_1069_v, n_1069_port_4);
  spice_transistor_nmos_vdd t2873(~n_1315_v[`W-1], n_381_v, n_381_port_3);
  spice_transistor_nmos_gnd t2871(notdor3_v, dor3_v, dor3_port_3);
  spice_transistor_nmos_gnd t1479(~op_T0_clc_sec_v[`W-1], n_889_v, n_889_port_1);
  spice_transistor_nmos_gnd t1478(~n_17_v[`W-1], n_646_v, n_646_port_2);
  spice_transistor_nmos_vdd t1477(~n_17_v[`W-1], clock1_v, clock1_port_40);
  spice_transistor_nmos_gnd t1474(~n_595_v[`W-1], n_992_v, n_992_port_0);
  spice_transistor_nmos_gnd t1470(~n_91_v[`W-1], n_1256_v, n_1256_port_0);
  spice_transistor_nmos_gnd t205(~n_999_v[`W-1], ab12_v, ab12_port_0);
  spice_transistor_nmos_vdd t3399(~n_1479_v[`W-1], ab1_v, ab1_port_1);
  spice_transistor_nmos_gnd t3427(~n_649_v[`W-1], A_B3_v, A_B3_port_1);
  spice_transistor_nmos t3391(~dpc6_SBS_v[`W-1], s7_v, sb7_v, s7_port_2, sb7_port_11);
  spice_transistor_nmos_gnd t3392(~n_642_v[`W-1], ab2_v, ab2_port_1);
  spice_transistor_nmos_gnd t3421(~aluanandb1_v[`W-1], n_936_v, n_936_port_4);
  spice_transistor_nmos_gnd t1864(~_C45_v[`W-1], DA_C45_v, DA_C45_port_1);
  spice_transistor_nmos_gnd t1865(~n_1194_v[`W-1], Pout3_v, Pout3_port_2);
  spice_transistor_nmos t1860(~dpc25_SBDB_v[`W-1], idb5_v, sb5_v, idb5_port_4, sb5_port_6);
  spice_transistor_nmos t1861(~dpc25_SBDB_v[`W-1], idb6_v, sb6_v, idb6_port_5, sb6_port_8);
  spice_transistor_nmos t1862(~dpc25_SBDB_v[`W-1], sb7_v, idb7_v, sb7_port_5, idb7_port_4);
  spice_transistor_nmos_gnd t1868(~VEC0_v[`W-1], n_728_v, n_728_port_0);
  spice_transistor_nmos_gnd t2654(~a0_v[`W-1], n_5_v, n_5_port_0);
  spice_transistor_nmos_gnd t1398(~op_T2_branch_v[`W-1], n_636_v, n_636_port_0);
  spice_transistor_nmos_gnd t1397(notalu1_v, alu1_v, alu1_port_1);
  spice_transistor_nmos_gnd t1395(n_675_v, n_888_v, n_888_port_0);
  spice_transistor_nmos t589(~dpc43_DL_DB_v[`W-1], idb4_v, n_1095_v, idb4_port_0, n_1095_port_1);
  spice_transistor_nmos_gnd t2110(~op_T0_cli_sei_v[`W-1], n_1065_v, n_1065_port_1);
  spice_transistor_nmos t587(~dpc43_DL_DB_v[`W-1], idb2_v, n_1424_v, idb2_port_1, n_1424_port_2);
  spice_transistor_nmos t586(~dpc43_DL_DB_v[`W-1], idb1_v, n_87_v, idb1_port_0, n_87_port_2);
  spice_transistor_nmos_gnd g_4468((~ir2_v[`W-1]|~ir4_v[`W-1]|~notir5_v[`W-1]|~ir7_v[`W-1]|~ir6_v[`W-1]|~irline3_v[`W-1]|~_t5_v[`W-1]|~ir3_v[`W-1]), op_T5_jsr_v, op_T5_jsr_port_10);
  spice_transistor_nmos_gnd g_4469((~_t2_v[`W-1]|~notir4_v[`W-1]|~notir0_v[`W-1]|~ir2_v[`W-1]|~ir3_v[`W-1]), op_T2_ind_y_v, op_T2_ind_y_port_8);
  spice_transistor_nmos_gnd g_4466((~_t3_v[`W-1]|~ir3_v[`W-1]|~notir4_v[`W-1]|~ir2_v[`W-1]|~notir0_v[`W-1]), x_op_T3_ind_y_v, x_op_T3_ind_y_port_7);
  spice_transistor_nmos_gnd g_4467((~_t2_v[`W-1]|~ir6_v[`W-1]|~ir2_v[`W-1]|~ir7_v[`W-1]|~notir5_v[`W-1]|~ir3_v[`W-1]|~irline3_v[`W-1]|~ir4_v[`W-1]), op_T2_jsr_v, op_T2_jsr_port_13);
  spice_transistor_nmos_gnd g_4464((n_1252_v|n_597_v), n_882_v, n_882_port_5);
  spice_transistor_nmos_gnd g_4465((~RnWstretched_v[`W-1]|~n_23_v[`W-1]), n_298_v, n_298_port_4);
  spice_transistor_nmos_gnd g_4462((~pd2_clearIR_v[`W-1]|~n_409_v[`W-1]|~pd4_clearIR_v[`W-1]|~n_1083_v[`W-1]), PD_xxx010x1_v, PD_xxx010x1_port_6);
  spice_transistor_nmos_gnd g_4463((~dpc22__DSA_v[`W-1]|~C34_v[`W-1]), n_1179_v, n_1179_port_4);
  spice_transistor_nmos_gnd g_4460((~n_641_v[`W-1]|~n_937_v[`W-1]|~dpc36_IPC_v[`W-1]|~n_783_v[`W-1]|~n_386_v[`W-1]|~n_1643_v[`W-1]|~n_232_v[`W-1]|~n_329_v[`W-1]|~n_249_v[`W-1]), dpc34_PCLC_v, dpc34_PCLC_port_14);
  spice_transistor_nmos_gnd g_4461((pipeUNK03_v|n_1177_v|~n_1111_v[`W-1]), n_1614_v, n_1614_port_5);
  spice_transistor_nmos t2278(~cclk_v[`W-1], n_927_v, notir4_v, n_927_port_1, notir4_port_24);
  spice_transistor_nmos_gnd t2279(~n_628_v[`W-1], n_1335_v, n_1335_port_0);
  spice_transistor_nmos_vdd t2270(~cclk_v[`W-1], idb5_v, idb5_port_6);
  spice_transistor_nmos_gnd t2274(~op_T3_branch_v[`W-1], n_1708_v, n_1708_port_3);
  spice_transistor_nmos_gnd t2276(~pclp4_v[`W-1], n_208_v, n_208_port_0);
  spice_transistor_nmos_vdd t466(~n_35_v[`W-1], dpc7_SS_v, dpc7_SS_port_7);
  spice_transistor_nmos_gnd t464(~n_378_v[`W-1], _t5_v, _t5_port_0);
  spice_transistor_nmos_gnd t465(~n_35_v[`W-1], n_71_v, n_71_port_0);
  spice_transistor_nmos_gnd t463(~a6_v[`W-1], n_1356_v, n_1356_port_0);
  spice_transistor_nmos_vdd t460(~abl3_v[`W-1], n_1041_v, n_1041_port_0);
  spice_transistor_nmos_gnd t461(pipeUNK11_v, n_1214_v, n_1214_port_0);
  spice_transistor_nmos_gnd t262(~op_T0_v[`W-1], n_638_v, n_638_port_0);
  spice_transistor_nmos_gnd t263(n_512_v, n_154_v, n_154_port_2);
  spice_transistor_nmos_gnd t265(~n_1427_v[`W-1], n_1448_v, n_1448_port_0);
  spice_transistor_nmos_gnd t266(n_223_v, n_1357_v, n_1357_port_0);
  spice_transistor_nmos_gnd t267(~n_1219_v[`W-1], n_1002_v, n_1002_port_1);
  spice_transistor_nmos t268(~H1x1_v[`W-1], idb0_v, Pout0_v, idb0_port_2, Pout0_port_0);
  spice_transistor_nmos_gnd g_4695((~fetch_v[`W-1]&~D1x1_v[`W-1]), clearIR_v, clearIR_port_18);
  spice_transistor_nmos g_4694((~ADL_ABL_v[`W-1]&~cp1_v[`W-1]), _ABL5_v, n_1094_v, _ABL5_port_3, n_1094_port_3);
  spice_transistor_nmos_gnd g_4697((~n_715_v[`W-1]&~n_1316_v[`W-1]), n_1386_v, n_1386_port_3);
  spice_transistor_nmos_gnd t1706(~ir1_v[`W-1], notir1_v, notir1_port_21);
  spice_transistor_nmos g_4690((~ADL_ABL_v[`W-1]&~cp1_v[`W-1]), _ABL6_v, n_1548_v, _ABL6_port_3, n_1548_port_3);
  spice_transistor_nmos g_4693((~ADL_ABL_v[`W-1]&~cp1_v[`W-1]), _ABL7_v, n_1046_v, _ABL7_port_3, n_1046_port_3);
  spice_transistor_nmos g_4692((~ADL_ABL_v[`W-1]&~cp1_v[`W-1]), _ABL4_v, n_1519_v, _ABL4_port_3, n_1519_port_3);
  spice_transistor_nmos_vdd t1701(~n_475_v[`W-1], ab12_v, ab12_port_1);
  spice_transistor_nmos_gnd t1700(~n_1708_v[`W-1], n_236_v, n_236_port_3);
  spice_transistor_nmos_gnd t1709(~n_1399_v[`W-1], n_1105_v, n_1105_port_2);
  spice_transistor_nmos_gnd t3404(~x3_v[`W-1], n_1521_v, n_1521_port_1);
  spice_transistor_nmos_gnd t3406(~n_355_v[`W-1], n_593_v, n_593_port_1);
  spice_transistor_nmos_vdd t3407(~n_355_v[`W-1], dpc4_SSB_v, dpc4_SSB_port_9);
  spice_transistor_nmos_gnd t1346(~y4_v[`W-1], n_565_v, n_565_port_0);
  spice_transistor_nmos_gnd t1806(~_t2_v[`W-1], op_T2_v, op_T2_port_0);
  spice_transistor_nmos_gnd t2827(~n_249_v[`W-1], n_163_v, n_163_port_2);
  spice_transistor_nmos_gnd t875(n_599_v, dpc22__DSA_v, dpc22__DSA_port_0);
  spice_transistor_nmos_vdd t877(~n_692_v[`W-1], dpc1_SBY_v, dpc1_SBY_port_3);
  spice_transistor_nmos_gnd t876(~n_692_v[`W-1], n_441_v, n_441_port_0);
  spice_transistor_nmos_vdd t870(~n_291_v[`W-1], dpc41_DL_ADL_v, dpc41_DL_ADL_port_0);
  spice_transistor_nmos_gnd t873(~n_278_v[`W-1], n_1488_v, n_1488_port_0);
  spice_transistor_nmos t2130(~H1x1_v[`W-1], p6_v, idb6_v, p6_port_0, idb6_port_6);
  spice_transistor_nmos_vdd t1118(~cclk_v[`W-1], sb3_v, sb3_port_3);
  spice_transistor_nmos t1110(~dpc17_SUMS_v[`W-1], __AxBxC_4_v, n_296_v, __AxBxC_4_port_2, n_296_port_1);
  spice_transistor_nmos t1111(~dpc17_SUMS_v[`W-1], __AxBxC_5_v, n_277_v, __AxBxC_5_port_1, n_277_port_2);
  spice_transistor_nmos t1112(~dpc17_SUMS_v[`W-1], n_722_v, __AxBxC_6_v, n_722_port_2, __AxBxC_6_port_1);
  spice_transistor_nmos t1113(~dpc17_SUMS_v[`W-1], n_304_v, __AxBxC_7_v, n_304_port_2, __AxBxC_7_port_0);
  spice_transistor_nmos_gnd g_4505((~DA_AxB2_v[`W-1]|~AxB1_v[`W-1]|~DA_C01_v[`W-1]|~n_936_v[`W-1]), n_388_v, n_388_port_6);
  spice_transistor_nmos_gnd g_4504((~n_862_v[`W-1]|~n_236_v[`W-1]|~n_646_v[`W-1]|~nnT2BR_v[`W-1]|~op_T2_abs_access_v[`W-1]|~op_T5_rts_v[`W-1]), n_272_v, n_272_port_9);
  spice_transistor_nmos_gnd g_4507((~n_1055_v[`W-1]|~op_T0_cmp_v[`W-1]|~op_T0_cpx_cpy_inx_iny_v[`W-1]), n_1560_v, n_1560_port_5);
  spice_transistor_nmos_gnd g_4506((~n_812_v[`W-1]|~n_31_v[`W-1]), n_1044_v, n_1044_port_4);
  spice_transistor_nmos_gnd g_4501((~cp1_v[`W-1]|~n_358_v[`W-1]), n_1129_v, n_1129_port_5);
  spice_transistor_nmos_gnd g_4500((~ir5_v[`W-1]|~notir3_v[`W-1]|~ir7_v[`W-1]|~irline3_v[`W-1]|~_t2_v[`W-1]|~notir6_v[`W-1]|~ir2_v[`W-1]|~ir4_v[`W-1]), op_T2_pha_v, op_T2_pha_port_10);
  spice_transistor_nmos_gnd g_4503((~notir3_v[`W-1]|~notir7_v[`W-1]|~notir6_v[`W-1]|~notir4_v[`W-1]|~irline3_v[`W-1]|~clock1_v[`W-1]|~ir2_v[`W-1]), op_T0_cld_sed_v, op_T0_cld_sed_port_9);
  spice_transistor_nmos_gnd g_4502((~n_1632_v[`W-1]|~n_647_v[`W-1]), AxB5_v, AxB5_port_7);
  spice_transistor_nmos_gnd g_4509((~n_739_v[`W-1]|~n_61_v[`W-1]), n_479_v, n_479_port_4);
  spice_transistor_nmos_gnd g_4508((~n_232_v[`W-1]|~n_344_v[`W-1]), n_1316_v, n_1316_port_7);
  spice_transistor_nmos_gnd t2011(n_666_v, n_862_v, n_862_port_4);
  spice_transistor_nmos_gnd t2012(~n_1323_v[`W-1], dpc37_PCLDB_v, dpc37_PCLDB_port_4);
  spice_transistor_nmos_gnd t2013(~pchp7_v[`W-1], n_1206_v, n_1206_port_0);
  spice_transistor_nmos t1507(~cclk_v[`W-1], n_146_v, a0_v, n_146_port_0, a0_port_0);
  spice_transistor_nmos_gnd t852(~ir7_v[`W-1], _op_branch_bit7_v, _op_branch_bit7_port_1);
  spice_transistor_nmos_gnd g_4440((~n_345_v[`W-1]|~n_432_v[`W-1]), n_1097_v, n_1097_port_4);
  spice_transistor_nmos_gnd g_4441((~n_790_v[`W-1]|~n_347_v[`W-1]|~notRdy0_v[`W-1]), n_191_v, n_191_port_5);
  spice_transistor_nmos_gnd g_4442((pipeUNK23_v|pipephi2Reset0_v), n_819_v, n_819_port_6);
  spice_transistor_nmos_gnd g_4443((~ir2_v[`W-1]|~notir6_v[`W-1]|~clock1_v[`W-1]|~ir4_v[`W-1]|~notir1_v[`W-1]|~notir3_v[`W-1]|~ir7_v[`W-1]), op_T0_shift_right_a_v, op_T0_shift_right_a_port_9);
  spice_transistor_nmos_gnd g_4444((~notir1_v[`W-1]|~notir6_v[`W-1]|~ir7_v[`W-1]), op_shift_right_v, op_shift_right_port_5);
  spice_transistor_nmos_gnd g_4445((~notir5_v[`W-1]|~notir1_v[`W-1]|~ir6_v[`W-1]|~ir7_v[`W-1]), op_rol_ror_v, op_rol_ror_port_7);
  spice_transistor_nmos_gnd g_4446((~notir1_v[`W-1]|~ir6_v[`W-1]|~ir7_v[`W-1]), op_shift_v, op_shift_port_5);
  spice_transistor_nmos_gnd g_4447((~clock2_v[`W-1]|~ir7_v[`W-1]|~ir2_v[`W-1]|~ir4_v[`W-1]|~notir1_v[`W-1]|~notir3_v[`W-1]), op_T__shift_a_v, op_T__shift_a_port_9);
  spice_transistor_nmos_gnd t1687(~op_xy_v[`W-1], n_1244_v, n_1244_port_1);
  spice_transistor_nmos_gnd t1503(pipeVectorA2_v, n_815_v, n_815_port_0);
  spice_transistor_nmos_gnd t1225(~n_384_v[`W-1], n_885_v, n_885_port_0);
  spice_transistor_nmos_gnd t3351(~adh7_v[`W-1], n_494_v, n_494_port_1);
  spice_transistor_nmos_gnd t3357(~n_184_v[`W-1], n_1531_v, n_1531_port_2);
  spice_transistor_nmos_gnd g_4448((~ir2_v[`W-1]|~notir3_v[`W-1]|~clock1_v[`W-1]|~ir5_v[`W-1]|~notir1_v[`W-1]|~ir6_v[`W-1]|~ir4_v[`W-1]|~notir7_v[`W-1]), op_T0_txa_v, op_T0_txa_port_11);
  spice_transistor_nmos_gnd g_4449((~pd0_clearIR_v[`W-1]|~n_1083_v[`W-1]|~pd2_clearIR_v[`W-1]), PD_xxxx10x0_v, PD_xxxx10x0_port_6);
  spice_transistor_nmos g_4818((~cp1_v[`W-1]&~ADH_ABH_v[`W-1]), n_1668_v, _ABH0_v, n_1668_port_3, _ABH0_port_3);
  spice_transistor_nmos_gnd t1566(~n_128_v[`W-1], n_1592_v, n_1592_port_1);
  spice_transistor_nmos_gnd t1561(~n_210_v[`W-1], ab5_v, ab5_port_0);
  spice_transistor_nmos t248(~dpc6_SBS_v[`W-1], s5_v, sb5_v, s5_port_0, sb5_port_1);
  spice_transistor_nmos t249(~dpc6_SBS_v[`W-1], s6_v, sb6_v, s6_port_0, sb6_port_3);
  spice_transistor_nmos t241(~cclk_v[`W-1], n_326_v, a6_v, n_326_port_0, a6_port_0);
  spice_transistor_nmos_gnd t2767(~n_1026_v[`W-1], n_322_v, n_322_port_2);
  spice_transistor_nmos_vdd t2764(~n_611_v[`W-1], dpc31_PCHPCH_v, dpc31_PCHPCH_port_11);
  spice_transistor_nmos_gnd t2763(~n_611_v[`W-1], n_255_v, n_255_port_1);
  spice_transistor_nmos_gnd t2760(~pd4_clearIR_v[`W-1], n_227_v, n_227_port_0);
  spice_transistor_nmos_gnd t3466(~D1x1_v[`W-1], n_1471_v, n_1471_port_1);
  spice_transistor_nmos_gnd t3467(~n_386_v[`W-1], n_392_v, n_392_port_2);
  spice_transistor_nmos_gnd t1828(~y7_v[`W-1], n_1640_v, n_1640_port_0);
  spice_transistor_nmos t1829(~cclk_v[`W-1], n_119_v, notir1_v, n_119_port_0, notir1_port_22);
  spice_transistor_nmos_gnd t1825(n_1679_v, n_1262_v, n_1262_port_2);
  spice_transistor_nmos t2482(~dpc31_PCHPCH_v[`W-1], pch1_v, n_209_v, pch1_port_2, n_209_port_0);
  spice_transistor_nmos t2481(~dpc31_PCHPCH_v[`W-1], pch0_v, n_1722_v, pch0_port_2, n_1722_port_1);
  spice_transistor_nmos t2480(~dpc31_PCHPCH_v[`W-1], pch3_v, n_141_v, pch3_port_2, n_141_port_1);
  spice_transistor_nmos_gnd t2487(~dpc29_0ADH17_v[`W-1], adh5_v, adh5_port_3);
  spice_transistor_nmos_gnd t2486(~dpc29_0ADH17_v[`W-1], adh2_v, adh2_port_5);
  spice_transistor_nmos_gnd t2485(~dpc29_0ADH17_v[`W-1], adh3_v, adh3_port_5);
  spice_transistor_nmos t2334(~dpc37_PCLDB_v[`W-1], idb4_v, n_208_v, idb4_port_7, n_208_port_1);
  spice_transistor_nmos_gnd t2488(~dpc29_0ADH17_v[`W-1], adh4_v, adh4_port_5);
  spice_transistor_nmos_gnd t2331(n_581_v, n_838_v, n_838_port_0);
  spice_transistor_nmos t1350(~cclk_v[`W-1], _ABL0_v, n_1100_v, _ABL0_port_2, n_1100_port_2);
  spice_transistor_nmos_vdd t2153(~n_1534_v[`W-1], dpc8_nDBADD_v, dpc8_nDBADD_port_6);
  spice_transistor_nmos_gnd t2152(~n_1534_v[`W-1], n_763_v, n_763_port_1);
  spice_transistor_nmos_gnd t2154(n_69_v, n_1045_v, n_1045_port_3);
  spice_transistor_nmos_vdd t2157(~n_417_v[`W-1], sync_v, sync_port_1);
  spice_transistor_nmos_gnd t1178(~a7_v[`W-1], n_128_v, n_128_port_0);
  spice_transistor_nmos_gnd t1176(~_ABL5_v[`W-1], abl5_v, abl5_port_0);
  spice_transistor_nmos_gnd g_4529((~dor0_v[`W-1]|~RnWstretched_v[`W-1]), n_1072_v, n_1072_port_4);
  spice_transistor_nmos_gnd g_4527((~ir5_v[`W-1]|~ir7_v[`W-1]|~ir6_v[`W-1]|~irline3_v[`W-1]|~ir4_v[`W-1]|~ir2_v[`W-1]|~ir3_v[`W-1]|~_t4_v[`W-1]), op_T4_brk_v, op_T4_brk_port_12);
  spice_transistor_nmos_gnd g_4526((~ir4_v[`W-1]|~ir7_v[`W-1]|~notir3_v[`W-1]|~irline3_v[`W-1]|~ir2_v[`W-1]), op_push_pull_v, op_push_pull_port_8);
  spice_transistor_nmos_gnd g_4525((~ir7_v[`W-1]|~notir3_v[`W-1]|~_t2_v[`W-1]|~ir5_v[`W-1]|~irline3_v[`W-1]|~ir2_v[`W-1]|~ir4_v[`W-1]), op_T2_php_pha_v, op_T2_php_pha_port_12);
  spice_transistor_nmos_gnd g_4524((~_t2_v[`W-1]|~irline3_v[`W-1]|~ir5_v[`W-1]|~ir2_v[`W-1]|~ir6_v[`W-1]|~ir4_v[`W-1]|~notir3_v[`W-1]|~ir7_v[`W-1]), op_T2_php_v, op_T2_php_port_10);
  spice_transistor_nmos_gnd g_4523((~_C45_v[`W-1]|~AxB5_v[`W-1]), __AxB5__C45_v, __AxB5__C45_port_4);
  spice_transistor_nmos_gnd g_4522((~n_218_v[`W-1]|~n_1258_v[`W-1]|~op_T3_branch_v[`W-1]|~n_510_v[`W-1]), n_1716_v, n_1716_port_6);
  spice_transistor_nmos_gnd g_4521((~_C23_v[`W-1]|~AxB3_v[`W-1]), __AxB3__C23_v, __AxB3__C23_port_4);
  spice_transistor_nmos_gnd g_4520((~n_604_v[`W-1]|~n_1377_v[`W-1]), n_385_v, n_385_port_4);
  spice_transistor_nmos_gnd g_4423((~RnWstretched_v[`W-1]|~dor4_v[`W-1]), n_1463_v, n_1463_port_5);
  spice_transistor_nmos_gnd g_4420((~n_781_v[`W-1]|~n_755_v[`W-1]), n_1170_v, n_1170_port_4);
  spice_transistor_nmos_gnd g_4421((~n_1214_v[`W-1]|~notRdy0_v[`W-1]), fetch_v, fetch_port_12);
  spice_transistor_nmos_gnd g_4426((~ir5_v[`W-1]|~notir6_v[`W-1]|~notir3_v[`W-1]|~notir7_v[`W-1]|~ir2_v[`W-1]|~notir1_v[`W-1]|~ir4_v[`W-1]|~clock1_v[`W-1]), op_T0_dex_v, op_T0_dex_port_11);
  spice_transistor_nmos_gnd g_4427((~_t2_v[`W-1]|~ir4_v[`W-1]|~ir3_v[`W-1]|~ir2_v[`W-1]|~notir0_v[`W-1]), op_T2_ind_x_v, op_T2_ind_x_port_8);
  spice_transistor_nmos_gnd g_4424((~RnWstretched_v[`W-1]|~dor4_v[`W-1]), n_147_v, n_147_port_4);
  spice_transistor_nmos_gnd g_4425((~ir5_v[`W-1]|~notir3_v[`W-1]|~clock2_v[`W-1]|~irline3_v[`W-1]|~ir4_v[`W-1]|~ir2_v[`W-1]|~notir7_v[`W-1]), op_T__iny_dey_v, op_T__iny_dey_port_9);
  spice_transistor_nmos_gnd g_4428((~ir2_v[`W-1]|~ir4_v[`W-1]|~notir3_v[`W-1]|~ir6_v[`W-1]|~clock1_v[`W-1]|~notir7_v[`W-1]|~ir5_v[`W-1]|~notir1_v[`W-1]), x_op_T0_txa_v, x_op_T0_txa_port_11);
  spice_transistor_nmos_gnd g_4429((~ir4_v[`W-1]|~irline3_v[`W-1]|~ir2_v[`W-1]|~notir3_v[`W-1]|~notir7_v[`W-1]|~ir5_v[`W-1]|~clock1_v[`W-1]), op_T0_iny_dey_v, op_T0_iny_dey_port_9);
  spice_transistor_nmos_gnd t1685(~n_476_v[`W-1], n_956_v, n_956_port_1);
  spice_transistor_nmos_vdd t1686(~n_476_v[`W-1], dpc12_0ADD_v, dpc12_0ADD_port_9);
  spice_transistor_nmos_gnd t1681(~s4_v[`W-1], n_973_v, n_973_port_1);
  spice_transistor_nmos_gnd t1682(~n_1471_v[`W-1], p4_v, p4_port_0);
  spice_transistor_nmos_gnd t1689(~idb5_v[`W-1], n_961_v, n_961_port_0);
  spice_transistor_nmos_vdd t382(~n_1076_v[`W-1], db4_v, db4_port_0);
  spice_transistor_nmos_gnd t386(~op_ror_v[`W-1], n_544_v, n_544_port_1);
  spice_transistor_nmos t385(~dpc4_SSB_v[`W-1], n_280_v, sb5_v, n_280_port_1, sb5_port_2);
  spice_transistor_nmos_gnd t3147(~abl4_v[`W-1], n_86_v, n_86_port_3);
  spice_transistor_nmos_gnd t3146(n_469_v, pchp5_v, pchp5_port_1);
  spice_transistor_nmos t3142(~dpc0_YSB_v[`W-1], n_767_v, sb1_v, n_767_port_2, sb1_port_11);
  spice_transistor_nmos_vdd t3149(~abl4_v[`W-1], n_634_v, n_634_port_1);
  spice_transistor_nmos_gnd t3148(~abl4_v[`W-1], n_1676_v, n_1676_port_2);
  spice_transistor_nmos_vdd t2818(~dor6_v[`W-1], n_7_v, n_7_port_2);
  spice_transistor_nmos_gnd t2819(~n_0_ADL0_v[`W-1], adl0_v, adl0_port_7);
  spice_transistor_nmos_gnd t1543(~n_1084_v[`W-1], n_803_v, n_803_port_0);
  spice_transistor_nmos_gnd t1540(~idb4_v[`W-1], n_797_v, n_797_port_1);
  spice_transistor_nmos_vdd t1548(~cclk_v[`W-1], sb7_v, sb7_port_3);
  spice_transistor_nmos_gnd t3448(~sb7_v[`W-1], n_852_v, n_852_port_2);
  spice_transistor_nmos_gnd t3336(~db7_v[`W-1], n_62_v, n_62_port_1);
  spice_transistor_nmos_gnd t3332(~pd1_clearIR_v[`W-1], n_1641_v, n_1641_port_1);
  spice_transistor_nmos_gnd t2667(~db6_v[`W-1], n_1638_v, n_1638_port_1);
  spice_transistor_nmos_gnd t2669(~n_206_v[`W-1], n_465_v, n_465_port_0);
  spice_transistor_nmos_gnd t2173(~_t4_v[`W-1], op_T4_v, op_T4_port_1);
  spice_transistor_nmos_gnd g_4549((~ir7_v[`W-1]|~irline3_v[`W-1]|~_t4_v[`W-1]|~ir2_v[`W-1]|~ir4_v[`W-1]|~ir5_v[`W-1]|~notir6_v[`W-1]|~ir3_v[`W-1]), x_op_T4_rti_v, x_op_T4_rti_port_10);
  spice_transistor_nmos_gnd g_4548((~_t2_v[`W-1]|~ir4_v[`W-1]|~notir2_v[`W-1]|~ir3_v[`W-1]), op_T2_mem_zp_v, op_T2_mem_zp_port_7);
  spice_transistor_nmos_gnd g_4541((~clock1_v[`W-1]|~ir6_v[`W-1]|~notir5_v[`W-1]|~notir7_v[`W-1]|~notir0_v[`W-1]), op_T0_lda_v, op_T0_lda_port_9);
  spice_transistor_nmos_gnd g_4540((~notir0_v[`W-1]|~clock1_v[`W-1]), op_T0_acc_v, op_T0_acc_port_4);
  spice_transistor_nmos_gnd g_4543((pipe_T0_v|~notRdy0_v[`W-1]), n_1180_v, n_1180_port_4);
  spice_transistor_nmos_gnd g_4545((~n_139_v[`W-1]|n_1624_v), n_169_v, n_169_port_4);
  spice_transistor_nmos_gnd g_4544((~n_225_v[`W-1]|~cclk_v[`W-1]|~n_1247_v[`W-1]), dpc9_DBADD_v, dpc9_DBADD_port_12);
  spice_transistor_nmos_gnd g_4547((~notir1_v[`W-1]|~notir3_v[`W-1]|~ir4_v[`W-1]|~ir2_v[`W-1]|~ir7_v[`W-1]|~clock1_v[`W-1]), op_T0_shift_a_v, op_T0_shift_a_port_11);
  spice_transistor_nmos_gnd g_4546((~ir6_v[`W-1]|~notir7_v[`W-1]|~ir4_v[`W-1]|~clock1_v[`W-1]|~notir5_v[`W-1]|~ir2_v[`W-1]|~irline3_v[`W-1]|~notir3_v[`W-1]), op_T0_tay_v, op_T0_tay_port_11);
  spice_transistor_nmos_gnd t1375(p1_v, n_318_v, n_318_port_1);
  spice_transistor_nmos_gnd t1372(n_1683_v, n_966_v, n_966_port_0);
  spice_transistor_nmos_gnd t1379(~pchp5_v[`W-1], n_1301_v, n_1301_port_0);
  spice_transistor_nmos_gnd g_4408((~ir6_v[`W-1]|~clock1_v[`W-1]|~irline3_v[`W-1]|~notir7_v[`W-1]|~ir4_v[`W-1]|~notir5_v[`W-1]), op_T0_tay_ldy_not_idx_v, op_T0_tay_ldy_not_idx_port_8);
  spice_transistor_nmos_gnd g_4409((~irline3_v[`W-1]|~notir7_v[`W-1]|~notir2_v[`W-1]|~notir5_v[`W-1]|~ir6_v[`W-1]|~clock1_v[`W-1]), op_T0_ldy_mem_v, op_T0_ldy_mem_port_8);
  spice_transistor_nmos_gnd g_4404((~_op_branch_bit7_v[`W-1]|~n_318_v[`W-1]|~_op_branch_bit6_v[`W-1]), n_1293_v, n_1293_port_6);
  spice_transistor_nmos_gnd g_4405((~n_236_v[`W-1]|~n_10_v[`W-1]), n_176_v, n_176_port_4);
  spice_transistor_nmos_gnd g_4406((~notir5_v[`W-1]|~irline3_v[`W-1]|~ir4_v[`W-1]|~ir6_v[`W-1]|~clock1_v[`W-1]|~ir3_v[`W-1]|~ir7_v[`W-1]|~ir2_v[`W-1]), op_T0_jsr_v, op_T0_jsr_port_12);
  spice_transistor_nmos_gnd g_4407((~ir2_v[`W-1]|~notir5_v[`W-1]|~clock2_v[`W-1]|~ir4_v[`W-1]|~irline3_v[`W-1]|~notir7_v[`W-1]|~notir6_v[`W-1]|~notir3_v[`W-1]), op_T__inx_v, op_T__inx_port_11);
  spice_transistor_nmos_gnd g_4400((~dor6_v[`W-1]|~RnWstretched_v[`W-1]), n_466_v, n_466_port_6);
  spice_transistor_nmos_gnd g_4401((~n_180_v[`W-1]|~n_819_v[`W-1]|~Reset0_v[`W-1]), n_501_v, n_501_port_5);
  spice_transistor_nmos_gnd g_4403((~op_T__dex_v[`W-1]|~op_T0_ldx_tax_tsx_v[`W-1]|~op_T__inx_v[`W-1]), n_844_v, n_844_port_6);
  spice_transistor_nmos_gnd t1388(notalu0_v, alu0_v, alu0_port_1);
  spice_transistor_nmos_gnd t199(n_982_v, n_1141_v, n_1141_port_1);
  spice_transistor_nmos_gnd t2780(n_1409_v, n_1231_v, n_1231_port_1);
  spice_transistor_nmos_gnd t2782(~sb5_v[`W-1], n_1135_v, n_1135_port_2);
  spice_transistor_nmos t2785(~cclk_v[`W-1], _ABL4_v, n_86_v, _ABL4_port_1, n_86_port_2);
  spice_transistor_nmos_gnd t2786(~n_70_v[`W-1], n_1117_v, n_1117_port_1);
  spice_transistor_nmos_gnd g_4398((~AxB1_v[`W-1]|~_C01_v[`W-1]), __AxB1__C01_v, __AxB1__C01_port_4);
  spice_transistor_nmos_gnd g_4399((~n_466_v[`W-1]|~RnWstretched_v[`W-1]), n_7_v, n_7_port_4);
  spice_transistor_nmos_gnd g_4394((~n_748_v[`W-1]|~n_1398_v[`W-1]), AxB7_v, AxB7_port_8);
  spice_transistor_nmos_gnd g_4395((~cclk_v[`W-1]|~n_491_v[`W-1]|~n_1247_v[`W-1]), dpc10_ADLADD_v, dpc10_ADLADD_port_12);
  spice_transistor_nmos_gnd g_4396((~ONEBYTE_v[`W-1]|pipeBRtaken_v|~notRdy0_v[`W-1]), n_1275_v, n_1275_port_5);
  spice_transistor_nmos_gnd g_4390((~n_347_v[`W-1]|~_op_store_v[`W-1]), n_335_v, n_335_port_10);
  spice_transistor_nmos_gnd g_4391((n_1162_v|~n_43_v[`W-1]), n_21_v, n_21_port_5);
  spice_transistor_nmos_gnd g_4392((~n_1449_v[`W-1]|n_759_v), n_944_v, n_944_port_4);
  spice_transistor_nmos_gnd g_4393((~n_544_v[`W-1]|n_785_v|~n_1175_v[`W-1]), n_267_v, n_267_port_5);
  spice_transistor_nmos_gnd t3163(~n_617_v[`W-1], n_1140_v, n_1140_port_2);
  spice_transistor_nmos_gnd t3161(~n_1398_v[`W-1], A_B7_v, A_B7_port_1);
  spice_transistor_nmos_gnd t3167(~x_op_T0_bit_v[`W-1], n_1379_v, n_1379_port_1);
  spice_transistor_nmos_gnd t3166(n_1625_v, n_90_v, n_90_port_3);
  spice_transistor_nmos_gnd t3164(n_1527_v, n_1295_v, n_1295_port_2);
  spice_transistor_nmos_gnd t994(~op_clv_v[`W-1], n_340_v, n_340_port_0);
  spice_transistor_nmos_gnd t992(~abh5_v[`W-1], n_869_v, n_869_port_1);
  spice_transistor_nmos t993(~dpc37_PCLDB_v[`W-1], idb2_v, n_481_v, idb2_port_3, n_481_port_1);
  spice_transistor_nmos_vdd t990(~abh5_v[`W-1], n_1608_v, n_1608_port_1);
  spice_transistor_nmos_gnd t991(~abh5_v[`W-1], n_1423_v, n_1423_port_0);
  spice_transistor_nmos_gnd t998(n_415_v, n_931_v, n_931_port_1);
  spice_transistor_nmos_gnd t999(n_88_v, n_1375_v, n_1375_port_0);
  spice_transistor_nmos t1529(~dpc3_SBX_v[`W-1], x5_v, sb5_v, x5_port_1, sb5_port_4);
  spice_transistor_nmos t1528(~dpc3_SBX_v[`W-1], sb6_v, x6_v, sb6_port_7, x6_port_1);
  spice_transistor_nmos_vdd t1521(~n_1677_v[`W-1], n_999_v, n_999_port_1);
  spice_transistor_nmos_gnd t1520(~n_1677_v[`W-1], n_475_v, n_475_port_0);
  spice_transistor_nmos t1525(~dpc3_SBX_v[`W-1], x2_v, sb2_v, x2_port_1, sb2_port_4);
  spice_transistor_nmos t1524(~dpc3_SBX_v[`W-1], x3_v, sb3_v, x3_port_1, sb3_port_6);
  spice_transistor_nmos_vdd t1527(~n_582_v[`W-1], ADH_ABH_v, ADH_ABH_port_4);
  spice_transistor_nmos_gnd t1526(~n_582_v[`W-1], n_1067_v, n_1067_port_0);
  spice_transistor_nmos_vdd t1344(~n_1715_v[`W-1], n_1105_v, n_1105_port_0);
  spice_transistor_nmos_gnd t1340(~alu6_v[`W-1], n_149_v, n_149_port_0);
  spice_transistor_nmos_gnd t3314(~s1_v[`W-1], n_1711_v, n_1711_port_1);
  spice_transistor_nmos t3316(~cclk_v[`W-1], y0_v, n_564_v, y0_port_2, n_564_port_2);
  spice_transistor_nmos t3317(~cclk_v[`W-1], n_659_v, _ABH7_v, n_659_port_3, _ABH7_port_2);
  spice_transistor_nmos_vdd t3313(~n_1463_v[`W-1], n_147_v, n_147_port_3);
  spice_transistor_nmos_vdd t176(~n_714_v[`W-1], dpc19_ADDSB7_v, dpc19_ADDSB7_port_0);
  spice_transistor_nmos t170(~cclk_v[`W-1], _ABL5_v, n_210_v, _ABL5_port_0, n_210_port_0);
  spice_transistor_nmos t2371(~dpc5_SADL_v[`W-1], adl1_v, n_694_v, adl1_port_4, n_694_port_3);
  spice_transistor_nmos t2370(~dpc24_ACSB_v[`W-1], n_1592_v, sb7_v, n_1592_port_3, sb7_port_9);
  spice_transistor_nmos_gnd t2373(pchp0_v, n_1722_v, n_1722_port_0);
  spice_transistor_nmos t2372(~cclk_v[`W-1], _ABL2_v, n_642_v, _ABL2_port_2, n_642_port_1);
  spice_transistor_nmos_gnd t505(pipeUNK21_v, n_572_v, n_572_port_0);
  spice_transistor_nmos_gnd t507(~n_1100_v[`W-1], ab0_v, ab0_port_0);
  spice_transistor_nmos_gnd t506(~sb6_v[`W-1], n_61_v, n_61_port_0);
  spice_transistor_nmos_gnd t501(~n_1676_v[`W-1], n_634_v, n_634_port_0);
  spice_transistor_nmos t503(~cclk_v[`W-1], notir0_v, n_310_v, notir0_port_1, n_310_port_0);
  spice_transistor_nmos_vdd t502(~n_1676_v[`W-1], n_86_v, n_86_port_0);
  spice_transistor_nmos t2199(~dpc27_SBADH_v[`W-1], adh2_v, sb2_v, adh2_port_4, sb2_port_8);
  spice_transistor_nmos t2198(~dpc27_SBADH_v[`W-1], adh3_v, sb3_v, adh3_port_3, sb3_port_9);
  spice_transistor_nmos_gnd t2195(~cp1_v[`W-1], n_1247_v, n_1247_port_13);
  spice_transistor_nmos_gnd t2194(~cp1_v[`W-1], n_38_v, n_38_port_1);
  spice_transistor_nmos t2191(~dpc27_SBADH_v[`W-1], sb6_v, adh6_v, sb6_port_9, adh6_port_3);
  spice_transistor_nmos t2190(~dpc27_SBADH_v[`W-1], adh7_v, sb7_v, adh7_port_3, sb7_port_7);
  spice_transistor_nmos t2193(~dpc27_SBADH_v[`W-1], adh0_v, sb0_v, adh0_port_2, sb0_port_9);
  spice_transistor_nmos t2192(~dpc1_SBY_v[`W-1], y0_v, sb0_v, y0_port_0, sb0_port_8);
  spice_transistor_nmos_gnd g_4563((~C12_v[`W-1]|~__AxB_2_v[`W-1]), _AxB_2__C12_v, _AxB_2__C12_port_4);
  spice_transistor_nmos_gnd g_4561((~n_453_v[`W-1]|~n_609_v[`W-1]), n_1213_v, n_1213_port_4);
  spice_transistor_nmos_gnd g_4560((n_1027_v|~n_43_v[`W-1]), n_476_v, n_476_port_5);
  spice_transistor_nmos_gnd g_4567((~AxB5_v[`W-1]|~DA_C45_v[`W-1]|~n_647_v[`W-1]|~n_122_v[`W-1]), n_570_v, n_570_port_6);
  spice_transistor_nmos_gnd g_4565((~irline3_v[`W-1]|~n_603_v[`W-1]|~ir2_v[`W-1]|~clock1_v[`W-1]|~ir3_v[`W-1]|~notir4_v[`W-1]), op_branch_done_v, op_branch_done_port_9);
  spice_transistor_nmos_gnd g_4564((~alub5_v[`W-1]|~alua5_v[`W-1]), n_1632_v, n_1632_port_7);
  spice_transistor_nmos_gnd g_4569((~n_440_v[`W-1]|~n_1258_v[`W-1]), n_813_v, n_813_port_4);
  spice_transistor_nmos_gnd g_4568((~n_992_v[`W-1]|~notRdy0_v[`W-1]), n_46_v, n_46_port_4);
  spice_transistor_nmos_gnd t1310(~idb1_v[`W-1], n_1474_v, n_1474_port_0);
  spice_transistor_nmos_gnd t1317(~so_v[`W-1], n_1650_v, n_1650_port_0);
  spice_transistor_nmos t1315(~cclk_v[`W-1], _ABL3_v, n_138_v, _ABL3_port_0, n_138_port_2);
  spice_transistor_nmos_gnd t1319(n_653_v, n_390_v, n_390_port_0);
  spice_transistor_nmos_gnd t1161(~n_236_v[`W-1], n_79_v, n_79_port_1);
  spice_transistor_nmos_gnd t1162(~C23_v[`W-1], _C23_v, _C23_port_2);
  spice_transistor_nmos t1165(~dpc8_nDBADD_v[`W-1], alub2_v, n_458_v, alub2_port_0, n_458_port_1);
  spice_transistor_nmos t1164(~dpc8_nDBADD_v[`W-1], alub4_v, n_478_v, alub4_port_0, n_478_port_0);
  spice_transistor_nmos_gnd t349(~ir0_v[`W-1], notir0_v, notir0_port_0);
  spice_transistor_nmos_gnd t347(~op_T3_jmp_v[`W-1], n_980_v, n_980_port_0);
  spice_transistor_nmos_vdd t345(~n_525_v[`W-1], dpc26_ACDB_v, dpc26_ACDB_port_0);
  spice_transistor_nmos_gnd t344(~n_525_v[`W-1], n_800_v, n_800_port_0);
  spice_transistor_nmos_gnd t343(~n_1305_v[`W-1], dpc17_SUMS_v, dpc17_SUMS_port_0);
  spice_transistor_nmos_gnd t340(n_1452_v, n_861_v, n_861_port_0);
  spice_transistor_nmos_gnd t2681(~a3_v[`W-1], n_947_v, n_947_port_1);
  spice_transistor_nmos_gnd g_4825((~alua7_v[`W-1]&~alub7_v[`W-1]), n_1318_v, n_1318_port_7);
  spice_transistor_nmos g_4822((~ADH_ABH_v[`W-1]&~cp1_v[`W-1]), _ABH2_v, n_168_v, _ABH2_port_3, n_168_port_3);
  spice_transistor_nmos_gnd g_4823((~n_681_v[`W-1]&~n_110_v[`W-1]), __AxB_2_v, __AxB_2_port_7);
  spice_transistor_nmos g_4820((~cp1_v[`W-1]&~fetch_v[`W-1]), n_227_v, n_927_v, n_227_port_3, n_927_port_3);
  spice_transistor_nmos_gnd g_4828((~n_813_v[`W-1]&~n_46_v[`W-1]), n_1101_v, n_1101_port_3);
  spice_transistor_nmos_gnd g_4829(((~n_83_v[`W-1]|~dpc35_PCHC_v[`W-1])&~n_523_v[`W-1]), n_1657_v, n_1657_port_3);
  spice_transistor_nmos_gnd t3103(~n_1254_v[`W-1], ab6_v, ab6_port_1);
  spice_transistor_nmos_gnd t3102(pipeUNK41_v, n_1497_v, n_1497_port_1);
  spice_transistor_nmos_gnd t978(~n_1585_v[`W-1], n_962_v, n_962_port_1);
  spice_transistor_nmos_gnd t974(~_ABL0_v[`W-1], abl0_v, abl0_port_3);
  spice_transistor_nmos t1508(~dpc0_YSB_v[`W-1], sb3_v, n_1531_v, sb3_port_5, n_1531_port_0);
  spice_transistor_nmos_gnd g_4619((~n_956_v[`W-1]|~cclk_v[`W-1]|~n_1247_v[`W-1]), dpc12_0ADD_v, dpc12_0ADD_port_12);
  spice_transistor_nmos_gnd g_4618((~n_1357_v[`W-1]|n_644_v), n_678_v, n_678_port_5);
  spice_transistor_nmos_gnd g_4615((~n_781_v[`W-1]|~n_1492_v[`W-1]), n_1457_v, n_1457_port_4);
  spice_transistor_nmos_gnd g_4614((~alub1_v[`W-1]|~alua1_v[`W-1]), aluanorb1_v, aluanorb1_port_7);
  spice_transistor_nmos_gnd g_4617((n_1606_v|~n_1357_v[`W-1]), n_188_v, n_188_port_5);
  spice_transistor_nmos_gnd g_4616((n_266_v|~cclk_v[`W-1]), n_525_v, n_525_port_5);
  spice_transistor_nmos_gnd g_4611((n_1360_v|~n_1357_v[`W-1]), n_1575_v, n_1575_port_5);
  spice_transistor_nmos_gnd g_4610((~n_1697_v[`W-1]|~n_773_v[`W-1]), n_275_v, n_275_port_4);
  spice_transistor_nmos_gnd g_4613((~n_1247_v[`W-1]|~cclk_v[`W-1]|~n_662_v[`W-1]), dpc3_SBX_v, dpc3_SBX_port_12);
  spice_transistor_nmos_gnd g_4612((~_t3_v[`W-1]|~ir4_v[`W-1]|~ir3_v[`W-1]|~ir2_v[`W-1]|~notir0_v[`W-1]), op_T3_ind_x_v, op_T3_ind_x_port_10);
  spice_transistor_nmos t3376(~dpc40_ADLPCL_v[`W-1], adl2_v, pcl2_v, adl2_port_8, pcl2_port_2);
  spice_transistor_nmos t3377(~dpc40_ADLPCL_v[`W-1], pcl5_v, adl5_v, pcl5_port_2, adl5_port_7);
  spice_transistor_nmos t3374(~dpc40_ADLPCL_v[`W-1], adl0_v, pcl0_v, adl0_port_8, pcl0_port_2);
  spice_transistor_nmos_gnd t2204(~y6_v[`W-1], n_1439_v, n_1439_port_1);
  spice_transistor_nmos t3378(~dpc40_ADLPCL_v[`W-1], adl4_v, pcl4_v, adl4_port_7, pcl4_port_2);
  spice_transistor_nmos t3379(~dpc40_ADLPCL_v[`W-1], adl6_v, pcl6_v, adl6_port_7, pcl6_port_2);
  spice_transistor_nmos_gnd t2759(~pcl2_v[`W-1], n_783_v, n_783_port_3);
  spice_transistor_nmos_gnd t153(~pch0_v[`W-1], n_1010_v, n_1010_port_0);
  spice_transistor_nmos_gnd t157(~_ABL7_v[`W-1], n_567_v, n_567_port_0);
  spice_transistor_nmos_vdd t154(~n_798_v[`W-1], db1_v, db1_port_1);
  spice_transistor_nmos_gnd t158(~adl6_v[`W-1], n_1548_v, n_1548_port_1);
  spice_transistor_nmos_gnd t1404(nots3_v, n_998_v, n_998_port_2);
  spice_transistor_nmos_gnd t1400(~db0_v[`W-1], n_93_v, n_93_port_0);
  spice_transistor_nmos_gnd t1401(~a2_v[`W-1], n_419_v, n_419_port_0);
  spice_transistor_nmos_gnd t2424(~n_1255_v[`W-1], dpc13_ORS_v, dpc13_ORS_port_5);
  spice_transistor_nmos_gnd t2427(n_897_v, n_1369_v, n_1369_port_2);
  spice_transistor_nmos_gnd t567(~__AxB_6_v[`W-1], n_122_v, n_122_port_0);
  spice_transistor_nmos_gnd t565(~n_664_v[`W-1], n_1697_v, n_1697_port_0);
  spice_transistor_nmos_gnd t569(~n_772_v[`W-1], n_1305_v, n_1305_port_1);
  spice_transistor_nmos_gnd g_4589((~cclk_v[`W-1]|~n_282_v[`W-1]|~n_1247_v[`W-1]), dpc6_SBS_v, dpc6_SBS_port_12);
  spice_transistor_nmos_gnd g_4588((~notir7_v[`W-1]|~ir5_v[`W-1]|~ir6_v[`W-1]), op_store_v, op_store_port_5);
  spice_transistor_nmos_gnd g_4585((~notir0_v[`W-1]|~notir5_v[`W-1]|~clock2_v[`W-1]|~notir6_v[`W-1]), x_op_T__adc_sbc_v, x_op_T__adc_sbc_port_8);
  spice_transistor_nmos_gnd g_4584((~alua4_v[`W-1]|~alub4_v[`W-1]), n_404_v, n_404_port_6);
  spice_transistor_nmos_gnd g_4587((~n_673_v[`W-1]|~op_T0_sbc_v[`W-1]), n_1304_v, n_1304_port_4);
  spice_transistor_nmos_gnd g_4586((n_1533_v|pipe_T0_v), n_964_v, n_964_port_7);
  spice_transistor_nmos_gnd g_4581((~notir7_v[`W-1]|~ir4_v[`W-1]|~irline3_v[`W-1]|~notir5_v[`W-1]|~clock1_v[`W-1]|~notir6_v[`W-1]), op_T0_cpx_inx_v, op_T0_cpx_inx_port_9);
  spice_transistor_nmos_gnd g_4580((~ir6_v[`W-1]|~notir5_v[`W-1]|~notir7_v[`W-1]|~notir1_v[`W-1]|~clock1_v[`W-1]), op_T0_ldx_tax_tsx_v, op_T0_ldx_tax_tsx_port_8);
  spice_transistor_nmos_gnd g_4583((~notir1_v[`W-1]|~ir6_v[`W-1]|~notir7_v[`W-1]), op_xy_v, op_xy_port_6);
  spice_transistor_nmos_gnd g_4582((~ir6_v[`W-1]|~ir5_v[`W-1]|~notir7_v[`W-1]|~notir1_v[`W-1]), op_from_x_v, op_from_x_port_7);
  spice_transistor_nmos_gnd t0(pipeVectorA0_v, n_0_ADL0_v, n_0_ADL0_port_0);
  spice_transistor_nmos t1338(~dpc3_SBX_v[`W-1], x1_v, sb1_v, x1_port_1, sb1_port_4);
  spice_transistor_nmos_gnd t1999(~n_1129_v[`W-1], n_1467_v, n_1467_port_1);
  spice_transistor_nmos t1331(~cclk_v[`W-1], n_831_v, a5_v, n_831_port_0, a5_port_0);
  spice_transistor_nmos_gnd t1996(~n_334_v[`W-1], n_118_v, n_118_port_1);
  spice_transistor_nmos t1333(~H1x1_v[`W-1], Pout1_v, idb1_v, Pout1_port_0, idb1_port_3);
  spice_transistor_nmos_gnd t1334(~n_172_v[`W-1], n_1633_v, n_1633_port_0);
  spice_transistor_nmos_vdd t1335(~n_172_v[`W-1], n_210_v, n_210_port_1);
  spice_transistor_nmos_gnd t1194(~_ABH3_v[`W-1], abh3_v, abh3_port_3);
  spice_transistor_nmos_gnd t1191(~_C34_v[`W-1], C34_v, C34_port_2);
  spice_transistor_nmos_vdd t367(~n_424_v[`W-1], notRdy0_v, notRdy0_port_3);
  spice_transistor_nmos_gnd t363(n_1333_v, n_906_v, n_906_port_0);
  spice_transistor_nmos_vdd t362(~n_1129_v[`W-1], cclk_v, cclk_port_28);
  spice_transistor_nmos_gnd t369(~n_198_v[`W-1], notRdy0_v, notRdy0_port_4);
  spice_transistor_nmos g_4802((~ADH_ABH_v[`W-1]&~cp1_v[`W-1]), _ABH5_v, n_254_v, _ABH5_port_3, n_254_port_3);
  spice_transistor_nmos_gnd g_4803((~n_462_v[`W-1]&~n_824_v[`W-1]), n_1642_v, n_1642_port_4);
  spice_transistor_nmos_gnd g_4805((~n_200_v[`W-1]&~n_1202_v[`W-1]), n_293_v, n_293_port_8);
  spice_transistor_nmos_gnd g_4807((~n_803_v[`W-1]&~n_336_v[`W-1]), __AxB_6_v, __AxB_6_port_11);
  spice_transistor_nmos_gnd g_4808((~alub0_v[`W-1]&~alua0_v[`W-1]), aluanandb0_v, aluanandb0_port_9);
  spice_transistor_nmos_gnd g_4809((~n_1542_v[`W-1]&(~n_1345_v[`W-1]|~n_1166_v[`W-1])), n_1099_v, n_1099_port_3);
  spice_transistor_nmos_gnd t3127(~n_1599_v[`W-1], n_538_v, n_538_port_1);
  spice_transistor_nmos_gnd t3125(~ir5_v[`W-1], notir5_v, notir5_port_36);
  spice_transistor_nmos_gnd t3123(~n_1719_v[`W-1], n_831_v, n_831_port_3);
  spice_transistor_nmos_vdd t3122(~n_224_v[`W-1], n_37_v, n_37_port_3);
  spice_transistor_nmos t3120(~dpc2_XSB_v[`W-1], n_436_v, sb4_v, n_436_port_2, sb4_port_12);
  spice_transistor_nmos_gnd t3129(~irq_v[`W-1], n_1599_v, n_1599_port_2);
  spice_transistor_nmos_gnd t2653(~n_1145_v[`W-1], op_ORS_v, op_ORS_port_2);
  spice_transistor_nmos_vdd t2651(~dor0_v[`W-1], n_1325_v, n_1325_port_2);
  spice_transistor_nmos_gnd t1078(~dpc12_0ADD_v[`W-1], alua0_v, alua0_port_1);
  spice_transistor_nmos_gnd t1627(~n_747_v[`W-1], n_1417_v, n_1417_port_2);
  spice_transistor_nmos t1621(~cclk_v[`W-1], n_1254_v, _ABL6_v, n_1254_port_1, _ABL6_port_1);
  spice_transistor_nmos_gnd g_4637((~n_645_v[`W-1]|~n_1374_v[`W-1]|~n_1578_v[`W-1]), n_1368_v, n_1368_port_5);
  spice_transistor_nmos_gnd g_4636((~n_440_v[`W-1]|~n_847_v[`W-1]|~nnT2BR_v[`W-1]|~op_T4_jmp_v[`W-1]|~n_275_v[`W-1]), n_104_v, n_104_port_7);
  spice_transistor_nmos_gnd g_4635((~notalucout_v[`W-1]|~n_1218_v[`W-1]), n_1257_v, n_1257_port_7);
  spice_transistor_nmos_gnd g_4634((~pd7_clearIR_v[`W-1]|~pd4_clearIR_v[`W-1]|~pd1_clearIR_v[`W-1]), PD_0xx0xx0x_v, PD_0xx0xx0x_port_5);
  spice_transistor_nmos_gnd g_4633((~n_771_v[`W-1]|~n_1708_v[`W-1]), n_1055_v, n_1055_port_5);
  spice_transistor_nmos_gnd g_4632((~n_1130_v[`W-1]|~n_267_v[`W-1]), n_80_v, n_80_port_4);
  spice_transistor_nmos_gnd g_4631((n_509_v|~n_43_v[`W-1]), n_1270_v, n_1270_port_5);
  spice_transistor_nmos_gnd g_4639((~n_708_v[`W-1]|~cclk_v[`W-1]|~n_1247_v[`W-1]), dpc11_SBADD_v, dpc11_SBADD_port_12);
  spice_transistor_nmos_gnd g_4638((~op_asl_rol_v[`W-1]|~op_lsr_ror_dec_inc_v[`W-1]), n_790_v, n_790_port_7);
  spice_transistor_nmos_gnd t3350(~n_310_v[`W-1], ir0_v, ir0_port_3);
  spice_transistor_nmos_vdd t3352(~cclk_v[`W-1], adh6_v, adh6_port_6);
  spice_transistor_nmos_vdd t3353(~cclk_v[`W-1], adl7_v, adl7_port_7);
  spice_transistor_nmos_gnd t3355(pclp1_v, n_976_v, n_976_port_3);
  spice_transistor_nmos_vdd t935(~n_1593_v[`W-1], dpc14_SRS_v, dpc14_SRS_port_1);
  spice_transistor_nmos_vdd t130(~n_1369_v[`W-1], dpc38_PCLADL_v, dpc38_PCLADL_port_0);
  spice_transistor_nmos t132(~dpc4_SSB_v[`W-1], n_721_v, sb7_v, n_721_port_0, sb7_port_0);
  spice_transistor_nmos t133(~dpc4_SSB_v[`W-1], n_618_v, sb6_v, n_618_port_0, sb6_port_2);
  spice_transistor_nmos_gnd t134(~n_818_v[`W-1], n_1043_v, n_1043_port_0);
  spice_transistor_nmos_vdd t135(~n_818_v[`W-1], dpc40_ADLPCL_v, dpc40_ADLPCL_port_0);
  spice_transistor_nmos t136(~dpc4_SSB_v[`W-1], n_3_v, sb4_v, n_3_port_0, sb4_port_3);
  spice_transistor_nmos_gnd t2890(~pchp1_v[`W-1], n_209_v, n_209_port_2);
  spice_transistor_nmos_gnd t2675(~abl5_v[`W-1], n_172_v, n_172_port_2);
  spice_transistor_nmos_vdd t2676(~abl5_v[`W-1], n_1633_v, n_1633_port_2);
  spice_transistor_nmos_gnd t540(~n_1635_v[`W-1], dpc29_0ADH17_v, dpc29_0ADH17_port_1);
  spice_transistor_nmos t546(~dpc13_ORS_v[`W-1], n_649_v, n_1071_v, n_649_port_0, n_1071_port_0);
  spice_transistor_nmos_vdd t1712(~n_1325_v[`W-1], db0_v, db0_port_1);
  spice_transistor_nmos_gnd t1718(~op_branch_done_v[`W-1], _op_branch_done_v, _op_branch_done_port_0);
  spice_transistor_nmos_gnd t301(~n_612_v[`W-1], db5_v, db5_port_0);
  spice_transistor_nmos_gnd t300(~n_730_v[`W-1], n_1724_v, n_1724_port_0);
  spice_transistor_nmos_gnd t309(~n_445_v[`W-1], n_417_v, n_417_port_0);
  spice_transistor_nmos_gnd t308(~n_445_v[`W-1], n_317_v, n_317_port_0);
  spice_transistor_nmos g_4790((~ADL_ABL_v[`W-1]&~cp1_v[`W-1]), _ABL2_v, n_935_v, _ABL2_port_3, n_935_port_3);
  spice_transistor_nmos_gnd g_4791((~n_918_v[`W-1]&~n_1063_v[`W-1]), __AxB_4_v, __AxB_4_port_6);
  spice_transistor_nmos_gnd g_4796((~Pout3_v[`W-1]&~op_T0_sbc_v[`W-1]), n_29_v, n_29_port_3);
  spice_transistor_nmos_gnd g_4798((~dpc35_PCHC_v[`W-1]&~n_83_v[`W-1]), n_523_v, n_523_port_6);
  spice_transistor_nmos_gnd g_4799((~alua2_v[`W-1]&~alub2_v[`W-1]), n_681_v, n_681_port_8);
  spice_transistor_nmos_gnd g_4868(((~n_523_v[`W-1]&~n_499_v[`W-1])|~n_743_v[`W-1]), n_875_v, n_875_port_5);
  spice_transistor_nmos_gnd g_4869((~n_936_v[`W-1]|(~C01_v[`W-1]&~A_B1_v[`W-1])), _C12_v, _C12_port_7);
  spice_transistor_nmos g_4862((~cp1_v[`W-1]&~fetch_v[`W-1]), n_1309_v, n_1675_v, n_1309_port_3, n_1675_port_3);
  spice_transistor_nmos g_4860((~cp1_v[`W-1]&~ADH_ABH_v[`W-1]), n_212_v, _ABH4_v, n_212_port_3, _ABH4_port_3);
  spice_transistor_nmos g_4861((~cp1_v[`W-1]&~fetch_v[`W-1]), n_928_v, n_1609_v, n_928_port_3, n_1609_port_3);
  spice_transistor_nmos_gnd g_4867((~aluanorb0_v[`W-1]|(~notalucin_v[`W-1]&~aluanandb0_v[`W-1])), DA_C01_v, DA_C01_port_8);
  spice_transistor_nmos g_4865((~cp1_v[`W-1]&~fetch_v[`W-1]), n_571_v, n_1300_v, n_571_port_3, n_1300_port_3);
  spice_transistor_nmos_gnd t2090(~n_981_v[`W-1], n_733_v, n_733_port_0);
  spice_transistor_nmos t2091(~cclk_v[`W-1], _ABL1_v, n_66_v, _ABL1_port_2, n_66_port_2);
  spice_transistor_nmos_vdd t2092(~abh4_v[`W-1], n_475_v, n_475_port_2);
  spice_transistor_nmos_gnd t2093(~abh4_v[`W-1], n_1677_v, n_1677_port_2);
  spice_transistor_nmos_gnd t2094(~abh4_v[`W-1], n_999_v, n_999_port_2);
  spice_transistor_nmos_gnd t2096(~C01_v[`W-1], _C01_v, _C01_port_2);
  spice_transistor_nmos_gnd t2098(n_1447_v, n_1175_v, n_1175_port_1);
  spice_transistor_nmos_gnd t2099(~_C78_v[`W-1], C78_v, C78_port_1);
  spice_transistor_nmos_gnd t1274(~n_1010_v[`W-1], n_311_v, n_311_port_2);
  spice_transistor_nmos t1273(~n_1446_v[`W-1], n_430_v, n_206_v, n_430_port_1, n_206_port_3);
  spice_transistor_nmos_gnd t932(~alu2_v[`W-1], _DA_ADD2_v, _DA_ADD2_port_2);
  spice_transistor_nmos_gnd t934(~n_1593_v[`W-1], n_1552_v, n_1552_port_0);
  spice_transistor_nmos_gnd t683(~pcl3_v[`W-1], n_249_v, n_249_port_0);
  spice_transistor_nmos t936(~dpc16_EORS_v[`W-1], __AxB_0_v, notaluoutmux0_v, __AxB_0_port_2, notaluoutmux0_port_0);
  spice_transistor_nmos t937(~dpc16_EORS_v[`W-1], notaluoutmux1_v, n_953_v, notaluoutmux1_port_0, n_953_port_0);
  spice_transistor_nmos t938(~dpc16_EORS_v[`W-1], __AxB_2_v, n_740_v, __AxB_2_port_0, n_740_port_1);
  spice_transistor_nmos t939(~dpc16_EORS_v[`W-1], n_884_v, n_1071_v, n_884_port_1, n_1071_port_2);
  spice_transistor_nmos_gnd t2678(~cp1_v[`W-1], n_43_v, n_43_port_13);
  spice_transistor_nmos_gnd t2674(~abl5_v[`W-1], n_210_v, n_210_port_3);
  spice_transistor_nmos_gnd t2892(~idb0_v[`W-1], n_1687_v, n_1687_port_1);
  spice_transistor_nmos_gnd t2677(~n_419_v[`W-1], n_1618_v, n_1618_port_2);
  spice_transistor_nmos_gnd t2894(~n_541_v[`W-1], ir7_v, ir7_port_59);
  spice_transistor_nmos t2895(~dpc20_ADDSB06_v[`W-1], alu1_v, sb1_v, alu1_port_3, sb1_port_10);
  spice_transistor_nmos_gnd t2896(pipeUNK12_v, n_587_v, n_587_port_1);
  spice_transistor_nmos t2897(~dpc20_ADDSB06_v[`W-1], alu0_v, sb0_v, alu0_port_2, sb0_port_11);
  spice_transistor_nmos_gnd t1011(~n_25_v[`W-1], n_674_v, n_674_port_0);
  spice_transistor_nmos t1010(~cclk_v[`W-1], n_1675_v, notir6_v, n_1675_port_0, notir6_port_1);
  spice_transistor_nmos t1015(~cclk_v[`W-1], n_929_v, a1_v, n_929_port_0, a1_port_0);
  spice_transistor_nmos_gnd t2339(nots0_v, n_332_v, n_332_port_2);
  spice_transistor_nmos_gnd g_4651((~_t2_v[`W-1]|~notir3_v[`W-1]|~op_push_pull_v[`W-1]), op_T2_abs_access_v, op_T2_abs_access_port_9);
  spice_transistor_nmos_gnd g_4650((~n_962_v[`W-1]|~cclk_v[`W-1]), _DBE_v, _DBE_port_5);
  spice_transistor_nmos_gnd g_4653((~n_8_v[`W-1]|~n_600_v[`W-1]), n_36_v, n_36_port_6);
  spice_transistor_nmos_gnd g_4652((~_t3_v[`W-1]|~notir3_v[`W-1]|~op_push_pull_v[`W-1]), op_T3_abs_idx_ind_v, op_T3_abs_idx_ind_port_6);
  spice_transistor_nmos_gnd g_4655((n_796_v|~n_43_v[`W-1]), n_35_v, n_35_port_5);
  spice_transistor_nmos_gnd g_4657((~n_1708_v[`W-1]|~n_770_v[`W-1]), n_19_v, n_19_port_4);
  spice_transistor_nmos_gnd g_4656((~op_T0_ora_v[`W-1]|~notRdy0_v[`W-1]), n_1145_v, n_1145_port_4);
  spice_transistor_nmos_gnd g_4659((~n_506_v[`W-1]|~n_933_v[`W-1]), n_877_v, n_877_port_5);
  spice_transistor_nmos_gnd g_4658((~RnWstretched_v[`W-1]|~dor0_v[`W-1]), n_769_v, n_769_port_6);
  spice_transistor_nmos_vdd t2336(~cclk_v[`W-1], adh3_v, adh3_port_4);
  spice_transistor_nmos_gnd t1352(~n_1380_v[`W-1], n_109_v, n_109_port_0);
  spice_transistor_nmos_gnd t115(notdor1_v, dor1_v, dor1_port_0);
  spice_transistor_nmos_gnd t112(~dpc12_0ADD_v[`W-1], alua3_v, alua3_port_1);
  spice_transistor_nmos_gnd t110(~abh3_v[`W-1], n_1346_v, n_1346_port_0);
  spice_transistor_nmos_gnd t111(~abh3_v[`W-1], n_359_v, n_359_port_0);
  spice_transistor_nmos_gnd t118(~_ABH7_v[`W-1], abh7_v, abh7_port_0);
  spice_transistor_nmos_gnd t2461(~AxB5_v[`W-1], n_1469_v, n_1469_port_1);
  spice_transistor_nmos_gnd t2462(~n_231_v[`W-1], ONEBYTE_v, ONEBYTE_port_1);
  spice_transistor_nmos_gnd t2467(~n_133_v[`W-1], n_602_v, n_602_port_0);
  spice_transistor_nmos_gnd t2466(~n_300_v[`W-1], n_847_v, n_847_port_1);
  spice_transistor_nmos_gnd t2469(~n_709_v[`W-1], dpc18__DAA_v, dpc18__DAA_port_2);
  spice_transistor_nmos_vdd t2468(~n_133_v[`W-1], dpc2_XSB_v, dpc2_XSB_port_2);
  spice_transistor_nmos_gnd t2565(~abl6_v[`W-1], n_1254_v, n_1254_port_2);
  spice_transistor_nmos_gnd t2566(~abl6_v[`W-1], n_1195_v, n_1195_port_2);
  spice_transistor_nmos_vdd t2567(~abl6_v[`W-1], n_1191_v, n_1191_port_2);
  spice_transistor_nmos_vdd t2560(~n_1041_v[`W-1], ab3_v, ab3_port_0);
  spice_transistor_nmos_vdd t2280(~n_628_v[`W-1], dpc24_ACSB_v, dpc24_ACSB_port_1);
  spice_transistor_nmos_gnd t331(n_1602_v, n_1596_v, n_1596_port_0);
  spice_transistor_nmos t1484(~dpc41_DL_ADL_v[`W-1], adl2_v, n_1424_v, adl2_port_2, n_1424_port_3);
  spice_transistor_nmos_vdd t1739(~cclk_v[`W-1], sb1_v, sb1_port_6);
  spice_transistor_nmos_gnd t1735(notidl7_v, idl7_v, idl7_port_0);
  spice_transistor_nmos t329(~dpc0_YSB_v[`W-1], n_564_v, sb0_v, n_564_port_0, sb0_port_1);
  spice_transistor_nmos t321(~dpc21_ADDADL_v[`W-1], alu2_v, adl2_v, alu2_port_0, adl2_port_0);
  spice_transistor_nmos t323(~dpc21_ADDADL_v[`W-1], adl0_v, alu0_v, adl0_port_0, alu0_port_0);
  spice_transistor_nmos t322(~dpc21_ADDADL_v[`W-1], adl1_v, alu1_v, adl1_port_0, alu1_port_0);
  spice_transistor_nmos_gnd g_4845((~n_1408_v[`W-1]&~n_980_v[`W-1]), n_473_v, n_473_port_3);
  spice_transistor_nmos g_4840((~cp1_v[`W-1]&~fetch_v[`W-1]), n_409_v, n_310_v, n_409_port_5, n_310_port_3);
  spice_transistor_nmos_gnd g_4843((~n_383_v[`W-1]&~n_1303_v[`W-1]), n_782_v, n_782_port_4);
  spice_transistor_nmos_gnd g_4849((n_1472_v&(n_1570_v|n_1581_v)), dpc36_IPC_v, dpc36_IPC_port_10);
  spice_transistor_nmos_gnd t2076(~abh0_v[`W-1], n_381_v, n_381_port_1);
  spice_transistor_nmos_gnd t2075(~abh0_v[`W-1], n_1315_v, n_1315_port_0);
  spice_transistor_nmos_gnd t1258(~n_1632_v[`W-1], A_B5_v, A_B5_port_1);
  spice_transistor_nmos_gnd t1253(~n_31_v[`W-1], Pout0_v, Pout0_port_1);
  spice_transistor_nmos_vdd t1254(~dor3_v[`W-1], n_42_v, n_42_port_0);
  spice_transistor_nmos_vdd t918(~n_1195_v[`W-1], n_1254_v, n_1254_port_0);
  spice_transistor_nmos_gnd t916(~n_726_v[`W-1], n_630_v, n_630_port_0);
  spice_transistor_nmos_gnd t917(~n_1195_v[`W-1], n_1191_v, n_1191_port_0);
  spice_transistor_nmos_gnd t914(nots7_v, n_721_v, n_721_port_2);
  spice_transistor_nmos_gnd t2618(notdor7_v, dor7_v, dor7_port_0);
  spice_transistor_nmos_gnd t2613(~n_1315_v[`W-1], n_826_v, n_826_port_2);
  spice_transistor_nmos_gnd t2611(~n_556_v[`W-1], n_1344_v, n_1344_port_2);
  spice_transistor_nmos t2616(~cclk_v[`W-1], n_733_v, y5_v, n_733_port_2, y5_port_1);
  spice_transistor_nmos_gnd t2614(~n_1265_v[`W-1], n_1202_v, n_1202_port_2);
  spice_transistor_nmos_vdd t1035(~n_358_v[`W-1], n_1467_v, n_1467_port_0);
  spice_transistor_nmos_gnd g_4679((~n_149_v[`W-1]|~n_761_v[`W-1]), n_762_v, n_762_port_4);
  spice_transistor_nmos_gnd g_4678((~n_499_v[`W-1]|~n_523_v[`W-1]), n_743_v, n_743_port_7);
  spice_transistor_nmos_gnd g_4673((~dor1_v[`W-1]|~RnWstretched_v[`W-1]), n_794_v, n_794_port_4);
  spice_transistor_nmos_gnd g_4672((~AxB7_v[`W-1]|~_C67_v[`W-1]), __AxB7__C67_v, __AxB7__C67_port_4);
  spice_transistor_nmos_gnd g_4671((~op_T4_brk_v[`W-1]|~op_T2_php_v[`W-1]), n_1391_v, n_1391_port_4);
  spice_transistor_nmos_gnd g_4670((~n_1070_v[`W-1]|~n_919_v[`W-1]), n_200_v, n_200_port_7);
  spice_transistor_nmos_gnd g_4677((~alua3_v[`W-1]|~alub3_v[`W-1]), n_649_v, n_649_port_7);
  spice_transistor_nmos_gnd g_4676((n_521_v|~n_43_v[`W-1]), n_6_v, n_6_port_5);
  spice_transistor_nmos_gnd g_4675((~alua6_v[`W-1]|~alub6_v[`W-1]), n_1084_v, n_1084_port_6);
  spice_transistor_nmos_gnd g_4674((~RnWstretched_v[`W-1]|~dor1_v[`W-1]), n_288_v, n_288_port_6);
  spice_transistor_nmos t2215(~dpc15_ANDS_v[`W-1], n_350_v, n_1071_v, n_350_port_3, n_1071_port_5);
  spice_transistor_nmos_gnd t2743(~n_519_v[`W-1], n_670_v, n_670_port_2);
  spice_transistor_nmos_gnd t2590(~_ABL4_v[`W-1], abl4_v, abl4_port_0);
  spice_transistor_nmos_gnd t2449(~n_754_v[`W-1], n_1595_v, n_1595_port_1);
  spice_transistor_nmos_gnd t2445(~op_SRS_v[`W-1], n_139_v, n_139_port_1);
  spice_transistor_nmos_gnd t2444(~op_store_v[`W-1], _op_store_v, _op_store_port_2);
  spice_transistor_nmos_gnd t2442(~dpc28_0ADH0_v[`W-1], adh0_v, adh0_port_3);
  spice_transistor_nmos_gnd t3066(~n_1462_v[`W-1], dpc38_PCLADL_v, dpc38_PCLADL_port_9);
  spice_transistor_nmos_gnd t3064(~adl2_v[`W-1], n_935_v, n_935_port_1);
  spice_transistor_nmos_gnd t3065(~n_5_v[`W-1], n_146_v, n_146_port_3);
  spice_transistor_nmos t2919(~cclk_v[`W-1], _ABH5_v, n_869_v, _ABH5_port_2, n_869_port_3);
  spice_transistor_nmos t2918(~dpc33_PCHDB_v[`W-1], idb7_v, n_1206_v, idb7_port_10, n_1206_port_3);
  spice_transistor_nmos t2915(~dpc33_PCHDB_v[`W-1], n_27_v, idb4_v, n_27_port_3, idb4_port_9);
  spice_transistor_nmos t2914(~dpc33_PCHDB_v[`W-1], n_141_v, idb3_v, n_141_port_3, idb3_port_10);
  spice_transistor_nmos t2917(~dpc33_PCHDB_v[`W-1], idb6_v, n_652_v, idb6_port_11, n_652_port_3);
  spice_transistor_nmos t2916(~dpc33_PCHDB_v[`W-1], n_1301_v, idb5_v, n_1301_port_3, idb5_port_9);
  spice_transistor_nmos t2911(~dpc33_PCHDB_v[`W-1], n_1722_v, idb0_v, n_1722_port_3, idb0_port_10);
  spice_transistor_nmos t2913(~dpc33_PCHDB_v[`W-1], idb2_v, n_1496_v, idb2_port_10, n_1496_port_3);
  spice_transistor_nmos t2912(~dpc33_PCHDB_v[`W-1], idb1_v, n_209_v, idb1_port_9, n_209_port_3);
  spice_transistor_nmos_gnd g_4354((~notir4_v[`W-1]|~_t2_v[`W-1]|~notir2_v[`W-1]), op_T2_idx_x_xy_v, op_T2_idx_x_xy_port_6);
  spice_transistor_nmos_gnd g_4355((~ir6_v[`W-1]|~ir2_v[`W-1]|~notir1_v[`W-1]|~ir5_v[`W-1]|~notir3_v[`W-1]|~notir4_v[`W-1]|~clock1_v[`W-1]|~notir7_v[`W-1]), op_T0_txs_v, op_T0_txs_port_12);
  spice_transistor_nmos_gnd t1939(~n_318_v[`W-1], Pout1_v, Pout1_port_1);
  spice_transistor_nmos_gnd t1937(~_ABH6_v[`W-1], abh6_v, abh6_port_3);
  spice_transistor_nmos_vdd t1934(~n_466_v[`W-1], n_471_v, n_471_port_3);
  spice_transistor_nmos_gnd g_4358((~op_T5_ind_x_v[`W-1]|~op_T0_jmp_v[`W-1]|~op_T5_rts_v[`W-1]|~op_T3_v[`W-1]|~op_T5_rti_v[`W-1]|~op_T4_v[`W-1]|~op_T0_brk_rti_v[`W-1]), n_256_v, n_256_port_9);
  spice_transistor_nmos_gnd g_4359((~n_838_v[`W-1]|~alucout_v[`W-1]), n_811_v, n_811_port_7);
  spice_transistor_nmos_gnd t495(~pd3_clearIR_v[`W-1], n_1083_v, n_1083_port_1);
  spice_transistor_nmos_gnd t492(~n_670_v[`W-1], n_747_v, n_747_port_0);
  spice_transistor_nmos_gnd t491(~adh6_v[`W-1], n_880_v, n_880_port_0);
  spice_transistor_nmos t490(~dpc7_SS_v[`W-1], s7_v, n_721_v, s7_port_0, n_721_port_1);
  spice_transistor_nmos t499(~dpc13_ORS_v[`W-1], n_722_v, n_1084_v, n_722_port_0, n_1084_port_0);
  spice_transistor_nmos t1752(~cp1_v[`W-1], n_1014_v, idl6_v, n_1014_port_3, idl6_port_1);
  spice_transistor_nmos_vdd t1750(~cclk_v[`W-1], adl2_v, adl2_port_4);
  spice_transistor_nmos_gnd t1756(n_1533_v, clock2_v, clock2_port_12);
  spice_transistor_nmos_vdd t1757(~n_373_v[`W-1], db5_v, db5_port_4);
  spice_transistor_nmos_gnd t1755(~n_905_v[`W-1], n_979_v, n_979_port_1);
  spice_transistor_nmos_gnd t92(~n_381_v[`W-1], ab8_v, ab8_port_1);
  spice_transistor_nmos t3181(~dpc27_SBADH_v[`W-1], adh5_v, sb5_v, adh5_port_5, sb5_port_11);
  spice_transistor_nmos t3180(~dpc39_PCLPCL_v[`W-1], pcl2_v, n_481_v, pcl2_port_1, n_481_port_3);
  spice_transistor_nmos_gnd t3183(~adh5_v[`W-1], n_254_v, n_254_port_1);
  spice_transistor_nmos t3182(~dpc5_SADL_v[`W-1], n_618_v, adl6_v, n_618_port_2, adl6_port_5);
  spice_transistor_nmos_gnd t3184(~n_336_v[`W-1], n_1038_v, n_1038_port_1);
  spice_transistor_nmos_gnd t3188(notidl1_v, idl1_v, idl1_port_1);
  spice_transistor_nmos_vdd t702(~abl2_v[`W-1], n_1152_v, n_1152_port_0);
  spice_transistor_nmos_gnd t701(~abl2_v[`W-1], n_951_v, n_951_port_0);
  spice_transistor_nmos_gnd t700(~abl2_v[`W-1], n_642_v, n_642_port_0);
  spice_transistor_nmos_gnd t709(~idb6_v[`W-1], n_351_v, n_351_port_0);
  spice_transistor_nmos_gnd t708(~AxB7_v[`W-1], n_177_v, n_177_port_0);
  spice_transistor_nmos_gnd t2588(~nmi_v[`W-1], n_1392_v, n_1392_port_2);
  spice_transistor_nmos_gnd t2583(pipeUNK22_v, n_533_v, n_533_port_1);
  spice_transistor_nmos_vdd t2586(~n_1423_v[`W-1], n_869_v, n_869_port_2);
  spice_transistor_nmos_gnd t2585(~n_1423_v[`W-1], n_1608_v, n_1608_port_2);
  spice_transistor_nmos_gnd t2635(~n_1157_v[`W-1], dpc41_DL_ADL_v, dpc41_DL_ADL_port_9);
  spice_transistor_nmos_gnd t2637(notdor5_v, dor5_v, dor5_port_3);
  spice_transistor_nmos t1615(~cclk_v[`W-1], n_436_v, x4_v, n_436_port_1, x4_port_1);
  spice_transistor_nmos_gnd t384(~pcl7_v[`W-1], n_641_v, n_641_port_0);
  spice_transistor_nmos_gnd t1619(~n_1045_v[`W-1], p7_v, p7_port_1);
  spice_transistor_nmos_gnd t1618(~db7_v[`W-1], n_588_v, n_588_port_0);
  spice_transistor_nmos_vdd t1587(~cclk_v[`W-1], sb0_v, sb0_port_4);
  spice_transistor_nmos_gnd t1580(pipedpc28_v, dpc28_0ADH0_v, dpc28_0ADH0_port_0);
  spice_transistor_nmos t924(~cclk_v[`W-1], n_359_v, _ABH3_v, n_359_port_1, _ABH3_port_1);
  spice_transistor_nmos_gnd t2658(~n_359_v[`W-1], ab11_v, ab11_port_1);
  spice_transistor_nmos_gnd t3450(~n_138_v[`W-1], ab3_v, ab3_port_1);
  spice_transistor_nmos_gnd t3049(n_993_v, pclp6_v, pclp6_port_0);
  spice_transistor_nmos_gnd t3046(~idb2_v[`W-1], n_1376_v, n_1376_port_1);
  spice_transistor_nmos_gnd t3047(~PD_0xx0xx0x_v[`W-1], PD_n_0xx0xx0x_v, PD_n_0xx0xx0x_port_0);
  spice_transistor_nmos_gnd t1917(n_663_v, pchp7_v, pchp7_port_0);
  spice_transistor_nmos_vdd t1911(~cclk_v[`W-1], adh2_v, adh2_port_3);
  spice_transistor_nmos_gnd t1919(~n_127_v[`W-1], n_135_v, n_135_port_2);
  spice_transistor_nmos_gnd t2119(~_ABH0_v[`W-1], abh0_v, abh0_port_3);
  spice_transistor_nmos_gnd t1773(~n_161_v[`W-1], n_969_v, n_969_port_0);
  spice_transistor_nmos_vdd t1774(~n_161_v[`W-1], dpc0_YSB_v, dpc0_YSB_port_3);
  spice_transistor_nmos_gnd t1775(~n_641_v[`W-1], n_715_v, n_715_port_2);
  spice_transistor_nmos t1779(~dpc1_SBY_v[`W-1], y5_v, sb5_v, y5_port_0, sb5_port_5);
  spice_transistor_nmos_gnd g_4738((~n_311_v[`W-1]&~dpc34_PCLC_v[`W-1]), n_919_v, n_919_port_6);
  spice_transistor_nmos_gnd g_4739((~_DA_ADD2_v[`W-1]&~_DA_ADD1_v[`W-1]), n_986_v, n_986_port_3);
  spice_transistor_nmos_gnd g_4732((~n_779_v[`W-1]&~n_604_v[`W-1]), n_1594_v, n_1594_port_3);
  spice_transistor_nmos_gnd g_4733((~n_1166_v[`W-1]&~n_1345_v[`W-1]), n_1542_v, n_1542_port_6);
  spice_transistor_nmos_gnd g_4731((~n_163_v[`W-1]&~n_1253_v[`W-1]), n_1184_v, n_1184_port_8);
  spice_transistor_nmos_gnd g_4888((~_AxB_4__C34_v[`W-1]|(~__AxB_4_v[`W-1]&~C34_v[`W-1])), __AxBxC_4_v, __AxBxC_4_port_5);
  spice_transistor_nmos_gnd g_4889(((~n_923_v[`W-1]&~n_293_v[`W-1])|~n_810_v[`W-1]), n_207_v, n_207_port_5);
  spice_transistor_nmos_gnd g_4880(((~op_from_x_v[`W-1]&~n_335_v[`W-1])|(~op_sty_cpy_mem_v[`W-1]&~n_335_v[`W-1])), n_1303_v, n_1303_port_7);
  spice_transistor_nmos_gnd g_4881(((~PD_n_0xx0xx0x_v[`W-1]&~PD_xxxx10x0_v[`W-1])|(~PD_xxx010x1_v[`W-1]|~PD_1xx000x0_v[`W-1])), _TWOCYCLE_v, _TWOCYCLE_port_7);
  spice_transistor_nmos_gnd g_4882((((~n_877_v[`W-1]|~n_1343_v[`W-1])&~n_79_v[`W-1])|~n_0_ADL0_v[`W-1]), n_696_v, n_696_port_5);
  spice_transistor_nmos_gnd g_4883((~n_1619_v[`W-1]|(~BRtaken_v[`W-1]&~nnT2BR_v[`W-1])), n_586_v, n_586_port_5);
  spice_transistor_nmos_gnd g_4884(((~_C56_v[`W-1]&~n_336_v[`W-1])|~n_1084_v[`W-1]), C67_v, C67_port_11);
  spice_transistor_nmos_gnd g_4885(((~notalucin_v[`W-1]&~aluanandb0_v[`W-1])|~aluanorb0_v[`W-1]), C01_v, C01_port_8);
  spice_transistor_nmos_gnd g_4886(((pipeUNK29_v&~n_1714_v[`W-1])|(~n_1511_v[`W-1]&pipeUNK28_v)), n_262_v, n_262_port_6);
  spice_transistor_nmos_gnd g_4887((~n_1159_v[`W-1]|(~n_1580_v[`W-1]&~n_613_v[`W-1])), dasb2_v, dasb2_port_5);
  spice_transistor_nmos t3210(~dpc10_ADLADD_v[`W-1], adl3_v, alub3_v, adl3_port_6, alub3_port_4);
  spice_transistor_nmos_gnd t3214(~db0_v[`W-1], n_718_v, n_718_port_1);
  spice_transistor_nmos_gnd t3217(~db2_v[`W-1], n_111_v, n_111_port_1);
  spice_transistor_nmos t3216(~cclk_v[`W-1], n_1618_v, a2_v, n_1618_port_3, a2_port_2);
  spice_transistor_nmos_gnd t3219(~db3_v[`W-1], n_896_v, n_896_port_1);
  spice_transistor_nmos t1485(~dpc41_DL_ADL_v[`W-1], adl0_v, n_719_v, adl0_port_3, n_719_port_3);
  spice_transistor_nmos t1482(~dpc41_DL_ADL_v[`W-1], adl4_v, n_1095_v, adl4_port_3, n_1095_port_2);
  spice_transistor_nmos t1483(~dpc41_DL_ADL_v[`W-1], adl1_v, n_87_v, adl1_port_2, n_87_port_3);
  spice_transistor_nmos t1481(~dpc41_DL_ADL_v[`W-1], adl3_v, n_1661_v, adl3_port_2, n_1661_port_2);
  spice_transistor_nmos_gnd t2033(~pd2_clearIR_v[`W-1], n_571_v, n_571_port_1);
  spice_transistor_nmos_gnd t2037(notidl4_v, idl4_v, idl4_port_0);
  spice_transistor_nmos t1211(~dpc20_ADDSB06_v[`W-1], alu3_v, sb3_v, alu3_port_1, sb3_port_4);
  spice_transistor_nmos t1210(~dpc20_ADDSB06_v[`W-1], sb4_v, alu4_v, sb4_port_5, alu4_port_2);
  spice_transistor_nmos_vdd t2326(~n_1566_v[`W-1], dpc43_DL_DB_v, dpc43_DL_DB_port_9);
  spice_transistor_nmos_gnd t2325(~n_1566_v[`W-1], n_1240_v, n_1240_port_1);
  spice_transistor_nmos_gnd t2490(~dpc29_0ADH17_v[`W-1], adh7_v, adh7_port_4);
  spice_transistor_nmos_gnd t2491(~dpc29_0ADH17_v[`W-1], adh6_v, adh6_port_4);
  spice_transistor_nmos t2320(~dpc37_PCLDB_v[`W-1], n_72_v, idb5_v, n_72_port_1, idb5_port_7);
  spice_transistor_nmos_gnd t1731(~pchp3_v[`W-1], n_141_v, n_141_port_0);
  spice_transistor_nmos_gnd g_4944(((~cclk_v[`W-1]&~n_538_v[`W-1])|~n_807_v[`W-1]), n_330_v, n_330_port_7);
  spice_transistor_nmos_gnd g_4946(((~n_862_v[`W-1]&~notRdy0_v[`W-1])|(((~nnT2BR_v[`W-1]&~BRtaken_v[`W-1])|~n_646_v[`W-1])&~n_372_v[`W-1])), n_1085_v, n_1085_port_6);
  spice_transistor_nmos_gnd g_4941(((~A_B5_v[`W-1]&~C45_v[`W-1])|~n_647_v[`W-1]), _C56_v, _C56_port_8);
  spice_transistor_nmos_gnd g_4940((~n_479_v[`W-1]|(~n_739_v[`W-1]&~n_61_v[`W-1])), dasb6_v, dasb6_port_5);
  spice_transistor_nmos_gnd g_4943((~__AxB3__C23_v[`W-1]|(~_C23_v[`W-1]&~AxB3_v[`W-1])), __AxBxC_3_v, __AxBxC_3_port_5);
  spice_transistor_nmos_gnd t2517(~_DA_ADD1_v[`W-1], n_1682_v, n_1682_port_1);
  spice_transistor_nmos_vdd t2516(~n_1613_v[`W-1], n_643_v, n_643_port_3);
  spice_transistor_nmos_gnd t791(notalu2_v, alu2_v, alu2_port_1);
  spice_transistor_nmos_gnd t3022(n_393_v, n_551_v, n_551_port_1);
  spice_transistor_nmos_gnd t3021(~adl1_v[`W-1], n_1016_v, n_1016_port_1);
  spice_transistor_nmos_gnd t1975(~n_119_v[`W-1], ir1_v, ir1_port_2);
  spice_transistor_nmos_gnd t1978(~n_188_v[`W-1], _t4_v, _t4_port_0);
  spice_transistor_nmos_vdd t2779(~abh1_v[`W-1], n_1140_v, n_1140_port_1);
  spice_transistor_nmos_vdd t2778(~n_842_v[`W-1], n_66_v, n_66_port_3);
  spice_transistor_nmos_gnd t1799(n_1565_v, n_1218_v, n_1218_port_1);
  spice_transistor_nmos_gnd t1797(~n_477_v[`W-1], n_647_v, n_647_port_3);
  spice_transistor_nmos_gnd t1792(~n_1501_v[`W-1], db7_v, db7_port_1);
  spice_transistor_nmos g_4711((~cp1_v[`W-1]&~fetch_v[`W-1]), n_1083_v, n_1620_v, n_1083_port_7, n_1620_port_3);
  spice_transistor_nmos g_4717((~ADH_ABH_v[`W-1]&~cp1_v[`W-1]), _ABH1_v, n_1267_v, _ABH1_port_3, n_1267_port_3);
  spice_transistor_nmos_gnd t52(~n_593_v[`W-1], dpc4_SSB_v, dpc4_SSB_port_0);
  spice_transistor_nmos t53(~dpc11_SBADD_v[`W-1], alua0_v, sb0_v, alua0_port_0, sb0_port_0);
  spice_transistor_nmos t55(~dpc11_SBADD_v[`W-1], alua5_v, sb5_v, alua5_port_0, sb5_port_0);
  spice_transistor_nmos t56(~dpc11_SBADD_v[`W-1], alua6_v, sb6_v, alua6_port_0, sb6_port_0);
  spice_transistor_nmos_gnd t57(~pch4_v[`W-1], n_1400_v, n_1400_port_0);
  spice_transistor_nmos_gnd t3237(~NMIP_v[`W-1], n_645_v, n_645_port_2);
  spice_transistor_nmos_gnd t3236(n_865_v, n_420_v, n_420_port_1);
  spice_transistor_nmos_gnd t3235(~n_1640_v[`W-1], n_1251_v, n_1251_port_2);
  spice_transistor_nmos_gnd t3234(~pch2_v[`W-1], n_1265_v, n_1265_port_2);
  spice_transistor_nmos t3233(~cclk_v[`W-1], a4_v, n_1344_v, a4_port_2, n_1344_port_3);
  spice_transistor_nmos_vdd t299(~cclk_v[`W-1], adh0_v, adh0_port_1);
  spice_transistor_nmos_gnd t295(~s6_v[`W-1], n_1187_v, n_1187_port_0);
  spice_transistor_nmos_gnd t297(~pd7_clearIR_v[`W-1], n_1605_v, n_1605_port_0);
  spice_transistor_nmos t296(~cp1_v[`W-1], n_719_v, idl0_v, n_719_port_1, idl0_port_0);
  spice_transistor_nmos_gnd t290(~_ABL6_v[`W-1], abl6_v, abl6_port_0);
  spice_transistor_nmos_gnd t293(~n_1413_v[`W-1], dpc32_PCHADH_v, dpc32_PCHADH_port_0);
  spice_transistor_nmos_vdd t3492(~n_6_v[`W-1], dpc6_SBS_v, dpc6_SBS_port_11);
  spice_transistor_nmos_gnd t3491(~n_6_v[`W-1], n_282_v, n_282_port_1);
  spice_transistor_nmos_gnd t3497(~n_678_v[`W-1], _t3_v, _t3_port_15);
  spice_transistor_nmos_gnd t3496(~x6_v[`W-1], n_730_v, n_730_port_1);
  spice_transistor_nmos_gnd t3495(~idb1_v[`W-1], n_583_v, n_583_port_1);
  spice_transistor_nmos_gnd t2018(~n_636_v[`W-1], nnT2BR_v, nnT2BR_port_5);
  spice_transistor_nmos_vdd t2019(~n_855_v[`W-1], ab0_v, ab0_port_1);
  spice_transistor_nmos t2548(~dpc32_PCHADH_v[`W-1], adh6_v, n_652_v, adh6_port_5, n_652_port_2);
  spice_transistor_nmos t2549(~dpc32_PCHADH_v[`W-1], adh5_v, n_1301_v, adh5_port_4, n_1301_port_2);
  spice_transistor_nmos t2547(~dpc32_PCHADH_v[`W-1], adh7_v, n_1206_v, adh7_port_5, n_1206_port_2);
  spice_transistor_nmos_vdd t2544(~n_839_v[`W-1], n_43_v, n_43_port_11);
  spice_transistor_nmos_gnd t2543(~adl3_v[`W-1], n_1507_v, n_1507_port_1);
  spice_transistor_nmos_gnd t2016(~idb7_v[`W-1], DBNeg_v, DBNeg_port_1);
  spice_transistor_nmos_gnd t2541(~n_1400_v[`W-1], n_83_v, n_83_port_0);
  spice_transistor_nmos_vdd t1894(~n_102_v[`W-1], rw_v, rw_port_0);
  spice_transistor_nmos_gnd t103(~y1_v[`W-1], n_1138_v, n_1138_port_0);
  spice_transistor_nmos t2733(~cclk_v[`W-1], _ABH2_v, n_994_v, _ABH2_port_2, n_994_port_2);
  spice_transistor_nmos_vdd t2227(~n_1499_v[`W-1], dpc18__DAA_v, dpc18__DAA_port_1);
  spice_transistor_nmos_vdd t196(~n_1720_v[`W-1], n_612_v, n_612_port_0);
  spice_transistor_nmos_vdd t197(~dor4_v[`W-1], n_1076_v, n_1076_port_0);
  spice_transistor_nmos_gnd t192(~pch7_v[`W-1], n_453_v, n_453_port_1);
  spice_transistor_nmos_gnd t190(~ir3_v[`W-1], notir3_v, notir3_port_0);
  spice_transistor_nmos t191(~cclk_v[`W-1], n_1609_v, notir5_v, n_1609_port_0, notir5_port_0);
  spice_transistor_nmos_gnd t3009(~n_312_v[`W-1], n_995_v, n_995_port_1);
  spice_transistor_nmos t1958(~dpc13_ORS_v[`W-1], aluanorb0_v, notaluoutmux0_v, aluanorb0_port_1, notaluoutmux0_port_3);
  spice_transistor_nmos_gnd t1959(~n_947_v[`W-1], n_1654_v, n_1654_port_1);
  spice_transistor_nmos_gnd t1955(~n_1230_v[`W-1], n_708_v, n_708_port_1);
  spice_transistor_nmos_vdd t1956(~n_1230_v[`W-1], dpc11_SBADD_v, dpc11_SBADD_port_9);
  spice_transistor_nmos t1957(~dpc13_ORS_v[`W-1], n_304_v, n_1398_v, n_304_port_3, n_1398_port_1);
  spice_transistor_nmos_gnd g_4349((~op_SRS_v[`W-1]|~n_781_v[`W-1]), n_160_v, n_160_port_4);
  spice_transistor_nmos_gnd g_4348((~op_T5_rti_rts_v[`W-1]|~op_T2_php_pha_v[`W-1]|~xx_op_T5_jsr_v[`W-1]|~x_op_T3_plp_pla_v[`W-1]|~op_T4_jmp_v[`W-1]|~op_T2_jmp_abs_v[`W-1]), n_368_v, n_368_port_8);
  spice_transistor_nmos_gnd g_4347((~_t4_v[`W-1]|~ir3_v[`W-1]|~notir4_v[`W-1]|~notir0_v[`W-1]|~ir2_v[`W-1]), x_op_T4_ind_y_v, x_op_T4_ind_y_port_10);
  spice_transistor_nmos_gnd g_4346((~ir3_v[`W-1]|~_t5_v[`W-1]|~notir0_v[`W-1]|~ir2_v[`W-1]|~ir4_v[`W-1]), op_T5_ind_x_v, op_T5_ind_x_port_9);
  spice_transistor_nmos_gnd g_4345((~_t2_v[`W-1]|~ir3_v[`W-1]|~ir2_v[`W-1]|~notir0_v[`W-1]), op_T2_ind_v, op_T2_ind_port_6);
  spice_transistor_nmos_gnd g_4344((~short_circuit_idx_add_v[`W-1]|~brk_done_v[`W-1]|~n_238_v[`W-1]), n_1215_v, n_1215_port_6);
  spice_transistor_nmos_gnd g_4341((~n_1109_v[`W-1]|~n_1002_v[`W-1]|~n_192_v[`W-1]|~n_1258_v[`W-1]|~n_862_v[`W-1]), n_1130_v, n_1130_port_8);
  spice_transistor_nmos_gnd g_4340((~RnWstretched_v[`W-1]|~dor2_v[`W-1]), n_37_v, n_37_port_4);
  spice_transistor_nmos_vdd t2752(~n_21_v[`W-1], dpc30_ADHPCH_v, dpc30_ADHPCH_port_10);
  spice_transistor_nmos_gnd t2751(~n_21_v[`W-1], n_228_v, n_228_port_0);
  spice_transistor_nmos_gnd t2209(~n_75_v[`W-1], dpc20_ADDSB06_v, dpc20_ADDSB06_port_5);
  spice_transistor_nmos_vdd t2208(~n_834_v[`W-1], n_102_v, n_102_port_2);
  spice_transistor_nmos_gnd t2754(notalu7_v, alu7_v, alu7_port_2);
  spice_transistor_nmos_gnd t1408(nots1_v, n_694_v, n_694_port_2);
  spice_transistor_nmos_gnd t1409(~n_321_v[`W-1], n_849_v, n_849_port_0);
  spice_transistor_nmos_gnd t1402(~ir7_v[`W-1], notir7_v, notir7_port_33);
  spice_transistor_nmos_gnd t1403(~n_1304_v[`W-1], n_1688_v, n_1688_port_0);
  spice_transistor_nmos_gnd g_4365((~ir7_v[`W-1]|~_t2_v[`W-1]|~ir4_v[`W-1]|~notir3_v[`W-1]|~notir2_v[`W-1]|~ir5_v[`W-1]|~irline3_v[`W-1]|~notir6_v[`W-1]), op_T2_jmp_abs_v, op_T2_jmp_abs_port_11);
  spice_transistor_nmos_gnd g_4364((~_t3_v[`W-1]|~notir3_v[`W-1]|~ir4_v[`W-1]|~notir2_v[`W-1]), op_T3_mem_abs_v, op_T3_mem_abs_port_7);
  spice_transistor_nmos_gnd g_4367((~_t3_v[`W-1]|~notir2_v[`W-1]|~ir3_v[`W-1]|~notir4_v[`W-1]), op_T3_mem_zp_idx_v, op_T3_mem_zp_idx_port_7);
  spice_transistor_nmos_gnd g_4366((~ir7_v[`W-1]|~irline3_v[`W-1]|~ir6_v[`W-1]|~clock2_v[`W-1]|~ir4_v[`W-1]|~notir2_v[`W-1]|~notir5_v[`W-1]), op_T__bit_v, op_T__bit_port_10);
  spice_transistor_nmos_gnd g_4361((~n_1184_v[`W-1]|~n_1643_v[`W-1]), n_410_v, n_410_port_6);
  spice_transistor_nmos_gnd g_4360((pd6_v|~clearIR_v[`W-1]), pd6_clearIR_v, pd6_clearIR_port_4);
  spice_transistor_nmos_gnd g_4363((~ir4_v[`W-1]|~notir3_v[`W-1]|~irline3_v[`W-1]|~notir6_v[`W-1]|~clock2_v[`W-1]|~notir7_v[`W-1]|~notir2_v[`W-1]), op_T__cpx_cpy_abs_v, op_T__cpx_cpy_abs_port_10);
  spice_transistor_nmos_gnd g_4362((~n_771_v[`W-1]|~n_850_v[`W-1]), n_1446_v, n_1446_port_4);
  spice_transistor_nmos_gnd g_4369((~_t2_v[`W-1]|~ir3_v[`W-1]|~notir2_v[`W-1]), op_T2_zp_zp_idx_v, op_T2_zp_zp_idx_port_5);
  spice_transistor_nmos_gnd g_4368((~irline3_v[`W-1]|~ir6_v[`W-1]|~notir5_v[`W-1]|~notir2_v[`W-1]|~ir7_v[`W-1]|~clock1_v[`W-1]|~ir4_v[`W-1]), x_op_T0_bit_v, x_op_T0_bit_port_9);
  spice_transistor_nmos_gnd g_4772((~alua6_v[`W-1]&~alub6_v[`W-1]), n_336_v, n_336_port_7);
  spice_transistor_nmos_gnd g_4776((~n_410_v[`W-1]&~n_392_v[`W-1]), n_344_v, n_344_port_8);
  spice_transistor_nmos_gnd g_4775((pipeUNK07_v&pipeUNK09_v), n_1111_v, n_1111_port_6);
  spice_transistor_nmos t72(~dpc1_SBY_v[`W-1], y6_v, sb6_v, y6_port_1, sb6_port_1);
  spice_transistor_nmos_vdd t76(~n_127_v[`W-1], clk2out_v, clk2out_port_0);
  spice_transistor_nmos t77(~dpc1_SBY_v[`W-1], y4_v, sb4_v, y4_port_0, sb4_port_2);
  spice_transistor_nmos_gnd t74(~n_1318_v[`W-1], n_748_v, n_748_port_0);
  spice_transistor_nmos_vdd t75(~dpc14_SRS_v[`W-1], n_304_v, n_304_port_0);
  spice_transistor_nmos_gnd t2569(~n_1541_v[`W-1], n_491_v, n_491_port_1);
  spice_transistor_nmos_gnd t8(~db2_v[`W-1], n_1199_v, n_1199_port_0);
  spice_transistor_nmos_vdd t4(~n_826_v[`W-1], ab8_v, ab8_port_0);
  spice_transistor_nmos_gnd t5(~db1_v[`W-1], n_1319_v, n_1319_port_0);
  spice_transistor_nmos_gnd t2(~notalucout_v[`W-1], alucout_v, alucout_port_0);
  spice_transistor_nmos_gnd g_4288((~n_979_v[`W-1]|~n_550_v[`W-1]|~n_782_v[`W-1]|~n_862_v[`W-1]|~nnT2BR_v[`W-1]|~op_T0_shift_a_v[`W-1]), n_1347_v, n_1347_port_8);
  spice_transistor_nmos_gnd g_4289((~notir7_v[`W-1]|~notir3_v[`W-1]|~ir4_v[`W-1]|~notir6_v[`W-1]|~clock2_v[`W-1]|~ir5_v[`W-1]|~notir1_v[`W-1]|~ir2_v[`W-1]), op_T__dex_v, op_T__dex_port_10);
  spice_transistor_nmos_gnd t880(~idb2_v[`W-1], n_458_v, n_458_port_0);
  spice_transistor_nmos_gnd t881(pchp4_v, n_27_v, n_27_port_0);
  spice_transistor_nmos_gnd t883(~pcl5_v[`W-1], n_386_v, n_386_port_0);
  spice_transistor_nmos_gnd t886(pipeUNK18_v, n_850_v, n_850_port_0);
  spice_transistor_nmos_vdd t1602(~cclk_v[`W-1], idb7_v, idb7_port_3);
  spice_transistor_nmos_gnd g_4909((~n_1115_v[`W-1]|(~n_270_v[`W-1]&~n_620_v[`W-1])), BRtaken_v, BRtaken_port_10);
  spice_transistor_nmos_gnd g_4908((~n_330_v[`W-1]|(~cclk_v[`W-1]&~n_1599_v[`W-1])), n_807_v, n_807_port_5);
  spice_transistor_nmos_gnd g_4901(((~op_T__cpx_cpy_imm_zp_v[`W-1]|~x_op_T__adc_sbc_v[`W-1]|~op_T__cpx_cpy_abs_v[`W-1]|~op_T__asl_rol_a_v[`W-1]|~op_T__cmp_v[`W-1])|(~op_asl_rol_v[`W-1]&~n_1258_v[`W-1])), _op_set_C_v, _op_set_C_port_10);
  spice_transistor_nmos_gnd g_4900(((~A_B3_v[`W-1]&~C23_v[`W-1])|(~DC34_v[`W-1]|~n_988_v[`W-1])), _C34_v, _C34_port_9);
  spice_transistor_nmos_gnd g_4903((~n_410_v[`W-1]|(~n_1184_v[`W-1]&~n_1643_v[`W-1])), n_474_v, n_474_port_5);
  spice_transistor_nmos_gnd g_4902(((~n_16_v[`W-1]&pipeT2out_v)|(pipeT3out_v&~notRdy0_v[`W-1])), n_428_v, n_428_port_6);
  spice_transistor_nmos_gnd g_4905(((pipeUNK05_v&~n_1614_v[`W-1])|(~n_1416_v[`W-1]&~n_1111_v[`W-1])|~n_587_v[`W-1]|(~n_1245_v[`W-1]&pipeUNK03_v)), n_299_v, n_299_port_9);
  spice_transistor_nmos_gnd g_4904(((~n_1398_v[`W-1]&~C67_v[`W-1])|~n_637_v[`W-1]), notaluvout_v, notaluvout_port_5);
  spice_transistor_nmos_gnd g_4907((~NMIP_v[`W-1]|(~n_1392_v[`W-1]&~cclk_v[`W-1])), n_297_v, n_297_port_5);
  spice_transistor_nmos_gnd g_4906(((~op_T3_ind_y_v[`W-1]|~x_op_T0_tya_v[`W-1]|~op_T0_cpy_iny_v[`W-1]|~op_T0_iny_dey_v[`W-1]|~op_T2_abs_y_v[`W-1])|(~n_335_v[`W-1]&~op_sty_cpy_mem_v[`W-1])|(~op_T2_idx_x_xy_v[`W-1]&~op_xy_v[`W-1])), n_1717_v, n_1717_port_12);
  spice_transistor_nmos_gnd t3440(n_1338_v, n_462_v, n_462_port_2);
  spice_transistor_nmos_vdd t3442(~n_7_v[`W-1], db6_v, db6_port_4);
  spice_transistor_nmos_gnd t3445(n_680_v, n_1526_v, n_1526_port_1);
  spice_transistor_nmos_vdd t3331(~cclk_v[`W-1], idb1_v, idb1_port_10);
  spice_transistor_nmos_gnd t2738(~n_1441_v[`W-1], dpc42_DL_ADH_v, dpc42_DL_ADH_port_8);
  spice_transistor_nmos_gnd t2228(~n_1549_v[`W-1], n_929_v, n_929_port_1);
  spice_transistor_nmos t2731(~cclk_v[`W-1], x5_v, n_578_v, x5_port_2, n_578_port_0);
  spice_transistor_nmos_vdd t2222(~n_1191_v[`W-1], ab6_v, ab6_port_0);
  spice_transistor_nmos_vdd t2221(~cclk_v[`W-1], adl1_v, adl1_port_3);
  spice_transistor_nmos_gnd t2732(~op_T0_tsx_v[`W-1], n_1586_v, n_1586_port_1);
  spice_transistor_nmos_gnd t2226(~n_1499_v[`W-1], n_709_v, n_709_port_0);
  spice_transistor_nmos_vdd t2736(~cclk_v[`W-1], adl0_v, adl0_port_6);
  spice_transistor_nmos_gnd t418(~idb5_v[`W-1], n_1383_v, n_1383_port_0);
  spice_transistor_nmos_vdd t416(~cclk_v[`W-1], sb6_v, sb6_port_4);
  spice_transistor_nmos t415(~dpc30_ADHPCH_v[`W-1], pch6_v, adh6_v, pch6_port_0, adh6_port_1);
  spice_transistor_nmos t414(~dpc30_ADHPCH_v[`W-1], pch7_v, adh7_v, pch7_port_1, adh7_port_1);
  spice_transistor_nmos t413(~dpc30_ADHPCH_v[`W-1], pch4_v, adh4_v, pch4_port_1, adh4_port_1);
  spice_transistor_nmos t412(~dpc30_ADHPCH_v[`W-1], pch5_v, adh5_v, pch5_port_0, adh5_port_1);
  spice_transistor_nmos t411(~dpc30_ADHPCH_v[`W-1], pch2_v, adh2_v, pch2_port_0, adh2_port_1);
  spice_transistor_nmos t410(~dpc30_ADHPCH_v[`W-1], pch3_v, adh3_v, pch3_port_1, adh3_port_2);
  spice_transistor_nmos_gnd g_4758((~alub4_v[`W-1]&~alua4_v[`W-1]), n_1063_v, n_1063_port_7);
  spice_transistor_nmos_gnd g_4754(((~n_743_v[`W-1]|~n_1488_v[`W-1])&~n_609_v[`W-1]), n_1192_v, n_1192_port_3);
  spice_transistor_nmos_gnd g_4750((~n_1044_v[`W-1]&(~op_rol_ror_v[`W-1]|~op_T0_adc_sbc_v[`W-1])), n_1408_v, n_1408_port_3);
  spice_transistor_nmos_gnd g_4753((~C34_v[`W-1]&~n_700_v[`W-1]), n_695_v, n_695_port_3);
  spice_transistor_nmos_vdd t15(~n_1140_v[`W-1], ab9_v, ab9_port_0);
  spice_transistor_nmos_gnd t10(n_190_v, n_220_v, n_220_port_0);
  spice_transistor_nmos_vdd t11(~n_38_v[`W-1], n_1247_v, n_1247_port_0);
  spice_transistor_nmos_gnd t789(~n_1300_v[`W-1], ir2_v, ir2_port_0);
  spice_transistor_nmos t1859(~dpc25_SBDB_v[`W-1], idb4_v, sb4_v, idb4_port_4, sb4_port_8);
  spice_transistor_nmos t1858(~dpc25_SBDB_v[`W-1], sb3_v, idb3_v, sb3_port_7, idb3_port_3);
  spice_transistor_nmos t1855(~dpc25_SBDB_v[`W-1], sb0_v, idb0_v, sb0_port_6, idb0_port_7);
  spice_transistor_nmos t1857(~dpc25_SBDB_v[`W-1], idb2_v, sb2_v, idb2_port_5, sb2_port_7);
  spice_transistor_nmos t1856(~dpc25_SBDB_v[`W-1], sb1_v, idb1_v, sb1_port_7, idb1_port_4);
  spice_transistor_nmos_gnd t1850(~n_251_v[`W-1], RnWstretched_v, RnWstretched_port_22);
  spice_transistor_nmos t1677(~dpc41_DL_ADL_v[`W-1], adl5_v, n_1387_v, adl5_port_2, n_1387_port_2);
  spice_transistor_nmos_gnd g_4923(((~dpc36_IPC_v[`W-1]&~n_937_v[`W-1])|~n_1345_v[`W-1]), n_1500_v, n_1500_port_5);
  spice_transistor_nmos_gnd g_4922(((~n_432_v[`W-1]&~n_345_v[`W-1])|~n_1097_v[`W-1]), dasb3_v, dasb3_port_5);
  spice_transistor_nmos_gnd g_4921(((~n_440_v[`W-1]&~op_inc_nop_v[`W-1])|(~op_T4_ind_y_v[`W-1]|~op_T3_ind_x_v[`W-1]|~op_T2_ind_y_v[`W-1]|~op_T3_abs_idx_v[`W-1]|~op_plp_pla_v[`W-1])), n_1107_v, n_1107_port_10);
  spice_transistor_nmos_gnd g_4920(((~n_1070_v[`W-1]&~n_919_v[`W-1])|~n_200_v[`W-1]), n_1486_v, n_1486_port_5);
  spice_transistor_nmos_gnd g_4927(((~n_243_v[`W-1]&~n_781_v[`W-1])|(~n_1170_v[`W-1]&pipeUNK14_v)|(~n_755_v[`W-1]&~_DBZ_v[`W-1])), n_566_v, n_566_port_8);
  spice_transistor_nmos_gnd g_4926((((~n_646_v[`W-1]|~nnT2BR_v[`W-1])&~n_480_v[`W-1])|n_50_v), n_629_v, n_629_port_5);
  spice_transistor_nmos_gnd g_4925(((~n_1056_v[`W-1]&~n_811_v[`W-1])|(~n_761_v[`W-1]&~n_1257_v[`W-1])), n_739_v, n_739_port_9);
  spice_transistor_nmos_gnd g_4924((~n_854_v[`W-1]|(~cclk_v[`W-1]&~n_995_v[`W-1])), n_975_v, n_975_port_6);
  spice_transistor_nmos_gnd g_4929((~n_1517_v[`W-1]|(~n_206_v[`W-1]&~n_853_v[`W-1])), n_916_v, n_916_port_7);
  spice_transistor_nmos_gnd g_4928((~op_T0_shift_right_a_v[`W-1]|(~n_440_v[`W-1]&~op_shift_right_v[`W-1])), n_366_v, n_366_port_5);
  spice_transistor_nmos t2503(~dpc8_nDBADD_v[`W-1], alub1_v, n_583_v, alub1_port_0, n_583_port_0);
  spice_transistor_nmos t528(~dpc21_ADDADL_v[`W-1], adl6_v, alu6_v, adl6_port_1, alu6_port_1);
  spice_transistor_nmos t527(~dpc21_ADDADL_v[`W-1], adl5_v, alu5_v, adl5_port_1, alu5_port_0);
  spice_transistor_nmos_gnd t2501(~adh0_v[`W-1], n_1668_v, n_1668_port_0);
  spice_transistor_nmos t526(~dpc21_ADDADL_v[`W-1], alu7_v, adl7_v, alu7_port_0, adl7_port_0);
  spice_transistor_nmos_gnd t524(~db5_v[`W-1], n_568_v, n_568_port_1);
  spice_transistor_nmos t2504(~dpc8_nDBADD_v[`W-1], alub3_v, n_1621_v, alub3_port_2, n_1621_port_0);
  spice_transistor_nmos t522(~dpc21_ADDADL_v[`W-1], adl4_v, alu4_v, adl4_port_1, alu4_port_1);
  spice_transistor_nmos_vdd t2179(~n_1399_v[`W-1], cp1_v, cp1_port_75);
  spice_transistor_nmos_gnd t2508(pipeUNK02_v, n_1492_v, n_1492_port_0);
  spice_transistor_nmos t2241(~dpc26_ACDB_v[`W-1], n_326_v, idb6_v, n_326_port_2, idb6_port_7);
  spice_transistor_nmos t2240(~dpc26_ACDB_v[`W-1], n_831_v, idb5_v, n_831_port_1, idb5_port_5);
  spice_transistor_nmos_gnd t2248(~s0_v[`W-1], n_983_v, n_983_port_1);
  spice_transistor_nmos_vdd t435(~n_1523_v[`W-1], n_635_v, n_635_port_0);
  spice_transistor_nmos_gnd t434(~n_1523_v[`W-1], n_963_v, n_963_port_1);
  spice_transistor_nmos_vdd t437(~n_1260_v[`W-1], dpc32_PCHADH_v, dpc32_PCHADH_port_1);
  spice_transistor_nmos_gnd t436(~n_1260_v[`W-1], n_1413_v, n_1413_port_1);
  spice_transistor_nmos t432(~dpc2_XSB_v[`W-1], n_1169_v, sb0_v, n_1169_port_0, sb0_port_2);
  spice_transistor_nmos_vdd t439(~n_220_v[`W-1], ADL_ABL_v, ADL_ABL_port_0);
  spice_transistor_nmos_gnd t438(~n_220_v[`W-1], n_130_v, n_130_port_0);
  spice_transistor_nmos_gnd g_4329((~idb6_v[`W-1]|~idb1_v[`W-1]|~idb0_v[`W-1]|~idb7_v[`W-1]|~idb3_v[`W-1]|~idb5_v[`W-1]|~idb4_v[`W-1]|~idb2_v[`W-1]), DBZ_v, DBZ_port_10);
  spice_transistor_nmos_gnd g_4328((~n_430_v[`W-1]|pipeUNK20_v), n_959_v, n_959_port_5);
  spice_transistor_nmos_gnd g_4321((~pd0_clearIR_v[`W-1]|~pd2_clearIR_v[`W-1]|~pd4_clearIR_v[`W-1]|~pd3_clearIR_v[`W-1]|~n_1605_v[`W-1]), PD_1xx000x0_v, PD_1xx000x0_port_7);
  spice_transistor_nmos_gnd g_4320((~n_882_v[`W-1]|n_562_v), n_1374_v, n_1374_port_5);
  spice_transistor_nmos_gnd g_4323((~op_T0_tya_v[`W-1]|~op_T__ora_and_eor_adc_v[`W-1]|~op_T__adc_sbc_v[`W-1]|~op_T0_txa_v[`W-1]|~op_T__shift_a_v[`W-1]|~op_T0_pla_v[`W-1]|~op_T0_lda_v[`W-1]), n_1455_v, n_1455_port_10);
  spice_transistor_nmos_gnd g_4322((~AxB7_v[`W-1]|~n_1038_v[`W-1]), n_269_v, n_269_port_4);
  spice_transistor_nmos_gnd g_4325((~C1x5Reset_v[`W-1]|pipe_WR_phi2_v|~notRdy0_v[`W-1]), notRnWprepad_v, notRnWprepad_port_7);
  spice_transistor_nmos_gnd g_4324((~n_630_v[`W-1]|~n_467_v[`W-1]), n_1705_v, n_1705_port_4);
  spice_transistor_nmos_gnd g_4327((~n_192_v[`W-1]|~n_236_v[`W-1]), n_506_v, n_506_port_5);
  spice_transistor_nmos_gnd g_4326((~n_1580_v[`W-1]|~n_613_v[`W-1]), n_1159_v, n_1159_port_4);
  spice_transistor_nmos_gnd t2867(~x4_v[`W-1], n_485_v, n_485_port_1);
  spice_transistor_nmos t2863(~cclk_v[`W-1], n_633_v, n_1059_v, n_633_port_0, n_1059_port_0);
  spice_transistor_nmos_gnd t2869(notdor4_v, dor4_v, dor4_port_3);
  spice_transistor_nmos_gnd t239(~op_T5_brk_v[`W-1], n_689_v, n_689_port_0);
  spice_transistor_nmos t238(~dpc42_DL_ADH_v[`W-1], adh7_v, n_1147_v, adh7_port_0, n_1147_port_0);
  spice_transistor_nmos t237(~dpc42_DL_ADH_v[`W-1], adh6_v, n_1014_v, adh6_port_0, n_1014_port_0);
  spice_transistor_nmos t236(~dpc42_DL_ADH_v[`W-1], adh5_v, n_1387_v, adh5_port_0, n_1387_port_0);
  spice_transistor_nmos t235(~dpc42_DL_ADH_v[`W-1], adh4_v, n_1095_v, adh4_port_0, n_1095_port_0);
  spice_transistor_nmos t234(~dpc42_DL_ADH_v[`W-1], adh3_v, n_1661_v, adh3_port_0, n_1661_port_0);
  spice_transistor_nmos t233(~dpc42_DL_ADH_v[`W-1], adh2_v, n_1424_v, adh2_port_0, n_1424_port_1);
  spice_transistor_nmos t232(~dpc42_DL_ADH_v[`W-1], adh1_v, n_87_v, adh1_port_0, n_87_port_0);
  spice_transistor_nmos t231(~dpc42_DL_ADH_v[`W-1], adh0_v, n_719_v, adh0_port_0, n_719_port_0);
  spice_transistor_nmos_vdd t36(~cclk_v[`W-1], sb4_v, sb4_port_0);
  spice_transistor_nmos t34(~cclk_v[`W-1], n_518_v, y6_v, n_518_port_0, y6_port_0);
  spice_transistor_nmos_gnd t35(p0_v, n_31_v, n_31_port_0);
  spice_transistor_nmos t2528(~dpc38_PCLADL_v[`W-1], n_1647_v, adl7_v, n_1647_port_1, adl7_port_5);
  spice_transistor_nmos t2529(~dpc38_PCLADL_v[`W-1], adl0_v, n_488_v, adl0_port_5, n_488_port_2);
  spice_transistor_nmos_gnd t2521(~notRdy0_v[`W-1], n_1718_v, n_1718_port_1);
  spice_transistor_nmos_vdd t2523(~n_747_v[`W-1], clk1out_v, clk1out_port_1);
  spice_transistor_nmos_gnd t2524(~n_358_v[`W-1], n_1715_v, n_1715_port_2);
  spice_transistor_nmos_gnd t3383(~res_v[`W-1], n_312_v, n_312_port_2);
  spice_transistor_nmos_gnd t3382(~n_1271_v[`W-1], dpc27_SBADH_v, dpc27_SBADH_port_9);
  spice_transistor_nmos_gnd t3439(~n_1017_v[`W-1], n_578_v, n_578_port_2);
  spice_transistor_nmos t3384(~dpc20_ADDSB06_v[`W-1], alu2_v, sb2_v, alu2_port_3, sb2_port_11);
  spice_transistor_nmos_gnd t3435(~sb3_v[`W-1], n_432_v, n_432_port_2);
  spice_transistor_nmos_vdd t3434(~n_1270_v[`W-1], dpc39_PCLPCL_v, dpc39_PCLPCL_port_11);
  spice_transistor_nmos_gnd t3437(~n_906_v[`W-1], n_714_v, n_714_port_1);
  spice_transistor_nmos_gnd t3388(nots6_v, n_618_v, n_618_port_3);
  spice_transistor_nmos_gnd t3433(~n_1270_v[`W-1], n_1518_v, n_1518_port_1);
  spice_transistor_nmos_gnd t3432(~cclk_v[`W-1], n_1585_v, n_1585_port_1);
  spice_transistor_nmos_gnd t1879(~n_1295_v[`W-1], n_1238_v, n_1238_port_1);
  spice_transistor_nmos_gnd t1873(~op_T0_cld_sed_v[`W-1], n_774_v, n_774_port_0);
  spice_transistor_nmos_gnd t1870(~_ABL3_v[`W-1], abl3_v, abl3_port_3);
  spice_transistor_nmos t1876(~dpc41_DL_ADL_v[`W-1], n_1147_v, adl7_v, n_1147_port_2, adl7_port_3);
  spice_transistor_nmos_gnd t1875(notdor6_v, dor6_v, dor6_port_2);
  spice_transistor_nmos_gnd t1874(~n_390_v[`W-1], n_1258_v, n_1258_port_4);
  spice_transistor_nmos_gnd t1385(~n_1356_v[`W-1], n_326_v, n_326_port_1);
  spice_transistor_nmos t1384(~dpc37_PCLDB_v[`W-1], n_1458_v, idb6_v, n_1458_port_0, idb6_port_3);
  spice_transistor_nmos t592(~dpc43_DL_DB_v[`W-1], idb7_v, n_1147_v, idb7_port_2, n_1147_port_1);
  spice_transistor_nmos t590(~dpc43_DL_DB_v[`W-1], idb5_v, n_1387_v, idb5_port_2, n_1387_port_1);
  spice_transistor_nmos t591(~dpc43_DL_DB_v[`W-1], idb6_v, n_1014_v, idb6_port_0, n_1014_port_1);
  spice_transistor_nmos_vdd t594(~n_322_v[`W-1], ab7_v, ab7_port_0);
  spice_transistor_nmos_gnd t1120(pclp5_v, n_72_v, n_72_port_0);
  spice_transistor_nmos_gnd t1123(~n_485_v[`W-1], n_436_v, n_436_port_0);
  spice_transistor_nmos_gnd t1650(~n_987_v[`W-1], n_1169_v, n_1169_port_1);
  spice_transistor_nmos t82(~H1x1_v[`W-1], p7_v, idb7_v, p7_port_0, idb7_port_0);
  spice_transistor_nmos_gnd g_4493((~ir2_v[`W-1]|~ir7_v[`W-1]|~_t5_v[`W-1]|~ir4_v[`W-1]|~notir6_v[`W-1]|~irline3_v[`W-1]|~ir3_v[`W-1]), op_T5_rti_rts_v, op_T5_rti_rts_port_10);
  spice_transistor_nmos_gnd g_4492((~ir3_v[`W-1]|~_t5_v[`W-1]|~notir0_v[`W-1]|~ir2_v[`W-1]), op_T5_mem_ind_idx_v, op_T5_mem_ind_idx_port_7);
  spice_transistor_nmos_gnd g_4491((~n_620_v[`W-1]|~n_270_v[`W-1]), n_1115_v, n_1115_port_4);
  spice_transistor_nmos_gnd g_4490((~clearIR_v[`W-1]|pd0_v), pd0_clearIR_v, pd0_clearIR_port_8);
  spice_transistor_nmos_gnd g_4497((~n_31_v[`W-1]|~_op_branch_bit7_v[`W-1]|~n_846_v[`W-1]), n_307_v, n_307_port_6);
  spice_transistor_nmos_gnd g_4496((~n_256_v[`W-1]|~n_192_v[`W-1]), n_25_v, n_25_port_4);
  spice_transistor_nmos_gnd g_4495((~ir3_v[`W-1]|~_t5_v[`W-1]|~notir0_v[`W-1]|~notir4_v[`W-1]|~ir2_v[`W-1]), op_T5_ind_y_v, op_T5_ind_y_port_8);
  spice_transistor_nmos_gnd g_4494((~ir3_v[`W-1]|~ir4_v[`W-1]|~ir2_v[`W-1]|~notir5_v[`W-1]|~irline3_v[`W-1]|~ir6_v[`W-1]|~_t5_v[`W-1]|~ir7_v[`W-1]), xx_op_T5_jsr_v, xx_op_T5_jsr_port_11);
  spice_transistor_nmos_gnd g_4499((~ir4_v[`W-1]|~ir7_v[`W-1]|~irline3_v[`W-1]|~notir2_v[`W-1]|~notir5_v[`W-1]|~clock1_v[`W-1]|~ir6_v[`W-1]), op_T0_bit_v, op_T0_bit_port_10);
  spice_transistor_nmos_gnd g_4498((~op_T0_bit_v[`W-1]|~op_T0_and_v[`W-1]), n_669_v, n_669_port_4);
  spice_transistor_nmos_gnd g_4339((~op_T4_mem_abs_idx_v[`W-1]|~op_T3_mem_abs_v[`W-1]|~op_T5_mem_ind_idx_v[`W-1]|~op_T3_mem_zp_idx_v[`W-1]|~op_T2_mem_zp_v[`W-1]), n_347_v, n_347_port_9);
  spice_transistor_nmos_gnd g_4332((pipephi2Reset0x_v|n_1132_v), n_717_v, n_717_port_5);
  spice_transistor_nmos_gnd g_4330((~notir7_v[`W-1]|~irline3_v[`W-1]|~clock2_v[`W-1]|~notir6_v[`W-1]|~ir4_v[`W-1]|~ir3_v[`W-1]), op_T__cpx_cpy_imm_zp_v, op_T__cpx_cpy_imm_zp_port_8);
  spice_transistor_nmos_gnd g_4331((~n_954_v[`W-1]|~n_507_v[`W-1]|~n_253_v[`W-1]), n_279_v, n_279_port_5);
  spice_transistor_nmos_gnd g_4336((~n_811_v[`W-1]|~n_1257_v[`W-1]), n_753_v, n_753_port_5);
  spice_transistor_nmos_gnd g_4337((~op_T2_v[`W-1]|~n_952_v[`W-1]|~n_630_v[`W-1]|~n_1002_v[`W-1]), n_152_v, n_152_port_6);
  spice_transistor_nmos_gnd t2266(~n_862_v[`W-1], n_445_v, n_445_port_3);
  spice_transistor_nmos_gnd t2264(~pch5_v[`W-1], n_499_v, n_499_port_0);
  spice_transistor_nmos t2263(~dpc0_YSB_v[`W-1], n_733_v, sb5_v, n_733_port_1, sb5_port_7);
  spice_transistor_nmos t2262(~dpc0_YSB_v[`W-1], n_518_v, sb6_v, n_518_port_2, sb6_port_10);
  spice_transistor_nmos_gnd t2261(n_47_v, n_603_v, n_603_port_1);
  spice_transistor_nmos t2260(~dpc0_YSB_v[`W-1], n_658_v, sb4_v, n_658_port_1, sb4_port_10);
  spice_transistor_nmos_gnd g_4303((n_459_v|~n_43_v[`W-1]), n_625_v, n_625_port_5);
  spice_transistor_nmos t450(~dpc9_DBADD_v[`W-1], alub0_v, idb0_v, alub0_port_3, idb0_port_4);
  spice_transistor_nmos_vdd t456(~cclk_v[`W-1], adh1_v, adh1_port_2);
  spice_transistor_nmos t455(~dpc2_XSB_v[`W-1], n_871_v, sb7_v, n_871_port_0, sb7_port_1);
  spice_transistor_nmos_gnd t459(~abl3_v[`W-1], n_990_v, n_990_port_0);
  spice_transistor_nmos_gnd t458(~abl3_v[`W-1], n_138_v, n_138_port_0);
  spice_transistor_nmos_gnd t1462(~_t3_v[`W-1], op_T3_v, op_T3_port_0);
  spice_transistor_nmos_gnd t215(~alucout_v[`W-1], n_206_v, n_206_port_0);
  spice_transistor_nmos_gnd t217(~n_241_v[`W-1], n_1033_v, n_1033_port_0);
  spice_transistor_nmos_gnd t213(~n_867_v[`W-1], n_876_v, n_876_port_0);
  spice_transistor_nmos_vdd t218(~n_241_v[`W-1], dpc21_ADDADL_v, dpc21_ADDADL_port_0);
  spice_transistor_nmos_gnd g_4686((~n_923_v[`W-1]|~n_293_v[`W-1]), n_810_v, n_810_port_4);
  spice_transistor_nmos_gnd g_4684((pd1_v|~clearIR_v[`W-1]), pd1_clearIR_v, pd1_clearIR_port_6);
  spice_transistor_nmos_gnd g_4682((~C67_v[`W-1]|~n_1318_v[`W-1]), n_637_v, n_637_port_4);
  spice_transistor_nmos_gnd g_4683((~ir6_v[`W-1]|~ir7_v[`W-1]|~notir1_v[`W-1]), op_asl_rol_v, op_asl_rol_port_7);
  spice_transistor_nmos_gnd g_4680((~op_T2_brk_v[`W-1]|~op_T3_jsr_v[`W-1]), n_824_v, n_824_port_6);
  spice_transistor_nmos_gnd g_4681((n_18_v|~n_1357_v[`W-1]), n_378_v, n_378_port_5);
  spice_transistor_nmos_gnd g_4689(((~n_1253_v[`W-1]|~n_163_v[`W-1])&~n_1184_v[`W-1]), n_1631_v, n_1631_port_3);
  spice_transistor_nmos_gnd t869(~n_291_v[`W-1], n_1157_v, n_1157_port_0);
  spice_transistor_nmos_gnd t3410(~n_794_v[`W-1], db1_v, db1_port_4);
  spice_transistor_nmos_vdd t1679(~n_42_v[`W-1], db3_v, db3_port_2);
  spice_transistor_nmos_gnd t2040(~n_196_v[`W-1], dpc5_SADL_v, dpc5_SADL_port_7);
  spice_transistor_nmos t2595(~dpc13_ORS_v[`W-1], n_1632_v, n_277_v, n_1632_port_4, n_277_port_5);
  spice_transistor_nmos t1676(~dpc41_DL_ADL_v[`W-1], adl6_v, n_1014_v, adl6_port_2, n_1014_port_2);
  spice_transistor_nmos_gnd t2107(~n_1138_v[`W-1], n_767_v, n_767_port_1);
  spice_transistor_nmos_gnd t2101(~n_171_v[`W-1], ab7_v, ab7_port_1);
  spice_transistor_nmos_gnd t860(~adl7_v[`W-1], n_1046_v, n_1046_port_0);
  spice_transistor_nmos_gnd t861(~n_1107_v[`W-1], n_389_v, n_389_port_1);
  spice_transistor_nmos_gnd t866(~y2_v[`W-1], n_1484_v, n_1484_port_0);
  spice_transistor_nmos t2108(~cp1_v[`W-1], n_1387_v, idl5_v, n_1387_port_3, idl5_port_0);
  spice_transistor_nmos_gnd t2109(~n_815_v[`W-1], n_0_ADL2_v, n_0_ADL2_port_0);
  spice_transistor_nmos t1103(~cclk_v[`W-1], n_1724_v, x6_v, n_1724_port_1, x6_port_0);
  spice_transistor_nmos_vdd t1101(~cclk_v[`W-1], adl3_v, adl3_port_1);
  spice_transistor_nmos t1107(~dpc17_SUMS_v[`W-1], __AxBxC_1_v, notaluoutmux1_v, __AxBxC_1_port_1, notaluoutmux1_port_1);
  spice_transistor_nmos t1106(~dpc17_SUMS_v[`W-1], __AxBxC_0_v, notaluoutmux0_v, __AxBxC_0_port_2, notaluoutmux0_port_1);
  spice_transistor_nmos_gnd t1105(~n_1238_v[`W-1], dpc25_SBDB_v, dpc25_SBDB_port_0);
  spice_transistor_nmos t1109(~dpc17_SUMS_v[`W-1], __AxBxC_3_v, n_1071_v, __AxBxC_3_port_1, n_1071_port_3);
  spice_transistor_nmos t1108(~dpc17_SUMS_v[`W-1], __AxBxC_2_v, n_740_v, __AxBxC_2_port_1, n_740_port_2);
  spice_transistor_nmos_gnd g_4516((~n_1518_v[`W-1]|~n_1247_v[`W-1]|~cclk_v[`W-1]), dpc39_PCLPCL_v, dpc39_PCLPCL_port_12);
  spice_transistor_nmos_gnd g_4517((~dor2_v[`W-1]|~RnWstretched_v[`W-1]), n_224_v, n_224_port_5);
  spice_transistor_nmos_gnd g_4514((~nnT2BR_v[`W-1]|~n_1286_v[`W-1]|~n_862_v[`W-1]|~n_1002_v[`W-1]|~op_T2_abs_access_v[`W-1]), n_1211_v, n_1211_port_9);
  spice_transistor_nmos_gnd g_4515((~brk_done_v[`W-1]|p2_v), n_334_v, n_334_port_6);
  spice_transistor_nmos_gnd g_4512((~brk_done_v[`W-1]|~n_717_v[`W-1]), n_1087_v, n_1087_port_4);
  spice_transistor_nmos_gnd g_4510((~n_1247_v[`W-1]|~n_1043_v[`W-1]|~cclk_v[`W-1]), dpc40_ADLPCL_v, dpc40_ADLPCL_port_12);
  spice_transistor_nmos_gnd g_4511((~clearIR_v[`W-1]|pd7_v), pd7_clearIR_v, pd7_clearIR_port_5);
  spice_transistor_nmos_gnd g_4518((~RnWstretched_v[`W-1]|~n_224_v[`W-1]), n_520_v, n_520_port_4);
  spice_transistor_nmos_gnd g_4519((~op_ANDS_v[`W-1]|~n_946_v[`W-1]|~n_1412_v[`W-1]|~n_1258_v[`W-1]), n_384_v, n_384_port_8);
  spice_transistor_nmos_gnd g_4479((~ir6_v[`W-1]|~notir0_v[`W-1]|~clock1_v[`W-1]|~ir7_v[`W-1]|~ir5_v[`W-1]), op_T0_ora_v, op_T0_ora_port_7);
  spice_transistor_nmos_gnd t679(~ir6_v[`W-1], _op_branch_bit6_v, _op_branch_bit6_port_0);
  spice_transistor_nmos_gnd g_4475((~notRdy0_v[`W-1]|~n_152_v[`W-1]), n_1343_v, n_1343_port_5);
  spice_transistor_nmos_gnd g_4474((~ir7_v[`W-1]|~clock1_v[`W-1]|~ir2_v[`W-1]|~ir5_v[`W-1]|~irline3_v[`W-1]|~ir4_v[`W-1]|~notir3_v[`W-1]), op_T0_php_pha_v, op_T0_php_pha_port_10);
  spice_transistor_nmos_gnd g_4477((~ir4_v[`W-1]|~ir7_v[`W-1]|~ir2_v[`W-1]|~irline3_v[`W-1]|~_t2_v[`W-1]), op_T2_stack_v, op_T2_stack_port_8);
  spice_transistor_nmos_gnd g_4471((~_t2_v[`W-1]|~ir4_v[`W-1]|~ir2_v[`W-1]|~ir7_v[`W-1]|~irline3_v[`W-1]), op_T2_stack_access_v, op_T2_stack_access_port_7);
  spice_transistor_nmos_gnd g_4470((~notir0_v[`W-1]|~ir4_v[`W-1]|~_t4_v[`W-1]|~ir2_v[`W-1]|~ir3_v[`W-1]), op_T4_ind_x_v, op_T4_ind_x_port_9);
  spice_transistor_nmos_gnd g_4473((~ir2_v[`W-1]|~_t5_v[`W-1]|~ir5_v[`W-1]|~ir6_v[`W-1]|~ir7_v[`W-1]|~ir3_v[`W-1]|~irline3_v[`W-1]|~ir4_v[`W-1]), op_T5_brk_v, op_T5_brk_port_12);
  spice_transistor_nmos_gnd g_4472((~irline3_v[`W-1]|~ir2_v[`W-1]|~notir3_v[`W-1]|~notir4_v[`W-1]|~clock1_v[`W-1]|~notir7_v[`W-1]|~ir5_v[`W-1]|~ir6_v[`W-1]), op_T0_tya_v, op_T0_tya_port_11);
  spice_transistor_nmos_gnd t1656(n_126_v, pchp1_v, pchp1_port_0);
  spice_transistor_nmos_gnd t475(~rdy_v[`W-1], n_958_v, n_958_port_0);
  spice_transistor_nmos_gnd t477(~n_1240_v[`W-1], dpc43_DL_DB_v, dpc43_DL_DB_port_0);
  spice_transistor_nmos_gnd t2829(~x2_v[`W-1], n_890_v, n_890_port_1);
  spice_transistor_nmos_gnd t2822(~a1_v[`W-1], n_1549_v, n_1549_port_1);
  spice_transistor_nmos_gnd t1651(n_95_v, n_531_v, n_531_port_0);
  spice_transistor_nmos_gnd t2826(~n_770_v[`W-1], n_853_v, n_853_port_2);
  spice_transistor_nmos_gnd t272(~n_1575_v[`W-1], _t2_v, _t2_port_0);
  spice_transistor_nmos_vdd t276(~n_631_v[`W-1], dpc37_PCLDB_v, dpc37_PCLDB_port_0);
  spice_transistor_nmos_gnd t275(~n_631_v[`W-1], n_1323_v, n_1323_port_0);
  spice_transistor_nmos_vdd t279(~cclk_v[`W-1], adl4_v, adl4_port_0);
  spice_transistor_nmos t2525(~dpc38_PCLADL_v[`W-1], adl4_v, n_208_v, adl4_port_5, n_208_port_2);
  spice_transistor_nmos_gnd t3470(~n_329_v[`W-1], n_1166_v, n_1166_port_2);
  spice_transistor_nmos_gnd t3473(~n_1072_v[`W-1], db0_v, db0_port_4);
  spice_transistor_nmos_gnd t1835(~idb6_v[`W-1], n_1684_v, n_1684_port_1);
  spice_transistor_nmos_gnd t1834(~n_503_v[`W-1], n_270_v, n_270_port_2);
  spice_transistor_nmos_gnd t1347(~pcl1_v[`W-1], n_329_v, n_329_port_0);
  spice_transistor_nmos_gnd t1341(~dpc12_0ADD_v[`W-1], alua7_v, alua7_port_0);
  spice_transistor_nmos_gnd t1342(~n_1715_v[`W-1], n_1399_v, n_1399_port_0);
  spice_transistor_nmos_gnd t2128(~db6_v[`W-1], n_374_v, n_374_port_1);
  spice_transistor_nmos t2129(~H1x1_v[`W-1], Pout3_v, idb3_v, Pout3_port_3, idb3_port_5);
  spice_transistor_nmos_gnd t2126(n_1579_v, n_221_v, n_221_port_1);
  spice_transistor_nmos t2127(~H1x1_v[`W-1], p4_v, idb4_v, p4_port_1, idb4_port_5);
  spice_transistor_nmos_gnd t2120(~clk0_v[`W-1], n_358_v, n_358_port_2);
  spice_transistor_nmos t2123(~dpc3_SBX_v[`W-1], x0_v, sb0_v, x0_port_0, sb0_port_7);
  spice_transistor_nmos_vdd t1169(~n_519_v[`W-1], n_135_v, n_135_port_1);
  spice_transistor_nmos_vdd t1699(~n_543_v[`W-1], dpc5_SADL_v, dpc5_SADL_port_0);
  spice_transistor_nmos_gnd t1698(~n_543_v[`W-1], n_196_v, n_196_port_0);
  spice_transistor_nmos_gnd t1693(n_1124_v, n_1662_v, n_1662_port_1);
  spice_transistor_nmos t1160(~dpc8_nDBADD_v[`W-1], alub0_v, n_624_v, alub0_port_4, n_624_port_1);
  spice_transistor_nmos_gnd t1697(n_226_v, n_1593_v, n_1593_port_2);
  spice_transistor_nmos_gnd t1694(n_1269_v, n_1401_v, n_1401_port_0);
  spice_transistor_nmos_gnd g_4530((~notRdy0_v[`W-1]|pipeUNK09_v), n_781_v, n_781_port_13);
  spice_transistor_nmos_gnd g_4531((~op_rmw_v[`W-1]|~n_347_v[`W-1]|~x_op_jmp_v[`W-1]), n_510_v, n_510_port_6);
  spice_transistor_nmos_gnd g_4532((~op_jsr_v[`W-1]|~x_op_jmp_v[`W-1]|~op_brk_rti_v[`W-1]), n_134_v, n_134_port_7);
  spice_transistor_nmos_gnd g_4533((~nnT2BR_v[`W-1]|~n_236_v[`W-1]), n_1427_v, n_1427_port_4);
  spice_transistor_nmos_gnd g_4534((~n_288_v[`W-1]|~RnWstretched_v[`W-1]), n_798_v, n_798_port_4);
  spice_transistor_nmos_gnd g_4535((~n_846_v[`W-1]|~n_1045_v[`W-1]|~n_201_v[`W-1]), n_1371_v, n_1371_port_6);
  spice_transistor_nmos_gnd g_4536((~notir0_v[`W-1]|~ir5_v[`W-1]|~ir6_v[`W-1]|~notir7_v[`W-1]), op_sta_cmp_v, op_sta_cmp_port_6);
  spice_transistor_nmos_gnd g_4537((~notir6_v[`W-1]|~clock2_v[`W-1]|~notir0_v[`W-1]|~notir5_v[`W-1]), op_T__adc_sbc_v, op_T__adc_sbc_port_7);
  spice_transistor_nmos_gnd g_4538((~notir0_v[`W-1]|~ir7_v[`W-1]|~clock2_v[`W-1]), op_T__ora_and_eor_adc_v, op_T__ora_and_eor_adc_port_6);
  spice_transistor_nmos_gnd g_4539((~notir5_v[`W-1]|~notir0_v[`W-1]|~ir6_v[`W-1]|~clock1_v[`W-1]|~ir7_v[`W-1]), op_T0_and_v, op_T0_and_port_8);
  spice_transistor_nmos_gnd g_4457((~n_1135_v[`W-1]|~n_753_v[`W-1]), n_1629_v, n_1629_port_4);
  spice_transistor_nmos_gnd g_4456((~dor7_v[`W-1]|~RnWstretched_v[`W-1]), n_23_v, n_23_port_5);
  spice_transistor_nmos_gnd g_4455((~cclk_v[`W-1]|~n_969_v[`W-1]|~n_1247_v[`W-1]), dpc0_YSB_v, dpc0_YSB_port_12);
  spice_transistor_nmos_gnd g_4454((~op_SRS_v[`W-1]|~op_ORS_v[`W-1]|~op_EORS_v[`W-1]|~op_ANDS_v[`W-1]), op_SUMS_v, op_SUMS_port_6);
  spice_transistor_nmos_gnd g_4453((~n_470_v[`W-1]|~n_134_v[`W-1]), n_467_v, n_467_port_6);
  spice_transistor_nmos_gnd g_4452((~n_1247_v[`W-1]|~cclk_v[`W-1]|~n_763_v[`W-1]), dpc8_nDBADD_v, dpc8_nDBADD_port_12);
  spice_transistor_nmos_gnd g_4451((~notRdy0_v[`W-1]|~n_861_v[`W-1]), brk_done_v, brk_done_port_12);
  spice_transistor_nmos_gnd g_4450((~cclk_v[`W-1]|n_1113_v), n_161_v, n_161_port_5);
  spice_transistor_nmos_gnd g_4459((~clearIR_v[`W-1]|pd4_v), pd4_clearIR_v, pd4_clearIR_port_8);
  spice_transistor_nmos_gnd g_4458((~clearIR_v[`W-1]|pd3_v), pd3_clearIR_v, pd3_clearIR_port_6);
  spice_transistor_nmos_gnd t512(nots4_v, n_3_v, n_3_port_2);
  spice_transistor_nmos_gnd t398(~dpc29_0ADH17_v[`W-1], adh1_v, adh1_port_1);
  spice_transistor_nmos_gnd t390(~notRdy0_v[`W-1], n_16_v, n_16_port_0);
  spice_transistor_nmos_gnd t391(~db1_v[`W-1], n_213_v, n_213_port_0);
  spice_transistor_nmos_gnd t392(pipeVectorA1_v, n_0_ADL1_v, n_0_ADL1_port_0);
  spice_transistor_nmos_gnd t393(nots5_v, n_280_v, n_280_port_2);
  spice_transistor_nmos t394(~cclk_v[`W-1], n_1654_v, a3_v, n_1654_port_0, a3_port_0);
  spice_transistor_nmos_vdd t397(~n_317_v[`W-1], n_417_v, n_417_port_1);
  spice_transistor_nmos t2804(~cclk_v[`W-1], n_871_v, x7_v, n_871_port_1, x7_port_2);
  spice_transistor_nmos_gnd t2803(~n_958_v[`W-1], n_1449_v, n_1449_port_1);
  spice_transistor_nmos_gnd t2802(~n_927_v[`W-1], ir4_v, ir4_port_68);
  spice_transistor_nmos t2800(~dpc8_nDBADD_v[`W-1], alub7_v, n_423_v, alub7_port_3, n_423_port_0);
  spice_transistor_nmos_gnd t2808(~n_1211_v[`W-1], n_1655_v, n_1655_port_1);
  spice_transistor_nmos t1576(~cclk_v[`W-1], y3_v, n_1531_v, y3_port_0, n_1531_port_1);
  spice_transistor_nmos_gnd t1573(n_15_v, pclp4_v, pclp4_port_0);
  spice_transistor_nmos_gnd t1570(~alucin_v[`W-1], notalucin_v, notalucin_port_2);
  spice_transistor_nmos t259(~cclk_v[`W-1], n_242_v, x3_v, n_242_port_0, x3_port_0);
  spice_transistor_nmos t251(~dpc6_SBS_v[`W-1], sb4_v, s4_v, sb4_port_4, s4_port_0);
  spice_transistor_nmos t250(~dpc6_SBS_v[`W-1], s3_v, sb3_v, s3_port_0, sb3_port_2);
  spice_transistor_nmos t253(~dpc6_SBS_v[`W-1], s2_v, sb2_v, s2_port_0, sb2_port_2);
  spice_transistor_nmos t252(~dpc6_SBS_v[`W-1], s1_v, sb1_v, s1_port_0, sb1_port_1);
  spice_transistor_nmos t1523(~dpc3_SBX_v[`W-1], sb4_v, x4_v, sb4_port_6, x4_port_0);
  spice_transistor_nmos_vdd t3458(~n_634_v[`W-1], ab4_v, ab4_port_1);
  spice_transistor_nmos_gnd t3457(~n_1358_v[`W-1], n_396_v, n_396_port_1);
  spice_transistor_nmos_gnd t3321(notalu3_v, alu3_v, alu3_port_2);
  spice_transistor_nmos_vdd t3323(~n_1277_v[`W-1], dpc42_DL_ADH_v, dpc42_DL_ADH_port_9);
  spice_transistor_nmos_gnd t3322(~n_1277_v[`W-1], n_1441_v, n_1441_port_1);
  spice_transistor_nmos_gnd t2328(~n_1133_v[`W-1], irline3_v, irline3_port_0);
  spice_transistor_nmos_gnd t2495(pipeUNK37_v, n_198_v, n_198_port_2);
  spice_transistor_nmos_gnd t2321(~aluanorb0_v[`W-1], aluaorb0_v, aluaorb0_port_1);
  spice_transistor_nmos_gnd t1369(notidl0_v, idl0_v, idl0_port_1);
  spice_transistor_nmos_gnd t1365(~idb4_v[`W-1], n_478_v, n_478_port_1);
  spice_transistor_nmos t2242(~dpc26_ACDB_v[`W-1], n_1592_v, idb7_v, n_1592_port_2, idb7_port_7);
  spice_transistor_nmos t538(~dpc13_ORS_v[`W-1], n_740_v, n_1691_v, n_740_port_0, n_1691_port_1);
  spice_transistor_nmos_gnd t534(~n_990_v[`W-1], n_1041_v, n_1041_port_1);
  spice_transistor_nmos_vdd t535(~n_990_v[`W-1], n_138_v, n_138_port_1);
  spice_transistor_nmos_gnd t2246(~n_1649_v[`W-1], n_795_v, n_795_port_0);
  spice_transistor_nmos_vdd t2148(~cclk_v[`W-1], adh5_v, adh5_port_2);
  spice_transistor_nmos_vdd t2149(~cclk_v[`W-1], adl6_v, adl6_port_3);
  spice_transistor_nmos_gnd t2143(~n_108_v[`W-1], dpc16_EORS_v, dpc16_EORS_port_8);
  spice_transistor_nmos_gnd t2140(notdor0_v, dor0_v, dor0_port_0);
  spice_transistor_nmos_gnd t2141(~aluvout_v[`W-1], n_1245_v, n_1245_port_1);
  spice_transistor_nmos t2146(~cclk_v[`W-1], n_1169_v, x0_v, n_1169_port_2, x0_port_1);
  spice_transistor_nmos_gnd t2145(~n_850_v[`W-1], n_430_v, n_430_port_2);
  spice_transistor_nmos_gnd g_4558((~_t4_v[`W-1]|~notir3_v[`W-1]|~notir4_v[`W-1]), op_T4_abs_idx_v, op_T4_abs_idx_port_6);
  spice_transistor_nmos_gnd g_4559((~alub2_v[`W-1]|~alua2_v[`W-1]), n_1691_v, n_1691_port_8);
  spice_transistor_nmos_gnd g_4552((~_DBE_v[`W-1]|~n_221_v[`W-1]), n_251_v, n_251_port_5);
  spice_transistor_nmos_gnd g_4553((~cclk_v[`W-1]|n_1404_v), n_133_v, n_133_port_5);
  spice_transistor_nmos_gnd g_4550((~RnWstretched_v[`W-1]|~dor5_v[`W-1]), n_612_v, n_612_port_4);
  spice_transistor_nmos_gnd g_4551((~ir4_v[`W-1]|~irline3_v[`W-1]|~_t3_v[`W-1]|~ir7_v[`W-1]), op_T3_stack_bit_jmp_v, op_T3_stack_bit_jmp_port_7);
  spice_transistor_nmos_gnd g_4556((~cclk_v[`W-1]|~n_1247_v[`W-1]|~n_1335_v[`W-1]), dpc24_ACSB_v, dpc24_ACSB_port_12);
  spice_transistor_nmos_gnd g_4557((~notir5_v[`W-1]|~ir4_v[`W-1]|~notir3_v[`W-1]|~ir2_v[`W-1]|~ir7_v[`W-1]|~irline3_v[`W-1]|~notir6_v[`W-1]|~clock1_v[`W-1]), op_T0_pla_v, op_T0_pla_port_11);
  spice_transistor_nmos_gnd g_4554((~cclk_v[`W-1]|~n_1247_v[`W-1]|~n_800_v[`W-1]), dpc26_ACDB_v, dpc26_ACDB_port_12);
  spice_transistor_nmos_gnd g_4555((~notir7_v[`W-1]|~irline3_v[`W-1]|~ir4_v[`W-1]|~ir5_v[`W-1]|~notir6_v[`W-1]|~clock1_v[`W-1]), op_T0_cpy_iny_v, op_T0_cpy_iny_port_9);
  spice_transistor_nmos_gnd g_4431((~n_389_v[`W-1]|~op_T2_abs_v[`W-1]|~op_T2_jsr_v[`W-1]|~brk_done_v[`W-1]|~n_1109_v[`W-1]|~op_rti_rts_v[`W-1]|~op_jmp_v[`W-1]|~notRdy0_v[`W-1]|~op_T4_ind_x_v[`W-1]), n_1649_v, n_1649_port_12);
  spice_transistor_nmos_gnd g_4430((~_DA_ADD1_v[`W-1]|~_DA_ADD2_v[`W-1]), n_867_v, n_867_port_4);
  spice_transistor_nmos_gnd g_4433((~alub7_v[`W-1]|~alua7_v[`W-1]), n_1398_v, n_1398_port_8);
  spice_transistor_nmos_gnd g_4432((n_1477_v|~n_43_v[`W-1]), n_1541_v, n_1541_port_5);
  spice_transistor_nmos_gnd g_4435((~n_1070_v[`W-1]|~n_1007_v[`W-1]|~n_923_v[`W-1]|~n_1265_v[`W-1]|~n_1010_v[`W-1]), dpc35_PCHC_v, dpc35_PCHC_port_8);
  spice_transistor_nmos_gnd g_4436((C78_phi2_v|DC78_phi2_v), notalucout_v, notalucout_port_5);
  spice_transistor_nmos_gnd g_4439((~aluanorb1_v[`W-1]|~n_936_v[`W-1]), AxB1_v, AxB1_port_8);
  spice_transistor_nmos_gnd g_4438((~__AxB_6_v[`W-1]|~C56_v[`W-1]), _AxB_6__C56_v, _AxB_6__C56_port_4);
  spice_transistor_nmos_vdd t1515(~n_288_v[`W-1], n_794_v, n_794_port_1);
  spice_transistor_nmos t2799(~dpc8_nDBADD_v[`W-1], alub6_v, n_351_v, alub6_port_3, n_351_port_1);
  spice_transistor_nmos t2798(~dpc8_nDBADD_v[`W-1], alub5_v, n_1383_v, alub5_port_3, n_1383_port_1);
  spice_transistor_nmos_gnd t2797(~n_565_v[`W-1], n_658_v, n_658_port_2);
  spice_transistor_nmos_gnd t3156(~PD_xxxx10x0_v[`W-1], n_231_v, n_231_port_1);
  spice_transistor_nmos_gnd t3157(~pclp6_v[`W-1], n_1458_v, n_1458_port_2);
  spice_transistor_nmos_gnd t3152(~n_681_v[`W-1], DA_AB2_v, DA_AB2_port_2);
  spice_transistor_nmos_gnd t3153(~n_130_v[`W-1], ADL_ABL_v, ADL_ABL_port_5);
  spice_transistor_nmos_gnd t3150(~n_1434_v[`W-1], n_1709_v, n_1709_port_1);
  spice_transistor_nmos_gnd t3151(nots2_v, n_1389_v, n_1389_port_3);
  spice_transistor_nmos_gnd t3158(~notRdy0_v[`W-1], n_1120_v, n_1120_port_1);
  spice_transistor_nmos_gnd t1554(~n_86_v[`W-1], ab4_v, ab4_port_0);
  spice_transistor_nmos_gnd t1552(~sb2_v[`W-1], n_1580_v, n_1580_port_0);
  spice_transistor_nmos_gnd t2056(~n_676_v[`W-1], ab9_v, ab9_port_1);
  spice_transistor_nmos_gnd t2050(~n_1346_v[`W-1], n_1296_v, n_1296_port_2);
  spice_transistor_nmos_gnd t1448(~op_implied_v[`W-1], n_664_v, n_664_port_1);
  spice_transistor_nmos_vdd t2051(~n_1346_v[`W-1], n_359_v, n_359_port_2);
  spice_transistor_nmos t2053(~dpc19_ADDSB7_v[`W-1], alu7_v, sb7_v, alu7_port_1, sb7_port_6);
  spice_transistor_nmos_gnd t3309(~n_1561_v[`W-1], n_871_v, n_871_port_2);
  spice_transistor_nmos_gnd t3056(~AxB1_v[`W-1], n_953_v, n_953_port_1);
  spice_transistor_nmos_gnd t518(~ir6_v[`W-1], notir6_v, notir6_port_0);
  spice_transistor_nmos_gnd t519(~n_1225_v[`W-1], n_1222_v, n_1222_port_0);
  spice_transistor_nmos_gnd t510(~op_T2_jsr_v[`W-1], n_383_v, n_383_port_0);
  spice_transistor_nmos_gnd t516(~n_1223_v[`W-1], n_225_v, n_225_port_0);
  spice_transistor_nmos_vdd t517(~n_1223_v[`W-1], dpc9_DBADD_v, dpc9_DBADD_port_1);
  spice_transistor_nmos_gnd t514(pipeUNK06_v, n_755_v, n_755_port_0);
  spice_transistor_nmos_gnd g_4574((pipeUNK32_v|pipeUNK33_v|pipeUNK31_v|pipeUNK30_v), n_1178_v, n_1178_port_6);
  spice_transistor_nmos_gnd g_4577((~AxB3_v[`W-1]|~DA_AB2_v[`W-1]), n_1610_v, n_1610_port_5);
  spice_transistor_nmos_gnd g_4570((~notRdy0_v[`W-1]|pipeUNK34_v), n_720_v, n_720_port_4);
  spice_transistor_nmos_gnd g_4571((~n_988_v[`W-1]|~n_649_v[`W-1]), AxB3_v, AxB3_port_8);
  spice_transistor_nmos_gnd g_4572((n_360_v|~n_43_v[`W-1]), n_1230_v, n_1230_port_5);
  spice_transistor_nmos_gnd g_4573((~RnWstretched_v[`W-1]|~dor7_v[`W-1]), n_1501_v, n_1501_port_4);
  spice_transistor_nmos_gnd g_4578((~n_1691_v[`W-1]|~DA_AB2_v[`W-1]), DA_AxB2_v, DA_AxB2_port_5);
  spice_transistor_nmos_gnd g_4579((~notir3_v[`W-1]|~ir4_v[`W-1]|~ir2_v[`W-1]|~irline3_v[`W-1]|~ir7_v[`W-1]), x_op_push_pull_v, x_op_push_pull_port_8);
  spice_transistor_nmos_gnd t1307(~adh2_v[`W-1], n_168_v, n_168_port_0);
  spice_transistor_nmos t1308(~dpc10_ADLADD_v[`W-1], adl2_v, alub2_v, adl2_port_1, alub2_port_1);
  spice_transistor_nmos_gnd g_4419((~notir2_v[`W-1]|~notir6_v[`W-1]|~irline3_v[`W-1]|~notir3_v[`W-1]|~ir4_v[`W-1]|~ir7_v[`W-1]|~_t3_v[`W-1]), op_T3_jmp_v, op_T3_jmp_port_9);
  spice_transistor_nmos_gnd g_4418((~notir0_v[`W-1]|~notir5_v[`W-1]|~clock1_v[`W-1]|~notir6_v[`W-1]), op_T0_adc_sbc_v, op_T0_adc_sbc_port_8);
  spice_transistor_nmos_gnd g_4413((~clock1_v[`W-1]|~notir6_v[`W-1]|~notir0_v[`W-1]|~notir5_v[`W-1]|~notir7_v[`W-1]), op_T0_sbc_v, op_T0_sbc_port_9);
  spice_transistor_nmos_gnd g_4412((~notir0_v[`W-1]|~clock1_v[`W-1]|~notir6_v[`W-1]|~ir5_v[`W-1]|~notir7_v[`W-1]), op_T0_cmp_v, op_T0_cmp_port_7);
  spice_transistor_nmos_gnd g_4411((~notir3_v[`W-1]|~notir5_v[`W-1]|~ir7_v[`W-1]|~irline3_v[`W-1]|~ir4_v[`W-1]|~ir2_v[`W-1]), op_plp_pla_v, op_plp_pla_port_9);
  spice_transistor_nmos_gnd g_4410((~notir5_v[`W-1]|~notir1_v[`W-1]|~notir7_v[`W-1]|~notir6_v[`W-1]), op_inc_nop_v, op_inc_nop_port_6);
  spice_transistor_nmos_gnd g_4417((~notir0_v[`W-1]|~notir6_v[`W-1]|~clock1_v[`W-1]|~ir5_v[`W-1]|~ir7_v[`W-1]), op_T0_eor_v, op_T0_eor_port_7);
  spice_transistor_nmos_gnd g_4416((~irline3_v[`W-1]|~_t4_v[`W-1]|~ir3_v[`W-1]|~ir5_v[`W-1]|~ir4_v[`W-1]|~notir6_v[`W-1]|~ir7_v[`W-1]|~ir2_v[`W-1]), op_T4_rti_v, op_T4_rti_port_10);
  spice_transistor_nmos_gnd g_4415((~clock1_v[`W-1]|~ir4_v[`W-1]|~irline3_v[`W-1]|~notir7_v[`W-1]|~notir6_v[`W-1]), op_T0_cpx_cpy_inx_iny_v, op_T0_cpx_cpy_inx_iny_port_7);
  spice_transistor_nmos_gnd g_4414((~ir4_v[`W-1]|~irline3_v[`W-1]|~ir7_v[`W-1]|~ir2_v[`W-1]|~ir3_v[`W-1]|~notir6_v[`W-1]), op_rti_rts_v, op_rti_rts_port_10);
  spice_transistor_nmos_gnd t358(~idb0_v[`W-1], n_1224_v, n_1224_port_0);
  spice_transistor_nmos_gnd t356(n_1341_v, n_600_v, n_600_port_1);
  spice_transistor_nmos_gnd t350(~n_66_v[`W-1], ab1_v, ab1_port_0);

  spice_pullup pullup_3285(n_91_v, n_91_port_3);
  spice_pullup pullup_3284(n_90_v, n_90_port_4);
  spice_pullup pullup_3287(dor0_v, dor0_port_4);
  spice_pullup pullup_3286(n_93_v, n_93_port_2);
  spice_pullup pullup_3281(n_83_v, n_83_port_3);
  spice_pullup pullup_3280(n_80_v, n_80_port_3);
  spice_pullup pullup_3283(rdy_v, rdy_port_2);
  spice_pullup pullup_3282(op_T2_ind_x_v, op_T2_ind_x_port_6);
  spice_pullup pullup_3289(n_105_v, n_105_port_3);
  spice_pullup pullup_3288(n_104_v, n_104_port_6);
  spice_pullup pullup_3476(n_397_v, n_397_port_2);
  spice_pullup pullup_4088(op_T0_lda_v, op_T0_lda_port_7);
  spice_pullup pullup_4089(Pout2_v, Pout2_port_2);
  spice_pullup pullup_4082(n_1412_v, n_1412_port_2);
  spice_pullup pullup_4083(n_1413_v, n_1413_port_2);
  spice_pullup pullup_4080(n_1408_v, n_1408_port_2);
  spice_pullup pullup_4081(pd7_clearIR_v, pd7_clearIR_port_4);
  spice_pullup pullup_4086(n_1416_v, n_1416_port_2);
  spice_pullup pullup_4087(op_T0_cld_sed_v, op_T0_cld_sed_port_8);
  spice_pullup pullup_4084(alu3_v, alu3_port_3);
  spice_pullup pullup_4085(dor6_v, dor6_port_4);
  spice_pullup pullup_3348(n_207_v, n_207_port_3);
  spice_pullup pullup_3349(n_208_v, n_208_port_4);
  spice_pullup pullup_3618(n_645_v, n_645_port_3);
  spice_pullup pullup_3619(n_646_v, n_646_port_8);
  spice_pullup pullup_3616(AxB3_v, AxB3_port_6);
  spice_pullup pullup_3617(n_641_v, n_641_port_3);
  spice_pullup pullup_3614(n_637_v, n_637_port_3);
  spice_pullup pullup_3615(n_638_v, n_638_port_2);
  spice_pullup pullup_3612(n_632_v, n_632_port_3);
  spice_pullup pullup_3613(n_636_v, n_636_port_2);
  spice_pullup pullup_3346(op_T2_ADL_ADD_v, op_T2_ADL_ADD_port_3);
  spice_pullup pullup_3347(n_206_v, n_206_port_5);
  spice_pullup pullup_3352(n_213_v, n_213_port_2);
  spice_pullup pullup_3350(n_209_v, n_209_port_4);
  spice_pullup pullup_3605(n_624_v, n_624_port_2);
  spice_pullup pullup_3604(DA_C01_v, DA_C01_port_4);
  spice_pullup pullup_3355(n_218_v, n_218_port_2);
  spice_pullup pullup_3354(n_0_ADL0_v, n_0_ADL0_port_3);
  spice_pullup pullup_3409(n_291_v, n_291_port_3);
  spice_pullup pullup_3408(n_288_v, n_288_port_4);
  spice_pullup pullup_3403(n_282_v, n_282_port_2);
  spice_pullup pullup_3402(op_T4_mem_abs_idx_v, op_T4_mem_abs_idx_port_4);
  spice_pullup pullup_3401(n_280_v, n_280_port_4);
  spice_pullup pullup_3400(n_279_v, n_279_port_4);
  spice_pullup pullup_3407(abh2_v, abh2_port_4);
  spice_pullup pullup_3406(op_T0_tay_ldy_not_idx_v, op_T0_tay_ldy_not_idx_port_7);
  spice_pullup pullup_3405(op_T2_zp_zp_idx_v, op_T2_zp_zp_idx_port_4);
  spice_pullup pullup_3404(n_284_v, n_284_port_2);
  spice_pullup pullup_3769(_DA_ADD1_v, _DA_ADD1_port_5);
  spice_pullup pullup_3362(n_228_v, n_228_port_2);
  spice_pullup pullup_3363(dpc28_0ADH0_v, dpc28_0ADH0_port_2);
  spice_pullup pullup_3360(n_225_v, n_225_port_2);
  spice_pullup pullup_3361(n_227_v, n_227_port_2);
  spice_pullup pullup_3366(n_233_v, n_233_port_2);
  spice_pullup pullup_3367(abl5_v, abl5_port_4);
  spice_pullup pullup_3364(n_231_v, n_231_port_2);
  spice_pullup pullup_3365(n_232_v, n_232_port_4);
  spice_pullup pullup_3368(n_236_v, n_236_port_7);
  spice_pullup pullup_3369(n_238_v, n_238_port_2);
  spice_pullup pullup_3968(n_1223_v, n_1223_port_4);
  spice_pullup pullup_3969(n_1224_v, n_1224_port_2);
  spice_pullup pullup_3960(n_1213_v, n_1213_port_3);
  spice_pullup pullup_3961(n_1214_v, n_1214_port_2);
  spice_pullup pullup_3962(n_1215_v, n_1215_port_5);
  spice_pullup pullup_3963(__AxB7__C67_v, __AxB7__C67_port_3);
  spice_pullup pullup_3964(n_1218_v, n_1218_port_2);
  spice_pullup pullup_3965(n_1219_v, n_1219_port_2);
  spice_pullup pullup_3966(AxB5_v, AxB5_port_6);
  spice_pullup pullup_3967(n_1222_v, n_1222_port_2);
  spice_pullup pullup_4235(n_1694_v, n_1694_port_3);
  spice_pullup pullup_4234(n_1691_v, n_1691_port_7);
  spice_pullup pullup_4237(dpc34_PCLC_v, dpc34_PCLC_port_12);
  spice_pullup pullup_3540(C12_v, C12_port_3);
  spice_pullup pullup_3237(n_3_v, n_3_port_4);
  spice_pullup pullup_3799(n_951_v, n_951_port_3);
  spice_pullup pullup_3798(op_T__cpx_cpy_abs_v, op_T__cpx_cpy_abs_port_8);
  spice_pullup pullup_3793(n_937_v, n_937_port_4);
  spice_pullup pullup_3792(n_936_v, n_936_port_5);
  spice_pullup pullup_3791(n_935_v, n_935_port_2);
  spice_pullup pullup_3790(op_SRS_v, op_SRS_port_6);
  spice_pullup pullup_3797(n_947_v, n_947_port_2);
  spice_pullup pullup_3796(n_946_v, n_946_port_2);
  spice_pullup pullup_3795(n_944_v, n_944_port_3);
  spice_pullup pullup_3794(aluvout_v, aluvout_port_2);
  spice_pullup pullup_3427(n_319_v, n_319_port_2);
  spice_pullup pullup_3426(n_318_v, n_318_port_4);
  spice_pullup pullup_3421(op_T2_jmp_abs_v, op_T2_jmp_abs_port_9);
  spice_pullup pullup_3420(__AxB_4_v, __AxB_4_port_4);
  spice_pullup pullup_3423(n_312_v, n_312_port_3);
  spice_pullup pullup_3422(n_311_v, n_311_port_3);
  spice_pullup pullup_3889(n_1091_v, n_1091_port_3);
  spice_pullup pullup_3888(n_1090_v, n_1090_port_3);
  spice_pullup pullup_3887(n_1089_v, n_1089_port_2);
  spice_pullup pullup_3886(dor4_v, dor4_port_4);
  spice_pullup pullup_3885(n_1087_v, n_1087_port_3);
  spice_pullup pullup_3884(op_T2_pha_v, op_T2_pha_port_9);
  spice_pullup pullup_3883(n_1085_v, n_1085_port_3);
  spice_pullup pullup_3882(n_1084_v, n_1084_port_5);
  spice_pullup pullup_3881(n_1083_v, n_1083_port_4);
  spice_pullup pullup_3880(n_1082_v, n_1082_port_5);
  spice_pullup pullup_3304(n_130_v, n_130_port_2);
  spice_pullup pullup_3305(op_T0_pla_v, op_T0_pla_port_9);
  spice_pullup pullup_3306(n_132_v, n_132_port_2);
  spice_pullup pullup_3307(n_133_v, n_133_port_4);
  spice_pullup pullup_3300(pchp3_v, pchp3_port_2);
  spice_pullup pullup_3301(PD_n_0xx0xx0x_v, PD_n_0xx0xx0x_port_2);
  spice_pullup pullup_3302(n_127_v, n_127_port_4);
  spice_pullup pullup_3303(n_128_v, n_128_port_2);
  spice_pullup pullup_3308(n_134_v, n_134_port_5);
  spice_pullup pullup_3309(n_139_v, n_139_port_2);
  spice_pullup pullup_3942(short_circuit_idx_add_v, short_circuit_idx_add_port_5);
  spice_pullup pullup_3943(n_1187_v, n_1187_port_2);
  spice_pullup pullup_3940(notir2_v, notir2_port_20);
  spice_pullup pullup_3941(n_1184_v, n_1184_port_4);
  spice_pullup pullup_3946(n_0_ADL2_v, n_0_ADL2_port_2);
  spice_pullup pullup_3947(n_1194_v, n_1194_port_3);
  spice_pullup pullup_3944(n_1190_v, n_1190_port_2);
  spice_pullup pullup_3945(n_1192_v, n_1192_port_2);
  spice_pullup pullup_3948(n_1195_v, n_1195_port_3);
  spice_pullup pullup_3949(op_SUMS_v, op_SUMS_port_5);
  spice_pullup pullup_3487(n_423_v, n_423_port_2);
  spice_pullup pullup_3486(abh3_v, abh3_port_4);
  spice_pullup pullup_3447(n_345_v, n_345_port_4);
  spice_pullup pullup_3446(n_344_v, n_344_port_4);
  spice_pullup pullup_3445(x_op_T3_ind_y_v, x_op_T3_ind_y_port_6);
  spice_pullup pullup_3444(op_T4_v, op_T4_port_2);
  spice_pullup pullup_3443(n_340_v, n_340_port_2);
  spice_pullup pullup_3442(ir6_v, ir6_port_43);
  spice_pullup pullup_3448(n_347_v, n_347_port_8);
  spice_pullup pullup_3328(_AxB_6__C56_v, _AxB_6__C56_port_3);
  spice_pullup pullup_3329(n_176_v, n_176_port_3);
  spice_pullup pullup_3326(n_169_v, n_169_port_3);
  spice_pullup pullup_3327(n_172_v, n_172_port_3);
  spice_pullup pullup_3324(op_T0_tax_v, op_T0_tax_port_9);
  spice_pullup pullup_3325(n_168_v, n_168_port_2);
  spice_pullup pullup_3322(n_161_v, n_161_port_4);
  spice_pullup pullup_3323(n_163_v, n_163_port_3);
  spice_pullup pullup_3320(op_T2_stack_access_v, op_T2_stack_access_port_6);
  spice_pullup pullup_3924(x_op_T__adc_sbc_v, x_op_T__adc_sbc_port_6);
  spice_pullup pullup_3925(n_1157_v, n_1157_port_2);
  spice_pullup pullup_3926(n_1159_v, n_1159_port_3);
  spice_pullup pullup_3927(op_clv_v, op_clv_port_8);
  spice_pullup pullup_3920(n_1145_v, n_1145_port_3);
  spice_pullup pullup_3921(alucout_v, alucout_port_3);
  spice_pullup pullup_3922(n_1153_v, n_1153_port_3);
  spice_pullup pullup_3923(n_1154_v, n_1154_port_3);
  spice_pullup pullup_3928(notalucin_v, notalucin_port_4);
  spice_pullup pullup_3929(n_1166_v, n_1166_port_3);
  spice_pullup pullup_3340(_AxB_2__C12_v, _AxB_2__C12_port_3);
  spice_pullup pullup_3341(notir0_v, notir0_port_28);
  spice_pullup pullup_3342(n_196_v, n_196_port_2);
  spice_pullup pullup_3343(n_198_v, n_198_port_3);
  spice_pullup pullup_3344(n_200_v, n_200_port_5);
  spice_pullup pullup_3345(n_201_v, n_201_port_3);
  spice_pullup pullup_3610(n_630_v, n_630_port_3);
  spice_pullup pullup_3611(n_631_v, n_631_port_3);
  spice_pullup pullup_3469(n_386_v, n_386_port_3);
  spice_pullup pullup_3461(n_374_v, n_374_port_2);
  spice_pullup pullup_3460(n_372_v, n_372_port_2);
  spice_pullup pullup_3463(n_378_v, n_378_port_4);
  spice_pullup pullup_3462(abl1_v, abl1_port_4);
  spice_pullup pullup_3465(op_T0_iny_dey_v, op_T0_iny_dey_port_8);
  spice_pullup pullup_3464(dpc36_IPC_v, dpc36_IPC_port_5);
  spice_pullup pullup_3467(n_384_v, n_384_port_6);
  spice_pullup pullup_3466(n_383_v, n_383_port_3);
  spice_pullup pullup_4118(n_1474_v, n_1474_port_2);
  spice_pullup pullup_4119(dasb3_v, dasb3_port_3);
  spice_pullup pullup_4110(pd6_clearIR_v, pd6_clearIR_port_3);
  spice_pullup pullup_4111(n_1462_v, n_1462_port_2);
  spice_pullup pullup_4112(n_1463_v, n_1463_port_4);
  spice_pullup pullup_4114(VEC0_v, VEC0_port_5);
  spice_pullup pullup_4115(op_rol_ror_v, op_rol_ror_port_5);
  spice_pullup pullup_4116(n_1469_v, n_1469_port_2);
  spice_pullup pullup_4117(n_1471_v, n_1471_port_2);
  spice_pullup pullup_3696(op_T5_jsr_v, op_T5_jsr_port_9);
  spice_pullup pullup_3697(ONEBYTE_v, ONEBYTE_port_2);
  spice_pullup pullup_3694(n_774_v, n_774_port_2);
  spice_pullup pullup_3695(abh5_v, abh5_port_4);
  spice_pullup pullup_3692(n_772_v, n_772_port_3);
  spice_pullup pullup_3693(n_773_v, n_773_port_3);
  spice_pullup pullup_3690(n_770_v, n_770_port_3);
  spice_pullup pullup_3691(n_771_v, n_771_port_4);
  spice_pullup pullup_3698(n_779_v, n_779_port_3);
  spice_pullup pullup_3699(n_781_v, n_781_port_9);
  spice_pullup pullup_3908(_C12_v, _C12_port_4);
  spice_pullup pullup_3909(notir3_v, notir3_port_51);
  spice_pullup pullup_3906(p4_v, p4_port_2);
  spice_pullup pullup_3907(n_1120_v, n_1120_port_2);
  spice_pullup pullup_3904(idl6_v, idl6_port_2);
  spice_pullup pullup_3905(n_1117_v, n_1117_port_2);
  spice_pullup pullup_3902(op_T0_clc_sec_v, op_T0_clc_sec_port_8);
  spice_pullup pullup_3903(n_1115_v, n_1115_port_3);
  spice_pullup pullup_3900(n_1111_v, n_1111_port_3);
  spice_pullup pullup_3901(ir4_v, ir4_port_70);
  spice_pullup pullup_4228(n_1677_v, n_1677_port_3);
  spice_pullup pullup_3483(notalucout_v, notalucout_port_4);
  spice_pullup pullup_3482(n_410_v, n_410_port_5);
  spice_pullup pullup_3481(n_409_v, n_409_port_3);
  spice_pullup pullup_3480(n_404_v, n_404_port_5);
  spice_pullup pullup_3484(n_419_v, n_419_port_2);
  spice_pullup pullup_3489(AxB1_v, AxB1_port_6);
  spice_pullup pullup_4132(n_1496_v, n_1496_port_4);
  spice_pullup pullup_4133(n_1497_v, n_1497_port_2);
  spice_pullup pullup_4130(dasb7_v, dasb7_port_3);
  spice_pullup pullup_4131(n_1495_v, n_1495_port_4);
  spice_pullup pullup_4136(abl2_v, abl2_port_4);
  spice_pullup pullup_4137(op_T0_and_v, op_T0_and_port_6);
  spice_pullup pullup_4134(n_1499_v, n_1499_port_3);
  spice_pullup pullup_4135(n_1500_v, n_1500_port_3);
  spice_pullup pullup_4138(_C01_v, _C01_port_3);
  spice_pullup pullup_4139(n_1507_v, n_1507_port_2);
  spice_pullup pullup_3496(n_440_v, n_440_port_10);
  spice_pullup pullup_3713(op_T4_brk_jsr_v, op_T4_brk_jsr_port_8);
  spice_pullup pullup_3712(n_803_v, n_803_port_2);
  spice_pullup pullup_3711(n_800_v, n_800_port_2);
  spice_pullup pullup_3710(n_797_v, n_797_port_2);
  spice_pullup pullup_3717(n_810_v, n_810_port_3);
  spice_pullup pullup_3716(pd1_clearIR_v, pd1_clearIR_port_4);
  spice_pullup pullup_3715(C78_v, C78_port_2);
  spice_pullup pullup_3714(n_807_v, n_807_port_3);
  spice_pullup pullup_3719(n_812_v, n_812_port_3);
  spice_pullup pullup_3718(n_811_v, n_811_port_5);
  spice_pullup pullup_4154(n_1541_v, n_1541_port_4);
  spice_pullup pullup_4155(n_1542_v, n_1542_port_4);
  spice_pullup pullup_4156(x_op_T0_txa_v, x_op_T0_txa_port_9);
  spice_pullup pullup_4157(BRtaken_v, BRtaken_port_4);
  spice_pullup pullup_4150(n_1526_v, n_1526_port_2);
  spice_pullup pullup_4151(n_1531_v, n_1531_port_3);
  spice_pullup pullup_4152(n_1534_v, n_1534_port_4);
  spice_pullup pullup_4153(op_from_x_v, op_from_x_port_6);
  spice_pullup pullup_4158(n_1548_v, n_1548_port_2);
  spice_pullup pullup_4159(n_1549_v, n_1549_port_2);
  spice_pullup pullup_3388(n_262_v, n_262_port_3);
  spice_pullup pullup_3389(dasb5_v, dasb5_port_3);
  spice_pullup pullup_3384(op_T2_idx_x_xy_v, op_T2_idx_x_xy_port_5);
  spice_pullup pullup_3385(op_jsr_v, op_jsr_port_8);
  spice_pullup pullup_3386(n_260_v, n_260_port_3);
  spice_pullup pullup_3387(n_261_v, n_261_port_3);
  spice_pullup pullup_3380(n_254_v, n_254_port_2);
  spice_pullup pullup_3381(n_255_v, n_255_port_2);
  spice_pullup pullup_3382(n_256_v, n_256_port_8);
  spice_pullup pullup_3383(op_T0_tya_v, op_T0_tya_port_9);
  spice_pullup pullup_3528(n_488_v, n_488_port_4);
  spice_pullup pullup_3529(abh7_v, abh7_port_4);
  spice_pullup pullup_3520(n_478_v, n_478_port_2);
  spice_pullup pullup_3521(n_479_v, n_479_port_3);
  spice_pullup pullup_3522(n_480_v, n_480_port_2);
  spice_pullup pullup_3523(n_481_v, n_481_port_4);
  spice_pullup pullup_3524(n_484_v, n_484_port_2);
  spice_pullup pullup_3525(n_485_v, n_485_port_2);
  spice_pullup pullup_3526(__AxBxC_5_v, __AxBxC_5_port_3);
  spice_pullup pullup_3527(op_T2_brk_v, op_T2_brk_port_9);
  spice_pullup pullup_3735(aluanandb1_v, aluanandb1_port_4);
  spice_pullup pullup_3734(_op_branch_bit6_v, _op_branch_bit6_port_4);
  spice_pullup pullup_3737(n_844_v, n_844_port_5);
  spice_pullup pullup_3736(n_842_v, n_842_port_3);
  spice_pullup pullup_3731(n_837_v, n_837_port_2);
  spice_pullup pullup_3730(n_834_v, n_834_port_4);
  spice_pullup pullup_3733(n_839_v, n_839_port_2);
  spice_pullup pullup_3732(n_838_v, n_838_port_2);
  spice_pullup pullup_3739(n_846_v, n_846_port_3);
  spice_pullup pullup_3738(n_845_v, n_845_port_4);
  spice_pullup pullup_4178(n_1588_v, n_1588_port_2);
  spice_pullup pullup_4176(n_1586_v, n_1586_port_2);
  spice_pullup pullup_4177(pd3_clearIR_v, pd3_clearIR_port_4);
  spice_pullup pullup_4174(op_T2_stack_v, op_T2_stack_port_7);
  spice_pullup pullup_4175(n_1585_v, n_1585_port_2);
  spice_pullup pullup_4172(n_1578_v, n_1578_port_2);
  spice_pullup pullup_4173(n_1580_v, n_1580_port_3);
  spice_pullup pullup_4170(n_1575_v, n_1575_port_4);
  spice_pullup pullup_4171(ir3_v, ir3_port_41);
  spice_pullup pullup_3502(x_op_T3_abs_idx_v, x_op_T3_abs_idx_port_4);
  spice_pullup pullup_3503(dasb2_v, dasb2_port_3);
  spice_pullup pullup_3500(n_445_v, n_445_port_4);
  spice_pullup pullup_3501(op_T5_rti_rts_v, op_T5_rti_rts_port_8);
  spice_pullup pullup_3506(n_458_v, n_458_port_2);
  spice_pullup pullup_3507(x_op_T4_ind_y_v, x_op_T4_ind_y_port_7);
  spice_pullup pullup_3504(n_453_v, n_453_port_3);
  spice_pullup pullup_3505(n_457_v, n_457_port_2);
  spice_pullup pullup_3508(n_462_v, n_462_port_3);
  spice_pullup pullup_3509(idl3_v, idl3_port_2);
  spice_pullup pullup_4250(n_1720_v, n_1720_port_4);
  spice_pullup pullup_3757(n_877_v, n_877_port_3);
  spice_pullup pullup_3756(n_876_v, n_876_port_2);
  spice_pullup pullup_3755(n_875_v, n_875_port_3);
  spice_pullup pullup_3754(alu1_v, alu1_port_4);
  spice_pullup pullup_3753(n_871_v, n_871_port_3);
  spice_pullup pullup_3752(idl1_v, idl1_port_2);
  spice_pullup pullup_3751(n_867_v, n_867_port_3);
  spice_pullup pullup_3750(n_862_v, n_862_port_9);
  spice_pullup pullup_3398(n_275_v, n_275_port_3);
  spice_pullup pullup_4190(n_1610_v, n_1610_port_3);
  spice_pullup pullup_4191(op_T4_rts_v, op_T4_rts_port_9);
  spice_pullup pullup_4194(n_1618_v, n_1618_port_4);
  spice_pullup pullup_4195(n_1619_v, n_1619_port_3);
  spice_pullup pullup_4196(n_1621_v, n_1621_port_2);
  spice_pullup pullup_4197(pd0_clearIR_v, pd0_clearIR_port_5);
  spice_pullup pullup_4198(op_T0_eor_v, op_T0_eor_port_6);
  spice_pullup pullup_4199(ir1_v, ir1_port_3);
  spice_pullup pullup_3564(n_550_v, n_550_port_3);
  spice_pullup pullup_3565(n_551_v, n_551_port_2);
  spice_pullup pullup_3566(op_T0_php_pha_v, op_T0_php_pha_port_8);
  spice_pullup pullup_3567(n_553_v, n_553_port_3);
  spice_pullup pullup_3560(n_543_v, n_543_port_3);
  spice_pullup pullup_3561(n_544_v, n_544_port_2);
  spice_pullup pullup_3562(op_shift_v, op_shift_port_4);
  spice_pullup pullup_3563(n_548_v, n_548_port_2);
  spice_pullup pullup_3568(_AxB_0__C0in_v, _AxB_0__C0in_port_3);
  spice_pullup pullup_3569(n_556_v, n_556_port_2);
  spice_pullup pullup_4039(n_1339_v, n_1339_port_2);
  spice_pullup pullup_4038(op_T0_cpx_cpy_inx_iny_v, op_T0_cpx_cpy_inx_iny_port_6);
  spice_pullup pullup_4033(_C78_v, _C78_port_3);
  spice_pullup pullup_4032(op_T__shift_a_v, op_T__shift_a_port_7);
  spice_pullup pullup_4031(n_1323_v, n_1323_port_2);
  spice_pullup pullup_4030(notir7_v, notir7_port_35);
  spice_pullup pullup_4037(n_1335_v, n_1335_port_2);
  spice_pullup pullup_4036(dpc35_PCHC_v, dpc35_PCHC_port_7);
  spice_pullup pullup_4035(ir5_v, ir5_port_33);
  spice_pullup pullup_4034(ir7_v, ir7_port_60);
  spice_pullup pullup_3986(n_1245_v, n_1245_port_2);
  spice_pullup pullup_3987(op_shift_right_v, op_shift_right_port_4);
  spice_pullup pullup_3984(op_T__ora_and_eor_adc_v, op_T__ora_and_eor_adc_port_4);
  spice_pullup pullup_3985(n_1244_v, n_1244_port_2);
  spice_pullup pullup_3982(n_1240_v, n_1240_port_2);
  spice_pullup pullup_3983(AxB7_v, AxB7_port_6);
  spice_pullup pullup_3980(n_1238_v, n_1238_port_2);
  spice_pullup pullup_3981(op_T2_branch_v, op_T2_branch_port_6);
  spice_pullup pullup_3988(abl3_v, abl3_port_4);
  spice_pullup pullup_3989(n_1251_v, n_1251_port_3);
  spice_pullup pullup_3771(n_905_v, n_905_port_2);
  spice_pullup pullup_3770(op_T3_mem_zp_idx_v, op_T3_mem_zp_idx_port_5);
  spice_pullup pullup_3773(_t5_v, _t5_port_10);
  spice_pullup pullup_3772(n_906_v, n_906_port_3);
  spice_pullup pullup_3775(n_913_v, n_913_port_2);
  spice_pullup pullup_3774(alucin_v, alucin_port_2);
  spice_pullup pullup_3777(n_917_v, n_917_port_3);
  spice_pullup pullup_3776(n_916_v, n_916_port_4);
  spice_pullup pullup_3779(n_919_v, n_919_port_4);
  spice_pullup pullup_3778(n_918_v, n_918_port_2);
  spice_pullup pullup_4200(aluanandb0_v, aluanandb0_port_5);
  spice_pullup pullup_4201(n_1629_v, n_1629_port_3);
  spice_pullup pullup_4202(n_1631_v, n_1631_port_2);
  spice_pullup pullup_4203(n_1632_v, n_1632_port_5);
  spice_pullup pullup_4204(dor2_v, dor2_port_4);
  spice_pullup pullup_4205(n_1635_v, n_1635_port_2);
  spice_pullup pullup_4207(n_1638_v, n_1638_port_2);
  spice_pullup pullup_3859(n_1046_v, n_1046_port_2);
  spice_pullup pullup_3855(H1x1_v, H1x1_port_8);
  spice_pullup pullup_3238(op_T0_tay_v, op_T0_tay_port_9);
  spice_pullup pullup_3239(n_5_v, n_5_port_2);
  spice_pullup pullup_3548(n_518_v, n_518_port_3);
  spice_pullup pullup_3549(n_519_v, n_519_port_4);
  spice_pullup pullup_3546(DA_AxB2_v, DA_AxB2_port_3);
  spice_pullup pullup_3547(op_store_v, op_store_port_4);
  spice_pullup pullup_3544(n_513_v, n_513_port_4);
  spice_pullup pullup_3545(n_515_v, n_515_port_3);
  spice_pullup pullup_3542(n_507_v, n_507_port_3);
  spice_pullup pullup_3543(n_510_v, n_510_port_4);
  spice_pullup pullup_3236(op_T5_rts_v, op_T5_rts_port_12);
  spice_pullup pullup_3541(n_506_v, n_506_port_4);
  spice_pullup pullup_4019(idl4_v, idl4_port_2);
  spice_pullup pullup_4018(n_1305_v, n_1305_port_2);
  spice_pullup pullup_4015(n_1301_v, n_1301_port_4);
  spice_pullup pullup_4014(n_1295_v, n_1295_port_3);
  spice_pullup pullup_4017(n_1304_v, n_1304_port_3);
  spice_pullup pullup_4016(n_1303_v, n_1303_port_3);
  spice_pullup pullup_4011(op_T0_cli_sei_v, op_T0_cli_sei_port_8);
  spice_pullup pullup_4010(n_1290_v, n_1290_port_3);
  spice_pullup pullup_4013(PD_1xx000x0_v, PD_1xx000x0_port_6);
  spice_pullup pullup_4012(n_1293_v, n_1293_port_4);
  spice_pullup pullup_3418(n_306_v, n_306_port_2);
  spice_pullup pullup_3419(n_307_v, n_307_port_4);
  spice_pullup pullup_3416(PD_xxx010x1_v, PD_xxx010x1_port_5);
  spice_pullup pullup_4229(n_1682_v, n_1682_port_2);
  spice_pullup pullup_4222(op_T__inx_v, op_T__inx_port_9);
  spice_pullup pullup_4223(op_T__asl_rol_a_v, op_T__asl_rol_a_port_8);
  spice_pullup pullup_4220(n_1660_v, n_1660_port_3);
  spice_pullup pullup_4221(n_1662_v, n_1662_port_3);
  spice_pullup pullup_4226(so_v, so_port_2);
  spice_pullup pullup_4227(n_1676_v, n_1676_port_3);
  spice_pullup pullup_4224(n_1668_v, n_1668_port_2);
  spice_pullup pullup_4225(pd2_clearIR_v, pd2_clearIR_port_6);
  spice_pullup pullup_4077(n_1400_v, n_1400_port_2);
  spice_pullup pullup_4076(n_1399_v, n_1399_port_3);
  spice_pullup pullup_4075(n_1398_v, n_1398_port_6);
  spice_pullup pullup_4074(op_T0_shift_a_v, op_T0_shift_a_port_8);
  spice_pullup pullup_4073(notir5_v, notir5_port_37);
  spice_pullup pullup_4072(n_1392_v, n_1392_port_3);
  spice_pullup pullup_4071(n_1391_v, n_1391_port_3);
  spice_pullup pullup_4070(n_1389_v, n_1389_port_4);
  spice_pullup pullup_4079(n_1402_v, n_1402_port_2);
  spice_pullup pullup_4078(n_1401_v, n_1401_port_2);
  spice_pullup pullup_3267(n_61_v, n_61_port_3);
  spice_pullup pullup_3594(alu4_v, alu4_port_3);
  spice_pullup pullup_3265(op_T3_abs_idx_v, op_T3_abs_idx_port_4);
  spice_pullup pullup_3264(op_lsr_ror_dec_inc_v, op_lsr_ror_dec_inc_port_3);
  spice_pullup pullup_3591(n_602_v, n_602_port_2);
  spice_pullup pullup_3590(n_600_v, n_600_port_4);
  spice_pullup pullup_3260(n_36_v, n_36_port_4);
  spice_pullup pullup_3858(n_1045_v, n_1045_port_4);
  spice_pullup pullup_3850(n_1034_v, n_1034_port_3);
  spice_pullup pullup_3851(_DBE_v, _DBE_port_3);
  spice_pullup pullup_3852(n_1037_v, n_1037_port_3);
  spice_pullup pullup_3853(n_1038_v, n_1038_port_2);
  spice_pullup pullup_3854(n_1039_v, n_1039_port_3);
  spice_pullup pullup_3856(n_1043_v, n_1043_port_2);
  spice_pullup pullup_3857(n_1044_v, n_1044_port_3);
  spice_pullup pullup_3669(n_732_v, n_732_port_4);
  spice_pullup pullup_3668(pclp6_v, pclp6_port_2);
  spice_pullup pullup_3663(n_723_v, n_723_port_4);
  spice_pullup pullup_3662(n_721_v, n_721_port_4);
  spice_pullup pullup_3661(n_720_v, n_720_port_3);
  spice_pullup pullup_3660(n_718_v, n_718_port_2);
  spice_pullup pullup_3667(n_730_v, n_730_port_2);
  spice_pullup pullup_3666(n_728_v, n_728_port_2);
  spice_pullup pullup_3665(n_726_v, n_726_port_5);
  spice_pullup pullup_3664(dpc22__DSA_v, dpc22__DSA_port_3);
  spice_pullup pullup_4248(n_1718_v, n_1718_port_2);
  spice_pullup pullup_4249(n_1719_v, n_1719_port_2);
  spice_pullup pullup_4244(n_1714_v, n_1714_port_2);
  spice_pullup pullup_4245(n_1715_v, n_1715_port_3);
  spice_pullup pullup_4246(n_1716_v, n_1716_port_5);
  spice_pullup pullup_4247(n_1717_v, n_1717_port_8);
  spice_pullup pullup_4240(n_1709_v, n_1709_port_3);
  spice_pullup pullup_4241(op_T__cpx_cpy_imm_zp_v, op_T__cpx_cpy_imm_zp_port_7);
  spice_pullup pullup_4242(n_1711_v, n_1711_port_2);
  spice_pullup pullup_4243(n_1712_v, n_1712_port_4);
  spice_pullup pullup_3588(op_T0_jmp_v, op_T0_jmp_port_8);
  spice_pullup pullup_3589(n_595_v, n_595_port_4);
  spice_pullup pullup_3582(n_583_v, n_583_port_2);
  spice_pullup pullup_3583(n_586_v, n_586_port_3);
  spice_pullup pullup_3580(op_T3_jsr_v, op_T3_jsr_port_9);
  spice_pullup pullup_3581(n_582_v, n_582_port_3);
  spice_pullup pullup_3586(_C67_v, _C67_port_3);
  spice_pullup pullup_3587(n_593_v, n_593_port_2);
  spice_pullup pullup_3584(n_587_v, n_587_port_2);
  spice_pullup pullup_3585(n_588_v, n_588_port_2);
  spice_pullup pullup_3274(n_72_v, n_72_port_4);
  spice_pullup pullup_3275(n_75_v, n_75_port_2);
  spice_pullup pullup_3276(op_T0_dex_v, op_T0_dex_port_9);
  spice_pullup pullup_3277(p6_v, p6_port_2);
  spice_pullup pullup_3270(_AxB_4__C34_v, _AxB_4__C34_port_3);
  spice_pullup pullup_3271(Reset0_v, Reset0_port_5);
  spice_pullup pullup_3273(n_71_v, n_71_port_2);
  spice_pullup pullup_3278(C34_v, C34_port_5);
  spice_pullup pullup_3279(n_79_v, n_79_port_2);
  spice_pullup pullup_4059(n_1375_v, n_1375_port_2);
  spice_pullup pullup_4058(n_1374_v, n_1374_port_4);
  spice_pullup pullup_4051(n_1358_v, n_1358_port_5);
  spice_pullup pullup_4050(n_1357_v, n_1357_port_5);
  spice_pullup pullup_4053(n_1368_v, n_1368_port_4);
  spice_pullup pullup_4052(n_1364_v, n_1364_port_3);
  spice_pullup pullup_4055(p7_v, p7_port_2);
  spice_pullup pullup_4054(n_1369_v, n_1369_port_3);
  spice_pullup pullup_4057(DC34_v, DC34_port_4);
  spice_pullup pullup_4056(n_1371_v, n_1371_port_4);
  spice_pullup pullup_3872(n_1069_v, n_1069_port_3);
  spice_pullup pullup_3873(n_1070_v, n_1070_port_4);
  spice_pullup pullup_3870(idl2_v, idl2_port_2);
  spice_pullup pullup_3871(n_1067_v, n_1067_port_2);
  spice_pullup pullup_3876(n_1075_v, n_1075_port_2);
  spice_pullup pullup_3877(clearIR_v, clearIR_port_9);
  spice_pullup pullup_3874(n_1073_v, n_1073_port_2);
  spice_pullup pullup_3875(op_T0_shift_right_a_v, op_T0_shift_right_a_port_8);
  spice_pullup pullup_3878(pclp2_v, pclp2_port_2);
  spice_pullup pullup_3879(n_1081_v, n_1081_port_3);
  spice_pullup pullup_3649(_DA_ADD2_v, _DA_ADD2_port_3);
  spice_pullup pullup_3648(n_696_v, n_696_port_3);
  spice_pullup pullup_3645(aluaorb0_v, aluaorb0_port_2);
  spice_pullup pullup_3644(n_692_v, n_692_port_4);
  spice_pullup pullup_3647(n_695_v, n_695_port_2);
  spice_pullup pullup_3646(n_694_v, n_694_port_4);
  spice_pullup pullup_3641(n_689_v, n_689_port_2);
  spice_pullup pullup_3640(Pout0_v, Pout0_port_2);
  spice_pullup pullup_3643(op_asl_rol_v, op_asl_rol_port_5);
  spice_pullup pullup_3642(_t4_v, _t4_port_13);
  spice_pullup pullup_3353(DA_AB2_v, DA_AB2_port_3);
  spice_pullup pullup_3351(n_212_v, n_212_port_2);
  spice_pullup pullup_4064(op_T3_jmp_v, op_T3_jmp_port_8);
  spice_pullup pullup_3258(n_34_v, n_34_port_2);
  spice_pullup pullup_3259(n_35_v, n_35_port_4);
  spice_pullup pullup_3256(n_31_v, n_31_port_6);
  spice_pullup pullup_3257(pchp5_v, pchp5_port_2);
  spice_pullup pullup_3254(n_27_v, n_27_port_4);
  spice_pullup pullup_3255(n_29_v, n_29_port_2);
  spice_pullup pullup_3252(n_25_v, n_25_port_3);
  spice_pullup pullup_3253(notir4_v, notir4_port_26);
  spice_pullup pullup_3250(__AxBxC_2_v, __AxBxC_2_port_3);
  spice_pullup pullup_3251(n_23_v, n_23_port_4);
  spice_pullup pullup_4160(n_1552_v, n_1552_port_2);
  spice_pullup pullup_4166(_t3_v, _t3_port_16);
  spice_pullup pullup_3429(n_321_v, n_321_port_3);
  spice_pullup pullup_3428(n_320_v, n_320_port_3);
  spice_pullup pullup_3425(n_317_v, n_317_port_2);
  spice_pullup pullup_3424(alu5_v, alu5_port_4);
  spice_pullup pullup_3814(n_973_v, n_973_port_2);
  spice_pullup pullup_3815(n_975_v, n_975_port_3);
  spice_pullup pullup_3816(n_976_v, n_976_port_4);
  spice_pullup pullup_3817(n_979_v, n_979_port_2);
  spice_pullup pullup_3810(n_966_v, n_966_port_3);
  spice_pullup pullup_3811(nnT2BR_v, nnT2BR_port_10);
  spice_pullup pullup_3812(n_969_v, n_969_port_2);
  spice_pullup pullup_3813(_t2_v, _t2_port_21);
  spice_pullup pullup_3818(n_980_v, n_980_port_2);
  spice_pullup pullup_3819(n_981_v, n_981_port_2);
  spice_pullup pullup_3627(n_664_v, n_664_port_2);
  spice_pullup pullup_3626(n_662_v, n_662_port_2);
  spice_pullup pullup_3625(op_T3_branch_v, op_T3_branch_port_7);
  spice_pullup pullup_3624(n_658_v, n_658_port_3);
  spice_pullup pullup_3623(n_652_v, n_652_port_4);
  spice_pullup pullup_3622(__AxBxC_4_v, __AxBxC_4_port_3);
  spice_pullup pullup_3621(n_649_v, n_649_port_5);
  spice_pullup pullup_3620(n_647_v, n_647_port_5);
  spice_pullup pullup_3629(pd5_clearIR_v, pd5_clearIR_port_3);
  spice_pullup pullup_3628(op_T0_ldy_mem_v, op_T0_ldy_mem_port_7);
  spice_pullup pullup_3485(n_420_v, n_420_port_2);
  spice_pullup pullup_3488(n_424_v, n_424_port_2);
  spice_pullup pullup_4099(n_1440_v, n_1440_port_2);
  spice_pullup pullup_4098(n_1439_v, n_1439_port_2);
  spice_pullup pullup_3272(n_70_v, n_70_port_3);
  spice_pullup pullup_3838(n_1017_v, n_1017_port_2);
  spice_pullup pullup_3839(n_1018_v, n_1018_port_2);
  spice_pullup pullup_3836(n_1010_v, n_1010_port_3);
  spice_pullup pullup_3837(n_1016_v, n_1016_port_2);
  spice_pullup pullup_3834(n_1007_v, n_1007_port_2);
  spice_pullup pullup_3835(dasb1_v, dasb1_port_3);
  spice_pullup pullup_3832(_C23_v, _C23_port_3);
  spice_pullup pullup_3833(op_implied_v, op_implied_port_5);
  spice_pullup pullup_3830(n_998_v, n_998_port_4);
  spice_pullup pullup_3831(n_1002_v, n_1002_port_5);
  spice_pullup pullup_3609(n_629_v, n_629_port_3);
  spice_pullup pullup_3608(n_628_v, n_628_port_4);
  spice_pullup pullup_3359(n_224_v, n_224_port_4);
  spice_pullup pullup_3358(n_221_v, n_221_port_2);
  spice_pullup pullup_3601(n_617_v, n_617_port_3);
  spice_pullup pullup_3600(n_616_v, n_616_port_5);
  spice_pullup pullup_3603(n_620_v, n_620_port_6);
  spice_pullup pullup_3602(n_618_v, n_618_port_4);
  spice_pullup pullup_3357(n_220_v, n_220_port_3);
  spice_pullup pullup_3356(op_T2_mem_zp_v, op_T2_mem_zp_port_5);
  spice_pullup pullup_3607(n_626_v, n_626_port_3);
  spice_pullup pullup_3606(n_625_v, n_625_port_4);
  spice_pullup pullup_3298(n_122_v, n_122_port_2);
  spice_pullup pullup_3299(n_123_v, n_123_port_2);
  spice_pullup pullup_3292(n_110_v, n_110_port_2);
  spice_pullup pullup_3293(n_111_v, n_111_port_2);
  spice_pullup pullup_3290(n_108_v, n_108_port_2);
  spice_pullup pullup_3291(n_109_v, n_109_port_2);
  spice_pullup pullup_3296(n_118_v, n_118_port_2);
  spice_pullup pullup_3297(op_T3_v, op_T3_port_2);
  spice_pullup pullup_3294(pchp1_v, pchp1_port_2);
  spice_pullup pullup_3295(A_B7_v, A_B7_port_2);
  spice_pullup pullup_3379(n_253_v, n_253_port_3);
  spice_pullup pullup_3378(_op_set_C_v, _op_set_C_port_7);
  spice_pullup pullup_3375(op_T0_txs_v, op_T0_txs_port_10);
  spice_pullup pullup_3374(op_ror_v, op_ror_port_5);
  spice_pullup pullup_3377(n_251_v, n_251_port_4);
  spice_pullup pullup_3376(n_249_v, n_249_port_3);
  spice_pullup pullup_3371(n_241_v, n_241_port_3);
  spice_pullup pullup_3370(idl5_v, idl5_port_2);
  spice_pullup pullup_3373(n_243_v, n_243_port_2);
  spice_pullup pullup_3372(n_242_v, n_242_port_3);
  spice_pullup pullup_3979(A_B5_v, A_B5_port_2);
  spice_pullup pullup_3978(op_T0_cpy_iny_v, op_T0_cpy_iny_port_7);
  spice_pullup pullup_3973(op_ANDS_v, op_ANDS_port_6);
  spice_pullup pullup_3972(pclp0_v, pclp0_port_2);
  spice_pullup pullup_3971(op_T0_plp_v, op_T0_plp_port_9);
  spice_pullup pullup_3970(n_1225_v, n_1225_port_5);
  spice_pullup pullup_3977(abl4_v, abl4_port_4);
  spice_pullup pullup_3976(n_1231_v, n_1231_port_2);
  spice_pullup pullup_3975(n_1230_v, n_1230_port_4);
  spice_pullup pullup_3974(n_1229_v, n_1229_port_2);
  spice_pullup pullup_4179(op_T4_jmp_v, op_T4_jmp_port_9);
  spice_pullup pullup_3410(n_293_v, n_293_port_4);
  spice_pullup pullup_3411(__AxB1__C01_v, __AxB1__C01_port_3);
  spice_pullup pullup_3412(n_297_v, n_297_port_3);
  spice_pullup pullup_3413(n_299_v, n_299_port_5);
  spice_pullup pullup_3414(n_300_v, n_300_port_7);
  spice_pullup pullup_3415(op_T__cmp_v, op_T__cmp_port_6);
  spice_pullup pullup_3417(op_T0_bit_v, op_T0_bit_port_8);
  spice_pullup pullup_3436(alu6_v, alu6_port_4);
  spice_pullup pullup_3437(n_332_v, n_332_port_4);
  spice_pullup pullup_3438(DC78_v, DC78_port_4);
  spice_pullup pullup_3439(n_334_v, n_334_port_5);
  spice_pullup pullup_3317(n_154_v, n_154_port_3);
  spice_pullup pullup_3316(n_152_v, n_152_port_5);
  spice_pullup pullup_3315(n_149_v, n_149_port_3);
  spice_pullup pullup_3314(n_146_v, n_146_port_4);
  spice_pullup pullup_3313(op_sta_cmp_v, op_sta_cmp_port_5);
  spice_pullup pullup_3312(aluanorb0_v, aluanorb0_port_6);
  spice_pullup pullup_3311(C45_v, C45_port_4);
  spice_pullup pullup_3310(n_141_v, n_141_port_4);
  spice_pullup pullup_3319(clock2_v, clock2_port_13);
  spice_pullup pullup_3318(aluanorb1_v, aluanorb1_port_5);
  spice_pullup pullup_3261(n_38_v, n_38_port_2);
  spice_pullup pullup_3959(n_1211_v, n_1211_port_8);
  spice_pullup pullup_3958(op_T5_ind_x_v, op_T5_ind_x_port_7);
  spice_pullup pullup_3955(n_1205_v, n_1205_port_4);
  spice_pullup pullup_3954(op_T2_ind_y_v, op_T2_ind_y_port_6);
  spice_pullup pullup_3957(n_1209_v, n_1209_port_3);
  spice_pullup pullup_3956(n_1206_v, n_1206_port_4);
  spice_pullup pullup_3951(n_1199_v, n_1199_port_2);
  spice_pullup pullup_3950(__AxBxC_6_v, __AxBxC_6_port_3);
  spice_pullup pullup_3953(n_1202_v, n_1202_port_3);
  spice_pullup pullup_3952(DBNeg_v, DBNeg_port_3);
  spice_pullup pullup_3788(op_T2_php_pha_v, op_T2_php_pha_port_9);
  spice_pullup pullup_3789(n_933_v, n_933_port_2);
  spice_pullup pullup_3780(n_920_v, n_920_port_2);
  spice_pullup pullup_3781(n_923_v, n_923_port_4);
  spice_pullup pullup_3782(_op_store_v, _op_store_port_3);
  spice_pullup pullup_3783(C1x5Reset_v, C1x5Reset_port_5);
  spice_pullup pullup_3784(n_928_v, n_928_port_2);
  spice_pullup pullup_3785(n_929_v, n_929_port_4);
  spice_pullup pullup_3786(n_930_v, n_930_port_3);
  spice_pullup pullup_3787(n_931_v, n_931_port_2);
  spice_pullup pullup_3432(n_327_v, n_327_port_3);
  spice_pullup pullup_3433(ir0_v, ir0_port_4);
  spice_pullup pullup_3430(op_inc_nop_v, op_inc_nop_port_5);
  spice_pullup pullup_3431(n_326_v, n_326_port_4);
  spice_pullup pullup_3434(n_329_v, n_329_port_3);
  spice_pullup pullup_3435(n_330_v, n_330_port_4);
  spice_pullup pullup_3898(n_1109_v, n_1109_port_5);
  spice_pullup pullup_3899(n_1110_v, n_1110_port_3);
  spice_pullup pullup_3894(n_1099_v, n_1099_port_2);
  spice_pullup pullup_3895(n_1101_v, n_1101_port_2);
  spice_pullup pullup_3896(n_1106_v, n_1106_port_8);
  spice_pullup pullup_3897(n_1107_v, n_1107_port_7);
  spice_pullup pullup_3890(n_1093_v, n_1093_port_2);
  spice_pullup pullup_3891(n_1094_v, n_1094_port_2);
  spice_pullup pullup_3892(abl0_v, abl0_port_4);
  spice_pullup pullup_3893(n_1097_v, n_1097_port_3);
  spice_pullup pullup_3339(n_192_v, n_192_port_4);
  spice_pullup pullup_3338(n_191_v, n_191_port_4);
  spice_pullup pullup_3331(abl6_v, abl6_port_4);
  spice_pullup pullup_3330(n_177_v, n_177_port_2);
  spice_pullup pullup_3333(n_180_v, n_180_port_3);
  spice_pullup pullup_3335(n_184_v, n_184_port_2);
  spice_pullup pullup_3334(n_182_v, n_182_port_7);
  spice_pullup pullup_3337(n_188_v, n_188_port_4);
  spice_pullup pullup_3336(notRnWprepad_v, notRnWprepad_port_6);
  spice_pullup pullup_3937(n_1179_v, n_1179_port_3);
  spice_pullup pullup_3936(n_1178_v, n_1178_port_5);
  spice_pullup pullup_3935(n_1175_v, n_1175_port_3);
  spice_pullup pullup_3934(_op_branch_bit7_v, _op_branch_bit7_port_4);
  spice_pullup pullup_3933(x_op_T0_tya_v, x_op_T0_tya_port_9);
  spice_pullup pullup_3932(n_1170_v, n_1170_port_3);
  spice_pullup pullup_3931(n_1169_v, n_1169_port_3);
  spice_pullup pullup_3939(n_1181_v, n_1181_port_3);
  spice_pullup pullup_3938(n_1180_v, n_1180_port_3);
  spice_pullup pullup_3727(D1x1_v, D1x1_port_5);
  spice_pullup pullup_3454(n_358_v, n_358_port_4);
  spice_pullup pullup_3455(PD_0xx0xx0x_v, PD_0xx0xx0x_port_4);
  spice_pullup pullup_3450(n_351_v, n_351_port_2);
  spice_pullup pullup_3451(op_T4_brk_v, op_T4_brk_port_10);
  spice_pullup pullup_3452(op_T4_abs_idx_v, op_T4_abs_idx_port_4);
  spice_pullup pullup_3453(n_355_v, n_355_port_3);
  spice_pullup pullup_3459(__AxBxC_0_v, __AxBxC_0_port_3);
  spice_pullup pullup_4109(__AxB_6_v, __AxB_6_port_6);
  spice_pullup pullup_4108(n_1458_v, n_1458_port_4);
  spice_pullup pullup_4103(n_1448_v, n_1448_port_2);
  spice_pullup pullup_4102(n_1446_v, n_1446_port_3);
  spice_pullup pullup_4101(Pout1_v, Pout1_port_2);
  spice_pullup pullup_4100(n_1441_v, n_1441_port_2);
  spice_pullup pullup_4107(n_1457_v, n_1457_port_3);
  spice_pullup pullup_4106(n_1455_v, n_1455_port_9);
  spice_pullup pullup_4105(dor5_v, dor5_port_4);
  spice_pullup pullup_4104(n_1449_v, n_1449_port_2);
  spice_pullup pullup_3681(n_755_v, n_755_port_3);
  spice_pullup pullup_3680(n_754_v, n_754_port_4);
  spice_pullup pullup_3683(n_761_v, n_761_port_5);
  spice_pullup pullup_3682(n_757_v, n_757_port_2);
  spice_pullup pullup_3685(n_763_v, n_763_port_2);
  spice_pullup pullup_3684(n_762_v, n_762_port_3);
  spice_pullup pullup_3687(alu7_v, alu7_port_3);
  spice_pullup pullup_3686(op_jmp_v, op_jmp_port_7);
  spice_pullup pullup_3689(n_769_v, n_769_port_4);
  spice_pullup pullup_3688(n_767_v, n_767_port_3);
  spice_pullup pullup_3919(DA_C45_v, DA_C45_port_3);
  spice_pullup pullup_3918(abh4_v, abh4_port_4);
  spice_pullup pullup_3911(n_1130_v, n_1130_port_7);
  spice_pullup pullup_3910(n_1129_v, n_1129_port_4);
  spice_pullup pullup_3913(_VEC_v, _VEC_port_5);
  spice_pullup pullup_3912(n_1133_v, n_1133_port_3);
  spice_pullup pullup_3915(n_1137_v, n_1137_port_2);
  spice_pullup pullup_3914(n_1135_v, n_1135_port_3);
  spice_pullup pullup_3917(n_1141_v, n_1141_port_2);
  spice_pullup pullup_3916(n_1138_v, n_1138_port_2);
  spice_pullup pullup_3332(op_T0_txa_v, op_T0_txa_port_9);
  spice_pullup pullup_3477(n_400_v, n_400_port_3);
  spice_pullup pullup_3474(n_392_v, n_392_port_3);
  spice_pullup pullup_3475(n_396_v, n_396_port_2);
  spice_pullup pullup_3472(n_390_v, n_390_port_2);
  spice_pullup pullup_3473(idl7_v, idl7_port_2);
  spice_pullup pullup_3470(n_388_v, n_388_port_5);
  spice_pullup pullup_3471(n_389_v, n_389_port_4);
  spice_pullup pullup_4129(n_1492_v, n_1492_port_3);
  spice_pullup pullup_4125(n_1486_v, n_1486_port_3);
  spice_pullup pullup_4124(n_1484_v, n_1484_port_2);
  spice_pullup pullup_4127(n_1488_v, n_1488_port_3);
  spice_pullup pullup_4126(op_T3_plp_pla_v, op_T3_plp_pla_port_8);
  spice_pullup pullup_4121(op_T0_brk_rti_v, op_T0_brk_rti_port_8);
  spice_pullup pullup_4120(x_op_T0_bit_v, x_op_T0_bit_port_8);
  spice_pullup pullup_4123(op_T__iny_dey_v, op_T__iny_dey_port_8);
  spice_pullup pullup_4122(VEC1_v, VEC1_port_4);
  spice_pullup pullup_3441(n_336_v, n_336_port_6);
  spice_pullup pullup_3440(n_335_v, n_335_port_8);
  spice_pullup pullup_3449(n_350_v, n_350_port_4);
  spice_pullup pullup_3490(_C56_v, _C56_port_4);
  spice_pullup pullup_3491(n_428_v, n_428_port_3);
  spice_pullup pullup_3492(n_432_v, n_432_port_3);
  spice_pullup pullup_3493(op_rmw_v, op_rmw_port_2);
  spice_pullup pullup_3494(n_436_v, n_436_port_3);
  spice_pullup pullup_3495(Pout3_v, Pout3_port_4);
  spice_pullup pullup_3497(n_441_v, n_441_port_2);
  spice_pullup pullup_3498(n_442_v, n_442_port_2);
  spice_pullup pullup_3499(dor3_v, dor3_port_4);
  spice_pullup pullup_4147(n_1523_v, n_1523_port_3);
  spice_pullup pullup_4146(n_1521_v, n_1521_port_2);
  spice_pullup pullup_4145(op_plp_pla_v, op_plp_pla_port_7);
  spice_pullup pullup_4144(n_1519_v, n_1519_port_2);
  spice_pullup pullup_4143(n_1518_v, n_1518_port_2);
  spice_pullup pullup_4142(n_1517_v, n_1517_port_3);
  spice_pullup pullup_4141(op_T2_abs_y_v, op_T2_abs_y_port_6);
  spice_pullup pullup_4140(n_1511_v, n_1511_port_2);
  spice_pullup pullup_4149(__AxB_0_v, __AxB_0_port_4);
  spice_pullup pullup_4148(op_T2_ind_v, op_T2_ind_port_5);
  spice_pullup pullup_3399(n_278_v, n_278_port_2);
  spice_pullup pullup_3397(__AxBxC_3_v, __AxBxC_3_port_3);
  spice_pullup pullup_3396(op_T2_abs_access_v, op_T2_abs_access_port_6);
  spice_pullup pullup_3395(n_272_v, n_272_port_8);
  spice_pullup pullup_3394(op_T0_jsr_v, op_T0_jsr_port_10);
  spice_pullup pullup_3393(n_270_v, n_270_port_6);
  spice_pullup pullup_3392(n_269_v, n_269_port_3);
  spice_pullup pullup_3391(n_267_v, n_267_port_4);
  spice_pullup pullup_3390(n_264_v, n_264_port_6);
  spice_pullup pullup_3539(n_504_v, n_504_port_2);
  spice_pullup pullup_3538(n_503_v, n_503_port_2);
  spice_pullup pullup_3533(n_494_v, n_494_port_2);
  spice_pullup pullup_3532(op_T4_ind_y_v, op_T4_ind_y_port_6);
  spice_pullup pullup_3531(n_491_v, n_491_port_2);
  spice_pullup pullup_3530(n_490_v, n_490_port_2);
  spice_pullup pullup_3537(n_501_v, n_501_port_4);
  spice_pullup pullup_3536(C56_v, C56_port_3);
  spice_pullup pullup_3535(n_499_v, n_499_port_3);
  spice_pullup pullup_3534(n_496_v, n_496_port_2);
  spice_pullup pullup_3930(op_T5_ind_y_v, op_T5_ind_y_port_6);
  spice_pullup pullup_3759(n_880_v, n_880_port_2);
  spice_pullup pullup_3758(fetch_v, fetch_port_11);
  spice_pullup pullup_3700(n_782_v, n_782_port_2);
  spice_pullup pullup_3701(n_783_v, n_783_port_4);
  spice_pullup pullup_3702(op_T5_rti_v, op_T5_rti_port_10);
  spice_pullup pullup_3703(op_T__dex_v, op_T__dex_port_9);
  spice_pullup pullup_3704(op_T0_sbc_v, op_T0_sbc_port_8);
  spice_pullup pullup_3705(op_T2_v, op_T2_port_2);
  spice_pullup pullup_3706(n_789_v, n_789_port_2);
  spice_pullup pullup_3707(n_790_v, n_790_port_5);
  spice_pullup pullup_3708(op_push_pull_v, op_push_pull_port_7);
  spice_pullup pullup_3709(n_795_v, n_795_port_2);
  spice_pullup pullup_4169(n_1573_v, n_1573_port_2);
  spice_pullup pullup_4168(_C45_v, _C45_port_4);
  spice_pullup pullup_4161(op_brk_rti_v, op_brk_rti_port_7);
  spice_pullup pullup_4163(n_1561_v, n_1561_port_2);
  spice_pullup pullup_4162(n_1560_v, n_1560_port_4);
  spice_pullup pullup_4165(n_1566_v, n_1566_port_3);
  spice_pullup pullup_4164(op_xy_v, op_xy_port_5);
  spice_pullup pullup_4167(x_op_T4_rti_v, x_op_T4_rti_port_9);
  spice_pullup pullup_3519(n_477_v, n_477_port_4);
  spice_pullup pullup_3518(n_476_v, n_476_port_4);
  spice_pullup pullup_3515(n_472_v, n_472_port_3);
  spice_pullup pullup_3514(n_470_v, n_470_port_3);
  spice_pullup pullup_3517(n_474_v, n_474_port_3);
  spice_pullup pullup_3516(n_473_v, n_473_port_2);
  spice_pullup pullup_3511(n_466_v, n_466_port_4);
  spice_pullup pullup_3510(n_465_v, n_465_port_2);
  spice_pullup pullup_3513(n_468_v, n_468_port_3);
  spice_pullup pullup_3512(n_467_v, n_467_port_4);
  spice_pullup pullup_4192(n_1613_v, n_1613_port_4);
  spice_pullup pullup_3728(n_830_v, n_830_port_4);
  spice_pullup pullup_3729(n_831_v, n_831_port_4);
  spice_pullup pullup_3722(__AxB5__C45_v, __AxB5__C45_port_3);
  spice_pullup pullup_3723(n_818_v, n_818_port_4);
  spice_pullup pullup_3720(n_813_v, n_813_port_3);
  spice_pullup pullup_3721(n_815_v, n_815_port_2);
  spice_pullup pullup_3726(n_824_v, n_824_port_5);
  spice_pullup pullup_3724(n_819_v, n_819_port_4);
  spice_pullup pullup_3725(op_T__adc_sbc_v, op_T__adc_sbc_port_5);
  spice_pullup pullup_3457(n_368_v, n_368_port_7);
  spice_pullup pullup_3458(op_T5_brk_v, op_T5_brk_port_10);
  spice_pullup pullup_4183(n_1595_v, n_1595_port_2);
  spice_pullup pullup_4182(n_1594_v, n_1594_port_2);
  spice_pullup pullup_4181(n_1593_v, n_1593_port_3);
  spice_pullup pullup_4180(n_1592_v, n_1592_port_4);
  spice_pullup pullup_4187(n_1600_v, n_1600_port_2);
  spice_pullup pullup_4186(n_1599_v, n_1599_port_3);
  spice_pullup pullup_4185(idl0_v, idl0_port_2);
  spice_pullup pullup_4184(n_1596_v, n_1596_port_3);
  spice_pullup pullup_4189(n_1605_v, n_1605_port_3);
  spice_pullup pullup_4188(op_sty_cpy_mem_v, op_sty_cpy_mem_port_7);
  spice_pullup pullup_3577(n_572_v, n_572_port_3);
  spice_pullup pullup_3576(n_571_v, n_571_port_2);
  spice_pullup pullup_3575(n_570_v, n_570_port_5);
  spice_pullup pullup_3574(n_568_v, n_568_port_2);
  spice_pullup pullup_3573(n_567_v, n_567_port_4);
  spice_pullup pullup_3572(n_566_v, n_566_port_4);
  spice_pullup pullup_3571(n_565_v, n_565_port_2);
  spice_pullup pullup_3570(n_564_v, n_564_port_3);
  spice_pullup pullup_3579(n_578_v, n_578_port_3);
  spice_pullup pullup_3578(op_T0_adc_sbc_v, op_T0_adc_sbc_port_6);
  spice_pullup pullup_3321(n_160_v, n_160_port_3);
  spice_pullup pullup_3991(n_1255_v, n_1255_port_2);
  spice_pullup pullup_3990(n_1253_v, n_1253_port_5);
  spice_pullup pullup_3993(n_1257_v, n_1257_port_5);
  spice_pullup pullup_3992(n_1256_v, n_1256_port_2);
  spice_pullup pullup_3995(op_T4_ind_x_v, op_T4_ind_x_port_7);
  spice_pullup pullup_3994(n_1258_v, n_1258_port_7);
  spice_pullup pullup_3997(n_1262_v, n_1262_port_3);
  spice_pullup pullup_3996(n_1260_v, n_1260_port_3);
  spice_pullup pullup_3999(n_1267_v, n_1267_port_2);
  spice_pullup pullup_3998(n_1265_v, n_1265_port_3);
  spice_pullup pullup_3748(__AxB3__C23_v, __AxB3__C23_port_3);
  spice_pullup pullup_3749(n_861_v, n_861_port_2);
  spice_pullup pullup_3744(n_852_v, n_852_port_3);
  spice_pullup pullup_3745(n_853_v, n_853_port_3);
  spice_pullup pullup_3746(n_854_v, n_854_port_4);
  spice_pullup pullup_3747(op_rti_rts_v, op_rti_rts_port_9);
  spice_pullup pullup_3740(n_847_v, n_847_port_2);
  spice_pullup pullup_3741(n_849_v, n_849_port_2);
  spice_pullup pullup_3742(n_850_v, n_850_port_3);
  spice_pullup pullup_3743(_TWOCYCLE_v, _TWOCYCLE_port_4);
  spice_pullup pullup_4213(n_1647_v, n_1647_port_4);
  spice_pullup pullup_4212(op_T__bit_v, op_T__bit_port_9);
  spice_pullup pullup_4211(n_1643_v, n_1643_port_4);
  spice_pullup pullup_4210(n_1642_v, n_1642_port_2);
  spice_pullup pullup_4215(n_1650_v, n_1650_port_2);
  spice_pullup pullup_4214(n_1649_v, n_1649_port_11);
  spice_pullup pullup_3559(pd4_clearIR_v, pd4_clearIR_port_6);
  spice_pullup pullup_3558(n_538_v, n_538_port_2);
  spice_pullup pullup_3551(n_523_v, n_523_port_4);
  spice_pullup pullup_3550(op_ORS_v, op_ORS_port_3);
  spice_pullup pullup_3553(xx_op_T5_jsr_v, xx_op_T5_jsr_port_9);
  spice_pullup pullup_3552(n_525_v, n_525_port_4);
  spice_pullup pullup_3555(__AxBxC_7_v, __AxBxC_7_port_3);
  spice_pullup pullup_3554(n_531_v, n_531_port_3);
  spice_pullup pullup_3557(pchp7_v, pchp7_port_2);
  spice_pullup pullup_3556(n_533_v, n_533_port_2);
  spice_pullup pullup_4028(n_1318_v, n_1318_port_5);
  spice_pullup pullup_4029(n_1319_v, n_1319_port_2);
  spice_pullup pullup_4020(notaluvout_v, notaluvout_port_3);
  spice_pullup pullup_4021(n_1309_v, n_1309_port_2);
  spice_pullup pullup_4022(op_T4_rti_v, op_T4_rti_port_9);
  spice_pullup pullup_4023(n_1312_v, n_1312_port_3);
  spice_pullup pullup_4024(A_B3_v, A_B3_port_2);
  spice_pullup pullup_4025(C67_v, C67_port_6);
  spice_pullup pullup_4026(n_1315_v, n_1315_port_3);
  spice_pullup pullup_4027(n_1316_v, n_1316_port_5);
  spice_pullup pullup_3766(n_890_v, n_890_port_2);
  spice_pullup pullup_3767(notir6_v, notir6_port_39);
  spice_pullup pullup_3764(n_888_v, n_888_port_2);
  spice_pullup pullup_3765(n_889_v, n_889_port_2);
  spice_pullup pullup_3762(n_884_v, n_884_port_2);
  spice_pullup pullup_3763(n_885_v, n_885_port_2);
  spice_pullup pullup_3760(n_882_v, n_882_port_3);
  spice_pullup pullup_3761(n_883_v, n_883_port_2);
  spice_pullup pullup_3768(n_896_v, n_896_port_2);
  spice_pullup pullup_4233(op_EORS_v, op_EORS_port_3);
  spice_pullup pullup_4232(n_1688_v, n_1688_port_2);
  spice_pullup pullup_4239(n_1708_v, n_1708_port_4);
  spice_pullup pullup_4238(n_1705_v, n_1705_port_3);
  spice_pullup pullup_4217(n_1655_v, n_1655_port_2);
  spice_pullup pullup_4216(n_1654_v, n_1654_port_4);
  spice_pullup pullup_4219(op_T0_cpx_inx_v, op_T0_cpx_inx_port_7);
  spice_pullup pullup_4218(n_1657_v, n_1657_port_2);
  spice_pullup pullup_4002(n_1271_v, n_1271_port_2);
  spice_pullup pullup_4003(op_T0_v, op_T0_port_2);
  spice_pullup pullup_4000(_DBZ_v, _DBZ_port_2);
  spice_pullup pullup_4001(n_1270_v, n_1270_port_4);
  spice_pullup pullup_4006(n_1281_v, n_1281_port_2);
  spice_pullup pullup_4007(C01_v, C01_port_4);
  spice_pullup pullup_4004(n_1275_v, n_1275_port_4);
  spice_pullup pullup_4005(n_1277_v, n_1277_port_3);
  spice_pullup pullup_4008(n_1286_v, n_1286_port_3);
  spice_pullup pullup_4009(n_1289_v, n_1289_port_2);
  spice_pullup pullup_3849(n_1033_v, n_1033_port_2);
  spice_pullup pullup_3848(NMIP_v, NMIP_port_4);
  spice_pullup pullup_3843(n_1024_v, n_1024_port_3);
  spice_pullup pullup_3842(C23_v, C23_port_4);
  spice_pullup pullup_3841(A_B1_v, A_B1_port_2);
  spice_pullup pullup_3840(PD_xxxx10x0_v, PD_xxxx10x0_port_5);
  spice_pullup pullup_3847(op_T3_stack_bit_jmp_v, op_T3_stack_bit_jmp_port_5);
  spice_pullup pullup_3846(n_1028_v, n_1028_port_2);
  spice_pullup pullup_3845(n_1026_v, n_1026_port_3);
  spice_pullup pullup_3844(n_1025_v, n_1025_port_2);
  spice_pullup pullup_4253(n_1724_v, n_1724_port_3);
  spice_pullup pullup_4252(n_1722_v, n_1722_port_4);
  spice_pullup pullup_4251(op_branch_done_v, op_branch_done_port_8);
  spice_pullup pullup_3595(op_T3_mem_abs_v, op_T3_mem_abs_port_5);
  spice_pullup pullup_3266(op_T3_ind_y_v, op_T3_ind_y_port_6);
  spice_pullup pullup_3597(n_609_v, n_609_port_4);
  spice_pullup pullup_3596(n_608_v, n_608_port_2);
  spice_pullup pullup_3263(n_46_v, n_46_port_3);
  spice_pullup pullup_3262(pclp4_v, pclp4_port_2);
  spice_pullup pullup_3593(n_604_v, n_604_port_10);
  spice_pullup pullup_3592(n_603_v, n_603_port_2);
  spice_pullup pullup_3599(n_613_v, n_613_port_4);
  spice_pullup pullup_3598(n_611_v, n_611_port_4);
  spice_pullup pullup_3269(dor7_v, dor7_port_4);
  spice_pullup pullup_3268(n_62_v, n_62_port_2);
  spice_pullup pullup_4065(brk_done_v, brk_done_port_9);
  spice_pullup pullup_4066(n_1383_v, n_1383_port_2);
  spice_pullup pullup_4067(ir2_v, ir2_port_72);
  spice_pullup pullup_4060(n_1376_v, n_1376_port_2);
  spice_pullup pullup_4061(n_1377_v, n_1377_port_2);
  spice_pullup pullup_4062(n_1379_v, n_1379_port_2);
  spice_pullup pullup_4063(n_1380_v, n_1380_port_4);
  spice_pullup pullup_4068(op_T5_mem_ind_idx_v, op_T5_mem_ind_idx_port_5);
  spice_pullup pullup_4069(n_1386_v, n_1386_port_2);
  spice_pullup pullup_3468(n_385_v, n_385_port_3);
  spice_pullup pullup_4128(n_1491_v, n_1491_port_3);
  spice_pullup pullup_4113(n_1464_v, n_1464_port_7);
  spice_pullup pullup_3869(n_1065_v, n_1065_port_2);
  spice_pullup pullup_3868(n_1063_v, n_1063_port_5);
  spice_pullup pullup_3865(n_1055_v, n_1055_port_3);
  spice_pullup pullup_3864(n_1054_v, n_1054_port_2);
  spice_pullup pullup_3867(op_T2_abs_v, op_T2_abs_port_5);
  spice_pullup pullup_3866(n_1056_v, n_1056_port_2);
  spice_pullup pullup_3861(_op_branch_done_v, _op_branch_done_port_2);
  spice_pullup pullup_3860(n_1047_v, n_1047_port_2);
  spice_pullup pullup_3863(x_op_jmp_v, x_op_jmp_port_8);
  spice_pullup pullup_3862(x_op_push_pull_v, x_op_push_pull_port_6);
  spice_pullup pullup_3678(op_T2_php_v, op_T2_php_port_9);
  spice_pullup pullup_3679(n_753_v, n_753_port_4);
  spice_pullup pullup_3670(n_733_v, n_733_port_3);
  spice_pullup pullup_3671(n_735_v, n_735_port_3);
  spice_pullup pullup_3672(n_739_v, n_739_port_4);
  spice_pullup pullup_3673(n_743_v, n_743_port_5);
  spice_pullup pullup_3674(DBZ_v, DBZ_port_9);
  spice_pullup pullup_3675(dor1_v, dor1_port_4);
  spice_pullup pullup_3676(n_747_v, n_747_port_3);
  spice_pullup pullup_3677(n_748_v, n_748_port_3);
  spice_pullup pullup_3456(n_366_v, n_366_port_3);
  spice_pullup pullup_3249(n_21_v, n_21_port_4);
  spice_pullup pullup_3248(n_20_v, n_20_port_3);
  spice_pullup pullup_3241(n_8_v, n_8_port_4);
  spice_pullup pullup_3240(n_6_v, n_6_port_4);
  spice_pullup pullup_3243(n_11_v, n_11_port_6);
  spice_pullup pullup_3242(n_10_v, n_10_port_4);
  spice_pullup pullup_3245(n_16_v, n_16_port_5);
  spice_pullup pullup_3244(n_14_v, n_14_port_4);
  spice_pullup pullup_3247(n_19_v, n_19_port_3);
  spice_pullup pullup_3246(n_17_v, n_17_port_5);
  spice_pullup pullup_4048(op_T0_cmp_v, op_T0_cmp_port_6);
  spice_pullup pullup_4049(n_1356_v, n_1356_port_2);
  spice_pullup pullup_4046(INTG_v, INTG_port_4);
  spice_pullup pullup_4047(_WR_v, _WR_port_7);
  spice_pullup pullup_4044(n_1346_v, n_1346_port_3);
  spice_pullup pullup_4045(n_1347_v, n_1347_port_7);
  spice_pullup pullup_4042(n_1344_v, n_1344_port_4);
  spice_pullup pullup_4043(n_1345_v, n_1345_port_5);
  spice_pullup pullup_4040(op_T0_acc_v, op_T0_acc_port_3);
  spice_pullup pullup_4041(n_1343_v, n_1343_port_3);
  spice_pullup pullup_4096(n_1433_v, n_1433_port_4);
  spice_pullup pullup_4090(n_1423_v, n_1423_port_3);
  spice_pullup pullup_4092(n_1427_v, n_1427_port_3);
  spice_pullup pullup_3807(n_962_v, n_962_port_2);
  spice_pullup pullup_3806(n_961_v, n_961_port_2);
  spice_pullup pullup_3805(n_959_v, n_959_port_4);
  spice_pullup pullup_3804(n_958_v, n_958_port_3);
  spice_pullup pullup_3803(n_956_v, n_956_port_2);
  spice_pullup pullup_3802(n_954_v, n_954_port_4);
  spice_pullup pullup_3801(n_953_v, n_953_port_2);
  spice_pullup pullup_3800(n_952_v, n_952_port_3);
  spice_pullup pullup_3809(__AxBxC_1_v, __AxBxC_1_port_3);
  spice_pullup pullup_3808(n_964_v, n_964_port_4);
  spice_pullup pullup_3652(notir1_v, notir1_port_23);
  spice_pullup pullup_3653(n_708_v, n_708_port_2);
  spice_pullup pullup_3650(n_700_v, n_700_port_3);
  spice_pullup pullup_3651(__AxB_2_v, __AxB_2_port_4);
  spice_pullup pullup_3656(abh1_v, abh1_port_4);
  spice_pullup pullup_3657(n_714_v, n_714_port_2);
  spice_pullup pullup_3654(n_709_v, n_709_port_2);
  spice_pullup pullup_3655(op_T2_jsr_v, op_T2_jsr_port_11);
  spice_pullup pullup_3658(n_715_v, n_715_port_3);
  spice_pullup pullup_3659(n_717_v, n_717_port_4);
  spice_pullup pullup_4095(x_op_T3_plp_pla_v, x_op_T3_plp_pla_port_8);
  spice_pullup pullup_4094(abh0_v, abh0_port_4);
  spice_pullup pullup_4097(n_1434_v, n_1434_port_2);
  spice_pullup pullup_4091(_C34_v, _C34_port_5);
  spice_pullup pullup_4093(op_T3_ind_x_v, op_T3_ind_x_port_7);
  spice_pullup pullup_4206(alu2_v, alu2_port_4);
  spice_pullup pullup_4208(n_1640_v, n_1640_port_2);
  spice_pullup pullup_4209(n_1641_v, n_1641_port_2);
  spice_pullup pullup_4193(n_1614_v, n_1614_port_4);
  spice_pullup pullup_3829(abh6_v, abh6_port_4);
  spice_pullup pullup_3828(irline3_v, irline3_port_64);
  spice_pullup pullup_3821(op_T0_ldx_tax_tsx_v, op_T0_ldx_tax_tsx_port_6);
  spice_pullup pullup_3820(n_983_v, n_983_port_2);
  spice_pullup pullup_3823(n_987_v, n_987_port_2);
  spice_pullup pullup_3822(n_986_v, n_986_port_2);
  spice_pullup pullup_3825(n_990_v, n_990_port_3);
  spice_pullup pullup_3824(n_988_v, n_988_port_3);
  spice_pullup pullup_3827(n_995_v, n_995_port_2);
  spice_pullup pullup_3826(n_992_v, n_992_port_2);
  spice_pullup pullup_4236(n_1697_v, n_1697_port_2);
  spice_pullup pullup_4231(n_1687_v, n_1687_port_2);
  spice_pullup pullup_4230(n_1684_v, n_1684_port_2);
  spice_pullup pullup_3634(op_T3_abs_idx_ind_v, op_T3_abs_idx_ind_port_4);
  spice_pullup pullup_3635(n_678_v, n_678_port_4);
  spice_pullup pullup_3636(dasb6_v, dasb6_port_3);
  spice_pullup pullup_3637(n_681_v, n_681_port_6);
  spice_pullup pullup_3630(n_669_v, n_669_port_3);
  spice_pullup pullup_3631(n_670_v, n_670_port_3);
  spice_pullup pullup_3632(n_673_v, n_673_port_2);
  spice_pullup pullup_3633(n_674_v, n_674_port_2);
  spice_pullup pullup_3638(op_T0_tsx_v, op_T0_tsx_port_9);
  spice_pullup pullup_3639(n_0_ADL1_v, n_0_ADL1_port_2);
  spice_pullup pullup_3478(alu0_v, alu0_port_3);
  spice_pullup pullup_3479(op_T0_ora_v, op_T0_ora_port_6);

  spice_latch latch_5130(eclk,ereset, ~cclk_v[`W-1], ~n_1101_v[`W-1], n_190_v);
  spice_latch latch_5131(eclk,ereset, ~cclk_v[`W-1], ~n_1110_v[`W-1], pipeUNK01_v);
  spice_latch latch_5132(eclk,ereset, ~cp1_v[`W-1], ~n_533_v[`W-1], n_599_v);
  spice_latch latch_5133(eclk,ereset, ~cp1_v[`W-1], ~n_920_v[`W-1], n_785_v);
  spice_latch latch_5134(eclk,ereset, ~cclk_v[`W-1], ~VEC1_v[`W-1], n_1452_v);
  spice_latch latch_5135(eclk,ereset, ~cclk_v[`W-1], ~n_896_v[`W-1], notidl3_v);
  spice_latch latch_5138(eclk,ereset, ~cclk_v[`W-1], ~n_1187_v[`W-1], nots6_v);
  spice_latch latch_5109(eclk,ereset, ~cclk_v[`W-1], ~n_722_v[`W-1], notalu6_v);
  spice_latch latch_5107(eclk,ereset, ~cp1_v[`W-1], ~n_566_v[`W-1], p1_v);
  spice_latch latch_5106(eclk,ereset, ~cp1_v[`W-1], ~notRnWprepad_v[`W-1], n_1579_v);
  spice_latch latch_5045(eclk,ereset, ~cclk_v[`W-1], ~n_440_v[`W-1], pipeUNK39_v);
  spice_latch latch_5047(eclk,ereset, ~cp1_v[`W-1], ~n_1526_v[`W-1], n_1450_v);
  spice_latch latch_4972(eclk,ereset, ~cclk_v[`W-1], ~n_862_v[`W-1], pipeT_SYNC_v);
  spice_latch latch_5088(eclk,ereset, ~cp1_v[`W-1], ~n_1497_v[`W-1], n_653_v);
  spice_latch latch_5089(eclk,ereset, ~cclk_v[`W-1], ~n_616_v[`W-1], n_460_v);
  spice_latch latch_5084(eclk,ereset, ~cclk_v[`W-1], ~n_1281_v[`W-1], pd3_v);
  spice_latch latch_5085(eclk,ereset, ~cclk_v[`W-1], ~n_1588_v[`W-1], pd5_v);
  spice_latch latch_5086(eclk,ereset, ~cclk_v[`W-1], ~n_1075_v[`W-1], pd4_v);
  spice_latch latch_5087(eclk,ereset, ~cclk_v[`W-1], ~n_1638_v[`W-1], notidl6_v);
  spice_latch latch_5080(eclk,ereset, ~cclk_v[`W-1], ~notaluoutmux0_v[`W-1], notalu0_v);
  spice_latch latch_5081(eclk,ereset, ~cclk_v[`W-1], ~n_296_v[`W-1], notalu4_v);
  spice_latch latch_5082(eclk,ereset, ~cclk_v[`W-1], ~n_340_v[`W-1], pipeUNK12_v);
  spice_latch latch_5083(eclk,ereset, ~cp1_v[`W-1], ~notRnWprepad_v[`W-1], n_759_v);
  spice_latch latch_5136(eclk,ereset, ~cp1_v[`W-1], ~n_720_v[`W-1], n_1338_v);
  spice_latch latch_5137(eclk,ereset, ~cclk_v[`W-1], ~n_1229_v[`W-1], pchp0_v);
  spice_latch latch_5139(eclk,ereset, ~cp1_v[`W-1], ~n_1082_v[`W-1], p0_v);
  spice_latch latch_5054(eclk,ereset, ~cclk_v[`W-1], ~n_34_v[`W-1], nots3_v);
  spice_latch latch_4959(eclk,ereset, ~cclk_v[`W-1], ~n_1194_v[`W-1], pipeUNK04_v);
  spice_latch latch_4958(eclk,ereset, ~cclk_v[`W-1], ~n_1106_v[`W-1], n_1404_v);
  spice_latch latch_4955(eclk,ereset, ~cp1_v[`W-1], ~n_1275_v[`W-1], n_1581_v);
  spice_latch latch_4954(eclk,ereset, ~cclk_v[`W-1], ~n_718_v[`W-1], notidl0_v);
  spice_latch latch_4957(eclk,ereset, ~cclk_v[`W-1], ~n_1391_v[`W-1], pipeUNK15_v);
  spice_latch latch_4956(eclk,ereset, ~cp1_v[`W-1], ~D1x1_v[`W-1], n_1472_v);
  spice_latch latch_4951(eclk,ereset, ~cclk_v[`W-1], ~n_548_v[`W-1], nots7_v);
  spice_latch latch_4950(eclk,ereset, ~cclk_v[`W-1], ~n_695_v[`W-1], n_1341_v);
  spice_latch latch_4953(eclk,ereset, ~cclk_v[`W-1], ~n_740_v[`W-1], notalu2_v);
  spice_latch latch_4952(eclk,ereset, ~cclk_v[`W-1], ~n_795_v[`W-1], n_360_v);
  spice_latch latch_4977(eclk,ereset, ~cclk_v[`W-1], ~n_490_v[`W-1], notidl4_v);
  spice_latch latch_4976(eclk,ereset, ~cclk_v[`W-1], ~n_182_v[`W-1], n_265_v);
  spice_latch latch_4975(eclk,ereset, ~cp1_v[`W-1], ~notRdy0_v[`W-1], n_902_v);
  spice_latch latch_4974(eclk,ereset, ~cp1_v[`W-1], ~n_789_v[`W-1], notdor7_v);
  spice_latch latch_4971(eclk,ereset, ~cclk_v[`W-1], ~n_862_v[`W-1], pipeUNK11_v);
  spice_latch latch_4970(eclk,ereset, ~cp1_v[`W-1], ~n_299_v[`W-1], n_1625_v);
  spice_latch latch_5022(eclk,ereset, ~cclk_v[`W-1], ~n_318_v[`W-1], pipeUNK14_v);
  spice_latch latch_5023(eclk,ereset, ~cclk_v[`W-1], ~n_188_v[`W-1], pipeT4out_v);
  spice_latch latch_5020(eclk,ereset, ~cclk_v[`W-1], ~n_462_v[`W-1], n_878_v);
  spice_latch latch_5021(eclk,ereset, ~cp1_v[`W-1], ~n_845_v[`W-1], p2_v);
  spice_latch latch_5026(eclk,ereset, ~cclk_v[`W-1], ~n_1090_v[`W-1], n_1683_v);
  spice_latch latch_5027(eclk,ereset, ~cclk_v[`W-1], ~n_586_v[`W-1], pipeBRtaken_v);
  spice_latch latch_5024(eclk,ereset, ~cp1_v[`W-1], ~n_1087_v[`W-1], n_1132_v);
  spice_latch latch_5025(eclk,ereset, ~cclk_v[`W-1], ~C78_v[`W-1], C78_phi2_v);
  spice_latch latch_5028(eclk,ereset, ~cclk_v[`W-1], ~n_983_v[`W-1], nots0_v);
  spice_latch latch_5029(eclk,ereset, ~cclk_v[`W-1], ~n_272_v[`W-1], n_1162_v);
  spice_latch latch_5123(eclk,ereset, ~cclk_v[`W-1], ~n_1175_v[`W-1], pipeUNK28_v);
  spice_latch latch_5122(eclk,ereset, ~cclk_v[`W-1], ~n_1085_v[`W-1], pipeUNK23_v);
  spice_latch latch_5129(eclk,ereset, ~cclk_v[`W-1], ~op_EORS_v[`W-1], n_982_v);
  spice_latch latch_5128(eclk,ereset, ~cclk_v[`W-1], ~n_484_v[`W-1], pclp7_v);
  spice_latch latch_5004(eclk,ereset, ~cp1_v[`W-1], ~n_1375_v[`W-1], n_95_v);
  spice_latch latch_5005(eclk,ereset, ~cp1_v[`W-1], ~n_1089_v[`W-1], n_1529_v);
  spice_latch latch_5006(eclk,ereset, ~cclk_v[`W-1], ~n_1631_v[`W-1], pclp3_v);
  spice_latch latch_5007(eclk,ereset, ~cp1_v[`W-1], ~brk_done_v[`W-1], n_1291_v);
  spice_latch latch_5000(eclk,ereset, ~cp1_v[`W-1], ~n_913_v[`W-1], n_1274_v);
  spice_latch latch_5001(eclk,ereset, ~cclk_v[`W-1], ~n_1688_v[`W-1], n_680_v);
  spice_latch latch_5002(eclk,ereset, ~cclk_v[`W-1], ~VEC0_v[`W-1], n_1126_v);
  spice_latch latch_5003(eclk,ereset, ~cclk_v[`W-1], ~_WR_v[`W-1], pipe_WR_phi2_v);
  spice_latch latch_5008(eclk,ereset, ~cp1_v[`W-1], ~n_428_v[`W-1], n_644_v);
  spice_latch latch_5009(eclk,ereset, ~cp1_v[`W-1], ~n_1474_v[`W-1], notdor1_v);
  spice_latch latch_5068(eclk,ereset, ~cclk_v[`W-1], ~n_1705_v[`W-1], n_1020_v);
  spice_latch latch_5069(eclk,ereset, ~cclk_v[`W-1], ~n_944_v[`W-1], pipeUNK37_v);
  spice_latch latch_5066(eclk,ereset, ~cp1_v[`W-1], ~INTG_v[`W-1], n_50_v);
  spice_latch latch_5067(eclk,ereset, ~cclk_v[`W-1], ~n_396_v[`W-1], n_796_v);
  spice_latch latch_5064(eclk,ereset, ~cclk_v[`W-1], ~op_ORS_v[`W-1], n_88_v);
  spice_latch latch_5065(eclk,ereset, ~cclk_v[`W-1], ~n_629_v[`W-1], n_760_v);
  spice_latch latch_5062(eclk,ereset, ~cclk_v[`W-1], ~n_515_v[`W-1], n_1411_v);
  spice_latch latch_5063(eclk,ereset, ~cclk_v[`W-1], ~n_1211_v[`W-1], n_897_v);
  spice_latch latch_5060(eclk,ereset, ~cclk_v[`W-1], ~n_504_v[`W-1], pipeUNK41_v);
  spice_latch latch_5061(eclk,ereset, ~cclk_v[`W-1], ~op_ANDS_v[`W-1], n_1574_v);
  spice_latch latch_5071(eclk,ereset, ~cclk_v[`W-1], ~n_17_v[`W-1], pipe_T0_v);
  spice_latch latch_5040(eclk,ereset, ~cp1_v[`W-1], ~n_1290_v[`W-1], n_698_v);
  spice_latch latch_5041(eclk,ereset, ~cclk_v[`W-1], ~n_374_v[`W-1], pd6_v);
  spice_latch latch_5042(eclk,ereset, ~cp1_v[`W-1], ~n_1718_v[`W-1], n_671_v);
  spice_latch latch_5043(eclk,ereset, ~cp1_v[`W-1], ~notRdy0_v[`W-1], n_1679_v);
  spice_latch latch_5044(eclk,ereset, ~cp1_v[`W-1], ~n_1215_v[`W-1], n_223_v);
  spice_latch latch_5046(eclk,ereset, ~cp1_v[`W-1], ~n_931_v[`W-1], n_1674_v);
  spice_latch latch_5048(eclk,ereset, ~cclk_v[`W-1], ~n_604_v[`W-1], n_1477_v);
  spice_latch latch_5049(eclk,ereset, ~cclk_v[`W-1], ~n_501_v[`W-1], pipeUNK35_v);
  spice_latch latch_5118(eclk,ereset, ~cclk_v[`W-1], ~n_80_v[`W-1], n_1333_v);
  spice_latch latch_4973(eclk,ereset, ~cclk_v[`W-1], ~n_213_v[`W-1], notidl1_v);
  spice_latch latch_4979(eclk,ereset, ~cclk_v[`W-1], ~n_513_v[`W-1], pipeUNK06_v);
  spice_latch latch_4978(eclk,ereset, ~cclk_v[`W-1], ~op_T__bit_v[`W-1], n_1673_v);
  spice_latch latch_5141(eclk,ereset, ~cclk_v[`W-1], ~n_844_v[`W-1], n_459_v);
  spice_latch latch_5140(eclk,ereset, ~cclk_v[`W-1], ~n_1486_v[`W-1], n_126_v);
  spice_latch latch_5143(eclk,ereset, ~cclk_v[`W-1], ~n_1575_v[`W-1], pipeT2out_v);
  spice_latch latch_5142(eclk,ereset, ~cclk_v[`W-1], ~n_474_v[`W-1], n_15_v);
  spice_latch latch_5145(eclk,ereset, ~cp1_v[`W-1], ~n_1339_v[`W-1], n_597_v);
  spice_latch latch_5144(eclk,ereset, ~cclk_v[`W-1], ~n_973_v[`W-1], nots4_v);
  spice_latch latch_5146(eclk,ereset, ~cp1_v[`W-1], ~notRnWprepad_v[`W-1], n_402_v);
  spice_latch latch_5157(eclk,ereset, ~cp1_v[`W-1], ~n_1650_v[`W-1], n_94_v);
  spice_latch latch_4988(eclk,ereset, ~cclk_v[`W-1], ~n_1192_v[`W-1], pchp6_v);
  spice_latch latch_4989(eclk,ereset, ~cclk_v[`W-1], ~n_632_v[`W-1], n_339_v);
  spice_latch latch_4980(eclk,ereset, ~cp1_v[`W-1], ~n_854_v[`W-1], n_1395_v);
  spice_latch latch_4981(eclk,ereset, ~cp1_v[`W-1], ~n_468_v[`W-1], n_18_v);
  spice_latch latch_4984(eclk,ereset, ~cclk_v[`W-1], ~nnT2BR_v[`W-1], n_1269_v);
  spice_latch latch_4985(eclk,ereset, ~cclk_v[`W-1], ~n_327_v[`W-1], pipeUNK09_v);
  spice_latch latch_5169(eclk,ereset, ~cclk_v[`W-1], ~n_588_v[`W-1], notidl7_v);
  spice_latch latch_5168(eclk,ereset, ~cp1_v[`W-1], ~n_1180_v[`W-1], n_1533_v);
  spice_latch latch_5163(eclk,ereset, ~cclk_v[`W-1], ~n_958_v[`W-1], n_865_v);
  spice_latch latch_5162(eclk,ereset, ~cclk_v[`W-1], ~n_889_v[`W-1], pipeUNK42_v);
  spice_latch latch_5161(eclk,ereset, ~cclk_v[`W-1], ~n_90_v[`W-1], pipeUNK05_v);
  spice_latch latch_5160(eclk,ereset, ~cp1_v[`W-1], ~n_472_v[`W-1], n_1606_v);
  spice_latch latch_5167(eclk,ereset, ~cclk_v[`W-1], ~n_1455_v[`W-1], n_1505_v);
  spice_latch latch_5166(eclk,ereset, ~cclk_v[`W-1], ~n_1037_v[`W-1], n_266_v);
  spice_latch latch_5165(eclk,ereset, ~cclk_v[`W-1], ~n_1649_v[`W-1], n_1027_v);
  spice_latch latch_5164(eclk,ereset, ~cclk_v[`W-1], ~Reset0_v[`W-1], pipephi2Reset0_v);
  spice_latch latch_5108(eclk,ereset, ~cclk_v[`W-1], ~n_306_v[`W-1], n_581_v);
  spice_latch latch_5105(eclk,ereset, ~cclk_v[`W-1], ~_op_set_C_v[`W-1], pipeUNK08_v);
  spice_latch latch_5104(eclk,ereset, ~cclk_v[`W-1], ~n_678_v[`W-1], pipeT3out_v);
  spice_latch latch_5101(eclk,ereset, ~cclk_v[`W-1], ~n_1225_v[`W-1], n_1121_v);
  spice_latch latch_5100(eclk,ereset, ~cclk_v[`W-1], ~n_1402_v[`W-1], pchp2_v);
  spice_latch latch_5103(eclk,ereset, ~cclk_v[`W-1], ~n_1024_v[`W-1], n_1699_v);
  spice_latch latch_5102(eclk,ereset, ~cclk_v[`W-1], ~n_277_v[`W-1], notalu5_v);
  spice_latch latch_5152(eclk,ereset, ~cclk_v[`W-1], ~x_op_T__adc_sbc_v[`W-1], pipeUNK03_v);
  spice_latch latch_5153(eclk,ereset, ~cclk_v[`W-1], ~DC78_v[`W-1], DC78_phi2_v);
  spice_latch latch_5150(eclk,ereset, ~cclk_v[`W-1], ~n_14_v[`W-1], pipeUNK20_v);
  spice_latch latch_5151(eclk,ereset, ~cclk_v[`W-1], ~n_696_v[`W-1], n_610_v);
  spice_latch latch_5156(eclk,ereset, ~cclk_v[`W-1], ~n_506_v[`W-1], n_1602_v);
  spice_latch latch_5154(eclk,ereset, ~cclk_v[`W-1], ~n_207_v[`W-1], n_1061_v);
  spice_latch latch_5155(eclk,ereset, ~cclk_v[`W-1], ~n_31_v[`W-1], pipeUNK16_v);
  spice_latch latch_5127(eclk,ereset, ~cclk_v[`W-1], ~n_1319_v[`W-1], pd1_v);
  spice_latch latch_5126(eclk,ereset, ~cclk_v[`W-1], ~n_93_v[`W-1], pd0_v);
  spice_latch latch_5125(eclk,ereset, ~cclk_v[`W-1], ~op_SRS_v[`W-1], pipeUNK27_v);
  spice_latch latch_5124(eclk,ereset, ~cclk_v[`W-1], ~n_160_v[`W-1], n_1049_v);
  spice_latch latch_5121(eclk,ereset, ~cclk_v[`W-1], ~n_378_v[`W-1], pipeT5out_v);
  spice_latch latch_5120(eclk,ereset, ~cp1_v[`W-1], ~n_1215_v[`W-1], n_1528_v);
  spice_latch latch_5149(eclk,ereset, ~cclk_v[`W-1], ~n_29_v[`W-1], pipeUNK22_v);
  spice_latch latch_5148(eclk,ereset, ~cclk_v[`W-1], ~n_1717_v[`W-1], n_1113_v);
  spice_latch latch_5093(eclk,ereset, ~cclk_v[`W-1], ~n_1069_v[`W-1], n_1177_v);
  spice_latch latch_5092(eclk,ereset, ~cclk_v[`W-1], ~n_1045_v[`W-1], pipeUNK13_v);
  spice_latch latch_5091(eclk,ereset, ~cclk_v[`W-1], ~n_728_v[`W-1], pipeVectorA0_v);
  spice_latch latch_5090(eclk,ereset, ~cp1_v[`W-1], ~n_109_v[`W-1], n_1161_v);
  spice_latch latch_5097(eclk,ereset, ~cclk_v[`W-1], ~n_1711_v[`W-1], nots1_v);
  spice_latch latch_5096(eclk,ereset, ~cclk_v[`W-1], ~n_1586_v[`W-1], n_621_v);
  spice_latch latch_5095(eclk,ereset, ~cclk_v[`W-1], ~n_1225_v[`W-1], pipedpc28_v);
  spice_latch latch_5094(eclk,ereset, ~cclk_v[`W-1], ~Reset0_v[`W-1], pipephi2Reset0x_v);
  spice_latch latch_5099(eclk,ereset, ~cclk_v[`W-1], ~n_1073_v[`W-1], pclp5_v);
  spice_latch latch_5098(eclk,ereset, ~cclk_v[`W-1], ~n_1358_v[`W-1], n_521_v);
  spice_latch latch_4948(eclk,ereset, ~cp1_v[`W-1], ~n_645_v[`W-1], n_562_v);
  spice_latch latch_4949(eclk,ereset, ~cp1_v[`W-1], ~n_262_v[`W-1], n_1447_v);
  spice_latch latch_4947(eclk,ereset, ~cclk_v[`W-1], ~n_11_v[`W-1], n_55_v);
  spice_latch latch_4960(eclk,ereset, ~cclk_v[`W-1], ~n_385_v[`W-1], pipeUNK30_v);
  spice_latch latch_4961(eclk,ereset, ~cclk_v[`W-1], ~n_442_v[`W-1], n_509_v);
  spice_latch latch_4962(eclk,ereset, ~cp1_v[`W-1], ~n_1368_v[`W-1], n_1149_v);
  spice_latch latch_4963(eclk,ereset, ~cclk_v[`W-1], ~n_1179_v[`W-1], n_393_v);
  spice_latch latch_4964(eclk,ereset, ~cp1_v[`W-1], ~n_430_v[`W-1], n_1570_v);
  spice_latch latch_4965(eclk,ereset, ~cclk_v[`W-1], ~_VEC_v[`W-1], pipe_VEC_v);
  spice_latch latch_4966(eclk,ereset, ~cclk_v[`W-1], ~n_261_v[`W-1], pipeUNK36_v);
  spice_latch latch_4967(eclk,ereset, ~cp1_v[`W-1], ~n_959_v[`W-1], n_323_v);
  spice_latch latch_4968(eclk,ereset, ~cclk_v[`W-1], ~n_169_v[`W-1], pipeUNK29_v);
  spice_latch latch_4969(eclk,ereset, ~cp1_v[`W-1], ~n_1687_v[`W-1], notdor0_v);
  spice_latch latch_5031(eclk,ereset, ~cclk_v[`W-1], ~n_191_v[`W-1], pipeUNK40_v);
  spice_latch latch_5030(eclk,ereset, ~cp1_v[`W-1], ~n_1495_v[`W-1], p3_v);
  spice_latch latch_5033(eclk,ereset, ~cclk_v[`W-1], ~n_264_v[`W-1], n_799_v);
  spice_latch latch_5032(eclk,ereset, ~cclk_v[`W-1], ~n_1500_v[`W-1], n_526_v);
  spice_latch latch_5035(eclk,ereset, ~cclk_v[`W-1], ~n_334_v[`W-1], pipeUNK17_v);
  spice_latch latch_5034(eclk,ereset, ~cclk_v[`W-1], ~n_264_v[`W-1], n_1693_v);
  spice_latch latch_5037(eclk,ereset, ~cclk_v[`W-1], ~n_1065_v[`W-1], n_1124_v);
  spice_latch latch_5036(eclk,ereset, ~cclk_v[`W-1], ~n_824_v[`W-1], n_398_v);
  spice_latch latch_5039(eclk,ereset, ~cclk_v[`W-1], ~n_62_v[`W-1], pd7_v);
  spice_latch latch_5038(eclk,ereset, ~cclk_v[`W-1], ~n_111_v[`W-1], pd2_v);
  spice_latch latch_5019(eclk,ereset, ~cclk_v[`W-1], ~notaluvout_v[`W-1], n_408_v);
  spice_latch latch_5018(eclk,ereset, ~cclk_v[`W-1], ~n_779_v[`W-1], n_805_v);
  spice_latch latch_5013(eclk,ereset, ~cclk_v[`W-1], ~n_1594_v[`W-1], n_688_v);
  spice_latch latch_5012(eclk,ereset, ~cclk_v[`W-1], ~n_1374_v[`W-1], n_1252_v);
  spice_latch latch_5011(eclk,ereset, ~cclk_v[`W-1], ~n_1347_v[`W-1], n_1527_v);
  spice_latch latch_5010(eclk,ereset, ~cp1_v[`W-1], ~n_1380_v[`W-1], n_666_v);
  spice_latch latch_5017(eclk,ereset, ~cp1_v[`W-1], ~n_1141_v[`W-1], n_101_v);
  spice_latch latch_5016(eclk,ereset, ~cclk_v[`W-1], ~n_132_v[`W-1], pipeUNK26_v);
  spice_latch latch_5015(eclk,ereset, ~cclk_v[`W-1], ~n_1209_v[`W-1], n_663_v);
  spice_latch latch_5014(eclk,ereset, ~cp1_v[`W-1], ~n_1181_v[`W-1], n_69_v);
  spice_latch latch_4982(eclk,ereset, ~cp1_v[`W-1], ~n_1039_v[`W-1], n_24_v);
  spice_latch latch_4983(eclk,ereset, ~cclk_v[`W-1], ~n_20_v[`W-1], n_993_v);
  spice_latch latch_4987(eclk,ereset, ~cp1_v[`W-1], ~n_1178_v[`W-1], n_590_v);
  spice_latch latch_5079(eclk,ereset, ~cclk_v[`W-1], ~n_1071_v[`W-1], notalu3_v);
  spice_latch latch_5078(eclk,ereset, ~cclk_v[`W-1], ~n_473_v[`W-1], pipeUNK33_v);
  spice_latch latch_5075(eclk,ereset, ~cclk_v[`W-1], ~n_1199_v[`W-1], notidl2_v);
  spice_latch latch_5074(eclk,ereset, ~cclk_v[`W-1], ~n_1081_v[`W-1], pipeUNK32_v);
  spice_latch latch_5077(eclk,ereset, ~cclk_v[`W-1], ~n_389_v[`W-1], pipeUNK31_v);
  spice_latch latch_5076(eclk,ereset, ~cclk_v[`W-1], ~n_824_v[`W-1], pipeUNK34_v);
  spice_latch latch_5070(eclk,ereset, ~cp1_v[`W-1], ~n_1684_v[`W-1], notdor6_v);
  spice_latch latch_5073(eclk,ereset, ~cclk_v[`W-1], ~notaluoutmux1_v[`W-1], notalu1_v);
  spice_latch latch_5072(eclk,ereset, ~cp1_v[`W-1], ~_TWOCYCLE_v[`W-1], _TWOCYCLE_phi1_v);
  spice_latch latch_5057(eclk,ereset, ~cp1_v[`W-1], ~n_797_v[`W-1], notdor4_v);
  spice_latch latch_5056(eclk,ereset, ~cclk_v[`W-1], ~n_1117_v[`W-1], pipeVectorA1_v);
  spice_latch latch_5055(eclk,ereset, ~cp1_v[`W-1], ~n_916_v[`W-1], n_1409_v);
  spice_latch latch_5053(eclk,ereset, ~cp1_v[`W-1], ~n_1376_v[`W-1], notdor2_v);
  spice_latch latch_5052(eclk,ereset, ~cclk_v[`W-1], ~n_952_v[`W-1], n_1509_v);
  spice_latch latch_5051(eclk,ereset, ~cp1_v[`W-1], ~n_961_v[`W-1], notdor5_v);
  spice_latch latch_5050(eclk,ereset, ~cp1_v[`W-1], ~notRdy0_v[`W-1], n_1276_v);
  spice_latch latch_5059(eclk,ereset, ~cp1_v[`W-1], ~n_1091_v[`W-1], n_1360_v);
  spice_latch latch_5058(eclk,ereset, ~cclk_v[`W-1], ~n_700_v[`W-1], n_1565_v);
  spice_latch latch_5158(eclk,ereset, ~cp1_v[`W-1], ~notRdy0_v[`W-1], n_1272_v);
  spice_latch latch_5159(eclk,ereset, ~cp1_v[`W-1], ~n_1093_v[`W-1], n_226_v);
  spice_latch latch_5147(eclk,ereset, ~cclk_v[`W-1], ~n_568_v[`W-1], notidl5_v);
  spice_latch latch_5119(eclk,ereset, ~cclk_v[`W-1], ~n_1657_v[`W-1], pchp4_v);
  spice_latch latch_5112(eclk,ereset, ~cp1_v[`W-1], ~n_626_v[`W-1], n_756_v);
  spice_latch latch_5113(eclk,ereset, ~cclk_v[`W-1], ~n_104_v[`W-1], n_1221_v);
  spice_latch latch_5170(eclk,ereset, ~cp1_v[`W-1], ~notRdy0_v[`W-1], n_1624_v);
  spice_latch latch_5171(eclk,ereset, ~cp1_v[`W-1], ~n_330_v[`W-1], n_675_v);
  spice_latch latch_5172(eclk,ereset, ~cclk_v[`W-1], ~n_1712_v[`W-1], pipeVectorA2_v);
  spice_latch latch_5173(eclk,ereset, ~cclk_v[`W-1], ~n_496_v[`W-1], nots5_v);
  spice_latch latch_4999(eclk,ereset, ~cclk_v[`W-1], ~n_875_v[`W-1], n_469_v);
  spice_latch latch_4998(eclk,ereset, ~cclk_v[`W-1], ~n_176_v[`W-1], n_598_v);
  spice_latch latch_4991(eclk,ereset, ~cclk_v[`W-1], ~n_1379_v[`W-1], pipeUNK07_v);
  spice_latch latch_4990(eclk,ereset, ~cclk_v[`W-1], ~n_1190_v[`W-1], nots2_v);
  spice_latch latch_4993(eclk,ereset, ~cclk_v[`W-1], ~n_1130_v[`W-1], n_512_v);
  spice_latch latch_4992(eclk,ereset, ~cclk_v[`W-1], ~n_1099_v[`W-1], pclp1_v);
  spice_latch latch_4995(eclk,ereset, ~cclk_v[`W-1], ~n_774_v[`W-1], pipeUNK02_v);
  spice_latch latch_4994(eclk,ereset, ~cclk_v[`W-1], ~n_674_v[`W-1], n_745_v);
  spice_latch latch_4997(eclk,ereset, ~cclk_v[`W-1], ~op_SUMS_v[`W-1], n_415_v);
  spice_latch latch_4996(eclk,ereset, ~cclk_v[`W-1], ~op_SRS_v[`W-1], n_968_v);
  spice_latch latch_5116(eclk,ereset, ~cclk_v[`W-1], ~n_19_v[`W-1], pipeUNK18_v);
  spice_latch latch_5117(eclk,ereset, ~cclk_v[`W-1], ~n_304_v[`W-1], notalu7_v);
  spice_latch latch_5114(eclk,ereset, ~cp1_v[`W-1], ~n_420_v[`W-1], n_47_v);
  spice_latch latch_5115(eclk,ereset, ~cclk_v[`W-1], ~n_1231_v[`W-1], pipeUNK21_v);
  spice_latch latch_5110(eclk,ereset, ~cclk_v[`W-1], ~n_608_v[`W-1], n_559_v);
  spice_latch latch_5111(eclk,ereset, ~cp1_v[`W-1], ~n_457_v[`W-1], notdor3_v);

  spice_node_2 n_dor5(eclk, ereset, dor5_port_3,dor5_port_4, dor5_v);
  spice_node_2 n_dor4(eclk, ereset, dor4_port_3,dor4_port_4, dor4_v);
  spice_node_2 n_dor7(eclk, ereset, dor7_port_0,dor7_port_4, dor7_v);
  spice_node_2 n_dor6(eclk, ereset, dor6_port_2,dor6_port_4, dor6_v);
  spice_node_2 n_dor1(eclk, ereset, dor1_port_0,dor1_port_4, dor1_v);
  spice_node_2 n_dor0(eclk, ereset, dor0_port_0,dor0_port_4, dor0_v);
  spice_node_2 n_dor3(eclk, ereset, dor3_port_3,dor3_port_4, dor3_v);
  spice_node_2 n_dor2(eclk, ereset, dor2_port_3,dor2_port_4, dor2_v);
  spice_node_2 n__DBZ(eclk, ereset, _DBZ_port_2,_DBZ_port_0, _DBZ_v);
  spice_node_2 n__DBE(eclk, ereset, _DBE_port_3,_DBE_port_5, _DBE_v);
  spice_node_2 n_n_1714(eclk, ereset, n_1714_port_2,n_1714_port_1, n_1714_v);
  spice_node_2 n_n_1715(eclk, ereset, n_1715_port_2,n_1715_port_3, n_1715_v);
  spice_node_2 n_n_1716(eclk, ereset, n_1716_port_6,n_1716_port_5, n_1716_v);
  spice_node_2 n_n_1717(eclk, ereset, n_1717_port_8,n_1717_port_12, n_1717_v);
  spice_node_2 n_n_1247(eclk, ereset, n_1247_port_13,n_1247_port_0, n_1247_v);
  spice_node_2 n_n_1244(eclk, ereset, n_1244_port_2,n_1244_port_1, n_1244_v);
  spice_node_2 n_n_1245(eclk, ereset, n_1245_port_2,n_1245_port_1, n_1245_v);
  spice_node_2 n_n_1718(eclk, ereset, n_1718_port_2,n_1718_port_1, n_1718_v);
  spice_node_2 n_n_1719(eclk, ereset, n_1719_port_2,n_1719_port_0, n_1719_v);
  spice_node_2 n__ABL7(eclk, ereset, _ABL7_port_3,_ABL7_port_1, _ABL7_v);
  spice_node_2 n__ABL6(eclk, ereset, _ABL6_port_3,_ABL6_port_1, _ABL6_v);
  spice_node_2 n__ABL5(eclk, ereset, _ABL5_port_3,_ABL5_port_0, _ABL5_v);
  spice_node_2 n__ABL3(eclk, ereset, _ABL3_port_3,_ABL3_port_0, _ABL3_v);
  spice_node_2 n__ABL2(eclk, ereset, _ABL2_port_2,_ABL2_port_3, _ABL2_v);
  spice_node_2 n__ABL1(eclk, ereset, _ABL1_port_2,_ABL1_port_3, _ABL1_v);
  spice_node_2 n__ABL0(eclk, ereset, _ABL0_port_2,_ABL0_port_3, _ABL0_v);
  spice_node_2 n_dpc5_SADL(eclk, ereset, dpc5_SADL_port_0,dpc5_SADL_port_7, dpc5_SADL_v);
  spice_node_2 n_n_604(eclk, ereset, n_604_port_10,n_604_port_15, n_604_v);
  spice_node_2 n_n_600(eclk, ereset, n_600_port_1,n_600_port_4, n_600_v);
  spice_node_2 n_n_602(eclk, ereset, n_602_port_2,n_602_port_0, n_602_v);
  spice_node_2 n_n_603(eclk, ereset, n_603_port_2,n_603_port_1, n_603_v);
  spice_node_2 n_n_608(eclk, ereset, n_608_port_2,n_608_port_0, n_608_v);
  spice_node_2 n_n_609(eclk, ereset, n_609_port_6,n_609_port_4, n_609_v);
  spice_node_2 n_pd6_clearIR(eclk, ereset, pd6_clearIR_port_3,pd6_clearIR_port_4, pd6_clearIR_v);
  spice_node_2 n_n_462(eclk, ereset, n_462_port_2,n_462_port_3, n_462_v);
  spice_node_3 n_n_465(eclk, ereset, n_465_port_2,n_465_port_0,n_465_port_1, n_465_v);
  spice_node_2 n_n_466(eclk, ereset, n_466_port_6,n_466_port_4, n_466_v);
  spice_node_2 n_n_467(eclk, ereset, n_467_port_6,n_467_port_4, n_467_v);
  spice_node_2 n_n_468(eclk, ereset, n_468_port_3,n_468_port_6, n_468_v);
  spice_node_2 n_op_T4_brk(eclk, ereset, op_T4_brk_port_10,op_T4_brk_port_12, op_T4_brk_v);
  spice_node_2 n_rw(eclk, ereset, rw_port_0,rw_port_1, rw_v);
  spice_node_2 n_x_op_T3_plp_pla(eclk, ereset, x_op_T3_plp_pla_port_8,x_op_T3_plp_pla_port_10, x_op_T3_plp_pla_v);
  spice_node_3 n_idl7(eclk, ereset, idl7_port_2,idl7_port_0,idl7_port_1, idl7_v);
  spice_node_3 n_idl6(eclk, ereset, idl6_port_2,idl6_port_0,idl6_port_1, idl6_v);
  spice_node_3 n_idl5(eclk, ereset, idl5_port_2,idl5_port_0,idl5_port_1, idl5_v);
  spice_node_3 n_idl4(eclk, ereset, idl4_port_2,idl4_port_0,idl4_port_1, idl4_v);
  spice_node_3 n_idl3(eclk, ereset, idl3_port_2,idl3_port_0,idl3_port_1, idl3_v);
  spice_node_3 n_idl2(eclk, ereset, idl2_port_2,idl2_port_0,idl2_port_1, idl2_v);
  spice_node_3 n_idl1(eclk, ereset, idl1_port_2,idl1_port_0,idl1_port_1, idl1_v);
  spice_node_3 n_idl0(eclk, ereset, idl0_port_2,idl0_port_0,idl0_port_1, idl0_v);
  spice_node_2 n_n_1523(eclk, ereset, n_1523_port_2,n_1523_port_3, n_1523_v);
  spice_node_2 n_n_1521(eclk, ereset, n_1521_port_2,n_1521_port_1, n_1521_v);
  spice_node_2 n_n_1526(eclk, ereset, n_1526_port_2,n_1526_port_1, n_1526_v);
  spice_node_4 n_n_733(eclk, ereset, n_733_port_2,n_733_port_3,n_733_port_0,n_733_port_1, n_733_v);
  spice_node_2 n_dpc20_ADDSB06(eclk, ereset, dpc20_ADDSB06_port_0,dpc20_ADDSB06_port_5, dpc20_ADDSB06_v);
  spice_node_5 n_n_1389(eclk, ereset, n_1389_port_2,n_1389_port_3,n_1389_port_0,n_1389_port_1,n_1389_port_4, n_1389_v);
  spice_node_4 n_n_1387(eclk, ereset, n_1387_port_2,n_1387_port_3,n_1387_port_0,n_1387_port_1, n_1387_v);
  spice_node_2 n_n_1386(eclk, ereset, n_1386_port_2,n_1386_port_3, n_1386_v);
  spice_node_3 n_n_1383(eclk, ereset, n_1383_port_2,n_1383_port_0,n_1383_port_1, n_1383_v);
  spice_node_2 n_n_1380(eclk, ereset, n_1380_port_4,n_1380_port_5, n_1380_v);
  spice_node_2 n_n_917(eclk, ereset, n_917_port_3,n_917_port_5, n_917_v);
  spice_node_2 n_x6(eclk, ereset, x6_port_0,x6_port_1, x6_v);
  spice_node_2 n_n_819(eclk, ereset, n_819_port_6,n_819_port_4, n_819_v);
  spice_node_2 n_n_818(eclk, ereset, n_818_port_4,n_818_port_5, n_818_v);
  spice_node_2 n_n_811(eclk, ereset, n_811_port_7,n_811_port_5, n_811_v);
  spice_node_2 n_n_810(eclk, ereset, n_810_port_3,n_810_port_4, n_810_v);
  spice_node_2 n_n_813(eclk, ereset, n_813_port_3,n_813_port_4, n_813_v);
  spice_node_2 n_n_812(eclk, ereset, n_812_port_3,n_812_port_4, n_812_v);
  spice_node_2 n_n_815(eclk, ereset, n_815_port_2,n_815_port_0, n_815_v);
  spice_node_1 n_irq(eclk, ereset, irq_port_2, irq_v);
  spice_node_2 n_ir0(eclk, ereset, ir0_port_3,ir0_port_4, ir0_v);
  spice_node_2 n_ir1(eclk, ereset, ir1_port_2,ir1_port_3, ir1_v);
  spice_node_2 n_ir2(eclk, ereset, ir2_port_72,ir2_port_0, ir2_v);
  spice_node_2 n_ir3(eclk, ereset, ir3_port_1,ir3_port_41, ir3_v);
  spice_node_2 n_ir4(eclk, ereset, ir4_port_70,ir4_port_68, ir4_v);
  spice_node_2 n_ir5(eclk, ereset, ir5_port_0,ir5_port_33, ir5_v);
  spice_node_2 n_ir6(eclk, ereset, ir6_port_42,ir6_port_43, ir6_v);
  spice_node_2 n_ir7(eclk, ereset, ir7_port_59,ir7_port_60, ir7_v);
  spice_node_3 n_n_1267(eclk, ereset, n_1267_port_2,n_1267_port_3,n_1267_port_0, n_1267_v);
  spice_node_2 n_n_1260(eclk, ereset, n_1260_port_2,n_1260_port_3, n_1260_v);
  spice_node_2 n_op_T__inx(eclk, ereset, op_T__inx_port_9,op_T__inx_port_11, op_T__inx_v);
  spice_node_2 n_n_5(eclk, ereset, n_5_port_2,n_5_port_0, n_5_v);
  spice_node_2 n_n_6(eclk, ereset, n_6_port_4,n_6_port_5, n_6_v);
  spice_node_2 n_n_7(eclk, ereset, n_7_port_2,n_7_port_4, n_7_v);
  spice_node_5 n_n_3(eclk, ereset, n_3_port_2,n_3_port_3,n_3_port_0,n_3_port_1,n_3_port_4, n_3_v);
  spice_node_3 n_aluanandb0(eclk, ereset, aluanandb0_port_9,aluanandb0_port_3,aluanandb0_port_5, aluanandb0_v);
  spice_node_4 n_aluanandb1(eclk, ereset, aluanandb1_port_0,aluanandb1_port_1,aluanandb1_port_4,aluanandb1_port_5, aluanandb1_v);
  spice_node_2 n_n_1240(eclk, ereset, n_1240_port_2,n_1240_port_1, n_1240_v);
  spice_node_2 n_n_1711(eclk, ereset, n_1711_port_2,n_1711_port_1, n_1711_v);
  spice_node_2 n_n_1712(eclk, ereset, n_1712_port_4,n_1712_port_5, n_1712_v);
  spice_node_2 n_op_T0_php_pha(eclk, ereset, op_T0_php_pha_port_8,op_T0_php_pha_port_10, op_T0_php_pha_v);
  spice_node_3 n_dasb6(eclk, ereset, dasb6_port_3,dasb6_port_0,dasb6_port_5, dasb6_v);
  spice_node_3 n_dasb5(eclk, ereset, dasb5_port_3,dasb5_port_1,dasb5_port_5, dasb5_v);
  spice_node_3 n_dasb3(eclk, ereset, dasb3_port_3,dasb3_port_1,dasb3_port_5, dasb3_v);
  spice_node_3 n_dasb2(eclk, ereset, dasb2_port_3,dasb2_port_1,dasb2_port_5, dasb2_v);
  spice_node_3 n_dasb1(eclk, ereset, dasb1_port_3,dasb1_port_0,dasb1_port_5, dasb1_v);
  spice_node_2 n_n_662(eclk, ereset, n_662_port_2,n_662_port_0, n_662_v);
  spice_node_2 n_n_664(eclk, ereset, n_664_port_2,n_664_port_1, n_664_v);
  spice_node_4 n_alu4(eclk, ereset, alu4_port_2,alu4_port_3,alu4_port_0,alu4_port_1, alu4_v);
  spice_node_4 n_alu5(eclk, ereset, alu5_port_3,alu5_port_0,alu5_port_1,alu5_port_4, alu5_v);
  spice_node_4 n_alu6(eclk, ereset, alu6_port_2,alu6_port_0,alu6_port_1,alu6_port_4, alu6_v);
  spice_node_4 n_alu7(eclk, ereset, alu7_port_2,alu7_port_3,alu7_port_0,alu7_port_1, alu7_v);
  spice_node_4 n_alu0(eclk, ereset, alu0_port_2,alu0_port_3,alu0_port_0,alu0_port_1, alu0_v);
  spice_node_4 n_alu1(eclk, ereset, alu1_port_3,alu1_port_0,alu1_port_1,alu1_port_4, alu1_v);
  spice_node_4 n_alu2(eclk, ereset, alu2_port_3,alu2_port_0,alu2_port_1,alu2_port_4, alu2_v);
  spice_node_4 n_alu3(eclk, ereset, alu3_port_2,alu3_port_3,alu3_port_0,alu3_port_1, alu3_v);
  spice_node_2 n__ABL4(eclk, ereset, _ABL4_port_3,_ABL4_port_1, _ABL4_v);
  spice_node_5 n_n_488(eclk, ereset, n_488_port_2,n_488_port_3,n_488_port_0,n_488_port_1,n_488_port_4, n_488_v);
  spice_node_2 n_n_484(eclk, ereset, n_484_port_2,n_484_port_3, n_484_v);
  spice_node_2 n_n_485(eclk, ereset, n_485_port_2,n_485_port_1, n_485_v);
  spice_node_2 n_n_480(eclk, ereset, n_480_port_2,n_480_port_4, n_480_v);
  spice_node_5 n_n_481(eclk, ereset, n_481_port_2,n_481_port_3,n_481_port_0,n_481_port_1,n_481_port_4, n_481_v);
  spice_node_2 n_PD_xxx010x1(eclk, ereset, PD_xxx010x1_port_6,PD_xxx010x1_port_5, PD_xxx010x1_v);
  spice_node_2 n_op_shift(eclk, ereset, op_shift_port_4,op_shift_port_5, op_shift_v);
  spice_node_2 n_op_xy(eclk, ereset, op_xy_port_6,op_xy_port_5, op_xy_v);
  spice_node_2 n_op_T0_cld_sed(eclk, ereset, op_T0_cld_sed_port_8,op_T0_cld_sed_port_9, op_T0_cld_sed_v);
  spice_node_2 n_n_327(eclk, ereset, n_327_port_3,n_327_port_4, n_327_v);
  spice_node_5 n_n_326(eclk, ereset, n_326_port_2,n_326_port_3,n_326_port_0,n_326_port_1,n_326_port_4, n_326_v);
  spice_node_2 n__AxB_0__C0in(eclk, ereset, _AxB_0__C0in_port_3,_AxB_0__C0in_port_4, _AxB_0__C0in_v);
  spice_node_2 n_n_321(eclk, ereset, n_321_port_2,n_321_port_3, n_321_v);
  spice_node_2 n_n_320(eclk, ereset, n_320_port_3,n_320_port_0, n_320_v);
  spice_node_2 n_n_1105(eclk, ereset, n_1105_port_2,n_1105_port_0, n_1105_v);
  spice_node_2 n_n_1107(eclk, ereset, n_1107_port_7,n_1107_port_10, n_1107_v);
  spice_node_2 n_n_1106(eclk, ereset, n_1106_port_8,n_1106_port_12, n_1106_v);
  spice_node_2 n_n_1101(eclk, ereset, n_1101_port_2,n_1101_port_3, n_1101_v);
  spice_node_3 n_n_1100(eclk, ereset, n_1100_port_2,n_1100_port_3,n_1100_port_0, n_1100_v);
  spice_node_2 n_n_1109(eclk, ereset, n_1109_port_9,n_1109_port_5, n_1109_v);
  spice_node_2 n_pd4_clearIR(eclk, ereset, pd4_clearIR_port_8,pd4_clearIR_port_6, pd4_clearIR_v);
  spice_node_2 n_op_ror(eclk, ereset, op_ror_port_6,op_ror_port_5, op_ror_v);
  spice_node_2 n_dpc6_SBS(eclk, ereset, dpc6_SBS_port_11,dpc6_SBS_port_12, dpc6_SBS_v);
  spice_node_2 n_n_345(eclk, ereset, n_345_port_4,n_345_port_10, n_345_v);
  spice_node_2 n_n_347(eclk, ereset, n_347_port_8,n_347_port_9, n_347_v);
  spice_node_2 n_n_340(eclk, ereset, n_340_port_2,n_340_port_0, n_340_v);
  spice_node_5 n_n_831(eclk, ereset, n_831_port_2,n_831_port_3,n_831_port_0,n_831_port_1,n_831_port_4, n_831_v);
  spice_node_2 n_n_830(eclk, ereset, n_830_port_4,n_830_port_5, n_830_v);
  spice_node_2 n_n_839(eclk, ereset, n_839_port_2,n_839_port_1, n_839_v);
  spice_node_2 n_n_838(eclk, ereset, n_838_port_2,n_838_port_0, n_838_v);
  spice_node_2 n_op_T0_ldy_mem(eclk, ereset, op_T0_ldy_mem_port_8,op_T0_ldy_mem_port_7, op_T0_ldy_mem_v);
  spice_node_2 n_D1x1(eclk, ereset, D1x1_port_6,D1x1_port_5, D1x1_v);
  spice_node_2 n_s3(eclk, ereset, s3_port_0,s3_port_1, s3_v);
  spice_node_2 n_s2(eclk, ereset, s2_port_0,s2_port_1, s2_v);
  spice_node_2 n_s1(eclk, ereset, s1_port_0,s1_port_1, s1_v);
  spice_node_2 n_s0(eclk, ereset, s0_port_0,s0_port_1, s0_v);
  spice_node_2 n_s7(eclk, ereset, s7_port_2,s7_port_0, s7_v);
  spice_node_2 n_s6(eclk, ereset, s6_port_0,s6_port_1, s6_v);
  spice_node_2 n_s5(eclk, ereset, s5_port_0,s5_port_1, s5_v);
  spice_node_2 n_s4(eclk, ereset, s4_port_0,s4_port_1, s4_v);
  spice_node_2 n_so(eclk, ereset, so_port_2,so_port_3, so_v);
  spice_node_2 n_dpc15_ANDS(eclk, ereset, dpc15_ANDS_port_9,dpc15_ANDS_port_0, dpc15_ANDS_v);
  spice_node_2 n_n_1585(eclk, ereset, n_1585_port_2,n_1585_port_1, n_1585_v);
  spice_node_2 n_n_1586(eclk, ereset, n_1586_port_2,n_1586_port_1, n_1586_v);
  spice_node_2 n__TWOCYCLE(eclk, ereset, _TWOCYCLE_port_7,_TWOCYCLE_port_4, _TWOCYCLE_v);
  spice_node_2 n_dpc27_SBADH(eclk, ereset, dpc27_SBADH_port_9,dpc27_SBADH_port_0, dpc27_SBADH_v);
  spice_node_2 n_pd3_clearIR(eclk, ereset, pd3_clearIR_port_6,pd3_clearIR_port_4, pd3_clearIR_v);
  spice_node_3 n_n_649(eclk, ereset, n_649_port_0,n_649_port_7,n_649_port_5, n_649_v);
  spice_node_3 n_n_138(eclk, ereset, n_138_port_2,n_138_port_0,n_138_port_1, n_138_v);
  spice_node_2 n_n_139(eclk, ereset, n_139_port_2,n_139_port_1, n_139_v);
  spice_node_2 n_n_641(eclk, ereset, n_641_port_3,n_641_port_0, n_641_v);
  spice_node_3 n_n_642(eclk, ereset, n_642_port_3,n_642_port_0,n_642_port_1, n_642_v);
  spice_node_2 n_n_643(eclk, ereset, n_643_port_3,n_643_port_4, n_643_v);
  spice_node_2 n_n_132(eclk, ereset, n_132_port_2,n_132_port_1, n_132_v);
  spice_node_2 n_n_645(eclk, ereset, n_645_port_2,n_645_port_3, n_645_v);
  spice_node_2 n_n_646(eclk, ereset, n_646_port_8,n_646_port_2, n_646_v);
  spice_node_2 n_n_647(eclk, ereset, n_647_port_3,n_647_port_5, n_647_v);
  spice_node_3 n_n_1632(eclk, ereset, n_1632_port_7,n_1632_port_4,n_1632_port_5, n_1632_v);
  spice_node_2 n_n_1635(eclk, ereset, n_1635_port_2,n_1635_port_1, n_1635_v);
  spice_node_2 n__AxB_6__C56(eclk, ereset, _AxB_6__C56_port_3,_AxB_6__C56_port_4, _AxB_6__C56_v);
  spice_node_2 n_pd0_clearIR(eclk, ereset, pd0_clearIR_port_8,pd0_clearIR_port_5, pd0_clearIR_v);
  spice_node_2 n_op_T0_shift_a(eclk, ereset, op_T0_shift_a_port_8,op_T0_shift_a_port_11, op_T0_shift_a_v);
  spice_node_2 n___AxB7__C67(eclk, ereset, __AxB7__C67_port_3,__AxB7__C67_port_4, __AxB7__C67_v);
  spice_node_2 n_n_1439(eclk, ereset, n_1439_port_2,n_1439_port_1, n_1439_v);
  spice_node_2 n__VEC(eclk, ereset, _VEC_port_8,_VEC_port_5, _VEC_v);
  spice_node_2 n_n_1129(eclk, ereset, n_1129_port_4,n_1129_port_5, n_1129_v);
  spice_node_2 n_n_1120(eclk, ereset, n_1120_port_2,n_1120_port_1, n_1120_v);
  spice_node_2 n_n_587(eclk, ereset, n_587_port_2,n_587_port_1, n_587_v);
  spice_node_2 n_n_586(eclk, ereset, n_586_port_3,n_586_port_5, n_586_v);
  spice_node_3 n_n_583(eclk, ereset, n_583_port_2,n_583_port_0,n_583_port_1, n_583_v);
  spice_node_2 n_n_582(eclk, ereset, n_582_port_2,n_582_port_3, n_582_v);
  spice_node_2 n_n_588(eclk, ereset, n_588_port_2,n_588_port_0, n_588_v);
  spice_node_2 n_op_rmw(eclk, ereset, op_rmw_port_2,op_rmw_port_0, op_rmw_v);
  spice_node_2 n_n_366(eclk, ereset, n_366_port_3,n_366_port_5, n_366_v);
  spice_node_2 n_n_368(eclk, ereset, n_368_port_8,n_368_port_7, n_368_v);
  spice_node_2 n_op_jmp(eclk, ereset, op_jmp_port_8,op_jmp_port_7, op_jmp_v);
  spice_node_2 n_C12(eclk, ereset, C12_port_2,C12_port_3, C12_v);
  spice_node_2 n_n_1433(eclk, ereset, n_1433_port_6,n_1433_port_4, n_1433_v);
  spice_node_2 n_op_shift_right(eclk, ereset, op_shift_right_port_4,op_shift_right_port_5, op_shift_right_v);
  spice_node_2 n_op_EORS(eclk, ereset, op_EORS_port_2,op_EORS_port_3, op_EORS_v);
  spice_node_2 n_x_op_T__adc_sbc(eclk, ereset, x_op_T__adc_sbc_port_8,x_op_T__adc_sbc_port_6, x_op_T__adc_sbc_v);
  spice_node_2 n_n_1631(eclk, ereset, n_1631_port_2,n_1631_port_3, n_1631_v);
  spice_node_3 n_notir0(eclk, ereset, notir0_port_0,notir0_port_1,notir0_port_28, notir0_v);
  spice_node_3 n_notir1(eclk, ereset, notir1_port_21,notir1_port_23,notir1_port_22, notir1_v);
  spice_node_3 n_notir2(eclk, ereset, notir2_port_19,notir2_port_0,notir2_port_20, notir2_v);
  spice_node_3 n_notir3(eclk, ereset, notir3_port_51,notir3_port_0,notir3_port_1, notir3_v);
  spice_node_3 n_notir4(eclk, ereset, notir4_port_25,notir4_port_24,notir4_port_26, notir4_v);
  spice_node_3 n_notir5(eclk, ereset, notir5_port_36,notir5_port_37,notir5_port_0, notir5_v);
  spice_node_3 n_notir6(eclk, ereset, notir6_port_0,notir6_port_1,notir6_port_39, notir6_v);
  spice_node_3 n_notir7(eclk, ereset, notir7_port_34,notir7_port_35,notir7_port_33, notir7_v);
  spice_node_2 n_n_93(eclk, ereset, n_93_port_2,n_93_port_0, n_93_v);
  spice_node_2 n_n_90(eclk, ereset, n_90_port_3,n_90_port_4, n_90_v);
  spice_node_2 n_n_91(eclk, ereset, n_91_port_3,n_91_port_0, n_91_v);
  spice_node_2 n_op_lsr_ror_dec_inc(eclk, ereset, op_lsr_ror_dec_inc_port_3,op_lsr_ror_dec_inc_port_4, op_lsr_ror_dec_inc_v);
  spice_node_2 n_n_110(eclk, ereset, n_110_port_2,n_110_port_1, n_110_v);
  spice_node_2 n_n_111(eclk, ereset, n_111_port_2,n_111_port_1, n_111_v);
  spice_node_2 n_n_118(eclk, ereset, n_118_port_2,n_118_port_1, n_118_v);
  spice_node_2 n_n_119(eclk, ereset, n_119_port_3,n_119_port_0, n_119_v);
  spice_node_2 n_cp1(eclk, ereset, cp1_port_75,cp1_port_50, cp1_v);
  spice_node_2 n_a3(eclk, ereset, a3_port_0,a3_port_1, a3_v);
  spice_node_2 n_a6(eclk, ereset, a6_port_2,a6_port_0, a6_v);
  spice_node_2 n_n_696(eclk, ereset, n_696_port_3,n_696_port_5, n_696_v);
  spice_node_2 n_n_1199(eclk, ereset, n_1199_port_2,n_1199_port_0, n_1199_v);
  spice_node_2 n_n_930(eclk, ereset, n_930_port_3,n_930_port_4, n_930_v);
  spice_node_2 n_DA_AxB2(eclk, ereset, DA_AxB2_port_3,DA_AxB2_port_5, DA_AxB2_v);
  spice_node_2 n_n_1479(eclk, ereset, n_1479_port_0,n_1479_port_1, n_1479_v);
  spice_node_2 n_sync(eclk, ereset, sync_port_0,sync_port_1, sync_v);
  spice_node_2 n_n_1499(eclk, ereset, n_1499_port_3,n_1499_port_0, n_1499_v);
  spice_node_2 n_n_1325(eclk, ereset, n_1325_port_2,n_1325_port_4, n_1325_v);
  spice_node_5 n_n_1496(eclk, ereset, n_1496_port_2,n_1496_port_3,n_1496_port_0,n_1496_port_1,n_1496_port_4, n_1496_v);
  spice_node_2 n_n_1495(eclk, ereset, n_1495_port_8,n_1495_port_4, n_1495_v);
  spice_node_2 n_n_1492(eclk, ereset, n_1492_port_3,n_1492_port_0, n_1492_v);
  spice_node_2 n_n_1323(eclk, ereset, n_1323_port_2,n_1323_port_0, n_1323_v);
  spice_node_2 n_n_1141(eclk, ereset, n_1141_port_2,n_1141_port_1, n_1141_v);
  spice_node_2 n_n_568(eclk, ereset, n_568_port_2,n_568_port_1, n_568_v);
  spice_node_2 n_n_565(eclk, ereset, n_565_port_2,n_565_port_0, n_565_v);
  spice_node_4 n_n_564(eclk, ereset, n_564_port_2,n_564_port_3,n_564_port_0,n_564_port_1, n_564_v);
  spice_node_2 n_n_567(eclk, ereset, n_567_port_0,n_567_port_4, n_567_v);
  spice_node_2 n_n_566(eclk, ereset, n_566_port_8,n_566_port_4, n_566_v);
  spice_node_3 n___AxBxC_6(eclk, ereset, __AxBxC_6_port_3,__AxBxC_6_port_1,__AxBxC_6_port_5, __AxBxC_6_v);
  spice_node_3 n___AxBxC_7(eclk, ereset, __AxBxC_7_port_3,__AxBxC_7_port_0,__AxBxC_7_port_5, __AxBxC_7_v);
  spice_node_3 n___AxBxC_4(eclk, ereset, __AxBxC_4_port_2,__AxBxC_4_port_3,__AxBxC_4_port_5, __AxBxC_4_v);
  spice_node_3 n___AxBxC_5(eclk, ereset, __AxBxC_5_port_3,__AxBxC_5_port_1,__AxBxC_5_port_5, __AxBxC_5_v);
  spice_node_3 n___AxBxC_2(eclk, ereset, __AxBxC_2_port_3,__AxBxC_2_port_1,__AxBxC_2_port_5, __AxBxC_2_v);
  spice_node_3 n___AxBxC_3(eclk, ereset, __AxBxC_3_port_3,__AxBxC_3_port_1,__AxBxC_3_port_5, __AxBxC_3_v);
  spice_node_3 n___AxBxC_0(eclk, ereset, __AxBxC_0_port_2,__AxBxC_0_port_3,__AxBxC_0_port_5, __AxBxC_0_v);
  spice_node_3 n___AxBxC_1(eclk, ereset, __AxBxC_1_port_3,__AxBxC_1_port_1,__AxBxC_1_port_5, __AxBxC_1_v);
  spice_node_2 n_n_300(eclk, ereset, n_300_port_8,n_300_port_7, n_300_v);
  spice_node_5 n_n_304(eclk, ereset, n_304_port_2,n_304_port_3,n_304_port_0,n_304_port_1,n_304_port_4, n_304_v);
  spice_node_2 n_n_307(eclk, ereset, n_307_port_6,n_307_port_4, n_307_v);
  spice_node_2 n_n_306(eclk, ereset, n_306_port_2,n_306_port_0, n_306_v);
  spice_node_2 n_aluaorb0(eclk, ereset, aluaorb0_port_2,aluaorb0_port_1, aluaorb0_v);
  spice_node_2 n_x_op_T0_tya(eclk, ereset, x_op_T0_tya_port_9,x_op_T0_tya_port_10, x_op_T0_tya_v);
  spice_node_2 n_x_op_T4_ind_y(eclk, ereset, x_op_T4_ind_y_port_7,x_op_T4_ind_y_port_10, x_op_T4_ind_y_v);
  spice_node_2 n_pclp0(eclk, ereset, pclp0_port_2,pclp0_port_1, pclp0_v);
  spice_node_2 n_pclp2(eclk, ereset, pclp2_port_2,pclp2_port_1, pclp2_v);
  spice_node_2 n_pclp4(eclk, ereset, pclp4_port_2,pclp4_port_0, pclp4_v);
  spice_node_2 n_pclp6(eclk, ereset, pclp6_port_2,pclp6_port_0, pclp6_v);
  spice_node_2 n_op_T3_branch(eclk, ereset, op_T3_branch_port_8,op_T3_branch_port_7, op_T3_branch_v);
  spice_node_2 n_ab12(eclk, ereset, ab12_port_0,ab12_port_1, ab12_v);
  spice_node_2 n_ab13(eclk, ereset, ab13_port_0,ab13_port_1, ab13_v);
  spice_node_2 n_ab10(eclk, ereset, ab10_port_0,ab10_port_1, ab10_v);
  spice_node_2 n_ab11(eclk, ereset, ab11_port_0,ab11_port_1, ab11_v);
  spice_node_2 n_n_79(eclk, ereset, n_79_port_2,n_79_port_1, n_79_v);
  spice_node_2 n_ab14(eclk, ereset, ab14_port_0,ab14_port_1, ab14_v);
  spice_node_2 n_ab15(eclk, ereset, ab15_port_0,ab15_port_1, ab15_v);
  spice_node_2 n_n_75(eclk, ereset, n_75_port_2,n_75_port_0, n_75_v);
  spice_node_2 n_n_70(eclk, ereset, n_70_port_3,n_70_port_4, n_70_v);
  spice_node_2 n_n_71(eclk, ereset, n_71_port_2,n_71_port_0, n_71_v);
  spice_node_5 n_n_72(eclk, ereset, n_72_port_2,n_72_port_3,n_72_port_0,n_72_port_1,n_72_port_4, n_72_v);
  spice_node_2 n_n_1705(eclk, ereset, n_1705_port_3,n_1705_port_4, n_1705_v);
  spice_node_2 n_n_1256(eclk, ereset, n_1256_port_2,n_1256_port_0, n_1256_v);
  spice_node_2 n_op_T0_tya(eclk, ereset, op_T0_tya_port_9,op_T0_tya_port_11, op_T0_tya_v);
  spice_node_2 n_n_172(eclk, ereset, n_172_port_2,n_172_port_3, n_172_v);
  spice_node_2 n_n_176(eclk, ereset, n_176_port_3,n_176_port_4, n_176_v);
  spice_node_3 n_n_177(eclk, ereset, n_177_port_2,n_177_port_0,n_177_port_1, n_177_v);
  spice_node_2 n_n_797(eclk, ereset, n_797_port_2,n_797_port_1, n_797_v);
  spice_node_2 n_n_794(eclk, ereset, n_794_port_1,n_794_port_4, n_794_v);
  spice_node_2 n_n_795(eclk, ereset, n_795_port_2,n_795_port_0, n_795_v);
  spice_node_2 n_n_790(eclk, ereset, n_790_port_7,n_790_port_5, n_790_v);
  spice_node_2 n_n_798(eclk, ereset, n_798_port_1,n_798_port_4, n_798_v);
  spice_node_2 n_n_1305(eclk, ereset, n_1305_port_2,n_1305_port_1, n_1305_v);
  spice_node_2 n_n_1304(eclk, ereset, n_1304_port_3,n_1304_port_4, n_1304_v);
  spice_node_2 n_n_1303(eclk, ereset, n_1303_port_3,n_1303_port_7, n_1303_v);
  spice_node_5 n_n_1301(eclk, ereset, n_1301_port_2,n_1301_port_3,n_1301_port_0,n_1301_port_1,n_1301_port_4, n_1301_v);
  spice_node_2 n_n_1300(eclk, ereset, n_1300_port_2,n_1300_port_3, n_1300_v);
  spice_node_3 n_n_1309(eclk, ereset, n_1309_port_2,n_1309_port_3,n_1309_port_1, n_1309_v);
  spice_node_2 n_n_330(eclk, ereset, n_330_port_7,n_330_port_4, n_330_v);
  spice_node_5 n_n_332(eclk, ereset, n_332_port_2,n_332_port_3,n_332_port_0,n_332_port_1,n_332_port_4, n_332_v);
  spice_node_2 n_n_1166(eclk, ereset, n_1166_port_2,n_1166_port_3, n_1166_v);
  spice_node_4 n_n_1169(eclk, ereset, n_1169_port_2,n_1169_port_3,n_1169_port_0,n_1169_port_1, n_1169_v);
  spice_node_2 n_PD_1xx000x0(eclk, ereset, PD_1xx000x0_port_6,PD_1xx000x0_port_7, PD_1xx000x0_v);
  spice_node_2 n_n_548(eclk, ereset, n_548_port_2,n_548_port_0, n_548_v);
  spice_node_2 n_op_T2_brk(eclk, ereset, op_T2_brk_port_9,op_T2_brk_port_10, op_T2_brk_v);
  spice_node_2 n_n_543(eclk, ereset, n_543_port_3,n_543_port_0, n_543_v);
  spice_node_2 n_n_541(eclk, ereset, n_541_port_3,n_541_port_1, n_541_v);
  spice_node_2 n_n_544(eclk, ereset, n_544_port_2,n_544_port_1, n_544_v);
  spice_node_2 n_C56(eclk, ereset, C56_port_3,C56_port_0, C56_v);
  spice_node_2 n_n_890(eclk, ereset, n_890_port_2,n_890_port_1, n_890_v);
  spice_node_2 n_n_322(eclk, ereset, n_322_port_2,n_322_port_1, n_322_v);
  spice_node_2 n_n_896(eclk, ereset, n_896_port_2,n_896_port_1, n_896_v);
  spice_node_2 n_n_329(eclk, ereset, n_329_port_3,n_329_port_0, n_329_v);
  spice_node_2 n_xx_op_T5_jsr(eclk, ereset, xx_op_T5_jsr_port_9,xx_op_T5_jsr_port_11, xx_op_T5_jsr_v);
  spice_node_2 n_PD_xxxx10x0(eclk, ereset, PD_xxxx10x0_port_6,PD_xxxx10x0_port_5, PD_xxxx10x0_v);
  spice_node_2 n_n_1028(eclk, ereset, n_1028_port_2,n_1028_port_0, n_1028_v);
  spice_node_2 n_dpc24_ACSB(eclk, ereset, dpc24_ACSB_port_1,dpc24_ACSB_port_12, dpc24_ACSB_v);
  spice_node_2 n_n_152(eclk, ereset, n_152_port_6,n_152_port_5, n_152_v);
  spice_node_2 n_n_154(eclk, ereset, n_154_port_2,n_154_port_3, n_154_v);
  spice_node_2 n_rdy(eclk, ereset, rdy_port_2,rdy_port_3, rdy_v);
  spice_node_2 n_n_1347(eclk, ereset, n_1347_port_8,n_1347_port_7, n_1347_v);
  spice_node_2 n_op_ORS(eclk, ereset, op_ORS_port_2,op_ORS_port_3, op_ORS_v);
  spice_node_2 n_n_1346(eclk, ereset, n_1346_port_3,n_1346_port_0, n_1346_v);
  spice_node_2 n__AxB_2__C12(eclk, ereset, _AxB_2__C12_port_3,_AxB_2__C12_port_4, _AxB_2__C12_v);
  spice_node_2 n_n_1364(eclk, ereset, n_1364_port_3,n_1364_port_0, n_1364_v);
  spice_node_2 n_n_1369(eclk, ereset, n_1369_port_2,n_1369_port_3, n_1369_v);
  spice_node_2 n_n_1368(eclk, ereset, n_1368_port_4,n_1368_port_5, n_1368_v);
  spice_node_2 n_clearIR(eclk, ereset, clearIR_port_9,clearIR_port_18, clearIR_v);
  spice_node_2 n_op_T__cpx_cpy_imm_zp(eclk, ereset, op_T__cpx_cpy_imm_zp_port_8,op_T__cpx_cpy_imm_zp_port_7, op_T__cpx_cpy_imm_zp_v);
  spice_node_2 n_n_1187(eclk, ereset, n_1187_port_2,n_1187_port_0, n_1187_v);
  spice_node_2 n_n_1181(eclk, ereset, n_1181_port_3,n_1181_port_6, n_1181_v);
  spice_node_2 n_n_1180(eclk, ereset, n_1180_port_3,n_1180_port_4, n_1180_v);
  spice_node_2 n_op_T5_mem_ind_idx(eclk, ereset, op_T5_mem_ind_idx_port_7,op_T5_mem_ind_idx_port_5, op_T5_mem_ind_idx_v);
  spice_node_2 n_n_520(eclk, ereset, n_520_port_0,n_520_port_4, n_520_v);
  spice_node_2 n_n_523(eclk, ereset, n_523_port_6,n_523_port_4, n_523_v);
  spice_node_2 n_n_525(eclk, ereset, n_525_port_4,n_525_port_5, n_525_v);
  spice_node_2 n_C78(eclk, ereset, C78_port_2,C78_port_1, C78_v);
  spice_node_2 n_dpc21_ADDADL(eclk, ereset, dpc21_ADDADL_port_9,dpc21_ADDADL_port_0, dpc21_ADDADL_v);
  spice_node_5 n_n_1592(eclk, ereset, n_1592_port_2,n_1592_port_3,n_1592_port_0,n_1592_port_1,n_1592_port_4, n_1592_v);
  spice_node_2 n_n_31(eclk, ereset, n_31_port_0,n_31_port_6, n_31_v);
  spice_node_2 n_n_34(eclk, ereset, n_34_port_2,n_34_port_1, n_34_v);
  spice_node_2 n_n_35(eclk, ereset, n_35_port_4,n_35_port_5, n_35_v);
  spice_node_2 n_n_36(eclk, ereset, n_36_port_6,n_36_port_4, n_36_v);
  spice_node_2 n_n_37(eclk, ereset, n_37_port_3,n_37_port_4, n_37_v);
  spice_node_3 n_db1(eclk, ereset, db1_port_1,db1_port_4,db1_port_5, db1_v);
  spice_node_3 n_db0(eclk, ereset, db0_port_1,db0_port_4,db0_port_5, db0_v);
  spice_node_3 n_db3(eclk, ereset, db3_port_2,db3_port_3,db3_port_5, db3_v);
  spice_node_3 n_db2(eclk, ereset, db2_port_2,db2_port_3,db2_port_5, db2_v);
  spice_node_3 n_db5(eclk, ereset, db5_port_0,db5_port_4,db5_port_5, db5_v);
  spice_node_3 n_db4(eclk, ereset, db4_port_3,db4_port_0,db4_port_5, db4_v);
  spice_node_3 n_db7(eclk, ereset, db7_port_3,db7_port_1,db7_port_5, db7_v);
  spice_node_3 n_db6(eclk, ereset, db6_port_0,db6_port_4,db6_port_5, db6_v);
  spice_node_2 n_pchp5(eclk, ereset, pchp5_port_2,pchp5_port_1, pchp5_v);
  spice_node_2 n_pchp7(eclk, ereset, pchp7_port_2,pchp7_port_0, pchp7_v);
  spice_node_2 n_pchp1(eclk, ereset, pchp1_port_2,pchp1_port_0, pchp1_v);
  spice_node_2 n_pchp3(eclk, ereset, pchp3_port_2,pchp3_port_0, pchp3_v);
  spice_node_2 n_clk1out(eclk, ereset, clk1out_port_0,clk1out_port_1, clk1out_v);
  spice_node_2 n__WR(eclk, ereset, _WR_port_8,_WR_port_7, _WR_v);
  spice_node_5 n_n_1647(eclk, ereset, n_1647_port_2,n_1647_port_3,n_1647_port_0,n_1647_port_1,n_1647_port_4, n_1647_v);
  spice_node_2 n_n_1642(eclk, ereset, n_1642_port_2,n_1642_port_4, n_1642_v);
  spice_node_2 n_n_1643(eclk, ereset, n_1643_port_3,n_1643_port_4, n_1643_v);
  spice_node_2 n_n_1640(eclk, ereset, n_1640_port_2,n_1640_port_0, n_1640_v);
  spice_node_3 n_n_1641(eclk, ereset, n_1641_port_2,n_1641_port_3,n_1641_port_1, n_1641_v);
  spice_node_2 n_n_1649(eclk, ereset, n_1649_port_11,n_1649_port_12, n_1649_v);
  spice_node_2 n__op_branch_bit6(eclk, ereset, _op_branch_bit6_port_0,_op_branch_bit6_port_4, _op_branch_bit6_v);
  spice_node_2 n__op_branch_bit7(eclk, ereset, _op_branch_bit7_port_1,_op_branch_bit7_port_4, _op_branch_bit7_v);
  spice_node_2 n_n_1184(eclk, ereset, n_1184_port_8,n_1184_port_4, n_1184_v);
  spice_node_2 n_op_rol_ror(eclk, ereset, op_rol_ror_port_7,op_rol_ror_port_5, op_rol_ror_v);
  spice_node_4 n_n_1491(eclk, ereset, n_1491_port_2,n_1491_port_3,n_1491_port_0,n_1491_port_1, n_1491_v);
  spice_node_2 n_n_201(eclk, ereset, n_201_port_3,n_201_port_1, n_201_v);
  spice_node_3 n_n_206(eclk, ereset, n_206_port_3,n_206_port_0,n_206_port_5, n_206_v);
  spice_node_2 n_clock1(eclk, ereset, clock1_port_68,clock1_port_40, clock1_v);
  spice_node_2 n_clock2(eclk, ereset, clock2_port_12,clock2_port_13, clock2_v);
  spice_node_2 n_n_1434(eclk, ereset, n_1434_port_2,n_1434_port_0, n_1434_v);
  spice_node_5 n_n_1344(eclk, ereset, n_1344_port_2,n_1344_port_3,n_1344_port_0,n_1344_port_1,n_1344_port_4, n_1344_v);
  spice_node_2 n_op_asl_rol(eclk, ereset, op_asl_rol_port_7,op_asl_rol_port_5, op_asl_rol_v);
  spice_node_2 n_short_circuit_idx_add(eclk, ereset, short_circuit_idx_add_port_7,short_circuit_idx_add_port_5, short_circuit_idx_add_v);
  spice_node_2 n_n_507(eclk, ereset, n_507_port_2,n_507_port_3, n_507_v);
  spice_node_2 n_n_506(eclk, ereset, n_506_port_4,n_506_port_5, n_506_v);
  spice_node_2 n_n_504(eclk, ereset, n_504_port_2,n_504_port_3, n_504_v);
  spice_node_2 n_n_503(eclk, ereset, n_503_port_2,n_503_port_0, n_503_v);
  spice_node_2 n_n_501(eclk, ereset, n_501_port_4,n_501_port_5, n_501_v);
  spice_node_2 n_x_op_T0_bit(eclk, ereset, x_op_T0_bit_port_8,x_op_T0_bit_port_9, x_op_T0_bit_v);
  spice_node_2 n_n_16(eclk, ereset, n_16_port_0,n_16_port_5, n_16_v);
  spice_node_2 n_n_17(eclk, ereset, n_17_port_6,n_17_port_5, n_17_v);
  spice_node_2 n_n_14(eclk, ereset, n_14_port_4,n_14_port_5, n_14_v);
  spice_node_2 n_n_10(eclk, ereset, n_10_port_6,n_10_port_4, n_10_v);
  spice_node_2 n_n_11(eclk, ereset, n_11_port_9,n_11_port_6, n_11_v);
  spice_node_3 n_n_1084(eclk, ereset, n_1084_port_0,n_1084_port_6,n_1084_port_5, n_1084_v);
  spice_node_2 n_n_1085(eclk, ereset, n_1085_port_3,n_1085_port_6, n_1085_v);
  spice_node_2 n_n_1087(eclk, ereset, n_1087_port_3,n_1087_port_4, n_1087_v);
  spice_node_2 n_n_1081(eclk, ereset, n_1081_port_2,n_1081_port_3, n_1081_v);
  spice_node_2 n_n_1082(eclk, ereset, n_1082_port_5,n_1082_port_10, n_1082_v);
  spice_node_3 n_n_1083(eclk, ereset, n_1083_port_1,n_1083_port_7,n_1083_port_4, n_1083_v);
  spice_node_2 n_n_1089(eclk, ereset, n_1089_port_2,n_1089_port_1, n_1089_v);
  spice_node_2 n_dpc35_PCHC(eclk, ereset, dpc35_PCHC_port_8,dpc35_PCHC_port_7, dpc35_PCHC_v);
  spice_node_2 n_n_1265(eclk, ereset, n_1265_port_2,n_1265_port_3, n_1265_v);
  spice_node_4 n_n_1661(eclk, ereset, n_1661_port_2,n_1661_port_3,n_1661_port_0,n_1661_port_1, n_1661_v);
  spice_node_2 n_n_1662(eclk, ereset, n_1662_port_3,n_1662_port_1, n_1662_v);
  spice_node_2 n_n_1262(eclk, ereset, n_1262_port_2,n_1262_port_3, n_1262_v);
  spice_node_3 n_n_1668(eclk, ereset, n_1668_port_2,n_1668_port_3,n_1668_port_0, n_1668_v);
  spice_node_2 n_op_T2_abs_y(eclk, ereset, op_T2_abs_y_port_6,op_T2_abs_y_port_7, op_T2_abs_y_v);
  spice_node_2 n_n_267(eclk, ereset, n_267_port_4,n_267_port_5, n_267_v);
  spice_node_2 n_n_264(eclk, ereset, n_264_port_8,n_264_port_6, n_264_v);
  spice_node_2 n_n_262(eclk, ereset, n_262_port_3,n_262_port_6, n_262_v);
  spice_node_2 n_n_260(eclk, ereset, n_260_port_3,n_260_port_4, n_260_v);
  spice_node_2 n_n_261(eclk, ereset, n_261_port_3,n_261_port_4, n_261_v);
  spice_node_2 n_n_269(eclk, ereset, n_269_port_3,n_269_port_4, n_269_v);
  spice_node_2 n_dpc32_PCHADH(eclk, ereset, dpc32_PCHADH_port_0,dpc32_PCHADH_port_1, dpc32_PCHADH_v);
  spice_node_8 n_idb1(eclk, ereset, idb1_port_8,idb1_port_9,idb1_port_3,idb1_port_0,idb1_port_7,idb1_port_4,idb1_port_5,idb1_port_10, idb1_v);
  spice_node_8 n_idb0(eclk, ereset, idb0_port_8,idb0_port_2,idb0_port_1,idb0_port_6,idb0_port_7,idb0_port_4,idb0_port_5,idb0_port_10, idb0_v);
  spice_node_8 n_idb3(eclk, ereset, idb3_port_8,idb3_port_9,idb3_port_3,idb3_port_0,idb3_port_1,idb3_port_6,idb3_port_5,idb3_port_10, idb3_v);
  spice_node_8 n_idb2(eclk, ereset, idb2_port_9,idb2_port_3,idb2_port_0,idb2_port_1,idb2_port_6,idb2_port_4,idb2_port_5,idb2_port_10, idb2_v);
  spice_node_7 n_idb5(eclk, ereset, idb5_port_8,idb5_port_9,idb5_port_2,idb5_port_6,idb5_port_7,idb5_port_4,idb5_port_5, idb5_v);
  spice_node_8 n_idb4(eclk, ereset, idb4_port_8,idb4_port_9,idb4_port_0,idb4_port_6,idb4_port_7,idb4_port_4,idb4_port_5,idb4_port_10, idb4_v);
  spice_node_8 n_idb7(eclk, ereset, idb7_port_8,idb7_port_9,idb7_port_2,idb7_port_3,idb7_port_0,idb7_port_7,idb7_port_4,idb7_port_10, idb7_v);
  spice_node_8 n_idb6(eclk, ereset, idb6_port_9,idb6_port_3,idb6_port_0,idb6_port_6,idb6_port_7,idb6_port_5,idb6_port_10,idb6_port_11, idb6_v);
  spice_node_2 n_n_8(eclk, ereset, n_8_port_1,n_8_port_4, n_8_v);
  spice_node_2 n_op_T3_mem_abs(eclk, ereset, op_T3_mem_abs_port_7,op_T3_mem_abs_port_5, op_T3_mem_abs_v);
  spice_node_2 n_op_T2_ADL_ADD(eclk, ereset, op_T2_ADL_ADD_port_3,op_T2_ADL_ADD_port_4, op_T2_ADL_ADD_v);
  spice_node_2 n_n_1417(eclk, ereset, n_1417_port_2,n_1417_port_0, n_1417_v);
  spice_node_2 n_n_1416(eclk, ereset, n_1416_port_2,n_1416_port_0, n_1416_v);
  spice_node_2 n_n_1413(eclk, ereset, n_1413_port_2,n_1413_port_1, n_1413_v);
  spice_node_2 n_n_1412(eclk, ereset, n_1412_port_2,n_1412_port_0, n_1412_v);
  spice_node_3 n_n_381(eclk, ereset, n_381_port_2,n_381_port_3,n_381_port_1, n_381_v);
  spice_node_2 n_n_383(eclk, ereset, n_383_port_3,n_383_port_0, n_383_v);
  spice_node_2 n_n_385(eclk, ereset, n_385_port_3,n_385_port_4, n_385_v);
  spice_node_2 n_n_384(eclk, ereset, n_384_port_8,n_384_port_6, n_384_v);
  spice_node_2 n_n_386(eclk, ereset, n_386_port_3,n_386_port_0, n_386_v);
  spice_node_2 n_n_389(eclk, ereset, n_389_port_1,n_389_port_4, n_389_v);
  spice_node_2 n_n_388(eclk, ereset, n_388_port_6,n_388_port_5, n_388_v);
  spice_node_2 n_op_T__shift_a(eclk, ereset, op_T__shift_a_port_9,op_T__shift_a_port_7, op_T__shift_a_v);
  spice_node_2 n_n_927(eclk, ereset, n_927_port_3,n_927_port_1, n_927_v);
  spice_node_2 n_n_920(eclk, ereset, n_920_port_2,n_920_port_1, n_920_v);
  spice_node_2 n_n_923(eclk, ereset, n_923_port_0,n_923_port_4, n_923_v);
  spice_node_3 n_n_928(eclk, ereset, n_928_port_2,n_928_port_3,n_928_port_1, n_928_v);
  spice_node_2 n_n_1039(eclk, ereset, n_1039_port_3,n_1039_port_5, n_1039_v);
  spice_node_3 n_alub2(eclk, ereset, alub2_port_0,alub2_port_1,alub2_port_4, alub2_v);
  spice_node_2 n_pch7(eclk, ereset, pch7_port_2,pch7_port_1, pch7_v);
  spice_node_2 n_pch6(eclk, ereset, pch6_port_2,pch6_port_0, pch6_v);
  spice_node_2 n_pch5(eclk, ereset, pch5_port_2,pch5_port_0, pch5_v);
  spice_node_2 n_pch4(eclk, ereset, pch4_port_2,pch4_port_1, pch4_v);
  spice_node_2 n_pch3(eclk, ereset, pch3_port_2,pch3_port_1, pch3_v);
  spice_node_2 n_pch2(eclk, ereset, pch2_port_0,pch2_port_1, pch2_v);
  spice_node_2 n_pch1(eclk, ereset, pch1_port_2,pch1_port_1, pch1_v);
  spice_node_2 n_pch0(eclk, ereset, pch0_port_2,pch0_port_1, pch0_v);
  spice_node_2 n_op_T3_mem_zp_idx(eclk, ereset, op_T3_mem_zp_idx_port_7,op_T3_mem_zp_idx_port_5, op_T3_mem_zp_idx_v);
  spice_node_2 n_notalucin(eclk, ereset, notalucin_port_2,notalucin_port_4, notalucin_v);
  spice_node_2 n_dpc13_ORS(eclk, ereset, dpc13_ORS_port_8,dpc13_ORS_port_5, dpc13_ORS_v);
  spice_node_2 n_n_1069(eclk, ereset, n_1069_port_3,n_1069_port_4, n_1069_v);
  spice_node_2 n_n_1067(eclk, ereset, n_1067_port_2,n_1067_port_0, n_1067_v);
  spice_node_2 n_n_1065(eclk, ereset, n_1065_port_2,n_1065_port_1, n_1065_v);
  spice_node_4 n_n_1063(eclk, ereset, n_1063_port_2,n_1063_port_7,n_1063_port_4,n_1063_port_5, n_1063_v);
  spice_node_2 n_op_T0_tay(eclk, ereset, op_T0_tay_port_9,op_T0_tay_port_11, op_T0_tay_v);
  spice_node_2 n_op_T0_tax(eclk, ereset, op_T0_tax_port_9,op_T0_tax_port_10, op_T0_tax_v);
  spice_node_2 n_n_1608(eclk, ereset, n_1608_port_2,n_1608_port_1, n_1608_v);
  spice_node_2 n_n_1609(eclk, ereset, n_1609_port_3,n_1609_port_0, n_1609_v);
  spice_node_3 n_n_1605(eclk, ereset, n_1605_port_3,n_1605_port_0,n_1605_port_5, n_1605_v);
  spice_node_2 n_op_T0_brk_rti(eclk, ereset, op_T0_brk_rti_port_8,op_T0_brk_rti_port_9, op_T0_brk_rti_v);
  spice_node_2 n_n_249(eclk, ereset, n_249_port_3,n_249_port_0, n_249_v);
  spice_node_2 n_n_718(eclk, ereset, n_718_port_2,n_718_port_1, n_718_v);
  spice_node_4 n_n_719(eclk, ereset, n_719_port_2,n_719_port_3,n_719_port_0,n_719_port_1, n_719_v);
  spice_node_2 n_n_717(eclk, ereset, n_717_port_4,n_717_port_5, n_717_v);
  spice_node_2 n_n_715(eclk, ereset, n_715_port_2,n_715_port_3, n_715_v);
  spice_node_2 n_n_241(eclk, ereset, n_241_port_2,n_241_port_3, n_241_v);
  spice_node_4 n_n_242(eclk, ereset, n_242_port_2,n_242_port_3,n_242_port_0,n_242_port_1, n_242_v);
  spice_node_2 n_n_243(eclk, ereset, n_243_port_2,n_243_port_1, n_243_v);
  spice_node_3 n_dasb7(eclk, ereset, dasb7_port_3,dasb7_port_1,dasb7_port_5, dasb7_v);
  spice_node_2 n_op_T5_rti_rts(eclk, ereset, op_T5_rti_rts_port_8,op_T5_rti_rts_port_10, op_T5_rti_rts_v);
  spice_node_2 n_n_669(eclk, ereset, n_669_port_3,n_669_port_4, n_669_v);
  spice_node_2 n__C23(eclk, ereset, _C23_port_2,_C23_port_3, _C23_v);
  spice_node_2 n_nnT2BR(eclk, ereset, nnT2BR_port_5,nnT2BR_port_10, nnT2BR_v);
  spice_node_2 n_n_1474(eclk, ereset, n_1474_port_2,n_1474_port_0, n_1474_v);
  spice_node_2 n_op_T4_ind_x(eclk, ereset, op_T4_ind_x_port_9,op_T4_ind_x_port_7, op_T4_ind_x_v);
  spice_node_2 n_op_T4_ind_y(eclk, ereset, op_T4_ind_y_port_8,op_T4_ind_y_port_6, op_T4_ind_y_v);
  spice_node_2 n_n_1295(eclk, ereset, n_1295_port_2,n_1295_port_3, n_1295_v);
  spice_node_2 n_n_1296(eclk, ereset, n_1296_port_2,n_1296_port_0, n_1296_v);
  spice_node_2 n_n_1290(eclk, ereset, n_1290_port_3,n_1290_port_5, n_1290_v);
  spice_node_2 n_n_1293(eclk, ereset, n_1293_port_6,n_1293_port_4, n_1293_v);
  spice_node_2 n_dpc7_SS(eclk, ereset, dpc7_SS_port_7,dpc7_SS_port_12, dpc7_SS_v);
  spice_node_2 n_op_T__iny_dey(eclk, ereset, op_T__iny_dey_port_8,op_T__iny_dey_port_9, op_T__iny_dey_v);
  spice_node_2 n_n_906(eclk, ereset, n_906_port_3,n_906_port_0, n_906_v);
  spice_node_2 n_n_905(eclk, ereset, n_905_port_2,n_905_port_3, n_905_v);
  spice_node_2 n_n_1356(eclk, ereset, n_1356_port_2,n_1356_port_0, n_1356_v);
  spice_node_2 n_n_1423(eclk, ereset, n_1423_port_3,n_1423_port_0, n_1423_v);
  spice_node_2 n_n_38(eclk, ereset, n_38_port_2,n_38_port_1, n_38_v);
  spice_node_2 n_n_1599(eclk, ereset, n_1599_port_2,n_1599_port_3, n_1599_v);
  spice_node_2 n_n_1041(eclk, ereset, n_1041_port_0,n_1041_port_1, n_1041_v);
  spice_node_2 n_n_1043(eclk, ereset, n_1043_port_2,n_1043_port_0, n_1043_v);
  spice_node_2 n_n_1596(eclk, ereset, n_1596_port_3,n_1596_port_0, n_1596_v);
  spice_node_2 n_n_1045(eclk, ereset, n_1045_port_3,n_1045_port_4, n_1045_v);
  spice_node_3 n_n_1046(eclk, ereset, n_1046_port_2,n_1046_port_3,n_1046_port_0, n_1046_v);
  spice_node_2 n_n_1595(eclk, ereset, n_1595_port_2,n_1595_port_1, n_1595_v);
  spice_node_2 n_n_1620(eclk, ereset, n_1620_port_3,n_1620_port_0, n_1620_v);
  spice_node_3 n_n_1621(eclk, ereset, n_1621_port_2,n_1621_port_0,n_1621_port_1, n_1621_v);
  spice_node_2 n_n_1629(eclk, ereset, n_1629_port_3,n_1629_port_4, n_1629_v);
  spice_node_2 n_n_228(eclk, ereset, n_228_port_2,n_228_port_0, n_228_v);
  spice_node_2 n_n_220(eclk, ereset, n_220_port_3,n_220_port_0, n_220_v);
  spice_node_2 n_n_221(eclk, ereset, n_221_port_2,n_221_port_1, n_221_v);
  spice_node_3 n_n_227(eclk, ereset, n_227_port_2,n_227_port_3,n_227_port_0, n_227_v);
  spice_node_2 n_n_224(eclk, ereset, n_224_port_4,n_224_port_5, n_224_v);
  spice_node_2 n_n_225(eclk, ereset, n_225_port_2,n_225_port_0, n_225_v);
  spice_node_2 n_op_T4_abs_idx(eclk, ereset, op_T4_abs_idx_port_6,op_T4_abs_idx_port_4, op_T4_abs_idx_v);
  spice_node_2 n_op_implied(eclk, ereset, op_implied_port_6,op_implied_port_5, op_implied_v);
  spice_node_2 n_n_735(eclk, ereset, n_735_port_3,n_735_port_4, n_735_v);
  spice_node_2 n_n_730(eclk, ereset, n_730_port_2,n_730_port_1, n_730_v);
  spice_node_2 n_n_732(eclk, ereset, n_732_port_8,n_732_port_4, n_732_v);
  spice_node_2 n_dpc22__DSA(eclk, ereset, dpc22__DSA_port_3,dpc22__DSA_port_0, dpc22__DSA_v);
  spice_node_2 n_n_739(eclk, ereset, n_739_port_9,n_739_port_4, n_739_v);
  spice_node_2 n_x2(eclk, ereset, x2_port_0,x2_port_1, x2_v);
  spice_node_2 n_x3(eclk, ereset, x3_port_0,x3_port_1, x3_v);
  spice_node_2 n_x0(eclk, ereset, x0_port_0,x0_port_1, x0_v);
  spice_node_2 n_x1(eclk, ereset, x1_port_0,x1_port_1, x1_v);
  spice_node_2 n_op_T__dex(eclk, ereset, op_T__dex_port_9,op_T__dex_port_10, op_T__dex_v);
  spice_node_2 n_x7(eclk, ereset, x7_port_2,x7_port_1, x7_v);
  spice_node_2 n_x4(eclk, ereset, x4_port_0,x4_port_1, x4_v);
  spice_node_2 n_x5(eclk, ereset, x5_port_2,x5_port_1, x5_v);
  spice_node_2 n__C01(eclk, ereset, _C01_port_2,_C01_port_3, _C01_v);
  spice_node_2 n_op_T0_sbc(eclk, ereset, op_T0_sbc_port_8,op_T0_sbc_port_9, op_T0_sbc_v);
  spice_node_2 n_n_410(eclk, ereset, n_410_port_6,n_410_port_5, n_410_v);
  spice_node_5 n_n_1458(eclk, ereset, n_1458_port_2,n_1458_port_3,n_1458_port_0,n_1458_port_1,n_1458_port_4, n_1458_v);
  spice_node_2 n_n_1457(eclk, ereset, n_1457_port_3,n_1457_port_4, n_1457_v);
  spice_node_2 n_n_1455(eclk, ereset, n_1455_port_9,n_1455_port_10, n_1455_v);
  spice_node_2 n_DA_AB2(eclk, ereset, DA_AB2_port_2,DA_AB2_port_3, DA_AB2_v);
  spice_node_2 n_n_692(eclk, ereset, n_692_port_4,n_692_port_5, n_692_v);
  spice_node_2 n_n_695(eclk, ereset, n_695_port_2,n_695_port_3, n_695_v);
  spice_node_5 n_n_694(eclk, ereset, n_694_port_2,n_694_port_3,n_694_port_0,n_694_port_1,n_694_port_4, n_694_v);
  spice_node_2 n_n_969(eclk, ereset, n_969_port_2,n_969_port_0, n_969_v);
  spice_node_2 n_n_961(eclk, ereset, n_961_port_2,n_961_port_0, n_961_v);
  spice_node_2 n_n_963(eclk, ereset, n_963_port_2,n_963_port_1, n_963_v);
  spice_node_2 n_n_962(eclk, ereset, n_962_port_2,n_962_port_1, n_962_v);
  spice_node_2 n_n_964(eclk, ereset, n_964_port_7,n_964_port_4, n_964_v);
  spice_node_2 n_n_966(eclk, ereset, n_966_port_3,n_966_port_0, n_966_v);
  spice_node_2 n_irline3(eclk, ereset, irline3_port_0,irline3_port_64, irline3_v);
  spice_node_2 n_pcl3(eclk, ereset, pcl3_port_2,pcl3_port_1, pcl3_v);
  spice_node_2 n_pcl2(eclk, ereset, pcl2_port_2,pcl2_port_1, pcl2_v);
  spice_node_2 n_pcl1(eclk, ereset, pcl1_port_2,pcl1_port_1, pcl1_v);
  spice_node_2 n_pcl0(eclk, ereset, pcl0_port_2,pcl0_port_1, pcl0_v);
  spice_node_2 n_pcl7(eclk, ereset, pcl7_port_2,pcl7_port_1, pcl7_v);
  spice_node_2 n_pcl6(eclk, ereset, pcl6_port_2,pcl6_port_1, pcl6_v);
  spice_node_2 n_pcl5(eclk, ereset, pcl5_port_2,pcl5_port_1, pcl5_v);
  spice_node_2 n_pcl4(eclk, ereset, pcl4_port_2,pcl4_port_1, pcl4_v);
  spice_node_2 n_dpc0_YSB(eclk, ereset, dpc0_YSB_port_3,dpc0_YSB_port_12, dpc0_YSB_v);
  spice_node_2 n_n_1026(eclk, ereset, n_1026_port_3,n_1026_port_0, n_1026_v);
  spice_node_2 n_n_1024(eclk, ereset, n_1024_port_3,n_1024_port_0, n_1024_v);
  spice_node_2 n_n_1025(eclk, ereset, n_1025_port_2,n_1025_port_1, n_1025_v);
  spice_node_2 n_alua6(eclk, ereset, alua6_port_0,alua6_port_1, alua6_v);
  spice_node_2 n_alua7(eclk, ereset, alua7_port_3,alua7_port_0, alua7_v);
  spice_node_2 n_alua4(eclk, ereset, alua4_port_0,alua4_port_1, alua4_v);
  spice_node_2 n_alua5(eclk, ereset, alua5_port_0,alua5_port_1, alua5_v);
  spice_node_2 n_alua2(eclk, ereset, alua2_port_0,alua2_port_1, alua2_v);
  spice_node_2 n_alua3(eclk, ereset, alua3_port_0,alua3_port_1, alua3_v);
  spice_node_2 n_alua0(eclk, ereset, alua0_port_0,alua0_port_1, alua0_v);
  spice_node_2 n_alua1(eclk, ereset, alua1_port_2,alua1_port_3, alua1_v);
  spice_node_2 n_n_1271(eclk, ereset, n_1271_port_2,n_1271_port_0, n_1271_v);
  spice_node_1 n_nmi(eclk, ereset, nmi_port_2, nmi_v);
  spice_node_2 n_op_T2_branch(eclk, ereset, op_T2_branch_port_6,op_T2_branch_port_7, op_T2_branch_v);
  spice_node_2 n_dpc41_DL_ADL(eclk, ereset, dpc41_DL_ADL_port_9,dpc41_DL_ADL_port_0, dpc41_DL_ADL_v);
  spice_node_2 n_n_200(eclk, ereset, n_200_port_7,n_200_port_5, n_200_v);
  spice_node_2 n_n_753(eclk, ereset, n_753_port_4,n_753_port_5, n_753_v);
  spice_node_2 n_n_757(eclk, ereset, n_757_port_2,n_757_port_5, n_757_v);
  spice_node_2 n_n_754(eclk, ereset, n_754_port_8,n_754_port_4, n_754_v);
  spice_node_2 n_n_207(eclk, ereset, n_207_port_3,n_207_port_5, n_207_v);
  spice_node_5 n_n_208(eclk, ereset, n_208_port_2,n_208_port_3,n_208_port_0,n_208_port_1,n_208_port_4, n_208_v);
  spice_node_5 n_n_209(eclk, ereset, n_209_port_2,n_209_port_3,n_209_port_0,n_209_port_1,n_209_port_4, n_209_v);
  spice_node_2 n__C67(eclk, ereset, _C67_port_3,_C67_port_0, _C67_v);
  spice_node_2 n_dpc37_PCLDB(eclk, ereset, dpc37_PCLDB_port_0,dpc37_PCLDB_port_4, dpc37_PCLDB_v);
  spice_node_2 n___AxB3__C23(eclk, ereset, __AxB3__C23_port_3,__AxB3__C23_port_4, __AxB3__C23_v);
  spice_node_2 n_pd5_clearIR(eclk, ereset, pd5_clearIR_port_3,pd5_clearIR_port_4, pd5_clearIR_v);
  spice_node_2 n_dpc12_0ADD(eclk, ereset, dpc12_0ADD_port_9,dpc12_0ADD_port_12, dpc12_0ADD_v);
  spice_node_2 n_dpc4_SSB(eclk, ereset, dpc4_SSB_port_9,dpc4_SSB_port_0, dpc4_SSB_v);
  spice_node_2 n_n_134(eclk, ereset, n_134_port_7,n_134_port_5, n_134_v);
  spice_node_2 n_n_947(eclk, ereset, n_947_port_2,n_947_port_1, n_947_v);
  spice_node_2 n_n_946(eclk, ereset, n_946_port_2,n_946_port_4, n_946_v);
  spice_node_2 n_n_417(eclk, ereset, n_417_port_0,n_417_port_1, n_417_v);
  spice_node_2 n_n_944(eclk, ereset, n_944_port_3,n_944_port_4, n_944_v);
  spice_node_2 n_op_T0_cpy_iny(eclk, ereset, op_T0_cpy_iny_port_9,op_T0_cpy_iny_port_7, op_T0_cpy_iny_v);
  spice_node_2 n_n_419(eclk, ereset, n_419_port_2,n_419_port_0, n_419_v);
  spice_node_2 n_y1(eclk, ereset, y1_port_2,y1_port_0, y1_v);
  spice_node_2 n_y0(eclk, ereset, y0_port_2,y0_port_0, y0_v);
  spice_node_2 n_y3(eclk, ereset, y3_port_2,y3_port_0, y3_v);
  spice_node_2 n_y2(eclk, ereset, y2_port_2,y2_port_0, y2_v);
  spice_node_2 n_y5(eclk, ereset, y5_port_0,y5_port_1, y5_v);
  spice_node_2 n_y4(eclk, ereset, y4_port_2,y4_port_0, y4_v);
  spice_node_2 n_y7(eclk, ereset, y7_port_0,y7_port_1, y7_v);
  spice_node_2 n_y6(eclk, ereset, y6_port_0,y6_port_1, y6_v);
  spice_node_2 n_n_1007(eclk, ereset, n_1007_port_2,n_1007_port_1, n_1007_v);
  spice_node_2 n_n_1002(eclk, ereset, n_1002_port_1,n_1002_port_5, n_1002_v);
  spice_node_2 n_abh5(eclk, ereset, abh5_port_3,abh5_port_4, abh5_v);
  spice_node_2 n_abh4(eclk, ereset, abh4_port_0,abh4_port_4, abh4_v);
  spice_node_2 n_abh7(eclk, ereset, abh7_port_0,abh7_port_4, abh7_v);
  spice_node_2 n_abh6(eclk, ereset, abh6_port_3,abh6_port_4, abh6_v);
  spice_node_2 n_abh1(eclk, ereset, abh1_port_3,abh1_port_4, abh1_v);
  spice_node_2 n_abh0(eclk, ereset, abh0_port_3,abh0_port_4, abh0_v);
  spice_node_2 n_abh3(eclk, ereset, abh3_port_3,abh3_port_4, abh3_v);
  spice_node_2 n_abh2(eclk, ereset, abh2_port_0,abh2_port_4, abh2_v);
  spice_node_2 n_n_1552(eclk, ereset, n_1552_port_2,n_1552_port_0, n_1552_v);
  spice_node_2 n_alucin(eclk, ereset, alucin_port_2,alucin_port_1, alucin_v);
  spice_node_2 n_x_op_push_pull(eclk, ereset, x_op_push_pull_port_8,x_op_push_pull_port_6, x_op_push_pull_v);
  spice_node_2 n_dpc11_SBADD(eclk, ereset, dpc11_SBADD_port_9,dpc11_SBADD_port_12, dpc11_SBADD_v);
  spice_node_2 n_dpc10_ADLADD(eclk, ereset, dpc10_ADLADD_port_5,dpc10_ADLADD_port_12, dpc10_ADLADD_v);
  spice_node_2 n_n_779(eclk, ereset, n_779_port_3,n_779_port_5, n_779_v);
  spice_node_2 n_n_770(eclk, ereset, n_770_port_3,n_770_port_1, n_770_v);
  spice_node_2 n_n_771(eclk, ereset, n_771_port_1,n_771_port_4, n_771_v);
  spice_node_2 n_n_772(eclk, ereset, n_772_port_2,n_772_port_3, n_772_v);
  spice_node_2 n_n_773(eclk, ereset, n_773_port_3,n_773_port_5, n_773_v);
  spice_node_2 n_n_774(eclk, ereset, n_774_port_2,n_774_port_0, n_774_v);
  spice_node_2 n_n_837(eclk, ereset, n_837_port_2,n_837_port_0, n_837_v);
  spice_node_2 n_op_T0_bit(eclk, ereset, op_T0_bit_port_8,op_T0_bit_port_10, op_T0_bit_v);
  spice_node_2 n_n_344(eclk, ereset, n_344_port_8,n_344_port_4, n_344_v);
  spice_node_2 n_n_834(eclk, ereset, n_834_port_2,n_834_port_4, n_834_v);
  spice_node_2 n_dpc29_0ADH17(eclk, ereset, dpc29_0ADH17_port_2,dpc29_0ADH17_port_1, dpc29_0ADH17_v);
  spice_node_2 n_dpc26_ACDB(eclk, ereset, dpc26_ACDB_port_0,dpc26_ACDB_port_12, dpc26_ACDB_v);
  spice_node_2 n__C45(eclk, ereset, _C45_port_1,_C45_port_4, _C45_v);
  spice_node_2 n_VEC0(eclk, ereset, VEC0_port_6,VEC0_port_5, VEC0_v);
  spice_node_2 n_VEC1(eclk, ereset, VEC1_port_3,VEC1_port_4, VEC1_v);
  spice_node_2 n_op_T4_rts(eclk, ereset, op_T4_rts_port_9,op_T4_rts_port_11, op_T4_rts_v);
  spice_node_3 n_n_430(eclk, ereset, n_430_port_2,n_430_port_3,n_430_port_1, n_430_v);
  spice_node_4 n_n_436(eclk, ereset, n_436_port_2,n_436_port_3,n_436_port_0,n_436_port_1, n_436_v);
  spice_node_2 n_op_T4_rti(eclk, ereset, op_T4_rti_port_9,op_T4_rti_port_10, op_T4_rti_v);
  spice_node_2 n_op_SRS(eclk, ereset, op_SRS_port_2,op_SRS_port_6, op_SRS_v);
  spice_node_2 n_n_1343(eclk, ereset, n_1343_port_3,n_1343_port_5, n_1343_v);
  spice_node_2 n_n_1345(eclk, ereset, n_1345_port_7,n_1345_port_5, n_1345_v);
  spice_node_2 n_n_1578(eclk, ereset, n_1578_port_2,n_1578_port_1, n_1578_v);
  spice_node_2 n_n_1573(eclk, ereset, n_1573_port_2,n_1573_port_0, n_1573_v);
  spice_node_2 n_DC78(eclk, ereset, DC78_port_7,DC78_port_4, DC78_v);
  spice_node_2 n_op_sta_cmp(eclk, ereset, op_sta_cmp_port_6,op_sta_cmp_port_5, op_sta_cmp_v);
  spice_node_2 n_op_SUMS(eclk, ereset, op_SUMS_port_6,op_SUMS_port_5, op_SUMS_v);
  spice_node_2 n_n_1688(eclk, ereset, n_1688_port_2,n_1688_port_0, n_1688_v);
  spice_node_3 n_n_404(eclk, ereset, n_404_port_2,n_404_port_6,n_404_port_5, n_404_v);
  spice_node_2 n_n_954(eclk, ereset, n_954_port_3,n_954_port_4, n_954_v);
  spice_node_2 n_n_400(eclk, ereset, n_400_port_2,n_400_port_3, n_400_v);
  spice_node_2 n_op_T4_brk_jsr(eclk, ereset, op_T4_brk_jsr_port_8,op_T4_brk_jsr_port_9, op_T4_brk_jsr_v);
  spice_node_2 n_n_1219(eclk, ereset, n_1219_port_2,n_1219_port_1, n_1219_v);
  spice_node_2 n_n_1215(eclk, ereset, n_1215_port_6,n_1215_port_5, n_1215_v);
  spice_node_2 n_n_1214(eclk, ereset, n_1214_port_2,n_1214_port_0, n_1214_v);
  spice_node_2 n_n_1211(eclk, ereset, n_1211_port_8,n_1211_port_9, n_1211_v);
  spice_node_2 n_n_1213(eclk, ereset, n_1213_port_3,n_1213_port_4, n_1213_v);
  spice_node_2 n_n_1655(eclk, ereset, n_1655_port_2,n_1655_port_1, n_1655_v);
  spice_node_2 n_pd2_clearIR(eclk, ereset, pd2_clearIR_port_6,pd2_clearIR_port_7, pd2_clearIR_v);
  spice_node_5 n_n_1654(eclk, ereset, n_1654_port_2,n_1654_port_3,n_1654_port_0,n_1654_port_1,n_1654_port_4, n_1654_v);
  spice_node_2 n_n_1657(eclk, ereset, n_1657_port_2,n_1657_port_3, n_1657_v);
  spice_node_2 n_n_1650(eclk, ereset, n_1650_port_2,n_1650_port_0, n_1650_v);
  spice_node_2 n_n_182(eclk, ereset, n_182_port_7,n_182_port_11, n_182_v);
  spice_node_2 n_n_180(eclk, ereset, n_180_port_3,n_180_port_5, n_180_v);
  spice_node_2 n_n_184(eclk, ereset, n_184_port_2,n_184_port_0, n_184_v);
  spice_node_3 n_n_635(eclk, ereset, n_635_port_3,n_635_port_0,n_635_port_1, n_635_v);
  spice_node_2 n_n_634(eclk, ereset, n_634_port_0,n_634_port_1, n_634_v);
  spice_node_2 n_n_637(eclk, ereset, n_637_port_3,n_637_port_4, n_637_v);
  spice_node_2 n_n_636(eclk, ereset, n_636_port_2,n_636_port_0, n_636_v);
  spice_node_2 n_n_631(eclk, ereset, n_631_port_2,n_631_port_3, n_631_v);
  spice_node_2 n_n_630(eclk, ereset, n_630_port_3,n_630_port_0, n_630_v);
  spice_node_1 n_n_633(eclk, ereset, n_633_port_0, n_633_v);
  spice_node_2 n_n_632(eclk, ereset, n_632_port_3,n_632_port_5, n_632_v);
  spice_node_3 n_n_458(eclk, ereset, n_458_port_2,n_458_port_0,n_458_port_1, n_458_v);
  spice_node_2 n_n_988(eclk, ereset, n_988_port_3,n_988_port_1, n_988_v);
  spice_node_2 n_n_983(eclk, ereset, n_983_port_2,n_983_port_1, n_983_v);
  spice_node_2 n_n_981(eclk, ereset, n_981_port_2,n_981_port_1, n_981_v);
  spice_node_2 n_n_987(eclk, ereset, n_987_port_2,n_987_port_1, n_987_v);
  spice_node_2 n_n_986(eclk, ereset, n_986_port_2,n_986_port_3, n_986_v);
  spice_node_2 n_n_457(eclk, ereset, n_457_port_2,n_457_port_1, n_457_v);
  spice_node_2 n_op_T0_lda(eclk, ereset, op_T0_lda_port_9,op_T0_lda_port_7, op_T0_lda_v);
  spice_node_2 n_abl1(eclk, ereset, abl1_port_3,abl1_port_4, abl1_v);
  spice_node_2 n_abl0(eclk, ereset, abl0_port_3,abl0_port_4, abl0_v);
  spice_node_2 n_abl4(eclk, ereset, abl4_port_0,abl4_port_4, abl4_v);
  spice_node_2 n_op_T3_plp_pla(eclk, ereset, op_T3_plp_pla_port_8,op_T3_plp_pla_port_10, op_T3_plp_pla_v);
  spice_node_2 n_n_1517(eclk, ereset, n_1517_port_3,n_1517_port_4, n_1517_v);
  spice_node_2 n_n_1518(eclk, ereset, n_1518_port_2,n_1518_port_1, n_1518_v);
  spice_node_3 n_n_1519(eclk, ereset, n_1519_port_2,n_1519_port_3,n_1519_port_0, n_1519_v);
  spice_node_2 n_n_279(eclk, ereset, n_279_port_4,n_279_port_5, n_279_v);
  spice_node_2 n_n_846(eclk, ereset, n_846_port_3,n_846_port_1, n_846_v);
  spice_node_2 n_n_847(eclk, ereset, n_847_port_2,n_847_port_1, n_847_v);
  spice_node_2 n_n_844(eclk, ereset, n_844_port_6,n_844_port_5, n_844_v);
  spice_node_2 n_n_845(eclk, ereset, n_845_port_8,n_845_port_4, n_845_v);
  spice_node_2 n_n_842(eclk, ereset, n_842_port_3,n_842_port_0, n_842_v);
  spice_node_2 n_op_T3_jmp(eclk, ereset, op_T3_jmp_port_8,op_T3_jmp_port_9, op_T3_jmp_v);
  spice_node_2 n_n_849(eclk, ereset, n_849_port_2,n_849_port_0, n_849_v);
  spice_node_2 n___AxB5__C45(eclk, ereset, __AxB5__C45_port_3,__AxB5__C45_port_4, __AxB5__C45_v);
  spice_node_2 n_dpc16_EORS(eclk, ereset, dpc16_EORS_port_8,dpc16_EORS_port_9, dpc16_EORS_v);
  spice_node_2 n_n_1231(eclk, ereset, n_1231_port_2,n_1231_port_1, n_1231_v);
  spice_node_2 n_n_1230(eclk, ereset, n_1230_port_4,n_1230_port_5, n_1230_v);
  spice_node_2 n_n_1238(eclk, ereset, n_1238_port_2,n_1238_port_1, n_1238_v);
  spice_node_5 n_n_1722(eclk, ereset, n_1722_port_2,n_1722_port_3,n_1722_port_0,n_1722_port_1,n_1722_port_4, n_1722_v);
  spice_node_2 n_op_branch_done(eclk, ereset, op_branch_done_port_8,op_branch_done_port_9, op_branch_done_v);
  spice_node_2 n_aluvout(eclk, ereset, aluvout_port_2,aluvout_port_0, aluvout_v);
  spice_node_5 n_n_618(eclk, ereset, n_618_port_2,n_618_port_3,n_618_port_0,n_618_port_1,n_618_port_4, n_618_v);
  spice_node_2 n_n_613(eclk, ereset, n_613_port_4,n_613_port_10, n_613_v);
  spice_node_2 n_n_612(eclk, ereset, n_612_port_0,n_612_port_4, n_612_v);
  spice_node_2 n_n_611(eclk, ereset, n_611_port_4,n_611_port_5, n_611_v);
  spice_node_2 n_n_617(eclk, ereset, n_617_port_3,n_617_port_0, n_617_v);
  spice_node_2 n_n_616(eclk, ereset, n_616_port_6,n_616_port_5, n_616_v);
  spice_node_2 n_n_1137(eclk, ereset, n_1137_port_2,n_1137_port_4, n_1137_v);
  spice_node_2 n_n_620(eclk, ereset, n_620_port_6,n_620_port_7, n_620_v);
  spice_node_3 n_n_884(eclk, ereset, n_884_port_2,n_884_port_0,n_884_port_1, n_884_v);
  spice_node_3 n_Pout0(eclk, ereset, Pout0_port_2,Pout0_port_0,Pout0_port_1, Pout0_v);
  spice_node_2 n_n_1545(eclk, ereset, n_1545_port_2,n_1545_port_1, n_1545_v);
  spice_node_2 n_n_1010(eclk, ereset, n_1010_port_3,n_1010_port_0, n_1010_v);
  spice_node_2 n_n_1017(eclk, ereset, n_1017_port_2,n_1017_port_0, n_1017_v);
  spice_node_2 n_n_1542(eclk, ereset, n_1542_port_6,n_1542_port_4, n_1542_v);
  spice_node_2 n_dpc19_ADDSB7(eclk, ereset, dpc19_ADDSB7_port_2,dpc19_ADDSB7_port_0, dpc19_ADDSB7_v);
  spice_node_4 n_n_477(eclk, ereset, n_477_port_3,n_477_port_1,n_477_port_4,n_477_port_5, n_477_v);
  spice_node_2 n_n_476(eclk, ereset, n_476_port_4,n_476_port_5, n_476_v);
  spice_node_2 n_n_475(eclk, ereset, n_475_port_2,n_475_port_0, n_475_v);
  spice_node_2 n_n_474(eclk, ereset, n_474_port_3,n_474_port_5, n_474_v);
  spice_node_2 n_n_473(eclk, ereset, n_473_port_2,n_473_port_3, n_473_v);
  spice_node_2 n_n_472(eclk, ereset, n_472_port_3,n_472_port_6, n_472_v);
  spice_node_2 n_n_471(eclk, ereset, n_471_port_3,n_471_port_4, n_471_v);
  spice_node_2 n_n_470(eclk, ereset, n_470_port_2,n_470_port_3, n_470_v);
  spice_node_2 n_n_479(eclk, ereset, n_479_port_3,n_479_port_4, n_479_v);
  spice_node_3 n_n_478(eclk, ereset, n_478_port_2,n_478_port_0,n_478_port_1, n_478_v);
  spice_node_2 n_brk_done(eclk, ereset, brk_done_port_9,brk_done_port_12, brk_done_v);
  spice_node_2 n_op_T0_txa(eclk, ereset, op_T0_txa_port_9,op_T0_txa_port_11, op_T0_txa_v);
  spice_node_3 n_p6(eclk, ereset, p6_port_2,p6_port_0,p6_port_1, p6_v);
  spice_node_3 n_p7(eclk, ereset, p7_port_2,p7_port_0,p7_port_1, p7_v);
  spice_node_2 n_DC34(eclk, ereset, DC34_port_9,DC34_port_4, DC34_v);
  spice_node_2 n_op_T2_stack(eclk, ereset, op_T2_stack_port_8,op_T2_stack_port_7, op_T2_stack_v);
  spice_node_2 n_n_1534(eclk, ereset, n_1534_port_4,n_1534_port_5, n_1534_v);
  spice_node_4 n_n_1531(eclk, ereset, n_1531_port_2,n_1531_port_3,n_1531_port_0,n_1531_port_1, n_1531_v);
  spice_node_2 n_n_1391(eclk, ereset, n_1391_port_3,n_1391_port_4, n_1391_v);
  spice_node_2 n_n_1392(eclk, ereset, n_1392_port_2,n_1392_port_3, n_1392_v);
  spice_node_3 n_n_1398(eclk, ereset, n_1398_port_8,n_1398_port_1,n_1398_port_6, n_1398_v);
  spice_node_2 n_n_1399(eclk, ereset, n_1399_port_3,n_1399_port_0, n_1399_v);
  spice_node_2 n_n_288(eclk, ereset, n_288_port_6,n_288_port_4, n_288_v);
  spice_node_5 n_n_280(eclk, ereset, n_280_port_2,n_280_port_3,n_280_port_0,n_280_port_1,n_280_port_4, n_280_v);
  spice_node_2 n_n_282(eclk, ereset, n_282_port_2,n_282_port_1, n_282_v);
  spice_node_2 n_n_284(eclk, ereset, n_284_port_2,n_284_port_0, n_284_v);
  spice_node_2 n_n_135(eclk, ereset, n_135_port_2,n_135_port_1, n_135_v);
  spice_node_2 n_n_133(eclk, ereset, n_133_port_4,n_133_port_5, n_133_v);
  spice_node_2 n_n_130(eclk, ereset, n_130_port_2,n_130_port_0, n_130_v);
  spice_node_3 n_n_869(eclk, ereset, n_869_port_2,n_869_port_3,n_869_port_1, n_869_v);
  spice_node_0 n_n_866(eclk, ereset,  n_866_v);
  spice_node_2 n_n_867(eclk, ereset, n_867_port_3,n_867_port_4, n_867_v);
  spice_node_2 n_n_861(eclk, ereset, n_861_port_2,n_861_port_0, n_861_v);
  spice_node_2 n_n_862(eclk, ereset, n_862_port_9,n_862_port_4, n_862_v);
  spice_node_4 n_n_350(eclk, ereset, n_350_port_3,n_350_port_1,n_350_port_4,n_350_port_5, n_350_v);
  spice_node_2 n_dpc17_SUMS(eclk, ereset, dpc17_SUMS_port_0,dpc17_SUMS_port_1, dpc17_SUMS_v);
  spice_node_2 n__op_branch_done(eclk, ereset, _op_branch_done_port_2,_op_branch_done_port_0, _op_branch_done_v);
  spice_node_2 n_op_T0_acc(eclk, ereset, op_T0_acc_port_3,op_T0_acc_port_4, op_T0_acc_v);
  spice_node_2 n_BRtaken(eclk, ereset, BRtaken_port_4,BRtaken_port_10, BRtaken_v);
  spice_node_4 n_n_1251(eclk, ereset, n_1251_port_2,n_1251_port_3,n_1251_port_0,n_1251_port_1, n_1251_v);
  spice_node_2 n_n_1253(eclk, ereset, n_1253_port_7,n_1253_port_5, n_1253_v);
  spice_node_2 n_n_1257(eclk, ereset, n_1257_port_7,n_1257_port_5, n_1257_v);
  spice_node_2 n_n_1258(eclk, ereset, n_1258_port_7,n_1258_port_4, n_1258_v);
  spice_node_4 n_n_1709(eclk, ereset, n_1709_port_2,n_1709_port_3,n_1709_port_0,n_1709_port_1, n_1709_v);
  spice_node_2 n_n_1708(eclk, ereset, n_1708_port_3,n_1708_port_4, n_1708_v);
  spice_node_2 n_dpc3_SBX(eclk, ereset, dpc3_SBX_port_9,dpc3_SBX_port_12, dpc3_SBX_v);
  spice_node_2 n_op_T2_php(eclk, ereset, op_T2_php_port_9,op_T2_php_port_10, op_T2_php_v);
  spice_node_2 n_op_T2_pha(eclk, ereset, op_T2_pha_port_9,op_T2_pha_port_10, op_T2_pha_v);
  spice_node_2 n_dpc31_PCHPCH(eclk, ereset, dpc31_PCHPCH_port_11,dpc31_PCHPCH_port_12, dpc31_PCHPCH_v);
  spice_node_2 n_n_670(eclk, ereset, n_670_port_2,n_670_port_3, n_670_v);
  spice_node_2 n_n_673(eclk, ereset, n_673_port_2,n_673_port_4, n_673_v);
  spice_node_2 n_n_674(eclk, ereset, n_674_port_2,n_674_port_0, n_674_v);
  spice_node_3 n_n_676(eclk, ereset, n_676_port_2,n_676_port_3,n_676_port_0, n_676_v);
  spice_node_2 n_n_678(eclk, ereset, n_678_port_4,n_678_port_5, n_678_v);
  spice_node_3 n_Pout1(eclk, ereset, Pout1_port_2,Pout1_port_0,Pout1_port_1, Pout1_v);
  spice_node_3 n_Pout3(eclk, ereset, Pout3_port_2,Pout3_port_3,Pout3_port_4, Pout3_v);
  spice_node_3 n_Pout2(eclk, ereset, Pout2_port_2,Pout2_port_0,Pout2_port_1, Pout2_v);
  spice_node_2 n_n_499(eclk, ereset, n_499_port_3,n_499_port_0, n_499_v);
  spice_node_3 n_n_494(eclk, ereset, n_494_port_2,n_494_port_3,n_494_port_1, n_494_v);
  spice_node_2 n_n_496(eclk, ereset, n_496_port_2,n_496_port_1, n_496_v);
  spice_node_2 n_n_491(eclk, ereset, n_491_port_2,n_491_port_1, n_491_v);
  spice_node_2 n_n_490(eclk, ereset, n_490_port_2,n_490_port_1, n_490_v);
  spice_node_2 n_pd7_clearIR(eclk, ereset, pd7_clearIR_port_4,pd7_clearIR_port_5, pd7_clearIR_v);
  spice_node_2 n_n_1401(eclk, ereset, n_1401_port_2,n_1401_port_0, n_1401_v);
  spice_node_2 n_op_T4_jmp(eclk, ereset, op_T4_jmp_port_9,op_T4_jmp_port_11, op_T4_jmp_v);
  spice_node_2 n_n_19(eclk, ereset, n_19_port_3,n_19_port_4, n_19_v);
  spice_node_2 n_n_1117(eclk, ereset, n_1117_port_2,n_1117_port_1, n_1117_v);
  spice_node_2 n_n_1115(eclk, ereset, n_1115_port_3,n_1115_port_4, n_1115_v);
  spice_node_2 n_n_1110(eclk, ereset, n_1110_port_3,n_1110_port_1, n_1110_v);
  spice_node_2 n_n_1111(eclk, ereset, n_1111_port_3,n_1111_port_6, n_1111_v);
  spice_node_2 n_n_803(eclk, ereset, n_803_port_2,n_803_port_0, n_803_v);
  spice_node_2 n_n_800(eclk, ereset, n_800_port_2,n_800_port_0, n_800_v);
  spice_node_0 n_n_806(eclk, ereset,  n_806_v);
  spice_node_2 n_n_807(eclk, ereset, n_807_port_3,n_807_port_5, n_807_v);
  spice_node_2 n_n_432(eclk, ereset, n_432_port_2,n_432_port_3, n_432_v);
  spice_node_2 n_n_1277(eclk, ereset, n_1277_port_3,n_1277_port_0, n_1277_v);
  spice_node_2 n_n_1275(eclk, ereset, n_1275_port_4,n_1275_port_5, n_1275_v);
  spice_node_2 n_n_1660(eclk, ereset, n_1660_port_3,n_1660_port_0, n_1660_v);
  spice_node_2 n_op_inc_nop(eclk, ereset, op_inc_nop_port_6,op_inc_nop_port_5, op_inc_nop_v);
  spice_node_2 n_n_128(eclk, ereset, n_128_port_2,n_128_port_0, n_128_v);
  spice_node_3 n_n_659(eclk, ereset, n_659_port_2,n_659_port_3,n_659_port_1, n_659_v);
  spice_node_4 n_n_658(eclk, ereset, n_658_port_2,n_658_port_3,n_658_port_0,n_658_port_1, n_658_v);
  spice_node_2 n_n_127(eclk, ereset, n_127_port_4,n_127_port_5, n_127_v);
  spice_node_5 n_n_652(eclk, ereset, n_652_port_2,n_652_port_3,n_652_port_0,n_652_port_1,n_652_port_4, n_652_v);
  spice_node_3 n_n_123(eclk, ereset, n_123_port_2,n_123_port_3,n_123_port_0, n_123_v);
  spice_node_2 n_n_122(eclk, ereset, n_122_port_2,n_122_port_0, n_122_v);
  spice_node_2 n_op_T0_shift_right_a(eclk, ereset, op_T0_shift_right_a_port_8,op_T0_shift_right_a_port_9, op_T0_shift_right_a_v);
  spice_node_2 n_op_T0_adc_sbc(eclk, ereset, op_T0_adc_sbc_port_8,op_T0_adc_sbc_port_6, op_T0_adc_sbc_v);
  spice_node_2 n_op_push_pull(eclk, ereset, op_push_pull_port_8,op_push_pull_port_7, op_push_pull_v);
  spice_node_2 n_n_1130(eclk, ereset, n_1130_port_8,n_1130_port_7, n_1130_v);
  spice_node_2 n_n_1133(eclk, ereset, n_1133_port_3,n_1133_port_4, n_1133_v);
  spice_node_2 n_n_1135(eclk, ereset, n_1135_port_2,n_1135_port_3, n_1135_v);
  spice_node_2 n_n_1138(eclk, ereset, n_1138_port_2,n_1138_port_0, n_1138_v);
  spice_node_2 n_op_T2_mem_zp(eclk, ereset, op_T2_mem_zp_port_7,op_T2_mem_zp_port_5, op_T2_mem_zp_v);
  spice_node_2 n_n_355(eclk, ereset, n_355_port_3,n_355_port_0, n_355_v);
  spice_node_2 n_n_824(eclk, ereset, n_824_port_6,n_824_port_5, n_824_v);
  spice_node_2 n_n_826(eclk, ereset, n_826_port_2,n_826_port_1, n_826_v);
  spice_node_3 n_n_351(eclk, ereset, n_351_port_2,n_351_port_0,n_351_port_1, n_351_v);
  spice_node_2 n_dpc9_DBADD(eclk, ereset, dpc9_DBADD_port_1,dpc9_DBADD_port_12, dpc9_DBADD_v);
  spice_node_2 n_n_358(eclk, ereset, n_358_port_2,n_358_port_4, n_358_v);
  spice_node_3 n_n_359(eclk, ereset, n_359_port_2,n_359_port_0,n_359_port_1, n_359_v);
  spice_node_2 n_dpc33_PCHDB(eclk, ereset, dpc33_PCHDB_port_0,dpc33_PCHDB_port_1, dpc33_PCHDB_v);
  spice_node_2 n_INTG(eclk, ereset, INTG_port_6,INTG_port_4, INTG_v);
  spice_node_2 n_n_755(eclk, ereset, n_755_port_3,n_755_port_0, n_755_v);
  spice_node_2 n_op_T2_ind(eclk, ereset, op_T2_ind_port_6,op_T2_ind_port_5, op_T2_ind_v);
  spice_node_2 n_op_rti_rts(eclk, ereset, op_rti_rts_port_9,op_rti_rts_port_10, op_rti_rts_v);
  spice_node_2 n_dpc8_nDBADD(eclk, ereset, dpc8_nDBADD_port_6,dpc8_nDBADD_port_12, dpc8_nDBADD_v);
  spice_node_2 n_n_109(eclk, ereset, n_109_port_2,n_109_port_0, n_109_v);
  spice_node_2 n_n_108(eclk, ereset, n_108_port_2,n_108_port_1, n_108_v);
  spice_node_2 n_n_102(eclk, ereset, n_102_port_2,n_102_port_0, n_102_v);
  spice_node_2 n_n_105(eclk, ereset, n_105_port_2,n_105_port_3, n_105_v);
  spice_node_2 n_n_104(eclk, ereset, n_104_port_6,n_104_port_7, n_104_v);
  spice_node_2 n_n_1575(eclk, ereset, n_1575_port_4,n_1575_port_5, n_1575_v);
  spice_node_2 n_dpc39_PCLPCL(eclk, ereset, dpc39_PCLPCL_port_11,dpc39_PCLPCL_port_12, dpc39_PCLPCL_v);
  spice_node_2 n_ADH_ABH(eclk, ereset, ADH_ABH_port_7,ADH_ABH_port_4, ADH_ABH_v);
  spice_node_2 n_Reset0(eclk, ereset, Reset0_port_4,Reset0_port_5, Reset0_v);
  spice_node_2 n_dpc25_SBDB(eclk, ereset, dpc25_SBDB_port_9,dpc25_SBDB_port_0, dpc25_SBDB_v);
  spice_node_2 n_n_1541(eclk, ereset, n_1541_port_4,n_1541_port_5, n_1541_v);
  spice_node_2 n_dpc23_SBAC(eclk, ereset, dpc23_SBAC_port_11,dpc23_SBAC_port_12, dpc23_SBAC_v);
  spice_node_2 n_n_1484(eclk, ereset, n_1484_port_2,n_1484_port_0, n_1484_v);
  spice_node_2 n_x_op_jmp(eclk, ereset, x_op_jmp_port_8,x_op_jmp_port_9, x_op_jmp_v);
  spice_node_2 n_n_1339(eclk, ereset, n_1339_port_2,n_1339_port_1, n_1339_v);
  spice_node_2 n_n_1488(eclk, ereset, n_1488_port_3,n_1488_port_0, n_1488_v);
  spice_node_2 n_n_1335(eclk, ereset, n_1335_port_2,n_1335_port_0, n_1335_v);
  spice_node_2 n_n_1159(eclk, ereset, n_1159_port_3,n_1159_port_4, n_1159_v);
  spice_node_2 n_n_1152(eclk, ereset, n_1152_port_2,n_1152_port_0, n_1152_v);
  spice_node_2 n_n_1157(eclk, ereset, n_1157_port_2,n_1157_port_0, n_1157_v);
  spice_node_2 n_n_1154(eclk, ereset, n_1154_port_3,n_1154_port_5, n_1154_v);
  spice_node_2 n__t2(eclk, ereset, _t2_port_0,_t2_port_21, _t2_v);
  spice_node_2 n__t3(eclk, ereset, _t3_port_15,_t3_port_16, _t3_v);
  spice_node_2 n_n_595(eclk, ereset, n_595_port_4,n_595_port_5, n_595_v);
  spice_node_2 n__t4(eclk, ereset, _t4_port_0,_t4_port_13, _t4_v);
  spice_node_2 n__t5(eclk, ereset, _t5_port_0,_t5_port_10, _t5_v);
  spice_node_2 n_n_1682(eclk, ereset, n_1682_port_2,n_1682_port_1, n_1682_v);
  spice_node_2 n_n_378(eclk, ereset, n_378_port_4,n_378_port_5, n_378_v);
  spice_node_2 n_n_374(eclk, ereset, n_374_port_2,n_374_port_1, n_374_v);
  spice_node_2 n_n_372(eclk, ereset, n_372_port_2,n_372_port_0, n_372_v);
  spice_node_2 n_n_373(eclk, ereset, n_373_port_0,n_373_port_4, n_373_v);
  spice_node_2 n_x_op_T0_txa(eclk, ereset, x_op_T0_txa_port_9,x_op_T0_txa_port_11, x_op_T0_txa_v);
  spice_node_2 n_C01(eclk, ereset, C01_port_8,C01_port_4, C01_v);
  spice_node_2 n_op_store(eclk, ereset, op_store_port_4,op_store_port_5, op_store_v);
  spice_node_2 n_n_1687(eclk, ereset, n_1687_port_2,n_1687_port_1, n_1687_v);
  spice_node_2 n_ab0(eclk, ereset, ab0_port_0,ab0_port_1, ab0_v);
  spice_node_2 n_ab1(eclk, ereset, ab1_port_0,ab1_port_1, ab1_v);
  spice_node_2 n_ab2(eclk, ereset, ab2_port_0,ab2_port_1, ab2_v);
  spice_node_2 n_ab3(eclk, ereset, ab3_port_0,ab3_port_1, ab3_v);
  spice_node_2 n_ab4(eclk, ereset, ab4_port_0,ab4_port_1, ab4_v);
  spice_node_2 n_ab5(eclk, ereset, ab5_port_0,ab5_port_1, ab5_v);
  spice_node_2 n_ab6(eclk, ereset, ab6_port_0,ab6_port_1, ab6_v);
  spice_node_2 n_ab7(eclk, ereset, ab7_port_0,ab7_port_1, ab7_v);
  spice_node_2 n_ab8(eclk, ereset, ab8_port_0,ab8_port_1, ab8_v);
  spice_node_2 n_ab9(eclk, ereset, ab9_port_0,ab9_port_1, ab9_v);
  spice_node_2 n_n_80(eclk, ereset, n_80_port_3,n_80_port_4, n_80_v);
  spice_node_2 n_n_83(eclk, ereset, n_83_port_3,n_83_port_0, n_83_v);
  spice_node_4 n_n_87(eclk, ereset, n_87_port_2,n_87_port_3,n_87_port_0,n_87_port_1, n_87_v);
  spice_node_3 n_n_86(eclk, ereset, n_86_port_2,n_86_port_3,n_86_port_0, n_86_v);
  spice_node_2 n_n_1684(eclk, ereset, n_1684_port_2,n_1684_port_1, n_1684_v);
  spice_node_2 n_n_161(eclk, ereset, n_161_port_4,n_161_port_5, n_161_v);
  spice_node_2 n_n_160(eclk, ereset, n_160_port_3,n_160_port_4, n_160_v);
  spice_node_2 n_n_163(eclk, ereset, n_163_port_2,n_163_port_3, n_163_v);
  spice_node_2 n_n_169(eclk, ereset, n_169_port_3,n_169_port_4, n_169_v);
  spice_node_3 n_n_168(eclk, ereset, n_168_port_2,n_168_port_3,n_168_port_0, n_168_v);
  spice_node_2 n_n_781(eclk, ereset, n_781_port_9,n_781_port_13, n_781_v);
  spice_node_2 n_n_783(eclk, ereset, n_783_port_3,n_783_port_4, n_783_v);
  spice_node_2 n_n_782(eclk, ereset, n_782_port_2,n_782_port_4, n_782_v);
  spice_node_2 n_n_789(eclk, ereset, n_789_port_2,n_789_port_0, n_789_v);
  spice_node_12 n_sb2(eclk, ereset, sb2_port_8,sb2_port_9,sb2_port_2,sb2_port_3,sb2_port_0,sb2_port_1,sb2_port_6,sb2_port_7,sb2_port_4,sb2_port_10,sb2_port_11,sb2_port_12, sb2_v);
  spice_node_12 n_sb3(eclk, ereset, sb3_port_8,sb3_port_9,sb3_port_2,sb3_port_3,sb3_port_0,sb3_port_1,sb3_port_6,sb3_port_7,sb3_port_4,sb3_port_5,sb3_port_10,sb3_port_11, sb3_v);
  spice_node_13 n_sb0(eclk, ereset, sb0_port_8,sb0_port_9,sb0_port_2,sb0_port_3,sb0_port_0,sb0_port_1,sb0_port_6,sb0_port_7,sb0_port_4,sb0_port_5,sb0_port_10,sb0_port_11,sb0_port_12, sb0_v);
  spice_node_12 n_sb1(eclk, ereset, sb1_port_8,sb1_port_9,sb1_port_2,sb1_port_0,sb1_port_1,sb1_port_6,sb1_port_7,sb1_port_4,sb1_port_5,sb1_port_10,sb1_port_11,sb1_port_12, sb1_v);
  spice_node_12 n_sb6(eclk, ereset, sb6_port_8,sb6_port_9,sb6_port_2,sb6_port_3,sb6_port_0,sb6_port_1,sb6_port_6,sb6_port_7,sb6_port_4,sb6_port_10,sb6_port_11,sb6_port_12, sb6_v);
  spice_node_12 n_sb7(eclk, ereset, sb7_port_8,sb7_port_9,sb7_port_2,sb7_port_3,sb7_port_0,sb7_port_1,sb7_port_6,sb7_port_7,sb7_port_4,sb7_port_5,sb7_port_10,sb7_port_11, sb7_v);
  spice_node_13 n_sb4(eclk, ereset, sb4_port_8,sb4_port_9,sb4_port_2,sb4_port_3,sb4_port_0,sb4_port_1,sb4_port_6,sb4_port_7,sb4_port_4,sb4_port_5,sb4_port_10,sb4_port_11,sb4_port_12, sb4_v);
  spice_node_12 n_sb5(eclk, ereset, sb5_port_8,sb5_port_2,sb5_port_3,sb5_port_0,sb5_port_1,sb5_port_6,sb5_port_7,sb5_port_4,sb5_port_5,sb5_port_10,sb5_port_11,sb5_port_12, sb5_v);
  spice_node_3 n___AxB_6(eclk, ereset, __AxB_6_port_2,__AxB_6_port_6,__AxB_6_port_11, __AxB_6_v);
  spice_node_3 n___AxB_4(eclk, ereset, __AxB_4_port_0,__AxB_4_port_6,__AxB_4_port_4, __AxB_4_v);
  spice_node_3 n___AxB_2(eclk, ereset, __AxB_2_port_0,__AxB_2_port_7,__AxB_2_port_4, __AxB_2_v);
  spice_node_3 n___AxB_0(eclk, ereset, __AxB_0_port_2,__AxB_0_port_6,__AxB_0_port_4, __AxB_0_v);
  spice_node_4 n_n_1318(eclk, ereset, n_1318_port_2,n_1318_port_3,n_1318_port_7,n_1318_port_5, n_1318_v);
  spice_node_2 n_n_1319(eclk, ereset, n_1319_port_2,n_1319_port_0, n_1319_v);
  spice_node_2 n_n_1312(eclk, ereset, n_1312_port_3,n_1312_port_5, n_1312_v);
  spice_node_2 n_n_1315(eclk, ereset, n_1315_port_3,n_1315_port_0, n_1315_v);
  spice_node_2 n_n_1316(eclk, ereset, n_1316_port_7,n_1316_port_5, n_1316_v);
  spice_node_2 n_dpc2_XSB(eclk, ereset, dpc2_XSB_port_2,dpc2_XSB_port_12, dpc2_XSB_v);
  spice_node_2 n_n_1175(eclk, ereset, n_1175_port_3,n_1175_port_1, n_1175_v);
  spice_node_2 n_n_1170(eclk, ereset, n_1170_port_3,n_1170_port_4, n_1170_v);
  spice_node_2 n_n_1178(eclk, ereset, n_1178_port_6,n_1178_port_5, n_1178_v);
  spice_node_2 n_n_1179(eclk, ereset, n_1179_port_3,n_1179_port_4, n_1179_v);
  spice_node_4 n_n_578(eclk, ereset, n_578_port_2,n_578_port_3,n_578_port_0,n_578_port_1, n_578_v);
  spice_node_2 n_n_572(eclk, ereset, n_572_port_3,n_572_port_0, n_572_v);
  spice_node_2 n_n_570(eclk, ereset, n_570_port_6,n_570_port_5, n_570_v);
  spice_node_3 n_n_571(eclk, ereset, n_571_port_2,n_571_port_3,n_571_port_1, n_571_v);
  spice_node_2 n_n_318(eclk, ereset, n_318_port_1,n_318_port_4, n_318_v);
  spice_node_2 n_n_319(eclk, ereset, n_319_port_2,n_319_port_4, n_319_v);
  spice_node_2 n_n_312(eclk, ereset, n_312_port_2,n_312_port_3, n_312_v);
  spice_node_2 n_n_310(eclk, ereset, n_310_port_3,n_310_port_0, n_310_v);
  spice_node_2 n_n_311(eclk, ereset, n_311_port_2,n_311_port_3, n_311_v);
  spice_node_2 n_n_317(eclk, ereset, n_317_port_2,n_317_port_0, n_317_v);
  spice_node_2 n_PD_n_0xx0xx0x(eclk, ereset, PD_n_0xx0xx0x_port_2,PD_n_0xx0xx0x_port_0, PD_n_0xx0xx0x_v);
  spice_node_2 n_C23(eclk, ereset, C23_port_7,C23_port_4, C23_v);
  spice_node_2 n_PD_0xx0xx0x(eclk, ereset, PD_0xx0xx0x_port_4,PD_0xx0xx0x_port_5, PD_0xx0xx0x_v);
  spice_node_2 n_op_T0_dex(eclk, ereset, op_T0_dex_port_9,op_T0_dex_port_11, op_T0_dex_v);
  spice_node_2 n_op_T__ora_and_eor_adc(eclk, ereset, op_T__ora_and_eor_adc_port_6,op_T__ora_and_eor_adc_port_4, op_T__ora_and_eor_adc_v);
  spice_node_2 n_dpc14_SRS(eclk, ereset, dpc14_SRS_port_2,dpc14_SRS_port_1, dpc14_SRS_v);
  spice_node_2 n_op_T2_ind_x(eclk, ereset, op_T2_ind_x_port_8,op_T2_ind_x_port_6, op_T2_ind_x_v);
  spice_node_2 n_op_T2_ind_y(eclk, ereset, op_T2_ind_y_port_8,op_T2_ind_y_port_6, op_T2_ind_y_v);
  spice_node_2 n_op_plp_pla(eclk, ereset, op_plp_pla_port_9,op_plp_pla_port_7, op_plp_pla_v);
  spice_node_2 n_op_T0_txs(eclk, ereset, op_T0_txs_port_10,op_T0_txs_port_12, op_T0_txs_v);
  spice_node_3 n_n_66(eclk, ereset, n_66_port_2,n_66_port_3,n_66_port_1, n_66_v);
  spice_node_2 n_n_62(eclk, ereset, n_62_port_2,n_62_port_1, n_62_v);
  spice_node_2 n_n_61(eclk, ereset, n_61_port_3,n_61_port_0, n_61_v);
  spice_node_2 n_n_149(eclk, ereset, n_149_port_3,n_149_port_0, n_149_v);
  spice_node_2 n_n_147(eclk, ereset, n_147_port_3,n_147_port_4, n_147_v);
  spice_node_5 n_n_146(eclk, ereset, n_146_port_2,n_146_port_3,n_146_port_0,n_146_port_1,n_146_port_4, n_146_v);
  spice_node_5 n_n_141(eclk, ereset, n_141_port_2,n_141_port_3,n_141_port_0,n_141_port_1,n_141_port_4, n_141_v);
  spice_node_2 n__op_set_C(eclk, ereset, _op_set_C_port_7,_op_set_C_port_10, _op_set_C_v);
  spice_node_2 n_op_T5_rti(eclk, ereset, op_T5_rti_port_10,op_T5_rti_port_13, op_T5_rti_v);
  spice_node_2 n_op_T5_ind_y(eclk, ereset, op_T5_ind_y_port_8,op_T5_ind_y_port_6, op_T5_ind_y_v);
  spice_node_2 n_op_T5_ind_x(eclk, ereset, op_T5_ind_x_port_9,op_T5_ind_x_port_7, op_T5_ind_x_v);
  spice_node_2 n_op_T3_jsr(eclk, ereset, op_T3_jsr_port_9,op_T3_jsr_port_10, op_T3_jsr_v);
  spice_node_2 n_op_T5_brk(eclk, ereset, op_T5_brk_port_10,op_T5_brk_port_12, op_T5_brk_v);
  spice_node_2 n_ADL_ABL(eclk, ereset, ADL_ABL_port_0,ADL_ABL_port_5, ADL_ABL_v);
  spice_node_2 n_n_1371(eclk, ereset, n_1371_port_6,n_1371_port_4, n_1371_v);
  spice_node_2 n_n_1376(eclk, ereset, n_1376_port_2,n_1376_port_1, n_1376_v);
  spice_node_2 n_n_1377(eclk, ereset, n_1377_port_2,n_1377_port_1, n_1377_v);
  spice_node_2 n_n_1374(eclk, ereset, n_1374_port_4,n_1374_port_5, n_1374_v);
  spice_node_2 n_n_1375(eclk, ereset, n_1375_port_2,n_1375_port_0, n_1375_v);
  spice_node_2 n_n_1379(eclk, ereset, n_1379_port_2,n_1379_port_1, n_1379_v);
  spice_node_4 n_n_1724(eclk, ereset, n_1724_port_2,n_1724_port_3,n_1724_port_0,n_1724_port_1, n_1724_v);
  spice_node_2 n_n_1194(eclk, ereset, n_1194_port_2,n_1194_port_3, n_1194_v);
  spice_node_2 n_n_1195(eclk, ereset, n_1195_port_2,n_1195_port_3, n_1195_v);
  spice_node_2 n_n_1192(eclk, ereset, n_1192_port_2,n_1192_port_3, n_1192_v);
  spice_node_2 n_n_1190(eclk, ereset, n_1190_port_2,n_1190_port_0, n_1190_v);
  spice_node_2 n_n_1191(eclk, ereset, n_1191_port_2,n_1191_port_0, n_1191_v);
  spice_node_2 n_n_708(eclk, ereset, n_708_port_2,n_708_port_1, n_708_v);
  spice_node_2 n_n_556(eclk, ereset, n_556_port_2,n_556_port_0, n_556_v);
  spice_node_2 n_n_550(eclk, ereset, n_550_port_3,n_550_port_5, n_550_v);
  spice_node_2 n_n_551(eclk, ereset, n_551_port_2,n_551_port_1, n_551_v);
  spice_node_2 n_n_553(eclk, ereset, n_553_port_3,n_553_port_4, n_553_v);
  spice_node_2 n_C45(eclk, ereset, C45_port_7,C45_port_4, C45_v);
  spice_node_2 n_x_op_T3_ind_y(eclk, ereset, x_op_T3_ind_y_port_6,x_op_T3_ind_y_port_7, x_op_T3_ind_y_v);
  spice_node_2 n_op_T__asl_rol_a(eclk, ereset, op_T__asl_rol_a_port_8,op_T__asl_rol_a_port_10, op_T__asl_rol_a_v);
  spice_node_2 n_n_882(eclk, ereset, n_882_port_3,n_882_port_5, n_882_v);
  spice_node_3 n_n_883(eclk, ereset, n_883_port_2,n_883_port_3,n_883_port_1, n_883_v);
  spice_node_3 n_n_880(eclk, ereset, n_880_port_2,n_880_port_3,n_880_port_0, n_880_v);
  spice_node_2 n_n_334(eclk, ereset, n_334_port_6,n_334_port_5, n_334_v);
  spice_node_2 n_n_335(eclk, ereset, n_335_port_8,n_335_port_10, n_335_v);
  spice_node_4 n_n_336(eclk, ereset, n_336_port_3,n_336_port_1,n_336_port_6,n_336_port_7, n_336_v);
  spice_node_2 n_n_885(eclk, ereset, n_885_port_2,n_885_port_0, n_885_v);
  spice_node_2 n_n_888(eclk, ereset, n_888_port_2,n_888_port_0, n_888_v);
  spice_node_2 n_n_889(eclk, ereset, n_889_port_2,n_889_port_1, n_889_v);
  spice_node_2 n__AxB_4__C34(eclk, ereset, _AxB_4__C34_port_3,_AxB_4__C34_port_4, _AxB_4__C34_v);
  spice_node_2 n_dpc28_0ADH0(eclk, ereset, dpc28_0ADH0_port_2,dpc28_0ADH0_port_0, dpc28_0ADH0_v);
  spice_node_2 n_fetch(eclk, ereset, fetch_port_11,fetch_port_12, fetch_v);
  spice_node_2 n_op_ANDS(eclk, ereset, op_ANDS_port_6,op_ANDS_port_5, op_ANDS_v);
  spice_node_2 n_n_46(eclk, ereset, n_46_port_3,n_46_port_4, n_46_v);
  spice_node_2 n_n_43(eclk, ereset, n_43_port_11,n_43_port_13, n_43_v);
  spice_node_2 n_n_42(eclk, ereset, n_42_port_0,n_42_port_4, n_42_v);
  spice_node_2 n_op_T__cpx_cpy_abs(eclk, ereset, op_T__cpx_cpy_abs_port_8,op_T__cpx_cpy_abs_port_10, op_T__cpx_cpy_abs_v);
  spice_node_2 n_n_1153(eclk, ereset, n_1153_port_3,n_1153_port_0, n_1153_v);
  spice_node_1 n_res(eclk, ereset, res_port_2, res_v);
  spice_node_7 n_adl7(eclk, ereset, adl7_port_2,adl7_port_3,adl7_port_0,adl7_port_6,adl7_port_7,adl7_port_4,adl7_port_5, adl7_v);
  spice_node_7 n_adl6(eclk, ereset, adl6_port_2,adl6_port_3,adl6_port_1,adl6_port_6,adl6_port_7,adl6_port_4,adl6_port_5, adl6_v);
  spice_node_7 n_adl5(eclk, ereset, adl5_port_2,adl5_port_3,adl5_port_0,adl5_port_1,adl5_port_7,adl5_port_4,adl5_port_5, adl5_v);
  spice_node_7 n_adl4(eclk, ereset, adl4_port_3,adl4_port_0,adl4_port_1,adl4_port_6,adl4_port_7,adl4_port_4,adl4_port_5, adl4_v);
  spice_node_7 n_adl3(eclk, ereset, adl3_port_2,adl3_port_3,adl3_port_0,adl3_port_1,adl3_port_6,adl3_port_7,adl3_port_4, adl3_v);
  spice_node_8 n_adl2(eclk, ereset, adl2_port_8,adl2_port_2,adl2_port_3,adl2_port_0,adl2_port_1,adl2_port_6,adl2_port_4,adl2_port_5, adl2_v);
  spice_node_8 n_adl1(eclk, ereset, adl1_port_8,adl1_port_2,adl1_port_3,adl1_port_0,adl1_port_1,adl1_port_7,adl1_port_4,adl1_port_5, adl1_v);
  spice_node_8 n_adl0(eclk, ereset, adl0_port_8,adl0_port_3,adl0_port_0,adl0_port_1,adl0_port_6,adl0_port_7,adl0_port_4,adl0_port_5, adl0_v);
  spice_node_4 n_n_1014(eclk, ereset, n_1014_port_2,n_1014_port_3,n_1014_port_0,n_1014_port_1, n_1014_v);
  spice_node_2 n_n_0_ADL1(eclk, ereset, n_0_ADL1_port_2,n_0_ADL1_port_0, n_0_ADL1_v);
  spice_node_2 n_n_0_ADL0(eclk, ereset, n_0_ADL0_port_3,n_0_ADL0_port_0, n_0_ADL0_v);
  spice_node_2 n_n_0_ADL2(eclk, ereset, n_0_ADL2_port_2,n_0_ADL2_port_0, n_0_ADL2_v);
  spice_node_2 n_op_T3_abs_idx(eclk, ereset, op_T3_abs_idx_port_6,op_T3_abs_idx_port_4, op_T3_abs_idx_v);
  spice_node_2 n_op_jsr(eclk, ereset, op_jsr_port_8,op_jsr_port_9, op_jsr_v);
  spice_node_2 n_dpc40_ADLPCL(eclk, ereset, dpc40_ADLPCL_port_0,dpc40_ADLPCL_port_12, dpc40_ADLPCL_v);
  spice_node_2 n_n_593(eclk, ereset, n_593_port_2,n_593_port_1, n_593_v);
  spice_node_5 n_n_929(eclk, ereset, n_929_port_2,n_929_port_3,n_929_port_0,n_929_port_1,n_929_port_4, n_929_v);
  spice_node_2 n_n_1255(eclk, ereset, n_1255_port_2,n_1255_port_1, n_1255_v);
  spice_node_2 n_n_1358(eclk, ereset, n_1358_port_6,n_1358_port_5, n_1358_v);
  spice_node_2 n_n_1427(eclk, ereset, n_1427_port_3,n_1427_port_4, n_1427_v);
  spice_node_4 n_n_1424(eclk, ereset, n_1424_port_2,n_1424_port_3,n_1424_port_0,n_1424_port_1, n_1424_v);
  spice_node_2 n_n_1357(eclk, ereset, n_1357_port_0,n_1357_port_5, n_1357_v);
  spice_node_5 n_notaluoutmux0(eclk, ereset, notaluoutmux0_port_2,notaluoutmux0_port_3,notaluoutmux0_port_0,notaluoutmux0_port_1,notaluoutmux0_port_5, notaluoutmux0_v);
  spice_node_5 n_notaluoutmux1(eclk, ereset, notaluoutmux1_port_2,notaluoutmux1_port_0,notaluoutmux1_port_1,notaluoutmux1_port_4,notaluoutmux1_port_5, notaluoutmux1_v);
  spice_node_2 n_n_533(eclk, ereset, n_533_port_2,n_533_port_1, n_533_v);
  spice_node_2 n_n_531(eclk, ereset, n_531_port_3,n_531_port_0, n_531_v);
  spice_node_2 n_n_538(eclk, ereset, n_538_port_2,n_538_port_1, n_538_v);
  spice_node_2 n_C67(eclk, ereset, C67_port_6,C67_port_11, C67_v);
  spice_node_2 n_C1x5Reset(eclk, ereset, C1x5Reset_port_2,C1x5Reset_port_5, C1x5Reset_v);
  spice_node_2 n_op_T__adc_sbc(eclk, ereset, op_T__adc_sbc_port_7,op_T__adc_sbc_port_5, op_T__adc_sbc_v);
  spice_node_2 n_op_T0_cmp(eclk, ereset, op_T0_cmp_port_6,op_T0_cmp_port_7, op_T0_cmp_v);
  spice_node_2 n_n_1218(eclk, ereset, n_1218_port_2,n_1218_port_1, n_1218_v);
  spice_node_2 n_dpc30_ADHPCH(eclk, ereset, dpc30_ADHPCH_port_10,dpc30_ADHPCH_port_12, dpc30_ADHPCH_v);
  spice_node_2 n_dpc43_DL_DB(eclk, ereset, dpc43_DL_DB_port_9,dpc43_DL_DB_port_0, dpc43_DL_DB_v);
  spice_node_2 n_n_23(eclk, ereset, n_23_port_4,n_23_port_5, n_23_v);
  spice_node_2 n_n_21(eclk, ereset, n_21_port_4,n_21_port_5, n_21_v);
  spice_node_2 n_n_20(eclk, ereset, n_20_port_3,n_20_port_5, n_20_v);
  spice_node_5 n_n_27(eclk, ereset, n_27_port_2,n_27_port_3,n_27_port_0,n_27_port_1,n_27_port_4, n_27_v);
  spice_node_3 n_aluanorb0(eclk, ereset, aluanorb0_port_1,aluanorb0_port_6,aluanorb0_port_7, aluanorb0_v);
  spice_node_2 n_n_25(eclk, ereset, n_25_port_3,n_25_port_4, n_25_v);
  spice_node_2 n_n_29(eclk, ereset, n_29_port_2,n_29_port_3, n_29_v);
  spice_node_4 n_n_1694(eclk, ereset, n_1694_port_2,n_1694_port_3,n_1694_port_0,n_1694_port_1, n_1694_v);
  spice_node_2 n_a1(eclk, ereset, a1_port_0,a1_port_1, a1_v);
  spice_node_2 n_a0(eclk, ereset, a0_port_0,a0_port_1, a0_v);
  spice_node_2 n_a2(eclk, ereset, a2_port_2,a2_port_1, a2_v);
  spice_node_2 n_a5(eclk, ereset, a5_port_2,a5_port_0, a5_v);
  spice_node_2 n_a4(eclk, ereset, a4_port_2,a4_port_0, a4_v);
  spice_node_2 n_a7(eclk, ereset, a7_port_2,a7_port_1, a7_v);
  spice_node_2 n_n_275(eclk, ereset, n_275_port_3,n_275_port_4, n_275_v);
  spice_node_5 n_n_277(eclk, ereset, n_277_port_2,n_277_port_3,n_277_port_1,n_277_port_4,n_277_port_5, n_277_v);
  spice_node_2 n_n_270(eclk, ereset, n_270_port_2,n_270_port_6, n_270_v);
  spice_node_2 n_n_272(eclk, ereset, n_272_port_8,n_272_port_9, n_272_v);
  spice_node_2 n_n_278(eclk, ereset, n_278_port_2,n_278_port_0, n_278_v);
  spice_node_2 n_n_1486(eclk, ereset, n_1486_port_3,n_1486_port_5, n_1486_v);
  spice_node_2 n_n_638(eclk, ereset, n_638_port_2,n_638_port_0, n_638_v);
  spice_node_2 n_n_1408(eclk, ereset, n_1408_port_2,n_1408_port_3, n_1408_v);
  spice_node_2 n_n_188(eclk, ereset, n_188_port_4,n_188_port_5, n_188_v);
  spice_node_2 n_n_1400(eclk, ereset, n_1400_port_2,n_1400_port_0, n_1400_v);
  spice_node_2 n_n_1402(eclk, ereset, n_1402_port_2,n_1402_port_3, n_1402_v);
  spice_node_2 n_op_T0_ora(eclk, ereset, op_T0_ora_port_6,op_T0_ora_port_7, op_T0_ora_v);
  spice_node_4 n_n_518(eclk, ereset, n_518_port_2,n_518_port_3,n_518_port_0,n_518_port_1, n_518_v);
  spice_node_2 n_n_519(eclk, ereset, n_519_port_2,n_519_port_4, n_519_v);
  spice_node_2 n_n_510(eclk, ereset, n_510_port_6,n_510_port_4, n_510_v);
  spice_node_2 n_n_513(eclk, ereset, n_513_port_4,n_513_port_5, n_513_v);
  spice_node_2 n_n_515(eclk, ereset, n_515_port_3,n_515_port_5, n_515_v);
  spice_node_2 n_n_1463(eclk, ereset, n_1463_port_4,n_1463_port_5, n_1463_v);
  spice_node_2 n_n_453(eclk, ereset, n_453_port_3,n_453_port_1, n_453_v);
  spice_node_2 n_n_1467(eclk, ereset, n_1467_port_0,n_1467_port_1, n_1467_v);
  spice_node_2 n_n_980(eclk, ereset, n_980_port_2,n_980_port_0, n_980_v);
  spice_node_2 n_n_1464(eclk, ereset, n_1464_port_8,n_1464_port_7, n_1464_v);
  spice_node_2 n_alucout(eclk, ereset, alucout_port_3,alucout_port_0, alucout_v);
  spice_node_2 n_op_brk_rti(eclk, ereset, op_brk_rti_port_8,op_brk_rti_port_7, op_brk_rti_v);
  spice_node_2 n_DBZ(eclk, ereset, DBZ_port_9,DBZ_port_10, DBZ_v);
  spice_node_2 n_n_1600(eclk, ereset, n_1600_port_2,n_1600_port_0, n_1600_v);
  spice_node_2 n_n_1093(eclk, ereset, n_1093_port_2,n_1093_port_1, n_1093_v);
  spice_node_2 n_n_1091(eclk, ereset, n_1091_port_3,n_1091_port_6, n_1091_v);
  spice_node_2 n_n_1090(eclk, ereset, n_1090_port_3,n_1090_port_4, n_1090_v);
  spice_node_2 n_n_1097(eclk, ereset, n_1097_port_3,n_1097_port_4, n_1097_v);
  spice_node_4 n_n_1095(eclk, ereset, n_1095_port_2,n_1095_port_3,n_1095_port_0,n_1095_port_1, n_1095_v);
  spice_node_3 n_n_1094(eclk, ereset, n_1094_port_2,n_1094_port_3,n_1094_port_1, n_1094_v);
  spice_node_2 n_n_1099(eclk, ereset, n_1099_port_2,n_1099_port_3, n_1099_v);
  spice_node_2 n_n_1677(eclk, ereset, n_1677_port_2,n_1677_port_3, n_1677_v);
  spice_node_2 n_n_1676(eclk, ereset, n_1676_port_2,n_1676_port_3, n_1676_v);
  spice_node_2 n_n_1675(eclk, ereset, n_1675_port_3,n_1675_port_0, n_1675_v);
  spice_node_6 n_adh3(eclk, ereset, adh3_port_2,adh3_port_3,adh3_port_0,adh3_port_6,adh3_port_4,adh3_port_5, adh3_v);
  spice_node_6 n_adh2(eclk, ereset, adh2_port_3,adh2_port_0,adh2_port_1,adh2_port_6,adh2_port_4,adh2_port_5, adh2_v);
  spice_node_6 n_adh1(eclk, ereset, adh1_port_2,adh1_port_0,adh1_port_1,adh1_port_6,adh1_port_4,adh1_port_5, adh1_v);
  spice_node_6 n_adh0(eclk, ereset, adh0_port_2,adh0_port_3,adh0_port_0,adh0_port_1,adh0_port_6,adh0_port_4, adh0_v);
  spice_node_6 n_adh7(eclk, ereset, adh7_port_2,adh7_port_3,adh7_port_0,adh7_port_1,adh7_port_4,adh7_port_5, adh7_v);
  spice_node_6 n_adh6(eclk, ereset, adh6_port_3,adh6_port_0,adh6_port_1,adh6_port_6,adh6_port_4,adh6_port_5, adh6_v);
  spice_node_6 n_adh5(eclk, ereset, adh5_port_2,adh5_port_3,adh5_port_0,adh5_port_1,adh5_port_4,adh5_port_5, adh5_v);
  spice_node_6 n_adh4(eclk, ereset, adh4_port_2,adh4_port_0,adh4_port_1,adh4_port_6,adh4_port_4,adh4_port_5, adh4_v);
  spice_node_2 n_op_T5_rts(eclk, ereset, op_T5_rts_port_12,op_T5_rts_port_14, op_T5_rts_v);
  spice_node_2 n_n_253(eclk, ereset, n_253_port_2,n_253_port_3, n_253_v);
  spice_node_2 n_n_251(eclk, ereset, n_251_port_4,n_251_port_5, n_251_v);
  spice_node_2 n_n_709(eclk, ereset, n_709_port_2,n_709_port_0, n_709_v);
  spice_node_2 n_n_256(eclk, ereset, n_256_port_8,n_256_port_9, n_256_v);
  spice_node_2 n_n_255(eclk, ereset, n_255_port_2,n_255_port_1, n_255_v);
  spice_node_3 n_n_254(eclk, ereset, n_254_port_2,n_254_port_3,n_254_port_1, n_254_v);
  spice_node_2 n_n_700(eclk, ereset, n_700_port_3,n_700_port_1, n_700_v);
  spice_node_2 n_n_1462(eclk, ereset, n_1462_port_2,n_1462_port_0, n_1462_v);
  spice_node_3 n_n_1469(eclk, ereset, n_1469_port_2,n_1469_port_0,n_1469_port_1, n_1469_v);
  spice_node_2 n_n_714(eclk, ereset, n_714_port_2,n_714_port_1, n_714_v);
  spice_node_2 n_n_1286(eclk, ereset, n_1286_port_3,n_1286_port_5, n_1286_v);
  spice_node_2 n_n_1281(eclk, ereset, n_1281_port_2,n_1281_port_0, n_1281_v);
  spice_node_2 n_n_1289(eclk, ereset, n_1289_port_2,n_1289_port_1, n_1289_v);
  spice_node_2 n_A_B7(eclk, ereset, A_B7_port_2,A_B7_port_1, A_B7_v);
  spice_node_2 n_A_B5(eclk, ereset, A_B5_port_2,A_B5_port_1, A_B5_v);
  spice_node_2 n_A_B3(eclk, ereset, A_B3_port_2,A_B3_port_1, A_B3_v);
  spice_node_2 n_A_B1(eclk, ereset, A_B1_port_2,A_B1_port_0, A_B1_v);
  spice_node_2 n_n_392(eclk, ereset, n_392_port_2,n_392_port_3, n_392_v);
  spice_node_2 n_n_390(eclk, ereset, n_390_port_2,n_390_port_0, n_390_v);
  spice_node_2 n_n_396(eclk, ereset, n_396_port_2,n_396_port_1, n_396_v);
  spice_node_2 n_n_397(eclk, ereset, n_397_port_2,n_397_port_0, n_397_v);
  spice_node_2 n_n_1497(eclk, ereset, n_1497_port_2,n_1497_port_1, n_1497_v);
  spice_node_2 n_n_936(eclk, ereset, n_936_port_4,n_936_port_5, n_936_v);
  spice_node_2 n_n_937(eclk, ereset, n_937_port_0,n_937_port_4, n_937_v);
  spice_node_3 n_n_935(eclk, ereset, n_935_port_2,n_935_port_3,n_935_port_1, n_935_v);
  spice_node_2 n_n_933(eclk, ereset, n_933_port_2,n_933_port_4, n_933_v);
  spice_node_2 n_n_931(eclk, ereset, n_931_port_2,n_931_port_1, n_931_v);
  spice_node_2 n_op_T2_php_pha(eclk, ereset, op_T2_php_pha_port_9,op_T2_php_pha_port_12, op_T2_php_pha_v);
  spice_node_2 n_ONEBYTE(eclk, ereset, ONEBYTE_port_2,ONEBYTE_port_1, ONEBYTE_v);
  spice_node_2 n_NMIP(eclk, ereset, NMIP_port_7,NMIP_port_4, NMIP_v);
  spice_node_2 n_n_1075(eclk, ereset, n_1075_port_2,n_1075_port_1, n_1075_v);
  spice_node_2 n_n_1076(eclk, ereset, n_1076_port_0,n_1076_port_4, n_1076_v);
  spice_node_5 n_n_1071(eclk, ereset, n_1071_port_2,n_1071_port_3,n_1071_port_0,n_1071_port_4,n_1071_port_5, n_1071_v);
  spice_node_2 n_n_1070(eclk, ereset, n_1070_port_3,n_1070_port_4, n_1070_v);
  spice_node_2 n_n_1073(eclk, ereset, n_1073_port_2,n_1073_port_3, n_1073_v);
  spice_node_2 n_n_1072(eclk, ereset, n_1072_port_2,n_1072_port_4, n_1072_v);
  spice_node_2 n_abl2(eclk, ereset, abl2_port_3,abl2_port_4, abl2_v);
  spice_node_2 n_abl5(eclk, ereset, abl5_port_0,abl5_port_4, abl5_v);
  spice_node_2 n_abl6(eclk, ereset, abl6_port_0,abl6_port_4, abl6_v);
  spice_node_2 n_n_1619(eclk, ereset, n_1619_port_3,n_1619_port_4, n_1619_v);
  spice_node_2 n_notaluvout(eclk, ereset, notaluvout_port_3,notaluvout_port_5, notaluvout_v);
  spice_node_2 n_n_1140(eclk, ereset, n_1140_port_2,n_1140_port_1, n_1140_v);
  spice_node_2 n_n_1614(eclk, ereset, n_1614_port_4,n_1614_port_5, n_1614_v);
  spice_node_2 n_n_1145(eclk, ereset, n_1145_port_3,n_1145_port_4, n_1145_v);
  spice_node_4 n_n_1147(eclk, ereset, n_1147_port_2,n_1147_port_3,n_1147_port_0,n_1147_port_1, n_1147_v);
  spice_node_2 n_dpc34_PCLC(eclk, ereset, dpc34_PCLC_port_12,dpc34_PCLC_port_14, dpc34_PCLC_v);
  spice_node_3 n_aluanorb1(eclk, ereset, aluanorb1_port_7,aluanorb1_port_4,aluanorb1_port_5, aluanorb1_v);
  spice_node_2 n_H1x1(eclk, ereset, H1x1_port_8,H1x1_port_4, H1x1_v);
  spice_node_2 n_n_238(eclk, ereset, n_238_port_2,n_238_port_1, n_238_v);
  spice_node_2 n_n_728(eclk, ereset, n_728_port_2,n_728_port_0, n_728_v);
  spice_node_5 n_n_723(eclk, ereset, n_723_port_2,n_723_port_3,n_723_port_0,n_723_port_1,n_723_port_4, n_723_v);
  spice_node_5 n_n_722(eclk, ereset, n_722_port_2,n_722_port_0,n_722_port_1,n_722_port_4,n_722_port_5, n_722_v);
  spice_node_5 n_n_721(eclk, ereset, n_721_port_2,n_721_port_3,n_721_port_0,n_721_port_1,n_721_port_4, n_721_v);
  spice_node_2 n_n_720(eclk, ereset, n_720_port_3,n_720_port_4, n_720_v);
  spice_node_2 n_n_726(eclk, ereset, n_726_port_6,n_726_port_5, n_726_v);
  spice_node_2 n_dpc1_SBY(eclk, ereset, dpc1_SBY_port_3,dpc1_SBY_port_12, dpc1_SBY_v);
  spice_node_2 n_op_T2_abs(eclk, ereset, op_T2_abs_port_7,op_T2_abs_port_5, op_T2_abs_v);
  spice_node_2 n_op_T0_plp(eclk, ereset, op_T0_plp_port_9,op_T0_plp_port_10, op_T0_plp_v);
  spice_node_2 n_op_T0_pla(eclk, ereset, op_T0_pla_port_9,op_T0_pla_port_11, op_T0_pla_v);
  spice_node_2 n_op_T2_jmp_abs(eclk, ereset, op_T2_jmp_abs_port_9,op_T2_jmp_abs_port_11, op_T2_jmp_abs_v);
  spice_node_2 n__C34(eclk, ereset, _C34_port_9,_C34_port_5, _C34_v);
  spice_node_2 n_DA_C01(eclk, ereset, DA_C01_port_8,DA_C01_port_4, DA_C01_v);
  spice_node_2 n_n_1448(eclk, ereset, n_1448_port_2,n_1448_port_0, n_1448_v);
  spice_node_2 n_n_1449(eclk, ereset, n_1449_port_2,n_1449_port_1, n_1449_v);
  spice_node_2 n_cclk(eclk, ereset, cclk_port_236,cclk_port_28, cclk_v);
  spice_node_2 n_n_1446(eclk, ereset, n_1446_port_3,n_1446_port_4, n_1446_v);
  spice_node_2 n_n_1440(eclk, ereset, n_1440_port_2,n_1440_port_1, n_1440_v);
  spice_node_2 n_n_1441(eclk, ereset, n_1441_port_2,n_1441_port_1, n_1441_v);
  spice_node_2 n_notRnWprepad(eclk, ereset, notRnWprepad_port_6,notRnWprepad_port_7, notRnWprepad_v);
  spice_node_2 n_n_1511(eclk, ereset, n_1511_port_2,n_1511_port_1, n_1511_v);
  spice_node_2 n_n_918(eclk, ereset, n_918_port_2,n_918_port_1, n_918_v);
  spice_node_2 n_n_919(eclk, ereset, n_919_port_6,n_919_port_4, n_919_v);
  spice_node_2 n_n_916(eclk, ereset, n_916_port_7,n_916_port_4, n_916_v);
  spice_node_2 n_RnWstretched(eclk, ereset, RnWstretched_port_23,RnWstretched_port_22, RnWstretched_v);
  spice_node_2 n_n_913(eclk, ereset, n_913_port_2,n_913_port_0, n_913_v);
  spice_node_2 n_op_T0_tay_ldy_not_idx(eclk, ereset, op_T0_tay_ldy_not_idx_port_8,op_T0_tay_ldy_not_idx_port_7, op_T0_tay_ldy_not_idx_v);
  spice_node_2 n_op_T0(eclk, ereset, op_T0_port_2,op_T0_port_1, op_T0_v);
  spice_node_2 n_op_T3(eclk, ereset, op_T3_port_2,op_T3_port_0, op_T3_v);
  spice_node_2 n_op_T2(eclk, ereset, op_T2_port_2,op_T2_port_0, op_T2_v);
  spice_node_2 n_op_T4(eclk, ereset, op_T4_port_2,op_T4_port_1, op_T4_v);
  spice_node_2 n_n_1224(eclk, ereset, n_1224_port_2,n_1224_port_0, n_1224_v);
  spice_node_2 n_op_T3_stack_bit_jmp(eclk, ereset, op_T3_stack_bit_jmp_port_7,op_T3_stack_bit_jmp_port_5, op_T3_stack_bit_jmp_v);
  spice_node_2 n_op_T5_jsr(eclk, ereset, op_T5_jsr_port_9,op_T5_jsr_port_10, op_T5_jsr_v);
  spice_node_2 n_op_T2_stack_access(eclk, ereset, op_T2_stack_access_port_6,op_T2_stack_access_port_7, op_T2_stack_access_v);
  spice_node_2 n_n_1056(eclk, ereset, n_1056_port_2,n_1056_port_0, n_1056_v);
  spice_node_2 n_n_1055(eclk, ereset, n_1055_port_3,n_1055_port_5, n_1055_v);
  spice_node_2 n_n_1054(eclk, ereset, n_1054_port_2,n_1054_port_0, n_1054_v);
  spice_node_2 n_op_T4_mem_abs_idx(eclk, ereset, op_T4_mem_abs_idx_port_6,op_T4_mem_abs_idx_port_4, op_T4_mem_abs_idx_v);
  spice_node_1 n_n_1059(eclk, ereset, n_1059_port_0, n_1059_v);
  spice_node_2 n_n_1588(eclk, ereset, n_1588_port_2,n_1588_port_1, n_1588_v);
  spice_node_2 n_n_1580(eclk, ereset, n_1580_port_3,n_1580_port_0, n_1580_v);
  spice_node_2 n_n_1633(eclk, ereset, n_1633_port_2,n_1633_port_0, n_1633_v);
  spice_node_2 n_n_1639(eclk, ereset, n_1639_port_2,n_1639_port_0, n_1639_v);
  spice_node_2 n_n_1638(eclk, ereset, n_1638_port_2,n_1638_port_1, n_1638_v);
  spice_node_2 n_C34(eclk, ereset, C34_port_2,C34_port_5, C34_v);
  spice_node_2 n__DA_ADD2(eclk, ereset, _DA_ADD2_port_2,_DA_ADD2_port_3, _DA_ADD2_v);
  spice_node_2 n__DA_ADD1(eclk, ereset, _DA_ADD1_port_0,_DA_ADD1_port_5, _DA_ADD1_v);
  spice_node_5 n_n_740(eclk, ereset, n_740_port_2,n_740_port_3,n_740_port_0,n_740_port_1,n_740_port_4, n_740_v);
  spice_node_2 n_n_743(eclk, ereset, n_743_port_7,n_743_port_5, n_743_v);
  spice_node_2 n_n_213(eclk, ereset, n_213_port_2,n_213_port_0, n_213_v);
  spice_node_3 n_n_212(eclk, ereset, n_212_port_2,n_212_port_3,n_212_port_1, n_212_v);
  spice_node_2 n_n_747(eclk, ereset, n_747_port_3,n_747_port_0, n_747_v);
  spice_node_3 n_n_210(eclk, ereset, n_210_port_3,n_210_port_0,n_210_port_1, n_210_v);
  spice_node_2 n_n_748(eclk, ereset, n_748_port_3,n_748_port_0, n_748_v);
  spice_node_2 n_n_218(eclk, ereset, n_218_port_2,n_218_port_0, n_218_v);
  spice_node_2 n_notRdy0(eclk, ereset, notRdy0_port_3,notRdy0_port_4, notRdy0_v);
  spice_node_2 n_notalucout(eclk, ereset, notalucout_port_4,notalucout_port_5, notalucout_v);
  spice_node_2 n_dpc36_IPC(eclk, ereset, dpc36_IPC_port_5,dpc36_IPC_port_10, dpc36_IPC_v);
  spice_node_2 n_op_T0_cpx_cpy_inx_iny(eclk, ereset, op_T0_cpx_cpy_inx_iny_port_6,op_T0_cpx_cpy_inx_iny_port_7, op_T0_cpx_cpy_inx_iny_v);
  spice_node_3 n_n_624(eclk, ereset, n_624_port_2,n_624_port_0,n_624_port_1, n_624_v);
  spice_node_2 n_op_T2_zp_zp_idx(eclk, ereset, op_T2_zp_zp_idx_port_4,op_T2_zp_zp_idx_port_5, op_T2_zp_zp_idx_v);
  spice_node_2 n__C12(eclk, ereset, _C12_port_7,_C12_port_4, _C12_v);
  spice_node_2 n_clk2out(eclk, ereset, clk2out_port_0,clk2out_port_1, clk2out_v);
  spice_node_2 n_n_689(eclk, ereset, n_689_port_2,n_689_port_0, n_689_v);
  spice_node_4 n_n_681(eclk, ereset, n_681_port_8,n_681_port_3,n_681_port_1,n_681_port_6, n_681_v);
  spice_node_2 n_n_1471(eclk, ereset, n_1471_port_2,n_1471_port_1, n_1471_v);
  spice_node_2 n_n_979(eclk, ereset, n_979_port_2,n_979_port_1, n_979_v);
  spice_node_2 n_n_973(eclk, ereset, n_973_port_2,n_973_port_1, n_973_v);
  spice_node_5 n_n_976(eclk, ereset, n_976_port_2,n_976_port_3,n_976_port_0,n_976_port_1,n_976_port_4, n_976_v);
  spice_node_2 n_n_975(eclk, ereset, n_975_port_3,n_975_port_6, n_975_v);
  spice_node_2 n_op_T__bit(eclk, ereset, op_T__bit_port_9,op_T__bit_port_10, op_T__bit_v);
  spice_node_2 n_op_T0_iny_dey(eclk, ereset, op_T0_iny_dey_port_8,op_T0_iny_dey_port_9, op_T0_iny_dey_v);
  spice_node_2 n_n_1270(eclk, ereset, n_1270_port_4,n_1270_port_5, n_1270_v);
  spice_node_2 n_op_T__cmp(eclk, ereset, op_T__cmp_port_8,op_T__cmp_port_6, op_T__cmp_v);
  spice_node_5 n_n_1618(eclk, ereset, n_1618_port_2,n_1618_port_3,n_1618_port_0,n_1618_port_1,n_1618_port_4, n_1618_v);
  spice_node_2 n_op_T0_jsr(eclk, ereset, op_T0_jsr_port_10,op_T0_jsr_port_12, op_T0_jsr_v);
  spice_node_2 n_n_1610(eclk, ereset, n_1610_port_3,n_1610_port_5, n_1610_v);
  spice_node_2 n_op_T2_abs_access(eclk, ereset, op_T2_abs_access_port_9,op_T2_abs_access_port_6, op_T2_abs_access_v);
  spice_node_2 n_n_1613(eclk, ereset, n_1613_port_4,n_1613_port_5, n_1613_v);
  spice_node_2 n_n_1033(eclk, ereset, n_1033_port_2,n_1033_port_0, n_1033_v);
  spice_node_2 n_n_1034(eclk, ereset, n_1034_port_3,n_1034_port_0, n_1034_v);
  spice_node_2 n_n_1037(eclk, ereset, n_1037_port_3,n_1037_port_5, n_1037_v);
  spice_node_3 n_alub3(eclk, ereset, alub3_port_2,alub3_port_3,alub3_port_4, alub3_v);
  spice_node_2 n_n_1038(eclk, ereset, n_1038_port_2,n_1038_port_1, n_1038_v);
  spice_node_3 n_alub1(eclk, ereset, alub1_port_0,alub1_port_1,alub1_port_4, alub1_v);
  spice_node_3 n_alub0(eclk, ereset, alub0_port_2,alub0_port_3,alub0_port_4, alub0_v);
  spice_node_3 n_alub7(eclk, ereset, alub7_port_3,alub7_port_0,alub7_port_4, alub7_v);
  spice_node_3 n_alub6(eclk, ereset, alub6_port_2,alub6_port_3,alub6_port_4, alub6_v);
  spice_node_3 n_alub5(eclk, ereset, alub5_port_2,alub5_port_3,alub5_port_4, alub5_v);
  spice_node_3 n_alub4(eclk, ereset, alub4_port_3,alub4_port_0,alub4_port_4, alub4_v);
  spice_node_2 n_x_op_T4_rti(eclk, ereset, x_op_T4_rti_port_9,x_op_T4_rti_port_10, x_op_T4_rti_v);
  spice_node_2 n_dpc42_DL_ADH(eclk, ereset, dpc42_DL_ADH_port_8,dpc42_DL_ADH_port_9, dpc42_DL_ADH_v);
  spice_node_2 n_n_769(eclk, ereset, n_769_port_6,n_769_port_4, n_769_v);
  spice_node_4 n_n_767(eclk, ereset, n_767_port_2,n_767_port_3,n_767_port_0,n_767_port_1, n_767_v);
  spice_node_2 n_n_763(eclk, ereset, n_763_port_2,n_763_port_1, n_763_v);
  spice_node_2 n_n_762(eclk, ereset, n_762_port_3,n_762_port_4, n_762_v);
  spice_node_2 n_n_761(eclk, ereset, n_761_port_4,n_761_port_5, n_761_v);
  spice_node_2 n_op_T3_abs_idx_ind(eclk, ereset, op_T3_abs_idx_ind_port_6,op_T3_abs_idx_ind_port_4, op_T3_abs_idx_ind_v);
  spice_node_2 n_op_T2_jsr(eclk, ereset, op_T2_jsr_port_11,op_T2_jsr_port_13, op_T2_jsr_v);
  spice_node_2 n_DA_C45(eclk, ereset, DA_C45_port_3,DA_C45_port_1, DA_C45_v);
  spice_node_2 n_n_231(eclk, ereset, n_231_port_2,n_231_port_1, n_231_v);
  spice_node_2 n__C78(eclk, ereset, _C78_port_3,_C78_port_5, _C78_v);
  spice_node_2 n_n_233(eclk, ereset, n_233_port_2,n_233_port_4, n_233_v);
  spice_node_2 n_n_232(eclk, ereset, n_232_port_0,n_232_port_4, n_232_v);
  spice_node_2 n_n_236(eclk, ereset, n_236_port_3,n_236_port_7, n_236_v);
  spice_node_2 n_n_951(eclk, ereset, n_951_port_3,n_951_port_0, n_951_v);
  spice_node_2 n_n_952(eclk, ereset, n_952_port_3,n_952_port_0, n_952_v);
  spice_node_3 n_n_953(eclk, ereset, n_953_port_2,n_953_port_0,n_953_port_1, n_953_v);
  spice_node_2 n_n_958(eclk, ereset, n_958_port_3,n_958_port_0, n_958_v);
  spice_node_2 n_n_959(eclk, ereset, n_959_port_4,n_959_port_5, n_959_v);
  spice_node_3 n_n_409(eclk, ereset, n_409_port_3,n_409_port_0,n_409_port_5, n_409_v);
  spice_node_2 n_op_T0_eor(eclk, ereset, op_T0_eor_port_6,op_T0_eor_port_7, op_T0_eor_v);
  spice_node_2 n_pd1_clearIR(eclk, ereset, pd1_clearIR_port_6,pd1_clearIR_port_4, pd1_clearIR_v);
  spice_node_2 n_abl3(eclk, ereset, abl3_port_3,abl3_port_4, abl3_v);
  spice_node_2 n_op_T0_jmp(eclk, ereset, op_T0_jmp_port_8,op_T0_jmp_port_9, op_T0_jmp_v);
  spice_node_2 n_n_1018(eclk, ereset, n_1018_port_2,n_1018_port_0, n_1018_v);
  spice_node_2 n_n_1549(eclk, ereset, n_1549_port_2,n_1549_port_1, n_1549_v);
  spice_node_3 n_n_1548(eclk, ereset, n_1548_port_2,n_1548_port_3,n_1548_port_1, n_1548_v);
  spice_node_3 n_n_1016(eclk, ereset, n_1016_port_2,n_1016_port_3,n_1016_port_1, n_1016_v);
  spice_node_3 n_p4(eclk, ereset, p4_port_2,p4_port_0,p4_port_1, p4_v);
  spice_node_2 n___AxB1__C01(eclk, ereset, __AxB1__C01_port_3,__AxB1__C01_port_4, __AxB1__C01_v);
  spice_node_2 n_op_T2_idx_x_xy(eclk, ereset, op_T2_idx_x_xy_port_6,op_T2_idx_x_xy_port_5, op_T2_idx_x_xy_v);
  spice_node_2 n_op_clv(eclk, ereset, op_clv_port_8,op_clv_port_9, op_clv_v);
  spice_node_2 n_op_T0_and(eclk, ereset, op_T0_and_port_8,op_T0_and_port_6, op_T0_and_v);
  spice_node_3 n_n_171(eclk, ereset, n_171_port_3,n_171_port_0,n_171_port_1, n_171_v);
  spice_node_1 n_clk0(eclk, ereset, clk0_port_3, clk0_v);
  spice_node_2 n_op_T0_clc_sec(eclk, ereset, op_T0_clc_sec_port_8,op_T0_clc_sec_port_9, op_T0_clc_sec_v);
  spice_node_2 n__C56(eclk, ereset, _C56_port_8,_C56_port_4, _C56_v);
  spice_node_2 n_n_1209(eclk, ereset, n_1209_port_3,n_1209_port_5, n_1209_v);
  spice_node_5 n_n_1206(eclk, ereset, n_1206_port_2,n_1206_port_3,n_1206_port_0,n_1206_port_1,n_1206_port_4, n_1206_v);
  spice_node_2 n_n_1205(eclk, ereset, n_1205_port_4,n_1205_port_10, n_1205_v);
  spice_node_2 n_n_1202(eclk, ereset, n_1202_port_2,n_1202_port_3, n_1202_v);
  spice_node_2 n_n_1500(eclk, ereset, n_1500_port_3,n_1500_port_5, n_1500_v);
  spice_node_2 n__ABH3(eclk, ereset, _ABH3_port_3,_ABH3_port_1, _ABH3_v);
  spice_node_2 n__ABH2(eclk, ereset, _ABH2_port_2,_ABH2_port_3, _ABH2_v);
  spice_node_2 n__ABH1(eclk, ereset, _ABH1_port_3,_ABH1_port_0, _ABH1_v);
  spice_node_2 n__ABH0(eclk, ereset, _ABH0_port_2,_ABH0_port_3, _ABH0_v);
  spice_node_2 n__ABH7(eclk, ereset, _ABH7_port_2,_ABH7_port_3, _ABH7_v);
  spice_node_2 n__ABH6(eclk, ereset, _ABH6_port_2,_ABH6_port_3, _ABH6_v);
  spice_node_2 n__ABH5(eclk, ereset, _ABH5_port_2,_ABH5_port_3, _ABH5_v);
  spice_node_2 n__ABH4(eclk, ereset, _ABH4_port_2,_ABH4_port_3, _ABH4_v);
  spice_node_3 n_n_1507(eclk, ereset, n_1507_port_2,n_1507_port_3,n_1507_port_1, n_1507_v);
  spice_node_2 n_n_428(eclk, ereset, n_428_port_3,n_428_port_6, n_428_v);
  spice_node_2 n_n_424(eclk, ereset, n_424_port_2,n_424_port_1, n_424_v);
  spice_node_2 n_n_420(eclk, ereset, n_420_port_2,n_420_port_1, n_420_v);
  spice_node_3 n_n_423(eclk, ereset, n_423_port_2,n_423_port_0,n_423_port_1, n_423_v);
  spice_node_2 n_op_sty_cpy_mem(eclk, ereset, op_sty_cpy_mem_port_8,op_sty_cpy_mem_port_7, op_sty_cpy_mem_v);
  spice_node_3 n_n_1254(eclk, ereset, n_1254_port_2,n_1254_port_0,n_1254_port_1, n_1254_v);
  spice_node_2 n_dpc18__DAA(eclk, ereset, dpc18__DAA_port_2,dpc18__DAA_port_1, dpc18__DAA_v);
  spice_node_2 n_n_1720(eclk, ereset, n_1720_port_4,n_1720_port_5, n_1720_v);
  spice_node_2 n_AxB5(eclk, ereset, AxB5_port_6,AxB5_port_7, AxB5_v);
  spice_node_2 n_AxB7(eclk, ereset, AxB7_port_8,AxB7_port_6, AxB7_v);
  spice_node_2 n_AxB1(eclk, ereset, AxB1_port_8,AxB1_port_6, AxB1_v);
  spice_node_2 n_AxB3(eclk, ereset, AxB3_port_8,AxB3_port_6, AxB3_v);
  spice_node_2 n_op_T3_ind_y(eclk, ereset, op_T3_ind_y_port_6,op_T3_ind_y_port_7, op_T3_ind_y_v);
  spice_node_2 n_op_T3_ind_x(eclk, ereset, op_T3_ind_x_port_7,op_T3_ind_x_port_10, op_T3_ind_x_v);
  spice_node_2 n_n_1566(eclk, ereset, n_1566_port_3,n_1566_port_0, n_1566_v);
  spice_node_2 n_n_1561(eclk, ereset, n_1561_port_2,n_1561_port_0, n_1561_v);
  spice_node_2 n_n_1560(eclk, ereset, n_1560_port_4,n_1560_port_5, n_1560_v);
  spice_node_2 n_dpc38_PCLADL(eclk, ereset, dpc38_PCLADL_port_9,dpc38_PCLADL_port_0, dpc38_PCLADL_v);
  spice_node_3 n_n_1691(eclk, ereset, n_1691_port_8,n_1691_port_1,n_1691_port_7, n_1691_v);
  spice_node_2 n_n_1697(eclk, ereset, n_1697_port_2,n_1697_port_0, n_1697_v);
  spice_node_2 n_n_1696(eclk, ereset, n_1696_port_0,n_1696_port_1, n_1696_v);
  spice_node_2 n_x_op_T3_abs_idx(eclk, ereset, x_op_T3_abs_idx_port_6,x_op_T3_abs_idx_port_4, x_op_T3_abs_idx_v);
  spice_node_2 n_op_from_x(eclk, ereset, op_from_x_port_6,op_from_x_port_7, op_from_x_v);
  spice_node_2 n_n_855(eclk, ereset, n_855_port_2,n_855_port_0, n_855_v);
  spice_node_2 n_n_854(eclk, ereset, n_854_port_6,n_854_port_4, n_854_v);
  spice_node_2 n_n_850(eclk, ereset, n_850_port_3,n_850_port_0, n_850_v);
  spice_node_2 n_n_853(eclk, ereset, n_853_port_2,n_853_port_3, n_853_v);
  spice_node_2 n_n_852(eclk, ereset, n_852_port_2,n_852_port_3, n_852_v);
  spice_node_2 n_op_T0_cli_sei(eclk, ereset, op_T0_cli_sei_port_8,op_T0_cli_sei_port_9, op_T0_cli_sei_v);
  spice_node_2 n_op_T0_ldx_tax_tsx(eclk, ereset, op_T0_ldx_tax_tsx_port_8,op_T0_ldx_tax_tsx_port_6, op_T0_ldx_tax_tsx_v);
  spice_node_2 n_n_1229(eclk, ereset, n_1229_port_2,n_1229_port_3, n_1229_v);
  spice_node_2 n_n_1593(eclk, ereset, n_1593_port_2,n_1593_port_3, n_1593_v);
  spice_node_2 n_n_1222(eclk, ereset, n_1222_port_2,n_1222_port_0, n_1222_v);
  spice_node_2 n_n_1223(eclk, ereset, n_1223_port_4,n_1223_port_5, n_1223_v);
  spice_node_2 n_n_1225(eclk, ereset, n_1225_port_6,n_1225_port_5, n_1225_v);
  spice_node_2 n_n_1044(eclk, ereset, n_1044_port_3,n_1044_port_4, n_1044_v);
  spice_node_2 n_n_1594(eclk, ereset, n_1594_port_2,n_1594_port_3, n_1594_v);
  spice_node_2 n_n_1047(eclk, ereset, n_1047_port_2,n_1047_port_1, n_1047_v);
  spice_node_2 n_n_198(eclk, ereset, n_198_port_2,n_198_port_3, n_198_v);
  spice_node_2 n_n_628(eclk, ereset, n_628_port_4,n_628_port_5, n_628_v);
  spice_node_2 n_n_629(eclk, ereset, n_629_port_3,n_629_port_5, n_629_v);
  spice_node_2 n_n_626(eclk, ereset, n_626_port_3,n_626_port_6, n_626_v);
  spice_node_2 n_n_196(eclk, ereset, n_196_port_2,n_196_port_0, n_196_v);
  spice_node_2 n_n_625(eclk, ereset, n_625_port_4,n_625_port_5, n_625_v);
  spice_node_2 n_n_191(eclk, ereset, n_191_port_4,n_191_port_5, n_191_v);
  spice_node_2 n_n_192(eclk, ereset, n_192_port_8,n_192_port_4, n_192_v);
  spice_node_2 n_n_442(eclk, ereset, n_442_port_2,n_442_port_0, n_442_v);
  spice_node_2 n_n_440(eclk, ereset, n_440_port_7,n_440_port_10, n_440_v);
  spice_node_2 n_n_441(eclk, ereset, n_441_port_2,n_441_port_0, n_441_v);
  spice_node_2 n_n_445(eclk, ereset, n_445_port_3,n_445_port_4, n_445_v);
  spice_node_2 n_DBNeg(eclk, ereset, DBNeg_port_3,DBNeg_port_1, DBNeg_v);
  spice_node_2 n_op_T0_tsx(eclk, ereset, op_T0_tsx_port_9,op_T0_tsx_port_10, op_T0_tsx_v);
  spice_node_3 n_n_994(eclk, ereset, n_994_port_2,n_994_port_3,n_994_port_1, n_994_v);
  spice_node_2 n_n_995(eclk, ereset, n_995_port_2,n_995_port_1, n_995_v);
  spice_node_2 n_n_990(eclk, ereset, n_990_port_3,n_990_port_0, n_990_v);
  spice_node_2 n_n_992(eclk, ereset, n_992_port_2,n_992_port_0, n_992_v);
  spice_node_5 n_n_998(eclk, ereset, n_998_port_2,n_998_port_3,n_998_port_0,n_998_port_1,n_998_port_4, n_998_v);
  spice_node_3 n_n_999(eclk, ereset, n_999_port_2,n_999_port_3,n_999_port_1, n_999_v);
  spice_node_2 n__op_store(eclk, ereset, _op_store_port_2,_op_store_port_3, _op_store_v);
  spice_node_2 n_n_1501(eclk, ereset, n_1501_port_1,n_1501_port_4, n_1501_v);
  spice_node_2 n_op_T0_cpx_inx(eclk, ereset, op_T0_cpx_inx_port_9,op_T0_cpx_inx_port_7, op_T0_cpx_inx_v);
  spice_node_2 n_n_299(eclk, ereset, n_299_port_9,n_299_port_5, n_299_v);
  spice_node_2 n_n_298(eclk, ereset, n_298_port_3,n_298_port_4, n_298_v);
  spice_node_2 n_n_297(eclk, ereset, n_297_port_3,n_297_port_5, n_297_v);
  spice_node_5 n_n_296(eclk, ereset, n_296_port_3,n_296_port_0,n_296_port_1,n_296_port_4,n_296_port_5, n_296_v);
  spice_node_2 n_n_293(eclk, ereset, n_293_port_8,n_293_port_4, n_293_v);
  spice_node_2 n_n_291(eclk, ereset, n_291_port_2,n_291_port_3, n_291_v);
  spice_node_4 n_n_871(eclk, ereset, n_871_port_2,n_871_port_3,n_871_port_0,n_871_port_1, n_871_v);
  spice_node_2 n_n_877(eclk, ereset, n_877_port_3,n_877_port_5, n_877_v);
  spice_node_2 n_n_876(eclk, ereset, n_876_port_2,n_876_port_0, n_876_v);
  spice_node_2 n_n_875(eclk, ereset, n_875_port_3,n_875_port_5, n_875_v);
  spice_node_2 n_n_956(eclk, ereset, n_956_port_2,n_956_port_1, n_956_v);

endmodule

module spice_node_0(input eclk,ereset, output signed [`W-1:0] v);
  assign v = 0;
endmodule

module spice_node_1(input eclk,ereset, input signed [`W-1:0] i0, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_2(input eclk,ereset, input signed [`W-1:0] i0,i1, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_3(input eclk,ereset, input signed [`W-1:0] i0,i1,i2, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_4(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_5(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_6(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_7(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_8(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6,i7, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6+i7;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_12(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6+i7+i8+i9+i10+i11;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_13(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6+i7+i8+i9+i10+i11+i12;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

