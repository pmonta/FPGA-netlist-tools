* SPICE3 file created from 6800.ext - technology: 6800-nmos

.option scale=0.001u

M1000 diff_617000_6170000# diff_83000_3098000# diff_83000_3098000# GND efet w=82000 l=12000
+ ad=-1.30187e+09 pd=3.17e+06 as=1.89415e+09 ps=5.24546e+08 
M1001 diff_1120000_5760000# diff_1278000_5968000# diff_83000_3098000# GND efet w=162500 l=8500
+ ad=1.22803e+09 pd=652000 as=0 ps=0 
M1002 diff_83000_3098000# diff_1278000_5968000# diff_1128000_5767000# GND efet w=325500 l=8500
+ ad=0 pd=0 as=9.73294e+08 ps=4.164e+06 
M1003 diff_83000_3098000# diff_1278000_5968000# diff_1128000_5767000# GND efet w=326500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1004 diff_1120000_5760000# diff_1278000_5968000# diff_83000_3098000# GND efet w=162500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1005 diff_1278000_5968000# diff_1586000_6057000# diff_83000_3098000# GND efet w=304500 l=8500
+ ad=-5.30967e+08 pd=438000 as=0 ps=0 
M1006 diff_83000_3098000# diff_1278000_5968000# diff_1128000_5767000# GND efet w=326500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1007 diff_1120000_5760000# diff_1278000_5968000# diff_83000_3098000# GND efet w=152500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M1008 diff_83000_3098000# diff_1278000_5968000# diff_1128000_5767000# GND efet w=326000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1009 diff_95000_5192000# diff_1120000_5760000# diff_1120000_5760000# GND efet w=39000 l=9000
+ ad=-3.89442e+08 pd=2.0134e+08 as=0 ps=0 
M1010 diff_1278000_5968000# diff_1278000_5968000# diff_95000_5192000# GND efet w=27000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1011 diff_514000_5774000# diff_744000_5834000# diff_83000_3098000# GND efet w=120500 l=8500
+ ad=-6.79967e+08 pd=674000 as=0 ps=0 
M1012 diff_774000_5785000# diff_68000_5288000# diff_744000_5834000# GND efet w=13000 l=11000
+ ad=3.8e+08 pd=84000 as=-6.61967e+08 ps=552000 
M1013 diff_896000_5771000# diff_72000_4515000# diff_774000_5785000# GND efet w=13000 l=11000
+ ad=1.814e+09 pd=330000 as=0 ps=0 
M1014 diff_514000_5774000# diff_68000_5288000# diff_509000_5593000# GND efet w=20000 l=12000
+ ad=0 pd=0 as=3.05e+08 ps=102000 
M1015 diff_83000_3098000# diff_774000_5785000# diff_514000_5774000# GND efet w=111500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1016 diff_744000_5834000# diff_514000_5774000# diff_83000_3098000# GND efet w=96000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1017 diff_83000_3098000# diff_836000_5746000# diff_744000_5834000# GND efet w=114500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1018 diff_836000_5746000# diff_68000_5288000# diff_83000_3098000# GND efet w=65000 l=9000
+ ad=1.437e+09 pd=308000 as=0 ps=0 
M1019 diff_83000_3098000# diff_896000_5771000# diff_836000_5746000# GND efet w=68000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1020 diff_235000_3317000# diff_509000_5593000# diff_83000_3098000# GND efet w=130500 l=8500
+ ad=-1.82497e+09 pd=404000 as=0 ps=0 
M1021 diff_95000_5192000# diff_235000_3317000# diff_235000_3317000# GND efet w=13000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M1022 diff_83000_3098000# diff_969000_5800000# diff_896000_5771000# GND efet w=83000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1023 diff_896000_5771000# diff_896000_5771000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M1024 diff_83000_3098000# diff_617000_6170000# diff_969000_5800000# GND efet w=126000 l=10000
+ ad=0 pd=0 as=1.567e+09 ps=344000 
M1025 diff_95000_5192000# diff_617000_6170000# diff_617000_6170000# GND efet w=70000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1026 diff_1128000_5767000# diff_1120000_5760000# diff_95000_5192000# GND efet w=266000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1027 diff_1128000_5767000# diff_1120000_5760000# diff_95000_5192000# GND efet w=260000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1028 diff_1128000_5767000# diff_1120000_5760000# diff_95000_5192000# GND efet w=227000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1029 diff_1128000_5767000# diff_1120000_5760000# diff_95000_5192000# GND efet w=226500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1030 diff_1128000_5767000# diff_1120000_5760000# diff_95000_5192000# GND efet w=228000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1031 diff_1128000_5767000# diff_1120000_5760000# diff_95000_5192000# GND efet w=228000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1032 diff_1128000_5767000# diff_1120000_5760000# diff_95000_5192000# GND efet w=228000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1033 diff_514000_5774000# diff_514000_5774000# diff_95000_5192000# GND efet w=13000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M1034 diff_744000_5834000# diff_744000_5834000# diff_95000_5192000# GND efet w=12000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M1035 diff_836000_5746000# diff_836000_5746000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M1036 diff_1586000_6057000# diff_1586000_5876000# diff_83000_3098000# GND efet w=260000 l=9000
+ ad=1.11607e+09 pd=1.29e+06 as=0 ps=0 
M1037 diff_83000_3098000# diff_88000_5400000# diff_1586000_6057000# GND efet w=228000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1038 diff_1586000_6057000# diff_1648000_5847000# diff_83000_3098000# GND efet w=227000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1039 diff_83000_3098000# diff_197000_5470000# diff_1586000_6057000# GND efet w=227000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1040 diff_1586000_6057000# diff_1586000_6057000# diff_95000_5192000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1041 diff_969000_5800000# diff_969000_5800000# diff_95000_5192000# GND efet w=13000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1042 diff_1748000_6170000# diff_83000_3098000# diff_83000_3098000# GND efet w=93500 l=13500
+ ad=-1.33869e+08 pd=3.486e+06 as=0 ps=0 
M1043 diff_83000_3098000# diff_95000_5192000# diff_2049000_5823000# GND efet w=70000 l=10000
+ ad=0 pd=0 as=1.436e+09 ps=316000 
M1044 diff_83000_3098000# diff_1748000_6170000# diff_301000_4194000# GND efet w=125000 l=10000
+ ad=0 pd=0 as=-3.06967e+08 ps=808000 
M1045 diff_95000_5192000# diff_301000_4194000# diff_301000_4194000# GND efet w=14000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1046 diff_571000_4610000# diff_68000_5288000# diff_1586000_5876000# GND efet w=15000 l=11000
+ ad=-6.20967e+08 pd=676000 as=2.74e+08 ps=92000 
M1047 diff_83000_3098000# diff_474000_5143000# diff_506000_5537000# GND efet w=95500 l=9500
+ ad=0 pd=0 as=-3.59935e+08 ps=1.082e+06 
M1048 diff_506000_5537000# diff_474000_5143000# diff_83000_3098000# GND efet w=94500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1049 diff_135000_5507000# diff_91000_5337000# diff_83000_3098000# GND efet w=213000 l=8000
+ ad=-1.73493e+09 pd=954000 as=0 ps=0 
M1050 diff_83000_3098000# diff_474000_5143000# diff_506000_5537000# GND efet w=105000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1051 diff_83000_3098000# diff_91000_5337000# diff_135000_5507000# GND efet w=76000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1052 diff_95000_5192000# diff_506000_5537000# diff_506000_5537000# GND efet w=28000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1053 diff_95000_5192000# diff_835000_5621000# diff_835000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-5.06967e+08 ps=852000 
M1054 diff_95000_5192000# diff_894000_5621000# diff_894000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-3.83967e+08 ps=868000 
M1055 diff_95000_5192000# diff_761000_5561000# diff_761000_5561000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-5.93967e+08 ps=788000 
M1056 diff_95000_5192000# diff_797000_5587000# diff_797000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-8.18967e+08 ps=754000 
M1057 diff_95000_5192000# diff_953000_5621000# diff_953000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-1.29673e+07 ps=900000 
M1058 diff_95000_5192000# diff_855000_5587000# diff_855000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-1.16297e+09 ps=720000 
M1059 diff_95000_5192000# diff_1012000_5621000# diff_1012000_5621000# GND efet w=11000 l=47000
+ ad=0 pd=0 as=-5.61967e+08 ps=858000 
M1060 diff_95000_5192000# diff_914000_5587000# diff_914000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-9.98967e+08 ps=736000 
M1061 diff_95000_5192000# diff_973000_5587000# diff_973000_5587000# GND efet w=14000 l=47000
+ ad=0 pd=0 as=-8.95967e+08 ps=746000 
M1062 diff_95000_5192000# diff_1032000_5587000# diff_1032000_5587000# GND efet w=14000 l=47000
+ ad=0 pd=0 as=-5.09967e+08 ps=786000 
M1063 diff_95000_5192000# diff_1110000_5621000# diff_1110000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-4.29967e+08 ps=858000 
M1064 diff_95000_5192000# diff_1169000_5621000# diff_1169000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-1.03967e+08 ps=890000 
M1065 diff_95000_5192000# diff_1228000_5621000# diff_1228000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-5.95967e+08 ps=848000 
M1066 diff_95000_5192000# diff_1130000_5587000# diff_1130000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-9.64967e+08 ps=740000 
M1067 diff_95000_5192000# diff_1286000_5621000# diff_1286000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-3.10967e+08 ps=870000 
M1068 diff_95000_5192000# diff_1188000_5587000# diff_1188000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-9.78967e+08 ps=738000 
M1069 diff_95000_5192000# diff_1346000_5621000# diff_1346000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-6.18967e+08 ps=846000 
M1070 diff_95000_5192000# diff_1248000_5587000# diff_1248000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-8.59967e+08 ps=750000 
M1071 diff_95000_5192000# diff_1404000_5621000# diff_1404000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-3.75967e+08 ps=864000 
M1072 diff_95000_5192000# diff_1306000_5587000# diff_1306000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-8.83967e+08 ps=748000 
M1073 diff_95000_5192000# diff_1464000_5621000# diff_1464000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-2.16967e+08 ps=886000 
M1074 diff_95000_5192000# diff_1366000_5587000# diff_1366000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-6.29967e+08 ps=774000 
M1075 diff_95000_5192000# diff_1522000_5621000# diff_1522000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=9.80327e+07 ps=912000 
M1076 diff_95000_5192000# diff_1424000_5587000# diff_1424000_5587000# GND efet w=14000 l=47000
+ ad=0 pd=0 as=-6.60967e+08 ps=770000 
M1077 diff_95000_5192000# diff_1484000_5587000# diff_1484000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-9.93967e+08 ps=736000 
M1078 diff_95000_5192000# diff_1542000_5587000# diff_1542000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-1.09897e+09 ps=728000 
M1079 diff_95000_5192000# diff_1619000_5621000# diff_1619000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-4.23967e+08 ps=866000 
M1080 diff_95000_5192000# diff_1678000_5621000# diff_1678000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-2.22967e+08 ps=880000 
M1081 diff_95000_5192000# diff_1737000_5621000# diff_1737000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-5.08967e+08 ps=856000 
M1082 diff_95000_5192000# diff_1639000_5587000# diff_1639000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-1.08497e+09 ps=728000 
M1083 diff_95000_5192000# diff_1795000_5621000# diff_1795000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-2.69967e+08 ps=874000 
M1084 diff_95000_5192000# diff_1698000_5587000# diff_1698000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-5.57967e+08 ps=782000 
M1085 diff_2071000_5823000# diff_72000_4515000# diff_2049000_5823000# GND efet w=12000 l=11000
+ ad=1.2e+08 pd=44000 as=0 ps=0 
M1086 diff_2092000_5823000# diff_68000_5288000# diff_2071000_5823000# GND efet w=12000 l=11000
+ ad=4.17e+08 pd=108000 as=0 ps=0 
M1087 diff_2092000_5823000# diff_1748000_6170000# diff_1748000_6170000# GND efet w=10000 l=74000
+ ad=0 pd=0 as=0 ps=0 
M1088 diff_83000_3098000# diff_83000_3098000# diff_83000_3098000# GND efet w=1000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M1089 diff_83000_3098000# diff_83000_3098000# diff_68000_5288000# GND efet w=78000 l=13000
+ ad=0 pd=0 as=-1.78693e+09 ps=708000 
M1090 diff_2157000_5726000# diff_2049000_5823000# diff_1748000_6170000# GND efet w=12000 l=11000
+ ad=1.8e+08 pd=54000 as=0 ps=0 
M1091 diff_2194000_5726000# diff_83000_3098000# diff_2157000_5726000# GND efet w=12000 l=22000
+ ad=-1.16787e+09 pd=3.336e+06 as=0 ps=0 
M1092 diff_83000_3098000# diff_83000_3098000# diff_2194000_5726000# GND efet w=80000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M1093 diff_2523000_5770000# diff_2194000_5726000# diff_83000_3098000# GND efet w=137000 l=10000
+ ad=-1.87997e+09 pd=458000 as=0 ps=0 
M1094 diff_2621000_5834000# diff_2613000_5827000# diff_83000_3098000# GND efet w=124000 l=8000
+ ad=1.903e+09 pd=430000 as=0 ps=0 
M1095 diff_83000_3098000# diff_1581000_4325000# diff_2748000_5772000# GND efet w=69500 l=8500
+ ad=0 pd=0 as=1.662e+09 ps=336000 
M1096 diff_2621000_5834000# diff_2621000_5834000# diff_95000_5192000# GND efet w=12000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M1097 diff_2613000_5827000# diff_68000_5288000# diff_2523000_5770000# GND efet w=12000 l=11000
+ ad=3.12e+08 pd=96000 as=0 ps=0 
M1098 diff_2523000_5770000# diff_2523000_5770000# diff_95000_5192000# GND efet w=13000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M1099 diff_83000_3098000# diff_2621000_5834000# diff_2748000_5772000# GND efet w=64000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1100 diff_2841000_5928000# diff_2833000_5761000# diff_83000_3098000# GND efet w=112000 l=9000
+ ad=-6.79673e+07 pd=792000 as=0 ps=0 
M1101 diff_83000_3098000# diff_94000_3551000# diff_2841000_5928000# GND efet w=109000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1102 diff_2841000_5928000# diff_2877000_5745000# diff_83000_3098000# GND efet w=111500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1103 diff_2877000_5745000# diff_2841000_5928000# diff_83000_3098000# GND efet w=126000 l=8000
+ ad=5.37033e+08 pd=902000 as=0 ps=0 
M1104 diff_2877000_5745000# diff_2983000_5746000# diff_83000_3098000# GND efet w=133500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M1105 diff_197000_5470000# diff_3099000_5787000# diff_83000_3098000# GND efet w=425500 l=7500
+ ad=1.66307e+09 pd=1.692e+06 as=0 ps=0 
M1106 diff_2748000_5772000# diff_2748000_5772000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M1107 diff_2833000_5761000# diff_72000_4515000# diff_2621000_5834000# GND efet w=13000 l=11000
+ ad=5.69e+08 pd=134000 as=0 ps=0 
M1108 diff_2841000_5928000# diff_2841000_5928000# diff_95000_5192000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M1109 diff_2877000_5745000# diff_68000_5288000# diff_2833000_5761000# GND efet w=14000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1110 diff_3099000_5787000# diff_68000_5288000# diff_2877000_5745000# GND efet w=34000 l=11000
+ ad=4.76e+08 pd=124000 as=0 ps=0 
M1111 diff_2748000_5772000# diff_72000_4515000# diff_2983000_5746000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=7.4e+08 ps=158000 
M1112 diff_2983000_5746000# diff_68000_5288000# diff_2841000_5928000# GND efet w=13000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1113 diff_197000_5470000# diff_94000_3551000# diff_83000_3098000# GND efet w=330000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M1114 diff_3583000_5810000# diff_3505000_5809000# diff_83000_3098000# GND efet w=122500 l=8500
+ ad=-1.69897e+09 pd=500000 as=0 ps=0 
M1115 diff_197000_5470000# diff_94000_3551000# diff_83000_3098000# GND efet w=24000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M1116 diff_197000_5470000# diff_94000_3551000# diff_83000_3098000# GND efet w=62000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M1117 diff_94000_3551000# diff_3505000_5809000# diff_95000_5192000# GND efet w=25000 l=7000
+ ad=1.15003e+09 pd=734000 as=0 ps=0 
M1118 diff_197000_5470000# diff_197000_5470000# diff_95000_5192000# GND efet w=25000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1119 diff_94000_3551000# diff_3505000_5809000# diff_95000_5192000# GND efet w=200500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M1120 diff_2877000_5745000# diff_2877000_5745000# diff_95000_5192000# GND efet w=12000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M1121 diff_95000_5192000# diff_1944000_5621000# diff_1944000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-4.46967e+08 ps=862000 
M1122 diff_95000_5192000# diff_1757000_5587000# diff_1757000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-6.21967e+08 ps=776000 
M1123 diff_95000_5192000# diff_2002000_5621000# diff_2002000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-4.41967e+08 ps=856000 
M1124 diff_95000_5192000# diff_1815000_5587000# diff_1815000_5587000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-9.55967e+08 ps=742000 
M1125 diff_95000_5192000# diff_2061000_5621000# diff_2061000_5621000# GND efet w=11000 l=47000
+ ad=0 pd=0 as=-2.87967e+08 ps=886000 
M1126 diff_95000_5192000# diff_1964000_5587000# diff_1964000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-9.20967e+08 ps=746000 
M1127 diff_95000_5192000# diff_2119000_5621000# diff_2119000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-9.89673e+07 ps=892000 
M1128 diff_95000_5192000# diff_2022000_5587000# diff_2022000_5587000# GND efet w=14000 l=47000
+ ad=0 pd=0 as=-8.98967e+08 ps=746000 
M1129 diff_95000_5192000# diff_2081000_5587000# diff_2081000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-9.53967e+08 ps=742000 
M1130 diff_95000_5192000# diff_2139000_5587000# diff_2139000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-6.91967e+08 ps=768000 
M1131 diff_95000_5192000# diff_2218000_5621000# diff_2218000_5621000# GND efet w=14000 l=47000
+ ad=0 pd=0 as=-3.03967e+08 ps=864000 
M1132 diff_95000_5192000# diff_2276000_5621000# diff_2276000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=9.50327e+07 ps=912000 
M1133 diff_95000_5192000# diff_2335000_5621000# diff_2335000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-2.54967e+08 ps=882000 
M1134 diff_95000_5192000# diff_2238000_5587000# diff_2238000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-8.59967e+08 ps=752000 
M1135 diff_95000_5192000# diff_2394000_5621000# diff_2394000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-4.42967e+08 ps=856000 
M1136 diff_95000_5192000# diff_2296000_5587000# diff_2296000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-1.01697e+09 ps=734000 
M1137 diff_94000_3551000# diff_3583000_5810000# diff_83000_3098000# GND efet w=366500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M1138 diff_1648000_5847000# diff_3695000_5841000# diff_3677000_5839000# GND efet w=106500 l=7500
+ ad=-1.70597e+09 pd=404000 as=3.30033e+08 ps=888000 
M1139 diff_3677000_5839000# diff_3695000_5841000# diff_1648000_5847000# GND efet w=159000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1140 diff_83000_3098000# diff_3757000_5782000# diff_3677000_5839000# GND efet w=149000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1141 diff_83000_3098000# diff_3757000_5782000# diff_3505000_5809000# GND efet w=182500 l=8500
+ ad=0 pd=0 as=2.127e+09 ps=426000 
M1142 diff_3583000_5810000# diff_3505000_5809000# diff_83000_3098000# GND efet w=32000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1143 diff_95000_5192000# diff_3583000_5810000# diff_3583000_5810000# GND efet w=12000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1144 diff_1648000_5847000# diff_1648000_5847000# diff_95000_5192000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1145 diff_3677000_5839000# diff_3757000_5782000# diff_83000_3098000# GND efet w=99000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1146 diff_83000_3098000# diff_3884000_5844000# diff_3872000_5819000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=1.52033e+08 ps=874000 
M1147 diff_3903000_5737000# diff_3872000_5819000# diff_83000_3098000# GND efet w=55000 l=8000
+ ad=-1.35897e+09 pd=516000 as=0 ps=0 
M1148 diff_83000_3098000# diff_3884000_5844000# diff_3872000_5819000# GND efet w=79000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1149 diff_83000_3098000# diff_3962000_5824000# diff_3903000_5737000# GND efet w=119000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1150 diff_83000_3098000# diff_3962000_5824000# diff_3884000_5844000# GND efet w=68500 l=8500
+ ad=0 pd=0 as=-2.02997e+09 ps=412000 
M1151 diff_3903000_5737000# diff_3872000_5819000# diff_83000_3098000# GND efet w=59500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M1152 diff_83000_3098000# diff_68000_5288000# diff_3884000_5844000# GND efet w=74500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M1153 diff_3872000_5819000# diff_3903000_5737000# diff_83000_3098000# GND efet w=115000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1154 diff_3884000_5844000# diff_3884000_5844000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M1155 diff_3962000_5824000# diff_68000_5288000# diff_3872000_5819000# GND efet w=28000 l=12000
+ ad=8.84e+08 pd=232000 as=0 ps=0 
M1156 diff_83000_3098000# diff_4198000_5803000# diff_3695000_5841000# GND efet w=102500 l=8500
+ ad=0 pd=0 as=2.132e+09 ps=466000 
M1157 diff_3505000_5809000# diff_3505000_5809000# diff_95000_5192000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1158 diff_3872000_5819000# diff_68000_5288000# diff_3757000_5782000# GND efet w=27000 l=11000
+ ad=0 pd=0 as=3.59e+08 ps=106000 
M1159 diff_3903000_5737000# diff_3903000_5737000# diff_95000_5192000# GND efet w=13000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M1160 diff_3695000_5841000# diff_72000_4515000# diff_3962000_5824000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1161 diff_83000_3098000# diff_4056000_6171000# diff_4198000_5803000# GND efet w=128500 l=10500
+ ad=0 pd=0 as=1.555e+09 ps=324000 
M1162 diff_4427000_5701000# diff_4356000_5717000# diff_83000_3098000# GND efet w=178500 l=9500
+ ad=1.776e+09 pd=280000 as=0 ps=0 
M1163 diff_95000_5192000# diff_3872000_5819000# diff_3872000_5819000# GND efet w=13000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M1164 diff_3695000_5841000# diff_3695000_5841000# diff_95000_5192000# GND efet w=12000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M1165 diff_4056000_6171000# diff_83000_3098000# diff_83000_3098000# GND efet w=79000 l=12000
+ ad=4.36098e+08 pd=2.726e+06 as=0 ps=0 
M1166 diff_88000_5400000# diff_4356000_5717000# diff_83000_3098000# GND efet w=188500 l=9500
+ ad=-1.58293e+09 pd=934000 as=0 ps=0 
M1167 diff_88000_5400000# diff_4356000_5717000# diff_83000_3098000# GND efet w=228500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1168 diff_95000_5192000# diff_4427000_5701000# diff_88000_5400000# GND efet w=319500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1169 diff_4198000_5803000# diff_4198000_5803000# diff_95000_5192000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1170 diff_4056000_6171000# diff_4056000_6171000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M1171 diff_95000_5192000# diff_4427000_5701000# diff_88000_5400000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1172 diff_4427000_5701000# diff_4427000_5701000# diff_95000_5192000# GND efet w=11000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1173 diff_4356000_5717000# diff_4356000_5717000# diff_95000_5192000# GND efet w=12000 l=12000
+ ad=1.693e+09 pd=324000 as=0 ps=0 
M1174 diff_83000_3098000# diff_4398000_6171000# diff_4356000_5717000# GND efet w=133500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M1175 diff_4398000_6171000# diff_83000_3098000# diff_83000_3098000# GND efet w=80000 l=12000
+ ad=1.4271e+09 pd=2.822e+06 as=0 ps=0 
M1176 diff_5087000_472000# diff_5406000_5992000# diff_83000_3098000# GND efet w=699000 l=8000
+ ad=6.28131e+08 pd=1.998e+06 as=0 ps=0 
M1177 diff_5087000_472000# diff_5406000_5992000# diff_83000_3098000# GND efet w=168000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1178 diff_83000_3098000# diff_5772000_6155000# diff_5761000_6140000# GND efet w=403500 l=8500
+ ad=0 pd=0 as=1.76307e+09 ps=1.47e+06 
M1179 diff_5430000_5898000# diff_5453000_5802000# diff_83000_3098000# GND efet w=204000 l=9000
+ ad=1.787e+09 pd=282000 as=0 ps=0 
M1180 diff_83000_3098000# diff_5406000_5992000# diff_5087000_472000# GND efet w=75500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M1181 diff_83000_3098000# diff_5406000_5992000# diff_5087000_472000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1182 diff_83000_3098000# diff_135000_5507000# diff_5761000_6140000# GND efet w=381500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1183 diff_5430000_5898000# diff_5430000_5898000# diff_95000_5192000# GND efet w=12000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1184 diff_5772000_6155000# diff_68000_5288000# diff_5507000_5789000# GND efet w=34000 l=13000
+ ad=4.27e+08 pd=116000 as=-1.20497e+09 ps=682000 
M1185 diff_5406000_5992000# diff_5173000_5735000# diff_83000_3098000# GND efet w=72500 l=9500
+ ad=1.696e+09 pd=334000 as=0 ps=0 
M1186 diff_5259000_5770000# diff_5430000_5898000# diff_5406000_5992000# GND efet w=74500 l=9500
+ ad=-1.73793e+09 pd=902000 as=0 ps=0 
M1187 diff_95000_5192000# diff_2483000_5621000# diff_2483000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-8.09673e+07 ps=900000 
M1188 diff_95000_5192000# diff_2355000_5587000# diff_2355000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-5.13967e+08 ps=786000 
M1189 diff_95000_5192000# diff_2541000_5621000# diff_2541000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-3.48967e+08 ps=866000 
M1190 diff_95000_5192000# diff_2414000_5587000# diff_2414000_5587000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-9.88967e+08 ps=738000 
M1191 diff_95000_5192000# diff_2600000_5621000# diff_2600000_5621000# GND efet w=11000 l=47000
+ ad=0 pd=0 as=-5.39967e+08 ps=852000 
M1192 diff_95000_5192000# diff_2503000_5587000# diff_2503000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-4.87967e+08 ps=788000 
M1193 diff_95000_5192000# diff_2659000_5621000# diff_2659000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-3.12967e+08 ps=870000 
M1194 diff_95000_5192000# diff_2561000_5587000# diff_2561000_5587000# GND efet w=14000 l=47000
+ ad=0 pd=0 as=-8.86967e+08 ps=748000 
M1195 diff_95000_5192000# diff_2620000_5587000# diff_2620000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-6.31967e+08 ps=774000 
M1196 diff_95000_5192000# diff_2679000_5587000# diff_2679000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-7.67967e+08 ps=760000 
M1197 diff_95000_5192000# diff_2757000_5621000# diff_2757000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-4.42967e+08 ps=856000 
M1198 diff_95000_5192000# diff_2815000_5621000# diff_2815000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-2.75967e+08 ps=874000 
M1199 diff_95000_5192000# diff_2874000_5621000# diff_2874000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-1.22967e+08 ps=896000 
M1200 diff_95000_5192000# diff_2777000_5587000# diff_2777000_5587000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-1.00597e+09 ps=738000 
M1201 diff_95000_5192000# diff_2933000_5621000# diff_2933000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-3.48967e+08 ps=866000 
M1202 diff_95000_5192000# diff_2835000_5587000# diff_2835000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-7.39967e+08 ps=764000 
M1203 diff_95000_5192000# diff_2992000_5621000# diff_2992000_5621000# GND efet w=11000 l=47000
+ ad=0 pd=0 as=-5.46967e+08 ps=860000 
M1204 diff_95000_5192000# diff_2894000_5587000# diff_2894000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-5.71967e+08 ps=780000 
M1205 diff_95000_5192000# diff_3051000_5621000# diff_3051000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-8.19673e+07 ps=900000 
M1206 diff_95000_5192000# diff_2953000_5587000# diff_2953000_5587000# GND efet w=14000 l=47000
+ ad=0 pd=0 as=-8.71967e+08 ps=748000 
M1207 diff_95000_5192000# diff_3110000_5621000# diff_3110000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-5.19967e+08 ps=850000 
M1208 diff_95000_5192000# diff_3012000_5587000# diff_3012000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-6.91967e+08 ps=768000 
M1209 diff_95000_5192000# diff_3169000_5621000# diff_3169000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-4.43967e+08 ps=862000 
M1210 diff_95000_5192000# diff_3071000_5587000# diff_3071000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-8.37967e+08 ps=752000 
M1211 diff_95000_5192000# diff_3130000_5587000# diff_3130000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-4.48967e+08 ps=794000 
M1212 diff_95000_5192000# diff_3189000_5587000# diff_3189000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-8.10967e+08 ps=756000 
M1213 diff_95000_5192000# diff_3266000_5621000# diff_3266000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-2.04967e+08 ps=882000 
M1214 diff_95000_5192000# diff_3324000_5621000# diff_3324000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-3.10967e+08 ps=876000 
M1215 diff_95000_5192000# diff_3383000_5621000# diff_3383000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-1.71967e+08 ps=892000 
M1216 diff_95000_5192000# diff_3286000_5587000# diff_3286000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-9.65967e+08 ps=740000 
M1217 diff_95000_5192000# diff_3442000_5621000# diff_3442000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-3.74967e+08 ps=864000 
M1218 diff_95000_5192000# diff_3344000_5587000# diff_3344000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-8.49967e+08 ps=752000 
M1219 diff_95000_5192000# diff_3501000_5621000# diff_3501000_5621000# GND efet w=11000 l=47000
+ ad=0 pd=0 as=-5.46967e+08 ps=860000 
M1220 diff_95000_5192000# diff_3403000_5587000# diff_3403000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-1.05097e+09 ps=732000 
M1221 diff_95000_5192000# diff_3560000_5621000# diff_3560000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=8.30327e+07 ps=910000 
M1222 diff_95000_5192000# diff_3462000_5587000# diff_3462000_5587000# GND efet w=14000 l=47000
+ ad=0 pd=0 as=-8.36967e+08 ps=754000 
M1223 diff_95000_5192000# diff_3619000_5621000# diff_3619000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-4.33967e+08 ps=858000 
M1224 diff_95000_5192000# diff_3521000_5587000# diff_3521000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-9.92967e+08 ps=738000 
M1225 diff_95000_5192000# diff_3678000_5621000# diff_3678000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-3.69673e+07 ps=898000 
M1226 diff_95000_5192000# diff_3580000_5587000# diff_3580000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-6.50967e+08 ps=772000 
M1227 diff_95000_5192000# diff_3639000_5587000# diff_3639000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-6.16967e+08 ps=776000 
M1228 diff_95000_5192000# diff_3698000_5587000# diff_3698000_5587000# GND efet w=14000 l=47000
+ ad=0 pd=0 as=-1.05397e+09 ps=728000 
M1229 diff_95000_5192000# diff_3776000_5621000# diff_3776000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-4.12967e+08 ps=860000 
M1230 diff_95000_5192000# diff_3834000_5621000# diff_3834000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-2.9673e+06 ps=902000 
M1231 diff_95000_5192000# diff_3893000_5621000# diff_3893000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-3.28967e+08 ps=876000 
M1232 diff_95000_5192000# diff_3796000_5587000# diff_3796000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-7.34967e+08 ps=764000 
M1233 diff_95000_5192000# diff_3952000_5621000# diff_3952000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-1.37967e+08 ps=888000 
M1234 diff_95000_5192000# diff_3854000_5587000# diff_3854000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-8.91967e+08 ps=748000 
M1235 diff_95000_5192000# diff_4011000_5621000# diff_4011000_5621000# GND efet w=11000 l=47000
+ ad=0 pd=0 as=-2.72967e+08 ps=888000 
M1236 diff_95000_5192000# diff_3913000_5587000# diff_3913000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-9.44967e+08 ps=742000 
M1237 diff_95000_5192000# diff_4070000_5621000# diff_4070000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-2.9673e+06 ps=908000 
M1238 diff_95000_5192000# diff_3972000_5587000# diff_3972000_5587000# GND efet w=14000 l=47000
+ ad=0 pd=0 as=-8.82967e+08 ps=748000 
M1239 diff_95000_5192000# diff_4129000_5621000# diff_4129000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-2.69967e+08 ps=876000 
M1240 diff_95000_5192000# diff_4031000_5587000# diff_4031000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-7.46967e+08 ps=762000 
M1241 diff_95000_5192000# diff_4188000_5621000# diff_4188000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-5.82967e+08 ps=848000 
M1242 diff_95000_5192000# diff_4090000_5587000# diff_4090000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-1.16297e+09 ps=720000 
M1243 diff_95000_5192000# diff_4149000_5587000# diff_4149000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-6.21967e+08 ps=776000 
M1244 diff_95000_5192000# diff_4208000_5587000# diff_4208000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-7.15967e+08 ps=766000 
M1245 diff_95000_5192000# diff_4288000_5621000# diff_4288000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-2.55967e+08 ps=882000 
M1246 diff_95000_5192000# diff_4346000_5621000# diff_4346000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-4.43967e+08 ps=864000 
M1247 diff_95000_5192000# diff_4405000_5621000# diff_4405000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-4.28967e+08 ps=864000 
M1248 diff_95000_5192000# diff_4307000_5587000# diff_4307000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-9.80967e+08 ps=738000 
M1249 diff_95000_5192000# diff_4464000_5621000# diff_4464000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-4.90967e+08 ps=852000 
M1250 diff_95000_5192000# diff_4366000_5587000# diff_4366000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-1.07597e+09 ps=728000 
M1251 diff_95000_5192000# diff_4523000_5621000# diff_4523000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-1.81967e+08 ps=890000 
M1252 diff_95000_5192000# diff_4425000_5587000# diff_4425000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-8.78967e+08 ps=750000 
M1253 diff_95000_5192000# diff_4582000_5621000# diff_4582000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-3.88967e+08 ps=870000 
M1254 diff_95000_5192000# diff_4484000_5587000# diff_4484000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-8.21967e+08 ps=756000 
M1255 diff_83000_3098000# diff_83000_3098000# diff_72000_4515000# GND efet w=80000 l=13000
+ ad=0 pd=0 as=8.48033e+08 ps=520000 
M1256 diff_5067000_5900000# diff_83000_3098000# diff_83000_3098000# GND efet w=81000 l=13000
+ ad=1.5361e+09 pd=2.764e+06 as=0 ps=0 
M1257 diff_83000_3098000# diff_5067000_5900000# diff_5173000_5735000# GND efet w=310500 l=8500
+ ad=0 pd=0 as=7.37033e+08 ps=804000 
M1258 diff_83000_3098000# diff_5173000_5735000# diff_5259000_5770000# GND efet w=379500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1259 diff_95000_5192000# diff_5173000_5735000# diff_5173000_5735000# GND efet w=24000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1260 diff_5402000_5747000# diff_5259000_5770000# diff_83000_3098000# GND efet w=247500 l=9500
+ ad=1.874e+09 pd=360000 as=0 ps=0 
M1261 diff_5087000_472000# diff_5402000_5747000# diff_95000_5192000# GND efet w=113000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1262 diff_5087000_472000# diff_5402000_5747000# diff_95000_5192000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1263 diff_95000_5192000# diff_5402000_5747000# diff_5087000_472000# GND efet w=275000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1264 diff_5928000_6128000# diff_5761000_6140000# diff_83000_3098000# GND efet w=838000 l=8000
+ ad=-2.03274e+09 pd=4.152e+06 as=0 ps=0 
M1265 diff_5928000_6128000# diff_5761000_6140000# diff_83000_3098000# GND efet w=597000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1266 diff_5928000_6128000# diff_5775000_5847000# diff_95000_5192000# GND efet w=481000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1267 diff_95000_5192000# diff_5761000_6140000# diff_5761000_6140000# GND efet w=35000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1268 diff_95000_5192000# diff_5775000_5847000# diff_5775000_5847000# GND efet w=41000 l=9000
+ ad=0 pd=0 as=-1.7559e+09 ps=1.596e+06 
M1269 diff_5775000_5847000# diff_5761000_6140000# diff_83000_3098000# GND efet w=493000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1270 diff_95000_5192000# diff_5775000_5847000# diff_5928000_6128000# GND efet w=238500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1271 diff_5775000_5847000# diff_135000_5507000# diff_83000_3098000# GND efet w=125000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1272 diff_95000_5192000# diff_5775000_5847000# diff_5928000_6128000# GND efet w=240500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M1273 diff_5775000_5847000# diff_135000_5507000# diff_83000_3098000# GND efet w=269000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1274 diff_5928000_6128000# diff_5775000_5847000# diff_95000_5192000# GND efet w=679000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1275 diff_5487000_5789000# diff_5402000_5747000# diff_5453000_5802000# GND efet w=35000 l=12000
+ ad=3.15e+08 pd=88000 as=5.74e+08 ps=124000 
M1276 diff_5507000_5789000# diff_68000_5288000# diff_5487000_5789000# GND efet w=35000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1277 diff_5402000_5747000# diff_5402000_5747000# diff_95000_5192000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1278 diff_5259000_5770000# diff_5259000_5770000# diff_95000_5192000# GND efet w=34000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1279 diff_4478000_4817000# diff_72000_4515000# diff_6105000_5745000# GND efet w=20000 l=12000
+ ad=1.12303e+09 pd=980000 as=3.36e+08 ps=112000 
M1280 diff_95000_5192000# diff_5507000_5789000# diff_5507000_5789000# GND efet w=13000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M1281 diff_5507000_5789000# diff_6105000_5745000# diff_83000_3098000# GND efet w=159000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1282 diff_95000_5192000# diff_4730000_5621000# diff_4730000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-1.91967e+08 ps=890000 
M1283 diff_95000_5192000# diff_4543000_5587000# diff_4543000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-1.06097e+09 ps=730000 
M1284 diff_95000_5192000# diff_4788000_5621000# diff_4788000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-4.99967e+08 ps=858000 
M1285 diff_95000_5192000# diff_4602000_5587000# diff_4602000_5587000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-9.11967e+08 ps=746000 
M1286 diff_95000_5192000# diff_4847000_5621000# diff_4847000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-1.51967e+08 ps=894000 
M1287 diff_95000_5192000# diff_4750000_5587000# diff_4750000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-9.00967e+08 ps=746000 
M1288 diff_95000_5192000# diff_4906000_5621000# diff_4906000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-1.89967e+08 ps=890000 
M1289 diff_95000_5192000# diff_4808000_5587000# diff_4808000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-8.47967e+08 ps=752000 
M1290 diff_95000_5192000# diff_4867000_5587000# diff_4867000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-6.43967e+08 ps=772000 
M1291 diff_95000_5192000# diff_4926000_5587000# diff_4926000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-7.22967e+08 ps=764000 
M1292 diff_95000_5192000# diff_5004000_5621000# diff_5004000_5621000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-4.96967e+08 ps=852000 
M1293 diff_95000_5192000# diff_5062000_5621000# diff_5062000_5621000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-5.70967e+08 ps=852000 
M1294 diff_775000_5479000# diff_775000_5479000# diff_95000_5192000# GND efet w=14000 l=8000
+ ad=5.30033e+08 pd=954000 as=0 ps=0 
M1295 diff_775000_5479000# diff_5252000_5062000# diff_83000_3098000# GND efet w=182000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1296 diff_775000_5479000# diff_5501000_5678000# diff_83000_3098000# GND efet w=189000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1297 diff_83000_3098000# diff_5502000_5646000# diff_5501000_5678000# GND efet w=101500 l=7500
+ ad=0 pd=0 as=-1.56097e+09 ps=708000 
M1298 diff_83000_3098000# diff_5252000_5062000# diff_775000_5448000# GND efet w=179500 l=8500
+ ad=0 pd=0 as=1.98103e+09 ps=954000 
M1299 diff_775000_5448000# diff_5502000_5646000# diff_83000_3098000# GND efet w=179000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1300 diff_95000_5192000# diff_5024000_5587000# diff_5024000_5587000# GND efet w=13000 l=47000
+ ad=0 pd=0 as=-1.10297e+09 ps=726000 
M1301 diff_95000_5192000# diff_775000_5448000# diff_775000_5448000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1302 diff_95000_5192000# diff_5082000_5587000# diff_5082000_5587000# GND efet w=12000 l=47000
+ ad=0 pd=0 as=-1.22297e+09 ps=712000 
M1303 diff_761000_5561000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1304 diff_797000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1305 diff_835000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1306 diff_855000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1307 diff_894000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=17000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1308 diff_914000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1309 diff_953000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1310 diff_973000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1311 diff_1012000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=17000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1312 diff_1032000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1313 diff_135000_5507000# diff_135000_5507000# diff_95000_5192000# GND efet w=25000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1314 diff_506000_5537000# diff_402000_4713000# diff_83000_3098000# GND efet w=140000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1315 diff_1110000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1316 diff_1130000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1317 diff_1169000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1318 diff_1188000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1319 diff_1228000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1320 diff_1248000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1321 diff_1286000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1322 diff_1306000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1323 diff_1346000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=17000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1324 diff_1366000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1325 diff_1404000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1326 diff_1424000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1327 diff_1464000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=17000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1328 diff_1484000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1329 diff_1522000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1330 diff_1542000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1331 diff_1619000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1332 diff_1639000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1333 diff_1678000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1334 diff_1698000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1335 diff_1737000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1336 diff_1757000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1337 diff_1795000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1338 diff_1815000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1339 diff_1944000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=17000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1340 diff_1964000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1341 diff_2002000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1342 diff_2022000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1343 diff_2061000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=17000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1344 diff_2081000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1345 diff_2119000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1346 diff_2139000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1347 diff_2218000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1348 diff_2238000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1349 diff_2276000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1350 diff_2296000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1351 diff_2335000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=17000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1352 diff_2355000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1353 diff_2394000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1354 diff_2414000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1355 diff_2483000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=17000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1356 diff_2503000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1357 diff_2541000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1358 diff_2561000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1359 diff_2600000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=17000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1360 diff_2620000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1361 diff_2659000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1362 diff_2679000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1363 diff_2757000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1364 diff_2777000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1365 diff_2815000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1366 diff_2835000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1367 diff_2874000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=17000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1368 diff_2894000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1369 diff_2933000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1370 diff_2953000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1371 diff_2992000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=17000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1372 diff_3012000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1373 diff_3051000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1374 diff_3071000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1375 diff_3110000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1376 diff_3130000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1377 diff_3169000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1378 diff_3189000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1379 diff_3266000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1380 diff_3286000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1381 diff_3324000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1382 diff_3344000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1383 diff_3383000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=17000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1384 diff_3403000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1385 diff_3442000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1386 diff_3462000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1387 diff_3501000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=17000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1388 diff_3521000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1389 diff_3560000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1390 diff_3580000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1391 diff_3619000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1392 diff_3639000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1393 diff_3678000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1394 diff_3698000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1395 diff_3776000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1396 diff_3796000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1397 diff_3834000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1398 diff_3854000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1399 diff_3893000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=17000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1400 diff_3913000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1401 diff_3952000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1402 diff_3972000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1403 diff_4011000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=17000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1404 diff_4031000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1405 diff_4070000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1406 diff_4090000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1407 diff_4129000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1408 diff_4149000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1409 diff_4188000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1410 diff_4208000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1411 diff_4288000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1412 diff_4307000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1413 diff_4346000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1414 diff_4366000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1415 diff_4405000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=17000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1416 diff_4425000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1417 diff_4464000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1418 diff_4484000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1419 diff_4523000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1420 diff_4543000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1421 diff_4582000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1422 diff_4602000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1423 diff_4730000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1424 diff_4750000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1425 diff_4788000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1426 diff_4808000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1427 diff_4847000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1428 diff_4867000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1429 diff_4906000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1430 diff_4926000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1431 diff_5004000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1432 diff_5024000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1433 diff_5062000_5621000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1434 diff_5082000_5587000# diff_474000_5143000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1435 diff_91000_5337000# diff_197000_5470000# diff_83000_3098000# GND efet w=232000 l=9000
+ ad=-1.99887e+09 pd=1.828e+06 as=0 ps=0 
M1436 diff_95000_5192000# diff_91000_5337000# diff_91000_5337000# GND efet w=43000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1437 diff_83000_3098000# diff_402000_4713000# diff_506000_5537000# GND efet w=140000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1438 diff_5501000_5678000# diff_5501000_5678000# diff_95000_5192000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M1439 diff_5501000_5678000# diff_5954000_5147000# diff_5700000_5646000# GND efet w=13000 l=11000
+ ad=0 pd=0 as=5.53e+08 ps=148000 
M1440 diff_5954000_5147000# diff_5954000_5147000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=1.221e+09 pd=316000 as=0 ps=0 
M1441 diff_5954000_5147000# diff_474000_5143000# diff_83000_3098000# GND efet w=64000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1442 diff_83000_3098000# diff_5700000_5646000# diff_5502000_5646000# GND efet w=101000 l=8000
+ ad=0 pd=0 as=-1.29497e+09 ps=624000 
M1443 diff_95000_5192000# diff_5502000_5646000# diff_5502000_5646000# GND efet w=13000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M1444 diff_5502000_5646000# diff_5502000_5646000# diff_5502000_5646000# GND efet w=500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1445 diff_5700000_5646000# diff_474000_5143000# diff_5972000_5632000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=-1.71397e+09 ps=528000 
M1446 diff_95000_5192000# diff_5972000_5632000# diff_5972000_5632000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M1447 diff_83000_3098000# diff_6062000_5632000# diff_5972000_5632000# GND efet w=115500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1448 diff_83000_3098000# diff_775000_5479000# diff_761000_5561000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1449 diff_83000_3098000# diff_775000_5479000# diff_894000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1450 diff_83000_3098000# diff_775000_5479000# diff_973000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1451 diff_83000_3098000# diff_775000_5479000# diff_1032000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1452 diff_83000_3098000# diff_775000_5479000# diff_1169000_5621000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1453 diff_83000_3098000# diff_775000_5479000# diff_1228000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1454 diff_83000_3098000# diff_775000_5479000# diff_1366000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1455 diff_83000_3098000# diff_775000_5479000# diff_1424000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1456 diff_83000_3098000# diff_775000_5479000# diff_1522000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1457 diff_83000_3098000# diff_775000_5479000# diff_1678000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1458 diff_83000_3098000# diff_775000_5479000# diff_2119000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1459 diff_83000_3098000# diff_775000_5479000# diff_2276000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1460 diff_83000_3098000# diff_775000_5479000# diff_2355000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1461 diff_83000_3098000# diff_775000_5479000# diff_2503000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1462 diff_83000_3098000# diff_775000_5479000# diff_2679000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1463 diff_83000_3098000# diff_775000_5479000# diff_2894000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1464 diff_83000_3098000# diff_775000_5479000# diff_3012000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1465 diff_83000_3098000# diff_775000_5479000# diff_3071000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1466 diff_83000_3098000# diff_775000_5479000# diff_3130000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1467 diff_83000_3098000# diff_775000_5479000# diff_3169000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1468 diff_83000_3098000# diff_775000_5479000# diff_3266000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1469 diff_83000_3098000# diff_775000_5479000# diff_3560000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1470 diff_83000_3098000# diff_775000_5479000# diff_3580000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1471 diff_83000_3098000# diff_775000_5479000# diff_3639000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1472 diff_83000_3098000# diff_775000_5479000# diff_3893000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1473 diff_83000_3098000# diff_775000_5479000# diff_3913000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1474 diff_83000_3098000# diff_775000_5479000# diff_4011000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1475 diff_83000_3098000# diff_775000_5479000# diff_4307000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1476 diff_83000_3098000# diff_775000_5479000# diff_4808000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1477 diff_83000_3098000# diff_775000_5479000# diff_5004000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1478 diff_83000_3098000# diff_88000_5400000# diff_91000_5337000# GND efet w=83000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1479 diff_83000_3098000# diff_88000_5400000# diff_91000_5337000# GND efet w=112000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1480 diff_91000_5337000# diff_197000_5470000# diff_83000_3098000# GND efet w=49500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1481 diff_91000_5337000# diff_88000_5400000# diff_83000_3098000# GND efet w=83000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1482 diff_402000_4713000# diff_402000_4713000# diff_95000_5192000# GND efet w=16000 l=12000
+ ad=5.68033e+08 pd=812000 as=0 ps=0 
M1483 diff_775000_5421000# diff_775000_5421000# diff_95000_5192000# GND efet w=14000 l=8000
+ ad=-1.99593e+09 pd=1.378e+06 as=0 ps=0 
M1484 diff_775000_5421000# diff_5252000_5062000# diff_83000_3098000# GND efet w=182000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1485 diff_775000_5421000# diff_5501000_5603000# diff_83000_3098000# GND efet w=189000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1486 diff_83000_3098000# diff_5502000_5571000# diff_5501000_5603000# GND efet w=101500 l=7500
+ ad=0 pd=0 as=-1.56097e+09 ps=708000 
M1487 diff_83000_3098000# diff_5252000_5062000# diff_775000_5390000# GND efet w=179500 l=8500
+ ad=0 pd=0 as=1.98103e+09 ps=954000 
M1488 diff_775000_5390000# diff_5502000_5571000# diff_83000_3098000# GND efet w=179000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1489 diff_95000_5192000# diff_775000_5390000# diff_775000_5390000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1490 diff_5501000_5603000# diff_5501000_5603000# diff_95000_5192000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M1491 diff_5501000_5603000# diff_5954000_5147000# diff_5700000_5571000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=5.4e+08 ps=146000 
M1492 diff_5972000_5632000# diff_6022000_5610000# diff_83000_3098000# GND efet w=101000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1493 diff_6174000_5604000# diff_72000_4515000# diff_6022000_5610000# GND efet w=20000 l=12000
+ ad=-1.65197e+09 pd=588000 as=3.35e+08 ps=88000 
M1494 diff_6174000_5604000# diff_6174000_5604000# diff_6174000_5604000# GND efet w=1000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M1495 diff_95000_5192000# diff_6174000_5604000# diff_6174000_5604000# GND efet w=12000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M1496 diff_6174000_5604000# diff_5619000_2893000# diff_83000_3098000# GND efet w=126000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1497 diff_83000_3098000# diff_5700000_5571000# diff_5502000_5571000# GND efet w=101000 l=8000
+ ad=0 pd=0 as=-1.29497e+09 ps=624000 
M1498 diff_95000_5192000# diff_5502000_5571000# diff_5502000_5571000# GND efet w=13000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M1499 diff_5502000_5571000# diff_5502000_5571000# diff_5502000_5571000# GND efet w=500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1500 diff_5700000_5571000# diff_474000_5143000# diff_5972000_5557000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=1.761e+09 ps=416000 
M1501 diff_95000_5192000# diff_5972000_5557000# diff_5972000_5557000# GND efet w=13000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M1502 diff_83000_3098000# diff_5619000_2172000# diff_6194000_5553000# GND efet w=128000 l=10000
+ ad=0 pd=0 as=-1.85397e+09 ps=544000 
M1503 diff_797000_5587000# diff_775000_5448000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1504 diff_1464000_5621000# diff_775000_5448000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1505 diff_1698000_5587000# diff_775000_5448000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1506 diff_2061000_5621000# diff_775000_5448000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1507 diff_2874000_5621000# diff_775000_5448000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1508 diff_3189000_5587000# diff_775000_5448000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1509 diff_3324000_5621000# diff_775000_5448000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1510 diff_3344000_5587000# diff_775000_5448000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1511 diff_3678000_5621000# diff_775000_5448000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1512 diff_3796000_5587000# diff_775000_5448000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1513 diff_3834000_5621000# diff_775000_5448000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1514 diff_4031000_5587000# diff_775000_5448000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1515 diff_4070000_5621000# diff_775000_5448000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1516 diff_4129000_5621000# diff_775000_5448000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1517 diff_4208000_5587000# diff_775000_5448000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1518 diff_4484000_5587000# diff_775000_5448000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1519 diff_83000_3098000# diff_94000_3551000# diff_402000_4713000# GND efet w=77000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1520 diff_91000_5337000# diff_88000_5400000# diff_83000_3098000# GND efet w=99000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1521 diff_91000_5337000# diff_197000_5470000# diff_83000_3098000# GND efet w=51500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M1522 diff_6194000_5553000# diff_72000_4515000# diff_6016000_5535000# GND efet w=21000 l=12000
+ ad=0 pd=0 as=3.38e+08 ps=88000 
M1523 diff_6194000_5553000# diff_6062000_5632000# diff_83000_3098000# GND efet w=121500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1524 diff_83000_3098000# diff_6016000_5535000# diff_5972000_5557000# GND efet w=104000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1525 diff_402000_4713000# diff_94000_3551000# diff_83000_3098000# GND efet w=69000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1526 diff_775000_5364000# diff_775000_5364000# diff_95000_5192000# GND efet w=14000 l=9000
+ ad=2.02803e+09 pd=1.372e+06 as=0 ps=0 
M1527 diff_775000_5364000# diff_5252000_5062000# diff_83000_3098000# GND efet w=182000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1528 diff_775000_5364000# diff_5501000_5528000# diff_83000_3098000# GND efet w=189000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1529 diff_83000_3098000# diff_775000_5421000# diff_761000_5561000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1530 diff_83000_3098000# diff_775000_5421000# diff_894000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1531 diff_83000_3098000# diff_775000_5421000# diff_1012000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1532 diff_83000_3098000# diff_775000_5421000# diff_1130000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1533 diff_83000_3098000# diff_775000_5421000# diff_1464000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1534 diff_83000_3098000# diff_775000_5421000# diff_1678000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1535 diff_83000_3098000# diff_775000_5421000# diff_1698000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1536 diff_83000_3098000# diff_775000_5421000# diff_2061000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1537 diff_83000_3098000# diff_775000_5421000# diff_2561000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1538 diff_83000_3098000# diff_775000_5421000# diff_2777000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1539 diff_83000_3098000# diff_775000_5421000# diff_2835000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1540 diff_83000_3098000# diff_775000_5421000# diff_2874000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1541 diff_83000_3098000# diff_775000_5421000# diff_2894000_5587000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1542 diff_83000_3098000# diff_775000_5421000# diff_2933000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1543 diff_83000_3098000# diff_775000_5421000# diff_3012000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1544 diff_83000_3098000# diff_775000_5421000# diff_3051000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1545 diff_83000_3098000# diff_775000_5421000# diff_3071000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1546 diff_83000_3098000# diff_775000_5421000# diff_3130000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1547 diff_83000_3098000# diff_775000_5421000# diff_3324000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1548 diff_83000_3098000# diff_775000_5421000# diff_3560000_5621000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1549 diff_83000_3098000# diff_775000_5421000# diff_3580000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1550 diff_83000_3098000# diff_775000_5421000# diff_3639000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1551 diff_83000_3098000# diff_775000_5421000# diff_3678000_5621000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1552 diff_83000_3098000# diff_775000_5421000# diff_3698000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1553 diff_83000_3098000# diff_775000_5421000# diff_3834000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1554 diff_83000_3098000# diff_775000_5421000# diff_3893000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1555 diff_83000_3098000# diff_775000_5421000# diff_3952000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1556 diff_83000_3098000# diff_775000_5421000# diff_4011000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1557 diff_83000_3098000# diff_775000_5421000# diff_4031000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1558 diff_83000_3098000# diff_775000_5421000# diff_4070000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1559 diff_83000_3098000# diff_775000_5421000# diff_4129000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1560 diff_83000_3098000# diff_775000_5421000# diff_4582000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1561 diff_83000_3098000# diff_775000_5421000# diff_4847000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1562 diff_83000_3098000# diff_775000_5421000# diff_4867000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1563 diff_83000_3098000# diff_775000_5421000# diff_4906000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1564 diff_83000_3098000# diff_775000_5421000# diff_5082000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1565 diff_83000_3098000# diff_197000_5470000# diff_402000_4713000# GND efet w=130000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1566 diff_83000_3098000# diff_5502000_5496000# diff_5501000_5528000# GND efet w=101000 l=7000
+ ad=0 pd=0 as=-1.46097e+09 ps=708000 
M1567 diff_83000_3098000# diff_5252000_5062000# diff_775000_5333000# GND efet w=179500 l=8500
+ ad=0 pd=0 as=1.95703e+09 ps=956000 
M1568 diff_775000_5333000# diff_5502000_5496000# diff_83000_3098000# GND efet w=179000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1569 diff_95000_5192000# diff_775000_5333000# diff_775000_5333000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1570 diff_5501000_5528000# diff_5501000_5528000# diff_95000_5192000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M1571 diff_5501000_5528000# diff_5954000_5147000# diff_5700000_5496000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=5.7e+08 ps=144000 
M1572 diff_83000_3098000# diff_6017000_5510000# diff_5972000_5482000# GND efet w=103000 l=9000
+ ad=0 pd=0 as=2.063e+09 ps=426000 
M1573 diff_83000_3098000# diff_5700000_5496000# diff_5502000_5496000# GND efet w=101000 l=8000
+ ad=0 pd=0 as=-1.06397e+09 ps=626000 
M1574 diff_95000_5192000# diff_5502000_5496000# diff_5502000_5496000# GND efet w=13000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M1575 diff_5502000_5496000# diff_5502000_5496000# diff_5502000_5496000# GND efet w=500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1576 diff_5700000_5496000# diff_474000_5143000# diff_5972000_5482000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1577 diff_5972000_5482000# diff_5972000_5482000# diff_95000_5192000# GND efet w=12000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M1578 diff_6194000_5553000# diff_6194000_5553000# diff_95000_5192000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1579 diff_6194000_5481000# diff_72000_4515000# diff_6017000_5510000# GND efet w=19000 l=12000
+ ad=-1.83897e+09 pd=536000 as=2.97e+08 ps=84000 
M1580 diff_95000_5192000# diff_6194000_5481000# diff_6194000_5481000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1581 diff_83000_3098000# diff_6062000_5632000# diff_6194000_5481000# GND efet w=122000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1582 diff_83000_3098000# diff_75000_5299000# diff_91000_5337000# GND efet w=223500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1583 diff_953000_5621000# diff_775000_5390000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1584 diff_1032000_5587000# diff_775000_5390000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1585 diff_1110000_5621000# diff_775000_5390000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1586 diff_1169000_5621000# diff_775000_5390000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1587 diff_1366000_5587000# diff_775000_5390000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1588 diff_1424000_5587000# diff_775000_5390000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1589 diff_1522000_5621000# diff_775000_5390000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1590 diff_1757000_5587000# diff_775000_5390000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1591 diff_2119000_5621000# diff_775000_5390000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1592 diff_2139000_5587000# diff_775000_5390000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1593 diff_2276000_5621000# diff_775000_5390000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1594 diff_2355000_5587000# diff_775000_5390000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1595 diff_2483000_5621000# diff_775000_5390000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1596 diff_2503000_5587000# diff_775000_5390000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1597 diff_2620000_5587000# diff_775000_5390000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1598 diff_2659000_5621000# diff_775000_5390000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1599 diff_3189000_5587000# diff_775000_5390000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1600 diff_3266000_5621000# diff_775000_5390000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1601 diff_3286000_5587000# diff_775000_5390000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1602 diff_3344000_5587000# diff_775000_5390000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1603 diff_3383000_5621000# diff_775000_5390000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1604 diff_3796000_5587000# diff_775000_5390000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1605 diff_3913000_5587000# diff_775000_5390000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1606 diff_4149000_5587000# diff_775000_5390000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1607 diff_4208000_5587000# diff_775000_5390000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1608 diff_4288000_5621000# diff_775000_5390000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1609 diff_4523000_5621000# diff_775000_5390000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1610 diff_4730000_5621000# diff_775000_5390000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1611 diff_4926000_5587000# diff_775000_5390000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1612 diff_402000_4713000# diff_473000_5333000# diff_83000_3098000# GND efet w=155500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1613 diff_83000_3098000# diff_197000_5470000# diff_91000_5337000# GND efet w=49500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1614 diff_83000_3098000# diff_775000_5364000# diff_761000_5561000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1615 diff_83000_3098000# diff_775000_5364000# diff_797000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1616 diff_83000_3098000# diff_775000_5364000# diff_894000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1617 diff_83000_3098000# diff_775000_5364000# diff_914000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1618 diff_83000_3098000# diff_775000_5364000# diff_1032000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1619 diff_83000_3098000# diff_775000_5364000# diff_1130000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1620 diff_83000_3098000# diff_775000_5364000# diff_1169000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1621 diff_83000_3098000# diff_775000_5364000# diff_1366000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1622 diff_83000_3098000# diff_775000_5364000# diff_1424000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1623 diff_83000_3098000# diff_775000_5364000# diff_1464000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1624 diff_83000_3098000# diff_775000_5364000# diff_1522000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1625 diff_83000_3098000# diff_775000_5364000# diff_1678000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1626 diff_83000_3098000# diff_775000_5364000# diff_1698000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1627 diff_83000_3098000# diff_775000_5364000# diff_2061000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1628 diff_83000_3098000# diff_775000_5364000# diff_2119000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1629 diff_83000_3098000# diff_775000_5364000# diff_2238000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1630 diff_83000_3098000# diff_775000_5364000# diff_2276000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1631 diff_83000_3098000# diff_775000_5364000# diff_2335000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1632 diff_83000_3098000# diff_775000_5364000# diff_2503000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1633 diff_83000_3098000# diff_775000_5364000# diff_2561000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1634 diff_83000_3098000# diff_775000_5364000# diff_2600000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1635 diff_83000_3098000# diff_775000_5364000# diff_2679000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1636 diff_83000_3098000# diff_775000_5364000# diff_2777000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1637 diff_83000_3098000# diff_775000_5364000# diff_2815000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1638 diff_83000_3098000# diff_775000_5364000# diff_2835000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1639 diff_83000_3098000# diff_775000_5364000# diff_2874000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1640 diff_83000_3098000# diff_775000_5364000# diff_2933000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1641 diff_83000_3098000# diff_775000_5364000# diff_2953000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1642 diff_83000_3098000# diff_775000_5364000# diff_3012000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1643 diff_83000_3098000# diff_775000_5364000# diff_3051000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1644 diff_83000_3098000# diff_775000_5364000# diff_3071000_5587000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1645 diff_83000_3098000# diff_775000_5364000# diff_3130000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1646 diff_83000_3098000# diff_775000_5364000# diff_3189000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1647 diff_83000_3098000# diff_775000_5364000# diff_3462000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1648 diff_83000_3098000# diff_775000_5364000# diff_3501000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1649 diff_83000_3098000# diff_775000_5364000# diff_3560000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1650 diff_83000_3098000# diff_775000_5364000# diff_3580000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1651 diff_83000_3098000# diff_775000_5364000# diff_3639000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1652 diff_83000_3098000# diff_775000_5364000# diff_3678000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1653 diff_83000_3098000# diff_775000_5364000# diff_3698000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1654 diff_83000_3098000# diff_775000_5364000# diff_3796000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1655 diff_83000_3098000# diff_775000_5364000# diff_3834000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1656 diff_83000_3098000# diff_775000_5364000# diff_3952000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1657 diff_83000_3098000# diff_775000_5364000# diff_4011000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1658 diff_83000_3098000# diff_775000_5364000# diff_4031000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1659 diff_83000_3098000# diff_775000_5364000# diff_4070000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1660 diff_83000_3098000# diff_775000_5364000# diff_4208000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1661 diff_83000_3098000# diff_775000_5364000# diff_4405000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1662 diff_83000_3098000# diff_775000_5364000# diff_4425000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1663 diff_83000_3098000# diff_775000_5364000# diff_4543000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1664 diff_83000_3098000# diff_775000_5364000# diff_4582000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1665 diff_83000_3098000# diff_775000_5364000# diff_4602000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1666 diff_83000_3098000# diff_775000_5364000# diff_4750000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1667 diff_83000_3098000# diff_775000_5364000# diff_4867000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1668 diff_83000_3098000# diff_775000_5364000# diff_4926000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1669 diff_83000_3098000# diff_775000_5364000# diff_5062000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1670 diff_775000_5306000# diff_775000_5306000# diff_95000_5192000# GND efet w=14000 l=9000
+ ad=-1.69493e+09 pd=1.464e+06 as=0 ps=0 
M1671 diff_775000_5306000# diff_5252000_5062000# diff_83000_3098000# GND efet w=182000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1672 diff_775000_5306000# diff_5501000_5453000# diff_83000_3098000# GND efet w=187500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1673 diff_83000_3098000# diff_5502000_5421000# diff_5501000_5453000# GND efet w=101000 l=7000
+ ad=0 pd=0 as=-1.33097e+09 ps=704000 
M1674 diff_83000_3098000# diff_5252000_5062000# diff_775000_5275000# GND efet w=178000 l=8000
+ ad=0 pd=0 as=1.89903e+09 ps=950000 
M1675 diff_83000_3098000# diff_5502000_5421000# diff_775000_5275000# GND efet w=177500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1676 diff_91000_5337000# diff_75000_5299000# diff_83000_3098000# GND efet w=187000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1677 diff_91000_5337000# diff_197000_5470000# diff_83000_3098000# GND efet w=49500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1678 diff_83000_3098000# diff_493000_5343000# diff_499000_5334000# GND efet w=138000 l=8000
+ ad=0 pd=0 as=1.732e+09 ps=382000 
M1679 diff_95000_5192000# diff_775000_5275000# diff_775000_5275000# GND efet w=14000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1680 diff_5501000_5453000# diff_5501000_5453000# diff_95000_5192000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M1681 diff_5501000_5453000# diff_5954000_5147000# diff_5700000_5421000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=5.7e+08 ps=144000 
M1682 diff_6194000_5481000# diff_5619000_2102000# diff_83000_3098000# GND efet w=130000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1683 diff_95000_5192000# diff_5972000_5406000# diff_5972000_5406000# GND efet w=12000 l=16000
+ ad=0 pd=0 as=1.857e+09 ps=454000 
M1684 diff_83000_3098000# diff_5700000_5421000# diff_5502000_5421000# GND efet w=101000 l=9000
+ ad=0 pd=0 as=-1.16597e+09 ps=624000 
M1685 diff_95000_5192000# diff_5502000_5421000# diff_5502000_5421000# GND efet w=13000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M1686 diff_83000_3098000# diff_5619000_1381000# diff_6170000_5416000# GND efet w=130000 l=10000
+ ad=0 pd=0 as=-1.49497e+09 ps=584000 
M1687 diff_83000_3098000# diff_6017000_5422000# diff_5972000_5406000# GND efet w=104500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1688 diff_5502000_5421000# diff_5502000_5421000# diff_5502000_5421000# GND efet w=500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1689 diff_5700000_5421000# diff_474000_5143000# diff_5972000_5406000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1690 diff_6170000_5416000# diff_72000_4515000# diff_6017000_5422000# GND efet w=21000 l=12000
+ ad=0 pd=0 as=3.25e+08 ps=90000 
M1691 diff_83000_3098000# diff_6062000_5632000# diff_6170000_5416000# GND efet w=121500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M1692 diff_75000_5299000# diff_68000_5288000# diff_64000_4639000# GND efet w=28000 l=11000
+ ad=3.61e+08 pd=104000 as=9.62033e+08 ps=824000 
M1693 diff_473000_5333000# diff_68000_5288000# diff_465000_5280000# GND efet w=11000 l=11000
+ ad=1.94e+08 pd=88000 as=-1.56897e+09 ps=398000 
M1694 diff_499000_5334000# diff_502000_5322000# diff_465000_5280000# GND efet w=147500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1695 diff_465000_5280000# diff_465000_5280000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M1696 diff_95000_5192000# diff_85000_5213000# diff_95000_5160000# GND efet w=234500 l=7500
+ ad=0 pd=0 as=8.93229e+08 ps=3.008e+06 
M1697 diff_502000_5322000# diff_72000_4515000# diff_100000_3992000# GND efet w=13000 l=11000
+ ad=2.44e+08 pd=94000 as=-5.63967e+08 ps=784000 
M1698 diff_953000_5621000# diff_775000_5333000# diff_83000_3098000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1699 diff_973000_5587000# diff_775000_5333000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1700 diff_1012000_5621000# diff_775000_5333000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1701 diff_1757000_5587000# diff_775000_5333000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1702 diff_2139000_5587000# diff_775000_5333000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1703 diff_2355000_5587000# diff_775000_5333000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1704 diff_2483000_5621000# diff_775000_5333000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1705 diff_2620000_5587000# diff_775000_5333000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1706 diff_2659000_5621000# diff_775000_5333000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1707 diff_2757000_5621000# diff_775000_5333000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1708 diff_2894000_5587000# diff_775000_5333000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1709 diff_3169000_5621000# diff_775000_5333000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1710 diff_3266000_5621000# diff_775000_5333000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1711 diff_3286000_5587000# diff_775000_5333000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1712 diff_3324000_5621000# diff_775000_5333000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1713 diff_3344000_5587000# diff_775000_5333000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1714 diff_3383000_5621000# diff_775000_5333000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1715 diff_3893000_5621000# diff_775000_5333000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1716 diff_4129000_5621000# diff_775000_5333000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1717 diff_4149000_5587000# diff_775000_5333000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1718 diff_4188000_5621000# diff_775000_5333000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1719 diff_4288000_5621000# diff_775000_5333000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1720 diff_4366000_5587000# diff_775000_5333000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1721 diff_4484000_5587000# diff_775000_5333000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1722 diff_4523000_5621000# diff_775000_5333000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1723 diff_4730000_5621000# diff_775000_5333000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1724 diff_4808000_5587000# diff_775000_5333000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1725 diff_4847000_5621000# diff_775000_5333000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1726 diff_4906000_5621000# diff_775000_5333000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1727 diff_83000_3098000# diff_775000_5306000# diff_797000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1728 diff_83000_3098000# diff_775000_5306000# diff_914000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1729 diff_83000_3098000# diff_775000_5306000# diff_953000_5621000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1730 diff_83000_3098000# diff_775000_5306000# diff_973000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1731 diff_83000_3098000# diff_775000_5306000# diff_1032000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1732 diff_83000_3098000# diff_775000_5306000# diff_1169000_5621000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1733 diff_83000_3098000# diff_775000_5306000# diff_1366000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1734 diff_83000_3098000# diff_775000_5306000# diff_1424000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1735 diff_83000_3098000# diff_775000_5306000# diff_1464000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1736 diff_83000_3098000# diff_775000_5306000# diff_1522000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1737 diff_83000_3098000# diff_775000_5306000# diff_1698000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1738 diff_83000_3098000# diff_775000_5306000# diff_1757000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1739 diff_83000_3098000# diff_775000_5306000# diff_2061000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1740 diff_83000_3098000# diff_775000_5306000# diff_2119000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1741 diff_83000_3098000# diff_775000_5306000# diff_2139000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1742 diff_83000_3098000# diff_775000_5306000# diff_2238000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1743 diff_83000_3098000# diff_775000_5306000# diff_2276000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1744 diff_83000_3098000# diff_775000_5306000# diff_2355000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1745 diff_83000_3098000# diff_775000_5306000# diff_2483000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1746 diff_83000_3098000# diff_775000_5306000# diff_2561000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1747 diff_83000_3098000# diff_775000_5306000# diff_2600000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1748 diff_83000_3098000# diff_775000_5306000# diff_2620000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1749 diff_83000_3098000# diff_775000_5306000# diff_2659000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1750 diff_83000_3098000# diff_775000_5306000# diff_2679000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1751 diff_83000_3098000# diff_775000_5306000# diff_2757000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1752 diff_83000_3098000# diff_775000_5306000# diff_2815000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1753 diff_83000_3098000# diff_775000_5306000# diff_2835000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1754 diff_83000_3098000# diff_775000_5306000# diff_2894000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1755 diff_83000_3098000# diff_775000_5306000# diff_2933000_5621000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1756 diff_83000_3098000# diff_775000_5306000# diff_2953000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1757 diff_83000_3098000# diff_775000_5306000# diff_3012000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1758 diff_83000_3098000# diff_775000_5306000# diff_3169000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1759 diff_83000_3098000# diff_775000_5306000# diff_3189000_5587000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1760 diff_83000_3098000# diff_775000_5306000# diff_3266000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1761 diff_83000_3098000# diff_775000_5306000# diff_3383000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1762 diff_83000_3098000# diff_775000_5306000# diff_3462000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1763 diff_83000_3098000# diff_775000_5306000# diff_3639000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1764 diff_83000_3098000# diff_775000_5306000# diff_3678000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1765 diff_83000_3098000# diff_775000_5306000# diff_3796000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1766 diff_83000_3098000# diff_775000_5306000# diff_4149000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1767 diff_83000_3098000# diff_775000_5306000# diff_4208000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1768 diff_83000_3098000# diff_775000_5306000# diff_4288000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1769 diff_83000_3098000# diff_775000_5306000# diff_4307000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1770 diff_83000_3098000# diff_775000_5306000# diff_4405000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1771 diff_83000_3098000# diff_775000_5306000# diff_4425000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1772 diff_83000_3098000# diff_775000_5306000# diff_4484000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1773 diff_83000_3098000# diff_775000_5306000# diff_4523000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1774 diff_83000_3098000# diff_775000_5306000# diff_4582000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1775 diff_83000_3098000# diff_775000_5306000# diff_4730000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1776 diff_83000_3098000# diff_775000_5306000# diff_4808000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1777 diff_83000_3098000# diff_775000_5306000# diff_4847000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1778 diff_83000_3098000# diff_775000_5306000# diff_4867000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1779 diff_83000_3098000# diff_775000_5306000# diff_4906000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1780 diff_83000_3098000# diff_775000_5306000# diff_4926000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1781 diff_83000_3098000# diff_775000_5306000# diff_5024000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1782 diff_775000_5249000# diff_775000_5249000# diff_95000_5192000# GND efet w=14000 l=8000
+ ad=1.83803e+09 pd=1.32e+06 as=0 ps=0 
M1783 diff_775000_5249000# diff_5252000_5062000# diff_83000_3098000# GND efet w=180500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1784 diff_775000_5249000# diff_5501000_5377000# diff_83000_3098000# GND efet w=188500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1785 diff_83000_3098000# diff_5502000_5346000# diff_5501000_5377000# GND efet w=101000 l=8000
+ ad=0 pd=0 as=-1.63397e+09 ps=670000 
M1786 diff_83000_3098000# diff_5252000_5062000# diff_775000_5218000# GND efet w=178500 l=8500
+ ad=0 pd=0 as=1.78303e+09 ps=952000 
M1787 diff_83000_3098000# diff_5502000_5346000# diff_775000_5218000# GND efet w=179000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1788 diff_95000_5192000# diff_775000_5218000# diff_775000_5218000# GND efet w=13000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1789 diff_5501000_5377000# diff_5501000_5377000# diff_95000_5192000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M1790 diff_5501000_5377000# diff_5954000_5147000# diff_5700000_5345000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=5.59e+08 ps=146000 
M1791 diff_6170000_5416000# diff_6170000_5416000# diff_95000_5192000# GND efet w=13000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M1792 diff_83000_3098000# diff_6012000_5360000# diff_5972000_5331000# GND efet w=104000 l=8000
+ ad=0 pd=0 as=2.142e+09 ps=420000 
M1793 diff_761000_5561000# diff_775000_5275000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1794 diff_835000_5621000# diff_775000_5275000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1795 diff_894000_5621000# diff_775000_5275000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1796 diff_1012000_5621000# diff_775000_5275000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1797 diff_1110000_5621000# diff_775000_5275000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1798 diff_1130000_5587000# diff_775000_5275000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1799 diff_2503000_5587000# diff_775000_5275000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1800 diff_2874000_5621000# diff_775000_5275000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1801 diff_3051000_5621000# diff_775000_5275000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1802 diff_3130000_5587000# diff_775000_5275000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1803 diff_3286000_5587000# diff_775000_5275000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1804 diff_3324000_5621000# diff_775000_5275000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1805 diff_3344000_5587000# diff_775000_5275000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1806 diff_3521000_5587000# diff_775000_5275000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1807 diff_3560000_5621000# diff_775000_5275000# diff_83000_3098000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1808 diff_3580000_5587000# diff_775000_5275000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1809 diff_3834000_5621000# diff_775000_5275000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1810 diff_3893000_5621000# diff_775000_5275000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1811 diff_3913000_5587000# diff_775000_5275000# diff_83000_3098000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1812 diff_3952000_5621000# diff_775000_5275000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1813 diff_4011000_5621000# diff_775000_5275000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1814 diff_4031000_5587000# diff_775000_5275000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1815 diff_4070000_5621000# diff_775000_5275000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1816 diff_4129000_5621000# diff_775000_5275000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1817 diff_4188000_5621000# diff_775000_5275000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1818 diff_4366000_5587000# diff_775000_5275000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1819 diff_4543000_5587000# diff_775000_5275000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1820 diff_4602000_5587000# diff_775000_5275000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1821 diff_4750000_5587000# diff_775000_5275000# diff_83000_3098000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1822 diff_83000_3098000# diff_5700000_5345000# diff_5502000_5346000# GND efet w=101000 l=9000
+ ad=0 pd=0 as=-1.16697e+09 ps=624000 
M1823 diff_95000_5192000# diff_5502000_5346000# diff_5502000_5346000# GND efet w=13000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M1824 diff_5502000_5346000# diff_5502000_5346000# diff_5502000_5346000# GND efet w=500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1825 diff_5700000_5345000# diff_474000_5143000# diff_5972000_5331000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1826 diff_5972000_5331000# diff_5972000_5331000# diff_95000_5192000# GND efet w=12000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M1827 diff_6170000_5342000# diff_72000_4515000# diff_6012000_5360000# GND efet w=22000 l=12000
+ ad=-1.55897e+09 pd=592000 as=3.49e+08 ps=92000 
M1828 diff_95000_5192000# diff_6170000_5342000# diff_6170000_5342000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1829 diff_83000_3098000# diff_6062000_5632000# diff_6170000_5342000# GND efet w=122000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1830 diff_83000_3098000# diff_5619000_1309000# diff_6170000_5342000# GND efet w=128000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1831 diff_493000_5343000# diff_72000_4515000# diff_514000_5204000# GND efet w=11000 l=12000
+ ad=3.5e+08 pd=104000 as=1.632e+09 ps=318000 
M1832 diff_83000_3098000# diff_775000_5249000# diff_1188000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1833 diff_83000_3098000# diff_775000_5249000# diff_1248000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1834 diff_83000_3098000# diff_775000_5249000# diff_1286000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1835 diff_83000_3098000# diff_775000_5249000# diff_1306000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1836 diff_83000_3098000# diff_775000_5249000# diff_1346000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1837 diff_83000_3098000# diff_775000_5249000# diff_1795000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1838 diff_83000_3098000# diff_775000_5249000# diff_1944000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1839 diff_83000_3098000# diff_775000_5249000# diff_2335000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1840 diff_83000_3098000# diff_775000_5249000# diff_2394000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1841 diff_83000_3098000# diff_775000_5249000# diff_2503000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1842 diff_83000_3098000# diff_775000_5249000# diff_2620000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1843 diff_83000_3098000# diff_775000_5249000# diff_2894000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1844 diff_83000_3098000# diff_775000_5249000# diff_3051000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1845 diff_83000_3098000# diff_775000_5249000# diff_3442000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1846 diff_83000_3098000# diff_775000_5249000# diff_3560000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1847 diff_83000_3098000# diff_775000_5249000# diff_3619000_5621000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1848 diff_83000_3098000# diff_775000_5249000# diff_3834000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1849 diff_83000_3098000# diff_775000_5249000# diff_3854000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1850 diff_83000_3098000# diff_775000_5249000# diff_4070000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1851 diff_83000_3098000# diff_775000_5249000# diff_4149000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1852 diff_83000_3098000# diff_775000_5249000# diff_4847000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1853 diff_775000_5192000# diff_775000_5192000# diff_95000_5192000# GND efet w=14000 l=8000
+ ad=1.49203e+09 pd=1.218e+06 as=0 ps=0 
M1854 diff_775000_5192000# diff_5252000_5062000# diff_83000_3098000# GND efet w=180500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1855 diff_95000_5160000# diff_85000_5213000# diff_95000_5192000# GND efet w=241000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1856 diff_514000_5204000# diff_514000_5204000# diff_95000_5192000# GND efet w=13000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M1857 diff_83000_3098000# diff_197000_5470000# diff_514000_5204000# GND efet w=82000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1858 diff_95000_5192000# diff_85000_5213000# diff_95000_5160000# GND efet w=241000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1859 diff_83000_3098000# diff_77000_4827000# diff_95000_5160000# GND efet w=220000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1860 diff_95000_5160000# diff_77000_4827000# diff_83000_3098000# GND efet w=220000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1861 diff_83000_3098000# diff_77000_4827000# diff_95000_5160000# GND efet w=220000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1862 diff_95000_5160000# diff_77000_4827000# diff_83000_3098000# GND efet w=220000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1863 diff_83000_3098000# diff_77000_4827000# diff_95000_5160000# GND efet w=220000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1864 diff_95000_5160000# diff_77000_4827000# diff_83000_3098000# GND efet w=220000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1865 diff_83000_3098000# diff_77000_4827000# diff_85000_5213000# GND efet w=252500 l=8500
+ ad=0 pd=0 as=-5.04967e+08 ps=552000 
M1866 diff_95000_5192000# diff_85000_5213000# diff_95000_5160000# GND efet w=269500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1867 diff_474000_5143000# diff_465000_5069000# diff_83000_3098000# GND efet w=193000 l=8000
+ ad=6.55033e+08 pd=814000 as=0 ps=0 
M1868 diff_474000_5143000# diff_465000_5069000# diff_83000_3098000# GND efet w=162000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M1869 diff_83000_3098000# diff_487000_5098000# diff_465000_5069000# GND efet w=130000 l=9000
+ ad=0 pd=0 as=-2.07097e+09 ps=356000 
M1870 diff_465000_5069000# diff_465000_5069000# diff_95000_5192000# GND efet w=12000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1871 diff_95000_5192000# diff_487000_5098000# diff_474000_5143000# GND efet w=145000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1872 diff_775000_5192000# diff_5501000_5302000# diff_83000_3098000# GND efet w=187500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1873 diff_83000_3098000# diff_5502000_5270000# diff_5501000_5302000# GND efet w=101000 l=8000
+ ad=0 pd=0 as=-1.63297e+09 ps=672000 
M1874 diff_83000_3098000# diff_5252000_5062000# diff_775000_5160000# GND efet w=178500 l=8500
+ ad=0 pd=0 as=1.67603e+09 ps=942000 
M1875 diff_775000_5160000# diff_5502000_5270000# diff_83000_3098000# GND efet w=178500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1876 diff_5501000_5302000# diff_5501000_5302000# diff_95000_5192000# GND efet w=12000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M1877 diff_95000_5192000# diff_775000_5160000# diff_775000_5160000# GND efet w=13000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1878 diff_953000_5621000# diff_775000_5218000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1879 diff_1169000_5621000# diff_775000_5218000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1880 diff_1404000_5621000# diff_775000_5218000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1881 diff_1484000_5587000# diff_775000_5218000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1882 diff_1522000_5621000# diff_775000_5218000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1883 diff_1639000_5587000# diff_775000_5218000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1884 diff_1757000_5587000# diff_775000_5218000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1885 diff_1815000_5587000# diff_775000_5218000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1886 diff_1964000_5587000# diff_775000_5218000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1887 diff_2022000_5587000# diff_775000_5218000# diff_83000_3098000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1888 diff_2081000_5587000# diff_775000_5218000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1889 diff_2139000_5587000# diff_775000_5218000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1890 diff_2276000_5621000# diff_775000_5218000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1891 diff_2296000_5587000# diff_775000_5218000# diff_83000_3098000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1892 diff_2355000_5587000# diff_775000_5218000# diff_83000_3098000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1893 diff_2414000_5587000# diff_775000_5218000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1894 diff_2483000_5621000# diff_775000_5218000# diff_83000_3098000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1895 diff_2541000_5621000# diff_775000_5218000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1896 diff_2874000_5621000# diff_775000_5218000# diff_83000_3098000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1897 diff_3130000_5587000# diff_775000_5218000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1898 diff_3383000_5621000# diff_775000_5218000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1899 diff_3952000_5621000# diff_775000_5218000# diff_83000_3098000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1900 diff_3972000_5587000# diff_775000_5218000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1901 diff_4346000_5621000# diff_775000_5218000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1902 diff_4788000_5621000# diff_775000_5218000# diff_83000_3098000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1903 diff_4867000_5587000# diff_775000_5218000# diff_83000_3098000# GND efet w=18000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1904 diff_4906000_5621000# diff_775000_5218000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1905 diff_4926000_5587000# diff_775000_5218000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1906 diff_83000_3098000# diff_5700000_5270000# diff_5502000_5270000# GND efet w=101000 l=9000
+ ad=0 pd=0 as=-1.26797e+09 ps=628000 
M1907 diff_5501000_5302000# diff_5954000_5147000# diff_5700000_5270000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=5.53e+08 ps=146000 
M1908 diff_95000_5192000# diff_5972000_5256000# diff_5972000_5256000# GND efet w=12000 l=15000
+ ad=0 pd=0 as=1.813e+09 ps=440000 
M1909 diff_95000_5192000# diff_5502000_5270000# diff_5502000_5270000# GND efet w=13000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M1910 diff_83000_3098000# diff_6012000_5272000# diff_5972000_5256000# GND efet w=103000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1911 diff_5502000_5270000# diff_5502000_5270000# diff_5502000_5270000# GND efet w=500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1912 diff_5700000_5270000# diff_474000_5143000# diff_5972000_5256000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1913 diff_6170000_5282000# diff_72000_4515000# diff_6012000_5272000# GND efet w=21000 l=11000
+ ad=-8.17967e+08 pd=660000 as=3.56e+08 ps=92000 
M1914 diff_83000_3098000# diff_775000_5192000# diff_1032000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1915 diff_83000_3098000# diff_775000_5192000# diff_1188000_5587000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1916 diff_83000_3098000# diff_775000_5192000# diff_1248000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1917 diff_83000_3098000# diff_775000_5192000# diff_1404000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1918 diff_83000_3098000# diff_775000_5192000# diff_1484000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1919 diff_83000_3098000# diff_775000_5192000# diff_1619000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1920 diff_83000_3098000# diff_775000_5192000# diff_1698000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1921 diff_83000_3098000# diff_775000_5192000# diff_1815000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1922 diff_83000_3098000# diff_775000_5192000# diff_1944000_5621000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1923 diff_83000_3098000# diff_775000_5192000# diff_2081000_5587000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1924 diff_83000_3098000# diff_775000_5192000# diff_2218000_5621000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1925 diff_83000_3098000# diff_775000_5192000# diff_2296000_5587000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1926 diff_83000_3098000# diff_775000_5192000# diff_2335000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1927 diff_83000_3098000# diff_775000_5192000# diff_2394000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1928 diff_83000_3098000# diff_775000_5192000# diff_2414000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1929 diff_83000_3098000# diff_775000_5192000# diff_2503000_5587000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1930 diff_83000_3098000# diff_775000_5192000# diff_2541000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1931 diff_83000_3098000# diff_775000_5192000# diff_2620000_5587000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1932 diff_83000_3098000# diff_775000_5192000# diff_2894000_5587000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1933 diff_83000_3098000# diff_775000_5192000# diff_2992000_5621000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1934 diff_83000_3098000# diff_775000_5192000# diff_3051000_5621000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1935 diff_83000_3098000# diff_775000_5192000# diff_3560000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1936 diff_83000_3098000# diff_775000_5192000# diff_4070000_5621000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1937 diff_775000_5134000# diff_775000_5134000# diff_95000_5192000# GND efet w=14000 l=8000
+ ad=1.88303e+09 pd=1.282e+06 as=0 ps=0 
M1938 diff_775000_5134000# diff_5252000_5062000# diff_83000_3098000# GND efet w=180000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1939 diff_775000_5134000# diff_5501000_5227000# diff_83000_3098000# GND efet w=186500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1940 diff_83000_3098000# diff_5502000_5195000# diff_5501000_5227000# GND efet w=101000 l=8000
+ ad=0 pd=0 as=-1.63197e+09 ps=670000 
M1941 diff_953000_5621000# diff_775000_5160000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1942 diff_1286000_5621000# diff_775000_5160000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1943 diff_1306000_5587000# diff_775000_5160000# diff_83000_3098000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1944 diff_1522000_5621000# diff_775000_5160000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1945 diff_1737000_5621000# diff_775000_5160000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1946 diff_1757000_5587000# diff_775000_5160000# diff_83000_3098000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1947 diff_1795000_5621000# diff_775000_5160000# diff_83000_3098000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1948 diff_1964000_5587000# diff_775000_5160000# diff_83000_3098000# GND efet w=22000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1949 diff_2002000_5621000# diff_775000_5160000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1950 diff_2022000_5587000# diff_775000_5160000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1951 diff_2139000_5587000# diff_775000_5160000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1952 diff_2276000_5621000# diff_775000_5160000# diff_83000_3098000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1953 diff_2355000_5587000# diff_775000_5160000# diff_83000_3098000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1954 diff_2483000_5621000# diff_775000_5160000# diff_83000_3098000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1955 diff_2874000_5621000# diff_775000_5160000# diff_83000_3098000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1956 diff_3130000_5587000# diff_775000_5160000# diff_83000_3098000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1957 diff_3383000_5621000# diff_775000_5160000# diff_83000_3098000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1958 diff_3442000_5621000# diff_775000_5160000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1959 diff_3619000_5621000# diff_775000_5160000# diff_83000_3098000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1960 diff_3834000_5621000# diff_775000_5160000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1961 diff_3854000_5587000# diff_775000_5160000# diff_83000_3098000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1962 diff_3952000_5621000# diff_775000_5160000# diff_83000_3098000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1963 diff_3972000_5587000# diff_775000_5160000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1964 diff_4031000_5587000# diff_775000_5160000# diff_83000_3098000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1965 diff_4149000_5587000# diff_775000_5160000# diff_83000_3098000# GND efet w=22000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1966 diff_4346000_5621000# diff_775000_5160000# diff_83000_3098000# GND efet w=22000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1967 diff_4464000_5621000# diff_775000_5160000# diff_83000_3098000# GND efet w=22000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1968 diff_4788000_5621000# diff_775000_5160000# diff_83000_3098000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1969 diff_4847000_5621000# diff_775000_5160000# diff_83000_3098000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1970 diff_4867000_5587000# diff_775000_5160000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1971 diff_4906000_5621000# diff_775000_5160000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1972 diff_4926000_5587000# diff_775000_5160000# diff_83000_3098000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1973 diff_83000_3098000# diff_5252000_5062000# diff_775000_5103000# GND efet w=178000 l=9000
+ ad=0 pd=0 as=1.63303e+09 ps=952000 
M1974 diff_775000_5103000# diff_5502000_5195000# diff_83000_3098000# GND efet w=179000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1975 diff_5501000_5227000# diff_5501000_5227000# diff_95000_5192000# GND efet w=12000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M1976 diff_5501000_5227000# diff_5954000_5147000# diff_5700000_5195000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=5.42e+08 ps=146000 
M1977 diff_95000_5192000# diff_6170000_5282000# diff_6170000_5282000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1978 diff_83000_3098000# diff_5600000_575000# diff_6170000_5282000# GND efet w=127500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M1979 diff_95000_5192000# diff_775000_5103000# diff_775000_5103000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M1980 diff_83000_3098000# diff_5700000_5195000# diff_5502000_5195000# GND efet w=101000 l=9000
+ ad=0 pd=0 as=-1.28597e+09 ps=630000 
M1981 diff_83000_3098000# diff_6062000_5632000# diff_5972000_5181000# GND efet w=103000 l=8000
+ ad=0 pd=0 as=-1.95597e+09 ps=538000 
M1982 diff_83000_3098000# diff_6062000_5632000# diff_6170000_5282000# GND efet w=121000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1983 diff_95000_5192000# diff_5502000_5195000# diff_5502000_5195000# GND efet w=13000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M1984 diff_5502000_5195000# diff_5502000_5195000# diff_5502000_5195000# GND efet w=500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M1985 diff_5700000_5195000# diff_474000_5143000# diff_5972000_5181000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1986 diff_83000_3098000# diff_6074000_5195000# diff_5972000_5181000# GND efet w=104000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1987 diff_5972000_5181000# diff_5972000_5181000# diff_95000_5192000# GND efet w=12000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M1988 diff_6226000_5191000# diff_72000_4515000# diff_6074000_5195000# GND efet w=19000 l=11000
+ ad=-1.62897e+09 pd=576000 as=3.16e+08 ps=86000 
M1989 diff_83000_3098000# diff_775000_5134000# diff_1032000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1990 diff_83000_3098000# diff_775000_5134000# diff_1464000_5621000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1991 diff_83000_3098000# diff_775000_5134000# diff_1619000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1992 diff_83000_3098000# diff_775000_5134000# diff_1698000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1993 diff_83000_3098000# diff_775000_5134000# diff_2061000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1994 diff_83000_3098000# diff_775000_5134000# diff_2218000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1995 diff_83000_3098000# diff_775000_5134000# diff_2679000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1996 diff_83000_3098000# diff_775000_5134000# diff_2992000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1997 diff_83000_3098000# diff_775000_5134000# diff_3501000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1998 diff_83000_3098000# diff_775000_5134000# diff_3521000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1999 diff_83000_3098000# diff_775000_5134000# diff_3580000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2000 diff_83000_3098000# diff_775000_5134000# diff_3639000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2001 diff_83000_3098000# diff_775000_5134000# diff_3678000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2002 diff_83000_3098000# diff_775000_5134000# diff_3776000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2003 diff_83000_3098000# diff_775000_5134000# diff_3854000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2004 diff_83000_3098000# diff_775000_5134000# diff_3972000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2005 diff_83000_3098000# diff_775000_5134000# diff_4288000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2006 diff_83000_3098000# diff_775000_5134000# diff_4523000_5621000# GND efet w=22000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2007 diff_83000_3098000# diff_775000_5134000# diff_4602000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2008 diff_83000_3098000# diff_775000_5134000# diff_4730000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2009 diff_83000_3098000# diff_775000_5134000# diff_4750000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2010 diff_83000_3098000# diff_6074000_5171000# diff_5972000_5106000# GND efet w=104000 l=8000
+ ad=0 pd=0 as=-1.71397e+09 ps=580000 
M2011 diff_775000_5076000# diff_775000_5076000# diff_95000_5192000# GND efet w=14000 l=8000
+ ad=1.77603e+09 pd=1.226e+06 as=0 ps=0 
M2012 diff_775000_5076000# diff_5252000_5062000# diff_83000_3098000# GND efet w=180500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2013 diff_775000_5076000# diff_5501000_5152000# diff_83000_3098000# GND efet w=187500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2014 diff_83000_3098000# diff_5502000_5120000# diff_5501000_5152000# GND efet w=101000 l=8000
+ ad=0 pd=0 as=-1.62597e+09 ps=682000 
M2015 diff_953000_5621000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2016 diff_1248000_5587000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2017 diff_1404000_5621000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2018 diff_1757000_5587000# diff_775000_5103000# diff_83000_3098000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2019 diff_1815000_5587000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2020 diff_2081000_5587000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2021 diff_2139000_5587000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2022 diff_2296000_5587000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2023 diff_2335000_5621000# diff_775000_5103000# diff_83000_3098000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2024 diff_2355000_5587000# diff_775000_5103000# diff_83000_3098000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2025 diff_2483000_5621000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2026 diff_2503000_5587000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2027 diff_2620000_5587000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2028 diff_2835000_5587000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2029 diff_2874000_5621000# diff_775000_5103000# diff_83000_3098000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2030 diff_2894000_5587000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2031 diff_3051000_5621000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2032 diff_3110000_5621000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2033 diff_3130000_5587000# diff_775000_5103000# diff_83000_3098000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2034 diff_3383000_5621000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2035 diff_3403000_5587000# diff_775000_5103000# diff_83000_3098000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2036 diff_3442000_5621000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2037 diff_3560000_5621000# diff_775000_5103000# diff_83000_3098000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2038 diff_3834000_5621000# diff_775000_5103000# diff_83000_3098000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2039 diff_3952000_5621000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2040 diff_4011000_5621000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2041 diff_4031000_5587000# diff_775000_5103000# diff_83000_3098000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2042 diff_4070000_5621000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2043 diff_4149000_5587000# diff_775000_5103000# diff_83000_3098000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2044 diff_4346000_5621000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2045 diff_4788000_5621000# diff_775000_5103000# diff_83000_3098000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2046 diff_4847000_5621000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2047 diff_4867000_5587000# diff_775000_5103000# diff_83000_3098000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2048 diff_4906000_5621000# diff_775000_5103000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2049 diff_4926000_5587000# diff_775000_5103000# diff_83000_3098000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2050 diff_83000_3098000# diff_5252000_5062000# diff_778000_5046000# GND efet w=179000 l=9000
+ ad=0 pd=0 as=2.01603e+09 ps=956000 
M2051 diff_778000_5046000# diff_5502000_5120000# diff_83000_3098000# GND efet w=178000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2052 diff_5501000_5152000# diff_5501000_5152000# diff_95000_5192000# GND efet w=12000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M2053 diff_5501000_5152000# diff_5954000_5147000# diff_5700000_5120000# GND efet w=13000 l=13000
+ ad=0 pd=0 as=5.28e+08 ps=144000 
M2054 diff_95000_5192000# diff_5972000_5106000# diff_5972000_5106000# GND efet w=11000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M2055 diff_6226000_5161000# diff_72000_4515000# diff_6074000_5171000# GND efet w=20000 l=11000
+ ad=-1.07497e+09 pd=628000 as=3.4e+08 ps=88000 
M2056 diff_6226000_5191000# diff_6226000_5191000# diff_95000_5192000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M2057 diff_83000_3098000# diff_775000_5076000# diff_761000_5561000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2058 diff_83000_3098000# diff_775000_5076000# diff_797000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2059 diff_83000_3098000# diff_775000_5076000# diff_1169000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2060 diff_83000_3098000# diff_775000_5076000# diff_1286000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2061 diff_83000_3098000# diff_775000_5076000# diff_1306000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2062 diff_83000_3098000# diff_775000_5076000# diff_1366000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2063 diff_83000_3098000# diff_775000_5076000# diff_1424000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2064 diff_83000_3098000# diff_775000_5076000# diff_1522000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2065 diff_83000_3098000# diff_775000_5076000# diff_1639000_5587000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2066 diff_83000_3098000# diff_775000_5076000# diff_1678000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2067 diff_83000_3098000# diff_775000_5076000# diff_1795000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2068 diff_83000_3098000# diff_775000_5076000# diff_1944000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2069 diff_83000_3098000# diff_775000_5076000# diff_1964000_5587000# GND efet w=22000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2070 diff_83000_3098000# diff_775000_5076000# diff_2022000_5587000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2071 diff_83000_3098000# diff_775000_5076000# diff_2119000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2072 diff_83000_3098000# diff_775000_5076000# diff_2238000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2073 diff_83000_3098000# diff_775000_5076000# diff_2276000_5621000# GND efet w=22000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2074 diff_83000_3098000# diff_775000_5076000# diff_2541000_5621000# GND efet w=22000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2075 diff_83000_3098000# diff_775000_5076000# diff_2815000_5621000# GND efet w=22000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2076 diff_83000_3098000# diff_775000_5076000# diff_2835000_5587000# GND efet w=22000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2077 diff_83000_3098000# diff_775000_5076000# diff_2953000_5587000# GND efet w=22000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2078 diff_83000_3098000# diff_775000_5076000# diff_3012000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2079 diff_83000_3098000# diff_775000_5076000# diff_3071000_5587000# GND efet w=22000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2080 diff_83000_3098000# diff_775000_5076000# diff_3324000_5621000# GND efet w=22000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2081 diff_83000_3098000# diff_775000_5076000# diff_3403000_5587000# GND efet w=22000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2082 diff_83000_3098000# diff_775000_5076000# diff_3462000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2083 diff_83000_3098000# diff_775000_5076000# diff_3580000_5587000# GND efet w=22000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2084 diff_83000_3098000# diff_775000_5076000# diff_3639000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2085 diff_83000_3098000# diff_775000_5076000# diff_3678000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2086 diff_83000_3098000# diff_775000_5076000# diff_3776000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2087 diff_83000_3098000# diff_775000_5076000# diff_3796000_5587000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2088 diff_83000_3098000# diff_775000_5076000# diff_4011000_5621000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2089 diff_83000_3098000# diff_775000_5076000# diff_4208000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2090 diff_83000_3098000# diff_775000_5076000# diff_4405000_5621000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2091 diff_83000_3098000# diff_775000_5076000# diff_4425000_5587000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2092 diff_83000_3098000# diff_775000_5076000# diff_4484000_5587000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2093 diff_83000_3098000# diff_775000_5076000# diff_4808000_5587000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2094 diff_487000_5098000# diff_487000_5098000# diff_95000_5192000# GND efet w=13000 l=14000
+ ad=1.775e+09 pd=376000 as=0 ps=0 
M2095 diff_376000_4961000# diff_68000_5288000# diff_95000_5192000# GND efet w=171500 l=9500
+ ad=1.81303e+09 pd=964000 as=0 ps=0 
M2096 diff_95000_5192000# diff_376000_4961000# diff_376000_4961000# GND efet w=11000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M2097 diff_487000_5098000# diff_376000_4961000# diff_83000_3098000# GND efet w=96500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2098 diff_474000_5143000# diff_487000_5098000# diff_95000_5192000# GND efet w=35000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2099 diff_95000_5192000# diff_778000_5046000# diff_778000_5046000# GND efet w=14000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2100 diff_83000_3098000# diff_5700000_5120000# diff_5502000_5120000# GND efet w=101000 l=9000
+ ad=0 pd=0 as=-1.28997e+09 ps=628000 
M2101 diff_83000_3098000# diff_6062000_5632000# diff_5972000_5106000# GND efet w=113500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2102 diff_95000_5192000# diff_5502000_5120000# diff_5502000_5120000# GND efet w=13000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M2103 diff_5502000_5120000# diff_5502000_5120000# diff_5502000_5120000# GND efet w=500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2104 diff_5700000_5120000# diff_474000_5143000# diff_5972000_5106000# GND efet w=12000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M2105 diff_6062000_5632000# diff_72000_4515000# diff_667000_3269000# GND efet w=55000 l=12000
+ ad=5.1e+08 pd=156000 as=7.89033e+08 ps=1.014e+06 
M2106 diff_83000_3098000# diff_5596000_414000# diff_6226000_5191000# GND efet w=149000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2107 diff_95000_5192000# diff_6226000_5161000# diff_6226000_5161000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2108 diff_83000_3098000# diff_4952000_396000# diff_6226000_5161000# GND efet w=148500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M2109 diff_5252000_5062000# diff_5252000_5062000# diff_95000_5192000# GND efet w=17000 l=8000
+ ad=-1.48797e+09 pd=592000 as=0 ps=0 
M2110 diff_83000_3098000# diff_376000_4961000# diff_5252000_5062000# GND efet w=208500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M2111 diff_855000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2112 diff_953000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2113 diff_1032000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2114 diff_1248000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2115 diff_1404000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2116 diff_1464000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2117 diff_1542000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2118 diff_1619000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2119 diff_1698000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2120 diff_1737000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2121 diff_1757000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2122 diff_1815000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2123 diff_2002000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2124 diff_2061000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2125 diff_2081000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2126 diff_2139000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2127 diff_2218000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2128 diff_2296000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2129 diff_2335000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2130 diff_2355000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2131 diff_2483000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2132 diff_2503000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2133 diff_2620000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2134 diff_2679000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2135 diff_2874000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2136 diff_2894000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2137 diff_2992000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2138 diff_3051000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2139 diff_3110000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2140 diff_3130000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2141 diff_3383000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2142 diff_3442000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2143 diff_3501000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2144 diff_3521000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2145 diff_3560000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2146 diff_3619000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2147 diff_3834000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2148 diff_3854000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2149 diff_3952000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2150 diff_3972000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2151 diff_4031000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2152 diff_4070000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2153 diff_4090000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2154 diff_4149000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2155 diff_4288000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2156 diff_4346000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2157 diff_4464000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2158 diff_4523000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2159 diff_4602000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2160 diff_4730000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2161 diff_4750000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2162 diff_4788000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2163 diff_4847000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2164 diff_4867000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2165 diff_4906000_5621000# diff_778000_5046000# diff_83000_3098000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2166 diff_4926000_5587000# diff_778000_5046000# diff_83000_3098000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2167 diff_83000_3098000# diff_506000_5537000# diff_953000_5621000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2168 diff_83000_3098000# diff_506000_5537000# diff_1188000_5587000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2169 diff_83000_3098000# diff_506000_5537000# diff_1248000_5587000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2170 diff_83000_3098000# diff_506000_5537000# diff_1286000_5621000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2171 diff_83000_3098000# diff_506000_5537000# diff_1306000_5587000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2172 diff_83000_3098000# diff_506000_5537000# diff_1484000_5587000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2173 diff_83000_3098000# diff_506000_5537000# diff_1522000_5621000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2174 diff_83000_3098000# diff_506000_5537000# diff_1737000_5621000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2175 diff_83000_3098000# diff_506000_5537000# diff_1795000_5621000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2176 diff_83000_3098000# diff_506000_5537000# diff_2002000_5621000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2177 diff_83000_3098000# diff_506000_5537000# diff_2022000_5587000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2178 diff_83000_3098000# diff_506000_5537000# diff_2335000_5621000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2179 diff_83000_3098000# diff_506000_5537000# diff_2355000_5587000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2180 diff_83000_3098000# diff_506000_5537000# diff_2414000_5587000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2181 diff_83000_3098000# diff_506000_5537000# diff_2483000_5621000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2182 diff_83000_3098000# diff_506000_5537000# diff_2503000_5587000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2183 diff_83000_3098000# diff_506000_5537000# diff_2874000_5621000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2184 diff_83000_3098000# diff_506000_5537000# diff_3051000_5621000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2185 diff_83000_3098000# diff_506000_5537000# diff_3130000_5587000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2186 diff_83000_3098000# diff_506000_5537000# diff_3560000_5621000# GND efet w=21000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2187 diff_83000_3098000# diff_506000_5537000# diff_4070000_5621000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2188 diff_83000_3098000# diff_506000_5537000# diff_4867000_5587000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2189 diff_83000_3098000# diff_446000_4910000# diff_376000_4961000# GND efet w=255500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2190 diff_376000_4961000# diff_68000_5288000# diff_95000_5192000# GND efet w=34000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2191 diff_376000_4961000# diff_446000_4910000# diff_83000_3098000# GND efet w=182000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2192 diff_85000_5213000# diff_85000_5213000# diff_95000_5192000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2193 diff_83000_3098000# diff_68000_5288000# diff_446000_4910000# GND efet w=172000 l=9000
+ ad=0 pd=0 as=1.64903e+09 ps=946000 
M2194 diff_761000_5561000# diff_376000_4961000# diff_700000_4694000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.27e+08 ps=88000 
M2195 diff_797000_5587000# diff_376000_4961000# diff_668000_4504000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2196 diff_835000_5621000# diff_376000_4961000# diff_764000_4721000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2197 diff_855000_5587000# diff_376000_4961000# diff_831000_4716000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.04e+08 ps=70000 
M2198 diff_894000_5621000# diff_376000_4961000# diff_861000_4716000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2199 diff_914000_5587000# diff_376000_4961000# diff_888000_4706000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.04e+08 ps=70000 
M2200 diff_953000_5621000# diff_376000_4961000# diff_886000_3953000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2201 diff_973000_5587000# diff_376000_4961000# diff_988000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2202 diff_1012000_5621000# diff_376000_4961000# diff_1018000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.14e+08 ps=86000 
M2203 diff_1032000_5587000# diff_376000_4961000# diff_984000_4377000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2204 diff_1110000_5621000# diff_376000_4961000# diff_1038000_4590000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.05e+08 ps=72000 
M2205 diff_1130000_5587000# diff_376000_4961000# diff_1146000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.2e+08 ps=86000 
M2206 diff_1169000_5621000# diff_376000_4961000# diff_1145000_4574000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2207 diff_1188000_5587000# diff_376000_4961000# diff_1204000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2208 diff_1228000_5621000# diff_376000_4961000# diff_1233000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.27e+08 ps=88000 
M2209 diff_1248000_5587000# diff_376000_4961000# diff_1263000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2210 diff_1286000_5621000# diff_376000_4961000# diff_1292000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.13e+08 ps=86000 
M2211 diff_1306000_5587000# diff_376000_4961000# diff_1322000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.2e+08 ps=84000 
M2212 diff_1346000_5621000# diff_376000_4961000# diff_1351000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.43e+08 ps=88000 
M2213 diff_1366000_5587000# diff_376000_4961000# diff_1381000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.43e+08 ps=86000 
M2214 diff_1404000_5621000# diff_376000_4961000# diff_1410000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.2e+08 ps=86000 
M2215 diff_1424000_5587000# diff_376000_4961000# diff_1440000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.2e+08 ps=86000 
M2216 diff_1464000_5621000# diff_376000_4961000# diff_1469000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2217 diff_1484000_5587000# diff_376000_4961000# diff_1499000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.43e+08 ps=88000 
M2218 diff_1522000_5621000# diff_376000_4961000# diff_1528000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2219 diff_1542000_5587000# diff_376000_4961000# diff_1557000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.43e+08 ps=88000 
M2220 diff_1619000_5621000# diff_376000_4961000# diff_1625000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2221 diff_1639000_5587000# diff_376000_4961000# diff_1655000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.2e+08 ps=86000 
M2222 diff_1678000_5621000# diff_376000_4961000# diff_1683000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2223 diff_1698000_5587000# diff_376000_4961000# diff_1713000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.04e+08 ps=86000 
M2224 diff_1737000_5621000# diff_376000_4961000# diff_1742000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2225 diff_1757000_5587000# diff_376000_4961000# diff_1772000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2226 diff_1795000_5621000# diff_376000_4961000# diff_1801000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2227 diff_1815000_5587000# diff_376000_4961000# diff_1831000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2228 diff_446000_4910000# diff_197000_5470000# diff_83000_3098000# GND efet w=173000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2229 diff_95000_5192000# diff_77000_4827000# diff_77000_4827000# GND efet w=34000 l=8000
+ ad=0 pd=0 as=2.14033e+08 ps=738000 
M2230 diff_83000_3098000# diff_78000_4695000# diff_77000_4827000# GND efet w=322500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2231 diff_446000_4910000# diff_409000_4783000# diff_83000_3098000# GND efet w=178000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2232 diff_83000_3098000# diff_88000_5400000# diff_78000_4695000# GND efet w=182000 l=8000
+ ad=0 pd=0 as=2.00903e+09 ps=1.054e+06 
M2233 diff_95000_5192000# diff_78000_4695000# diff_78000_4695000# GND efet w=12000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2234 diff_83000_3098000# diff_201000_4774000# diff_78000_4695000# GND efet w=178000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2235 diff_83000_3098000# diff_85000_4683000# diff_78000_4695000# GND efet w=178000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2236 diff_231000_4715000# diff_205000_4722000# diff_83000_3098000# GND efet w=75500 l=8500
+ ad=1.352e+09 pd=274000 as=0 ps=0 
M2237 diff_409000_4783000# diff_100000_3992000# diff_83000_3098000# GND efet w=68000 l=8000
+ ad=1.172e+09 pd=222000 as=0 ps=0 
M2238 diff_95000_5192000# diff_409000_4783000# diff_409000_4783000# GND efet w=11000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2239 diff_446000_4910000# diff_446000_4910000# diff_95000_5192000# GND efet w=13000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2240 diff_201000_4774000# diff_72000_4515000# diff_231000_4715000# GND efet w=17000 l=11000
+ ad=3.54e+08 pd=100000 as=0 ps=0 
M2241 diff_205000_4722000# diff_68000_5288000# diff_121000_4669000# GND efet w=13000 l=11000
+ ad=2.34e+08 pd=78000 as=1.8e+09 ps=330000 
M2242 diff_231000_4715000# diff_231000_4715000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2243 diff_83000_3098000# diff_85000_4683000# diff_121000_4669000# GND efet w=64000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2244 diff_95000_5192000# diff_121000_4669000# diff_121000_4669000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2245 diff_85000_4683000# diff_85000_4683000# diff_95000_5192000# GND efet w=13000 l=14000
+ ad=-8.22967e+08 pd=640000 as=0 ps=0 
M2246 diff_85000_4683000# diff_64000_4639000# diff_83000_3098000# GND efet w=105000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2247 diff_85000_4683000# diff_197000_5470000# diff_83000_3098000# GND efet w=106000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2248 diff_64000_4639000# diff_230000_4601000# diff_83000_3098000# GND efet w=107500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2249 diff_83000_3098000# diff_81000_4527000# diff_64000_4639000# GND efet w=104000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2250 diff_95000_5192000# diff_64000_4639000# diff_64000_4639000# GND efet w=13000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M2251 diff_83000_3098000# diff_106000_4536000# diff_64000_4639000# GND efet w=114000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2252 diff_64000_4639000# diff_216000_4574000# diff_83000_3098000# GND efet w=104000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2253 diff_153000_4530000# diff_169000_4545000# diff_83000_3098000# GND efet w=103500 l=8500
+ ad=1.73e+09 pd=314000 as=0 ps=0 
M2254 diff_153000_4530000# diff_72000_4515000# diff_106000_4536000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=2.28e+08 ps=70000 
M2255 diff_81000_4527000# diff_72000_4515000# diff_74000_3122000# GND efet w=21000 l=12000
+ ad=3.82e+08 pd=104000 as=-1.97197e+09 ps=456000 
M2256 diff_153000_4530000# diff_153000_4530000# diff_95000_5192000# GND efet w=14000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M2257 diff_216000_4574000# diff_72000_4515000# diff_337000_4528000# GND efet w=13000 l=12000
+ ad=2.13e+08 pd=68000 as=-1.30897e+09 ps=610000 
M2258 diff_571000_4610000# diff_559000_4358000# diff_83000_3098000# GND efet w=197500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2259 diff_83000_3098000# diff_700000_4694000# diff_642000_4583000# GND efet w=42000 l=8000
+ ad=0 pd=0 as=1.524e+09 ps=320000 
M2260 diff_83000_3098000# diff_65000_4220000# diff_83000_4448000# GND efet w=65000 l=8000
+ ad=0 pd=0 as=-2.03797e+09 ps=436000 
M2261 diff_83000_3098000# diff_167000_4461000# diff_83000_4448000# GND efet w=64000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2262 diff_83000_4448000# diff_72000_4515000# diff_81000_4321000# GND efet w=18000 l=12000
+ ad=0 pd=0 as=1.01e+09 ps=274000 
M2263 diff_95000_5192000# diff_83000_4448000# diff_83000_4448000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2264 diff_83000_3098000# diff_81000_4321000# diff_109000_4359000# GND efet w=75000 l=8000
+ ad=0 pd=0 as=1.117e+09 ps=234000 
M2265 diff_95000_5192000# diff_109000_4359000# diff_109000_4359000# GND efet w=11000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2266 diff_83000_3098000# diff_109000_4359000# diff_88000_4249000# GND efet w=64500 l=9500
+ ad=0 pd=0 as=1.256e+09 ps=284000 
M2267 diff_88000_4249000# diff_68000_5288000# diff_81000_4321000# GND efet w=18000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2268 diff_95000_5192000# diff_88000_4249000# diff_88000_4249000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2269 diff_95000_5192000# diff_480000_4480000# diff_480000_4480000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=-1.30897e+09 ps=528000 
M2270 diff_83000_3098000# diff_531000_4622000# diff_520000_4360000# GND efet w=129000 l=7000
+ ad=0 pd=0 as=-1.22597e+09 ps=632000 
M2271 diff_571000_4610000# diff_571000_4610000# diff_95000_5192000# GND efet w=12000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2272 diff_96000_4258000# diff_88000_4249000# diff_78000_4235000# GND efet w=103500 l=8500
+ ad=-2.01397e+09 pd=482000 as=6.33033e+08 ps=776000 
M2273 diff_83000_3098000# diff_106000_4268000# diff_96000_4258000# GND efet w=206000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2274 diff_314000_4258000# diff_314000_4258000# diff_95000_5192000# GND efet w=12000 l=14000
+ ad=2.021e+09 pd=388000 as=0 ps=0 
M2275 diff_78000_4235000# diff_88000_4249000# diff_96000_4258000# GND efet w=121000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2276 diff_314000_4258000# diff_72000_4515000# diff_106000_4268000# GND efet w=25000 l=11000
+ ad=0 pd=0 as=3.93e+08 ps=114000 
M2277 diff_83000_3098000# diff_101000_4084000# diff_78000_4235000# GND efet w=131500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M2278 diff_95000_5192000# diff_78000_4235000# diff_78000_4235000# GND efet w=12000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M2279 diff_167000_4461000# diff_167000_4461000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=-1.56597e+09 pd=530000 as=0 ps=0 
M2280 diff_83000_3098000# diff_354000_4247000# diff_314000_4258000# GND efet w=108000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2281 diff_520000_4360000# diff_512000_4352000# diff_480000_4480000# GND efet w=133500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2282 diff_83000_3098000# diff_530000_4372000# diff_520000_4360000# GND efet w=147000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2283 diff_642000_4583000# diff_642000_4583000# diff_95000_5192000# GND efet w=13000 l=35000
+ ad=0 pd=0 as=0 ps=0 
M2284 diff_83000_3098000# diff_668000_4504000# diff_642000_4583000# GND efet w=43000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2285 diff_95000_5192000# diff_578000_4447000# diff_578000_4447000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=1.521e+09 ps=320000 
M2286 diff_83000_3098000# diff_583000_4388000# diff_578000_4447000# GND efet w=67500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2287 diff_739000_4508000# diff_725000_4490000# diff_686000_4521000# GND efet w=214500 l=7500
+ ad=2.10503e+09 pd=1.088e+06 as=-1.09197e+09 ps=684000 
M2288 diff_782000_4737000# diff_782000_4737000# diff_95000_5192000# GND efet w=11000 l=36000
+ ad=1.061e+09 pd=256000 as=0 ps=0 
M2289 diff_83000_3098000# diff_831000_4716000# diff_782000_4737000# GND efet w=43000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M2290 diff_861000_4692000# diff_861000_4716000# diff_83000_3098000# GND efet w=43000 l=8000
+ ad=1.373e+09 pd=278000 as=0 ps=0 
M2291 diff_1014000_4730000# diff_988000_4962000# diff_83000_3098000# GND efet w=139500 l=8500
+ ad=3.09033e+08 pd=734000 as=0 ps=0 
M2292 diff_83000_3098000# diff_888000_4706000# diff_861000_4692000# GND efet w=41000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2293 diff_95000_5192000# diff_686000_4521000# diff_686000_4521000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2294 diff_654000_4324000# diff_72000_4515000# diff_625000_4565000# GND efet w=12000 l=11000
+ ad=4.43e+08 pd=138000 as=-2.03097e+09 ps=482000 
M2295 diff_861000_4692000# diff_861000_4692000# diff_95000_5192000# GND efet w=13000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M2296 diff_793000_4433000# diff_764000_4721000# diff_725000_4490000# GND efet w=132000 l=8000
+ ad=1.191e+09 pd=282000 as=9.80327e+07 ps=786000 
M2297 diff_83000_3098000# diff_530000_4372000# diff_793000_4433000# GND efet w=132000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2298 diff_836000_4491000# diff_782000_4737000# diff_83000_3098000# GND efet w=206500 l=7500
+ ad=1.952e+09 pd=432000 as=0 ps=0 
M2299 diff_853000_4510000# diff_791000_4022000# diff_836000_4491000# GND efet w=207500 l=8500
+ ad=1.948e+09 pd=432000 as=0 ps=0 
M2300 diff_725000_4490000# diff_861000_4692000# diff_853000_4510000# GND efet w=206500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2301 diff_1014000_4730000# diff_597000_3013000# diff_936000_4586000# GND efet w=129000 l=8000
+ ad=0 pd=0 as=1.928e+09 ps=472000 
M2302 diff_83000_3098000# diff_1018000_4962000# diff_1014000_4730000# GND efet w=130000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2303 diff_936000_4586000# diff_936000_4586000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2304 diff_95000_5192000# diff_725000_4490000# diff_725000_4490000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2305 diff_583000_4388000# diff_72000_4515000# diff_480000_4480000# GND efet w=12000 l=11000
+ ad=2.68e+08 pd=94000 as=0 ps=0 
M2306 diff_167000_4461000# diff_301000_4194000# diff_83000_3098000# GND efet w=67000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2307 diff_222000_4165000# diff_68000_5288000# diff_101000_4084000# GND efet w=14000 l=10000
+ ad=3.38e+08 pd=104000 as=-8.95967e+08 ps=678000 
M2308 diff_83000_3098000# diff_222000_4165000# diff_167000_4461000# GND efet w=73000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2309 diff_83000_3098000# diff_128000_4097000# diff_101000_4084000# GND efet w=118500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2310 diff_354000_4247000# diff_68000_5288000# diff_128000_4097000# GND efet w=19000 l=12000
+ ad=3.31e+08 pd=78000 as=1.978e+09 ps=408000 
M2311 diff_83000_3098000# diff_578000_4447000# diff_559000_4358000# GND efet w=65000 l=8000
+ ad=0 pd=0 as=2.00003e+09 ps=1.184e+06 
M2312 diff_559000_4358000# diff_654000_4324000# diff_83000_3098000# GND efet w=77000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2313 diff_83000_3098000# diff_680000_4314000# diff_559000_4358000# GND efet w=60000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2314 diff_95000_5192000# diff_101000_4084000# diff_101000_4084000# GND efet w=12000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M2315 diff_101000_4084000# diff_78000_4235000# diff_83000_3098000# GND efet w=104000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2316 diff_282000_4044000# diff_282000_4044000# diff_95000_5192000# GND efet w=12000 l=15000
+ ad=2.037e+09 pd=384000 as=0 ps=0 
M2317 diff_282000_4044000# diff_169000_4545000# diff_83000_3098000# GND efet w=91000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2318 diff_282000_4044000# diff_169000_4545000# diff_83000_3098000# GND efet w=15000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2319 diff_83000_3098000# diff_282000_4044000# diff_130000_3949000# GND efet w=115000 l=8000
+ ad=0 pd=0 as=2.048e+09 ps=366000 
M2320 diff_83000_3098000# diff_100000_3992000# diff_106000_3785000# GND efet w=107500 l=7500
+ ad=0 pd=0 as=-1.82497e+09 ps=380000 
M2321 diff_95000_5192000# diff_106000_3785000# diff_106000_3785000# GND efet w=11000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M2322 diff_130000_3949000# diff_130000_3949000# diff_95000_5192000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M2323 diff_83000_3098000# diff_130000_3949000# diff_106000_3785000# GND efet w=116000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2324 diff_130000_3949000# diff_230000_4601000# diff_83000_3098000# GND efet w=100000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2325 diff_101000_4084000# diff_68000_5288000# diff_132000_3835000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.56e+08 ps=92000 
M2326 diff_337000_4528000# diff_232000_3858000# diff_83000_3098000# GND efet w=110500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2327 diff_139000_3844000# diff_132000_3835000# diff_83000_3098000# GND efet w=158000 l=8000
+ ad=-1.56897e+09 pd=550000 as=0 ps=0 
M2328 diff_232000_3858000# diff_232000_3858000# diff_95000_5192000# GND efet w=11000 l=21000
+ ad=1.783e+09 pd=378000 as=0 ps=0 
M2329 diff_232000_3858000# diff_94000_3753000# diff_139000_3844000# GND efet w=169500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2330 diff_337000_4528000# diff_337000_4528000# diff_95000_5192000# GND efet w=12000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M2331 diff_139000_3844000# diff_74000_3122000# diff_83000_3098000# GND efet w=25000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2332 diff_139000_3844000# diff_74000_3122000# diff_83000_3098000# GND efet w=104000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2333 diff_725000_4204000# diff_642000_4583000# diff_83000_3098000# GND efet w=200500 l=7500
+ ad=9.06033e+08 pd=984000 as=0 ps=0 
M2334 diff_739000_4508000# diff_668000_4504000# diff_725000_4204000# GND efet w=198500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2335 diff_725000_4204000# diff_757000_4475000# diff_739000_4508000# GND efet w=201000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2336 diff_95000_5192000# diff_559000_4358000# diff_559000_4358000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2337 diff_83000_3098000# diff_637000_4100000# diff_559000_4358000# GND efet w=77500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2338 diff_559000_4358000# diff_659000_4117000# diff_83000_3098000# GND efet w=75000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2339 diff_83000_3098000# diff_691000_4135000# diff_559000_4358000# GND efet w=64000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2340 diff_83000_3098000# diff_773000_4078000# diff_725000_4204000# GND efet w=199500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2341 diff_1024000_4536000# diff_519000_3032000# diff_83000_3098000# GND efet w=157500 l=8500
+ ad=1.30327e+07 pd=788000 as=0 ps=0 
M2342 diff_1076000_4557000# diff_1076000_4557000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=1.985e+09 pd=486000 as=0 ps=0 
M2343 diff_1158000_4673000# diff_519000_3032000# diff_1076000_4557000# GND efet w=130000 l=8000
+ ad=1.3e+09 pd=280000 as=0 ps=0 
M2344 diff_83000_3098000# diff_1146000_4962000# diff_1158000_4673000# GND efet w=130000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2345 diff_1177000_4478000# diff_1145000_4574000# diff_83000_3098000# GND efet w=42000 l=8000
+ ad=1.115e+09 pd=224000 as=0 ps=0 
M2346 diff_991000_4386000# diff_984000_4377000# diff_975000_4364000# GND efet w=145500 l=7500
+ ad=1.447e+09 pd=312000 as=-1.94397e+09 ps=552000 
M2347 diff_83000_3098000# diff_1001000_4394000# diff_991000_4386000# GND efet w=145500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2348 diff_1024000_4536000# diff_597000_3013000# diff_83000_3098000# GND efet w=162500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2349 diff_1053000_4267000# diff_1038000_4590000# diff_1024000_4536000# GND efet w=149500 l=8500
+ ad=-1.67497e+09 pd=558000 as=0 ps=0 
M2350 diff_531000_4622000# diff_72000_4515000# diff_1126000_4459000# GND efet w=11000 l=10000
+ ad=-1.18293e+09 pd=1.112e+06 as=2.73e+08 ps=104000 
M2351 diff_83000_3098000# diff_106000_3785000# diff_94000_3753000# GND efet w=104000 l=8000
+ ad=0 pd=0 as=-8.49967e+08 ps=624000 
M2352 diff_95000_5192000# diff_94000_3753000# diff_94000_3753000# GND efet w=13000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M2353 diff_83000_3098000# diff_92000_3714000# diff_94000_3753000# GND efet w=108000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2354 diff_94000_3753000# diff_197000_5470000# diff_83000_3098000# GND efet w=104500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2355 diff_83000_3098000# diff_118000_3658000# diff_92000_3714000# GND efet w=195000 l=8000
+ ad=0 pd=0 as=-1.99493e+09 ps=1.116e+06 
M2356 diff_92000_3714000# diff_94000_3551000# diff_83000_3098000# GND efet w=173500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2357 diff_185000_3712000# diff_68000_5288000# diff_118000_3658000# GND efet w=12000 l=11000
+ ad=1.213e+09 pd=250000 as=2.17e+08 ps=70000 
M2358 diff_95000_5192000# diff_185000_3712000# diff_185000_3712000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2359 diff_185000_3712000# diff_182000_3691000# diff_83000_3098000# GND efet w=72000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2360 diff_197000_5470000# diff_72000_4515000# diff_182000_3691000# GND efet w=13000 l=11000
+ ad=0 pd=0 as=2.32e+08 ps=82000 
M2361 diff_83000_3098000# diff_197000_5470000# diff_92000_3714000# GND efet w=63000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2362 diff_92000_3714000# diff_197000_5470000# diff_83000_3098000# GND efet w=101500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M2363 diff_92000_3714000# diff_92000_3714000# diff_95000_5192000# GND efet w=12000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2364 diff_650000_3859000# diff_608000_3765000# diff_83000_3098000# GND efet w=139500 l=8500
+ ad=1.28e+09 pd=298000 as=0 ps=0 
M2365 diff_635000_3800000# diff_660000_3853000# diff_650000_3859000# GND efet w=139500 l=8500
+ ad=1.19903e+09 pd=954000 as=0 ps=0 
M2366 diff_660000_3853000# diff_72000_4515000# diff_732000_3738000# GND efet w=14000 l=13000
+ ad=2.39e+08 pd=78000 as=-1.18697e+09 ps=568000 
M2367 diff_695000_3858000# diff_687000_3826000# diff_635000_3800000# GND efet w=130000 l=8000
+ ad=1.17e+09 pd=278000 as=0 ps=0 
M2368 diff_83000_3098000# diff_230000_4601000# diff_695000_3858000# GND efet w=130000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2369 diff_732000_3738000# diff_230000_4601000# diff_83000_3098000# GND efet w=97500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M2370 diff_83000_3098000# diff_752000_3797000# diff_732000_3738000# GND efet w=64000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2371 diff_635000_3800000# diff_635000_3800000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2372 diff_687000_3826000# diff_72000_4515000# diff_169000_4545000# GND efet w=12000 l=11000
+ ad=4.42e+08 pd=134000 as=-1.59497e+09 ps=580000 
M2373 diff_608000_3765000# diff_72000_4515000# diff_337000_4528000# GND efet w=11000 l=11000
+ ad=7.55e+08 pd=204000 as=0 ps=0 
M2374 diff_809000_3854000# diff_570000_3597000# diff_792000_3825000# GND efet w=142500 l=7500
+ ad=1.441e+09 pd=304000 as=-8.61967e+08 ps=708000 
M2375 diff_83000_3098000# diff_660000_3853000# diff_809000_3854000# GND efet w=142000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2376 diff_975000_4364000# diff_975000_4364000# diff_95000_5192000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M2377 diff_1053000_4267000# diff_1053000_4267000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2378 diff_1177000_4478000# diff_1177000_4478000# diff_95000_5192000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M2379 diff_1944000_5621000# diff_376000_4961000# diff_1949000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2380 diff_1964000_5587000# diff_376000_4961000# diff_1979000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.2e+08 ps=86000 
M2381 diff_2002000_5621000# diff_376000_4961000# diff_2007000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2382 diff_2022000_5587000# diff_376000_4961000# diff_2037000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2383 diff_2061000_5621000# diff_376000_4961000# diff_2067000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2384 diff_2081000_5587000# diff_376000_4961000# diff_2097000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.13e+08 ps=86000 
M2385 diff_2119000_5621000# diff_376000_4961000# diff_2125000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.2e+08 ps=86000 
M2386 diff_2139000_5587000# diff_376000_4961000# diff_2155000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.04e+08 ps=86000 
M2387 diff_2218000_5621000# diff_376000_4961000# diff_2223000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.27e+08 ps=88000 
M2388 diff_2238000_5587000# diff_376000_4961000# diff_2253000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2389 diff_2276000_5621000# diff_376000_4961000# diff_2282000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2390 diff_2296000_5587000# diff_376000_4961000# diff_2312000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2391 diff_2335000_5621000# diff_376000_4961000# diff_2341000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2392 diff_2355000_5587000# diff_376000_4961000# diff_2371000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2393 diff_2394000_5621000# diff_376000_4961000# diff_2399000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2394 diff_2414000_5587000# diff_376000_4961000# diff_2429000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2395 diff_2483000_5621000# diff_376000_4961000# diff_2488000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2396 diff_2503000_5587000# diff_376000_4961000# diff_2518000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2397 diff_2541000_5621000# diff_376000_4961000# diff_2547000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2398 diff_2561000_5587000# diff_376000_4961000# diff_2577000_4949000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=1.96e+08 ps=72000 
M2399 diff_2600000_5621000# diff_376000_4961000# diff_2606000_4947000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.04e+08 ps=70000 
M2400 diff_2620000_5587000# diff_376000_4961000# diff_2636000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2401 diff_2659000_5621000# diff_376000_4961000# diff_2664000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.28e+08 ps=90000 
M2402 diff_2679000_5587000# diff_376000_4961000# diff_2694000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2403 diff_2757000_5621000# diff_376000_4961000# diff_2762000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2404 diff_2777000_5587000# diff_376000_4961000# diff_2792000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.43e+08 ps=88000 
M2405 diff_2815000_5621000# diff_376000_4961000# diff_2821000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2406 diff_2835000_5587000# diff_376000_4961000# diff_2851000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=1.217e+09 ps=338000 
M2407 diff_2874000_5621000# diff_376000_4961000# diff_2880000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2408 diff_2894000_5587000# diff_376000_4961000# diff_2910000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.2e+08 ps=86000 
M2409 diff_2933000_5621000# diff_376000_4961000# diff_2849000_2986000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.27e+08 ps=88000 
M2410 diff_2953000_5587000# diff_376000_4961000# diff_2968000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2411 diff_2992000_5621000# diff_376000_4961000# diff_2998000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2412 diff_3012000_5587000# diff_376000_4961000# diff_3028000_4947000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.05e+08 ps=72000 
M2413 diff_3051000_5621000# diff_376000_4961000# diff_3056000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.27e+08 ps=88000 
M2414 diff_3071000_5587000# diff_376000_4961000# diff_3086000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2415 diff_3110000_5621000# diff_376000_4961000# diff_3116000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2416 diff_3130000_5587000# diff_376000_4961000# diff_3106000_3438000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=70000 
M2417 diff_3169000_5621000# diff_376000_4961000# diff_3174000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.43e+08 ps=88000 
M2418 diff_3189000_5587000# diff_376000_4961000# diff_3204000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.43e+08 ps=88000 
M2419 diff_3266000_5621000# diff_376000_4961000# diff_3271000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.43e+08 ps=88000 
M2420 diff_3286000_5587000# diff_376000_4961000# diff_3301000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2421 diff_3324000_5621000# diff_376000_4961000# diff_3330000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2422 diff_3344000_5587000# diff_376000_4961000# diff_3360000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.2e+08 ps=86000 
M2423 diff_3383000_5621000# diff_376000_4961000# diff_3389000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.2e+08 ps=86000 
M2424 diff_3403000_5587000# diff_376000_4961000# diff_3419000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=1.96e+08 ps=88000 
M2425 diff_3442000_5621000# diff_376000_4961000# diff_3447000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.29e+08 ps=90000 
M2426 diff_3462000_5587000# diff_376000_4961000# diff_3477000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2427 diff_3501000_5621000# diff_376000_4961000# diff_3507000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2428 diff_3521000_5587000# diff_376000_4961000# diff_3537000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.05e+08 ps=88000 
M2429 diff_3560000_5621000# diff_376000_4961000# diff_3565000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.27e+08 ps=90000 
M2430 diff_3580000_5587000# diff_376000_4961000# diff_3595000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.28e+08 ps=90000 
M2431 diff_3619000_5621000# diff_376000_4961000# diff_3625000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2432 diff_3639000_5587000# diff_376000_4961000# diff_3654000_3515000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2433 diff_3678000_5621000# diff_376000_4961000# diff_3683000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.43e+08 ps=88000 
M2434 diff_3698000_5587000# diff_376000_4961000# diff_3713000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.36e+08 ps=90000 
M2435 diff_3776000_5621000# diff_376000_4961000# diff_3781000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.27e+08 ps=88000 
M2436 diff_3796000_5587000# diff_376000_4961000# diff_3811000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2437 diff_3834000_5621000# diff_376000_4961000# diff_3840000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2438 diff_3854000_5587000# diff_376000_4961000# diff_3870000_4934000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.04e+08 ps=70000 
M2439 diff_3893000_5621000# diff_376000_4961000# diff_3899000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.04e+08 ps=88000 
M2440 diff_3913000_5587000# diff_376000_4961000# diff_3929000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2441 diff_3952000_5621000# diff_376000_4961000# diff_3957000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.19e+08 ps=90000 
M2442 diff_3972000_5587000# diff_376000_4961000# diff_3987000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.43e+08 ps=88000 
M2443 diff_4011000_5621000# diff_376000_4961000# diff_4017000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.04e+08 ps=88000 
M2444 diff_4031000_5587000# diff_376000_4961000# diff_4047000_4930000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=1.97e+08 ps=72000 
M2445 diff_4070000_5621000# diff_376000_4961000# diff_4075000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.27e+08 ps=88000 
M2446 diff_4090000_5587000# diff_376000_4961000# diff_4105000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.2e+08 ps=90000 
M2447 diff_4129000_5621000# diff_376000_4961000# diff_4135000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.2e+08 ps=86000 
M2448 diff_4149000_5587000# diff_376000_4961000# diff_4165000_4929000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.05e+08 ps=72000 
M2449 diff_4188000_5621000# diff_376000_4961000# diff_4193000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.28e+08 ps=90000 
M2450 diff_4208000_5587000# diff_376000_4961000# diff_4223000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.27e+08 ps=90000 
M2451 diff_4288000_5621000# diff_376000_4961000# diff_4293000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.04e+08 ps=88000 
M2452 diff_4307000_5587000# diff_376000_4961000# diff_4323000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.04e+08 ps=88000 
M2453 diff_4346000_5621000# diff_376000_4961000# diff_4351000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.27e+08 ps=88000 
M2454 diff_4366000_5587000# diff_376000_4961000# diff_4381000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2455 diff_4405000_5621000# diff_376000_4961000# diff_4411000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.13e+08 ps=88000 
M2456 diff_4425000_5587000# diff_376000_4961000# diff_4319000_4839000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.04e+08 ps=88000 
M2457 diff_4464000_5621000# diff_376000_4961000# diff_4469000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.18e+08 ps=90000 
M2458 diff_4484000_5587000# diff_376000_4961000# diff_4499000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.36e+08 ps=90000 
M2459 diff_4523000_5621000# diff_376000_4961000# diff_4529000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=6.98e+08 ps=286000 
M2460 diff_4543000_5587000# diff_376000_4961000# diff_4559000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2461 diff_4582000_5621000# diff_376000_4961000# diff_4587000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.27e+08 ps=90000 
M2462 diff_4602000_5587000# diff_376000_4961000# diff_4617000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.28e+08 ps=90000 
M2463 diff_4730000_5621000# diff_376000_4961000# diff_4735000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.27e+08 ps=88000 
M2464 diff_4750000_5587000# diff_376000_4961000# diff_4428000_3813000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.27e+08 ps=90000 
M2465 diff_4788000_5621000# diff_376000_4961000# diff_4770000_4458000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2466 diff_4808000_5587000# diff_376000_4961000# diff_4824000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M2467 diff_4847000_5621000# diff_376000_4961000# diff_4843000_4668000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.05e+08 ps=88000 
M2468 diff_4867000_5587000# diff_376000_4961000# diff_4883000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=4.47e+08 ps=152000 
M2469 diff_4906000_5621000# diff_376000_4961000# diff_4902000_4754000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=4.54e+08 ps=168000 
M2470 diff_4926000_5587000# diff_376000_4961000# diff_4920000_4772000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=1.338e+09 ps=354000 
M2471 diff_5004000_5621000# diff_376000_4961000# diff_5009000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.19e+08 ps=90000 
M2472 diff_5024000_5587000# diff_376000_4961000# diff_5039000_4962000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.28e+08 ps=90000 
M2473 diff_5062000_5621000# diff_376000_4961000# diff_5068000_4962000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.04e+08 ps=88000 
M2474 diff_5082000_5587000# diff_376000_4961000# diff_5098000_4894000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.04e+08 ps=70000 
M2475 diff_83000_3098000# diff_1233000_4962000# diff_94000_3158000# GND efet w=64000 l=8000
+ ad=0 pd=0 as=1.271e+09 ps=264000 
M2476 diff_807000_3040000# diff_1263000_4962000# diff_83000_3098000# GND efet w=64000 l=8000
+ ad=1.563e+09 pd=308000 as=0 ps=0 
M2477 diff_83000_3098000# diff_1292000_4962000# diff_991000_3076000# GND efet w=100000 l=7000
+ ad=0 pd=0 as=-1.83797e+09 ps=434000 
M2478 diff_94000_3158000# diff_94000_3158000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2479 diff_807000_3040000# diff_807000_3040000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2480 diff_1197000_3119000# diff_72000_4515000# diff_1200000_4480000# GND efet w=13000 l=12000
+ ad=-2.81967e+08 pd=806000 as=2.51e+08 ps=100000 
M2481 diff_1149000_4301000# diff_1126000_4459000# diff_83000_3098000# GND efet w=131000 l=8000
+ ad=1.747e+09 pd=320000 as=0 ps=0 
M2482 diff_1163000_4605000# diff_1145000_4574000# diff_1149000_4301000# GND efet w=130000 l=8000
+ ad=-4.69967e+08 pd=690000 as=0 ps=0 
M2483 diff_1195000_4346000# diff_1177000_4478000# diff_1163000_4605000# GND efet w=135000 l=8000
+ ad=1.359e+09 pd=292000 as=0 ps=0 
M2484 diff_83000_3098000# diff_1200000_4480000# diff_1195000_4346000# GND efet w=136000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2485 diff_1262000_4413000# diff_1253000_4407000# diff_1235000_4461000# GND efet w=131000 l=9000
+ ad=1.048e+09 pd=278000 as=-1.46997e+09 ps=578000 
M2486 diff_83000_3098000# diff_1204000_4962000# diff_1262000_4413000# GND efet w=131000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2487 diff_1448000_4598000# diff_1322000_4962000# diff_83000_3098000# GND efet w=64000 l=9000
+ ad=1.501e+09 pd=306000 as=0 ps=0 
M2488 diff_991000_3076000# diff_991000_3076000# diff_95000_5192000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M2489 diff_1235000_4461000# diff_1235000_4461000# diff_95000_5192000# GND efet w=13000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M2490 diff_1448000_4598000# diff_1448000_4598000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2491 diff_95000_5192000# diff_1180000_3099000# diff_1180000_3099000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=1.287e+09 ps=358000 
M2492 diff_680000_4314000# diff_68000_5288000# diff_997000_3891000# GND efet w=13000 l=13000
+ ad=-1.92897e+09 pd=564000 as=2.42e+08 ps=94000 
M2493 diff_873000_3938000# diff_72000_4515000# diff_929000_3956000# GND efet w=14000 l=11000
+ ad=5.90327e+07 pd=852000 as=2.72e+08 ps=92000 
M2494 diff_792000_3825000# diff_68000_5288000# diff_752000_3797000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=2.04e+08 ps=78000 
M2495 diff_95000_5192000# diff_792000_3825000# diff_792000_3825000# GND efet w=11000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2496 diff_732000_3738000# diff_732000_3738000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2497 diff_101000_3535000# diff_94000_3551000# diff_83000_3098000# GND efet w=121500 l=8500
+ ad=-3.52967e+08 pd=656000 as=0 ps=0 
M2498 diff_95000_5192000# diff_101000_3535000# diff_101000_3535000# GND efet w=13000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M2499 diff_83000_3098000# diff_124000_3549000# diff_101000_3535000# GND efet w=111000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2500 diff_83000_3098000# diff_608000_3765000# diff_570000_3597000# GND efet w=81000 l=8000
+ ad=0 pd=0 as=-9.52967e+08 ps=660000 
M2501 diff_83000_3098000# diff_94000_3551000# diff_635000_3800000# GND efet w=64000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2502 diff_95000_5192000# diff_230000_4601000# diff_230000_4601000# GND efet w=11000 l=22000
+ ad=0 pd=0 as=1.325e+09 ps=282000 
M2503 diff_101000_3535000# diff_88000_3357000# diff_83000_3098000# GND efet w=102000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2504 diff_101000_3535000# diff_72000_4515000# diff_104000_3496000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=3.11e+08 ps=96000 
M2505 diff_124000_3549000# diff_72000_4515000# diff_104000_3450000# GND efet w=20000 l=13000
+ ad=2.82e+08 pd=100000 as=-1.18597e+09 ps=564000 
M2506 diff_83000_3098000# diff_104000_3496000# diff_104000_3450000# GND efet w=105500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2507 diff_83000_3098000# diff_111000_3412000# diff_104000_3450000# GND efet w=126500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2508 diff_95000_5192000# diff_104000_3450000# diff_104000_3450000# GND efet w=13000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M2509 diff_74000_3122000# diff_104000_3450000# diff_83000_3098000# GND efet w=115000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2510 diff_95000_5192000# diff_74000_3122000# diff_74000_3122000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M2511 diff_83000_3098000# diff_94000_3551000# diff_570000_3597000# GND efet w=79000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2512 diff_792000_3825000# diff_787000_3667000# diff_83000_3098000# GND efet w=69000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2513 diff_1163000_4605000# diff_1163000_4605000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2514 diff_83000_3098000# diff_886000_3953000# diff_873000_3938000# GND efet w=40000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2515 diff_680000_4314000# diff_929000_3956000# diff_83000_3098000# GND efet w=70000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2516 diff_936000_4586000# diff_72000_4515000# diff_1055000_3959000# GND efet w=14000 l=12000
+ ad=0 pd=0 as=2.71e+08 ps=94000 
M2517 diff_975000_4364000# diff_72000_4515000# diff_1079000_3958000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.42e+08 ps=94000 
M2518 diff_987000_3874000# diff_997000_3891000# diff_83000_3098000# GND efet w=65000 l=9000
+ ad=1.326e+09 pd=294000 as=0 ps=0 
M2519 diff_1029000_3949000# diff_72000_4515000# diff_987000_3874000# GND efet w=14000 l=11000
+ ad=3.89e+08 pd=116000 as=0 ps=0 
M2520 diff_1053000_4267000# diff_72000_4515000# diff_1134000_3807000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=3.03e+08 ps=92000 
M2521 diff_1076000_4557000# diff_72000_4515000# diff_1152000_3809000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.44e+08 ps=82000 
M2522 diff_873000_3938000# diff_873000_3938000# diff_95000_5192000# GND efet w=12000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M2523 diff_987000_3874000# diff_987000_3874000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2524 diff_680000_4314000# diff_680000_4314000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2525 diff_787000_3667000# diff_72000_4515000# diff_784000_3633000# GND efet w=12000 l=12000
+ ad=2.34e+08 pd=78000 as=2.22033e+08 ps=810000 
M2526 diff_792000_3825000# diff_68000_5288000# diff_731000_3544000# GND efet w=13000 l=13000
+ ad=0 pd=0 as=2.56e+08 ps=92000 
M2527 diff_83000_3098000# diff_94000_3158000# diff_230000_4601000# GND efet w=67000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2528 diff_1048000_3792000# diff_1029000_3949000# diff_691000_4135000# GND efet w=131000 l=8000
+ ad=1.31e+09 pd=282000 as=-2.07297e+09 ps=440000 
M2529 diff_83000_3098000# diff_1055000_3959000# diff_1048000_3792000# GND efet w=131000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M2530 diff_637000_4100000# diff_1079000_3958000# diff_83000_3098000# GND efet w=64000 l=8000
+ ad=1.744e+09 pd=338000 as=0 ps=0 
M2531 diff_637000_4100000# diff_637000_4100000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2532 diff_1142000_3814000# diff_1134000_3807000# diff_659000_4117000# GND efet w=132000 l=8000
+ ad=1.32e+09 pd=284000 as=-1.46197e+09 ps=606000 
M2533 diff_83000_3098000# diff_1152000_3809000# diff_1142000_3814000# GND efet w=132000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2534 diff_659000_4117000# diff_659000_4117000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2535 diff_95000_5192000# diff_691000_4135000# diff_691000_4135000# GND efet w=11000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2536 diff_635000_3800000# diff_68000_5288000# diff_906000_3511000# GND efet w=20000 l=12000
+ ad=0 pd=0 as=3.12e+08 ps=106000 
M2537 diff_111000_3412000# diff_68000_5288000# diff_111000_3358000# GND efet w=21000 l=12000
+ ad=3.05e+08 pd=96000 as=-7.49673e+07 ps=658000 
M2538 diff_128000_3343000# diff_206000_3372000# diff_83000_3098000# GND efet w=84500 l=8500
+ ad=1.14e+09 pd=224000 as=0 ps=0 
M2539 diff_235000_3317000# diff_72000_4515000# diff_206000_3372000# GND efet w=14000 l=12000
+ ad=0 pd=0 as=2.49e+08 ps=80000 
M2540 diff_83000_3098000# diff_128000_3343000# diff_111000_3358000# GND efet w=110000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2541 diff_95000_5192000# diff_128000_3343000# diff_128000_3343000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2542 diff_95000_5192000# diff_111000_3358000# diff_111000_3358000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M2543 diff_111000_3358000# diff_88000_3357000# diff_83000_3098000# GND efet w=103000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2544 diff_111000_3358000# diff_235000_3317000# diff_83000_3098000# GND efet w=100000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2545 diff_83000_3098000# diff_731000_3544000# diff_169000_4545000# GND efet w=126000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2546 diff_95000_5192000# diff_65000_4220000# diff_65000_4220000# GND efet w=16000 l=8000
+ ad=0 pd=0 as=9.39033e+08 ps=1.06e+06 
M2547 diff_65000_4220000# diff_906000_3511000# diff_83000_3098000# GND efet w=255000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2548 diff_1581000_4325000# diff_860000_2987000# diff_83000_3098000# GND efet w=116000 l=8000
+ ad=-1.4349e+09 pd=1.906e+06 as=0 ps=0 
M2549 diff_83000_3098000# diff_1410000_4962000# diff_1541000_4610000# GND efet w=41000 l=10000
+ ad=0 pd=0 as=-1.64797e+09 ps=428000 
M2550 diff_1541000_4610000# diff_1440000_4962000# diff_83000_3098000# GND efet w=41000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2551 diff_83000_3098000# diff_1469000_4962000# diff_1541000_4610000# GND efet w=44000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2552 diff_83000_3098000# diff_1674000_4606000# diff_1581000_4325000# GND efet w=100000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2553 diff_1541000_4610000# diff_1541000_4610000# diff_95000_5192000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M2554 diff_83000_3098000# diff_1448000_4598000# diff_1180000_3099000# GND efet w=70000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2555 diff_169000_4545000# diff_169000_4545000# diff_95000_5192000# GND efet w=11000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M2556 diff_570000_3597000# diff_570000_3597000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2557 diff_88000_3357000# diff_68000_5288000# diff_90000_3265000# GND efet w=14000 l=12000
+ ad=2.59e+08 pd=84000 as=1.991e+09 ps=396000 
M2558 diff_90000_3265000# diff_111000_3254000# diff_83000_3098000# GND efet w=85000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2559 diff_95000_5192000# diff_90000_3265000# diff_90000_3265000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2560 diff_102000_3167000# diff_72000_4515000# diff_111000_3254000# GND efet w=12000 l=11000
+ ad=-1.14897e+09 pd=576000 as=2.68e+08 ps=86000 
M2561 diff_102000_3167000# diff_94000_3158000# diff_83000_3148000# GND efet w=213500 l=8500
+ ad=0 pd=0 as=-1.92997e+09 ps=486000 
M2562 diff_95000_5192000# diff_102000_3167000# diff_102000_3167000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2563 diff_83000_3148000# diff_65000_4220000# diff_83000_3131000# GND efet w=198000 l=8000
+ ad=0 pd=0 as=1.782e+09 ps=414000 
M2564 diff_83000_3131000# diff_74000_3122000# diff_83000_3098000# GND efet w=198000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2565 diff_83000_3098000# diff_534000_2989000# diff_519000_3032000# GND efet w=142000 l=8000
+ ad=0 pd=0 as=-1.50097e+09 ps=732000 
M2566 diff_519000_3032000# diff_519000_3032000# diff_95000_5192000# GND efet w=12000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M2567 diff_557000_2988000# diff_68000_5288000# diff_534000_2989000# GND efet w=13000 l=11000
+ ad=-1.85397e+09 pd=462000 as=5e+08 ps=146000 
M2568 diff_95000_5192000# diff_1595000_4502000# diff_1595000_4502000# GND efet w=13000 l=36000
+ ad=0 pd=0 as=1.276e+09 ps=250000 
M2569 diff_1549000_4377000# diff_1523000_4349000# diff_83000_3098000# GND efet w=103500 l=8500
+ ad=9.31e+08 pd=224000 as=0 ps=0 
M2570 diff_856000_3301000# diff_1381000_4962000# diff_1549000_4377000# GND efet w=103500 l=8500
+ ad=-1.55597e+09 pd=516000 as=0 ps=0 
M2571 diff_1595000_4502000# diff_1541000_4610000# diff_83000_3098000# GND efet w=60500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2572 diff_1740000_4513000# diff_1692000_4497000# diff_83000_3098000# GND efet w=199500 l=7500
+ ad=2.042e+09 pd=432000 as=0 ps=0 
M2573 diff_1000000_2990000# diff_68000_5288000# diff_1692000_4497000# GND efet w=13000 l=10000
+ ad=1.96503e+09 pd=1.336e+06 as=3e+08 ps=96000 
M2574 diff_83000_3098000# diff_640000_3020000# diff_557000_2988000# GND efet w=75000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2575 diff_667000_3269000# diff_669000_2930000# diff_83000_3098000# GND efet w=198000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2576 diff_83000_3098000# diff_687000_3101000# diff_667000_3269000# GND efet w=218500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2577 diff_1523000_4349000# diff_72000_4515000# diff_1477000_3932000# GND efet w=12000 l=12000
+ ad=3.6e+08 pd=102000 as=-1.94897e+09 ps=512000 
M2578 diff_1581000_4325000# diff_1581000_4325000# diff_95000_5192000# GND efet w=13000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M2579 diff_1406000_3519000# diff_72000_4515000# diff_531000_4622000# GND efet w=13000 l=11000
+ ad=1.281e+09 pd=332000 as=0 ps=0 
M2580 diff_1419000_3778000# diff_1351000_4962000# diff_83000_3098000# GND efet w=147000 l=8000
+ ad=1.431e+09 pd=314000 as=0 ps=0 
M2581 diff_1436000_3778000# diff_1406000_3519000# diff_1419000_3778000# GND efet w=148000 l=8000
+ ad=-2.09997e+09 pd=500000 as=0 ps=0 
M2582 diff_856000_3301000# diff_856000_3301000# diff_95000_5192000# GND efet w=11000 l=27000
+ ad=0 pd=0 as=0 ps=0 
M2583 diff_1581000_4325000# diff_1469000_4962000# diff_1740000_4513000# GND efet w=204000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2584 diff_1691000_4259000# diff_1595000_4502000# diff_83000_3098000# GND efet w=223500 l=8500
+ ad=-1.83097e+09 pd=466000 as=0 ps=0 
M2585 diff_1508000_3890000# diff_1237000_3461000# diff_1477000_3932000# GND efet w=101000 l=8000
+ ad=8.57e+08 pd=218000 as=0 ps=0 
M2586 diff_83000_3098000# diff_1516000_3900000# diff_1508000_3890000# GND efet w=100500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M2587 diff_1339000_3691000# diff_72000_4515000# diff_1235000_4461000# GND efet w=11000 l=11000
+ ad=4.13e+08 pd=130000 as=0 ps=0 
M2588 diff_687000_3101000# diff_100000_3992000# diff_83000_3098000# GND efet w=91500 l=8500
+ ad=-2.00897e+09 pd=424000 as=0 ps=0 
M2589 diff_1000000_2990000# diff_68000_5288000# diff_1272000_3500000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.71e+08 ps=98000 
M2590 diff_1237000_3461000# diff_1272000_3500000# diff_83000_3098000# GND efet w=47000 l=8000
+ ad=1.194e+09 pd=252000 as=0 ps=0 
M2591 diff_856000_3301000# diff_68000_5288000# diff_823000_3289000# GND efet w=13000 l=11000
+ ad=0 pd=0 as=3.63e+08 ps=114000 
M2592 diff_1237000_3461000# diff_1237000_3461000# diff_95000_5192000# GND efet w=11000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M2593 diff_95000_5192000# diff_1000000_2990000# diff_1000000_2990000# GND efet w=11000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M2594 diff_1000000_2990000# diff_1339000_3691000# diff_83000_3098000# GND efet w=145000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2595 diff_95000_5192000# diff_1436000_3778000# diff_1436000_3778000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2596 diff_597000_3013000# diff_94000_3551000# diff_83000_3098000# GND efet w=162000 l=8000
+ ad=1.09303e+09 pd=900000 as=0 ps=0 
M2597 diff_640000_3020000# diff_72000_4515000# diff_597000_3013000# GND efet w=12000 l=11000
+ ad=3.17e+08 pd=92000 as=0 ps=0 
M2598 diff_95000_5192000# diff_557000_2988000# diff_557000_2988000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2599 diff_83000_3098000# diff_94000_3158000# diff_743000_2974000# GND efet w=83000 l=8000
+ ad=0 pd=0 as=1.521e+09 ps=300000 
M2600 diff_687000_3101000# diff_687000_3101000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2601 diff_815000_3048000# diff_807000_3040000# diff_597000_3013000# GND efet w=336500 l=8500
+ ad=-1.04597e+09 pd=692000 as=0 ps=0 
M2602 diff_83000_3098000# diff_823000_3289000# diff_815000_3048000# GND efet w=336500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2603 diff_1477000_3932000# diff_1477000_3932000# diff_95000_5192000# GND efet w=13000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M2604 diff_1581000_4325000# diff_1483000_3488000# diff_1691000_4259000# GND efet w=216500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2605 diff_83000_3098000# diff_1276000_3285000# diff_625000_4565000# GND efet w=133500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M2606 diff_1966000_4584000# diff_1713000_4962000# diff_83000_3098000# GND efet w=42000 l=9000
+ ad=1.143e+09 pd=258000 as=0 ps=0 
M2607 diff_83000_3098000# diff_1742000_4962000# diff_2005000_4584000# GND efet w=67500 l=8500
+ ad=0 pd=0 as=1.02e+09 ps=256000 
M2608 diff_1674000_4606000# diff_2005000_4584000# diff_83000_3098000# GND efet w=68000 l=8000
+ ad=1.608e+09 pd=310000 as=0 ps=0 
M2609 diff_83000_3098000# diff_1772000_4962000# diff_1674000_4606000# GND efet w=65000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2610 diff_625000_4565000# diff_625000_4565000# diff_95000_5192000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M2611 diff_1966000_4584000# diff_1966000_4584000# diff_95000_5192000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M2612 diff_2005000_4584000# diff_2005000_4584000# diff_95000_5192000# GND efet w=11000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M2613 diff_83000_3098000# diff_686000_4521000# diff_1581000_4325000# GND efet w=97000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M2614 diff_1516000_3900000# diff_1499000_4962000# diff_83000_3098000# GND efet w=67000 l=8000
+ ad=1.284e+09 pd=276000 as=0 ps=0 
M2615 diff_83000_3098000# diff_1528000_4962000# diff_1516000_3900000# GND efet w=76500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2616 diff_1516000_3900000# diff_1516000_3900000# diff_95000_5192000# GND efet w=11000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2617 diff_1163000_4605000# diff_68000_5288000# diff_1589000_4012000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.74e+08 ps=96000 
M2618 diff_1097000_3119000# diff_1589000_4012000# diff_83000_3098000# GND efet w=112000 l=8000
+ ad=-2.08397e+09 pd=482000 as=0 ps=0 
M2619 diff_83000_3098000# diff_94000_3551000# diff_1097000_3119000# GND efet w=114500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M2620 diff_1197000_3119000# diff_1516000_3900000# diff_83000_3098000# GND efet w=221000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2621 diff_1581000_4325000# diff_72000_4515000# diff_1741000_4000000# GND efet w=14000 l=10000
+ ad=0 pd=0 as=2.56e+08 ps=94000 
M2622 diff_1097000_3119000# diff_1097000_3119000# diff_95000_5192000# GND efet w=13000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M2623 diff_83000_3098000# diff_1713000_3885000# diff_1646000_3414000# GND efet w=110000 l=8000
+ ad=0 pd=0 as=2.17033e+08 ps=862000 
M2624 diff_1713000_3885000# diff_1741000_4000000# diff_83000_3098000# GND efet w=64000 l=9000
+ ad=1.561e+09 pd=340000 as=0 ps=0 
M2625 diff_83000_3098000# diff_94000_3551000# diff_1713000_3885000# GND efet w=82000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2626 diff_1436000_3778000# diff_68000_5288000# diff_1459000_3632000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.43e+08 ps=86000 
M2627 diff_95000_5192000# diff_946000_3261000# diff_946000_3261000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=-1.94897e+09 ps=552000 
M2628 diff_946000_3261000# diff_1459000_3632000# diff_83000_3098000# GND efet w=105500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M2629 diff_1197000_3119000# diff_1197000_3119000# diff_95000_5192000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2630 diff_83000_3098000# diff_94000_3551000# diff_1406000_3519000# GND efet w=68000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2631 diff_95000_5192000# diff_1561000_3639000# diff_1561000_3639000# GND efet w=11000 l=35000
+ ad=0 pd=0 as=1.525e+09 ps=314000 
M2632 diff_1713000_3885000# diff_1713000_3885000# diff_95000_5192000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2633 diff_1097000_3119000# diff_72000_4515000# diff_1539000_3467000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=9.77e+08 ps=238000 
M2634 diff_95000_5192000# diff_100000_3992000# diff_100000_3992000# GND efet w=15000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M2635 diff_1646000_3414000# diff_92000_3714000# diff_83000_3098000# GND efet w=100000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2636 diff_95000_5192000# diff_1483000_3488000# diff_1483000_3488000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=1.423e+09 ps=282000 
M2637 diff_83000_3098000# diff_1539000_3467000# diff_1561000_3639000# GND efet w=46000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M2638 diff_1561000_3639000# diff_68000_5288000# diff_1475000_3480000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=2.87e+08 ps=96000 
M2639 diff_1483000_3488000# diff_1475000_3480000# diff_83000_3098000# GND efet w=69000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2640 diff_83000_3098000# diff_1622000_3414000# diff_100000_3992000# GND efet w=211500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2641 diff_1674000_4606000# diff_1674000_4606000# diff_95000_5192000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2642 diff_1000000_2990000# diff_68000_5288000# diff_2060000_4467000# GND efet w=13000 l=13000
+ ad=0 pd=0 as=2.27e+08 ps=88000 
M2643 diff_83000_3098000# diff_1801000_4962000# diff_2063000_4304000# GND efet w=63000 l=8000
+ ad=0 pd=0 as=-1.68197e+09 ps=558000 
M2644 diff_83000_3098000# diff_2187000_4495000# diff_791000_4022000# GND efet w=307000 l=8000
+ ad=0 pd=0 as=6.77098e+08 ps=2.446e+06 
M2645 diff_83000_3098000# diff_2007000_4962000# diff_2187000_4495000# GND efet w=110000 l=9000
+ ad=0 pd=0 as=1.78503e+09 ps=1.122e+06 
M2646 diff_2187000_4495000# diff_2037000_4962000# diff_83000_3098000# GND efet w=113000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2647 diff_791000_4022000# diff_2067000_4962000# diff_83000_3098000# GND efet w=315000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2648 diff_83000_3098000# diff_2097000_4962000# diff_791000_4022000# GND efet w=315000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2649 diff_791000_4022000# diff_2125000_4962000# diff_83000_3098000# GND efet w=322500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2650 diff_83000_3098000# diff_94000_3551000# diff_791000_4022000# GND efet w=325000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2651 diff_2063000_4304000# diff_2060000_4467000# diff_83000_3098000# GND efet w=66000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2652 diff_83000_3098000# diff_1483000_3488000# diff_2063000_4304000# GND efet w=66000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2653 diff_2063000_4304000# diff_2063000_4304000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2654 diff_1902000_3917000# diff_1655000_4962000# diff_83000_3098000# GND efet w=131000 l=8000
+ ad=1.31e+09 pd=282000 as=0 ps=0 
M2655 diff_1276000_3285000# diff_531000_4622000# diff_1902000_3917000# GND efet w=131000 l=8000
+ ad=1.53707e+09 pd=1.806e+06 as=0 ps=0 
M2656 diff_2187000_4495000# diff_2194000_4240000# diff_83000_3098000# GND efet w=108000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2657 diff_2173000_3038000# diff_2135000_4721000# diff_83000_3098000# GND efet w=66500 l=8500
+ ad=1.00033e+08 pd=822000 as=0 ps=0 
M2658 diff_2173000_3038000# diff_2371000_4962000# diff_83000_3098000# GND efet w=64500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M2659 diff_791000_4022000# diff_791000_4022000# diff_95000_5192000# GND efet w=26000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M2660 diff_83000_3098000# diff_2155000_4962000# diff_2405000_4387000# GND efet w=44500 l=8500
+ ad=0 pd=0 as=-2.07997e+09 ps=522000 
M2661 diff_2566000_3500000# diff_2488000_4962000# diff_83000_3098000# GND efet w=78000 l=8000
+ ad=-9.39673e+07 pd=762000 as=0 ps=0 
M2662 diff_83000_3098000# diff_2518000_4962000# diff_2566000_3500000# GND efet w=65000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2663 diff_2173000_3038000# diff_2341000_4962000# diff_83000_3098000# GND efet w=66500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2664 diff_2198000_3000000# diff_2282000_4962000# diff_83000_3098000# GND efet w=69000 l=9000
+ ad=1.274e+09 pd=272000 as=0 ps=0 
M2665 diff_2405000_4387000# diff_2223000_4962000# diff_83000_3098000# GND efet w=43000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2666 diff_83000_3098000# diff_2253000_4962000# diff_2405000_4387000# GND efet w=44500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2667 diff_83000_3098000# diff_2312000_4962000# diff_2198000_3000000# GND efet w=69000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2668 diff_2187000_4495000# diff_2187000_4495000# diff_95000_5192000# GND efet w=13000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M2669 diff_1976000_3921000# diff_1953000_3750000# diff_83000_3098000# GND efet w=196000 l=9000
+ ad=1.764e+09 pd=410000 as=0 ps=0 
M2670 diff_1993000_3921000# diff_1625000_4962000# diff_1976000_3921000# GND efet w=196000 l=8000
+ ad=1.764e+09 pd=410000 as=0 ps=0 
M2671 diff_1465000_3204000# diff_1966000_4584000# diff_1993000_3921000# GND efet w=196000 l=9000
+ ad=6.11033e+08 pd=1e+06 as=0 ps=0 
M2672 diff_1646000_3414000# diff_1646000_3414000# diff_95000_5192000# GND efet w=13000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M2673 diff_1276000_3285000# diff_1276000_3285000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2674 diff_95000_5192000# diff_512000_4352000# diff_512000_4352000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=1.855e+09 ps=450000 
M2675 diff_1944000_3756000# diff_1683000_4962000# diff_1276000_3285000# GND efet w=143500 l=8500
+ ad=1.296e+09 pd=306000 as=0 ps=0 
M2676 diff_83000_3098000# diff_1953000_3750000# diff_1944000_3756000# GND efet w=144000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2677 diff_2093000_3973000# diff_1483000_3488000# diff_83000_3098000# GND efet w=211000 l=8000
+ ad=2.038e+09 pd=440000 as=0 ps=0 
M2678 diff_2111000_3992000# diff_1831000_4962000# diff_2093000_3973000# GND efet w=210000 l=8000
+ ad=1.98e+09 pd=440000 as=0 ps=0 
M2679 diff_2129000_4009000# diff_2120000_4001000# diff_2111000_3992000# GND efet w=210500 l=8500
+ ad=2.03203e+09 pd=1.092e+06 as=0 ps=0 
M2680 diff_2194000_4240000# diff_68000_5288000# diff_2222000_4172000# GND efet w=20000 l=12000
+ ad=3.6e+08 pd=90000 as=-1.95897e+09 ps=440000 
M2681 diff_2154000_3995000# diff_531000_4622000# diff_2129000_4009000# GND efet w=147500 l=8500
+ ad=-5.29673e+07 pd=634000 as=0 ps=0 
M2682 diff_83000_3098000# diff_1949000_4962000# diff_2154000_3995000# GND efet w=131000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2683 diff_2154000_3995000# diff_1979000_4962000# diff_83000_3098000# GND efet w=146000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2684 diff_773000_4078000# diff_1001000_4394000# diff_83000_3098000# GND efet w=63000 l=8000
+ ad=1.407e+09 pd=330000 as=0 ps=0 
M2685 diff_2405000_4387000# diff_2405000_4387000# diff_95000_5192000# GND efet w=13000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M2686 diff_2198000_3000000# diff_2198000_3000000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2687 diff_2568000_4388000# diff_2399000_4962000# diff_2173000_3038000# GND efet w=131000 l=9000
+ ad=1.179e+09 pd=280000 as=0 ps=0 
M2688 diff_83000_3098000# diff_531000_4622000# diff_2568000_4388000# GND efet w=131000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2689 diff_773000_4078000# diff_773000_4078000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2690 diff_2063000_4304000# diff_72000_4515000# diff_2256000_3932000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.35e+08 ps=88000 
M2691 diff_791000_4022000# diff_72000_4515000# diff_2337000_4018000# GND efet w=14000 l=12000
+ ad=0 pd=0 as=3.42e+08 ps=104000 
M2692 diff_2173000_3038000# diff_2173000_3038000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2693 diff_83000_3098000# diff_2256000_3932000# diff_2222000_4172000# GND efet w=78000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2694 diff_83000_3098000# diff_2063000_4304000# diff_1953000_3750000# GND efet w=68000 l=8000
+ ad=0 pd=0 as=-2.00197e+09 ps=450000 
M2695 diff_2324000_3768000# diff_2337000_4018000# diff_83000_3098000# GND efet w=64500 l=8500
+ ad=1.812e+09 pd=396000 as=0 ps=0 
M2696 diff_2073000_3806000# diff_68000_5288000# diff_2050000_3807000# GND efet w=12000 l=11000
+ ad=4.59e+08 pd=136000 as=-1.37097e+09 ps=550000 
M2697 diff_1465000_3204000# diff_1465000_3204000# diff_95000_5192000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2698 diff_83000_3098000# diff_1557000_4962000# diff_512000_4352000# GND efet w=64000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M2699 diff_83000_3098000# diff_94000_3551000# diff_1539000_3467000# GND efet w=26000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2700 diff_946000_3261000# diff_72000_4515000# diff_946000_3225000# GND efet w=14000 l=12000
+ ad=0 pd=0 as=3.45e+08 ps=108000 
M2701 diff_906000_3226000# diff_72000_4515000# diff_917000_3186000# GND efet w=13000 l=12000
+ ad=-7.37967e+08 pd=726000 as=2.58e+08 ps=88000 
M2702 diff_1834000_3561000# diff_791000_4022000# diff_83000_3098000# GND efet w=130000 l=8000
+ ad=1.17e+09 pd=278000 as=0 ps=0 
M2703 diff_1276000_3285000# diff_1625000_4962000# diff_1834000_3561000# GND efet w=130000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2704 diff_1276000_3285000# diff_1097000_3119000# diff_83000_3098000# GND efet w=63000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2705 diff_83000_3098000# diff_1197000_3119000# diff_1276000_3285000# GND efet w=62000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2706 diff_83000_3098000# diff_875000_3125000# diff_860000_2987000# GND efet w=122000 l=9000
+ ad=0 pd=0 as=-1.12097e+09 ps=576000 
M2707 diff_95000_5192000# diff_667000_3269000# diff_667000_3269000# GND efet w=16000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2708 diff_743000_2974000# diff_743000_2974000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2709 diff_597000_3013000# diff_597000_3013000# diff_95000_5192000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2710 diff_912000_3048000# diff_917000_3186000# diff_83000_3098000# GND efet w=85500 l=8500
+ ad=-1.66697e+09 pd=504000 as=0 ps=0 
M2711 diff_962000_3082000# diff_946000_3225000# diff_912000_3048000# GND efet w=131000 l=8000
+ ad=1.31e+09 pd=282000 as=0 ps=0 
M2712 diff_83000_3098000# diff_512000_4352000# diff_962000_3082000# GND efet w=131000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2713 diff_967000_2989000# diff_991000_3076000# diff_83000_3098000# GND efet w=93500 l=8500
+ ad=-1.35697e+09 pd=506000 as=0 ps=0 
M2714 diff_912000_3048000# diff_68000_5288000# diff_875000_3125000# GND efet w=13000 l=11000
+ ad=0 pd=0 as=2.82e+08 ps=78000 
M2715 diff_860000_2987000# diff_860000_2987000# diff_95000_5192000# GND efet w=13000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M2716 diff_95000_5192000# diff_669000_2930000# diff_669000_2930000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=1.699e+09 ps=320000 
M2717 diff_669000_2930000# diff_337000_4528000# diff_83000_3098000# GND efet w=127500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2718 diff_912000_3048000# diff_912000_3048000# diff_95000_5192000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2719 diff_83000_3098000# diff_1048000_3119000# diff_1028000_3008000# GND efet w=76000 l=9000
+ ad=0 pd=0 as=-1.77897e+09 ps=552000 
M2720 diff_83000_3098000# diff_1097000_3119000# diff_1048000_3119000# GND efet w=100000 l=8000
+ ad=0 pd=0 as=2.01065e+08 ps=1.514e+06 
M2721 diff_1048000_3119000# diff_65000_4220000# diff_83000_3098000# GND efet w=95000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M2722 diff_83000_3098000# diff_1148000_3109000# diff_1048000_3119000# GND efet w=117500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M2723 diff_1028000_3008000# diff_1028000_3008000# diff_95000_5192000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2724 diff_967000_2989000# diff_967000_2989000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2725 diff_83000_3098000# diff_967000_2989000# diff_1048000_3119000# GND efet w=100000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2726 diff_1188000_3107000# diff_1180000_3099000# diff_83000_3098000# GND efet w=65000 l=8000
+ ad=2.07033e+08 pd=752000 as=0 ps=0 
M2727 diff_83000_3098000# diff_1197000_3119000# diff_1188000_3107000# GND efet w=93000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2728 diff_1276000_3285000# diff_72000_4515000# diff_1276000_3249000# GND efet w=14000 l=12000
+ ad=0 pd=0 as=2.72e+08 ps=92000 
M2729 diff_1646000_3414000# diff_68000_5288000# diff_1622000_3414000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=6.6e+08 ps=168000 
M2730 diff_83000_3098000# diff_169000_4545000# diff_1276000_3285000# GND efet w=65000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2731 diff_1979000_3617000# diff_1502000_2925000# diff_1556000_2817000# GND efet w=221000 l=8000
+ ad=2.061e+09 pd=488000 as=-1.09997e+09 ps=580000 
M2732 diff_83000_3098000# diff_1659000_2818000# diff_1979000_3617000# GND efet w=218000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2733 diff_2129000_4009000# diff_2129000_4009000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2734 diff_2222000_4172000# diff_2222000_4172000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2735 diff_2182000_3681000# diff_2174000_3677000# diff_2129000_4009000# GND efet w=130000 l=8000
+ ad=5.37033e+08 pd=794000 as=0 ps=0 
M2736 diff_2324000_3768000# diff_2324000_3768000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2737 diff_1953000_3750000# diff_1953000_3750000# diff_95000_5192000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2738 diff_2174000_3677000# diff_2174000_3677000# diff_95000_5192000# GND efet w=12000 l=37000
+ ad=2.02e+09 pd=414000 as=0 ps=0 
M2739 diff_2647000_4397000# diff_2429000_4962000# diff_83000_3098000# GND efet w=131000 l=8000
+ ad=1.31e+09 pd=282000 as=0 ps=0 
M2740 diff_2566000_3500000# diff_1253000_4407000# diff_2647000_4397000# GND efet w=131000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2741 diff_2642000_3475000# diff_2636000_4962000# diff_83000_3098000# GND efet w=42000 l=9000
+ ad=1.034e+09 pd=220000 as=0 ps=0 
M2742 diff_2642000_3475000# diff_2642000_3475000# diff_95000_5192000# GND efet w=12000 l=35000
+ ad=0 pd=0 as=0 ps=0 
M2743 diff_2687000_4368000# diff_2547000_4962000# diff_2566000_3500000# GND efet w=133500 l=8500
+ ad=1.188e+09 pd=284000 as=0 ps=0 
M2744 diff_83000_3098000# diff_531000_4622000# diff_2687000_4368000# GND efet w=132500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2745 diff_773000_4078000# diff_72000_4515000# diff_2471000_3862000# GND efet w=13000 l=13000
+ ad=0 pd=0 as=2.49e+08 ps=92000 
M2746 diff_2405000_4387000# diff_72000_4515000# diff_2490000_3879000# GND efet w=13000 l=13000
+ ad=0 pd=0 as=4.84e+08 ps=122000 
M2747 diff_2566000_3500000# diff_2566000_3500000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2748 diff_2050000_3807000# diff_2471000_3862000# diff_83000_3098000# GND efet w=66000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2749 diff_83000_3098000# diff_2490000_3879000# diff_2050000_3807000# GND efet w=78000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2750 diff_2135000_4721000# diff_2509000_3809000# diff_83000_3098000# GND efet w=74000 l=8000
+ ad=2.142e+09 pd=392000 as=0 ps=0 
M2751 diff_2915000_4682000# diff_2906000_4658000# diff_2878000_4622000# GND efet w=86000 l=9000
+ ad=6.88e+08 pd=188000 as=-2.02097e+09 ps=532000 
M2752 diff_83000_3098000# diff_2762000_4962000# diff_2915000_4682000# GND efet w=86000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2753 diff_2931000_4557000# diff_2792000_4962000# diff_83000_3098000# GND efet w=64000 l=7000
+ ad=-1.45197e+09 pd=560000 as=0 ps=0 
M2754 diff_83000_3098000# diff_2821000_4962000# diff_2931000_4557000# GND efet w=66500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2755 diff_2878000_4622000# diff_2878000_4622000# diff_95000_5192000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M2756 diff_95000_5192000# diff_2860000_4570000# diff_2860000_4570000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=1.362e+09 ps=322000 
M2757 diff_83000_3098000# diff_2971000_4656000# diff_2931000_4557000# GND efet w=68000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2758 diff_95000_5192000# diff_2931000_4557000# diff_2931000_4557000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2759 diff_3009000_4523000# diff_2880000_4962000# diff_83000_3098000# GND efet w=70500 l=8500
+ ad=-1.51597e+09 pd=598000 as=0 ps=0 
M2760 diff_3062000_4310000# diff_2910000_4962000# diff_3009000_4523000# GND efet w=134500 l=8500
+ ad=-8.82967e+08 pd=604000 as=0 ps=0 
M2761 diff_83000_3098000# diff_2877000_4437000# diff_2860000_4570000# GND efet w=85000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2762 diff_2877000_4437000# diff_72000_4515000# diff_2913000_4304000# GND efet w=12000 l=11000
+ ad=2.51e+08 pd=80000 as=-2.03397e+09 ps=472000 
M2763 diff_95000_5192000# diff_3009000_4523000# diff_3009000_4523000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2764 diff_2906000_4658000# diff_72000_4515000# diff_530000_4372000# GND efet w=13000 l=9000
+ ad=1.88e+09 pd=392000 as=7.85033e+08 ps=974000 
M2765 diff_2895000_4350000# diff_2694000_4962000# diff_83000_3098000# GND efet w=108500 l=8500
+ ad=1.029e+09 pd=236000 as=0 ps=0 
M2766 diff_2913000_4304000# diff_1001000_4394000# diff_2895000_4350000# GND efet w=87000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2767 diff_83000_3098000# diff_94000_3551000# diff_2906000_4658000# GND efet w=72000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M2768 diff_83000_3098000# diff_2570000_3912000# diff_2559000_3889000# GND efet w=146500 l=8500
+ ad=0 pd=0 as=-1.00693e+09 ps=1.318e+06 
M2769 diff_2559000_3889000# diff_946000_3261000# diff_83000_3098000# GND efet w=128500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M2770 diff_83000_3098000# diff_531000_4622000# diff_2559000_3889000# GND efet w=145500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2771 diff_2559000_3889000# diff_530000_4372000# diff_83000_3098000# GND efet w=139000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2772 diff_2913000_4304000# diff_2913000_4304000# diff_95000_5192000# GND efet w=11000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M2773 diff_83000_3098000# diff_2851000_4962000# diff_3012000_4154000# GND efet w=130000 l=9000
+ ad=0 pd=0 as=-9.79967e+08 ps=630000 
M2774 diff_3062000_4310000# diff_530000_4372000# diff_83000_3098000# GND efet w=129000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M2775 diff_3227000_4780000# diff_3056000_4962000# diff_83000_3098000# GND efet w=66000 l=9000
+ ad=1.70603e+09 pd=1.214e+06 as=0 ps=0 
M2776 diff_3227000_4780000# diff_2135000_4721000# diff_83000_3098000# GND efet w=80000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2777 diff_3033000_4154000# diff_791000_4022000# diff_3012000_4154000# GND efet w=131000 l=9000
+ ad=-2.00097e+09 pd=442000 as=0 ps=0 
M2778 diff_1253000_4407000# diff_3116000_4962000# diff_83000_3098000# GND efet w=67500 l=8500
+ ad=1.753e+09 pd=366000 as=0 ps=0 
M2779 diff_1253000_4407000# diff_1253000_4407000# diff_95000_5192000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2780 diff_83000_3098000# diff_2998000_4962000# diff_3184000_4336000# GND efet w=130000 l=8000
+ ad=0 pd=0 as=-5.27967e+08 ps=784000 
M2781 diff_3184000_4336000# diff_3028000_4947000# diff_83000_3098000# GND efet w=176500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2782 diff_3227000_4780000# diff_1001000_4394000# diff_3184000_4336000# GND efet w=152500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2783 diff_3359000_4501000# diff_3204000_4962000# diff_83000_3098000# GND efet w=82000 l=9000
+ ad=2.11065e+08 pd=1.792e+06 as=0 ps=0 
M2784 diff_83000_3098000# diff_3301000_4962000# diff_3359000_4501000# GND efet w=65000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2785 diff_3430000_4645000# diff_3421000_4638000# diff_3359000_4501000# GND efet w=145500 l=8500
+ ad=1.385e+09 pd=310000 as=0 ps=0 
M2786 diff_83000_3098000# diff_3330000_4962000# diff_3430000_4645000# GND efet w=147500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2787 diff_95000_5192000# diff_3359000_4501000# diff_3359000_4501000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2788 diff_3272000_4383000# diff_3086000_4962000# diff_3227000_4780000# GND efet w=149000 l=8000
+ ad=1.567e+09 pd=330000 as=0 ps=0 
M2789 diff_83000_3098000# diff_791000_4022000# diff_3272000_4383000# GND efet w=155000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2790 diff_3488000_4662000# diff_3488000_4662000# diff_95000_5192000# GND efet w=12000 l=36000
+ ad=1.491e+09 pd=364000 as=0 ps=0 
M2791 diff_3539000_4683000# diff_3389000_4962000# diff_3488000_4662000# GND efet w=87000 l=8000
+ ad=8.7e+08 pd=194000 as=0 ps=0 
M2792 diff_83000_3098000# diff_1001000_4394000# diff_3539000_4683000# GND efet w=87000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2793 diff_3700000_4748000# diff_2570000_3912000# diff_83000_3098000# GND efet w=42000 l=8000
+ ad=-1.86697e+09 pd=482000 as=0 ps=0 
M2794 diff_83000_3098000# diff_3565000_4962000# diff_3700000_4748000# GND efet w=42000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2795 diff_3754000_4644000# diff_3595000_4962000# diff_83000_3098000# GND efet w=85000 l=9000
+ ad=-1.86397e+09 pd=434000 as=0 ps=0 
M2796 diff_2799000_4040000# diff_2799000_4040000# diff_95000_5192000# GND efet w=12000 l=35000
+ ad=-1.23597e+09 pd=518000 as=0 ps=0 
M2797 diff_2799000_4040000# diff_2664000_4962000# diff_2853000_4056000# GND efet w=86000 l=9000
+ ad=0 pd=0 as=7.74e+08 ps=190000 
M2798 diff_2853000_4056000# diff_519000_3032000# diff_83000_3098000# GND efet w=86000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2799 diff_2799000_4040000# diff_72000_4515000# diff_2912000_3918000# GND efet w=14000 l=10000
+ ad=0 pd=0 as=5.12e+08 ps=140000 
M2800 diff_95000_5192000# diff_1001000_4394000# diff_1001000_4394000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=-9.71967e+08 ps=522000 
M2801 diff_2050000_3807000# diff_94000_3551000# diff_83000_3098000# GND efet w=64000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2802 diff_2135000_4721000# diff_2135000_4721000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2803 diff_2324000_3768000# diff_68000_5288000# diff_2340000_3697000# GND efet w=19000 l=10000
+ ad=0 pd=0 as=3.08e+08 ps=98000 
M2804 diff_2028000_3555000# diff_2028000_3555000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=1.578e+09 pd=270000 as=0 ps=0 
M2805 diff_757000_4475000# diff_757000_4475000# diff_95000_5192000# GND efet w=12000 l=14000
+ ad=1.761e+09 pd=338000 as=0 ps=0 
M2806 diff_1188000_3107000# diff_100000_3992000# diff_83000_3098000# GND efet w=66500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2807 diff_83000_3098000# diff_1251000_3051000# diff_1188000_3107000# GND efet w=79000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M2808 diff_1281000_3071000# diff_1276000_3249000# diff_83000_3098000# GND efet w=42000 l=8000
+ ad=-2.64967e+08 pd=728000 as=0 ps=0 
M2809 diff_1328000_3051000# diff_669000_2930000# diff_83000_3098000# GND efet w=245000 l=9000
+ ad=-5.43967e+08 pd=788000 as=0 ps=0 
M2810 diff_83000_3098000# diff_687000_3101000# diff_1328000_3051000# GND efet w=204500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2811 diff_1281000_3071000# diff_68000_5288000# diff_1411000_3066000# GND efet w=13000 l=11000
+ ad=0 pd=0 as=2.84e+08 ps=90000 
M2812 diff_1048000_3119000# diff_860000_2987000# diff_83000_3098000# GND efet w=113500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2813 diff_1188000_3107000# diff_1188000_3107000# diff_95000_5192000# GND efet w=14000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2814 diff_1281000_3071000# diff_1281000_3071000# diff_95000_5192000# GND efet w=14000 l=35000
+ ad=0 pd=0 as=0 ps=0 
M2815 diff_1334000_2958000# diff_1340000_3008000# diff_1328000_3051000# GND efet w=237000 l=8000
+ ad=-2.08997e+09 pd=412000 as=0 ps=0 
M2816 diff_1148000_3109000# diff_68000_5288000# diff_1000000_2990000# GND efet w=13000 l=11000
+ ad=2.33e+08 pd=78000 as=0 ps=0 
M2817 diff_1048000_3119000# diff_1048000_3119000# diff_95000_5192000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M2818 diff_1251000_3051000# diff_68000_5288000# diff_1000000_2990000# GND efet w=12000 l=10000
+ ad=2.34e+08 pd=82000 as=0 ps=0 
M2819 diff_1482000_3103000# diff_72000_4515000# diff_1465000_3204000# GND efet w=13000 l=11000
+ ad=5.46e+08 pd=152000 as=0 ps=0 
M2820 diff_1340000_3008000# diff_1411000_3066000# diff_83000_3098000# GND efet w=118500 l=8500
+ ad=-5.80967e+08 pd=656000 as=0 ps=0 
M2821 diff_83000_3098000# diff_197000_5470000# diff_1340000_3008000# GND efet w=121500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2822 diff_1459000_2943000# diff_1482000_3103000# diff_83000_3098000# GND efet w=56000 l=8000
+ ad=-1.90297e+09 pd=474000 as=0 ps=0 
M2823 diff_132000_2382000# diff_123000_2595000# diff_95000_5192000# GND efet w=860000 l=9000
+ ad=2.26163e+06 pd=4.268e+06 as=0 ps=0 
M2824 diff_83000_3098000# diff_553000_1211000# diff_123000_2595000# GND efet w=413500 l=8500
+ ad=0 pd=0 as=-9.37902e+08 ps=1.372e+06 
M2825 diff_95000_5192000# diff_123000_2595000# diff_132000_2382000# GND efet w=342000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2826 diff_95000_5192000# diff_123000_2595000# diff_132000_2382000# GND efet w=238500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M2827 diff_83000_3098000# diff_123000_2374000# diff_123000_2595000# GND efet w=269000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2828 diff_83000_3098000# diff_123000_2374000# diff_123000_2595000# GND efet w=181000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2829 diff_553000_1211000# diff_91000_5337000# diff_83000_3098000# GND efet w=304500 l=8500
+ ad=-7.18365e+07 pd=2.282e+06 as=0 ps=0 
M2830 diff_95000_5192000# diff_123000_2595000# diff_132000_2382000# GND efet w=238500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2831 diff_123000_2595000# diff_123000_2595000# diff_95000_5192000# GND efet w=41000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2832 diff_132000_2382000# diff_123000_2374000# diff_83000_3098000# GND efet w=879000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2833 diff_83000_3098000# diff_123000_2374000# diff_132000_2382000# GND efet w=240000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2834 diff_95000_5192000# diff_123000_2374000# diff_123000_2374000# GND efet w=35000 l=8000
+ ad=0 pd=0 as=1.96607e+09 ps=1.272e+06 
M2835 diff_719000_2538000# diff_680000_1019000# diff_582000_2472000# GND efet w=34000 l=11000
+ ad=-2.69673e+07 pd=920000 as=5.79e+08 ps=108000 
M2836 diff_83000_3098000# diff_582000_2472000# diff_123000_2374000# GND efet w=412500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2837 diff_83000_3098000# diff_91000_5337000# diff_553000_1211000# GND efet w=295000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2838 diff_553000_1211000# diff_91000_5337000# diff_83000_3098000# GND efet w=295000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2839 diff_95000_5192000# diff_938000_2548000# diff_553000_1211000# GND efet w=34000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2840 diff_938000_2548000# diff_938000_2548000# diff_95000_5192000# GND efet w=26000 l=7000
+ ad=-1.23697e+09 pd=568000 as=0 ps=0 
M2841 diff_83000_3098000# diff_91000_5337000# diff_938000_2548000# GND efet w=260500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2842 diff_95000_5192000# diff_938000_2548000# diff_553000_1211000# GND efet w=138000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2843 diff_95000_5192000# diff_938000_2548000# diff_553000_1211000# GND efet w=301000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2844 diff_1334000_2958000# diff_1334000_2958000# diff_95000_5192000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M2845 diff_83000_3098000# diff_1405000_2969000# diff_1340000_3008000# GND efet w=128500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M2846 diff_1659000_2818000# diff_2028000_3555000# diff_83000_3098000# GND efet w=99500 l=7500
+ ad=3.50327e+07 pd=834000 as=0 ps=0 
M2847 diff_1556000_2817000# diff_1556000_2817000# diff_95000_5192000# GND efet w=13000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M2848 diff_83000_3098000# diff_2073000_3806000# diff_757000_4475000# GND efet w=100000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2849 diff_83000_3098000# diff_2129000_4009000# diff_2028000_3555000# GND efet w=63000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M2850 diff_2182000_3681000# diff_686000_4521000# diff_83000_3098000# GND efet w=132000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2851 diff_83000_3098000# diff_1674000_4606000# diff_2182000_3681000# GND efet w=132500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M2852 diff_83000_3098000# diff_1979000_4962000# diff_2174000_3677000# GND efet w=42000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2853 diff_1001000_4394000# diff_2340000_3697000# diff_83000_3098000# GND efet w=278500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M2854 diff_95000_5192000# diff_2050000_3807000# diff_2050000_3807000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M2855 diff_2509000_3809000# diff_2577000_4949000# diff_2559000_3889000# GND efet w=149500 l=8500
+ ad=-2.11397e+09 pd=462000 as=0 ps=0 
M2856 diff_2559000_3889000# diff_784000_3633000# diff_83000_3098000# GND efet w=146000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M2857 diff_2697000_3827000# diff_519000_3032000# diff_2509000_3809000# GND efet w=130500 l=9500
+ ad=1.095e+09 pd=278000 as=0 ps=0 
M2858 diff_83000_3098000# diff_2606000_4947000# diff_2697000_3827000# GND efet w=129500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2859 diff_95000_5192000# diff_2509000_3809000# diff_2509000_3809000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M2860 diff_2270000_3390000# diff_743000_2974000# diff_83000_3098000# GND efet w=65000 l=7000
+ ad=-6.50967e+08 pd=590000 as=0 ps=0 
M2861 diff_906000_3226000# diff_94000_3551000# diff_83000_3098000# GND efet w=125500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2862 diff_83000_3098000# diff_2868000_3892000# diff_906000_3226000# GND efet w=132000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2863 diff_83000_3098000# diff_2912000_3918000# diff_2904000_3862000# GND efet w=80000 l=8000
+ ad=0 pd=0 as=1.497e+09 ps=324000 
M2864 diff_2909000_3804000# diff_2904000_3862000# diff_83000_3098000# GND efet w=66000 l=9000
+ ad=-1.56197e+09 pd=624000 as=0 ps=0 
M2865 diff_83000_3098000# diff_2965000_3936000# diff_2909000_3804000# GND efet w=63000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2866 diff_2965000_3936000# diff_72000_4515000# diff_3009000_3950000# GND efet w=13000 l=12000
+ ad=2.38e+08 pd=82000 as=7.81e+08 ps=188000 
M2867 diff_95000_5192000# diff_3033000_4154000# diff_3033000_4154000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2868 diff_2821000_3543000# diff_72000_4515000# diff_2938000_3467000# GND efet w=20000 l=11000
+ ad=2.106e+09 pd=502000 as=2.124e+09 ps=498000 
M2869 diff_3009000_3950000# diff_3009000_3950000# diff_95000_5192000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M2870 diff_83000_3098000# diff_3024000_3904000# diff_3009000_3950000# GND efet w=42000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2871 diff_83000_3098000# diff_2882000_3711000# diff_2909000_3804000# GND efet w=70500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M2872 diff_83000_3098000# diff_2270000_3390000# diff_2219000_3479000# GND efet w=175000 l=8000
+ ad=0 pd=0 as=2.103e+09 ps=484000 
M2873 diff_1716000_2866000# diff_65000_4220000# diff_83000_3098000# GND efet w=81000 l=9000
+ ad=-1.96297e+09 pd=464000 as=0 ps=0 
M2874 diff_2219000_3479000# diff_65000_4220000# diff_1733000_2883000# GND efet w=143500 l=8500
+ ad=0 pd=0 as=-1.44297e+09 ps=594000 
M2875 diff_1659000_2818000# diff_1659000_2818000# diff_95000_5192000# GND efet w=12000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M2876 diff_83000_3098000# diff_65000_4220000# diff_1502000_2925000# GND efet w=125500 l=7500
+ ad=0 pd=0 as=-1.69346e+07 ps=1.49e+06 
M2877 diff_1502000_2925000# diff_597000_3013000# diff_83000_3098000# GND efet w=110500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2878 diff_83000_3098000# diff_1604000_3123000# diff_1502000_2925000# GND efet w=104000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2879 diff_1028000_3008000# diff_72000_4515000# diff_955000_2507000# GND efet w=28000 l=11000
+ ad=0 pd=0 as=9.44e+08 ps=204000 
M2880 diff_1048000_3119000# diff_72000_4515000# diff_1157000_2480000# GND efet w=27000 l=11000
+ ad=0 pd=0 as=1.092e+09 ps=222000 
M2881 diff_83000_3098000# diff_955000_2507000# diff_877000_1128000# GND efet w=343500 l=8500
+ ad=0 pd=0 as=8.64065e+08 ps=1.288e+06 
M2882 diff_95000_5192000# diff_877000_1128000# diff_877000_1128000# GND efet w=24000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2883 diff_901000_991000# diff_901000_991000# diff_95000_5192000# GND efet w=24000 l=8000
+ ad=9.86065e+08 pd=1.34e+06 as=0 ps=0 
M2884 diff_83000_3098000# diff_72000_4515000# diff_877000_1128000# GND efet w=334500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M2885 diff_83000_3098000# diff_123000_2374000# diff_132000_2382000# GND efet w=305500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2886 diff_901000_991000# diff_72000_4515000# diff_83000_3098000# GND efet w=292000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2887 diff_123000_2374000# diff_553000_1211000# diff_83000_3098000# GND efet w=414500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2888 diff_83000_3098000# diff_1157000_2480000# diff_901000_991000# GND efet w=338500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M2889 diff_1259000_2792000# diff_68000_5288000# diff_1259000_2736000# GND efet w=13000 l=11000
+ ad=-1.09497e+09 pd=616000 as=8.87e+08 ps=172000 
M2890 diff_1459000_2943000# diff_1459000_2943000# diff_95000_5192000# GND efet w=13000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M2891 diff_1340000_3008000# diff_1340000_3008000# diff_95000_5192000# GND efet w=14000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M2892 diff_83000_3098000# diff_967000_2989000# diff_1502000_2925000# GND efet w=118000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2893 diff_1502000_2925000# diff_860000_2987000# diff_83000_3098000# GND efet w=123500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2894 diff_83000_3098000# diff_1586000_2912000# diff_1502000_2925000# GND efet w=124000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2895 diff_1502000_2925000# diff_1502000_2925000# diff_95000_5192000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M2896 diff_1459000_2943000# diff_68000_5288000# diff_1405000_2969000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=5.82e+08 ps=130000 
M2897 diff_1000000_2990000# diff_68000_5288000# diff_1586000_2912000# GND efet w=14000 l=11000
+ ad=0 pd=0 as=4.69e+08 ps=134000 
M2898 diff_83000_3098000# diff_94000_3551000# diff_2270000_3390000# GND efet w=61000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2899 diff_1817000_2934000# diff_94000_3551000# diff_83000_3098000# GND efet w=64500 l=8500
+ ad=1.385e+09 pd=308000 as=0 ps=0 
M2900 diff_1817000_2934000# diff_1817000_2934000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2901 diff_95000_5192000# diff_1716000_2866000# diff_1716000_2866000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2902 diff_95000_5192000# diff_1733000_2883000# diff_1733000_2883000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2903 diff_2270000_3390000# diff_2270000_3390000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2904 diff_2904000_3862000# diff_2904000_3862000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2905 diff_3005000_3816000# diff_68000_5288000# diff_3024000_3904000# GND efet w=11000 l=11000
+ ad=1.142e+09 pd=250000 as=3.34e+08 ps=128000 
M2906 diff_906000_3226000# diff_906000_3226000# diff_906000_3226000# GND efet w=1000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M2907 diff_2909000_3804000# diff_68000_5288000# diff_2868000_3892000# GND efet w=13000 l=10000
+ ad=0 pd=0 as=6.45e+08 ps=176000 
M2908 diff_95000_5192000# diff_906000_3226000# diff_906000_3226000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M2909 diff_2909000_3804000# diff_2909000_3804000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2910 diff_83000_3098000# diff_3032000_3774000# diff_3005000_3816000# GND efet w=43000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2911 diff_3005000_3816000# diff_3005000_3816000# diff_95000_5192000# GND efet w=13000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M2912 diff_519000_3032000# diff_72000_4515000# diff_2660000_3493000# GND efet w=14000 l=13000
+ ad=0 pd=0 as=1.988e+09 ps=452000 
M2913 diff_2772000_3402000# diff_72000_4515000# diff_3032000_3774000# GND efet w=12000 l=12000
+ ad=-1.98997e+09 pd=534000 as=4.6e+08 ps=136000 
M2914 diff_83000_3098000# diff_2566000_3500000# diff_1604000_3123000# GND efet w=183000 l=8000
+ ad=0 pd=0 as=-1.20097e+09 ps=610000 
M2915 diff_83000_3098000# diff_2598000_3304000# diff_530000_4372000# GND efet w=291000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2916 diff_65000_4220000# diff_72000_4515000# diff_2882000_3711000# GND efet w=14000 l=10000
+ ad=0 pd=0 as=8.52e+08 ps=238000 
M2917 diff_530000_4372000# diff_530000_4372000# diff_95000_5192000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2918 diff_2651000_3482000# diff_2642000_3475000# diff_83000_3098000# GND efet w=134500 l=8500
+ ad=1.284e+09 pd=288000 as=0 ps=0 
M2919 diff_2633000_3304000# diff_2660000_3493000# diff_2651000_3482000# GND efet w=134000 l=8000
+ ad=-7.84967e+08 pd=662000 as=0 ps=0 
M2920 diff_83000_3098000# diff_94000_3551000# diff_2660000_3493000# GND efet w=65000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M2921 diff_3227000_4780000# diff_3227000_4780000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2922 diff_3048000_3539000# diff_68000_5288000# diff_2878000_4622000# GND efet w=13000 l=11000
+ ad=4.5e+08 pd=134000 as=0 ps=0 
M2923 diff_83000_3098000# diff_1840000_3083000# diff_1826000_2942000# GND efet w=184500 l=7500
+ ad=0 pd=0 as=2.08033e+08 ps=878000 
M2924 diff_1751000_2974000# diff_1751000_2974000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=-1.58597e+09 pd=568000 as=0 ps=0 
M2925 diff_1808000_2942000# diff_65000_4220000# diff_1751000_2974000# GND efet w=175000 l=9000
+ ad=1.575e+09 pd=368000 as=0 ps=0 
M2926 diff_1826000_2942000# diff_1817000_2934000# diff_1808000_2942000# GND efet w=175000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2927 diff_83000_3098000# diff_743000_2974000# diff_1826000_2942000# GND efet w=25000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2928 diff_83000_3098000# diff_74000_3122000# diff_1840000_3083000# GND efet w=78500 l=8500
+ ad=0 pd=0 as=1.794e+09 ps=386000 
M2929 diff_1935000_3038000# diff_817000_909000# diff_83000_3098000# GND efet w=115500 l=8500
+ ad=-8.61967e+08 pd=626000 as=0 ps=0 
M2930 diff_1962000_3117000# diff_68000_5288000# diff_2004000_3055000# GND efet w=12000 l=12000
+ ad=2.7e+08 pd=76000 as=-1.35897e+09 ps=568000 
M2931 diff_1998000_3198000# diff_72000_4515000# diff_1698000_2848000# GND efet w=13000 l=12000
+ ad=3.93e+08 pd=108000 as=-5.92967e+08 ps=812000 
M2932 diff_83000_3098000# diff_743000_2974000# diff_1826000_2942000# GND efet w=155500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2933 diff_1840000_3083000# diff_1840000_3083000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2934 diff_1556000_2817000# diff_72000_4515000# diff_1554000_2586000# GND efet w=20000 l=12000
+ ad=0 pd=0 as=8.81e+08 ps=156000 
M2935 diff_1188000_3107000# diff_72000_4515000# diff_1610000_2779000# GND efet w=21000 l=13000
+ ad=0 pd=0 as=8.58e+08 ps=152000 
M2936 diff_1659000_2818000# diff_72000_4515000# diff_1659000_2777000# GND efet w=21000 l=13000
+ ad=0 pd=0 as=9.44e+08 ps=154000 
M2937 diff_83000_3098000# diff_1962000_3117000# diff_1963000_2987000# GND efet w=69000 l=8000
+ ad=0 pd=0 as=2.011e+09 ps=422000 
M2938 diff_2004000_3055000# diff_1998000_3198000# diff_83000_3098000# GND efet w=63000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2939 diff_2110000_2945000# diff_72000_4515000# diff_2082000_3201000# GND efet w=13000 l=11000
+ ad=-1.16497e+09 pd=576000 as=5.9e+08 ps=142000 
M2940 diff_95000_5192000# diff_1604000_3123000# diff_1604000_3123000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2941 diff_2633000_3304000# diff_2633000_3304000# diff_95000_5192000# GND efet w=13000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M2942 diff_2633000_3304000# diff_68000_5288000# diff_2598000_3304000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=4.75e+08 ps=98000 
M2943 diff_2066000_3013000# diff_2004000_3055000# diff_83000_3098000# GND efet w=115000 l=9000
+ ad=-1.97097e+09 pd=502000 as=0 ps=0 
M2944 diff_83000_3098000# diff_2082000_3201000# diff_2066000_3013000# GND efet w=115500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M2945 diff_2134000_3060000# diff_1097000_3119000# diff_83000_3098000# GND efet w=65000 l=8000
+ ad=-1.38997e+09 pd=554000 as=0 ps=0 
M2946 diff_2004000_3055000# diff_2004000_3055000# diff_95000_5192000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M2947 diff_95000_5192000# diff_1963000_2987000# diff_1963000_2987000# GND efet w=11000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M2948 diff_95000_5192000# diff_1935000_3038000# diff_1935000_3038000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M2949 diff_2066000_3013000# diff_2066000_3013000# diff_95000_5192000# GND efet w=13000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M2950 diff_2134000_3060000# diff_2134000_3060000# diff_95000_5192000# GND efet w=11000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M2951 diff_83000_3098000# diff_2198000_3000000# diff_2293000_3174000# GND efet w=152500 l=7500
+ ad=0 pd=0 as=-6.13967e+08 ps=744000 
M2952 diff_83000_3098000# diff_2198000_3000000# diff_2182000_3046000# GND efet w=40000 l=9000
+ ad=0 pd=0 as=1.14033e+08 ps=874000 
M2953 diff_2182000_3046000# diff_2134000_3060000# diff_83000_3098000# GND efet w=130000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2954 diff_83000_3098000# diff_2248000_3126000# diff_2182000_3046000# GND efet w=146000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2955 diff_2182000_3046000# diff_2173000_3038000# diff_2110000_2945000# GND efet w=153000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2956 diff_83000_3098000# diff_2198000_3000000# diff_2182000_3046000# GND efet w=103000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2957 diff_2293000_3174000# diff_2248000_3126000# diff_83000_3098000# GND efet w=143000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2958 diff_2356000_3007000# diff_2351000_3074000# diff_2293000_3174000# GND efet w=133000 l=8000
+ ad=-1.50997e+09 pd=428000 as=0 ps=0 
M2959 diff_2390000_3201000# diff_72000_4515000# diff_2356000_3007000# GND efet w=13000 l=12000
+ ad=2.69e+08 pd=96000 as=0 ps=0 
M2960 diff_2134000_3060000# diff_72000_4515000# diff_2420000_3102000# GND efet w=13000 l=11000
+ ad=0 pd=0 as=2.27e+08 ps=72000 
M2961 diff_2400000_2876000# diff_2390000_3201000# diff_83000_3098000# GND efet w=78000 l=9000
+ ad=1.513e+09 pd=316000 as=0 ps=0 
M2962 diff_83000_3098000# diff_2420000_3102000# diff_2400000_2876000# GND efet w=83000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2963 diff_83000_3098000# diff_2464000_2895000# diff_1259000_2792000# GND efet w=120000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2964 diff_1935000_3038000# diff_68000_5288000# diff_2248000_3126000# GND efet w=13000 l=11000
+ ad=0 pd=0 as=1.82e+08 ps=54000 
M2965 diff_2110000_2945000# diff_2110000_2945000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M2966 diff_1698000_2848000# diff_72000_4515000# diff_1712000_2778000# GND efet w=20000 l=13000
+ ad=0 pd=0 as=9.56e+08 ps=154000 
M2967 diff_1716000_2866000# diff_72000_4515000# diff_1776000_2770000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=1.05e+09 ps=160000 
M2968 diff_1733000_2883000# diff_72000_4515000# diff_1816000_2509000# GND efet w=14000 l=11000
+ ad=0 pd=0 as=1.141e+09 ps=164000 
M2969 diff_1751000_2974000# diff_72000_4515000# diff_1874000_2769000# GND efet w=14000 l=11000
+ ad=0 pd=0 as=1.037e+09 ps=160000 
M2970 diff_95000_5192000# diff_1276000_2574000# diff_1276000_2574000# GND efet w=13000 l=9000
+ ad=0 pd=0 as=1.63033e+08 ps=552000 
M2971 diff_95000_5192000# diff_1318000_2487000# diff_1318000_2487000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=1.327e+09 ps=326000 
M2972 diff_1276000_2574000# diff_1259000_2736000# diff_83000_3098000# GND efet w=116000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2973 diff_1281000_2492000# diff_1150000_1007000# diff_1276000_2574000# GND efet w=203500 l=8500
+ ad=-1.80497e+09 pd=470000 as=0 ps=0 
M2974 diff_132000_2005000# diff_123000_2207000# diff_83000_3098000# GND efet w=880500 l=8500
+ ad=-1.36738e+08 pd=4.268e+06 as=0 ps=0 
M2975 diff_83000_3098000# diff_123000_2207000# diff_132000_2005000# GND efet w=305000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2976 diff_83000_3098000# diff_553000_1211000# diff_123000_2207000# GND efet w=414500 l=8500
+ ad=0 pd=0 as=-2.0919e+09 ps=1.276e+06 
M2977 diff_83000_3098000# diff_1318000_2487000# diff_1281000_2492000# GND efet w=198000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2978 diff_1393000_2558000# diff_1393000_2558000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=-1.16097e+09 pd=580000 as=0 ps=0 
M2979 diff_95000_5192000# diff_1176000_1643000# diff_1176000_1643000# GND efet w=13000 l=9000
+ ad=0 pd=0 as=1.7061e+09 ps=2.726e+06 
M2980 diff_83000_3098000# diff_1334000_2958000# diff_1318000_2487000# GND efet w=77500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M2981 diff_1393000_2558000# diff_1334000_2958000# diff_83000_3098000# GND efet w=72500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2982 diff_83000_3098000# diff_1237000_1921000# diff_1393000_2558000# GND efet w=81000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2983 diff_83000_3098000# diff_1393000_2558000# diff_1252000_2261000# GND efet w=148500 l=9500
+ ad=0 pd=0 as=-2.10393e+09 ps=1.024e+06 
M2984 diff_1176000_1643000# diff_1334000_2958000# diff_83000_3098000# GND efet w=160000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2985 diff_95000_5192000# diff_1487000_841000# diff_1487000_841000# GND efet w=21000 l=7000
+ ad=0 pd=0 as=-2.14935e+08 ps=1.268e+06 
M2986 diff_1547000_932000# diff_1547000_932000# diff_95000_5192000# GND efet w=15000 l=8000
+ ad=1.41203e+09 pd=1.102e+06 as=0 ps=0 
M2987 diff_83000_3098000# diff_1237000_1921000# diff_1176000_1643000# GND efet w=188000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2988 diff_83000_3098000# diff_582000_2217000# diff_123000_2207000# GND efet w=413500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2989 diff_83000_3098000# diff_123000_2207000# diff_132000_2005000# GND efet w=240000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2990 diff_856000_2349000# diff_848000_2342000# diff_83000_3098000# GND efet w=132000 l=8000
+ ad=1.733e+09 pd=330000 as=0 ps=0 
M2991 diff_95000_5192000# diff_856000_2349000# diff_856000_2349000# GND efet w=12000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2992 diff_817000_2342000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=103000
+ ad=-1.63784e+09 pd=3.958e+06 as=0 ps=0 
M2993 diff_95000_5192000# diff_914000_2210000# diff_914000_2210000# GND efet w=13000 l=7000
+ ad=0 pd=0 as=2.018e+09 ps=432000 
M2994 diff_719000_2538000# diff_889000_2284000# diff_83000_3098000# GND efet w=104500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M2995 diff_83000_3098000# diff_817000_2342000# diff_914000_2210000# GND efet w=143000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2996 diff_95000_5192000# diff_719000_2538000# diff_719000_2538000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M2997 diff_1064000_2211000# diff_1064000_2211000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=-1.72397e+09 pd=452000 as=0 ps=0 
M2998 diff_889000_2284000# diff_877000_1128000# diff_856000_2349000# GND efet w=19000 l=11000
+ ad=4.18e+08 pd=82000 as=0 ps=0 
M2999 diff_914000_2210000# diff_901000_991000# diff_889000_2284000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3000 diff_95000_5192000# diff_123000_1997000# diff_132000_2005000# GND efet w=238500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3001 diff_123000_2207000# diff_123000_2207000# diff_95000_5192000# GND efet w=35000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3002 diff_582000_2217000# diff_680000_1019000# diff_719000_2180000# GND efet w=34000 l=11000
+ ad=5.18e+08 pd=102000 as=-8.69967e+08 ps=714000 
M3003 diff_95000_5192000# diff_123000_1997000# diff_123000_1997000# GND efet w=41000 l=9000
+ ad=0 pd=0 as=-1.2499e+09 ps=1.366e+06 
M3004 diff_132000_2005000# diff_123000_1997000# diff_95000_5192000# GND efet w=855000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3005 diff_95000_5192000# diff_123000_1997000# diff_132000_2005000# GND efet w=238500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3006 diff_83000_3098000# diff_123000_2207000# diff_123000_1997000# GND efet w=179000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3007 diff_95000_5192000# diff_123000_1997000# diff_132000_2005000# GND efet w=342500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3008 diff_83000_3098000# diff_123000_2207000# diff_123000_1997000# GND efet w=269000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3009 diff_123000_1997000# diff_553000_1211000# diff_83000_3098000# GND efet w=413000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3010 diff_132000_1628000# diff_123000_1841000# diff_95000_5192000# GND efet w=859000 l=9000
+ ad=-5.27738e+08 pd=4.268e+06 as=0 ps=0 
M3011 diff_83000_3098000# diff_553000_1211000# diff_123000_1841000# GND efet w=413500 l=8500
+ ad=0 pd=0 as=-1.0199e+09 ps=1.376e+06 
M3012 diff_95000_5192000# diff_123000_1841000# diff_132000_1628000# GND efet w=342500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3013 diff_83000_3098000# diff_123000_1620000# diff_123000_1841000# GND efet w=270000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3014 diff_95000_5192000# diff_123000_1841000# diff_132000_1628000# GND efet w=238500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3015 diff_83000_3098000# diff_123000_1620000# diff_123000_1841000# GND efet w=181000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3016 diff_95000_5192000# diff_123000_1841000# diff_132000_1628000# GND efet w=238500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3017 diff_123000_1841000# diff_123000_1841000# diff_95000_5192000# GND efet w=42000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3018 diff_95000_5192000# diff_95000_5192000# diff_817000_2040000# GND efet w=12000 l=103000
+ ad=0 pd=0 as=-2.89836e+08 ps=4.278e+06 
M3019 diff_856000_2022000# diff_848000_2016000# diff_83000_3098000# GND efet w=130000 l=8000
+ ad=1.722e+09 pd=332000 as=0 ps=0 
M3020 diff_1010000_2204000# diff_889000_2284000# diff_83000_3098000# GND efet w=36000 l=8000
+ ad=1.607e+09 pd=358000 as=0 ps=0 
M3021 diff_719000_2538000# diff_889000_2284000# diff_83000_3098000# GND efet w=47000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3022 diff_1010000_2204000# diff_889000_2284000# diff_83000_3098000# GND efet w=77500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3023 diff_1064000_2211000# diff_1037000_877000# diff_1010000_2204000# GND efet w=121000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3024 diff_1085000_2211000# diff_719000_2538000# diff_1064000_2211000# GND efet w=73500 l=8500
+ ad=1.506e+09 pd=340000 as=0 ps=0 
M3025 diff_83000_3098000# diff_1094000_1020000# diff_1085000_2211000# GND efet w=139000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3026 diff_1085000_2211000# diff_719000_2538000# diff_1064000_2211000# GND efet w=45000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3027 diff_1150000_1007000# diff_1064000_2211000# diff_83000_3098000# GND efet w=84000 l=8000
+ ad=-2.20836e+08 pd=3.454e+06 as=0 ps=0 
M3028 diff_1150000_1007000# diff_1064000_2211000# diff_83000_3098000# GND efet w=43000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M3029 diff_83000_3098000# diff_817000_2040000# diff_914000_2134000# GND efet w=141000 l=8000
+ ad=0 pd=0 as=2.019e+09 ps=430000 
M3030 diff_889000_2094000# diff_877000_1128000# diff_856000_2022000# GND efet w=19000 l=11000
+ ad=4.18e+08 pd=82000 as=0 ps=0 
M3031 diff_914000_2134000# diff_901000_991000# diff_889000_2094000# GND efet w=19000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M3032 diff_719000_2180000# diff_889000_2094000# diff_83000_3098000# GND efet w=47000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3033 diff_1010000_2185000# diff_889000_2094000# diff_83000_3098000# GND efet w=80000 l=8000
+ ad=1.537e+09 pd=360000 as=0 ps=0 
M3034 diff_719000_2180000# diff_889000_2094000# diff_83000_3098000# GND efet w=102000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3035 diff_95000_5192000# diff_856000_2022000# diff_856000_2022000# GND efet w=12000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3036 diff_856000_1972000# diff_848000_1965000# diff_83000_3098000# GND efet w=132000 l=8000
+ ad=1.782e+09 pd=330000 as=0 ps=0 
M3037 diff_95000_5192000# diff_856000_1972000# diff_856000_1972000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3038 diff_817000_1965000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=103000
+ ad=-6.19869e+08 pd=3.332e+06 as=0 ps=0 
M3039 diff_95000_5192000# diff_914000_2134000# diff_914000_2134000# GND efet w=13000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M3040 diff_1010000_2185000# diff_889000_2094000# diff_83000_3098000# GND efet w=37000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3041 diff_1064000_2064000# diff_1037000_877000# diff_1010000_2185000# GND efet w=121000 l=9000
+ ad=-1.67197e+09 pd=460000 as=0 ps=0 
M3042 diff_1085000_2099000# diff_719000_2180000# diff_1064000_2064000# GND efet w=44000 l=9000
+ ad=1.54e+09 pd=334000 as=0 ps=0 
M3043 diff_83000_3098000# diff_1094000_1020000# diff_1085000_2099000# GND efet w=137000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3044 diff_1085000_2099000# diff_719000_2180000# diff_1064000_2064000# GND efet w=72000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3045 diff_1150000_1007000# diff_1064000_2064000# diff_83000_3098000# GND efet w=43000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M3046 diff_95000_5192000# diff_719000_2180000# diff_719000_2180000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3047 diff_95000_5192000# diff_914000_1833000# diff_914000_1833000# GND efet w=13000 l=7000
+ ad=0 pd=0 as=2.042e+09 ps=430000 
M3048 diff_719000_1784000# diff_889000_1907000# diff_83000_3098000# GND efet w=104500 l=8500
+ ad=-9.30967e+08 pd=704000 as=0 ps=0 
M3049 diff_83000_3098000# diff_817000_1965000# diff_914000_1833000# GND efet w=142000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3050 diff_95000_5192000# diff_719000_1784000# diff_719000_1784000# GND efet w=12000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3051 diff_1064000_2064000# diff_1064000_2064000# diff_95000_5192000# GND efet w=14000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3052 diff_1064000_1834000# diff_1064000_1834000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=-1.71897e+09 pd=454000 as=0 ps=0 
M3053 diff_1150000_1007000# diff_1064000_2064000# diff_83000_3098000# GND efet w=84000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3054 diff_889000_1907000# diff_877000_1128000# diff_856000_1972000# GND efet w=19000 l=10000
+ ad=4.18e+08 pd=82000 as=0 ps=0 
M3055 diff_914000_1833000# diff_901000_991000# diff_889000_1907000# GND efet w=19000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M3056 diff_132000_1628000# diff_123000_1620000# diff_83000_3098000# GND efet w=877000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3057 diff_83000_3098000# diff_123000_1620000# diff_132000_1628000# GND efet w=240000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3058 diff_95000_5192000# diff_123000_1620000# diff_123000_1620000# GND efet w=35000 l=8000
+ ad=0 pd=0 as=2.02807e+09 ps=1.272e+06 
M3059 diff_719000_1784000# diff_680000_1019000# diff_582000_1718000# GND efet w=34000 l=11000
+ ad=0 pd=0 as=5.9e+08 ps=108000 
M3060 diff_83000_3098000# diff_582000_1718000# diff_123000_1620000# GND efet w=412500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3061 diff_83000_3098000# diff_123000_1620000# diff_132000_1628000# GND efet w=305000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3062 diff_123000_1620000# diff_553000_1211000# diff_83000_3098000# GND efet w=415500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3063 diff_95000_5192000# diff_95000_5192000# diff_817000_1663000# GND efet w=12000 l=104000
+ ad=0 pd=0 as=1.51113e+09 ps=3.796e+06 
M3064 diff_856000_1645000# diff_848000_1639000# diff_83000_3098000# GND efet w=130000 l=8000
+ ad=1.713e+09 pd=330000 as=0 ps=0 
M3065 diff_1010000_1827000# diff_889000_1907000# diff_83000_3098000# GND efet w=37000 l=8000
+ ad=1.648e+09 pd=360000 as=0 ps=0 
M3066 diff_719000_1784000# diff_889000_1907000# diff_83000_3098000# GND efet w=48000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3067 diff_1010000_1827000# diff_889000_1907000# diff_83000_3098000# GND efet w=77000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3068 diff_1064000_1834000# diff_1037000_877000# diff_1010000_1827000# GND efet w=122000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3069 diff_1085000_1834000# diff_719000_1784000# diff_1064000_1834000# GND efet w=74500 l=8500
+ ad=1.497e+09 pd=340000 as=0 ps=0 
M3070 diff_83000_3098000# diff_1094000_1020000# diff_1085000_1834000# GND efet w=140500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3071 diff_1085000_1834000# diff_719000_1784000# diff_1064000_1834000# GND efet w=45000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3072 diff_1150000_1007000# diff_1064000_1834000# diff_83000_3098000# GND efet w=84000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3073 diff_1150000_1007000# diff_1064000_1834000# diff_83000_3098000# GND efet w=43000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M3074 diff_83000_3098000# diff_817000_1663000# diff_914000_1757000# GND efet w=141000 l=8000
+ ad=0 pd=0 as=2.019e+09 ps=430000 
M3075 diff_888000_1717000# diff_877000_1128000# diff_856000_1645000# GND efet w=19000 l=10000
+ ad=4.18e+08 pd=82000 as=0 ps=0 
M3076 diff_914000_1757000# diff_901000_991000# diff_888000_1717000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M3077 diff_719000_1426000# diff_888000_1717000# diff_83000_3098000# GND efet w=47000 l=8000
+ ad=2.24033e+08 pd=940000 as=0 ps=0 
M3078 diff_1010000_1808000# diff_888000_1717000# diff_83000_3098000# GND efet w=80000 l=8000
+ ad=1.536e+09 pd=360000 as=0 ps=0 
M3079 diff_719000_1426000# diff_888000_1717000# diff_83000_3098000# GND efet w=101500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3080 diff_132000_1251000# diff_123000_1453000# diff_83000_3098000# GND efet w=882500 l=8500
+ ad=-6.52738e+08 pd=4.276e+06 as=0 ps=0 
M3081 diff_83000_3098000# diff_123000_1453000# diff_132000_1251000# GND efet w=305000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3082 diff_83000_3098000# diff_553000_1211000# diff_123000_1453000# GND efet w=414500 l=8500
+ ad=0 pd=0 as=-2.0929e+09 ps=1.276e+06 
M3083 diff_95000_5192000# diff_856000_1645000# diff_856000_1645000# GND efet w=11000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3084 diff_83000_3098000# diff_582000_1463000# diff_123000_1453000# GND efet w=413500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3085 diff_83000_3098000# diff_123000_1453000# diff_132000_1251000# GND efet w=240500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3086 diff_856000_1595000# diff_848000_1588000# diff_83000_3098000# GND efet w=132000 l=8000
+ ad=1.763e+09 pd=328000 as=0 ps=0 
M3087 diff_95000_5192000# diff_856000_1595000# diff_856000_1595000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3088 diff_817000_1588000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=103000
+ ad=1.38213e+09 pd=3.708e+06 as=0 ps=0 
M3089 diff_95000_5192000# diff_914000_1757000# diff_914000_1757000# GND efet w=13000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M3090 diff_1010000_1808000# diff_888000_1717000# diff_83000_3098000# GND efet w=37000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3091 diff_1064000_1687000# diff_1037000_877000# diff_1010000_1808000# GND efet w=121000 l=9000
+ ad=-1.70597e+09 pd=456000 as=0 ps=0 
M3092 diff_1085000_1723000# diff_719000_1426000# diff_1064000_1687000# GND efet w=44000 l=9000
+ ad=1.525e+09 pd=336000 as=0 ps=0 
M3093 diff_83000_3098000# diff_1094000_1020000# diff_1085000_1723000# GND efet w=138000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3094 diff_1085000_1723000# diff_719000_1426000# diff_1064000_1687000# GND efet w=72000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3095 diff_1150000_1007000# diff_1064000_1687000# diff_83000_3098000# GND efet w=43000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M3096 diff_95000_5192000# diff_719000_1426000# diff_719000_1426000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3097 diff_95000_5192000# diff_914000_1456000# diff_914000_1456000# GND efet w=13000 l=7000
+ ad=0 pd=0 as=2.042e+09 ps=430000 
M3098 diff_719000_1030000# diff_889000_1530000# diff_83000_3098000# GND efet w=104500 l=8500
+ ad=3.50327e+07 pd=928000 as=0 ps=0 
M3099 diff_83000_3098000# diff_817000_1588000# diff_914000_1456000# GND efet w=142000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3100 diff_95000_5192000# diff_719000_1030000# diff_719000_1030000# GND efet w=12000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3101 diff_1064000_1687000# diff_1064000_1687000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3102 diff_1063000_1457000# diff_1063000_1457000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=-1.59697e+09 pd=456000 as=0 ps=0 
M3103 diff_1150000_1007000# diff_1064000_1687000# diff_83000_3098000# GND efet w=84000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3104 diff_95000_5192000# diff_1189000_2359000# diff_1189000_2359000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=1.401e+09 ps=284000 
M3105 diff_1487000_841000# diff_1554000_2586000# diff_83000_3098000# GND efet w=295500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3106 diff_83000_3098000# diff_72000_4515000# diff_1487000_841000# GND efet w=253000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3107 diff_1547000_932000# diff_72000_4515000# diff_83000_3098000# GND efet w=231500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3108 diff_83000_3098000# diff_1610000_2779000# diff_1547000_932000# GND efet w=255500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3109 diff_1643000_833000# diff_1659000_2777000# diff_83000_3098000# GND efet w=246000 l=9000
+ ad=2.18033e+08 pd=894000 as=0 ps=0 
M3110 diff_95000_5192000# diff_1643000_833000# diff_1643000_833000# GND efet w=17000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3111 diff_1696000_986000# diff_1696000_986000# diff_95000_5192000# GND efet w=17000 l=8000
+ ad=9.59033e+08 pd=906000 as=0 ps=0 
M3112 diff_83000_3098000# diff_72000_4515000# diff_1643000_833000# GND efet w=201000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3113 diff_1696000_986000# diff_72000_4515000# diff_83000_3098000# GND efet w=201000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3114 diff_83000_3098000# diff_1712000_2778000# diff_1696000_986000# GND efet w=246500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3115 diff_95000_5192000# diff_1728000_2245000# diff_1728000_2245000# GND efet w=13000 l=15000
+ ad=0 pd=0 as=-1.70097e+09 ps=536000 
M3116 diff_95000_5192000# diff_1931000_2739000# diff_1931000_2739000# GND efet w=12000 l=15000
+ ad=0 pd=0 as=1.371e+09 ps=274000 
M3117 diff_1728000_2245000# diff_72000_4515000# diff_83000_3098000# GND efet w=102000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3118 diff_83000_3098000# diff_1776000_2770000# diff_1728000_2245000# GND efet w=119500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3119 diff_95000_5192000# diff_68000_5288000# diff_680000_1019000# GND efet w=12000 l=10000
+ ad=0 pd=0 as=-9.62967e+08 ps=452000 
M3120 diff_95000_5192000# diff_1729000_2091000# diff_1729000_2091000# GND efet w=11000 l=14000
+ ad=0 pd=0 as=-2.13097e+09 ps=506000 
M3121 diff_1729000_1868000# diff_1729000_1868000# diff_95000_5192000# GND efet w=11000 l=14000
+ ad=-1.76897e+09 pd=484000 as=0 ps=0 
M3122 diff_1931000_2739000# diff_68000_5288000# diff_83000_3098000# GND efet w=121500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3123 diff_680000_1019000# diff_72000_4515000# diff_83000_3098000# GND efet w=164500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3124 diff_83000_3098000# diff_1931000_2739000# diff_680000_1019000# GND efet w=176500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3125 diff_1729000_2091000# diff_1816000_2509000# diff_83000_3098000# GND efet w=107500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3126 diff_83000_3098000# diff_72000_4515000# diff_1729000_2091000# GND efet w=108000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3127 diff_1729000_1868000# diff_72000_4515000# diff_83000_3098000# GND efet w=107000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3128 diff_83000_3098000# diff_1874000_2769000# diff_1729000_1868000# GND efet w=107500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3129 diff_2356000_3007000# diff_2356000_3007000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3130 diff_2400000_2876000# diff_2400000_2876000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3131 diff_1963000_2987000# diff_72000_4515000# diff_2060000_2777000# GND efet w=21000 l=13000
+ ad=0 pd=0 as=9.53e+08 ps=154000 
M3132 diff_1259000_2792000# diff_1259000_2792000# diff_95000_5192000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M3133 diff_2561000_3213000# diff_72000_4515000# diff_2521000_3105000# GND efet w=14000 l=12000
+ ad=-1.83967e+08 pd=762000 as=2.72e+08 ps=92000 
M3134 diff_2464000_2895000# diff_2521000_3105000# diff_83000_3098000# GND efet w=80000 l=8000
+ ad=1.598e+09 pd=338000 as=0 ps=0 
M3135 diff_83000_3098000# diff_2400000_2876000# diff_2464000_2895000# GND efet w=79500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3136 diff_2561000_3213000# diff_2573000_3039000# diff_83000_3098000# GND efet w=70000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3137 diff_2464000_2895000# diff_2464000_2895000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3138 diff_83000_3098000# diff_2198000_3000000# diff_2561000_3213000# GND efet w=65000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3139 diff_3017000_3539000# diff_72000_4515000# diff_3014000_3475000# GND efet w=12000 l=11000
+ ad=4e+08 pd=136000 as=-1.04797e+09 ps=692000 
M3140 diff_83000_3098000# diff_2790000_3479000# diff_2772000_3402000# GND efet w=77500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3141 diff_83000_3098000# diff_94000_3551000# diff_2821000_3543000# GND efet w=65000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3142 diff_83000_3098000# diff_2821000_3543000# diff_2810000_3352000# GND efet w=42000 l=9000
+ ad=0 pd=0 as=-1.55397e+09 ps=586000 
M3143 diff_3380000_4294000# diff_1253000_4407000# diff_3359000_4501000# GND efet w=199500 l=7500
+ ad=2.102e+09 pd=420000 as=0 ps=0 
M3144 diff_3399000_4294000# diff_3271000_4962000# diff_3380000_4294000# GND efet w=199500 l=8500
+ ad=1.863e+09 pd=420000 as=0 ps=0 
M3145 diff_83000_3098000# diff_3408000_4288000# diff_3399000_4294000# GND efet w=201500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3146 diff_3421000_4638000# diff_3408000_4288000# diff_83000_3098000# GND efet w=42000 l=9000
+ ad=1.802e+09 pd=474000 as=0 ps=0 
M3147 diff_3494000_4370000# diff_3360000_4962000# diff_83000_3098000# GND efet w=148500 l=8500
+ ad=1.792e+09 pd=318000 as=0 ps=0 
M3148 diff_3401000_3461000# diff_519000_3032000# diff_3494000_4370000# GND efet w=142000 l=8000
+ ad=-1.60597e+09 pd=598000 as=0 ps=0 
M3149 diff_3535000_4387000# diff_3389000_4962000# diff_3401000_3461000# GND efet w=148000 l=8000
+ ad=1.663e+09 pd=320000 as=0 ps=0 
M3150 diff_83000_3098000# diff_1001000_4394000# diff_3535000_4387000# GND efet w=150500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3151 diff_3421000_4638000# diff_3421000_4638000# diff_95000_5192000# GND efet w=13000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M3152 diff_3272000_3283000# diff_3360000_4962000# diff_83000_3098000# GND efet w=49500 l=7500
+ ad=8.65e+08 pd=220000 as=0 ps=0 
M3153 diff_2772000_3402000# diff_2772000_3402000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3154 diff_3272000_3283000# diff_3272000_3283000# diff_95000_5192000# GND efet w=12000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M3155 diff_530000_4372000# diff_72000_4515000# diff_3339000_4042000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.12e+08 ps=86000 
M3156 diff_3348000_3929000# diff_3339000_4042000# diff_3325000_3886000# GND efet w=144000 l=8000
+ ad=1.44e+09 pd=308000 as=-2.03697e+09 ps=472000 
M3157 diff_83000_3098000# diff_2606000_4947000# diff_3348000_3929000# GND efet w=144000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3158 diff_2790000_3479000# diff_68000_5288000# diff_2810000_3352000# GND efet w=14000 l=11000
+ ad=2.58e+08 pd=80000 as=0 ps=0 
M3159 diff_2810000_3352000# diff_2810000_3352000# diff_95000_5192000# GND efet w=13000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M3160 diff_2561000_3213000# diff_2134000_3060000# diff_83000_3098000# GND efet w=67500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3161 diff_83000_3098000# diff_2351000_3074000# diff_2561000_3213000# GND efet w=76500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3162 diff_2678000_3055000# diff_906000_3226000# diff_83000_3098000# GND efet w=72000 l=8000
+ ad=1.908e+09 pd=420000 as=0 ps=0 
M3163 diff_83000_3098000# diff_402000_4713000# diff_2678000_3055000# GND efet w=81000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3164 diff_1935000_3038000# diff_68000_5288000# diff_2573000_3039000# GND efet w=13000 l=11000
+ ad=0 pd=0 as=3.03e+08 ps=92000 
M3165 diff_2561000_3213000# diff_2561000_3213000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3166 diff_2678000_3055000# diff_2678000_3055000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3167 diff_1659000_2818000# diff_72000_4515000# diff_2113000_2778000# GND efet w=21000 l=13000
+ ad=0 pd=0 as=9.66e+08 ps=156000 
M3168 diff_2066000_3013000# diff_68000_5288000# diff_2208000_2717000# GND efet w=18000 l=12000
+ ad=0 pd=0 as=9.03e+08 ps=246000 
M3169 diff_1837000_1364000# diff_2060000_2777000# diff_83000_3098000# GND efet w=246000 l=8000
+ ad=9.26033e+08 pd=1.034e+06 as=0 ps=0 
M3170 diff_95000_5192000# diff_1837000_1364000# diff_1837000_1364000# GND efet w=18000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3171 diff_1858000_1019000# diff_1858000_1019000# diff_95000_5192000# GND efet w=18000 l=7000
+ ad=8.89033e+08 pd=964000 as=0 ps=0 
M3172 diff_83000_3098000# diff_72000_4515000# diff_1837000_1364000# GND efet w=201500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3173 diff_1858000_1019000# diff_72000_4515000# diff_83000_3098000# GND efet w=202500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3174 diff_83000_3098000# diff_2113000_2778000# diff_1858000_1019000# GND efet w=244500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3175 diff_1037000_877000# diff_1037000_877000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=-1.68967e+08 pd=718000 as=0 ps=0 
M3176 diff_1094000_1020000# diff_1094000_1020000# diff_95000_5192000# GND efet w=19000 l=9000
+ ad=-1.08297e+09 pd=620000 as=0 ps=0 
M3177 diff_83000_3098000# diff_1037000_877000# diff_1094000_1020000# GND efet w=199500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3178 diff_1037000_877000# diff_2208000_2717000# diff_83000_3098000# GND efet w=222000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3179 diff_1252000_2261000# diff_1237000_1921000# diff_95000_5192000# GND efet w=12000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3180 diff_83000_3098000# diff_1064000_2211000# diff_1176000_1643000# GND efet w=154500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3181 diff_1189000_2359000# diff_1064000_2211000# diff_83000_3098000# GND efet w=59000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3182 diff_1345000_2360000# diff_1345000_2360000# diff_95000_5192000# GND efet w=11000 l=20000
+ ad=-1.72697e+09 pd=542000 as=0 ps=0 
M3183 diff_1245000_2015000# diff_1189000_2359000# diff_1252000_2261000# GND efet w=51000 l=10000
+ ad=2.48033e+08 pd=814000 as=0 ps=0 
M3184 diff_95000_5192000# diff_1305000_2339000# diff_1305000_2339000# GND efet w=12000 l=24000
+ ad=0 pd=0 as=1.428e+09 ps=310000 
M3185 diff_1437000_2361000# diff_72000_4515000# diff_1345000_2360000# GND efet w=21000 l=11000
+ ad=2.52e+08 pd=66000 as=0 ps=0 
M3186 diff_1460000_2361000# diff_1438000_786000# diff_1437000_2361000# GND efet w=21000 l=11000
+ ad=3.91e+08 pd=112000 as=0 ps=0 
M3187 diff_1390000_2312000# diff_719000_2538000# diff_1345000_2360000# GND efet w=78500 l=7500
+ ad=1.334e+09 pd=296000 as=0 ps=0 
M3188 diff_83000_3098000# diff_1064000_2064000# diff_1176000_1643000# GND efet w=155500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3189 diff_1245000_2015000# diff_1189000_2359000# diff_1252000_2261000# GND efet w=54000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3190 diff_1305000_2339000# diff_1252000_2261000# diff_83000_3098000# GND efet w=63000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3191 diff_83000_3098000# diff_719000_2538000# diff_1305000_2339000# GND efet w=62500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3192 diff_1345000_2360000# diff_1305000_2339000# diff_83000_3098000# GND efet w=50000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3193 diff_1390000_2312000# diff_719000_2538000# diff_1345000_2360000# GND efet w=24000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3194 diff_83000_3098000# diff_1252000_2261000# diff_1390000_2312000# GND efet w=104000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3195 diff_1189000_2023000# diff_1064000_2064000# diff_83000_3098000# GND efet w=60000 l=8000
+ ad=1.319e+09 pd=274000 as=0 ps=0 
M3196 diff_1189000_2023000# diff_1189000_2023000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3197 diff_1245000_1992000# diff_1189000_2023000# diff_1245000_2015000# GND efet w=35000 l=10000
+ ad=3.86033e+08 pd=798000 as=0 ps=0 
M3198 diff_1305000_2038000# diff_1245000_2015000# diff_83000_3098000# GND efet w=62000 l=8000
+ ad=1.418e+09 pd=312000 as=0 ps=0 
M3199 diff_83000_3098000# diff_719000_2180000# diff_1305000_2038000# GND efet w=62500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3200 diff_1345000_2016000# diff_1305000_2038000# diff_83000_3098000# GND efet w=50000 l=8000
+ ad=-1.76497e+09 pd=546000 as=0 ps=0 
M3201 diff_1390000_2052000# diff_719000_2180000# diff_1345000_2016000# GND efet w=25000 l=8000
+ ad=1.328e+09 pd=292000 as=0 ps=0 
M3202 diff_83000_3098000# diff_1245000_2015000# diff_1390000_2052000# GND efet w=104000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3203 diff_1245000_2015000# diff_1237000_1921000# diff_95000_5192000# GND efet w=14000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3204 diff_1245000_1992000# diff_1189000_2023000# diff_1245000_2015000# GND efet w=71000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3205 diff_1390000_2052000# diff_719000_2180000# diff_1345000_2016000# GND efet w=75500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3206 diff_1305000_2038000# diff_1305000_2038000# diff_95000_5192000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3207 diff_95000_5192000# diff_1189000_1979000# diff_1189000_1979000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=1.423e+09 ps=276000 
M3208 diff_1245000_1992000# diff_1237000_1921000# diff_95000_5192000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3209 diff_1477000_2222000# diff_1460000_2361000# diff_83000_3098000# GND efet w=195500 l=7500
+ ad=-7.53967e+08 pd=692000 as=0 ps=0 
M3210 diff_95000_5192000# diff_1477000_2222000# diff_1477000_2222000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3211 diff_95000_5192000# diff_95000_5192000# diff_1576000_2220000# GND efet w=13000 l=33000
+ ad=0 pd=0 as=9.13e+08 ps=190000 
M3212 diff_1583000_2229000# diff_95000_5192000# diff_1556000_2304000# GND efet w=12500 l=74500
+ ad=-2.95967e+08 pd=728000 as=5.13e+08 ps=176000 
M3213 diff_95000_5192000# diff_95000_5192000# diff_1583000_2229000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3214 diff_1477000_2222000# diff_1487000_841000# diff_848000_2342000# GND efet w=108500 l=10500
+ ad=0 pd=0 as=1.51403e+09 ps=1.208e+06 
M3215 diff_1556000_2304000# diff_1547000_932000# diff_1477000_2222000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3216 diff_1477000_2074000# diff_1460000_2015000# diff_83000_3098000# GND efet w=203500 l=7500
+ ad=-7.01967e+08 pd=692000 as=0 ps=0 
M3217 diff_1477000_2074000# diff_1487000_841000# diff_848000_2016000# GND efet w=109500 l=9500
+ ad=0 pd=0 as=1.46403e+09 ps=1.2e+06 
M3218 diff_848000_2342000# diff_1643000_833000# diff_1583000_2229000# GND efet w=102500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3219 diff_1576000_2220000# diff_1556000_2304000# diff_83000_3098000# GND efet w=70500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3220 diff_1583000_2229000# diff_1576000_2220000# diff_83000_3098000# GND efet w=209000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3221 diff_817000_2342000# diff_1696000_986000# diff_1583000_2229000# GND efet w=104000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3222 diff_1583000_2155000# diff_1576000_2146000# diff_83000_3098000# GND efet w=209000 l=8000
+ ad=-2.88967e+08 pd=718000 as=0 ps=0 
M3223 diff_1576000_2146000# diff_1556000_2076000# diff_83000_3098000# GND efet w=78500 l=7500
+ ad=9.41e+08 pd=188000 as=0 ps=0 
M3224 diff_1556000_2076000# diff_1547000_932000# diff_1477000_2074000# GND efet w=18000 l=9000
+ ad=5.41e+08 pd=162000 as=0 ps=0 
M3225 diff_1345000_2016000# diff_1345000_2016000# diff_95000_5192000# GND efet w=11000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M3226 diff_1437000_2015000# diff_72000_4515000# diff_1345000_2016000# GND efet w=21000 l=12000
+ ad=2.52e+08 pd=66000 as=0 ps=0 
M3227 diff_1460000_2015000# diff_1438000_786000# diff_1437000_2015000# GND efet w=21000 l=11000
+ ad=3.96e+08 pd=102000 as=0 ps=0 
M3228 diff_83000_3098000# diff_1064000_1834000# diff_1176000_1643000# GND efet w=152500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3229 diff_1189000_1979000# diff_1064000_1834000# diff_83000_3098000# GND efet w=58000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3230 diff_1345000_1983000# diff_1345000_1983000# diff_95000_5192000# GND efet w=12000 l=20000
+ ad=-1.74497e+09 pd=540000 as=0 ps=0 
M3231 diff_1265000_1694000# diff_1189000_1979000# diff_1245000_1992000# GND efet w=53000 l=10000
+ ad=-4.81967e+08 pd=664000 as=0 ps=0 
M3232 diff_95000_5192000# diff_1305000_1962000# diff_1305000_1962000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=1.443e+09 ps=312000 
M3233 diff_1437000_1984000# diff_72000_4515000# diff_1345000_1983000# GND efet w=21000 l=12000
+ ad=2.52e+08 pd=66000 as=0 ps=0 
M3234 diff_1460000_1984000# diff_1438000_786000# diff_1437000_1984000# GND efet w=21000 l=11000
+ ad=3.92e+08 pd=112000 as=0 ps=0 
M3235 diff_1390000_1935000# diff_719000_1784000# diff_1345000_1983000# GND efet w=77500 l=7500
+ ad=1.323e+09 pd=294000 as=0 ps=0 
M3236 diff_83000_3098000# diff_1064000_1687000# diff_1176000_1643000# GND efet w=125500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3237 diff_1265000_1694000# diff_1189000_1979000# diff_1245000_1992000# GND efet w=55000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3238 diff_1202000_1633000# diff_1176000_1643000# diff_83000_3098000# GND efet w=167500 l=9500
+ ad=3.57033e+08 pd=778000 as=0 ps=0 
M3239 diff_83000_3098000# diff_1064000_1687000# diff_1176000_1643000# GND efet w=31000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M3240 diff_1305000_1962000# diff_1245000_1992000# diff_83000_3098000# GND efet w=63000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3241 diff_83000_3098000# diff_719000_1784000# diff_1305000_1962000# GND efet w=63500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3242 diff_1345000_1983000# diff_1305000_1962000# diff_83000_3098000# GND efet w=50000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3243 diff_1390000_1935000# diff_719000_1784000# diff_1345000_1983000# GND efet w=24000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3244 diff_83000_3098000# diff_1245000_1992000# diff_1390000_1935000# GND efet w=104000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3245 diff_1305000_1661000# diff_1265000_1694000# diff_83000_3098000# GND efet w=62000 l=8000
+ ad=1.416e+09 pd=310000 as=0 ps=0 
M3246 diff_83000_3098000# diff_719000_1426000# diff_1305000_1661000# GND efet w=62500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3247 diff_1345000_1639000# diff_1305000_1661000# diff_83000_3098000# GND efet w=50000 l=8000
+ ad=-1.72297e+09 pd=546000 as=0 ps=0 
M3248 diff_1390000_1674000# diff_719000_1426000# diff_1345000_1639000# GND efet w=25000 l=8000
+ ad=1.336e+09 pd=294000 as=0 ps=0 
M3249 diff_83000_3098000# diff_1265000_1694000# diff_1390000_1674000# GND efet w=104000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3250 diff_1265000_1694000# diff_1237000_1921000# diff_95000_5192000# GND efet w=12000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3251 diff_1390000_1674000# diff_719000_1426000# diff_1345000_1639000# GND efet w=76500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3252 diff_1305000_1661000# diff_1305000_1661000# diff_95000_5192000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3253 diff_95000_5192000# diff_1237000_1921000# diff_1202000_1633000# GND efet w=12000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3254 diff_889000_1530000# diff_877000_1128000# diff_856000_1595000# GND efet w=19000 l=11000
+ ad=4.18e+08 pd=82000 as=0 ps=0 
M3255 diff_914000_1456000# diff_901000_991000# diff_889000_1530000# GND efet w=19000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M3256 diff_95000_5192000# diff_123000_1243000# diff_132000_1251000# GND efet w=238500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3257 diff_123000_1453000# diff_123000_1453000# diff_95000_5192000# GND efet w=35000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3258 diff_582000_1463000# diff_680000_1019000# diff_719000_1426000# GND efet w=34000 l=11000
+ ad=5.18e+08 pd=102000 as=0 ps=0 
M3259 diff_95000_5192000# diff_123000_1243000# diff_123000_1243000# GND efet w=42000 l=9000
+ ad=0 pd=0 as=-1.2619e+09 ps=1.368e+06 
M3260 diff_132000_1251000# diff_123000_1243000# diff_95000_5192000# GND efet w=857000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3261 diff_95000_5192000# diff_123000_1243000# diff_132000_1251000# GND efet w=238500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3262 diff_83000_3098000# diff_123000_1453000# diff_123000_1243000# GND efet w=178000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3263 diff_95000_5192000# diff_123000_1243000# diff_132000_1251000# GND efet w=342000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3264 diff_83000_3098000# diff_123000_1453000# diff_123000_1243000# GND efet w=269000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3265 diff_123000_1243000# diff_553000_1211000# diff_83000_3098000# GND efet w=413500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3266 diff_95000_5192000# diff_95000_5192000# diff_817000_1286000# GND efet w=12000 l=103000
+ ad=0 pd=0 as=-1.79384e+09 ps=3.924e+06 
M3267 diff_856000_1267000# diff_848000_1262000# diff_83000_3098000# GND efet w=131000 l=8000
+ ad=1.734e+09 pd=334000 as=0 ps=0 
M3268 diff_1010000_1450000# diff_889000_1530000# diff_83000_3098000# GND efet w=37000 l=8000
+ ad=1.648e+09 pd=360000 as=0 ps=0 
M3269 diff_719000_1030000# diff_889000_1530000# diff_83000_3098000# GND efet w=47000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3270 diff_1010000_1450000# diff_889000_1530000# diff_83000_3098000# GND efet w=77000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3271 diff_1063000_1457000# diff_1037000_877000# diff_1010000_1450000# GND efet w=122000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3272 diff_1085000_1457000# diff_719000_1030000# diff_1063000_1457000# GND efet w=74500 l=8500
+ ad=1.499e+09 pd=340000 as=0 ps=0 
M3273 diff_83000_3098000# diff_1094000_1020000# diff_1085000_1457000# GND efet w=140000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3274 diff_1085000_1457000# diff_719000_1030000# diff_1063000_1457000# GND efet w=45000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3275 diff_1150000_1007000# diff_1063000_1457000# diff_83000_3098000# GND efet w=84000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3276 diff_95000_5192000# diff_1196000_1522000# diff_1196000_1522000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=1.139e+09 ps=228000 
M3277 diff_1477000_1846000# diff_1460000_1984000# diff_83000_3098000# GND efet w=195500 l=7500
+ ad=-7.01967e+08 pd=686000 as=0 ps=0 
M3278 diff_1477000_2074000# diff_1477000_2074000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3279 diff_95000_5192000# diff_1477000_1846000# diff_1477000_1846000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3280 diff_848000_2016000# diff_1643000_833000# diff_1583000_2155000# GND efet w=99000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3281 diff_83000_3098000# diff_1728000_2245000# diff_817000_2342000# GND efet w=88000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M3282 diff_817000_2040000# diff_1696000_986000# diff_1583000_2155000# GND efet w=104000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3283 diff_1576000_2146000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=33000
+ ad=0 pd=0 as=0 ps=0 
M3284 diff_1583000_2155000# diff_95000_5192000# diff_1556000_2076000# GND efet w=12500 l=79500
+ ad=0 pd=0 as=0 ps=0 
M3285 diff_1583000_2155000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3286 diff_95000_5192000# diff_95000_5192000# diff_1576000_1843000# GND efet w=13000 l=33000
+ ad=0 pd=0 as=9e+08 ps=188000 
M3287 diff_1583000_1852000# diff_95000_5192000# diff_1556000_1927000# GND efet w=12500 l=76500
+ ad=-2.42967e+08 pd=722000 as=5.21e+08 ps=174000 
M3288 diff_95000_5192000# diff_95000_5192000# diff_1583000_1852000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3289 diff_1477000_1846000# diff_1487000_841000# diff_848000_1965000# GND efet w=108500 l=10500
+ ad=0 pd=0 as=1.40403e+09 ps=1.208e+06 
M3290 diff_1556000_1927000# diff_1547000_932000# diff_1477000_1846000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3291 diff_1477000_1697000# diff_1460000_1638000# diff_83000_3098000# GND efet w=204500 l=7500
+ ad=-6.00967e+08 pd=696000 as=0 ps=0 
M3292 diff_1477000_1697000# diff_1487000_841000# diff_848000_1639000# GND efet w=109500 l=9500
+ ad=0 pd=0 as=1.40703e+09 ps=1.2e+06 
M3293 diff_83000_3098000# diff_1729000_2091000# diff_817000_2040000# GND efet w=87000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3294 diff_848000_1965000# diff_1643000_833000# diff_1583000_1852000# GND efet w=102000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3295 diff_1576000_1843000# diff_1556000_1927000# diff_83000_3098000# GND efet w=71500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3296 diff_1583000_1852000# diff_1576000_1843000# diff_83000_3098000# GND efet w=209000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3297 diff_817000_1965000# diff_1696000_986000# diff_1583000_1852000# GND efet w=103000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3298 diff_1583000_1778000# diff_1576000_1768000# diff_83000_3098000# GND efet w=209000 l=8000
+ ad=-2.11967e+08 pd=716000 as=0 ps=0 
M3299 diff_1576000_1768000# diff_1556000_1698000# diff_83000_3098000# GND efet w=78500 l=7500
+ ad=9.26e+08 pd=186000 as=0 ps=0 
M3300 diff_1556000_1698000# diff_1547000_932000# diff_1477000_1697000# GND efet w=19000 l=9000
+ ad=5.32e+08 pd=164000 as=0 ps=0 
M3301 diff_1345000_1639000# diff_1345000_1639000# diff_95000_5192000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M3302 diff_1437000_1638000# diff_72000_4515000# diff_1345000_1639000# GND efet w=21000 l=11000
+ ad=2.52e+08 pd=66000 as=0 ps=0 
M3303 diff_1460000_1638000# diff_1438000_786000# diff_1437000_1638000# GND efet w=21000 l=11000
+ ad=3.97e+08 pd=102000 as=0 ps=0 
M3304 diff_1202000_1633000# diff_1196000_1522000# diff_1236000_1424000# GND efet w=120000 l=10000
+ ad=0 pd=0 as=-3.09967e+08 ps=650000 
M3305 diff_1150000_1007000# diff_1063000_1457000# diff_83000_3098000# GND efet w=43000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M3306 diff_83000_3098000# diff_817000_1286000# diff_914000_1380000# GND efet w=141000 l=8000
+ ad=0 pd=0 as=2.042e+09 ps=434000 
M3307 diff_889000_1340000# diff_877000_1128000# diff_856000_1267000# GND efet w=19000 l=11000
+ ad=4.18e+08 pd=82000 as=0 ps=0 
M3308 diff_914000_1380000# diff_901000_991000# diff_889000_1340000# GND efet w=19000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M3309 diff_752000_680000# diff_889000_1340000# diff_83000_3098000# GND efet w=47000 l=8000
+ ad=-1.36297e+09 pd=632000 as=0 ps=0 
M3310 diff_1010000_1431000# diff_889000_1340000# diff_83000_3098000# GND efet w=80000 l=8000
+ ad=1.536e+09 pd=360000 as=0 ps=0 
M3311 diff_752000_680000# diff_889000_1340000# diff_83000_3098000# GND efet w=101500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3312 diff_132000_874000# diff_123000_1087000# diff_95000_5192000# GND efet w=858500 l=8500
+ ad=-6.78738e+08 pd=4.268e+06 as=0 ps=0 
M3313 diff_83000_3098000# diff_553000_1211000# diff_123000_1087000# GND efet w=413000 l=9000
+ ad=0 pd=0 as=-1.2839e+09 ps=1.37e+06 
M3314 diff_95000_5192000# diff_123000_1087000# diff_132000_874000# GND efet w=343000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3315 diff_95000_5192000# diff_856000_1267000# diff_856000_1267000# GND efet w=12000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3316 diff_95000_5192000# diff_123000_1087000# diff_132000_874000# GND efet w=238500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3317 diff_83000_3098000# diff_123000_866000# diff_123000_1087000# GND efet w=269000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3318 diff_83000_3098000# diff_123000_866000# diff_123000_1087000# GND efet w=180500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3319 diff_95000_5192000# diff_123000_1087000# diff_132000_874000# GND efet w=239000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3320 diff_123000_1087000# diff_123000_1087000# diff_95000_5192000# GND efet w=43000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3321 diff_856000_1218000# diff_848000_1211000# diff_83000_3098000# GND efet w=131000 l=8000
+ ad=1.733e+09 pd=324000 as=0 ps=0 
M3322 diff_95000_5192000# diff_856000_1218000# diff_856000_1218000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3323 diff_817000_1211000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=103000
+ ad=-7.65869e+08 pd=3.384e+06 as=0 ps=0 
M3324 diff_95000_5192000# diff_914000_1380000# diff_914000_1380000# GND efet w=14000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M3325 diff_1010000_1431000# diff_889000_1340000# diff_83000_3098000# GND efet w=37000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3326 diff_1063000_1310000# diff_1037000_877000# diff_1010000_1431000# GND efet w=121000 l=8000
+ ad=-1.55897e+09 pd=462000 as=0 ps=0 
M3327 diff_1085000_1346000# diff_752000_680000# diff_1063000_1310000# GND efet w=44000 l=9000
+ ad=1.514e+09 pd=334000 as=0 ps=0 
M3328 diff_83000_3098000# diff_1094000_1020000# diff_1085000_1346000# GND efet w=137500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3329 diff_1196000_1522000# diff_1063000_1457000# diff_83000_3098000# GND efet w=52000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3330 diff_1085000_1346000# diff_752000_680000# diff_1063000_1310000# GND efet w=72000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3331 diff_1150000_1007000# diff_1063000_1310000# diff_83000_3098000# GND efet w=43000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M3332 diff_1236000_1424000# diff_1188000_1277000# diff_1236000_1245000# GND efet w=119500 l=9500
+ ad=0 pd=0 as=-1.99967e+08 ps=764000 
M3333 diff_95000_5192000# diff_752000_680000# diff_752000_680000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3334 diff_95000_5192000# diff_914000_1079000# diff_914000_1079000# GND efet w=13000 l=7000
+ ad=0 pd=0 as=2.056e+09 ps=430000 
M3335 diff_709000_308000# diff_889000_1153000# diff_83000_3098000# GND efet w=104500 l=8500
+ ad=-1.07897e+09 pd=664000 as=0 ps=0 
M3336 diff_83000_3098000# diff_817000_1211000# diff_914000_1079000# GND efet w=142000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3337 diff_95000_5192000# diff_709000_308000# diff_709000_308000# GND efet w=12000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3338 diff_1063000_1310000# diff_1063000_1310000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3339 diff_1064000_1080000# diff_1064000_1080000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=-1.71897e+09 pd=454000 as=0 ps=0 
M3340 diff_1150000_1007000# diff_1063000_1310000# diff_83000_3098000# GND efet w=84000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3341 diff_889000_1153000# diff_877000_1128000# diff_856000_1218000# GND efet w=19000 l=12000
+ ad=4.18e+08 pd=82000 as=0 ps=0 
M3342 diff_914000_1079000# diff_901000_991000# diff_889000_1153000# GND efet w=19000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M3343 diff_132000_874000# diff_123000_866000# diff_83000_3098000# GND efet w=876500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3344 diff_83000_3098000# diff_123000_866000# diff_132000_874000# GND efet w=240500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3345 diff_95000_5192000# diff_123000_866000# diff_123000_866000# GND efet w=35000 l=9000
+ ad=0 pd=0 as=1.92807e+09 ps=1.272e+06 
M3346 diff_719000_1030000# diff_680000_1019000# diff_582000_964000# GND efet w=34000 l=12000
+ ad=0 pd=0 as=5.56e+08 ps=106000 
M3347 diff_83000_3098000# diff_582000_964000# diff_123000_866000# GND efet w=415000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3348 diff_83000_3098000# diff_123000_866000# diff_132000_874000# GND efet w=305500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3349 diff_123000_866000# diff_553000_1211000# diff_83000_3098000# GND efet w=415000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3350 diff_95000_5192000# diff_95000_5192000# diff_817000_909000# GND efet w=12000 l=104000
+ ad=0 pd=0 as=1.33213e+09 ps=3.646e+06 
M3351 diff_856000_890000# diff_848000_885000# diff_83000_3098000# GND efet w=131000 l=8000
+ ad=1.754e+09 pd=332000 as=0 ps=0 
M3352 diff_1010000_1073000# diff_889000_1153000# diff_83000_3098000# GND efet w=38000 l=8000
+ ad=1.621e+09 pd=360000 as=0 ps=0 
M3353 diff_709000_308000# diff_889000_1153000# diff_83000_3098000# GND efet w=48000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3354 diff_1010000_1073000# diff_889000_1153000# diff_83000_3098000# GND efet w=77500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3355 diff_1064000_1080000# diff_1037000_877000# diff_1010000_1073000# GND efet w=122000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3356 diff_1085000_1080000# diff_709000_308000# diff_1064000_1080000# GND efet w=74500 l=8500
+ ad=1.498e+09 pd=340000 as=0 ps=0 
M3357 diff_83000_3098000# diff_1094000_1020000# diff_1085000_1080000# GND efet w=140500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3358 diff_1085000_1080000# diff_709000_308000# diff_1064000_1080000# GND efet w=45000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3359 diff_1150000_1007000# diff_1064000_1080000# diff_83000_3098000# GND efet w=84000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3360 diff_1150000_1007000# diff_1064000_1080000# diff_83000_3098000# GND efet w=43000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M3361 diff_83000_3098000# diff_817000_909000# diff_914000_1003000# GND efet w=141000 l=8000
+ ad=0 pd=0 as=2.091e+09 ps=432000 
M3362 diff_889000_963000# diff_877000_1128000# diff_856000_890000# GND efet w=19000 l=11000
+ ad=4.18e+08 pd=82000 as=0 ps=0 
M3363 diff_914000_1003000# diff_901000_991000# diff_889000_963000# GND efet w=19000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M3364 diff_970000_884000# diff_889000_963000# diff_83000_3098000# GND efet w=47000 l=8000
+ ad=4.68033e+08 pd=954000 as=0 ps=0 
M3365 diff_1010000_1054000# diff_889000_963000# diff_83000_3098000# GND efet w=80000 l=8000
+ ad=1.536e+09 pd=360000 as=0 ps=0 
M3366 diff_970000_884000# diff_889000_963000# diff_83000_3098000# GND efet w=102000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3367 diff_95000_5192000# diff_856000_890000# diff_856000_890000# GND efet w=12000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3368 diff_132000_496000# diff_123000_700000# diff_83000_3098000# GND efet w=879500 l=8500
+ ad=-1.01674e+09 pd=4.216e+06 as=0 ps=0 
M3369 diff_83000_3098000# diff_123000_700000# diff_132000_496000# GND efet w=304500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3370 diff_83000_3098000# diff_553000_1211000# diff_123000_700000# GND efet w=407000 l=9000
+ ad=0 pd=0 as=2.05007e+09 ps=1.266e+06 
M3371 diff_95000_5192000# diff_914000_1003000# diff_914000_1003000# GND efet w=13000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M3372 diff_1010000_1054000# diff_889000_963000# diff_83000_3098000# GND efet w=37000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3373 diff_1064000_933000# diff_1037000_877000# diff_1010000_1054000# GND efet w=121000 l=9000
+ ad=-1.71897e+09 pd=460000 as=0 ps=0 
M3374 diff_1085000_969000# diff_970000_884000# diff_1064000_933000# GND efet w=44000 l=9000
+ ad=1.513e+09 pd=334000 as=0 ps=0 
M3375 diff_83000_3098000# diff_1094000_1020000# diff_1085000_969000# GND efet w=137000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3376 diff_1085000_969000# diff_970000_884000# diff_1064000_933000# GND efet w=72000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3377 diff_1150000_1007000# diff_1064000_933000# diff_83000_3098000# GND efet w=43000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M3378 diff_1188000_1277000# diff_1063000_1310000# diff_83000_3098000# GND efet w=50500 l=7500
+ ad=1.754e+09 pd=396000 as=0 ps=0 
M3379 diff_1188000_1277000# diff_1188000_1277000# diff_95000_5192000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M3380 diff_1345000_1606000# diff_1345000_1606000# diff_95000_5192000# GND efet w=12000 l=20000
+ ad=-1.71897e+09 pd=542000 as=0 ps=0 
M3381 diff_95000_5192000# diff_1305000_1585000# diff_1305000_1585000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=1.449e+09 ps=312000 
M3382 diff_1437000_1607000# diff_72000_4515000# diff_1345000_1606000# GND efet w=21000 l=11000
+ ad=2.52e+08 pd=66000 as=0 ps=0 
M3383 diff_1460000_1607000# diff_1438000_786000# diff_1437000_1607000# GND efet w=21000 l=11000
+ ad=4e+08 pd=110000 as=0 ps=0 
M3384 diff_1390000_1558000# diff_719000_1030000# diff_1345000_1606000# GND efet w=77500 l=7500
+ ad=1.323e+09 pd=294000 as=0 ps=0 
M3385 diff_1305000_1585000# diff_1202000_1633000# diff_83000_3098000# GND efet w=63000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3386 diff_83000_3098000# diff_719000_1030000# diff_1305000_1585000# GND efet w=62500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3387 diff_1345000_1606000# diff_1305000_1585000# diff_83000_3098000# GND efet w=49000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3388 diff_1390000_1558000# diff_719000_1030000# diff_1345000_1606000# GND efet w=24000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3389 diff_83000_3098000# diff_1202000_1633000# diff_1390000_1558000# GND efet w=104000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3390 diff_1305000_1284000# diff_1236000_1424000# diff_83000_3098000# GND efet w=62000 l=8000
+ ad=1.416e+09 pd=310000 as=0 ps=0 
M3391 diff_83000_3098000# diff_752000_680000# diff_1305000_1284000# GND efet w=62500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3392 diff_1345000_1262000# diff_1305000_1284000# diff_83000_3098000# GND efet w=49000 l=8000
+ ad=-1.74397e+09 pd=546000 as=0 ps=0 
M3393 diff_1390000_1297000# diff_752000_680000# diff_1345000_1262000# GND efet w=25000 l=8000
+ ad=1.337e+09 pd=294000 as=0 ps=0 
M3394 diff_83000_3098000# diff_1236000_1424000# diff_1390000_1297000# GND efet w=104000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3395 diff_1390000_1297000# diff_752000_680000# diff_1345000_1262000# GND efet w=76500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3396 diff_1236000_1424000# diff_1237000_1921000# diff_95000_5192000# GND efet w=13000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3397 diff_1305000_1284000# diff_1305000_1284000# diff_95000_5192000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3398 diff_95000_5192000# diff_1237000_1921000# diff_1236000_1245000# GND efet w=12000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3399 diff_1477000_1468000# diff_1460000_1607000# diff_83000_3098000# GND efet w=195500 l=7500
+ ad=-7.69967e+08 pd=688000 as=0 ps=0 
M3400 diff_1477000_1697000# diff_1477000_1697000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3401 diff_95000_5192000# diff_1477000_1468000# diff_1477000_1468000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3402 diff_848000_1639000# diff_1643000_833000# diff_1583000_1778000# GND efet w=98500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3403 diff_83000_3098000# diff_1729000_1868000# diff_817000_1965000# GND efet w=87000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3404 diff_817000_1663000# diff_1696000_986000# diff_1583000_1778000# GND efet w=105000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3405 diff_1576000_1768000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=34000
+ ad=0 pd=0 as=0 ps=0 
M3406 diff_1583000_1778000# diff_95000_5192000# diff_1556000_1698000# GND efet w=12500 l=81500
+ ad=0 pd=0 as=0 ps=0 
M3407 diff_1583000_1778000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3408 diff_95000_5192000# diff_95000_5192000# diff_1576000_1466000# GND efet w=13000 l=32000
+ ad=0 pd=0 as=9.13e+08 ps=190000 
M3409 diff_1583000_1475000# diff_95000_5192000# diff_1557000_1550000# GND efet w=12500 l=74500
+ ad=-2.18967e+08 pd=726000 as=5.1e+08 ps=172000 
M3410 diff_95000_5192000# diff_95000_5192000# diff_1583000_1475000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3411 diff_1477000_1468000# diff_1487000_841000# diff_848000_1588000# GND efet w=108000 l=10000
+ ad=0 pd=0 as=1.55403e+09 ps=1.208e+06 
M3412 diff_1557000_1550000# diff_1547000_932000# diff_1477000_1468000# GND efet w=18000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3413 diff_1477000_1320000# diff_1460000_1261000# diff_83000_3098000# GND efet w=203500 l=7500
+ ad=-6.88967e+08 pd=694000 as=0 ps=0 
M3414 diff_1477000_1320000# diff_1487000_841000# diff_848000_1262000# GND efet w=110500 l=9500
+ ad=0 pd=0 as=1.50503e+09 ps=1.2e+06 
M3415 diff_848000_1588000# diff_1643000_833000# diff_1583000_1475000# GND efet w=102000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3416 diff_1576000_1466000# diff_1557000_1550000# diff_83000_3098000# GND efet w=71500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3417 diff_1583000_1475000# diff_1576000_1466000# diff_83000_3098000# GND efet w=209000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3418 diff_817000_1588000# diff_1696000_986000# diff_1583000_1475000# GND efet w=103000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3419 diff_1583000_1401000# diff_1576000_1391000# diff_83000_3098000# GND efet w=209000 l=8000
+ ad=-1.52967e+08 pd=716000 as=0 ps=0 
M3420 diff_1576000_1391000# diff_1557000_1321000# diff_83000_3098000# GND efet w=78500 l=7500
+ ad=9.26e+08 pd=186000 as=0 ps=0 
M3421 diff_1557000_1321000# diff_1547000_932000# diff_1477000_1320000# GND efet w=19000 l=10000
+ ad=5.14e+08 pd=162000 as=0 ps=0 
M3422 diff_1345000_1262000# diff_1345000_1262000# diff_95000_5192000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M3423 diff_1437000_1261000# diff_72000_4515000# diff_1345000_1262000# GND efet w=21000 l=12000
+ ad=2.52e+08 pd=66000 as=0 ps=0 
M3424 diff_1460000_1261000# diff_1438000_786000# diff_1437000_1261000# GND efet w=21000 l=11000
+ ad=3.96e+08 pd=102000 as=0 ps=0 
M3425 diff_95000_5192000# diff_1188000_1219000# diff_1188000_1219000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=1.316e+09 ps=280000 
M3426 diff_1345000_1229000# diff_1345000_1229000# diff_95000_5192000# GND efet w=11000 l=20000
+ ad=-1.73997e+09 pd=540000 as=0 ps=0 
M3427 diff_1188000_1219000# diff_1064000_1080000# diff_83000_3098000# GND efet w=49000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3428 diff_1236000_1245000# diff_1188000_1219000# diff_1238000_975000# GND efet w=114000 l=9000
+ ad=0 pd=0 as=-1.91397e+09 ps=508000 
M3429 diff_95000_5192000# diff_1305000_1208000# diff_1305000_1208000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=1.448e+09 ps=312000 
M3430 diff_1437000_1230000# diff_72000_4515000# diff_1345000_1229000# GND efet w=21000 l=12000
+ ad=2.52e+08 pd=66000 as=0 ps=0 
M3431 diff_1460000_1230000# diff_1438000_786000# diff_1437000_1230000# GND efet w=21000 l=11000
+ ad=3.99e+08 pd=110000 as=0 ps=0 
M3432 diff_95000_5192000# diff_970000_884000# diff_970000_884000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3433 diff_83000_3098000# diff_582000_709000# diff_123000_700000# GND efet w=414000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3434 diff_83000_3098000# diff_123000_700000# diff_132000_496000# GND efet w=240500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3435 diff_95000_5192000# diff_123000_488000# diff_132000_496000# GND efet w=239000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3436 diff_123000_700000# diff_123000_700000# diff_95000_5192000# GND efet w=36000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3437 diff_752000_680000# diff_680000_1019000# diff_582000_709000# GND efet w=35000 l=11000
+ ad=0 pd=0 as=4.9e+08 ps=112000 
M3438 diff_95000_5192000# diff_123000_488000# diff_123000_488000# GND efet w=41000 l=9000
+ ad=0 pd=0 as=-1.1129e+09 ps=1.406e+06 
M3439 diff_83000_3098000# diff_72000_4515000# diff_877000_1128000# GND efet w=77000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3440 diff_901000_991000# diff_72000_4515000# diff_83000_3098000# GND efet w=77000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3441 diff_1064000_933000# diff_1064000_933000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3442 diff_1150000_1007000# diff_1064000_933000# diff_83000_3098000# GND efet w=84000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3443 diff_95000_5192000# diff_1150000_1007000# diff_1150000_1007000# GND efet w=12000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M3444 diff_95000_5192000# diff_123000_488000# diff_132000_496000# GND efet w=238000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3445 diff_83000_3098000# diff_553000_1211000# diff_123000_488000# GND efet w=364500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3446 diff_132000_496000# diff_123000_488000# diff_95000_5192000# GND efet w=828500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3447 diff_95000_5192000# diff_123000_488000# diff_132000_496000# GND efet w=343000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3448 diff_123000_488000# diff_553000_1211000# diff_83000_3098000# GND efet w=38000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3449 diff_123000_488000# diff_123000_700000# diff_83000_3098000# GND efet w=81000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3450 diff_83000_3098000# diff_553000_1211000# diff_792000_356000# GND efet w=401500 l=7500
+ ad=0 pd=0 as=4.71065e+08 ps=1.348e+06 
M3451 diff_83000_3098000# diff_906000_615000# diff_792000_356000# GND efet w=407500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3452 diff_83000_3098000# diff_123000_700000# diff_123000_488000# GND efet w=381000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M3453 diff_970000_884000# diff_680000_1019000# diff_906000_615000# GND efet w=34000 l=12000
+ ad=0 pd=0 as=5e+08 ps=130000 
M3454 diff_1390000_1180000# diff_709000_308000# diff_1345000_1229000# GND efet w=77500 l=7500
+ ad=1.336e+09 pd=296000 as=0 ps=0 
M3455 diff_1305000_1208000# diff_1236000_1245000# diff_83000_3098000# GND efet w=63000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3456 diff_83000_3098000# diff_709000_308000# diff_1305000_1208000# GND efet w=62500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3457 diff_1345000_1229000# diff_1305000_1208000# diff_83000_3098000# GND efet w=49000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3458 diff_1390000_1180000# diff_709000_308000# diff_1345000_1229000# GND efet w=25000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3459 diff_83000_3098000# diff_1236000_1245000# diff_1390000_1180000# GND efet w=105000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3460 diff_95000_5192000# diff_1237000_1921000# diff_1238000_975000# GND efet w=13000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3461 diff_1305000_907000# diff_1238000_975000# diff_83000_3098000# GND efet w=62000 l=8000
+ ad=1.432e+09 pd=314000 as=0 ps=0 
M3462 diff_83000_3098000# diff_970000_884000# diff_1305000_907000# GND efet w=62500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3463 diff_1345000_885000# diff_1305000_907000# diff_83000_3098000# GND efet w=49000 l=8000
+ ad=-1.80297e+09 pd=548000 as=0 ps=0 
M3464 diff_1390000_920000# diff_970000_884000# diff_1345000_885000# GND efet w=24000 l=8000
+ ad=1.328e+09 pd=292000 as=0 ps=0 
M3465 diff_83000_3098000# diff_1238000_975000# diff_1390000_920000# GND efet w=103000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3466 diff_1390000_920000# diff_970000_884000# diff_1345000_885000# GND efet w=76500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3467 diff_1305000_907000# diff_1305000_907000# diff_95000_5192000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3468 diff_1477000_1091000# diff_1460000_1230000# diff_83000_3098000# GND efet w=194500 l=7500
+ ad=-7.88967e+08 pd=686000 as=0 ps=0 
M3469 diff_1477000_1320000# diff_1477000_1320000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3470 diff_95000_5192000# diff_1477000_1091000# diff_1477000_1091000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3471 diff_848000_1262000# diff_1643000_833000# diff_1583000_1401000# GND efet w=98500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3472 diff_817000_1286000# diff_1696000_986000# diff_1583000_1401000# GND efet w=105000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3473 diff_1576000_1391000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=34000
+ ad=0 pd=0 as=0 ps=0 
M3474 diff_1583000_1401000# diff_95000_5192000# diff_1557000_1321000# GND efet w=12500 l=80500
+ ad=0 pd=0 as=0 ps=0 
M3475 diff_1583000_1401000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3476 diff_95000_5192000# diff_95000_5192000# diff_1576000_1089000# GND efet w=13000 l=32000
+ ad=0 pd=0 as=9.14e+08 ps=190000 
M3477 diff_1583000_1098000# diff_95000_5192000# diff_1556000_1173000# GND efet w=12500 l=75500
+ ad=-2.37967e+08 pd=724000 as=5.33e+08 ps=176000 
M3478 diff_95000_5192000# diff_95000_5192000# diff_1583000_1098000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3479 diff_1477000_1091000# diff_1487000_841000# diff_848000_1211000# GND efet w=108000 l=10000
+ ad=0 pd=0 as=1.51203e+09 ps=1.204e+06 
M3480 diff_1556000_1173000# diff_1547000_932000# diff_1477000_1091000# GND efet w=18000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3481 diff_1477000_942000# diff_1460000_884000# diff_83000_3098000# GND efet w=202500 l=7500
+ ad=-6.95967e+08 pd=694000 as=0 ps=0 
M3482 diff_1477000_942000# diff_1487000_841000# diff_848000_885000# GND efet w=110000 l=10000
+ ad=0 pd=0 as=1.46203e+09 ps=1.2e+06 
M3483 diff_848000_1211000# diff_1643000_833000# diff_1583000_1098000# GND efet w=100500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3484 diff_1576000_1089000# diff_1556000_1173000# diff_83000_3098000# GND efet w=71500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3485 diff_1583000_1098000# diff_1576000_1089000# diff_83000_3098000# GND efet w=208000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3486 diff_817000_1211000# diff_1696000_986000# diff_1583000_1098000# GND efet w=103000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3487 diff_1583000_1024000# diff_1576000_1014000# diff_83000_3098000# GND efet w=209000 l=8000
+ ad=-1.37967e+08 pd=722000 as=0 ps=0 
M3488 diff_1576000_1014000# diff_1556000_944000# diff_83000_3098000# GND efet w=78500 l=7500
+ ad=9.38e+08 pd=188000 as=0 ps=0 
M3489 diff_1556000_944000# diff_1547000_932000# diff_1477000_942000# GND efet w=18000 l=9000
+ ad=5.37e+08 pd=160000 as=0 ps=0 
M3490 diff_1345000_885000# diff_1345000_885000# diff_95000_5192000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M3491 diff_1437000_884000# diff_72000_4515000# diff_1345000_885000# GND efet w=20000 l=11000
+ ad=2.4e+08 pd=64000 as=0 ps=0 
M3492 diff_1460000_884000# diff_1438000_786000# diff_1437000_884000# GND efet w=20000 l=11000
+ ad=3.9e+08 pd=98000 as=0 ps=0 
M3493 diff_1477000_942000# diff_1477000_942000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3494 diff_1237000_1921000# diff_72000_4515000# diff_83000_3098000# GND efet w=72000 l=10000
+ ad=-1.33593e+09 pd=1.116e+06 as=0 ps=0 
M3495 diff_848000_885000# diff_1643000_833000# diff_1583000_1024000# GND efet w=99000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3496 diff_817000_909000# diff_1696000_986000# diff_1583000_1024000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3497 diff_1576000_1014000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=32000
+ ad=0 pd=0 as=0 ps=0 
M3498 diff_1583000_1024000# diff_95000_5192000# diff_1556000_944000# GND efet w=12500 l=79500
+ ad=0 pd=0 as=0 ps=0 
M3499 diff_1583000_1024000# diff_95000_5192000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3500 diff_1438000_786000# diff_1386000_841000# diff_83000_3098000# GND efet w=72000 l=9000
+ ad=1.81807e+09 pd=1.662e+06 as=0 ps=0 
M3501 diff_83000_3098000# diff_72000_4515000# diff_1487000_841000# GND efet w=75000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3502 diff_1547000_932000# diff_72000_4515000# diff_83000_3098000# GND efet w=75000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3503 diff_83000_3098000# diff_72000_4515000# diff_1643000_833000# GND efet w=70000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3504 diff_1696000_986000# diff_72000_4515000# diff_83000_3098000# GND efet w=70000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3505 diff_1237000_1921000# diff_1237000_1921000# diff_95000_5192000# GND efet w=17000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3506 diff_95000_5192000# diff_2288000_2488000# diff_2288000_2488000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=2.135e+09 ps=404000 
M3507 diff_95000_5192000# diff_2304000_1746000# diff_2304000_1746000# GND efet w=12000 l=8000
+ ad=0 pd=0 as=-3.07869e+08 ps=2.872e+06 
M3508 diff_83000_3098000# diff_2288000_2488000# diff_2127000_2299000# GND efet w=135000 l=10000
+ ad=0 pd=0 as=1.04703e+09 ps=1.004e+06 
M3509 diff_2288000_2488000# diff_1237000_1921000# diff_83000_3098000# GND efet w=67500 l=6500
+ ad=0 pd=0 as=0 ps=0 
M3510 diff_83000_3098000# diff_1276000_2574000# diff_2288000_2488000# GND efet w=68000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3511 diff_2304000_1746000# diff_1276000_2574000# diff_83000_3098000# GND efet w=179500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3512 diff_83000_3098000# diff_1237000_1921000# diff_2304000_1746000# GND efet w=172000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3513 diff_1237000_1921000# diff_72000_4515000# diff_83000_3098000# GND efet w=199000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3514 diff_991000_3076000# diff_72000_4515000# diff_2529000_2777000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=9.43e+08 ps=154000 
M3515 diff_83000_3098000# diff_2962000_3296000# diff_2938000_3467000# GND efet w=62000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3516 diff_83000_3098000# diff_3017000_3539000# diff_2986000_3296000# GND efet w=42000 l=9000
+ ad=0 pd=0 as=-1.70797e+09 ps=576000 
M3517 diff_3014000_3475000# diff_3048000_3539000# diff_83000_3098000# GND efet w=79000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3518 diff_531000_4622000# diff_531000_4622000# diff_531000_4622000# GND efet w=2000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M3519 diff_3325000_3886000# diff_68000_5288000# diff_3212000_3556000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=7.75e+08 ps=222000 
M3520 diff_95000_5192000# diff_531000_4622000# diff_531000_4622000# GND efet w=24000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M3521 diff_3325000_3886000# diff_3325000_3886000# diff_95000_5192000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3522 diff_3413000_3852000# diff_2606000_4947000# diff_1698000_2848000# GND efet w=203000 l=8000
+ ad=1.827e+09 pd=424000 as=0 ps=0 
M3523 diff_83000_3098000# diff_597000_3013000# diff_3413000_3852000# GND efet w=203000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3524 diff_1698000_2848000# diff_1698000_2848000# diff_95000_5192000# GND efet w=12000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M3525 diff_83000_3098000# diff_3212000_3556000# diff_531000_4622000# GND efet w=268500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3526 diff_2938000_3467000# diff_2938000_3467000# diff_95000_5192000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M3527 diff_3401000_3461000# diff_3401000_3461000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3528 diff_3014000_3475000# diff_3014000_3475000# diff_95000_5192000# GND efet w=12000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M3529 diff_2986000_3296000# diff_2986000_3296000# diff_95000_5192000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M3530 diff_83000_3098000# diff_3033000_4154000# diff_2988000_3091000# GND efet w=72000 l=8000
+ ad=0 pd=0 as=1.363e+09 ps=308000 
M3531 diff_3113000_3386000# diff_3106000_3438000# diff_83000_3098000# GND efet w=67000 l=9000
+ ad=1.403e+09 pd=296000 as=0 ps=0 
M3532 diff_83000_3098000# diff_784000_3633000# diff_3113000_3386000# GND efet w=79000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3533 diff_3754000_4644000# diff_791000_4022000# diff_3700000_4748000# GND efet w=83000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M3534 diff_83000_3098000# diff_3625000_4962000# diff_3754000_4644000# GND efet w=89000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3535 diff_3664000_4488000# diff_3507000_4962000# diff_83000_3098000# GND efet w=148000 l=8000
+ ad=2.46033e+08 pd=820000 as=0 ps=0 
M3536 diff_3700000_4748000# diff_3700000_4748000# diff_95000_5192000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M3537 diff_95000_5192000# diff_3667000_4701000# diff_3667000_4701000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=-2.13997e+09 ps=476000 
M3538 diff_3664000_4488000# diff_791000_4022000# diff_3667000_4701000# GND efet w=151500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M3539 diff_3607000_4424000# diff_3419000_4962000# diff_83000_3098000# GND efet w=159000 l=8000
+ ad=-5.81967e+08 pd=720000 as=0 ps=0 
M3540 diff_83000_3098000# diff_3447000_4962000# diff_3607000_4424000# GND efet w=154500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3541 diff_83000_3098000# diff_3537000_4962000# diff_3664000_4488000# GND efet w=134500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3542 diff_83000_3098000# diff_3477000_4962000# diff_3658000_4142000# GND efet w=60500 l=8500
+ ad=0 pd=0 as=1.092e+09 ps=266000 
M3543 diff_3658000_4142000# diff_3658000_4142000# diff_95000_5192000# GND efet w=13000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M3544 diff_3666000_4149000# diff_3658000_4142000# diff_3607000_4424000# GND efet w=132000 l=8000
+ ad=1.32e+09 pd=284000 as=0 ps=0 
M3545 diff_3666000_4069000# diff_791000_4022000# diff_3666000_4149000# GND efet w=132000 l=8000
+ ad=-1.89097e+09 pd=478000 as=0 ps=0 
M3546 diff_95000_5192000# diff_3666000_4069000# diff_3666000_4069000# GND efet w=13000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M3547 diff_3535000_3825000# diff_68000_5288000# diff_3583000_4085000# GND efet w=13000 l=12000
+ ad=-8.39967e+08 pd=752000 as=2.4e+08 ps=92000 
M3548 diff_83000_3098000# diff_3448000_3517000# diff_3535000_3825000# GND efet w=65500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3549 diff_784000_3633000# diff_3583000_4085000# diff_83000_3098000# GND efet w=101000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3550 diff_3448000_3517000# diff_72000_4515000# diff_2570000_3912000# GND efet w=19000 l=11000
+ ad=-1.91097e+09 pd=492000 as=-4.47967e+08 ps=804000 
M3551 diff_946000_3261000# diff_72000_4515000# diff_3677000_3847000# GND efet w=13000 l=10000
+ ad=0 pd=0 as=2.75e+08 ps=90000 
M3552 diff_83000_3098000# diff_3623000_3886000# diff_2570000_3912000# GND efet w=64000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3553 diff_3668000_3852000# diff_3532000_3485000# diff_3619000_3826000# GND efet w=144000 l=8000
+ ad=1.383e+09 pd=308000 as=2.037e+09 ps=472000 
M3554 diff_2988000_3091000# diff_2988000_3091000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3555 diff_3113000_3386000# diff_3113000_3386000# diff_95000_5192000# GND efet w=14000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3556 diff_2735000_2818000# diff_2744000_3026000# diff_83000_3098000# GND efet w=85000 l=8000
+ ad=1.986e+09 pd=466000 as=0 ps=0 
M3557 diff_83000_3098000# diff_860000_2987000# diff_2735000_2818000# GND efet w=77000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3558 diff_2819000_3094000# diff_531000_4622000# diff_83000_3098000# GND efet w=132000 l=9000
+ ad=1.056e+09 pd=280000 as=0 ps=0 
M3559 diff_2808000_2818000# diff_512000_4352000# diff_2819000_3094000# GND efet w=132000 l=9000
+ ad=-1.66797e+09 pd=528000 as=0 ps=0 
M3560 diff_2744000_3026000# diff_68000_5288000# diff_1000000_2990000# GND efet w=12000 l=11000
+ ad=2.58e+08 pd=82000 as=0 ps=0 
M3561 diff_2735000_2818000# diff_2735000_2818000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3562 diff_2808000_2818000# diff_2808000_2818000# diff_95000_5192000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3563 diff_2986000_3296000# diff_68000_5288000# diff_2962000_3296000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=4.44e+08 ps=124000 
M3564 diff_2907000_3149000# diff_68000_5288000# diff_2874000_3145000# GND efet w=12000 l=12000
+ ad=1.641e+09 pd=344000 as=2.46e+08 ps=90000 
M3565 diff_83000_3098000# diff_2874000_3145000# diff_2602000_2818000# GND efet w=72000 l=8000
+ ad=0 pd=0 as=-2.09397e+09 ps=496000 
M3566 diff_2911000_2818000# diff_72000_4515000# diff_2922000_3078000# GND efet w=13000 l=11000
+ ad=-1.45497e+09 pd=606000 as=2.3e+08 ps=70000 
M3567 diff_83000_3098000# diff_2922000_3078000# diff_2907000_3149000# GND efet w=67500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3568 diff_2978000_3080000# diff_743000_2974000# diff_2911000_2818000# GND efet w=136000 l=8000
+ ad=1.552e+09 pd=338000 as=0 ps=0 
M3569 diff_83000_3098000# diff_2988000_3091000# diff_2978000_3080000# GND efet w=140500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3570 diff_3024000_3075000# diff_94000_3158000# diff_83000_3098000# GND efet w=134500 l=8500
+ ad=1.125e+09 pd=286000 as=0 ps=0 
M3571 diff_2907000_3149000# diff_2907000_3149000# diff_95000_5192000# GND efet w=13000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M3572 diff_2632000_2818000# diff_2988000_3091000# diff_3024000_3075000# GND efet w=133500 l=8500
+ ad=-7.01967e+08 pd=684000 as=0 ps=0 
M3573 diff_3072000_3193000# diff_72000_4515000# diff_2632000_2818000# GND efet w=13000 l=12000
+ ad=2.61e+08 pd=88000 as=0 ps=0 
M3574 diff_3122000_3080000# diff_68000_5288000# diff_3061000_3052000# GND efet w=12000 l=11000
+ ad=5.65e+08 pd=134000 as=-2.02397e+09 ps=414000 
M3575 diff_3061000_3052000# diff_3072000_3193000# diff_83000_3098000# GND efet w=63000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3576 diff_3535000_3825000# diff_3535000_3825000# diff_95000_5192000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M3577 diff_83000_3098000# diff_3677000_3847000# diff_3668000_3852000# GND efet w=144000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3578 diff_3619000_3826000# diff_68000_5288000# diff_3623000_3886000# GND efet w=11000 l=11000
+ ad=0 pd=0 as=4.33e+08 ps=130000 
M3579 diff_4020000_4533000# diff_3840000_4962000# diff_83000_3098000# GND efet w=88500 l=8500
+ ad=-1.80497e+09 pd=478000 as=0 ps=0 
M3580 diff_83000_3098000# diff_3870000_4934000# diff_4020000_4533000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3581 diff_95000_5192000# diff_3981000_4517000# diff_3981000_4517000# GND efet w=13000 l=36000
+ ad=0 pd=0 as=1.66903e+09 ps=1.266e+06 
M3582 diff_3981000_4517000# diff_1001000_4394000# diff_4020000_4533000# GND efet w=89500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3583 diff_3887000_4604000# diff_68000_5288000# diff_3909000_4369000# GND efet w=14000 l=11000
+ ad=2.48e+08 pd=76000 as=1.75e+09 ps=434000 
M3584 diff_784000_3633000# diff_784000_3633000# diff_95000_5192000# GND efet w=12000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M3585 diff_3619000_3826000# diff_3619000_3826000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3586 diff_95000_5192000# diff_2570000_3912000# diff_2570000_3912000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3587 diff_83000_3098000# diff_94000_3551000# diff_3448000_3517000# GND efet w=65500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M3588 diff_3645000_3521000# diff_791000_4022000# diff_3444000_3167000# GND efet w=146000 l=9000
+ ad=1.314e+09 pd=310000 as=-1.64297e+09 ps=570000 
M3589 diff_83000_3098000# diff_3569000_3530000# diff_3532000_3485000# GND efet w=81500 l=8500
+ ad=0 pd=0 as=1.567e+09 ps=272000 
M3590 diff_3444000_3167000# diff_3444000_3167000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3591 diff_83000_3098000# diff_3654000_3515000# diff_3645000_3521000# GND efet w=146000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3592 diff_3488000_4662000# diff_72000_4515000# diff_3702000_3518000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.43e+08 ps=88000 
M3593 diff_83000_3098000# diff_3887000_4604000# diff_3981000_4517000# GND efet w=43500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3594 diff_83000_3098000# diff_3014000_3475000# diff_3981000_4517000# GND efet w=42000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3595 diff_4126000_4460000# diff_3957000_4962000# diff_83000_3098000# GND efet w=149500 l=9500
+ ad=-9.35967e+08 pd=658000 as=0 ps=0 
M3596 diff_4175000_4495000# diff_4017000_4962000# diff_83000_3098000# GND efet w=135000 l=9000
+ ad=-4.59967e+08 pd=752000 as=0 ps=0 
M3597 diff_83000_3098000# diff_4047000_4930000# diff_4175000_4495000# GND efet w=134000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3598 diff_4125000_2818000# diff_4075000_4962000# diff_83000_3098000# GND efet w=67000 l=10000
+ ad=6.18033e+08 pd=848000 as=0 ps=0 
M3599 diff_83000_3098000# diff_4323000_4962000# diff_4382000_4593000# GND efet w=59500 l=8500
+ ad=0 pd=0 as=1.798e+09 ps=344000 
M3600 diff_83000_3098000# diff_4293000_4962000# diff_4382000_4593000# GND efet w=42000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3601 diff_83000_3098000# diff_3987000_4962000# diff_4126000_4460000# GND efet w=140500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3602 diff_4175000_4495000# diff_3987000_4962000# diff_83000_3098000# GND efet w=148500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3603 diff_4066000_4315000# diff_3899000_4962000# diff_83000_3098000# GND efet w=86500 l=8500
+ ad=1.095e+09 pd=222000 as=0 ps=0 
M3604 diff_3981000_4517000# diff_530000_4372000# diff_4066000_4315000# GND efet w=85000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3605 diff_3939000_3886000# diff_791000_4022000# diff_2971000_4656000# GND efet w=130000 l=8000
+ ad=1.17e+09 pd=278000 as=-9.77967e+08 ps=626000 
M3606 diff_83000_3098000# diff_3781000_4962000# diff_3939000_3886000# GND efet w=130000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3607 diff_3909000_4369000# diff_3944000_3772000# diff_83000_3098000# GND efet w=45500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3608 diff_2971000_4656000# diff_2971000_4656000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3609 diff_3909000_4369000# diff_3909000_4369000# diff_95000_5192000# GND efet w=12000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M3610 diff_3944000_3772000# diff_72000_4515000# diff_2971000_4656000# GND efet w=13000 l=11000
+ ad=2.25e+08 pd=80000 as=0 ps=0 
M3611 diff_83000_3098000# diff_2860000_4570000# diff_2351000_3074000# GND efet w=205000 l=9000
+ ad=0 pd=0 as=-8.13935e+08 ps=1.306e+06 
M3612 diff_3791000_3500000# diff_3683000_4962000# diff_83000_3098000# GND efet w=143000 l=9000
+ ad=1.594e+09 pd=310000 as=0 ps=0 
M3613 diff_83000_3098000# diff_3122000_3080000# diff_2941000_2818000# GND efet w=64000 l=8000
+ ad=0 pd=0 as=1.445e+09 ps=368000 
M3614 diff_3050000_2818000# diff_3113000_3386000# diff_83000_3098000# GND efet w=79500 l=7500
+ ad=2.109e+09 pd=460000 as=0 ps=0 
M3615 diff_3231000_3142000# diff_530000_4372000# diff_3014000_2818000# GND efet w=131000 l=9000
+ ad=1.179e+09 pd=280000 as=-2.61935e+08 ps=1.442e+06 
M3616 diff_83000_3098000# diff_512000_4352000# diff_3231000_3142000# GND efet w=131000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3617 diff_3282000_3144000# diff_3272000_3283000# diff_83000_3098000# GND efet w=129000 l=7000
+ ad=1.29e+09 pd=278000 as=0 ps=0 
M3618 diff_3014000_2818000# diff_519000_3032000# diff_3282000_3144000# GND efet w=129000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3619 diff_83000_3098000# diff_3174000_4962000# diff_3187000_3099000# GND efet w=144500 l=8500
+ ad=0 pd=0 as=1.856e+09 ps=424000 
M3620 diff_3187000_3099000# diff_906000_3226000# diff_3014000_2818000# GND efet w=140000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3621 diff_95000_5192000# diff_2602000_2818000# diff_2602000_2818000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3622 diff_3061000_3052000# diff_3061000_3052000# diff_95000_5192000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M3623 diff_2941000_2818000# diff_2941000_2818000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3624 diff_2632000_2818000# diff_2632000_2818000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3625 diff_95000_5192000# diff_2911000_2818000# diff_2911000_2818000# GND efet w=14000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3626 diff_3050000_2818000# diff_3050000_2818000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3627 diff_2602000_2818000# diff_72000_4515000# diff_2581000_2777000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=9.44e+08 ps=154000 
M3628 diff_2632000_2818000# diff_72000_4515000# diff_2632000_2777000# GND efet w=20000 l=13000
+ ad=0 pd=0 as=9.39e+08 ps=154000 
M3629 diff_2678000_3055000# diff_72000_4515000# diff_2684000_2777000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=9.34e+08 ps=154000 
M3630 diff_2735000_2818000# diff_72000_4515000# diff_2735000_2777000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=9.34e+08 ps=154000 
M3631 diff_3014000_2818000# diff_169000_4545000# diff_83000_3098000# GND efet w=64000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3632 diff_3532000_3485000# diff_3532000_3485000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3633 diff_3551000_3277000# diff_94000_3551000# diff_83000_3098000# GND efet w=62000 l=7000
+ ad=-4.84967e+08 pd=798000 as=0 ps=0 
M3634 diff_83000_3098000# diff_3702000_3518000# diff_3551000_3277000# GND efet w=78500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3635 diff_3551000_3277000# diff_3551000_3277000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3636 diff_3551000_3277000# diff_68000_5288000# diff_3517000_3179000# GND efet w=13000 l=14000
+ ad=0 pd=0 as=2.81e+08 ps=96000 
M3637 diff_3014000_2818000# diff_3014000_2818000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3638 diff_3355000_3022000# diff_597000_3013000# diff_2838000_2818000# GND efet w=130000 l=8000
+ ad=1.274e+09 pd=278000 as=-1.39697e+09 ps=600000 
M3639 diff_83000_3098000# diff_3365000_3033000# diff_3355000_3022000# GND efet w=129500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3640 diff_83000_3098000# diff_1604000_3123000# diff_3365000_3033000# GND efet w=77500 l=8500
+ ad=0 pd=0 as=2.012e+09 ps=378000 
M3641 diff_2838000_2818000# diff_2838000_2818000# diff_95000_5192000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M3642 diff_3365000_3033000# diff_3365000_3033000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3643 diff_2808000_2818000# diff_72000_4515000# diff_2788000_2777000# GND efet w=20000 l=13000
+ ad=0 pd=0 as=9.39e+08 ps=154000 
M3644 diff_2838000_2818000# diff_72000_4515000# diff_2838000_2777000# GND efet w=20000 l=13000
+ ad=0 pd=0 as=9.39e+08 ps=154000 
M3645 diff_2911000_2818000# diff_72000_4515000# diff_2891000_2777000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=9.2e+08 ps=152000 
M3646 diff_2941000_2818000# diff_72000_4515000# diff_2941000_2777000# GND efet w=20000 l=13000
+ ad=0 pd=0 as=9.48e+08 ps=154000 
M3647 diff_3014000_2818000# diff_72000_4515000# diff_2994000_2777000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=9.11e+08 ps=152000 
M3648 diff_3050000_2818000# diff_72000_4515000# diff_3047000_2783000# GND efet w=20000 l=13000
+ ad=0 pd=0 as=9.7e+08 ps=180000 
M3649 diff_2838000_2818000# diff_72000_4515000# diff_3115000_2777000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=9.43e+08 ps=154000 
M3650 diff_3188000_2818000# diff_72000_4515000# diff_3168000_2777000# GND efet w=19000 l=13000
+ ad=-1.31967e+08 pd=822000 as=9.11e+08 ps=152000 
M3651 diff_95000_5192000# diff_1438000_786000# diff_1438000_786000# GND efet w=25000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3652 diff_2448000_2717000# diff_2448000_2717000# diff_95000_5192000# GND efet w=18000 l=9000
+ ad=-2.20967e+08 pd=894000 as=0 ps=0 
M3653 diff_1438000_786000# diff_2448000_2717000# diff_83000_3098000# GND efet w=447000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3654 diff_83000_3098000# diff_1438000_786000# diff_1237000_1921000# GND efet w=214000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3655 diff_83000_3098000# diff_72000_4515000# diff_2448000_2717000# GND efet w=217500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3656 diff_1850000_2290000# diff_1837000_1364000# diff_817000_2342000# GND efet w=102000 l=10000
+ ad=-1.92967e+08 pd=730000 as=0 ps=0 
M3657 diff_1932000_2308000# diff_95000_5192000# diff_1850000_2290000# GND efet w=13000 l=79000
+ ad=8.94e+08 pd=206000 as=0 ps=0 
M3658 diff_95000_5192000# diff_95000_5192000# diff_1850000_2290000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3659 diff_95000_5192000# diff_95000_5192000# diff_1881000_2203000# GND efet w=13000 l=32000
+ ad=0 pd=0 as=1.107e+09 ps=212000 
M3660 diff_1850000_2290000# diff_1858000_1019000# diff_1399000_598000# GND efet w=105500 l=10500
+ ad=0 pd=0 as=3.04065e+08 ps=1.764e+06 
M3661 diff_95000_5192000# diff_1997000_2222000# diff_1997000_2222000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=-1.30597e+09 ps=670000 
M3662 diff_1997000_2222000# diff_1547000_932000# diff_1932000_2308000# GND efet w=20000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3663 diff_2102000_2360000# diff_1438000_786000# diff_2050000_2211000# GND efet w=22000 l=13000
+ ad=1.54e+08 pd=58000 as=3.68e+08 ps=100000 
M3664 diff_2122000_2360000# diff_72000_4515000# diff_2102000_2360000# GND efet w=22000 l=12500
+ ad=-1.30297e+09 pd=438000 as=0 ps=0 
M3665 diff_1399000_598000# diff_1487000_841000# diff_1997000_2222000# GND efet w=120000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3666 diff_83000_3098000# diff_1881000_2203000# diff_1850000_2290000# GND efet w=198500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3667 diff_1881000_2203000# diff_1932000_2308000# diff_83000_3098000# GND efet w=61000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3668 diff_1850000_2072000# diff_1858000_1019000# diff_1757000_739000# GND efet w=106000 l=10000
+ ad=-1.96967e+08 pd=726000 as=2.28065e+08 ps=1.764e+06 
M3669 diff_83000_3098000# diff_1881000_2171000# diff_1850000_2072000# GND efet w=197500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3670 diff_1850000_2072000# diff_1837000_1364000# diff_817000_2040000# GND efet w=103000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3671 diff_1881000_2171000# diff_1932000_2082000# diff_83000_3098000# GND efet w=62000 l=8000
+ ad=1.147e+09 pd=208000 as=0 ps=0 
M3672 diff_1850000_1913000# diff_1837000_1364000# diff_817000_1965000# GND efet w=102000 l=10000
+ ad=-6.89673e+07 pd=730000 as=0 ps=0 
M3673 diff_1997000_2222000# diff_2050000_2211000# diff_83000_3098000# GND efet w=185500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3674 diff_1757000_739000# diff_1487000_841000# diff_1997000_2116000# GND efet w=116500 l=10500
+ ad=0 pd=0 as=-1.20997e+09 ps=668000 
M3675 diff_1997000_2116000# diff_2050000_2147000# diff_83000_3098000# GND efet w=183500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3676 diff_1997000_2116000# diff_1547000_932000# diff_1932000_2082000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=8.32e+08 ps=202000 
M3677 diff_1850000_2072000# diff_95000_5192000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3678 diff_1932000_2082000# diff_95000_5192000# diff_1850000_2072000# GND efet w=12500 l=79500
+ ad=0 pd=0 as=0 ps=0 
M3679 diff_1881000_2171000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=32000
+ ad=0 pd=0 as=0 ps=0 
M3680 diff_1932000_1931000# diff_95000_5192000# diff_1850000_1913000# GND efet w=13000 l=79000
+ ad=8.73e+08 pd=204000 as=0 ps=0 
M3681 diff_95000_5192000# diff_95000_5192000# diff_1850000_1913000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3682 diff_95000_5192000# diff_95000_5192000# diff_1881000_1826000# GND efet w=13000 l=32000
+ ad=0 pd=0 as=1.112e+09 ps=212000 
M3683 diff_1850000_1913000# diff_1858000_1019000# diff_1774000_760000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=3.99065e+08 ps=1.766e+06 
M3684 diff_1997000_2116000# diff_1997000_2116000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3685 diff_95000_5192000# diff_1997000_1845000# diff_1997000_1845000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=-1.30597e+09 ps=668000 
M3686 diff_1997000_1845000# diff_1547000_932000# diff_1932000_1931000# GND efet w=19000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3687 diff_95000_5192000# diff_2122000_2360000# diff_2122000_2360000# GND efet w=11000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3688 diff_2122000_2360000# diff_2130000_2350000# diff_2137000_2334000# GND efet w=66000 l=7000
+ ad=0 pd=0 as=1.856e+09 ps=382000 
M3689 diff_95000_5192000# diff_2184000_2248000# diff_2184000_2248000# GND efet w=12000 l=19000
+ ad=0 pd=0 as=1.618e+09 ps=344000 
M3690 diff_2534000_2492000# diff_2529000_2777000# diff_83000_3098000# GND efet w=244000 l=8000
+ ad=3.85033e+08 pd=874000 as=0 ps=0 
M3691 diff_95000_5192000# diff_2534000_2492000# diff_2534000_2492000# GND efet w=17000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3692 diff_2583000_2725000# diff_2583000_2725000# diff_95000_5192000# GND efet w=17000 l=8000
+ ad=3.02033e+08 pd=870000 as=0 ps=0 
M3693 diff_83000_3098000# diff_72000_4515000# diff_2534000_2492000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3694 diff_2583000_2725000# diff_72000_4515000# diff_83000_3098000# GND efet w=204000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3695 diff_83000_3098000# diff_2581000_2777000# diff_2583000_2725000# GND efet w=244000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3696 diff_2638000_2492000# diff_2632000_2777000# diff_83000_3098000# GND efet w=244500 l=8500
+ ad=2.77033e+08 pd=870000 as=0 ps=0 
M3697 diff_95000_5192000# diff_2638000_2492000# diff_2638000_2492000# GND efet w=17000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M3698 diff_2641000_934000# diff_2641000_934000# diff_95000_5192000# GND efet w=17000 l=8000
+ ad=1.63033e+08 pd=870000 as=0 ps=0 
M3699 diff_83000_3098000# diff_72000_4515000# diff_2638000_2492000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3700 diff_2641000_934000# diff_72000_4515000# diff_83000_3098000# GND efet w=203000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3701 diff_83000_3098000# diff_2684000_2777000# diff_2641000_934000# GND efet w=244500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3702 diff_2713000_822000# diff_2735000_2777000# diff_83000_3098000# GND efet w=244500 l=8500
+ ad=2.19033e+08 pd=866000 as=0 ps=0 
M3703 diff_95000_5192000# diff_2713000_822000# diff_2713000_822000# GND efet w=17000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3704 diff_2775000_765000# diff_2775000_765000# diff_95000_5192000# GND efet w=17000 l=8000
+ ad=1.14203e+09 pd=966000 as=0 ps=0 
M3705 diff_83000_3098000# diff_72000_4515000# diff_2713000_822000# GND efet w=203000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3706 diff_2775000_765000# diff_72000_4515000# diff_83000_3098000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3707 diff_83000_3098000# diff_2788000_2777000# diff_2775000_765000# GND efet w=244000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3708 diff_2843000_1950000# diff_2838000_2777000# diff_83000_3098000# GND efet w=244500 l=8500
+ ad=4.22033e+08 pd=872000 as=0 ps=0 
M3709 diff_95000_5192000# diff_2843000_1950000# diff_2843000_1950000# GND efet w=17000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3710 diff_2893000_2725000# diff_2893000_2725000# diff_95000_5192000# GND efet w=17000 l=8000
+ ad=5.81033e+08 pd=882000 as=0 ps=0 
M3711 diff_83000_3098000# diff_72000_4515000# diff_2843000_1950000# GND efet w=203000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3712 diff_2893000_2725000# diff_72000_4515000# diff_83000_3098000# GND efet w=203000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3713 diff_83000_3098000# diff_2891000_2777000# diff_2893000_2725000# GND efet w=245000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3714 diff_2939000_824000# diff_2941000_2777000# diff_83000_3098000# GND efet w=245000 l=8000
+ ad=1.97033e+08 pd=852000 as=0 ps=0 
M3715 diff_95000_5192000# diff_2939000_824000# diff_2939000_824000# GND efet w=17000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3716 diff_2996000_2725000# diff_2996000_2725000# diff_95000_5192000# GND efet w=17000 l=7000
+ ad=4.36033e+08 pd=880000 as=0 ps=0 
M3717 diff_83000_3098000# diff_72000_4515000# diff_2939000_824000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3718 diff_2996000_2725000# diff_72000_4515000# diff_83000_3098000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3719 diff_83000_3098000# diff_2994000_2777000# diff_2996000_2725000# GND efet w=244500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3720 diff_95000_5192000# diff_3043000_2723000# diff_3043000_2723000# GND efet w=13000 l=11000
+ ad=0 pd=0 as=-2.96967e+08 ps=690000 
M3721 diff_3120000_2492000# diff_3115000_2777000# diff_83000_3098000# GND efet w=244000 l=8000
+ ad=2.50033e+08 pd=880000 as=0 ps=0 
M3722 diff_95000_5192000# diff_3120000_2492000# diff_3120000_2492000# GND efet w=18000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3723 diff_3171000_2725000# diff_3171000_2725000# diff_95000_5192000# GND efet w=18000 l=8000
+ ad=5.16033e+08 pd=856000 as=0 ps=0 
M3724 diff_83000_3098000# diff_72000_4515000# diff_3120000_2492000# GND efet w=202500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3725 diff_95000_5192000# diff_2281000_2195000# diff_2281000_2195000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=1.317e+09 ps=312000 
M3726 diff_95000_5192000# diff_1237000_1921000# diff_2127000_2299000# GND efet w=13000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3727 diff_2137000_2334000# diff_2127000_2299000# diff_83000_3098000# GND efet w=125500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3728 diff_2122000_2360000# diff_2130000_2350000# diff_2137000_2334000# GND efet w=72500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3729 diff_83000_3098000# diff_2184000_2248000# diff_2122000_2360000# GND efet w=57000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3730 diff_2184000_2248000# diff_2130000_2350000# diff_83000_3098000# GND efet w=64000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3731 diff_83000_3098000# diff_2127000_2299000# diff_2184000_2248000# GND efet w=72000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3732 diff_2137000_2050000# diff_2127000_2082000# diff_83000_3098000# GND efet w=129000 l=8000
+ ad=1.932e+09 pd=382000 as=0 ps=0 
M3733 diff_2122000_2014000# diff_2130000_2043000# diff_2137000_2050000# GND efet w=76000 l=8000
+ ad=-1.18897e+09 pd=466000 as=0 ps=0 
M3734 diff_2137000_2050000# diff_2130000_2043000# diff_2122000_2014000# GND efet w=62500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3735 diff_83000_3098000# diff_2184000_2056000# diff_2122000_2014000# GND efet w=56000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3736 diff_2184000_2056000# diff_2130000_2043000# diff_83000_3098000# GND efet w=64000 l=8000
+ ad=1.615e+09 pd=340000 as=0 ps=0 
M3737 diff_83000_3098000# diff_2127000_2082000# diff_2184000_2056000# GND efet w=72000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3738 diff_2184000_2056000# diff_2184000_2056000# diff_95000_5192000# GND efet w=12000 l=18000
+ ad=0 pd=0 as=0 ps=0 
M3739 diff_2102000_2014000# diff_1438000_786000# diff_2050000_2147000# GND efet w=21000 l=14000
+ ad=1.47e+08 pd=56000 as=3.56e+08 ps=90000 
M3740 diff_2122000_2014000# diff_72000_4515000# diff_2102000_2014000# GND efet w=21000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M3741 diff_95000_5192000# diff_2122000_2014000# diff_2122000_2014000# GND efet w=11000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3742 diff_95000_5192000# diff_2320000_2261000# diff_2320000_2261000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=-1.92397e+09 ps=430000 
M3743 diff_95000_5192000# diff_2130000_2350000# diff_2130000_2350000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=1.368e+09 ps=312000 
M3744 diff_2320000_2261000# diff_1094000_1020000# diff_2406000_2323000# GND efet w=150500 l=8500
+ ad=0 pd=0 as=1.535e+09 ps=306000 
M3745 diff_2127000_2299000# diff_2281000_2195000# diff_2127000_2082000# GND efet w=117500 l=9500
+ ad=0 pd=0 as=-1.49997e+09 ps=594000 
M3746 diff_83000_3098000# diff_2320000_2261000# diff_2281000_2195000# GND efet w=55500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3747 diff_2304000_1746000# diff_2320000_2261000# diff_83000_3098000# GND efet w=152000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3748 diff_2406000_2323000# diff_2130000_2350000# diff_83000_3098000# GND efet w=120000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3749 diff_2127000_1922000# diff_2281000_2086000# diff_2127000_2082000# GND efet w=137000 l=9000
+ ad=-7.44967e+08 pd=662000 as=0 ps=0 
M3750 diff_2304000_1746000# diff_2320000_2130000# diff_83000_3098000# GND efet w=154500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3751 diff_83000_3098000# diff_2320000_2130000# diff_2281000_2086000# GND efet w=62000 l=8000
+ ad=0 pd=0 as=1.247e+09 ps=306000 
M3752 diff_2102000_1984000# diff_1438000_786000# diff_2050000_1834000# GND efet w=20000 l=14000
+ ad=1.4e+08 pd=54000 as=3.17e+08 ps=92000 
M3753 diff_2122000_1984000# diff_72000_4515000# diff_2102000_1984000# GND efet w=20000 l=13000
+ ad=-1.33597e+09 pd=438000 as=0 ps=0 
M3754 diff_1774000_760000# diff_1487000_841000# diff_1997000_1845000# GND efet w=120000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3755 diff_83000_3098000# diff_1881000_1826000# diff_1850000_1913000# GND efet w=198500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3756 diff_1881000_1826000# diff_1932000_1931000# diff_83000_3098000# GND efet w=61000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3757 diff_1851000_1695000# diff_1858000_1019000# diff_1791000_798000# GND efet w=106000 l=10000
+ ad=-2.61967e+08 pd=722000 as=3.52065e+08 ps=1.768e+06 
M3758 diff_83000_3098000# diff_1881000_1794000# diff_1851000_1695000# GND efet w=198500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3759 diff_1851000_1695000# diff_1837000_1364000# diff_817000_1663000# GND efet w=101000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3760 diff_1881000_1794000# diff_1932000_1705000# diff_83000_3098000# GND efet w=62000 l=8000
+ ad=1.146e+09 pd=208000 as=0 ps=0 
M3761 diff_1997000_1845000# diff_2050000_1834000# diff_83000_3098000# GND efet w=184500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3762 diff_1997000_1739000# diff_2050000_1770000# diff_83000_3098000# GND efet w=185500 l=8500
+ ad=-1.21097e+09 pd=668000 as=0 ps=0 
M3763 diff_1791000_798000# diff_1487000_841000# diff_1997000_1739000# GND efet w=117000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3764 diff_1850000_1535000# diff_1837000_1364000# diff_817000_1588000# GND efet w=103000 l=10000
+ ad=-4.99673e+07 pd=732000 as=0 ps=0 
M3765 diff_1997000_1739000# diff_1547000_932000# diff_1932000_1705000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=8.15e+08 ps=198000 
M3766 diff_1851000_1695000# diff_95000_5192000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3767 diff_1932000_1705000# diff_95000_5192000# diff_1851000_1695000# GND efet w=12500 l=80500
+ ad=0 pd=0 as=0 ps=0 
M3768 diff_1881000_1794000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=32000
+ ad=0 pd=0 as=0 ps=0 
M3769 diff_1932000_1554000# diff_95000_5192000# diff_1850000_1535000# GND efet w=13000 l=78000
+ ad=8.52e+08 pd=202000 as=0 ps=0 
M3770 diff_95000_5192000# diff_95000_5192000# diff_1850000_1535000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3771 diff_95000_5192000# diff_95000_5192000# diff_1881000_1450000# GND efet w=13000 l=32000
+ ad=0 pd=0 as=1.062e+09 ps=210000 
M3772 diff_1850000_1535000# diff_1858000_1019000# diff_1851000_1456000# GND efet w=105500 l=10500
+ ad=0 pd=0 as=5.06065e+08 ps=1.78e+06 
M3773 diff_1997000_1739000# diff_1997000_1739000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3774 diff_95000_5192000# diff_1997000_1468000# diff_1997000_1468000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=-1.29797e+09 ps=668000 
M3775 diff_1997000_1468000# diff_1547000_932000# diff_1932000_1554000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3776 diff_95000_5192000# diff_2122000_1984000# diff_2122000_1984000# GND efet w=10000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3777 diff_2127000_2082000# diff_1237000_1921000# diff_95000_5192000# GND efet w=12000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3778 diff_2460000_2210000# diff_1037000_877000# diff_2320000_2261000# GND efet w=151000 l=8000
+ ad=1.672e+09 pd=328000 as=0 ps=0 
M3779 diff_817000_2342000# diff_1438000_786000# diff_95000_5192000# GND efet w=87500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3780 diff_83000_3098000# diff_2471000_2205000# diff_2460000_2210000# GND efet w=123500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3781 diff_2130000_2350000# diff_2471000_2205000# diff_83000_3098000# GND efet w=58000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M3782 diff_95000_5192000# diff_2532000_2233000# diff_2532000_2233000# GND efet w=11000 l=15000
+ ad=0 pd=0 as=1.573e+09 ps=342000 
M3783 diff_95000_5192000# diff_95000_5192000# diff_2674000_2207000# GND efet w=11000 l=31000
+ ad=0 pd=0 as=9.18e+08 ps=196000 
M3784 diff_2683000_2215000# diff_95000_5192000# diff_2651000_2299000# GND efet w=12000 l=74000
+ ad=-1.66967e+08 pd=732000 as=5.26e+08 ps=186000 
M3785 diff_95000_5192000# diff_95000_5192000# diff_2683000_2215000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3786 diff_2651000_2299000# diff_2641000_934000# diff_817000_2342000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3787 diff_83000_3098000# diff_1399000_598000# diff_2532000_2233000# GND efet w=84000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3788 diff_2532000_2233000# diff_2448000_2717000# diff_2471000_2205000# GND efet w=20000 l=13000
+ ad=0 pd=0 as=3.31e+08 ps=92000 
M3789 diff_2281000_2086000# diff_2281000_2086000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3790 diff_2127000_1922000# diff_1237000_1921000# diff_95000_5192000# GND efet w=10000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3791 diff_2122000_1984000# diff_2130000_1972000# diff_2137000_1957000# GND efet w=65500 l=7500
+ ad=0 pd=0 as=1.843e+09 ps=380000 
M3792 diff_95000_5192000# diff_2184000_1871000# diff_2184000_1871000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=1.631e+09 ps=342000 
M3793 diff_2137000_1957000# diff_2127000_1922000# diff_83000_3098000# GND efet w=125500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3794 diff_2122000_1984000# diff_2130000_1972000# diff_2137000_1957000# GND efet w=73000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3795 diff_83000_3098000# diff_2184000_1871000# diff_2122000_1984000# GND efet w=56000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3796 diff_2184000_1871000# diff_2130000_1972000# diff_83000_3098000# GND efet w=64000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3797 diff_83000_3098000# diff_2127000_1922000# diff_2184000_1871000# GND efet w=72000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3798 diff_2137000_1673000# diff_2127000_1705000# diff_83000_3098000# GND efet w=129000 l=8000
+ ad=1.936e+09 pd=382000 as=0 ps=0 
M3799 diff_2122000_1637000# diff_2130000_1666000# diff_2137000_1673000# GND efet w=75500 l=8500
+ ad=-1.20297e+09 pd=464000 as=0 ps=0 
M3800 diff_2137000_1673000# diff_2130000_1666000# diff_2122000_1637000# GND efet w=62500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3801 diff_83000_3098000# diff_2184000_1679000# diff_2122000_1637000# GND efet w=57000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3802 diff_2184000_1679000# diff_2130000_1666000# diff_83000_3098000# GND efet w=64000 l=8000
+ ad=1.628e+09 pd=338000 as=0 ps=0 
M3803 diff_83000_3098000# diff_2127000_1705000# diff_2184000_1679000# GND efet w=71000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3804 diff_2127000_1922000# diff_2281000_1866000# diff_2127000_1705000# GND efet w=117000 l=10000
+ ad=0 pd=0 as=-8.13967e+08 ps=602000 
M3805 diff_95000_5192000# diff_2281000_1866000# diff_2281000_1866000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=1.432e+09 ps=318000 
M3806 diff_2407000_2069000# diff_2130000_2043000# diff_83000_3098000# GND efet w=115500 l=8500
+ ad=1.514e+09 pd=296000 as=0 ps=0 
M3807 diff_2320000_2130000# diff_1094000_1020000# diff_2407000_2069000# GND efet w=146500 l=8500
+ ad=-1.92197e+09 pd=418000 as=0 ps=0 
M3808 diff_2460000_2101000# diff_1037000_877000# diff_2320000_2130000# GND efet w=150000 l=8000
+ ad=1.668e+09 pd=326000 as=0 ps=0 
M3809 diff_83000_3098000# diff_2471000_2112000# diff_2460000_2101000# GND efet w=123500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3810 diff_95000_5192000# diff_1438000_786000# diff_1399000_598000# GND efet w=85500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3811 diff_848000_2342000# diff_1438000_786000# diff_95000_5192000# GND efet w=71000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3812 diff_2674000_2207000# diff_2651000_2299000# diff_83000_3098000# GND efet w=63000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3813 diff_95000_5192000# diff_95000_5192000# diff_2829000_2242000# GND efet w=11000 l=22000
+ ad=0 pd=0 as=2.0327e+06 ps=736000 
M3814 diff_2915000_2318000# diff_95000_5192000# diff_2829000_2242000# GND efet w=12000 l=72000
+ ad=1.236e+09 pd=312000 as=0 ps=0 
M3815 diff_95000_5192000# diff_95000_5192000# diff_2876000_2205000# GND efet w=12000 l=30000
+ ad=0 pd=0 as=8.6e+08 ps=188000 
M3816 diff_3079000_2441000# diff_1237000_1921000# diff_3043000_2723000# GND efet w=244000 l=8000
+ ad=-2.02197e+09 pd=516000 as=0 ps=0 
M3817 diff_83000_3098000# diff_3047000_2783000# diff_3079000_2441000# GND efet w=248500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3818 diff_3171000_2725000# diff_72000_4515000# diff_83000_3098000# GND efet w=202000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3819 diff_83000_3098000# diff_3168000_2777000# diff_3171000_2725000# GND efet w=245500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3820 diff_95000_5192000# diff_3256000_1459000# diff_3256000_1459000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=-8.30967e+08 ps=642000 
M3821 diff_95000_5192000# diff_3283000_1426000# diff_3283000_1426000# GND efet w=13000 l=16000
+ ad=0 pd=0 as=-1.72297e+09 ps=516000 
M3822 diff_3283000_1426000# diff_3283000_1426000# diff_3283000_1426000# GND efet w=1000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3823 diff_3256000_1459000# diff_3254000_2509000# diff_83000_3098000# GND efet w=102000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3824 diff_3487000_3126000# diff_2849000_2986000# diff_83000_3098000# GND efet w=129000 l=9000
+ ad=1.161e+09 pd=276000 as=0 ps=0 
M3825 diff_3433000_2818000# diff_531000_4622000# diff_3487000_3126000# GND efet w=129000 l=9000
+ ad=-1.17097e+09 pd=644000 as=0 ps=0 
M3826 diff_83000_3098000# diff_3517000_3179000# diff_3433000_2818000# GND efet w=75500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3827 diff_83000_3098000# diff_3517000_3070000# diff_3433000_2818000# GND efet w=64000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3828 diff_3188000_2818000# diff_3188000_2818000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3829 diff_3188000_2818000# diff_791000_4022000# diff_3791000_3500000# GND efet w=143500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3830 diff_83000_3098000# diff_2772000_3402000# diff_3188000_2818000# GND efet w=64000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3831 diff_4126000_4460000# diff_1001000_4394000# diff_4136000_4237000# GND efet w=139000 l=9000
+ ad=0 pd=0 as=2.038e+09 ps=410000 
M3832 diff_4125000_2818000# diff_791000_4022000# diff_4175000_4495000# GND efet w=130000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3833 diff_4247000_4333000# diff_4105000_4962000# diff_4125000_2818000# GND efet w=131000 l=9000
+ ad=1.179e+09 pd=280000 as=0 ps=0 
M3834 diff_83000_3098000# diff_946000_3261000# diff_4247000_4333000# GND efet w=131000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3835 diff_4382000_4593000# diff_4382000_4593000# diff_95000_5192000# GND efet w=12000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M3836 diff_83000_3098000# diff_4381000_4962000# diff_4467000_4516000# GND efet w=42000 l=8000
+ ad=0 pd=0 as=8.08e+08 ps=208000 
M3837 diff_4318000_4212000# diff_4319000_4839000# diff_83000_3098000# GND efet w=77000 l=9000
+ ad=-1.01593e+09 pd=1.636e+06 as=0 ps=0 
M3838 diff_4125000_2818000# diff_4125000_2818000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3839 diff_4467000_4516000# diff_4467000_4516000# diff_95000_5192000# GND efet w=13000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M3840 diff_83000_3098000# diff_4559000_4962000# diff_4647000_4721000# GND efet w=40000 l=9000
+ ad=0 pd=0 as=-2.07297e+09 ps=434000 
M3841 diff_4647000_4721000# diff_4587000_4962000# diff_83000_3098000# GND efet w=44000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3842 diff_4647000_4721000# diff_4647000_4721000# diff_95000_5192000# GND efet w=12000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M3843 diff_83000_3098000# diff_4617000_4962000# diff_4694000_4601000# GND efet w=44000 l=8000
+ ad=0 pd=0 as=1.656e+09 ps=412000 
M3844 diff_4694000_4601000# diff_4735000_4962000# diff_83000_3098000# GND efet w=49500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3845 diff_4318000_4212000# diff_4351000_4962000# diff_83000_3098000# GND efet w=65000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3846 diff_83000_3098000# diff_4382000_4593000# diff_4318000_4212000# GND efet w=61000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3847 diff_4469000_4450000# diff_4351000_4962000# diff_83000_3098000# GND efet w=42000 l=8000
+ ad=-3.23967e+08 pd=834000 as=0 ps=0 
M3848 diff_83000_3098000# diff_4467000_4516000# diff_4469000_4450000# GND efet w=41000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3849 diff_4524000_4435000# diff_1001000_4394000# diff_83000_3098000# GND efet w=89000 l=8000
+ ad=8.33e+08 pd=196000 as=0 ps=0 
M3850 diff_95000_5192000# diff_4136000_4237000# diff_4136000_4237000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3851 diff_4169000_3959000# diff_72000_4515000# diff_4143000_3861000# GND efet w=13000 l=12000
+ ad=2.9e+08 pd=100000 as=-1.15897e+09 ps=704000 
M3852 diff_83000_3098000# diff_3929000_4962000# diff_4214000_3933000# GND efet w=43000 l=9000
+ ad=0 pd=0 as=-1.14197e+09 ps=586000 
M3853 diff_4143000_3861000# diff_3666000_4069000# diff_83000_3098000# GND efet w=40000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3854 diff_83000_3098000# diff_4169000_3959000# diff_4163000_3767000# GND efet w=53500 l=8500
+ ad=0 pd=0 as=1.876e+09 ps=458000 
M3855 diff_3188000_2818000# diff_72000_4515000# diff_3621000_3188000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=5.04e+08 ps=140000 
M3856 diff_3604000_3007000# diff_68000_5288000# diff_3579000_3164000# GND efet w=12000 l=12000
+ ad=1.761e+09 pd=344000 as=2.32e+08 ps=96000 
M3857 diff_3517000_3070000# diff_3444000_3167000# diff_83000_3098000# GND efet w=64000 l=8000
+ ad=1.339e+09 pd=282000 as=0 ps=0 
M3858 diff_83000_3098000# diff_3579000_3164000# diff_3506000_2818000# GND efet w=80000 l=8000
+ ad=0 pd=0 as=-1.42697e+09 ps=554000 
M3859 diff_3433000_2818000# diff_3433000_2818000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3860 diff_3517000_3070000# diff_3517000_3070000# diff_95000_5192000# GND efet w=13000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M3861 diff_83000_3098000# diff_3621000_3188000# diff_3604000_3007000# GND efet w=64000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3862 diff_3604000_3007000# diff_3604000_3007000# diff_95000_5192000# GND efet w=13000 l=35000
+ ad=0 pd=0 as=0 ps=0 
M3863 diff_3819000_3049000# diff_3713000_4962000# diff_83000_3098000# GND efet w=80000 l=9000
+ ad=1.532e+09 pd=316000 as=0 ps=0 
M3864 diff_83000_3098000# diff_3666000_4069000# diff_3819000_3049000# GND efet w=78500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3865 diff_4218000_3818000# diff_4187000_3788000# diff_83000_3098000# GND efet w=85000 l=9000
+ ad=9.83e+08 pd=216000 as=0 ps=0 
M3866 diff_4214000_3933000# diff_4136000_4237000# diff_4218000_3818000# GND efet w=85000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3867 diff_4187000_3788000# diff_68000_5288000# diff_4163000_3767000# GND efet w=12000 l=12000
+ ad=2.31e+08 pd=78000 as=0 ps=0 
M3868 diff_4163000_3767000# diff_4163000_3767000# diff_95000_5192000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M3869 diff_4214000_3933000# diff_4214000_3933000# diff_95000_5192000# GND efet w=12000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M3870 diff_95000_5192000# diff_4143000_3861000# diff_4143000_3861000# GND efet w=11000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M3871 diff_4044000_3493000# diff_791000_4022000# diff_3609000_2818000# GND efet w=134000 l=9000
+ ad=1.281e+09 pd=286000 as=-1.62997e+09 ps=630000 
M3872 diff_83000_3098000# diff_3811000_4962000# diff_4044000_3493000# GND efet w=134500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3873 diff_3639000_2818000# diff_1197000_3119000# diff_83000_3098000# GND efet w=65000 l=8000
+ ad=-5.62967e+08 pd=598000 as=0 ps=0 
M3874 diff_83000_3098000# diff_1604000_3123000# diff_3536000_2818000# GND efet w=77500 l=7500
+ ad=0 pd=0 as=1.638e+09 ps=380000 
M3875 diff_3639000_2818000# diff_1604000_3123000# diff_83000_3098000# GND efet w=78000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3876 diff_83000_3098000# diff_531000_4622000# diff_3639000_2818000# GND efet w=64000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3877 diff_83000_3098000# diff_2931000_4557000# diff_3712000_2818000# GND efet w=79500 l=8500
+ ad=0 pd=0 as=1.872e+09 ps=430000 
M3878 diff_3819000_3049000# diff_3819000_3049000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3879 diff_3551000_3277000# diff_68000_5288000# diff_3917000_3246000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=3.73e+08 ps=110000 
M3880 diff_3867000_3072000# diff_72000_4515000# diff_3609000_2818000# GND efet w=11000 l=11000
+ ad=4.49e+08 pd=140000 as=0 ps=0 
M3881 diff_3742000_2818000# diff_3819000_3049000# diff_83000_3098000# GND efet w=80000 l=9000
+ ad=-1.62897e+09 pd=544000 as=0 ps=0 
M3882 diff_95000_5192000# diff_3506000_2818000# diff_3506000_2818000# GND efet w=13000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M3883 diff_3536000_2818000# diff_3536000_2818000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3884 diff_3639000_2818000# diff_3639000_2818000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3885 diff_3712000_2818000# diff_3712000_2818000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3886 diff_3742000_2818000# diff_3742000_2818000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3887 diff_3867000_2981000# diff_3867000_3072000# diff_83000_3098000# GND efet w=65000 l=8000
+ ad=1.792e+09 pd=386000 as=0 ps=0 
M3888 diff_3815000_2818000# diff_3917000_3246000# diff_83000_3098000# GND efet w=63000 l=8000
+ ad=-1.35197e+09 pd=586000 as=0 ps=0 
M3889 diff_4003000_3074000# diff_3700000_4748000# diff_83000_3098000# GND efet w=55000 l=9000
+ ad=1.191e+09 pd=278000 as=0 ps=0 
M3890 diff_83000_3098000# diff_3840000_4962000# diff_4003000_3074000# GND efet w=50000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M3891 diff_4028000_3054000# diff_3981000_4517000# diff_83000_3098000# GND efet w=42000 l=8000
+ ad=-9.03967e+08 pd=752000 as=0 ps=0 
M3892 diff_83000_3098000# diff_4423000_4318000# diff_4318000_4212000# GND efet w=63000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3893 diff_83000_3098000# diff_4423000_4318000# diff_4469000_4450000# GND efet w=42000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3894 diff_4527000_4142000# diff_4411000_4962000# diff_4524000_4435000# GND efet w=89500 l=8500
+ ad=1.911e+09 pd=428000 as=0 ps=0 
M3895 diff_4694000_4601000# diff_4694000_4601000# diff_95000_5192000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M3896 diff_4527000_4142000# diff_4527000_4142000# diff_95000_5192000# GND efet w=12000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M3897 diff_4318000_4212000# diff_4318000_4212000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3898 diff_4469000_4450000# diff_4469000_4450000# diff_95000_5192000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M3899 diff_4374000_4012000# diff_3408000_4288000# diff_4318000_4212000# GND efet w=130000 l=9000
+ ad=1.04e+09 pd=276000 as=0 ps=0 
M3900 diff_83000_3098000# diff_4165000_4929000# diff_4374000_4012000# GND efet w=130000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3901 diff_83000_3098000# diff_4824000_4962000# diff_4788000_4476000# GND efet w=52500 l=8500
+ ad=0 pd=0 as=-2.11197e+09 ps=478000 
M3902 diff_83000_3098000# diff_4843000_4668000# diff_4788000_4476000# GND efet w=41000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3903 diff_95000_5192000# diff_5220000_4035000# diff_5220000_4035000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=1.509e+09 ps=280000 
M3904 diff_5296000_4764000# diff_72000_4515000# diff_4902000_4754000# GND efet w=13000 l=12000
+ ad=3.08e+08 pd=72000 as=0 ps=0 
M3905 diff_6029000_4913000# diff_72000_4515000# diff_2351000_3074000# GND efet w=14000 l=12000
+ ad=2.46e+08 pd=94000 as=0 ps=0 
M3906 diff_5220000_4035000# diff_6029000_4913000# diff_83000_3098000# GND efet w=81500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3907 diff_6029000_4890000# diff_72000_4515000# diff_4318000_4212000# GND efet w=13000 l=12000
+ ad=3.17e+08 pd=102000 as=0 ps=0 
M3908 diff_83000_3098000# diff_6029000_4913000# diff_6078000_4885000# GND efet w=131000 l=8000
+ ad=0 pd=0 as=1.179e+09 ps=280000 
M3909 diff_6078000_4885000# diff_6029000_4890000# diff_5601000_3945000# GND efet w=131000 l=10000
+ ad=0 pd=0 as=9.40654e+07 ps=1.138e+06 
M3910 diff_6029000_4851000# diff_72000_4515000# diff_4469000_4450000# GND efet w=14000 l=12000
+ ad=2.64e+08 pd=94000 as=0 ps=0 
M3911 diff_5601000_3945000# diff_6029000_4851000# diff_6078000_4836000# GND efet w=131000 l=8000
+ ad=0 pd=0 as=1.179e+09 ps=280000 
M3912 diff_83000_3098000# diff_5488000_4745000# diff_5413000_4658000# GND efet w=51500 l=7500
+ ad=0 pd=0 as=-1.36897e+09 ps=634000 
M3913 diff_4318000_4212000# diff_72000_4515000# diff_5488000_4745000# GND efet w=14000 l=12000
+ ad=0 pd=0 as=2.54e+08 ps=84000 
M3914 diff_4469000_4450000# diff_72000_4515000# diff_5489000_4718000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=6.27e+08 ps=142000 
M3915 diff_6078000_4836000# diff_5220000_4035000# diff_83000_3098000# GND efet w=131000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3916 diff_83000_3098000# diff_5489000_4718000# diff_5413000_4658000# GND efet w=52500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3917 diff_83000_3098000# diff_5641000_4717000# diff_6078000_4787000# GND efet w=131000 l=9000
+ ad=0 pd=0 as=1.179e+09 ps=280000 
M3918 diff_5641000_4717000# diff_68000_5288000# diff_817000_2342000# GND efet w=13000 l=13000
+ ad=2.43e+08 pd=88000 as=0 ps=0 
M3919 diff_6078000_4787000# diff_4927000_3400000# diff_5601000_3945000# GND efet w=131000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3920 diff_5601000_3945000# diff_4265000_3070000# diff_6078000_4738000# GND efet w=131000 l=8000
+ ad=0 pd=0 as=1.31e+09 ps=282000 
M3921 diff_5991000_4719000# diff_72000_4515000# diff_4920000_4772000# GND efet w=13000 l=13000
+ ad=3.96e+08 pd=104000 as=0 ps=0 
M3922 diff_6078000_4738000# diff_5991000_4719000# diff_83000_3098000# GND efet w=131000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3923 diff_4920000_4669000# diff_72000_4515000# diff_3009000_4523000# GND efet w=12000 l=12000
+ ad=2.34e+08 pd=72000 as=0 ps=0 
M3924 diff_4927000_3400000# diff_4920000_4669000# diff_83000_3098000# GND efet w=163000 l=9000
+ ad=-1.98097e+09 pd=506000 as=0 ps=0 
M3925 diff_4788000_4476000# diff_4788000_4476000# diff_95000_5192000# GND efet w=12000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M3926 diff_95000_5192000# diff_4927000_3400000# diff_4927000_3400000# GND efet w=13000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M3927 diff_5413000_4658000# diff_5413000_4658000# diff_95000_5192000# GND efet w=11000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M3928 diff_83000_3098000# diff_4751000_4352000# diff_5127000_4637000# GND efet w=80000 l=9000
+ ad=0 pd=0 as=6.4e+08 ps=176000 
M3929 diff_5601000_3945000# diff_5337000_4602000# diff_83000_3098000# GND efet w=74500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3930 diff_5127000_4637000# diff_4694000_4601000# diff_5127000_4617000# GND efet w=80000 l=9000
+ ad=0 pd=0 as=1.934e+09 ps=356000 
M3931 diff_83000_3098000# diff_5476000_4643000# diff_5413000_4658000# GND efet w=47000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3932 diff_4920000_4772000# diff_72000_4515000# diff_5476000_4643000# GND efet w=14000 l=11000
+ ad=0 pd=0 as=2.3e+08 ps=74000 
M3933 diff_5413000_4658000# diff_5296000_4530000# diff_83000_3098000# GND efet w=43000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3934 diff_5413000_4658000# diff_4927000_3400000# diff_83000_3098000# GND efet w=45000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3935 diff_95000_5192000# diff_5601000_3945000# diff_5601000_3945000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3936 diff_95000_5192000# diff_4806000_4501000# diff_4806000_4501000# GND efet w=13000 l=37000
+ ad=0 pd=0 as=-1.12897e+09 ps=656000 
M3937 diff_95000_5192000# diff_5127000_4617000# diff_5127000_4617000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M3938 diff_5337000_4602000# diff_5337000_4602000# diff_95000_5192000# GND efet w=11000 l=37000
+ ad=-2.05497e+09 pd=472000 as=0 ps=0 
M3939 diff_5160000_4311000# diff_72000_4515000# diff_5127000_4617000# GND efet w=11000 l=11000
+ ad=3.45e+08 pd=88000 as=0 ps=0 
M3940 diff_5096000_4554000# diff_4694000_4601000# diff_83000_3098000# GND efet w=58000 l=9000
+ ad=1.759e+09 pd=326000 as=0 ps=0 
M3941 diff_5601000_3945000# diff_5413000_4658000# diff_6079000_4659000# GND efet w=130000 l=9000
+ ad=0 pd=0 as=1.17e+09 ps=278000 
M3942 diff_6079000_4659000# diff_6049000_4641000# diff_83000_3098000# GND efet w=130000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3943 diff_6049000_4641000# diff_72000_4515000# diff_3408000_4288000# GND efet w=11000 l=12000
+ ad=3.17e+08 pd=98000 as=-1.90597e+09 ps=510000 
M3944 diff_95000_5192000# diff_3408000_4288000# diff_3408000_4288000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M3945 diff_3408000_4288000# diff_5711000_4528000# diff_83000_3098000# GND efet w=116000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3946 diff_5096000_4554000# diff_5074000_4506000# diff_83000_3098000# GND efet w=42000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3947 diff_5229000_4554000# diff_72000_4515000# diff_5096000_4554000# GND efet w=12000 l=11000
+ ad=5.27e+08 pd=100000 as=0 ps=0 
M3948 diff_83000_3098000# diff_1001000_4394000# diff_5074000_4506000# GND efet w=64000 l=8000
+ ad=0 pd=0 as=1.394e+09 ps=260000 
M3949 diff_5337000_4569000# diff_5337000_4569000# diff_95000_5192000# GND efet w=10000 l=37000
+ ad=1.859e+09 pd=418000 as=0 ps=0 
M3950 diff_4751000_4352000# diff_4770000_4458000# diff_83000_3098000# GND efet w=70500 l=8500
+ ad=1.767e+09 pd=420000 as=0 ps=0 
M3951 diff_83000_3098000# diff_4423000_4318000# diff_4751000_4352000# GND efet w=79500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M3952 diff_4806000_4501000# diff_4788000_4476000# diff_83000_3098000# GND efet w=44500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3953 diff_83000_3098000# diff_4423000_4318000# diff_4806000_4501000# GND efet w=43000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3954 diff_5096000_4554000# diff_5096000_4554000# diff_95000_5192000# GND efet w=12000 l=35000
+ ad=0 pd=0 as=0 ps=0 
M3955 diff_5337000_4602000# diff_5457000_4544000# diff_83000_3098000# GND efet w=40000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3956 diff_5296000_4530000# diff_5296000_4530000# diff_95000_5192000# GND efet w=12000 l=36000
+ ad=1.326e+09 pd=212000 as=0 ps=0 
M3957 diff_4751000_4352000# diff_4751000_4352000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3958 diff_4374000_3894000# diff_4165000_4929000# diff_4358000_3758000# GND efet w=134500 l=8500
+ ad=1.206e+09 pd=286000 as=-1.83397e+09 ps=548000 
M3959 diff_83000_3098000# diff_791000_4022000# diff_4374000_3894000# GND efet w=134500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3960 diff_4419000_3822000# diff_791000_4022000# diff_83000_3098000# GND efet w=132500 l=8500
+ ad=1.191e+09 pd=282000 as=0 ps=0 
M3961 diff_4415000_3774000# diff_4428000_3813000# diff_4419000_3822000# GND efet w=132000 l=8000
+ ad=-1.10697e+09 pd=670000 as=0 ps=0 
M3962 diff_83000_3098000# diff_4193000_4962000# diff_4458000_3837000# GND efet w=140500 l=8500
+ ad=0 pd=0 as=-7.70967e+08 ps=752000 
M3963 diff_4458000_3837000# diff_4223000_4962000# diff_83000_3098000# GND efet w=146500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M3964 diff_4462000_3008000# diff_4516000_3837000# diff_4458000_3837000# GND efet w=131000 l=8000
+ ad=-9.87967e+08 pd=692000 as=0 ps=0 
M3965 diff_83000_3098000# diff_1197000_3119000# diff_4516000_3837000# GND efet w=71000 l=8000
+ ad=0 pd=0 as=-1.04797e+09 ps=682000 
M3966 diff_95000_5192000# diff_4358000_3758000# diff_4358000_3758000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3967 diff_4415000_3774000# diff_4415000_3774000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3968 diff_95000_5192000# diff_4462000_3008000# diff_4462000_3008000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3969 diff_4516000_3837000# diff_4516000_3837000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M3970 diff_83000_3098000# diff_4214000_3933000# diff_4022000_2818000# GND efet w=72500 l=7500
+ ad=0 pd=0 as=3.80327e+07 ps=822000 
M3971 diff_83000_3098000# diff_3929000_4962000# diff_4028000_3054000# GND efet w=43000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3972 diff_4028000_3054000# diff_2968000_4962000# diff_83000_3098000# GND efet w=43000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3973 diff_3609000_2818000# diff_3609000_2818000# diff_95000_5192000# GND efet w=11000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3974 diff_4022000_2818000# diff_2938000_3467000# diff_83000_3098000# GND efet w=63000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3975 diff_4304000_3505000# diff_4135000_4962000# diff_4022000_2818000# GND efet w=131000 l=8000
+ ad=1.179e+09 pd=280000 as=0 ps=0 
M3976 diff_83000_3098000# diff_530000_4372000# diff_4304000_3505000# GND efet w=131000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3977 diff_4003000_3074000# diff_4003000_3074000# diff_95000_5192000# GND efet w=13000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M3978 diff_4028000_3054000# diff_4028000_3054000# diff_95000_5192000# GND efet w=13000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M3979 diff_4022000_2818000# diff_4022000_2818000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3980 diff_3815000_2818000# diff_3904000_3049000# diff_83000_3098000# GND efet w=64000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3981 diff_83000_3098000# diff_1604000_3123000# diff_3815000_2818000# GND efet w=89000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3982 diff_3904000_3049000# diff_68000_5288000# diff_3867000_2981000# GND efet w=12000 l=11000
+ ad=2.74e+08 pd=78000 as=0 ps=0 
M3983 diff_3867000_2981000# diff_3867000_2981000# diff_95000_5192000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M3984 diff_3815000_2818000# diff_3815000_2818000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3985 diff_4297000_3178000# diff_4265000_3070000# diff_83000_3098000# GND efet w=69000 l=9000
+ ad=1.655e+09 pd=332000 as=0 ps=0 
M3986 diff_83000_3098000# diff_4003000_3074000# diff_3846000_2818000# GND efet w=67000 l=8000
+ ad=0 pd=0 as=-1.59997e+09 ps=596000 
M3987 diff_3949000_2818000# diff_4028000_3054000# diff_83000_3098000# GND efet w=79000 l=8000
+ ad=1.878e+09 pd=406000 as=0 ps=0 
M3988 diff_3949000_2818000# diff_3949000_2818000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3989 diff_3846000_2818000# diff_3846000_2818000# diff_95000_5192000# GND efet w=11000 l=19000
+ ad=0 pd=0 as=0 ps=0 
M3990 diff_3444000_3167000# diff_72000_4515000# diff_4095000_3085000# GND efet w=13000 l=11000
+ ad=0 pd=0 as=4.25e+08 ps=126000 
M3991 diff_4087000_3165000# diff_68000_5288000# diff_4068000_3124000# GND efet w=11000 l=12000
+ ad=4.85e+08 pd=122000 as=-2.09897e+09 ps=470000 
M3992 diff_83000_3098000# diff_4095000_3085000# diff_4068000_3124000# GND efet w=41000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3993 diff_4052000_2818000# diff_4087000_3165000# diff_83000_3098000# GND efet w=68000 l=8000
+ ad=-1.59497e+09 pd=554000 as=0 ps=0 
M3994 diff_4068000_3124000# diff_4068000_3124000# diff_95000_5192000# GND efet w=13000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M3995 diff_4154000_3010000# diff_2849000_2986000# diff_4052000_2818000# GND efet w=131000 l=8000
+ ad=1.51e+09 pd=320000 as=0 ps=0 
M3996 diff_83000_3098000# diff_530000_4372000# diff_4154000_3010000# GND efet w=150000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M3997 diff_4052000_2818000# diff_4052000_2818000# diff_95000_5192000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M3998 diff_4297000_3178000# diff_4297000_3178000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M3999 diff_83000_3098000# diff_1935000_3038000# diff_4225000_2934000# GND efet w=79000 l=8000
+ ad=0 pd=0 as=-1.71297e+09 ps=476000 
M4000 diff_4306000_3185000# diff_4297000_3178000# diff_83000_3098000# GND efet w=114000 l=9000
+ ad=1.026e+09 pd=246000 as=0 ps=0 
M4001 diff_4262000_2987000# diff_3408000_4288000# diff_4306000_3185000# GND efet w=114500 l=8500
+ ad=2.61033e+08 pd=834000 as=0 ps=0 
M4002 diff_83000_3098000# diff_1097000_3119000# diff_4495000_3314000# GND efet w=82000 l=9000
+ ad=0 pd=0 as=-9.87967e+08 ps=668000 
M4003 diff_83000_3098000# diff_1001000_4394000# diff_4423000_4318000# GND efet w=104000 l=8000
+ ad=0 pd=0 as=1.296e+09 ps=318000 
M4004 diff_95000_5192000# diff_5074000_4506000# diff_5074000_4506000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M4005 diff_5601000_3945000# diff_68000_5288000# diff_5711000_4528000# GND efet w=14000 l=12000
+ ad=0 pd=0 as=2.84e+08 ps=100000 
M4006 diff_5337000_4569000# diff_72000_4515000# diff_5457000_4544000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=2.4e+08 ps=82000 
M4007 diff_5337000_4569000# diff_5296000_4530000# diff_5391000_4498000# GND efet w=126000 l=9000
+ ad=0 pd=0 as=1.417e+09 ps=312000 
M4008 diff_5397000_4487000# diff_68000_5288000# diff_817000_2342000# GND efet w=19000 l=12000
+ ad=5e+08 pd=146000 as=0 ps=0 
M4009 diff_6153000_4534000# diff_5098000_4894000# diff_83000_3098000# GND efet w=42000 l=8000
+ ad=1.843e+09 pd=394000 as=0 ps=0 
M4010 diff_6153000_4534000# diff_5980000_4397000# diff_83000_3098000# GND efet w=45000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4011 diff_95000_5192000# diff_6153000_4534000# diff_6153000_4534000# GND efet w=12000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M4012 diff_4182000_2528000# diff_5740000_4460000# diff_83000_3098000# GND efet w=80000 l=9000
+ ad=1.718e+09 pd=352000 as=0 ps=0 
M4013 diff_83000_3098000# diff_5397000_4487000# diff_5391000_4498000# GND efet w=129500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4014 diff_5022000_4457000# diff_72000_4515000# diff_4995000_4438000# GND efet w=12000 l=11000
+ ad=4.49e+08 pd=152000 as=1.249e+09 ps=290000 
M4015 diff_5296000_4530000# diff_5022000_4457000# diff_83000_3098000# GND efet w=42000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4016 diff_83000_3098000# diff_4927000_3400000# diff_5258000_4376000# GND efet w=43000 l=9000
+ ad=0 pd=0 as=-1.66697e+09 ps=458000 
M4017 diff_4995000_4438000# diff_4984000_4430000# diff_83000_3098000# GND efet w=59000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4018 diff_95000_5192000# diff_4995000_4438000# diff_4995000_4438000# GND efet w=12000 l=35000
+ ad=0 pd=0 as=0 ps=0 
M4019 diff_5740000_4460000# diff_68000_5288000# diff_5389000_4406000# GND efet w=12000 l=11000
+ ad=2.79e+08 pd=88000 as=1.45307e+09 ps=1.87e+06 
M4020 diff_6223000_4302000# diff_5980000_4397000# diff_83000_3098000# GND efet w=41000 l=9000
+ ad=1.419e+09 pd=246000 as=0 ps=0 
M4021 diff_95000_5192000# diff_6223000_4302000# diff_6223000_4302000# GND efet w=12000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M4022 diff_83000_3098000# diff_4303000_2657000# diff_5949000_4452000# GND efet w=86000 l=9000
+ ad=0 pd=0 as=-1.90397e+09 ps=434000 
M4023 diff_83000_3098000# diff_4182000_2528000# diff_5949000_4452000# GND efet w=86000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4024 diff_5949000_4452000# diff_5826000_4381000# diff_5980000_4397000# GND efet w=88000 l=8000
+ ad=0 pd=0 as=1.748e+09 ps=330000 
M4025 diff_5056000_4359000# diff_68000_5288000# diff_4984000_4430000# GND efet w=14000 l=11000
+ ad=9.69e+08 pd=238000 as=2.66e+08 ps=74000 
M4026 diff_95000_5192000# diff_5056000_4359000# diff_5056000_4359000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M4027 diff_5389000_4406000# diff_5346000_4399000# diff_5389000_4389000# GND efet w=130000 l=7000
+ ad=0 pd=0 as=1.3e+09 ps=280000 
M4028 diff_5258000_4376000# diff_5258000_4376000# diff_95000_5192000# GND efet w=11000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M4029 diff_83000_3098000# diff_5561000_4418000# diff_5569000_4409000# GND efet w=129000 l=9000
+ ad=0 pd=0 as=1.161e+09 ps=276000 
M4030 diff_4182000_2528000# diff_72000_4515000# diff_5561000_4418000# GND efet w=13000 l=11000
+ ad=0 pd=0 as=2.2e+08 ps=80000 
M4031 diff_5569000_4409000# diff_5258000_4376000# diff_5389000_4406000# GND efet w=129000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4032 diff_83000_3098000# diff_5229000_4554000# diff_5258000_4376000# GND efet w=58000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4033 diff_5389000_4389000# diff_5229000_4554000# diff_83000_3098000# GND efet w=130000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4034 diff_95000_5192000# diff_5389000_4406000# diff_5389000_4406000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4035 diff_5056000_4359000# diff_4981000_4331000# diff_83000_3098000# GND efet w=51000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4036 diff_5169000_4319000# diff_5160000_4311000# diff_83000_3098000# GND efet w=45000 l=9000
+ ad=8.44e+08 pd=176000 as=0 ps=0 
M4037 diff_95000_5192000# diff_5169000_4319000# diff_5169000_4319000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M4038 diff_4981000_4331000# diff_72000_4515000# diff_4415000_3774000# GND efet w=13000 l=12000
+ ad=2.19e+08 pd=74000 as=0 ps=0 
M4039 diff_6187000_3965000# diff_6153000_4534000# diff_83000_3098000# GND efet w=48500 l=8500
+ ad=1.563e+09 pd=296000 as=0 ps=0 
M4040 diff_5980000_4397000# diff_5980000_4397000# diff_95000_5192000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M4041 diff_95000_5192000# diff_6187000_3965000# diff_6187000_3965000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M4042 diff_6187000_3965000# diff_5098000_4894000# diff_6146000_4381000# GND efet w=87000 l=8000
+ ad=0 pd=0 as=-1.91297e+09 ps=516000 
M4043 diff_83000_3098000# diff_5296000_4764000# diff_5603000_4344000# GND efet w=129000 l=8000
+ ad=0 pd=0 as=1.29e+09 ps=278000 
M4044 diff_5826000_4381000# diff_5826000_4381000# diff_95000_5192000# GND efet w=12000 l=36000
+ ad=9.11e+08 pd=240000 as=0 ps=0 
M4045 diff_6146000_4381000# diff_4241000_2640000# diff_83000_3098000# GND efet w=86000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4046 diff_6146000_4381000# diff_6223000_4302000# diff_83000_3098000# GND efet w=43000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4047 diff_6146000_4381000# diff_6223000_4302000# diff_83000_3098000# GND efet w=40000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M4048 diff_83000_3098000# diff_5296000_4764000# diff_5258000_4376000# GND efet w=42000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4049 diff_5603000_4344000# diff_4265000_3070000# diff_5389000_4406000# GND efet w=129000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4050 diff_4423000_4318000# diff_4423000_4318000# diff_95000_5192000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M4051 diff_5055000_4275000# diff_72000_4515000# diff_4697000_3226000# GND efet w=13000 l=11000
+ ad=2.56e+08 pd=88000 as=8.70327e+07 ps=954000 
M4052 diff_95000_5192000# diff_5091000_4257000# diff_5091000_4257000# GND efet w=11000 l=20000
+ ad=0 pd=0 as=1.587e+09 ps=332000 
M4053 diff_5258000_4376000# diff_5169000_4319000# diff_83000_3098000# GND efet w=42000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4054 diff_83000_3098000# diff_5055000_4275000# diff_5091000_4257000# GND efet w=64000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4055 diff_5389000_4406000# diff_4927000_3400000# diff_5603000_4298000# GND efet w=138500 l=9500
+ ad=0 pd=0 as=1.267e+09 ps=312000 
M4056 diff_5603000_4298000# diff_5376000_4257000# diff_83000_3098000# GND efet w=147000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4057 diff_5091000_4257000# diff_68000_5288000# diff_5164000_4226000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=4.72e+08 ps=132000 
M4058 diff_5376000_4257000# diff_68000_5288000# diff_817000_2040000# GND efet w=14000 l=12000
+ ad=4.18e+08 pd=112000 as=0 ps=0 
M4059 diff_5826000_4381000# diff_4182000_2528000# diff_6031000_4330000# GND efet w=86000 l=9000
+ ad=0 pd=0 as=8.6e+08 ps=192000 
M4060 diff_6031000_4330000# diff_4303000_2657000# diff_83000_3098000# GND efet w=86000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4061 diff_83000_3098000# diff_5068000_4962000# diff_5956000_4224000# GND efet w=43500 l=8500
+ ad=0 pd=0 as=7.69e+08 ps=162000 
M4062 diff_83000_3098000# diff_4241000_2640000# diff_6145000_4251000# GND efet w=42000 l=8000
+ ad=0 pd=0 as=-2.03197e+09 ps=434000 
M4063 diff_83000_3098000# diff_6223000_4302000# diff_6145000_4251000# GND efet w=41000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4064 diff_95000_5192000# diff_6145000_4251000# diff_6145000_4251000# GND efet w=13000 l=35000
+ ad=0 pd=0 as=0 ps=0 
M4065 diff_5575000_4252000# diff_5169000_4319000# diff_83000_3098000# GND efet w=134000 l=8000
+ ad=1.277e+09 pd=288000 as=0 ps=0 
M4066 diff_5575000_4252000# diff_5567000_4243000# diff_5389000_4406000# GND efet w=135000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4067 diff_95000_5192000# diff_4182000_2528000# diff_4182000_2528000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4068 diff_5956000_4224000# diff_5956000_4224000# diff_95000_5192000# GND efet w=11000 l=35000
+ ad=0 pd=0 as=0 ps=0 
M4069 diff_4715000_3889000# diff_791000_4022000# diff_4697000_3226000# GND efet w=143000 l=8000
+ ad=1.296e+09 pd=304000 as=0 ps=0 
M4070 diff_83000_3098000# diff_4499000_4962000# diff_4715000_3889000# GND efet w=143000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4071 diff_4527000_4142000# diff_72000_4515000# diff_5004000_4150000# GND efet w=12000 l=13000
+ ad=0 pd=0 as=2.07e+08 ps=72000 
M4072 diff_95000_5192000# diff_5028000_4156000# diff_5028000_4156000# GND efet w=12000 l=37000
+ ad=0 pd=0 as=1.267e+09 ps=272000 
M4073 diff_5028000_4156000# diff_5004000_4150000# diff_83000_3098000# GND efet w=42000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4074 diff_4778000_3875000# diff_4529000_4962000# diff_4762000_3821000# GND efet w=141000 l=8000
+ ad=1.378e+09 pd=300000 as=-1.88397e+09 ps=584000 
M4075 diff_83000_3098000# diff_4516000_3837000# diff_4778000_3875000# GND efet w=139500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4076 diff_5028000_4156000# diff_68000_5288000# diff_5019000_4116000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=4.15e+08 ps=116000 
M4077 diff_83000_3098000# diff_5019000_4116000# diff_5029000_4064000# GND efet w=41000 l=9000
+ ad=0 pd=0 as=1.319e+09 ps=278000 
M4078 diff_95000_5192000# diff_5114000_4071000# diff_5114000_4071000# GND efet w=12000 l=37000
+ ad=0 pd=0 as=1.717e+09 ps=386000 
M4079 diff_5567000_4243000# diff_72000_4515000# diff_5674000_4156000# GND efet w=11000 l=12000
+ ad=1.81e+08 pd=62000 as=-1.67197e+09 ps=544000 
M4080 diff_95000_5192000# diff_5674000_4156000# diff_5674000_4156000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M4081 diff_6158000_4260000# diff_6145000_4251000# diff_6158000_4243000# GND efet w=86000 l=9000
+ ad=-2.08497e+09 pd=386000 as=6.88e+08 ps=188000 
M4082 diff_95000_5192000# diff_6158000_4260000# diff_6158000_4260000# GND efet w=13000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M4083 diff_6158000_4243000# diff_5098000_4894000# diff_83000_3098000# GND efet w=86000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4084 diff_6158000_4260000# diff_6179000_4193000# diff_83000_3098000# GND efet w=42000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4085 diff_5674000_4156000# diff_5387000_800000# diff_83000_3098000# GND efet w=67000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4086 diff_5674000_4156000# diff_5164000_4226000# diff_83000_3098000# GND efet w=67000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4087 diff_95000_5192000# diff_5029000_4064000# diff_5029000_4064000# GND efet w=12000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M4088 diff_5055000_4064000# diff_72000_4515000# diff_5029000_4064000# GND efet w=12000 l=11000
+ ad=2.31e+08 pd=88000 as=0 ps=0 
M4089 diff_5114000_4071000# diff_5055000_4064000# diff_83000_3098000# GND efet w=52000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4090 diff_6179000_4193000# diff_5098000_4894000# diff_83000_3098000# GND efet w=50500 l=8500
+ ad=1.671e+09 pd=364000 as=0 ps=0 
M4091 diff_83000_3098000# diff_6223000_4302000# diff_6179000_4193000# GND efet w=43000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4092 diff_83000_3098000# diff_5918000_4120000# diff_2120000_4001000# GND efet w=79500 l=8500
+ ad=0 pd=0 as=-1.46967e+08 ps=710000 
M4093 diff_5356000_4071000# diff_5331000_4062000# diff_5356000_4053000# GND efet w=143500 l=8500
+ ad=-5.99346e+07 pd=1.698e+06 as=1.287e+09 ps=304000 
M4094 diff_5356000_4053000# diff_5220000_4035000# diff_5356000_4035000# GND efet w=143500 l=8500
+ ad=0 pd=0 as=1.24e+09 ps=304000 
M4095 diff_5356000_4035000# diff_5008000_3739000# diff_83000_3098000# GND efet w=142500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4096 diff_83000_3098000# diff_3408000_4288000# diff_5850000_3991000# GND efet w=42000 l=8000
+ ad=0 pd=0 as=2.059e+09 ps=448000 
M4097 diff_5612000_4010000# diff_5601000_3945000# diff_83000_3098000# GND efet w=118500 l=8500
+ ad=-9.12967e+08 pd=698000 as=0 ps=0 
M4098 diff_5850000_3991000# diff_5850000_3991000# diff_95000_5192000# GND efet w=12000 l=35000
+ ad=0 pd=0 as=0 ps=0 
M4099 diff_5612000_4010000# diff_5371000_3654000# diff_83000_3098000# GND efet w=132000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4100 diff_4716000_3243000# diff_4647000_4721000# diff_83000_3098000# GND efet w=73000 l=8000
+ ad=-1.73097e+09 pd=584000 as=0 ps=0 
M4101 diff_83000_3098000# diff_4428000_3813000# diff_4716000_3243000# GND efet w=71500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4102 diff_4697000_3226000# diff_4697000_3226000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4103 diff_4762000_3821000# diff_4762000_3821000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4104 diff_4716000_3243000# diff_4716000_3243000# diff_95000_5192000# GND efet w=13000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M4105 diff_83000_3098000# diff_1197000_3119000# diff_4716000_3243000# GND efet w=64000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4106 diff_83000_3098000# diff_3359000_4501000# diff_4814000_3335000# GND efet w=63000 l=9000
+ ad=0 pd=0 as=-1.73697e+09 ps=616000 
M4107 diff_83000_3098000# diff_1197000_3119000# diff_4814000_3335000# GND efet w=63000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M4108 diff_4751000_4352000# diff_72000_4515000# diff_5061000_3959000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=4.3e+08 ps=128000 
M4109 diff_83000_3098000# diff_5061000_3959000# diff_5274000_3953000# GND efet w=76500 l=8500
+ ad=0 pd=0 as=-1.02797e+09 ps=598000 
M4110 diff_5080000_3926000# diff_68000_5288000# diff_3551000_3277000# GND efet w=13000 l=12000
+ ad=4.74e+08 pd=148000 as=0 ps=0 
M4111 diff_5356000_4071000# diff_5331000_4062000# diff_5274000_3953000# GND efet w=161000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4112 diff_83000_3098000# diff_5080000_3926000# diff_5067000_3914000# GND efet w=45000 l=10000
+ ad=0 pd=0 as=1.115e+09 ps=230000 
M4113 diff_5274000_3953000# diff_5264000_3945000# diff_5263000_3933000# GND efet w=142500 l=7500
+ ad=0 pd=0 as=1.244e+09 ps=300000 
M4114 diff_5067000_3914000# diff_72000_4515000# diff_4975000_3889000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=3.58e+08 ps=110000 
M4115 diff_5263000_3933000# diff_5114000_4071000# diff_83000_3098000# GND efet w=122000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4116 diff_83000_3098000# diff_4975000_3889000# diff_4973000_3872000# GND efet w=42000 l=10000
+ ad=0 pd=0 as=1.246e+09 ps=274000 
M4117 diff_95000_5192000# diff_5067000_3914000# diff_5067000_3914000# GND efet w=12000 l=35000
+ ad=0 pd=0 as=0 ps=0 
M4118 diff_83000_3098000# diff_5114000_4071000# diff_5228000_3879000# GND efet w=41000 l=8000
+ ad=0 pd=0 as=-1.76967e+08 ps=794000 
M4119 diff_83000_3098000# diff_4927000_3400000# diff_5228000_3879000# GND efet w=49000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4120 diff_4973000_3872000# diff_68000_5288000# diff_4973000_3834000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=2.68e+08 ps=92000 
M4121 diff_95000_5192000# diff_4973000_3872000# diff_4973000_3872000# GND efet w=13000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M4122 diff_83000_3098000# diff_4973000_3834000# diff_4997000_3824000# GND efet w=44500 l=8500
+ ad=0 pd=0 as=1.174e+09 ps=254000 
M4123 diff_5346000_4399000# diff_5625000_3954000# diff_5612000_4010000# GND efet w=159000 l=8000
+ ad=-1.59797e+09 pd=436000 as=0 ps=0 
M4124 diff_95000_5192000# diff_5346000_4399000# diff_5346000_4399000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4125 diff_5850000_3991000# diff_3569000_3530000# diff_83000_3098000# GND efet w=42000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4126 diff_5850000_3991000# diff_4241000_2640000# diff_83000_3098000# GND efet w=41000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4127 diff_95000_5192000# diff_6179000_4193000# diff_6179000_4193000# GND efet w=11000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M4128 diff_5996000_3977000# diff_3569000_3530000# diff_83000_3098000# GND efet w=132000 l=8000
+ ad=1.90033e+08 pd=784000 as=0 ps=0 
M4129 diff_83000_3098000# diff_5850000_3991000# diff_5996000_3977000# GND efet w=131000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4130 diff_6196000_3985000# diff_6187000_3965000# diff_83000_3098000# GND efet w=87000 l=9000
+ ad=-1.39197e+09 pd=646000 as=0 ps=0 
M4131 diff_5918000_4120000# diff_5009000_4962000# diff_6196000_3985000# GND efet w=95500 l=8500
+ ad=-1.28197e+09 pd=566000 as=0 ps=0 
M4132 diff_95000_5192000# diff_5918000_4120000# diff_5918000_4120000# GND efet w=13000 l=33000
+ ad=0 pd=0 as=0 ps=0 
M4133 diff_5918000_4120000# diff_5956000_4224000# diff_83000_3098000# GND efet w=39000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4134 diff_83000_3098000# diff_5763000_4184000# diff_5918000_4120000# GND efet w=40000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4135 diff_6196000_3985000# diff_6158000_4260000# diff_5918000_4120000# GND efet w=113000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4136 diff_83000_3098000# diff_5696000_3194000# diff_6196000_3985000# GND efet w=93000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4137 diff_6196000_3985000# diff_5696000_3194000# diff_83000_3098000# GND efet w=32000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4138 diff_5996000_3977000# diff_5988000_3969000# diff_2120000_4001000# GND efet w=154500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4139 diff_5625000_3954000# diff_5601000_3945000# diff_5625000_3936000# GND efet w=130000 l=9000
+ ad=-2.07197e+09 pd=456000 as=1.17e+09 ps=278000 
M4140 diff_2120000_4001000# diff_2120000_4001000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M4141 diff_5625000_3936000# diff_5371000_3654000# diff_83000_3098000# GND efet w=130000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4142 diff_95000_5192000# diff_5625000_3954000# diff_5625000_3954000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4143 diff_2120000_4001000# diff_5983000_3917000# diff_83000_3098000# GND efet w=63000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4144 diff_2120000_4001000# diff_6076000_3942000# diff_83000_3098000# GND efet w=64000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4145 diff_5763000_4184000# diff_5763000_4184000# diff_95000_5192000# GND efet w=13000 l=37000
+ ad=9.8e+08 pd=218000 as=0 ps=0 
M4146 diff_4997000_3824000# diff_72000_4515000# diff_4994000_3787000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.53e+08 ps=102000 
M4147 diff_95000_5192000# diff_4997000_3824000# diff_4997000_3824000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M4148 diff_4627000_3380000# diff_1698000_2848000# diff_83000_3098000# GND efet w=211000 l=9000
+ ad=1.926e+09 pd=438000 as=0 ps=0 
M4149 diff_4478000_4817000# diff_3227000_4780000# diff_4627000_3380000# GND efet w=209500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4150 diff_83000_3098000# diff_4511000_3502000# diff_4495000_3314000# GND efet w=70000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4151 diff_4511000_3502000# diff_4319000_4839000# diff_83000_3098000# GND efet w=78000 l=9000
+ ad=1.458e+09 pd=316000 as=0 ps=0 
M4152 diff_83000_3098000# diff_4423000_4318000# diff_4511000_3502000# GND efet w=64000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4153 diff_4511000_3502000# diff_4511000_3502000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4154 diff_4495000_3314000# diff_4495000_3314000# diff_95000_5192000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4155 diff_4478000_4817000# diff_4478000_4817000# diff_95000_5192000# GND efet w=12000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M4156 diff_83000_3098000# diff_4265000_3070000# diff_4278000_3058000# GND efet w=107500 l=8500
+ ad=0 pd=0 as=1.236e+09 ps=274000 
M4157 diff_4262000_2987000# diff_4225000_2934000# diff_4278000_3058000# GND efet w=100000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4158 diff_4262000_2987000# diff_4262000_2987000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M4159 diff_95000_5192000# diff_4225000_2934000# diff_4225000_2934000# GND efet w=11000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M4160 diff_4363000_2478000# diff_4262000_2987000# diff_83000_3098000# GND efet w=178000 l=8000
+ ad=-1.11797e+09 pd=578000 as=0 ps=0 
M4161 diff_83000_3098000# diff_3569000_3530000# diff_4363000_2478000# GND efet w=169000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4162 diff_4435000_3015000# diff_4358000_3758000# diff_83000_3098000# GND efet w=196000 l=8000
+ ad=1.96e+09 pd=412000 as=0 ps=0 
M4163 diff_4453000_3015000# diff_4415000_3774000# diff_4435000_3015000# GND efet w=196000 l=8000
+ ad=1.764e+09 pd=410000 as=0 ps=0 
M4164 diff_4462000_2971000# diff_4462000_3008000# diff_4453000_3015000# GND efet w=196000 l=9000
+ ad=-2.81967e+08 pd=622000 as=0 ps=0 
M4165 diff_4591000_3170000# diff_4478000_4817000# diff_83000_3098000# GND efet w=64000 l=9000
+ ad=9.30327e+07 pd=704000 as=0 ps=0 
M4166 diff_83000_3098000# diff_4469000_4962000# diff_4591000_3170000# GND efet w=63000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4167 diff_4814000_3335000# diff_4814000_3335000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4168 diff_95000_5192000# diff_5008000_3739000# diff_5008000_3739000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=8.98e+08 ps=214000 
M4169 diff_5228000_3879000# diff_5228000_3879000# diff_95000_5192000# GND efet w=13000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M4170 diff_83000_3098000# diff_5061000_3959000# diff_5228000_3879000# GND efet w=59000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4171 diff_5008000_3739000# diff_4994000_3787000# diff_83000_3098000# GND efet w=52000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4172 diff_95000_5192000# diff_128000_4097000# diff_128000_4097000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4173 diff_128000_4097000# diff_5048000_3693000# diff_5039000_3682000# GND efet w=48500 l=8500
+ ad=0 pd=0 as=1.997e+09 ps=418000 
M4174 diff_5039000_3682000# diff_5048000_3693000# diff_128000_4097000# GND efet w=79500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4175 diff_5264000_3945000# diff_72000_4515000# diff_4241000_2640000# GND efet w=12000 l=11000
+ ad=2.14e+08 pd=68000 as=-2.01197e+09 ps=470000 
M4176 diff_5763000_4184000# diff_5039000_4962000# diff_83000_3098000# GND efet w=41000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4177 diff_5983000_3917000# diff_5763000_4184000# diff_83000_3098000# GND efet w=49500 l=7500
+ ad=2.056e+09 pd=364000 as=0 ps=0 
M4178 diff_95000_5192000# diff_5983000_3917000# diff_5983000_3917000# GND efet w=13000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M4179 diff_5501000_3807000# diff_4927000_3400000# diff_83000_3098000# GND efet w=102000 l=8000
+ ad=9.18e+08 pd=222000 as=0 ps=0 
M4180 diff_5501000_3807000# diff_5321000_3744000# diff_5356000_4071000# GND efet w=102500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4181 diff_95000_5192000# diff_5356000_4071000# diff_5356000_4071000# GND efet w=13000 l=35000
+ ad=0 pd=0 as=0 ps=0 
M4182 diff_5356000_4071000# diff_5228000_3879000# diff_5501000_3768000# GND efet w=104000 l=9000
+ ad=0 pd=0 as=9.43e+08 ps=226000 
M4183 diff_5356000_4071000# diff_68000_5288000# diff_5678000_3740000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=2.86e+08 ps=70000 
M4184 diff_5983000_3917000# diff_5068000_4962000# diff_83000_3098000# GND efet w=56000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4185 diff_6161000_3828000# diff_6151000_3839000# diff_5983000_3917000# GND efet w=89000 l=9000
+ ad=2.066e+09 pd=436000 as=0 ps=0 
M4186 diff_6161000_3828000# diff_3569000_3530000# diff_83000_3098000# GND efet w=89000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4187 diff_6161000_3828000# diff_6155000_3762000# diff_83000_3098000# GND efet w=86000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4188 diff_5228000_3879000# diff_5008000_3739000# diff_83000_3098000# GND efet w=49000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4189 diff_5501000_3768000# diff_5491000_3760000# diff_83000_3098000# GND efet w=103500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4190 diff_3569000_3530000# diff_3569000_3530000# diff_95000_5192000# GND efet w=13000 l=23000
+ ad=9.36e+08 pd=144000 as=0 ps=0 
M4191 diff_4241000_2640000# diff_72000_4515000# diff_5491000_3760000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=2.49e+08 ps=84000 
M4192 diff_95000_5192000# diff_5043000_3671000# diff_5043000_3671000# GND efet w=11000 l=37000
+ ad=0 pd=0 as=8.87e+08 ps=188000 
M4193 diff_83000_3098000# diff_5043000_3671000# diff_5039000_3682000# GND efet w=136000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4194 diff_5043000_3671000# diff_4927000_3400000# diff_83000_3098000# GND efet w=41000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4195 diff_5321000_3744000# diff_68000_5288000# diff_817000_1965000# GND efet w=12000 l=12000
+ ad=2.69e+08 pd=68000 as=0 ps=0 
M4196 diff_95000_5192000# diff_4241000_2640000# diff_4241000_2640000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M4197 diff_4241000_2640000# diff_5678000_3740000# diff_83000_3098000# GND efet w=65000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4198 diff_83000_3098000# diff_5098000_4894000# diff_3569000_3530000# GND efet w=68500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4199 diff_5293000_3706000# diff_68000_5288000# diff_817000_1663000# GND efet w=12000 l=11000
+ ad=3.26e+08 pd=98000 as=0 ps=0 
M4200 diff_83000_3098000# diff_5293000_3706000# diff_5397000_3688000# GND efet w=97000 l=8000
+ ad=0 pd=0 as=8.92e+08 ps=212000 
M4201 diff_83000_3098000# diff_5009000_4962000# diff_6155000_3780000# GND efet w=86000 l=8000
+ ad=0 pd=0 as=7.74e+08 ps=190000 
M4202 diff_6155000_3780000# diff_4303000_2657000# diff_6155000_3762000# GND efet w=86000 l=8000
+ ad=0 pd=0 as=1.713e+09 ps=334000 
M4203 diff_6155000_3762000# diff_6146000_3754000# diff_83000_3098000# GND efet w=45000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4204 diff_95000_5192000# diff_6155000_3762000# diff_6155000_3762000# GND efet w=13000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M4205 diff_6146000_3754000# diff_4303000_2657000# diff_83000_3098000# GND efet w=44000 l=8000
+ ad=1.902e+09 pd=412000 as=0 ps=0 
M4206 diff_95000_5192000# diff_6146000_3754000# diff_6146000_3754000# GND efet w=11000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M4207 diff_6146000_3754000# diff_5009000_4962000# diff_83000_3098000# GND efet w=40000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4208 diff_5397000_3688000# diff_4927000_3400000# diff_5397000_3662000# GND efet w=96500 l=8500
+ ad=0 pd=0 as=1.91033e+08 ps=850000 
M4209 diff_4871000_3351000# diff_4927000_3400000# diff_83000_3098000# GND efet w=47500 l=8500
+ ad=-1.91497e+09 pd=414000 as=0 ps=0 
M4210 diff_83000_3098000# diff_5022000_3615000# diff_4871000_3351000# GND efet w=43000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M4211 diff_5022000_3615000# diff_72000_4515000# diff_4806000_4501000# GND efet w=12000 l=12000
+ ad=3.95e+08 pd=128000 as=0 ps=0 
M4212 diff_95000_5192000# diff_5228000_3587000# diff_5228000_3587000# GND efet w=13000 l=36000
+ ad=0 pd=0 as=-1.09097e+09 ps=742000 
M4213 diff_95000_5192000# diff_5397000_3662000# diff_5397000_3662000# GND efet w=13000 l=38000
+ ad=0 pd=0 as=0 ps=0 
M4214 diff_5397000_3662000# diff_5371000_3654000# diff_5397000_3644000# GND efet w=97000 l=8000
+ ad=0 pd=0 as=8.69e+08 ps=210000 
M4215 diff_5397000_3662000# diff_5228000_3587000# diff_5513000_3639000# GND efet w=55000 l=8000
+ ad=0 pd=0 as=1.261e+09 ps=300000 
M4216 diff_5397000_3644000# diff_5061000_3959000# diff_83000_3098000# GND efet w=96500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4217 diff_5228000_3587000# diff_5061000_3959000# diff_83000_3098000# GND efet w=42000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4218 diff_5513000_3639000# diff_5504000_3630000# diff_83000_3098000# GND efet w=115500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4219 diff_5397000_3662000# diff_68000_5288000# diff_5660000_3640000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=3.18e+08 ps=110000 
M4220 diff_5397000_3662000# diff_5228000_3587000# diff_5513000_3639000# GND efet w=26000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4221 diff_4303000_2657000# diff_5660000_3640000# diff_83000_3098000# GND efet w=62000 l=8000
+ ad=1.855e+09 pd=398000 as=0 ps=0 
M4222 diff_83000_3098000# diff_4927000_3400000# diff_5228000_3587000# GND efet w=41000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4223 diff_95000_5192000# diff_4871000_3351000# diff_4871000_3351000# GND efet w=12000 l=35000
+ ad=0 pd=0 as=0 ps=0 
M4224 diff_6151000_3839000# diff_3569000_3530000# diff_6185000_3575000# GND efet w=144000 l=9000
+ ad=-2.01297e+09 pd=446000 as=-1.81497e+09 ps=484000 
M4225 diff_4303000_2657000# diff_72000_4515000# diff_5504000_3630000# GND efet w=13000 l=11000
+ ad=0 pd=0 as=2.38e+08 ps=70000 
M4226 diff_95000_5192000# diff_4303000_2657000# diff_4303000_2657000# GND efet w=11000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4227 diff_6017000_3581000# diff_6017000_3581000# diff_95000_5192000# GND efet w=12000 l=35000
+ ad=1.666e+09 pd=342000 as=0 ps=0 
M4228 diff_83000_3098000# diff_5009000_4962000# diff_6185000_3600000# GND efet w=143500 l=8500
+ ad=0 pd=0 as=1.287e+09 ps=304000 
M4229 diff_83000_3098000# diff_4182000_2528000# diff_6017000_3581000# GND efet w=42000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4230 diff_6185000_3600000# diff_4182000_2528000# diff_6185000_3575000# GND efet w=143000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4231 diff_6017000_3581000# diff_5009000_4962000# diff_83000_3098000# GND efet w=41000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4232 diff_6185000_3575000# diff_6017000_3581000# diff_83000_3098000# GND efet w=71000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4233 diff_6151000_3839000# diff_6151000_3839000# diff_95000_5192000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M4234 diff_83000_3098000# diff_4927000_3400000# diff_5357000_3322000# GND efet w=43000 l=9000
+ ad=0 pd=0 as=-8.06967e+08 ps=674000 
M4235 diff_83000_3098000# diff_4927000_3400000# diff_5472000_3486000# GND efet w=94000 l=9000
+ ad=0 pd=0 as=7.52e+08 ps=204000 
M4236 diff_5472000_3486000# diff_5294000_3449000# diff_5048000_3693000# GND efet w=94000 l=9000
+ ad=0 pd=0 as=-1.88893e+09 ps=1.254e+06 
M4237 diff_6112000_3388000# diff_4241000_2640000# diff_6160000_3507000# GND efet w=87000 l=8000
+ ad=-9.07967e+08 pd=730000 as=6.96e+08 ps=190000 
M4238 diff_6160000_3507000# diff_5098000_4894000# diff_83000_3098000# GND efet w=87000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4239 diff_5294000_3449000# diff_68000_5288000# diff_817000_1588000# GND efet w=14000 l=11000
+ ad=2.5e+08 pd=98000 as=0 ps=0 
M4240 diff_5048000_3693000# diff_5432000_3451000# diff_5439000_3442000# GND efet w=97000 l=9000
+ ad=0 pd=0 as=8.73e+08 ps=212000 
M4241 diff_5048000_3693000# diff_68000_5288000# diff_5578000_3393000# GND efet w=13000 l=11000
+ ad=0 pd=0 as=3.32e+08 ps=80000 
M4242 diff_95000_5192000# diff_5048000_3693000# diff_5048000_3693000# GND efet w=12000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M4243 diff_95000_5192000# diff_6112000_3388000# diff_6112000_3388000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M4244 diff_83000_3098000# diff_3408000_4288000# diff_6160000_3457000# GND efet w=90500 l=8500
+ ad=0 pd=0 as=8.28e+08 ps=200000 
M4245 diff_4591000_3170000# diff_531000_4622000# diff_83000_3098000# GND efet w=67000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4246 diff_83000_3098000# diff_65000_4220000# diff_4591000_3170000# GND efet w=77500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4247 diff_4779000_3198000# diff_72000_4515000# diff_4697000_3226000# GND efet w=12000 l=11000
+ ad=5.25e+08 pd=146000 as=0 ps=0 
M4248 diff_83000_3098000# diff_3043000_2723000# diff_3256000_1459000# GND efet w=123500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4249 diff_3283000_1426000# diff_3043000_2723000# diff_83000_3098000# GND efet w=100000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4250 diff_83000_3098000# diff_3321000_2527000# diff_3283000_1426000# GND efet w=126000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4251 diff_3401000_3461000# diff_72000_4515000# diff_3383000_2778000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=9.01e+08 ps=148000 
M4252 diff_3433000_2818000# diff_72000_4515000# diff_3433000_2778000# GND efet w=20000 l=13000
+ ad=0 pd=0 as=9.36e+08 ps=150000 
M4253 diff_3506000_2818000# diff_72000_4515000# diff_3486000_2778000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=9.01e+08 ps=148000 
M4254 diff_3536000_2818000# diff_72000_4515000# diff_3536000_2778000# GND efet w=20000 l=13000
+ ad=0 pd=0 as=9.28e+08 ps=150000 
M4255 diff_3609000_2818000# diff_72000_4515000# diff_3589000_2778000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=9.09e+08 ps=148000 
M4256 diff_3639000_2818000# diff_72000_4515000# diff_3639000_2778000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=9.24e+08 ps=150000 
M4257 diff_3712000_2818000# diff_72000_4515000# diff_3692000_2778000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=9.01e+08 ps=148000 
M4258 diff_3742000_2818000# diff_72000_4515000# diff_3742000_2778000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=9.24e+08 ps=150000 
M4259 diff_3815000_2818000# diff_72000_4515000# diff_3794000_2778000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=9.31e+08 ps=150000 
M4260 diff_3846000_2818000# diff_72000_4515000# diff_3846000_2778000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=9.01e+08 ps=148000 
M4261 diff_3667000_4701000# diff_72000_4515000# diff_3898000_2778000# GND efet w=20000 l=13000
+ ad=0 pd=0 as=9.36e+08 ps=150000 
M4262 diff_3949000_2818000# diff_72000_4515000# diff_3949000_2778000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=9.23e+08 ps=150000 
M4263 diff_4022000_2818000# diff_72000_4515000# diff_4001000_2778000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=9.24e+08 ps=150000 
M4264 diff_4052000_2818000# diff_72000_4515000# diff_4052000_2778000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=9.24e+08 ps=150000 
M4265 diff_4125000_2818000# diff_72000_4515000# diff_4104000_2778000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=9.23e+08 ps=150000 
M4266 diff_3354000_2409000# diff_3354000_2409000# diff_95000_5192000# GND efet w=17000 l=8000
+ ad=1.29103e+09 pd=1.114e+06 as=0 ps=0 
M4267 diff_3354000_2409000# diff_72000_4515000# diff_83000_3098000# GND efet w=203000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4268 diff_83000_3098000# diff_3383000_2778000# diff_3354000_2409000# GND efet w=244500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4269 diff_3439000_2492000# diff_3433000_2778000# diff_83000_3098000# GND efet w=244000 l=8000
+ ad=8.13033e+08 pd=888000 as=0 ps=0 
M4270 diff_95000_5192000# diff_3439000_2492000# diff_3439000_2492000# GND efet w=18000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4271 diff_3489000_2725000# diff_3489000_2725000# diff_95000_5192000# GND efet w=18000 l=8000
+ ad=7.28033e+08 pd=886000 as=0 ps=0 
M4272 diff_83000_3098000# diff_72000_4515000# diff_3439000_2492000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4273 diff_2683000_2215000# diff_2674000_2207000# diff_83000_3098000# GND efet w=218500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4274 diff_1399000_598000# diff_2713000_822000# diff_2683000_2215000# GND efet w=103000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4275 diff_2532000_2143000# diff_2448000_2717000# diff_2471000_2112000# GND efet w=21000 l=12000
+ ad=1.589e+09 pd=340000 as=3.22e+08 ps=80000 
M4276 diff_2130000_2043000# diff_2471000_2112000# diff_83000_3098000# GND efet w=58000 l=7000
+ ad=1.394e+09 pd=304000 as=0 ps=0 
M4277 diff_83000_3098000# diff_1757000_739000# diff_2532000_2143000# GND efet w=78500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4278 diff_95000_5192000# diff_1438000_786000# diff_1757000_739000# GND efet w=86500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4279 diff_848000_2016000# diff_1438000_786000# diff_95000_5192000# GND efet w=71000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4280 diff_817000_2342000# diff_2775000_765000# diff_2683000_2215000# GND efet w=107000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4281 diff_2829000_2242000# diff_2583000_2725000# diff_817000_2342000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4282 diff_2915000_2318000# diff_2939000_824000# diff_817000_2342000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4283 diff_2915000_2318000# diff_2915000_2318000# diff_2915000_2318000# GND efet w=1000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4284 diff_2829000_2242000# diff_2843000_1950000# diff_848000_2342000# GND efet w=106500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4285 diff_2683000_2153000# diff_2674000_2144000# diff_83000_3098000# GND efet w=218500 l=8500
+ ad=-2.45967e+08 pd=718000 as=0 ps=0 
M4286 diff_2674000_2144000# diff_2651000_2077000# diff_83000_3098000# GND efet w=66000 l=8000
+ ad=8.86e+08 pd=194000 as=0 ps=0 
M4287 diff_1757000_739000# diff_2713000_822000# diff_2683000_2153000# GND efet w=103000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4288 diff_2532000_2143000# diff_2532000_2143000# diff_95000_5192000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M4289 diff_2320000_2130000# diff_2320000_2130000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4290 diff_95000_5192000# diff_2320000_1883000# diff_2320000_1883000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=-1.94197e+09 ps=426000 
M4291 diff_2130000_2043000# diff_2130000_2043000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4292 diff_95000_5192000# diff_2130000_1972000# diff_2130000_1972000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=1.403e+09 ps=310000 
M4293 diff_2320000_1883000# diff_1094000_1020000# diff_2406000_1946000# GND efet w=150500 l=8500
+ ad=0 pd=0 as=1.525e+09 ps=306000 
M4294 diff_83000_3098000# diff_2320000_1883000# diff_2281000_1866000# GND efet w=56000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M4295 diff_2304000_1746000# diff_2320000_1883000# diff_83000_3098000# GND efet w=152500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4296 diff_2406000_1946000# diff_2130000_1972000# diff_83000_3098000# GND efet w=120000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4297 diff_2304000_1746000# diff_2330000_1775000# diff_83000_3098000# GND efet w=151000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4298 diff_83000_3098000# diff_2304000_1746000# diff_2127000_1545000# GND efet w=161500 l=7500
+ ad=0 pd=0 as=1.31033e+08 ps=784000 
M4299 diff_2127000_1705000# diff_1237000_1921000# diff_95000_5192000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4300 diff_2184000_1679000# diff_2184000_1679000# diff_95000_5192000# GND efet w=12000 l=18000
+ ad=0 pd=0 as=0 ps=0 
M4301 diff_2102000_1637000# diff_1438000_786000# diff_2050000_1770000# GND efet w=21000 l=13000
+ ad=1.47e+08 pd=56000 as=3.84e+08 ps=90000 
M4302 diff_2122000_1637000# diff_72000_4515000# diff_2102000_1637000# GND efet w=21000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M4303 diff_95000_5192000# diff_2122000_1637000# diff_2122000_1637000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M4304 diff_2102000_1607000# diff_1438000_786000# diff_2050000_1457000# GND efet w=21000 l=13000
+ ad=1.47e+08 pd=56000 as=3.57e+08 ps=96000 
M4305 diff_2122000_1607000# diff_72000_4515000# diff_2102000_1607000# GND efet w=21000 l=13000
+ ad=-1.35397e+09 pd=438000 as=0 ps=0 
M4306 diff_1851000_1456000# diff_1487000_841000# diff_1997000_1468000# GND efet w=120000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4307 diff_83000_3098000# diff_1881000_1450000# diff_1850000_1535000# GND efet w=198500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4308 diff_1881000_1450000# diff_1932000_1554000# diff_83000_3098000# GND efet w=59000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4309 diff_1851000_1317000# diff_1858000_1019000# diff_1851000_1376000# GND efet w=105000 l=10000
+ ad=-1.29967e+08 pd=724000 as=9.99065e+08 ps=1.896e+06 
M4310 diff_83000_3098000# diff_1881000_1418000# diff_1851000_1317000# GND efet w=198500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4311 diff_1851000_1317000# diff_1837000_1364000# diff_817000_1286000# GND efet w=102500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4312 diff_1881000_1418000# diff_1932000_1328000# diff_83000_3098000# GND efet w=64000 l=8000
+ ad=1.198e+09 pd=210000 as=0 ps=0 
M4313 diff_1997000_1468000# diff_2050000_1457000# diff_83000_3098000# GND efet w=183500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4314 diff_1851000_1376000# diff_1487000_841000# diff_1997000_1362000# GND efet w=117000 l=10000
+ ad=0 pd=0 as=-1.21797e+09 ps=668000 
M4315 diff_1997000_1362000# diff_2050000_1393000# diff_83000_3098000# GND efet w=185500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4316 diff_1850000_1158000# diff_1837000_1364000# diff_817000_1211000# GND efet w=102500 l=9500
+ ad=-1.01967e+08 pd=736000 as=0 ps=0 
M4317 diff_1997000_1362000# diff_1547000_932000# diff_1932000_1328000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=8.35e+08 ps=200000 
M4318 diff_1851000_1317000# diff_95000_5192000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M4319 diff_1932000_1328000# diff_95000_5192000# diff_1851000_1317000# GND efet w=12500 l=80500
+ ad=0 pd=0 as=0 ps=0 
M4320 diff_1881000_1418000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=31000
+ ad=0 pd=0 as=0 ps=0 
M4321 diff_1932000_1177000# diff_95000_5192000# diff_1850000_1158000# GND efet w=13000 l=76000
+ ad=8.85e+08 pd=212000 as=0 ps=0 
M4322 diff_95000_5192000# diff_95000_5192000# diff_1850000_1158000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M4323 diff_95000_5192000# diff_95000_5192000# diff_1881000_1073000# GND efet w=13000 l=32000
+ ad=0 pd=0 as=1.074e+09 ps=212000 
M4324 diff_1850000_1158000# diff_1858000_1019000# diff_1851000_1079000# GND efet w=104500 l=10500
+ ad=0 pd=0 as=1.22907e+09 ps=1.978e+06 
M4325 diff_1997000_1362000# diff_1997000_1362000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4326 diff_95000_5192000# diff_1997000_1091000# diff_1997000_1091000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=-1.31697e+09 ps=664000 
M4327 diff_1997000_1091000# diff_1547000_932000# diff_1932000_1177000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4328 diff_95000_5192000# diff_2122000_1607000# diff_2122000_1607000# GND efet w=10000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M4329 diff_2122000_1607000# diff_2130000_1595000# diff_2137000_1580000# GND efet w=65000 l=8000
+ ad=0 pd=0 as=1.845e+09 ps=380000 
M4330 diff_95000_5192000# diff_2184000_1494000# diff_2184000_1494000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=1.595e+09 ps=340000 
M4331 diff_2137000_1580000# diff_2127000_1545000# diff_83000_3098000# GND efet w=126500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4332 diff_2122000_1607000# diff_2130000_1595000# diff_2137000_1580000# GND efet w=73500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4333 diff_83000_3098000# diff_2184000_1494000# diff_2122000_1607000# GND efet w=57000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4334 diff_2184000_1494000# diff_2130000_1595000# diff_83000_3098000# GND efet w=63000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4335 diff_83000_3098000# diff_2127000_1545000# diff_2184000_1494000# GND efet w=71000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4336 diff_2137000_1296000# diff_2127000_1328000# diff_83000_3098000# GND efet w=128000 l=8000
+ ad=1.93e+09 pd=382000 as=0 ps=0 
M4337 diff_2121000_1261000# diff_2130000_1289000# diff_2137000_1296000# GND efet w=76000 l=8000
+ ad=-1.22397e+09 pd=466000 as=0 ps=0 
M4338 diff_2137000_1296000# diff_2130000_1289000# diff_2121000_1261000# GND efet w=62500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4339 diff_83000_3098000# diff_2184000_1302000# diff_2121000_1261000# GND efet w=57000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4340 diff_2184000_1302000# diff_2130000_1289000# diff_83000_3098000# GND efet w=63000 l=8000
+ ad=1.617e+09 pd=336000 as=0 ps=0 
M4341 diff_83000_3098000# diff_2127000_1328000# diff_2184000_1302000# GND efet w=71000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4342 diff_2184000_1302000# diff_2184000_1302000# diff_95000_5192000# GND efet w=12000 l=18000
+ ad=0 pd=0 as=0 ps=0 
M4343 diff_2102000_1261000# diff_1438000_786000# diff_2050000_1393000# GND efet w=20000 l=13000
+ ad=1.4e+08 pd=54000 as=3.64e+08 ps=88000 
M4344 diff_2121000_1261000# diff_72000_4515000# diff_2102000_1261000# GND efet w=20000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4345 diff_95000_5192000# diff_2121000_1261000# diff_2121000_1261000# GND efet w=11000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M4346 diff_2460000_1833000# diff_1037000_877000# diff_2320000_1883000# GND efet w=151000 l=8000
+ ad=1.685e+09 pd=328000 as=0 ps=0 
M4347 diff_817000_2040000# diff_1438000_786000# diff_95000_5192000# GND efet w=87500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4348 diff_2651000_2077000# diff_2641000_934000# diff_817000_2040000# GND efet w=20000 l=10000
+ ad=5.15e+08 pd=178000 as=0 ps=0 
M4349 diff_817000_2040000# diff_2775000_765000# diff_2683000_2153000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4350 diff_83000_3098000# diff_2876000_2205000# diff_2829000_2242000# GND efet w=215500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4351 diff_2876000_2205000# diff_2915000_2318000# diff_83000_3098000# GND efet w=59500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4352 diff_817000_1965000# diff_1438000_786000# diff_95000_5192000# GND efet w=88500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4353 diff_83000_3098000# diff_2471000_1828000# diff_2460000_1833000# GND efet w=124500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4354 diff_2130000_1972000# diff_2471000_1828000# diff_83000_3098000# GND efet w=59000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M4355 diff_95000_5192000# diff_2531000_1855000# diff_2531000_1855000# GND efet w=11000 l=14000
+ ad=0 pd=0 as=1.641e+09 ps=346000 
M4356 diff_2674000_2144000# diff_95000_5192000# diff_95000_5192000# GND efet w=11000 l=31000
+ ad=0 pd=0 as=0 ps=0 
M4357 diff_2683000_2153000# diff_95000_5192000# diff_2651000_2077000# GND efet w=12500 l=80500
+ ad=0 pd=0 as=0 ps=0 
M4358 diff_2683000_2153000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4359 diff_95000_5192000# diff_95000_5192000# diff_2674000_1831000# GND efet w=11000 l=30000
+ ad=0 pd=0 as=9.06e+08 ps=196000 
M4360 diff_2683000_1839000# diff_95000_5192000# diff_2650000_1921000# GND efet w=12000 l=72000
+ ad=-2.25967e+08 pd=738000 as=5.56e+08 ps=192000 
M4361 diff_95000_5192000# diff_95000_5192000# diff_2683000_1839000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4362 diff_2650000_1921000# diff_2641000_934000# diff_817000_1965000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4363 diff_2829000_2070000# diff_2583000_2725000# diff_817000_2040000# GND efet w=86000 l=10000
+ ad=-1.32967e+08 pd=720000 as=0 ps=0 
M4364 diff_2829000_2070000# diff_2843000_1950000# diff_848000_2016000# GND efet w=106500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4365 diff_83000_3098000# diff_2876000_2170000# diff_2829000_2070000# GND efet w=214500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4366 diff_2876000_2170000# diff_2914000_2058000# diff_83000_3098000# GND efet w=68500 l=7500
+ ad=8.9e+08 pd=182000 as=0 ps=0 
M4367 diff_817000_2342000# diff_2638000_2492000# diff_3029000_2300000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=1.619e+09 ps=392000 
M4368 diff_95000_5192000# diff_95000_5192000# diff_3099000_2319000# GND efet w=12000 l=30000
+ ad=0 pd=0 as=9.79e+08 ps=200000 
M4369 diff_3117000_2217000# diff_95000_5192000# diff_3029000_2300000# GND efet w=12000 l=72000
+ ad=-3.04967e+08 pd=706000 as=0 ps=0 
M4370 diff_95000_5192000# diff_95000_5192000# diff_3117000_2217000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4371 diff_848000_2342000# diff_2996000_2725000# diff_2915000_2318000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4372 diff_3029000_2300000# diff_2996000_2725000# diff_1399000_598000# GND efet w=19000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4373 diff_3029000_2041000# diff_2996000_2725000# diff_1757000_739000# GND efet w=19000 l=10000
+ ad=1.548e+09 pd=370000 as=0 ps=0 
M4374 diff_848000_2016000# diff_2996000_2725000# diff_2914000_2058000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=1.224e+09 ps=306000 
M4375 diff_2829000_2070000# diff_95000_5192000# diff_95000_5192000# GND efet w=11000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4376 diff_2914000_2058000# diff_95000_5192000# diff_2829000_2070000# GND efet w=12500 l=80500
+ ad=0 pd=0 as=0 ps=0 
M4377 diff_2876000_2170000# diff_95000_5192000# diff_95000_5192000# GND efet w=11000 l=31000
+ ad=0 pd=0 as=0 ps=0 
M4378 diff_2914000_2058000# diff_2939000_824000# diff_817000_2040000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4379 diff_95000_5192000# diff_95000_5192000# diff_2829000_1865000# GND efet w=11000 l=22000
+ ad=0 pd=0 as=-8.9673e+06 ps=738000 
M4380 diff_2915000_1942000# diff_95000_5192000# diff_2829000_1865000# GND efet w=12000 l=71000
+ ad=1.226e+09 pd=312000 as=0 ps=0 
M4381 diff_95000_5192000# diff_95000_5192000# diff_2876000_1829000# GND efet w=12000 l=29000
+ ad=0 pd=0 as=8.52e+08 ps=188000 
M4382 diff_83000_3098000# diff_1774000_760000# diff_2531000_1855000# GND efet w=83500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4383 diff_2531000_1855000# diff_2448000_2717000# diff_2471000_1828000# GND efet w=21000 l=11000
+ ad=0 pd=0 as=3.71e+08 ps=96000 
M4384 diff_2407000_1692000# diff_2130000_1666000# diff_83000_3098000# GND efet w=115500 l=8500
+ ad=1.515e+09 pd=296000 as=0 ps=0 
M4385 diff_2330000_1775000# diff_1094000_1020000# diff_2407000_1692000# GND efet w=146500 l=8500
+ ad=-1.91097e+09 pd=416000 as=0 ps=0 
M4386 diff_2460000_1725000# diff_1037000_877000# diff_2330000_1775000# GND efet w=150000 l=8000
+ ad=1.659e+09 pd=326000 as=0 ps=0 
M4387 diff_83000_3098000# diff_2471000_1736000# diff_2460000_1725000# GND efet w=123500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4388 diff_95000_5192000# diff_1438000_786000# diff_1774000_760000# GND efet w=85500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4389 diff_848000_1965000# diff_1438000_786000# diff_95000_5192000# GND efet w=71000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4390 diff_2674000_1831000# diff_2650000_1921000# diff_83000_3098000# GND efet w=61000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4391 diff_2683000_1839000# diff_2674000_1831000# diff_83000_3098000# GND efet w=217500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4392 diff_1774000_760000# diff_2713000_822000# diff_2683000_1839000# GND efet w=103000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4393 diff_2531000_1766000# diff_2448000_2717000# diff_2471000_1736000# GND efet w=21000 l=11000
+ ad=1.606e+09 pd=340000 as=3.21e+08 ps=80000 
M4394 diff_2127000_1545000# diff_1237000_1921000# diff_95000_5192000# GND efet w=12000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4395 diff_2127000_1328000# diff_2291000_1482000# diff_2127000_1545000# GND efet w=122000 l=10000
+ ad=2.33033e+08 pd=702000 as=0 ps=0 
M4396 diff_95000_5192000# diff_2291000_1482000# diff_2291000_1482000# GND efet w=13000 l=20000
+ ad=0 pd=0 as=1.057e+09 ps=214000 
M4397 diff_2130000_1666000# diff_2471000_1736000# diff_83000_3098000# GND efet w=58000 l=7000
+ ad=1.387e+09 pd=302000 as=0 ps=0 
M4398 diff_83000_3098000# diff_1791000_798000# diff_2531000_1766000# GND efet w=79000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4399 diff_95000_5192000# diff_1438000_786000# diff_1791000_798000# GND efet w=86500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4400 diff_848000_1639000# diff_1438000_786000# diff_95000_5192000# GND efet w=72000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4401 diff_817000_1965000# diff_2775000_765000# diff_2683000_1839000# GND efet w=107500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4402 diff_2829000_1865000# diff_2583000_2725000# diff_817000_1965000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4403 diff_2915000_1942000# diff_2939000_824000# diff_817000_1965000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4404 diff_2915000_1942000# diff_2915000_1942000# diff_2915000_1942000# GND efet w=500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4405 diff_2829000_1865000# diff_2843000_1950000# diff_848000_1965000# GND efet w=107000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4406 diff_2683000_1777000# diff_2674000_1768000# diff_83000_3098000# GND efet w=219500 l=8500
+ ad=-3.11967e+08 pd=722000 as=0 ps=0 
M4407 diff_2674000_1768000# diff_2651000_1700000# diff_83000_3098000# GND efet w=69000 l=8000
+ ad=9.14e+08 pd=196000 as=0 ps=0 
M4408 diff_1791000_798000# diff_2713000_822000# diff_2683000_1777000# GND efet w=103500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4409 diff_2531000_1766000# diff_2531000_1766000# diff_95000_5192000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M4410 diff_2330000_1775000# diff_2330000_1775000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4411 diff_95000_5192000# diff_2335000_1514000# diff_2335000_1514000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=-1.84397e+09 ps=426000 
M4412 diff_2130000_1666000# diff_2130000_1666000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4413 diff_95000_5192000# diff_2130000_1595000# diff_2130000_1595000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=1.378e+09 ps=310000 
M4414 diff_2335000_1514000# diff_1094000_1020000# diff_2407000_1569000# GND efet w=150000 l=8000
+ ad=0 pd=0 as=1.52e+09 ps=304000 
M4415 diff_83000_3098000# diff_2335000_1514000# diff_2291000_1482000# GND efet w=59000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4416 diff_2407000_1569000# diff_2130000_1595000# diff_83000_3098000# GND efet w=119000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4417 diff_2459000_1456000# diff_1037000_877000# diff_2335000_1514000# GND efet w=151500 l=7500
+ ad=1.764e+09 pd=330000 as=0 ps=0 
M4418 diff_817000_1663000# diff_1438000_786000# diff_95000_5192000# GND efet w=87500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4419 diff_2651000_1700000# diff_2641000_934000# diff_817000_1663000# GND efet w=20000 l=10000
+ ad=5.23e+08 pd=158000 as=0 ps=0 
M4420 diff_817000_1663000# diff_2775000_765000# diff_2683000_1777000# GND efet w=106500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4421 diff_83000_3098000# diff_2876000_1829000# diff_2829000_1865000# GND efet w=213500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4422 diff_2876000_1829000# diff_2915000_1942000# diff_83000_3098000# GND efet w=59500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4423 diff_817000_1588000# diff_1438000_786000# diff_95000_5192000# GND efet w=87500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4424 diff_83000_3098000# diff_2471000_1451000# diff_2459000_1456000# GND efet w=124500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4425 diff_2130000_1595000# diff_2471000_1451000# diff_83000_3098000# GND efet w=59000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M4426 diff_95000_5192000# diff_2531000_1479000# diff_2531000_1479000# GND efet w=11000 l=15000
+ ad=0 pd=0 as=1.614e+09 ps=346000 
M4427 diff_2674000_1768000# diff_95000_5192000# diff_95000_5192000# GND efet w=11000 l=31000
+ ad=0 pd=0 as=0 ps=0 
M4428 diff_2683000_1777000# diff_95000_5192000# diff_2651000_1700000# GND efet w=12500 l=81500
+ ad=0 pd=0 as=0 ps=0 
M4429 diff_2683000_1777000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4430 diff_95000_5192000# diff_95000_5192000# diff_2674000_1454000# GND efet w=11000 l=31000
+ ad=0 pd=0 as=9.03e+08 ps=196000 
M4431 diff_2683000_1461000# diff_95000_5192000# diff_2651000_1545000# GND efet w=12000 l=74000
+ ad=-3.24967e+08 pd=736000 as=5.23e+08 ps=190000 
M4432 diff_95000_5192000# diff_95000_5192000# diff_2683000_1461000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4433 diff_2651000_1545000# diff_2641000_934000# diff_817000_1588000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4434 diff_2829000_1693000# diff_2583000_2725000# diff_817000_1663000# GND efet w=86000 l=10000
+ ad=-1.30967e+08 pd=718000 as=0 ps=0 
M4435 diff_2829000_1693000# diff_2843000_1950000# diff_848000_1639000# GND efet w=104500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4436 diff_83000_3098000# diff_2876000_1793000# diff_2829000_1693000# GND efet w=212500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4437 diff_2876000_1793000# diff_2914000_1681000# diff_83000_3098000# GND efet w=69500 l=7500
+ ad=9.13e+08 pd=184000 as=0 ps=0 
M4438 diff_83000_3098000# diff_2534000_2492000# diff_1399000_598000# GND efet w=106500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4439 diff_3099000_2319000# diff_3029000_2300000# diff_83000_3098000# GND efet w=60500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4440 diff_3117000_2217000# diff_3099000_2319000# diff_83000_3098000# GND efet w=213500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4441 diff_1399000_598000# diff_3120000_2492000# diff_3117000_2217000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4442 diff_817000_2342000# diff_2893000_2725000# diff_3117000_2217000# GND efet w=86000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4443 diff_83000_3098000# diff_2534000_2492000# diff_1757000_739000# GND efet w=106500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4444 diff_3117000_2154000# diff_3099000_2059000# diff_83000_3098000# GND efet w=212500 l=7500
+ ad=-4.81967e+08 pd=684000 as=0 ps=0 
M4445 diff_3099000_2059000# diff_3029000_2041000# diff_83000_3098000# GND efet w=68500 l=8500
+ ad=9.22e+08 pd=196000 as=0 ps=0 
M4446 diff_817000_2040000# diff_2638000_2492000# diff_3029000_2041000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4447 diff_817000_1965000# diff_2638000_2492000# diff_3029000_1923000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=1.616e+09 ps=392000 
M4448 diff_1757000_739000# diff_3120000_2492000# diff_3117000_2154000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4449 diff_817000_2040000# diff_2893000_2725000# diff_3117000_2154000# GND efet w=86000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4450 diff_3099000_2059000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=32000
+ ad=0 pd=0 as=0 ps=0 
M4451 diff_3117000_2154000# diff_95000_5192000# diff_3029000_2041000# GND efet w=12000 l=83000
+ ad=0 pd=0 as=0 ps=0 
M4452 diff_3117000_2154000# diff_95000_5192000# diff_95000_5192000# GND efet w=11000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4453 diff_95000_5192000# diff_95000_5192000# diff_3099000_1943000# GND efet w=12000 l=30000
+ ad=0 pd=0 as=9.76e+08 ps=200000 
M4454 diff_3117000_1841000# diff_95000_5192000# diff_3029000_1923000# GND efet w=12000 l=70000
+ ad=-2.87967e+08 pd=710000 as=0 ps=0 
M4455 diff_95000_5192000# diff_95000_5192000# diff_3117000_1841000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4456 diff_848000_1965000# diff_2996000_2725000# diff_2915000_1942000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4457 diff_3029000_1923000# diff_2996000_2725000# diff_1774000_760000# GND efet w=19000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4458 diff_3029000_1664000# diff_2996000_2725000# diff_1791000_798000# GND efet w=19000 l=10000
+ ad=1.547e+09 pd=370000 as=0 ps=0 
M4459 diff_848000_1639000# diff_2996000_2725000# diff_2914000_1681000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=1.221e+09 ps=310000 
M4460 diff_2829000_1693000# diff_95000_5192000# diff_95000_5192000# GND efet w=11000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4461 diff_2914000_1681000# diff_95000_5192000# diff_2829000_1693000# GND efet w=12500 l=80500
+ ad=0 pd=0 as=0 ps=0 
M4462 diff_2876000_1793000# diff_95000_5192000# diff_95000_5192000# GND efet w=11000 l=31000
+ ad=0 pd=0 as=0 ps=0 
M4463 diff_2914000_1681000# diff_2939000_824000# diff_817000_1663000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4464 diff_95000_5192000# diff_95000_5192000# diff_2829000_1488000# GND efet w=11000 l=22000
+ ad=0 pd=0 as=-5.59673e+07 ps=732000 
M4465 diff_2915000_1565000# diff_95000_5192000# diff_2829000_1488000# GND efet w=12000 l=73000
+ ad=1.221e+09 pd=310000 as=0 ps=0 
M4466 diff_95000_5192000# diff_95000_5192000# diff_2876000_1451000# GND efet w=12000 l=30000
+ ad=0 pd=0 as=8.62e+08 ps=188000 
M4467 diff_83000_3098000# diff_1851000_1456000# diff_2531000_1479000# GND efet w=83000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4468 diff_2531000_1479000# diff_2448000_2717000# diff_2471000_1451000# GND efet w=20000 l=12000
+ ad=0 pd=0 as=3.31e+08 ps=92000 
M4469 diff_2127000_1169000# diff_2290000_1294000# diff_2127000_1328000# GND efet w=123000 l=10000
+ ad=-5.54967e+08 pd=732000 as=0 ps=0 
M4470 diff_2102000_1230000# diff_1438000_786000# diff_2050000_1081000# GND efet w=21000 l=13000
+ ad=1.47e+08 pd=56000 as=3.49e+08 ps=98000 
M4471 diff_2121000_1230000# diff_72000_4515000# diff_2102000_1230000# GND efet w=21000 l=12000
+ ad=-1.30597e+09 pd=440000 as=0 ps=0 
M4472 diff_1851000_1079000# diff_1487000_841000# diff_1997000_1091000# GND efet w=120000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4473 diff_83000_3098000# diff_1881000_1073000# diff_1850000_1158000# GND efet w=197500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4474 diff_1881000_1073000# diff_1932000_1177000# diff_83000_3098000# GND efet w=59000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4475 diff_1850000_941000# diff_1858000_1019000# diff_1851000_999000# GND efet w=105000 l=10000
+ ad=-2.15967e+08 pd=720000 as=4.21065e+08 ps=1.768e+06 
M4476 diff_83000_3098000# diff_1881000_1041000# diff_1850000_941000# GND efet w=197500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4477 diff_1850000_941000# diff_1837000_1364000# diff_817000_909000# GND efet w=101500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4478 diff_1881000_1041000# diff_1931000_949000# diff_83000_3098000# GND efet w=63000 l=8000
+ ad=1.166e+09 pd=208000 as=0 ps=0 
M4479 diff_1997000_1091000# diff_2050000_1081000# diff_83000_3098000# GND efet w=181500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4480 diff_1851000_999000# diff_1487000_841000# diff_1997000_985000# GND efet w=116500 l=9500
+ ad=0 pd=0 as=-1.18797e+09 ps=670000 
M4481 diff_1997000_985000# diff_2050000_1017000# diff_83000_3098000# GND efet w=186500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4482 diff_1997000_985000# diff_1547000_932000# diff_1931000_949000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=8.3e+08 ps=198000 
M4483 diff_1850000_941000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4484 diff_1931000_949000# diff_95000_5192000# diff_1850000_941000# GND efet w=11500 l=83500
+ ad=0 pd=0 as=0 ps=0 
M4485 diff_1881000_1041000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=32000
+ ad=0 pd=0 as=0 ps=0 
M4486 diff_1997000_985000# diff_1997000_985000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M4487 diff_95000_5192000# diff_2121000_1230000# diff_2121000_1230000# GND efet w=11000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M4488 diff_2127000_1328000# diff_1237000_1921000# diff_95000_5192000# GND efet w=12000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4489 diff_95000_5192000# diff_1237000_1921000# diff_2127000_1169000# GND efet w=12000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4490 diff_2121000_1230000# diff_2130000_1219000# diff_2137000_1204000# GND efet w=65500 l=7500
+ ad=0 pd=0 as=1.807e+09 ps=380000 
M4491 diff_95000_5192000# diff_2184000_1118000# diff_2184000_1118000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=1.6e+09 ps=340000 
M4492 diff_2137000_1204000# diff_2127000_1169000# diff_83000_3098000# GND efet w=126000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4493 diff_2121000_1230000# diff_2130000_1219000# diff_2137000_1204000# GND efet w=73500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4494 diff_83000_3098000# diff_2184000_1118000# diff_2121000_1230000# GND efet w=57000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4495 diff_2184000_1118000# diff_2130000_1219000# diff_83000_3098000# GND efet w=64000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4496 diff_83000_3098000# diff_2127000_1169000# diff_2184000_1118000# GND efet w=72000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4497 diff_2137000_920000# diff_2127000_952000# diff_83000_3098000# GND efet w=129500 l=8500
+ ad=1.877e+09 pd=380000 as=0 ps=0 
M4498 diff_2121000_884000# diff_2130000_913000# diff_2137000_920000# GND efet w=75500 l=8500
+ ad=-1.20397e+09 pd=464000 as=0 ps=0 
M4499 diff_2137000_920000# diff_2130000_913000# diff_2121000_884000# GND efet w=62500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4500 diff_83000_3098000# diff_2184000_926000# diff_2121000_884000# GND efet w=57000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4501 diff_2184000_926000# diff_2130000_913000# diff_83000_3098000# GND efet w=64000 l=8000
+ ad=1.598e+09 pd=334000 as=0 ps=0 
M4502 diff_83000_3098000# diff_2127000_952000# diff_2184000_926000# GND efet w=72000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4503 diff_83000_3098000# diff_2335000_1372000# diff_2290000_1294000# GND efet w=63500 l=7500
+ ad=0 pd=0 as=1.206e+09 ps=222000 
M4504 diff_2406000_1315000# diff_2130000_1289000# diff_83000_3098000# GND efet w=116500 l=8500
+ ad=1.527e+09 pd=298000 as=0 ps=0 
M4505 diff_2335000_1372000# diff_1094000_1020000# diff_2406000_1315000# GND efet w=147000 l=8000
+ ad=-1.80997e+09 pd=416000 as=0 ps=0 
M4506 diff_2459000_1348000# diff_1037000_877000# diff_2335000_1372000# GND efet w=151000 l=8000
+ ad=1.756e+09 pd=330000 as=0 ps=0 
M4507 diff_83000_3098000# diff_2471000_1358000# diff_2459000_1348000# GND efet w=124500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4508 diff_95000_5192000# diff_1438000_786000# diff_1851000_1456000# GND efet w=86500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4509 diff_848000_1588000# diff_1438000_786000# diff_95000_5192000# GND efet w=71000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4510 diff_2674000_1454000# diff_2651000_1545000# diff_83000_3098000# GND efet w=60000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4511 diff_2683000_1461000# diff_2674000_1454000# diff_83000_3098000# GND efet w=217500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4512 diff_1851000_1456000# diff_2713000_822000# diff_2683000_1461000# GND efet w=102500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4513 diff_2531000_1389000# diff_2448000_2717000# diff_2471000_1358000# GND efet w=21000 l=11000
+ ad=1.616e+09 pd=342000 as=3.22e+08 ps=80000 
M4514 diff_2290000_1294000# diff_2290000_1294000# diff_95000_5192000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4515 diff_95000_5192000# diff_2290000_1091000# diff_2290000_1091000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=1.33e+09 ps=242000 
M4516 diff_2127000_952000# diff_2290000_1091000# diff_2127000_1169000# GND efet w=121000 l=10000
+ ad=-1.23297e+09 pd=552000 as=0 ps=0 
M4517 diff_2130000_1289000# diff_2471000_1358000# diff_83000_3098000# GND efet w=59000 l=8000
+ ad=1.316e+09 pd=302000 as=0 ps=0 
M4518 diff_83000_3098000# diff_1851000_1376000# diff_2531000_1389000# GND efet w=79000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4519 diff_95000_5192000# diff_1438000_786000# diff_1851000_1376000# GND efet w=85500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4520 diff_848000_1262000# diff_1438000_786000# diff_95000_5192000# GND efet w=71000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4521 diff_817000_1588000# diff_2775000_765000# diff_2683000_1461000# GND efet w=107500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4522 diff_2829000_1488000# diff_2583000_2725000# diff_817000_1588000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4523 diff_2915000_1565000# diff_2939000_824000# diff_817000_1588000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4524 diff_2915000_1565000# diff_2915000_1565000# diff_2915000_1565000# GND efet w=500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4525 diff_2829000_1488000# diff_2843000_1950000# diff_848000_1588000# GND efet w=105500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4526 diff_2683000_1400000# diff_2674000_1391000# diff_83000_3098000# GND efet w=218500 l=8500
+ ad=-3.98967e+08 pd=720000 as=0 ps=0 
M4527 diff_2674000_1391000# diff_2650000_1323000# diff_83000_3098000# GND efet w=68000 l=8000
+ ad=8.98e+08 pd=194000 as=0 ps=0 
M4528 diff_1851000_1376000# diff_2713000_822000# diff_2683000_1400000# GND efet w=103500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4529 diff_2531000_1389000# diff_2531000_1389000# diff_95000_5192000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M4530 diff_2335000_1372000# diff_2335000_1372000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4531 diff_95000_5192000# diff_2335000_1127000# diff_2335000_1127000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=-2.02697e+09 ps=426000 
M4532 diff_2130000_1289000# diff_2130000_1289000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4533 diff_95000_5192000# diff_2130000_1219000# diff_2130000_1219000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=1.377e+09 ps=310000 
M4534 diff_2335000_1127000# diff_1094000_1020000# diff_2406000_1192000# GND efet w=151500 l=9500
+ ad=0 pd=0 as=1.527e+09 ps=304000 
M4535 diff_2406000_1192000# diff_2130000_1219000# diff_83000_3098000# GND efet w=120000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4536 diff_83000_3098000# diff_2335000_1127000# diff_2290000_1091000# GND efet w=60000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4537 diff_2460000_1079000# diff_1037000_877000# diff_2335000_1127000# GND efet w=150500 l=8500
+ ad=1.671e+09 pd=328000 as=0 ps=0 
M4538 diff_817000_1286000# diff_1438000_786000# diff_95000_5192000# GND efet w=88500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4539 diff_2650000_1323000# diff_2641000_934000# diff_817000_1286000# GND efet w=21000 l=9000
+ ad=5.56e+08 pd=180000 as=0 ps=0 
M4540 diff_817000_1286000# diff_2775000_765000# diff_2683000_1400000# GND efet w=107500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4541 diff_83000_3098000# diff_2876000_1451000# diff_2829000_1488000# GND efet w=214500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4542 diff_2876000_1451000# diff_2915000_1565000# diff_83000_3098000# GND efet w=61500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4543 diff_817000_1211000# diff_1438000_786000# diff_95000_5192000# GND efet w=88500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4544 diff_83000_3098000# diff_2471000_1074000# diff_2460000_1079000# GND efet w=123500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4545 diff_2130000_1219000# diff_2471000_1074000# diff_83000_3098000# GND efet w=58000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4546 diff_95000_5192000# diff_2531000_1102000# diff_2531000_1102000# GND efet w=11000 l=16000
+ ad=0 pd=0 as=1.627e+09 ps=342000 
M4547 diff_2674000_1391000# diff_95000_5192000# diff_95000_5192000# GND efet w=11000 l=31000
+ ad=0 pd=0 as=0 ps=0 
M4548 diff_2683000_1400000# diff_95000_5192000# diff_2650000_1323000# GND efet w=12500 l=81500
+ ad=0 pd=0 as=0 ps=0 
M4549 diff_2683000_1400000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4550 diff_95000_5192000# diff_95000_5192000# diff_2674000_1077000# GND efet w=11000 l=31000
+ ad=0 pd=0 as=9.05e+08 ps=196000 
M4551 diff_2683000_1084000# diff_95000_5192000# diff_2651000_1168000# GND efet w=12000 l=74000
+ ad=-1.98967e+08 pd=736000 as=5.3e+08 ps=188000 
M4552 diff_95000_5192000# diff_95000_5192000# diff_2683000_1084000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4553 diff_2651000_1168000# diff_2641000_934000# diff_817000_1211000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4554 diff_83000_3098000# diff_1851000_1079000# diff_2531000_1102000# GND efet w=82500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4555 diff_2531000_1102000# diff_2448000_2717000# diff_2471000_1074000# GND efet w=21000 l=12000
+ ad=0 pd=0 as=3.35e+08 ps=80000 
M4556 diff_83000_3098000# diff_2409000_958000# diff_2130000_913000# GND efet w=64000 l=8000
+ ad=0 pd=0 as=1.616e+09 ps=356000 
M4557 diff_95000_5192000# diff_1438000_786000# diff_1851000_1079000# GND efet w=85500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4558 diff_848000_1211000# diff_1438000_786000# diff_95000_5192000# GND efet w=71000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4559 diff_2674000_1077000# diff_2651000_1168000# diff_83000_3098000# GND efet w=61000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4560 diff_2829000_1316000# diff_2583000_2725000# diff_817000_1286000# GND efet w=86000 l=10000
+ ad=-1.64967e+08 pd=722000 as=0 ps=0 
M4561 diff_2829000_1316000# diff_2843000_1950000# diff_848000_1262000# GND efet w=105500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4562 diff_83000_3098000# diff_2876000_1416000# diff_2829000_1316000# GND efet w=212500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4563 diff_2876000_1416000# diff_2914000_1304000# diff_83000_3098000# GND efet w=67500 l=7500
+ ad=8.92e+08 pd=182000 as=0 ps=0 
M4564 diff_83000_3098000# diff_2534000_2492000# diff_1774000_760000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4565 diff_3099000_1943000# diff_3029000_1923000# diff_83000_3098000# GND efet w=60500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4566 diff_3117000_1841000# diff_3099000_1943000# diff_83000_3098000# GND efet w=211500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4567 diff_1774000_760000# diff_3120000_2492000# diff_3117000_1841000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4568 diff_817000_1965000# diff_2893000_2725000# diff_3117000_1841000# GND efet w=87000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4569 diff_83000_3098000# diff_2534000_2492000# diff_1791000_798000# GND efet w=107000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4570 diff_3117000_1777000# diff_3099000_1681000# diff_83000_3098000# GND efet w=212500 l=7500
+ ad=-4.05967e+08 pd=686000 as=0 ps=0 
M4571 diff_3099000_1681000# diff_3029000_1664000# diff_83000_3098000# GND efet w=67500 l=8500
+ ad=9.44e+08 pd=198000 as=0 ps=0 
M4572 diff_817000_1663000# diff_2638000_2492000# diff_3029000_1664000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4573 diff_817000_1588000# diff_2638000_2492000# diff_3029000_1546000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=1.624e+09 ps=392000 
M4574 diff_1791000_798000# diff_3120000_2492000# diff_3117000_1777000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4575 diff_817000_1663000# diff_2893000_2725000# diff_3117000_1777000# GND efet w=86000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4576 diff_3099000_1681000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=31000
+ ad=0 pd=0 as=0 ps=0 
M4577 diff_3117000_1777000# diff_95000_5192000# diff_3029000_1664000# GND efet w=12000 l=81000
+ ad=0 pd=0 as=0 ps=0 
M4578 diff_3117000_1777000# diff_95000_5192000# diff_95000_5192000# GND efet w=11000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4579 diff_95000_5192000# diff_95000_5192000# diff_3099000_1566000# GND efet w=12000 l=30000
+ ad=0 pd=0 as=9.78e+08 ps=200000 
M4580 diff_3117000_1464000# diff_95000_5192000# diff_3029000_1546000# GND efet w=12000 l=72000
+ ad=-3.27967e+08 pd=708000 as=0 ps=0 
M4581 diff_95000_5192000# diff_95000_5192000# diff_3117000_1464000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4582 diff_848000_1588000# diff_2996000_2725000# diff_2915000_1565000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4583 diff_3029000_1546000# diff_2996000_2725000# diff_1851000_1456000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4584 diff_3029000_1287000# diff_2996000_2725000# diff_1851000_1376000# GND efet w=19000 l=10000
+ ad=1.547e+09 pd=370000 as=0 ps=0 
M4585 diff_848000_1262000# diff_2996000_2725000# diff_2914000_1304000# GND efet w=19000 l=10000
+ ad=0 pd=0 as=1.205e+09 ps=308000 
M4586 diff_2829000_1316000# diff_95000_5192000# diff_95000_5192000# GND efet w=11000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4587 diff_2914000_1304000# diff_95000_5192000# diff_2829000_1316000# GND efet w=12500 l=80500
+ ad=0 pd=0 as=0 ps=0 
M4588 diff_2876000_1416000# diff_95000_5192000# diff_95000_5192000# GND efet w=11000 l=31000
+ ad=0 pd=0 as=0 ps=0 
M4589 diff_2914000_1304000# diff_2939000_824000# diff_817000_1286000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4590 diff_95000_5192000# diff_95000_5192000# diff_2829000_1111000# GND efet w=11000 l=22000
+ ad=0 pd=0 as=-5.79673e+07 ps=732000 
M4591 diff_2915000_1188000# diff_95000_5192000# diff_2829000_1111000# GND efet w=12000 l=74000
+ ad=1.204e+09 pd=306000 as=0 ps=0 
M4592 diff_95000_5192000# diff_95000_5192000# diff_2876000_1074000# GND efet w=12000 l=30000
+ ad=0 pd=0 as=8.62e+08 ps=188000 
M4593 diff_817000_1211000# diff_2775000_765000# diff_2683000_1084000# GND efet w=108500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4594 diff_2683000_1084000# diff_2674000_1077000# diff_83000_3098000# GND efet w=218500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4595 diff_1851000_1079000# diff_2713000_822000# diff_2683000_1084000# GND efet w=102000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4596 diff_83000_3098000# diff_1851000_999000# diff_2531000_969000# GND efet w=80000 l=8000
+ ad=0 pd=0 as=1.711e+09 ps=340000 
M4597 diff_95000_5192000# diff_1438000_786000# diff_1851000_999000# GND efet w=86500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4598 diff_2127000_952000# diff_1237000_1921000# diff_95000_5192000# GND efet w=12000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4599 diff_2184000_926000# diff_2184000_926000# diff_95000_5192000# GND efet w=12000 l=19000
+ ad=0 pd=0 as=0 ps=0 
M4600 diff_2102000_884000# diff_1438000_786000# diff_2050000_1017000# GND efet w=20000 l=12000
+ ad=1.4e+08 pd=54000 as=4.06e+08 ps=92000 
M4601 diff_2121000_884000# diff_72000_4515000# diff_2102000_884000# GND efet w=20000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M4602 diff_95000_5192000# diff_2121000_884000# diff_2121000_884000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M4603 diff_83000_3098000# diff_72000_4515000# diff_1837000_1364000# GND efet w=70000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4604 diff_1858000_1019000# diff_72000_4515000# diff_83000_3098000# GND efet w=70000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4605 diff_83000_3098000# diff_72000_4515000# diff_1547000_932000# GND efet w=72000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4606 diff_1487000_841000# diff_72000_4515000# diff_83000_3098000# GND efet w=79500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4607 diff_83000_3098000# diff_1386000_841000# diff_1438000_786000# GND efet w=72000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4608 diff_1237000_1921000# diff_72000_4515000# diff_83000_3098000# GND efet w=72000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4609 diff_2531000_969000# diff_2448000_2717000# diff_2409000_958000# GND efet w=22000 l=12000
+ ad=0 pd=0 as=3.94e+08 ps=80000 
M4610 diff_848000_885000# diff_1438000_786000# diff_95000_5192000# GND efet w=72000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4611 diff_2829000_1111000# diff_2583000_2725000# diff_817000_1211000# GND efet w=86000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4612 diff_2915000_1188000# diff_2939000_824000# diff_817000_1211000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4613 diff_2915000_1188000# diff_2915000_1188000# diff_2915000_1188000# GND efet w=500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4614 diff_2829000_1111000# diff_2843000_1950000# diff_848000_1211000# GND efet w=106500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4615 diff_2683000_1022000# diff_2674000_1013000# diff_83000_3098000# GND efet w=218500 l=8500
+ ad=-2.13967e+08 pd=722000 as=0 ps=0 
M4616 diff_95000_5192000# diff_2130000_913000# diff_2130000_913000# GND efet w=14000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4617 diff_1386000_841000# diff_72000_4515000# diff_83000_3098000# GND efet w=102000 l=8000
+ ad=-2.02597e+09 pd=322000 as=0 ps=0 
M4618 diff_95000_5192000# diff_1386000_841000# diff_1386000_841000# GND efet w=14000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M4619 diff_2448000_2717000# diff_72000_4515000# diff_83000_3098000# GND efet w=72000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4620 diff_2674000_1013000# diff_2650000_947000# diff_83000_3098000# GND efet w=68000 l=8000
+ ad=9.11e+08 pd=194000 as=0 ps=0 
M4621 diff_1851000_999000# diff_2713000_822000# diff_2683000_1022000# GND efet w=103500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4622 diff_2531000_969000# diff_2531000_969000# diff_95000_5192000# GND efet w=13000 l=16000
+ ad=0 pd=0 as=0 ps=0 
M4623 diff_817000_909000# diff_1438000_786000# diff_95000_5192000# GND efet w=87500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4624 diff_2650000_947000# diff_2641000_934000# diff_817000_909000# GND efet w=20000 l=9000
+ ad=5.32e+08 pd=176000 as=0 ps=0 
M4625 diff_817000_909000# diff_2775000_765000# diff_2683000_1022000# GND efet w=108000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4626 diff_83000_3098000# diff_2876000_1074000# diff_2829000_1111000# GND efet w=213500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4627 diff_2876000_1074000# diff_2915000_1188000# diff_83000_3098000# GND efet w=61500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4628 diff_2674000_1013000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=32000
+ ad=0 pd=0 as=0 ps=0 
M4629 diff_2683000_1022000# diff_95000_5192000# diff_2650000_947000# GND efet w=12500 l=80500
+ ad=0 pd=0 as=0 ps=0 
M4630 diff_2683000_1022000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4631 diff_2829000_939000# diff_2583000_2725000# diff_817000_909000# GND efet w=86000 l=11000
+ ad=-1.57967e+08 pd=722000 as=0 ps=0 
M4632 diff_2829000_939000# diff_2843000_1950000# diff_848000_885000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4633 diff_83000_3098000# diff_2876000_1039000# diff_2829000_939000# GND efet w=212500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4634 diff_2876000_1039000# diff_2915000_927000# diff_83000_3098000# GND efet w=66500 l=7500
+ ad=8.91e+08 pd=182000 as=0 ps=0 
M4635 diff_1438000_786000# diff_1386000_841000# diff_83000_3098000# GND efet w=72000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4636 diff_83000_3098000# diff_72000_4515000# diff_2641000_934000# GND efet w=71000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4637 diff_83000_3098000# diff_2534000_2492000# diff_1851000_1456000# GND efet w=107000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4638 diff_3099000_1566000# diff_3029000_1546000# diff_83000_3098000# GND efet w=61500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4639 diff_3489000_2725000# diff_72000_4515000# diff_83000_3098000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4640 diff_83000_3098000# diff_3486000_2778000# diff_3489000_2725000# GND efet w=244500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4641 diff_3474000_792000# diff_3536000_2778000# diff_83000_3098000# GND efet w=244500 l=8500
+ ad=1.28103e+09 pd=974000 as=0 ps=0 
M4642 diff_95000_5192000# diff_3474000_792000# diff_3474000_792000# GND efet w=18000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M4643 diff_3567000_785000# diff_3567000_785000# diff_95000_5192000# GND efet w=18000 l=7000
+ ad=4.27033e+08 pd=936000 as=0 ps=0 
M4644 diff_83000_3098000# diff_72000_4515000# diff_3474000_792000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4645 diff_3567000_785000# diff_72000_4515000# diff_83000_3098000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4646 diff_83000_3098000# diff_3589000_2778000# diff_3567000_785000# GND efet w=245000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4647 diff_3596000_2395000# diff_3639000_2778000# diff_83000_3098000# GND efet w=244500 l=8500
+ ad=6.30033e+08 pd=858000 as=0 ps=0 
M4648 diff_95000_5192000# diff_3596000_2395000# diff_3596000_2395000# GND efet w=18000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4649 diff_3695000_2725000# diff_3695000_2725000# diff_95000_5192000# GND efet w=18000 l=8000
+ ad=1.00603e+09 pd=978000 as=0 ps=0 
M4650 diff_83000_3098000# diff_72000_4515000# diff_3596000_2395000# GND efet w=203000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4651 diff_3695000_2725000# diff_72000_4515000# diff_83000_3098000# GND efet w=203000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4652 diff_83000_3098000# diff_3692000_2778000# diff_3695000_2725000# GND efet w=244500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4653 diff_3749000_2434000# diff_3742000_2778000# diff_83000_3098000# GND efet w=245000 l=9000
+ ad=3.10327e+07 pd=858000 as=0 ps=0 
M4654 diff_95000_5192000# diff_3749000_2434000# diff_3749000_2434000# GND efet w=18000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4655 diff_3739000_826000# diff_3739000_826000# diff_95000_5192000# GND efet w=18000 l=8000
+ ad=8.17033e+08 pd=918000 as=0 ps=0 
M4656 diff_83000_3098000# diff_72000_4515000# diff_3749000_2434000# GND efet w=204000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4657 diff_3739000_826000# diff_72000_4515000# diff_83000_3098000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4658 diff_83000_3098000# diff_3794000_2778000# diff_3739000_826000# GND efet w=244000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4659 diff_3830000_787000# diff_3846000_2778000# diff_83000_3098000# GND efet w=244500 l=8500
+ ad=7.37033e+08 pd=922000 as=0 ps=0 
M4660 diff_95000_5192000# diff_3830000_787000# diff_3830000_787000# GND efet w=18000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4661 diff_3901000_2725000# diff_3901000_2725000# diff_95000_5192000# GND efet w=18000 l=8000
+ ad=3.02033e+08 pd=876000 as=0 ps=0 
M4662 diff_83000_3098000# diff_72000_4515000# diff_3830000_787000# GND efet w=204000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4663 diff_3901000_2725000# diff_72000_4515000# diff_83000_3098000# GND efet w=204000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4664 diff_83000_3098000# diff_3898000_2778000# diff_3901000_2725000# GND efet w=244000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4665 diff_3922000_786000# diff_3949000_2778000# diff_83000_3098000# GND efet w=244500 l=8500
+ ad=7.41033e+08 pd=940000 as=0 ps=0 
M4666 diff_95000_5192000# diff_3922000_786000# diff_3922000_786000# GND efet w=18000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4667 diff_4004000_2725000# diff_4004000_2725000# diff_95000_5192000# GND efet w=18000 l=8000
+ ad=8.78033e+08 pd=878000 as=0 ps=0 
M4668 diff_83000_3098000# diff_72000_4515000# diff_3922000_786000# GND efet w=203000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4669 diff_4004000_2725000# diff_72000_4515000# diff_83000_3098000# GND efet w=203000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4670 diff_83000_3098000# diff_4001000_2778000# diff_4004000_2725000# GND efet w=244500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4671 diff_3117000_1464000# diff_3099000_1566000# diff_83000_3098000# GND efet w=212500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4672 diff_1851000_1456000# diff_3120000_2492000# diff_3117000_1464000# GND efet w=85000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4673 diff_817000_1588000# diff_2893000_2725000# diff_3117000_1464000# GND efet w=87000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4674 diff_83000_3098000# diff_3256000_1459000# diff_817000_1588000# GND efet w=91000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4675 diff_95000_5192000# diff_95000_5192000# diff_95000_5192000# GND efet w=500 l=4500
+ ad=0 pd=0 as=0 ps=0 
M4676 diff_95000_5192000# diff_95000_5192000# diff_1399000_598000# GND efet w=12000 l=104000
+ ad=0 pd=0 as=0 ps=0 
M4677 diff_95000_5192000# diff_95000_5192000# diff_3427000_2321000# GND efet w=12000 l=32000
+ ad=0 pd=0 as=9.5e+08 ps=192000 
M4678 diff_3436000_2231000# diff_95000_5192000# diff_3374000_2284000# GND efet w=12000 l=74000
+ ad=-2.59673e+07 pd=728000 as=1.504e+09 ps=368000 
M4679 diff_95000_5192000# diff_95000_5192000# diff_3436000_2231000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4680 diff_817000_2342000# diff_3171000_2725000# diff_3374000_2284000# GND efet w=19000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4681 diff_3436000_2231000# diff_3439000_2492000# diff_817000_2342000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4682 diff_3577000_2265000# diff_3567000_785000# diff_3436000_2231000# GND efet w=109000 l=10000
+ ad=-2.13193e+09 pd=1.356e+06 as=0 ps=0 
M4683 diff_3374000_2284000# diff_3354000_2409000# diff_1399000_598000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4684 diff_3374000_2060000# diff_3354000_2409000# diff_1757000_739000# GND efet w=20000 l=10000
+ ad=1.521e+09 pd=382000 as=0 ps=0 
M4685 diff_1757000_739000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=102000
+ ad=0 pd=0 as=0 ps=0 
M4686 diff_3427000_2321000# diff_3374000_2284000# diff_83000_3098000# GND efet w=66000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4687 diff_3436000_2231000# diff_3427000_2321000# diff_83000_3098000# GND efet w=204500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4688 diff_1399000_598000# diff_3474000_792000# diff_3436000_2231000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4689 diff_3436000_2160000# diff_3428000_2064000# diff_83000_3098000# GND efet w=205500 l=7500
+ ad=-5.49673e+07 pd=720000 as=0 ps=0 
M4690 diff_3428000_2064000# diff_3374000_2060000# diff_83000_3098000# GND efet w=72000 l=8000
+ ad=9.43e+08 pd=192000 as=0 ps=0 
M4691 diff_1757000_739000# diff_3474000_792000# diff_3436000_2160000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4692 diff_848000_2342000# diff_3596000_2395000# diff_3577000_2265000# GND efet w=119000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4693 diff_3800000_830000# diff_4052000_2778000# diff_83000_3098000# GND efet w=244500 l=8500
+ ad=9.01033e+08 pd=924000 as=0 ps=0 
M4694 diff_95000_5192000# diff_3800000_830000# diff_3800000_830000# GND efet w=18000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4695 diff_4108000_2725000# diff_4108000_2725000# diff_95000_5192000# GND efet w=18000 l=8000
+ ad=2.61033e+08 pd=882000 as=0 ps=0 
M4696 diff_83000_3098000# diff_72000_4515000# diff_3800000_830000# GND efet w=203000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4697 diff_4108000_2725000# diff_72000_4515000# diff_83000_3098000# GND efet w=203000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4698 diff_83000_3098000# diff_4104000_2778000# diff_4108000_2725000# GND efet w=245500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4699 diff_4224000_2739000# diff_4224000_2739000# diff_95000_5192000# GND efet w=12000 l=14000
+ ad=3.93033e+08 pd=866000 as=0 ps=0 
M4700 diff_4277000_2781000# diff_4277000_2781000# diff_95000_5192000# GND efet w=14000 l=13000
+ ad=-7.27967e+08 pd=820000 as=0 ps=0 
M4701 diff_95000_5192000# diff_4363000_2478000# diff_4363000_2478000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4702 diff_83000_3098000# diff_4241000_2640000# diff_4224000_2739000# GND efet w=128500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4703 diff_95000_5192000# diff_4155000_2676000# diff_4155000_2676000# GND efet w=13000 l=16000
+ ad=0 pd=0 as=-8.37967e+08 ps=640000 
M4704 diff_4155000_2676000# diff_3043000_2723000# diff_83000_3098000# GND efet w=100000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M4705 diff_83000_3098000# diff_4182000_2528000# diff_4155000_2676000# GND efet w=117500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4706 diff_817000_2342000# diff_3489000_2725000# diff_3632000_2301000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=9.81e+08 ps=234000 
M4707 diff_95000_5192000# diff_95000_5192000# diff_3686000_2317000# GND efet w=13000 l=32000
+ ad=0 pd=0 as=1.066e+09 ps=202000 
M4708 diff_3696000_2230000# diff_95000_5192000# diff_3632000_2301000# GND efet w=12000 l=72000
+ ad=-2.80967e+08 pd=722000 as=0 ps=0 
M4709 diff_95000_5192000# diff_95000_5192000# diff_3696000_2230000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4710 diff_3632000_2301000# diff_3354000_2409000# diff_848000_2342000# GND efet w=19000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4711 diff_817000_2040000# diff_3171000_2725000# diff_3374000_2060000# GND efet w=19000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4712 diff_95000_5192000# diff_95000_5192000# diff_1774000_760000# GND efet w=12000 l=104000
+ ad=0 pd=0 as=0 ps=0 
M4713 diff_3428000_2064000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=32000
+ ad=0 pd=0 as=0 ps=0 
M4714 diff_3436000_2160000# diff_95000_5192000# diff_3374000_2060000# GND efet w=12500 l=79500
+ ad=0 pd=0 as=0 ps=0 
M4715 diff_3436000_2160000# diff_95000_5192000# diff_95000_5192000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4716 diff_95000_5192000# diff_95000_5192000# diff_3427000_1944000# GND efet w=12000 l=32000
+ ad=0 pd=0 as=9.45e+08 ps=192000 
M4717 diff_3436000_1854000# diff_95000_5192000# diff_3374000_1907000# GND efet w=12000 l=72000
+ ad=-6.19673e+07 pd=726000 as=1.503e+09 ps=368000 
M4718 diff_95000_5192000# diff_95000_5192000# diff_3436000_1854000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4719 diff_817000_1965000# diff_3171000_2725000# diff_3374000_1907000# GND efet w=19000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4720 diff_3436000_2160000# diff_3439000_2492000# diff_817000_2040000# GND efet w=105500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4721 diff_3577000_2123000# diff_3567000_785000# diff_3436000_2160000# GND efet w=109000 l=10000
+ ad=2.08703e+09 pd=1.35e+06 as=0 ps=0 
M4722 diff_848000_2016000# diff_3596000_2395000# diff_3577000_2123000# GND efet w=120000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4723 diff_3632000_2078000# diff_3354000_2409000# diff_848000_2016000# GND efet w=19000 l=11000
+ ad=9.89e+08 pd=240000 as=0 ps=0 
M4724 diff_3436000_1854000# diff_3439000_2492000# diff_817000_1965000# GND efet w=105500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4725 diff_3577000_1888000# diff_3567000_785000# diff_3436000_1854000# GND efet w=109000 l=10000
+ ad=2.14103e+09 pd=1.36e+06 as=0 ps=0 
M4726 diff_3374000_1907000# diff_3354000_2409000# diff_1774000_760000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4727 diff_3374000_1683000# diff_3354000_2409000# diff_1791000_798000# GND efet w=20000 l=10000
+ ad=1.539e+09 pd=384000 as=0 ps=0 
M4728 diff_1791000_798000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=102000
+ ad=0 pd=0 as=0 ps=0 
M4729 diff_3427000_1944000# diff_3374000_1907000# diff_83000_3098000# GND efet w=66000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4730 diff_3436000_1854000# diff_3427000_1944000# diff_83000_3098000# GND efet w=204500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4731 diff_1774000_760000# diff_3474000_792000# diff_3436000_1854000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4732 diff_3436000_1783000# diff_3428000_1687000# diff_83000_3098000# GND efet w=205500 l=7500
+ ad=-1.78967e+08 pd=718000 as=0 ps=0 
M4733 diff_3428000_1687000# diff_3374000_1683000# diff_83000_3098000# GND efet w=72000 l=8000
+ ad=9.55e+08 pd=194000 as=0 ps=0 
M4734 diff_1791000_798000# diff_3474000_792000# diff_3436000_1783000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4735 diff_848000_1965000# diff_3596000_2395000# diff_3577000_1888000# GND efet w=120000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4736 diff_817000_2342000# diff_3800000_830000# diff_3696000_2230000# GND efet w=102000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4737 diff_3846000_2258000# diff_3830000_787000# diff_817000_2342000# GND efet w=102000 l=10000
+ ad=-1.59967e+08 pd=720000 as=0 ps=0 
M4738 diff_3686000_2317000# diff_3632000_2301000# diff_83000_3098000# GND efet w=65500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4739 diff_3696000_2230000# diff_3686000_2317000# diff_83000_3098000# GND efet w=202000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4740 diff_3577000_2265000# diff_3739000_826000# diff_3696000_2230000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4741 diff_95000_5192000# diff_95000_5192000# diff_3846000_2258000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4742 diff_3938000_2317000# diff_95000_5192000# diff_3846000_2258000# GND efet w=12000 l=72000
+ ad=7.83e+08 pd=254000 as=0 ps=0 
M4743 diff_95000_5192000# diff_95000_5192000# diff_3902000_2206000# GND efet w=13000 l=32000
+ ad=0 pd=0 as=1.038e+09 ps=194000 
M4744 diff_83000_3098000# diff_4303000_2657000# diff_4277000_2781000# GND efet w=103000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4745 diff_83000_3098000# diff_3043000_2723000# diff_4224000_2739000# GND efet w=115000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4746 diff_83000_3098000# diff_3043000_2723000# diff_4277000_2781000# GND efet w=123500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4747 diff_3696000_2160000# diff_3687000_2066000# diff_83000_3098000# GND efet w=203000 l=8000
+ ad=-4.18967e+08 pd=712000 as=0 ps=0 
M4748 diff_3687000_2066000# diff_3632000_2078000# diff_83000_3098000# GND efet w=70500 l=8500
+ ad=1.014e+09 pd=200000 as=0 ps=0 
M4749 diff_3577000_2123000# diff_3739000_826000# diff_3696000_2160000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4750 diff_3846000_2258000# diff_3695000_2725000# diff_3577000_2265000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4751 diff_817000_2342000# diff_3922000_786000# diff_3938000_2317000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4752 diff_4037000_2327000# diff_4004000_2725000# diff_817000_2342000# GND efet w=20000 l=11000
+ ad=8.53e+08 pd=258000 as=0 ps=0 
M4753 diff_95000_5192000# diff_95000_5192000# diff_4057000_2222000# GND efet w=13000 l=32000
+ ad=0 pd=0 as=9.82e+08 ps=190000 
M4754 diff_4066000_2230000# diff_95000_5192000# diff_4037000_2327000# GND efet w=12500 l=72500
+ ad=-3.55967e+08 pd=696000 as=0 ps=0 
M4755 diff_95000_5192000# diff_95000_5192000# diff_4066000_2230000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4756 diff_83000_3098000# diff_3902000_2206000# diff_3846000_2258000# GND efet w=203000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4757 diff_3902000_2206000# diff_3938000_2317000# diff_83000_3098000# GND efet w=61500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4758 diff_817000_2040000# diff_3489000_2725000# diff_3632000_2078000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4759 diff_3687000_2066000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=32000
+ ad=0 pd=0 as=0 ps=0 
M4760 diff_3696000_2160000# diff_95000_5192000# diff_3632000_2078000# GND efet w=12500 l=79500
+ ad=0 pd=0 as=0 ps=0 
M4761 diff_3696000_2160000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4762 diff_817000_1965000# diff_3489000_2725000# diff_3632000_1923000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=9.94e+08 ps=234000 
M4763 diff_95000_5192000# diff_95000_5192000# diff_3686000_1940000# GND efet w=13000 l=32000
+ ad=0 pd=0 as=1.075e+09 ps=202000 
M4764 diff_3696000_1853000# diff_95000_5192000# diff_3632000_1923000# GND efet w=12000 l=73000
+ ad=-2.19967e+08 pd=722000 as=0 ps=0 
M4765 diff_95000_5192000# diff_95000_5192000# diff_3696000_1853000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4766 diff_3632000_1923000# diff_3354000_2409000# diff_848000_1965000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4767 diff_817000_1663000# diff_3171000_2725000# diff_3374000_1683000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4768 diff_83000_3098000# diff_2534000_2492000# diff_1851000_1376000# GND efet w=107000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4769 diff_3117000_1400000# diff_3099000_1304000# diff_83000_3098000# GND efet w=210500 l=7500
+ ad=-4.23967e+08 pd=688000 as=0 ps=0 
M4770 diff_3099000_1304000# diff_3029000_1287000# diff_83000_3098000# GND efet w=67500 l=8500
+ ad=9.43e+08 pd=198000 as=0 ps=0 
M4771 diff_817000_1286000# diff_2638000_2492000# diff_3029000_1287000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4772 diff_817000_1211000# diff_2638000_2492000# diff_3029000_1168000# GND efet w=21000 l=9000
+ ad=0 pd=0 as=1.611e+09 ps=390000 
M4773 diff_1851000_1376000# diff_3120000_2492000# diff_3117000_1400000# GND efet w=85000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4774 diff_817000_1286000# diff_3283000_1426000# diff_83000_3098000# GND efet w=89000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4775 diff_95000_5192000# diff_95000_5192000# diff_1851000_1456000# GND efet w=12000 l=104000
+ ad=0 pd=0 as=0 ps=0 
M4776 diff_3428000_1687000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=32000
+ ad=0 pd=0 as=0 ps=0 
M4777 diff_3436000_1783000# diff_95000_5192000# diff_3374000_1683000# GND efet w=12500 l=78500
+ ad=0 pd=0 as=0 ps=0 
M4778 diff_3436000_1783000# diff_95000_5192000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4779 diff_95000_5192000# diff_95000_5192000# diff_3427000_1566000# GND efet w=12000 l=32000
+ ad=0 pd=0 as=9.27e+08 ps=190000 
M4780 diff_3436000_1476000# diff_95000_5192000# diff_3374000_1530000# GND efet w=12000 l=74000
+ ad=-1.26967e+08 pd=724000 as=1.51e+09 ps=368000 
M4781 diff_95000_5192000# diff_95000_5192000# diff_3436000_1476000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4782 diff_817000_1588000# diff_3171000_2725000# diff_3374000_1530000# GND efet w=19000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4783 diff_3436000_1783000# diff_3439000_2492000# diff_817000_1663000# GND efet w=105000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4784 diff_3577000_1746000# diff_3567000_785000# diff_3436000_1783000# GND efet w=108000 l=10000
+ ad=-2.11093e+09 pd=1.354e+06 as=0 ps=0 
M4785 diff_848000_1639000# diff_3596000_2395000# diff_3577000_1746000# GND efet w=120000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4786 diff_3632000_1701000# diff_3354000_2409000# diff_848000_1639000# GND efet w=19000 l=10000
+ ad=1.015e+09 pd=244000 as=0 ps=0 
M4787 diff_3436000_1476000# diff_3439000_2492000# diff_817000_1588000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4788 diff_3577000_1511000# diff_3567000_785000# diff_3436000_1476000# GND efet w=109000 l=10000
+ ad=2.13503e+09 pd=1.34e+06 as=0 ps=0 
M4789 diff_817000_1286000# diff_2893000_2725000# diff_3117000_1400000# GND efet w=86000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4790 diff_3099000_1304000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=31000
+ ad=0 pd=0 as=0 ps=0 
M4791 diff_3117000_1400000# diff_95000_5192000# diff_3029000_1287000# GND efet w=12000 l=79000
+ ad=0 pd=0 as=0 ps=0 
M4792 diff_3117000_1400000# diff_95000_5192000# diff_95000_5192000# GND efet w=11000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4793 diff_95000_5192000# diff_95000_5192000# diff_3099000_1189000# GND efet w=12000 l=30000
+ ad=0 pd=0 as=9.85e+08 ps=200000 
M4794 diff_3117000_1087000# diff_95000_5192000# diff_3029000_1168000# GND efet w=12000 l=74000
+ ad=-2.66967e+08 pd=704000 as=0 ps=0 
M4795 diff_95000_5192000# diff_95000_5192000# diff_3117000_1087000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4796 diff_848000_1211000# diff_2996000_2725000# diff_2915000_1188000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M4797 diff_3029000_1168000# diff_2996000_2725000# diff_1851000_1079000# GND efet w=19000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4798 diff_3029000_910000# diff_2996000_2725000# diff_1851000_999000# GND efet w=19000 l=10000
+ ad=1.59e+09 pd=378000 as=0 ps=0 
M4799 diff_848000_885000# diff_2996000_2725000# diff_2915000_927000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=1.21e+09 ps=302000 
M4800 diff_2829000_939000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4801 diff_2915000_927000# diff_95000_5192000# diff_2829000_939000# GND efet w=12500 l=81500
+ ad=0 pd=0 as=0 ps=0 
M4802 diff_2876000_1039000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=31000
+ ad=0 pd=0 as=0 ps=0 
M4803 diff_2915000_927000# diff_2939000_824000# diff_817000_909000# GND efet w=19000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4804 diff_83000_3098000# diff_2534000_2492000# diff_1851000_1079000# GND efet w=106500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4805 diff_3099000_1189000# diff_3029000_1168000# diff_83000_3098000# GND efet w=62500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4806 diff_3374000_1530000# diff_3354000_2409000# diff_1851000_1456000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4807 diff_3374000_1306000# diff_3354000_2409000# diff_1851000_1376000# GND efet w=20000 l=10000
+ ad=1.526e+09 pd=382000 as=0 ps=0 
M4808 diff_1851000_1376000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=102000
+ ad=0 pd=0 as=0 ps=0 
M4809 diff_3427000_1566000# diff_3374000_1530000# diff_83000_3098000# GND efet w=65000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4810 diff_3436000_1476000# diff_3427000_1566000# diff_83000_3098000# GND efet w=203500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4811 diff_1851000_1456000# diff_3474000_792000# diff_3436000_1476000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4812 diff_3436000_1405000# diff_3428000_1309000# diff_83000_3098000# GND efet w=204500 l=7500
+ ad=-1.29967e+08 pd=716000 as=0 ps=0 
M4813 diff_3428000_1309000# diff_3374000_1306000# diff_83000_3098000# GND efet w=70000 l=8000
+ ad=9.3e+08 pd=192000 as=0 ps=0 
M4814 diff_1851000_1376000# diff_3474000_792000# diff_3436000_1405000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4815 diff_848000_1588000# diff_3596000_2395000# diff_3577000_1511000# GND efet w=120000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4816 diff_817000_2040000# diff_3800000_830000# diff_3696000_2160000# GND efet w=102000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4817 diff_3846000_2078000# diff_3830000_787000# diff_817000_2040000# GND efet w=102500 l=9500
+ ad=-1.86967e+08 pd=716000 as=0 ps=0 
M4818 diff_3846000_2078000# diff_3695000_2725000# diff_3577000_2123000# GND efet w=85000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4819 diff_83000_3098000# diff_3902000_2172000# diff_3846000_2078000# GND efet w=204000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4820 diff_3902000_2172000# diff_3939000_2058000# diff_83000_3098000# GND efet w=63000 l=8000
+ ad=1.034e+09 pd=192000 as=0 ps=0 
M4821 diff_817000_1965000# diff_3800000_830000# diff_3696000_1853000# GND efet w=102500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4822 diff_3846000_1881000# diff_3830000_787000# diff_817000_1965000# GND efet w=102500 l=9500
+ ad=-1.28967e+08 pd=720000 as=0 ps=0 
M4823 diff_3686000_1940000# diff_3632000_1923000# diff_83000_3098000# GND efet w=66500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4824 diff_3696000_1853000# diff_3686000_1940000# diff_83000_3098000# GND efet w=203000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4825 diff_3577000_1888000# diff_3739000_826000# diff_3696000_1853000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4826 diff_4057000_2222000# diff_4037000_2327000# diff_83000_3098000# GND efet w=59500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4827 diff_4066000_2230000# diff_4057000_2222000# diff_83000_3098000# GND efet w=202500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4828 diff_817000_2342000# diff_4108000_2725000# diff_4066000_2230000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4829 diff_3577000_2265000# diff_3749000_2434000# diff_4066000_2230000# GND efet w=85000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4830 diff_4066000_2160000# diff_4057000_2151000# diff_83000_3098000# GND efet w=204500 l=7500
+ ad=-3.80967e+08 pd=692000 as=0 ps=0 
M4831 diff_83000_3098000# diff_4036000_2051000# diff_4057000_2151000# GND efet w=60500 l=8500
+ ad=0 pd=0 as=9.37e+08 ps=184000 
M4832 diff_817000_2040000# diff_4108000_2725000# diff_4066000_2160000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4833 diff_83000_3098000# diff_3901000_2725000# diff_3577000_2265000# GND efet w=106000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4834 diff_83000_3098000# diff_3901000_2725000# diff_3577000_2123000# GND efet w=104000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4835 diff_817000_2040000# diff_4155000_2676000# diff_83000_3098000# GND efet w=89000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4836 diff_3846000_2078000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4837 diff_3939000_2058000# diff_95000_5192000# diff_3846000_2078000# GND efet w=12500 l=78500
+ ad=8.17e+08 pd=232000 as=0 ps=0 
M4838 diff_3902000_2172000# diff_95000_5192000# diff_95000_5192000# GND efet w=13000 l=32000
+ ad=0 pd=0 as=0 ps=0 
M4839 diff_817000_2040000# diff_3922000_786000# diff_3939000_2058000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4840 diff_4036000_2051000# diff_4004000_2725000# diff_817000_2040000# GND efet w=20000 l=10000
+ ad=8.55e+08 pd=220000 as=0 ps=0 
M4841 diff_3938000_1940000# diff_95000_5192000# diff_3846000_1881000# GND efet w=12000 l=74000
+ ad=8.01e+08 pd=256000 as=0 ps=0 
M4842 diff_95000_5192000# diff_95000_5192000# diff_3846000_1881000# GND efet w=11000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4843 diff_95000_5192000# diff_95000_5192000# diff_3902000_1829000# GND efet w=13000 l=32000
+ ad=0 pd=0 as=1.05e+09 ps=194000 
M4844 diff_4057000_2151000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=32000
+ ad=0 pd=0 as=0 ps=0 
M4845 diff_4066000_2160000# diff_95000_5192000# diff_4036000_2051000# GND efet w=12000 l=79000
+ ad=0 pd=0 as=0 ps=0 
M4846 diff_4066000_2160000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4847 diff_817000_1965000# diff_3922000_786000# diff_3938000_1940000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4848 diff_4036000_1950000# diff_4004000_2725000# diff_817000_1965000# GND efet w=20000 l=10000
+ ad=8.46e+08 pd=238000 as=0 ps=0 
M4849 diff_95000_5192000# diff_95000_5192000# diff_4057000_1845000# GND efet w=13000 l=32000
+ ad=0 pd=0 as=9.92e+08 ps=190000 
M4850 diff_4066000_1853000# diff_95000_5192000# diff_4036000_1950000# GND efet w=12000 l=74000
+ ad=-3.14967e+08 pd=698000 as=0 ps=0 
M4851 diff_3577000_2123000# diff_3749000_2434000# diff_4066000_2160000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4852 diff_95000_5192000# diff_95000_5192000# diff_4066000_1853000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4853 diff_3696000_1783000# diff_3687000_1689000# diff_83000_3098000# GND efet w=204000 l=8000
+ ad=-3.21967e+08 pd=718000 as=0 ps=0 
M4854 diff_3687000_1689000# diff_3632000_1701000# diff_83000_3098000# GND efet w=70500 l=8500
+ ad=1.025e+09 pd=202000 as=0 ps=0 
M4855 diff_3577000_1746000# diff_3739000_826000# diff_3696000_1783000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4856 diff_3846000_1881000# diff_3695000_2725000# diff_3577000_1888000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4857 diff_83000_3098000# diff_3902000_1829000# diff_3846000_1881000# GND efet w=204000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4858 diff_3902000_1829000# diff_3938000_1940000# diff_83000_3098000# GND efet w=62500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4859 diff_817000_1663000# diff_3489000_2725000# diff_3632000_1701000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4860 diff_3687000_1689000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=32000
+ ad=0 pd=0 as=0 ps=0 
M4861 diff_3696000_1783000# diff_95000_5192000# diff_3632000_1701000# GND efet w=12500 l=78500
+ ad=0 pd=0 as=0 ps=0 
M4862 diff_3696000_1783000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4863 diff_817000_1588000# diff_3489000_2725000# diff_3632000_1546000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=9.87e+08 ps=234000 
M4864 diff_95000_5192000# diff_95000_5192000# diff_3686000_1562000# GND efet w=13000 l=32000
+ ad=0 pd=0 as=1.05e+09 ps=200000 
M4865 diff_3696000_1475000# diff_95000_5192000# diff_3632000_1546000# GND efet w=12000 l=74000
+ ad=-2.82967e+08 pd=716000 as=0 ps=0 
M4866 diff_95000_5192000# diff_95000_5192000# diff_3696000_1475000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4867 diff_3632000_1546000# diff_3354000_2409000# diff_848000_1588000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4868 diff_817000_1286000# diff_3171000_2725000# diff_3374000_1306000# GND efet w=19000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4869 diff_3117000_1087000# diff_3099000_1189000# diff_83000_3098000# GND efet w=212500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4870 diff_1851000_1079000# diff_3120000_2492000# diff_3117000_1087000# GND efet w=86000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4871 diff_817000_1211000# diff_2893000_2725000# diff_3117000_1087000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4872 diff_83000_3098000# diff_2534000_2492000# diff_1851000_999000# GND efet w=106500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M4873 diff_3117000_1023000# diff_3099000_927000# diff_83000_3098000# GND efet w=213500 l=7500
+ ad=-3.94967e+08 pd=692000 as=0 ps=0 
M4874 diff_3099000_927000# diff_3029000_910000# diff_83000_3098000# GND efet w=67500 l=8500
+ ad=9.82e+08 pd=198000 as=0 ps=0 
M4875 diff_817000_909000# diff_2638000_2492000# diff_3029000_910000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4876 diff_1851000_999000# diff_3120000_2492000# diff_3117000_1023000# GND efet w=86000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4877 diff_817000_909000# diff_2893000_2725000# diff_3117000_1023000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4878 diff_3099000_927000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=32000
+ ad=0 pd=0 as=0 ps=0 
M4879 diff_3117000_1023000# diff_95000_5192000# diff_3029000_910000# GND efet w=12000 l=81000
+ ad=0 pd=0 as=0 ps=0 
M4880 diff_3117000_1023000# diff_95000_5192000# diff_95000_5192000# GND efet w=11000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M4881 diff_83000_3098000# diff_72000_4515000# diff_2713000_822000# GND efet w=71000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4882 diff_2775000_765000# diff_72000_4515000# diff_83000_3098000# GND efet w=71000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4883 diff_83000_3098000# diff_72000_4515000# diff_2583000_2725000# GND efet w=70000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4884 diff_2843000_1950000# diff_72000_4515000# diff_83000_3098000# GND efet w=70000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4885 diff_83000_3098000# diff_72000_4515000# diff_2939000_824000# GND efet w=71000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4886 diff_2996000_2725000# diff_72000_4515000# diff_83000_3098000# GND efet w=71000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4887 diff_83000_3098000# diff_72000_4515000# diff_2638000_2492000# GND efet w=71000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4888 diff_2534000_2492000# diff_72000_4515000# diff_83000_3098000# GND efet w=71000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4889 diff_83000_3098000# diff_792000_356000# diff_969000_456000# GND efet w=506500 l=8500
+ ad=0 pd=0 as=1.76307e+09 ps=1.502e+06 
M4890 diff_95000_5192000# diff_792000_356000# diff_792000_356000# GND efet w=33000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4891 diff_969000_456000# diff_969000_456000# diff_95000_5192000# GND efet w=42000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4892 diff_969000_456000# diff_553000_1211000# diff_83000_3098000# GND efet w=331000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4893 diff_969000_456000# diff_553000_1211000# diff_83000_3098000# GND efet w=63000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4894 diff_135000_355000# diff_126000_347000# diff_95000_5192000# GND efet w=691500 l=8500
+ ad=-1.41774e+09 pd=4.186e+06 as=0 ps=0 
M4895 diff_801000_364000# diff_792000_356000# diff_83000_3098000# GND efet w=233000 l=9000
+ ad=-1.60771e+09 pd=4.316e+06 as=0 ps=0 
M4896 diff_83000_3098000# diff_553000_1211000# diff_126000_347000# GND efet w=275500 l=8500
+ ad=0 pd=0 as=-2.1289e+09 ps=1.608e+06 
M4897 diff_95000_5192000# diff_126000_347000# diff_135000_355000# GND efet w=244500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4898 diff_83000_3098000# diff_792000_356000# diff_801000_364000# GND efet w=195500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4899 diff_83000_3098000# diff_792000_356000# diff_801000_364000# GND efet w=195500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4900 diff_95000_5192000# diff_969000_456000# diff_801000_364000# GND efet w=351000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4901 diff_83000_3098000# diff_553000_1211000# diff_1204000_546000# GND efet w=440000 l=8000
+ ad=0 pd=0 as=-4.21902e+08 ps=1.994e+06 
M4902 diff_83000_3098000# diff_1277000_568000# diff_1204000_546000# GND efet w=486500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4903 diff_95000_5192000# diff_1204000_546000# diff_1204000_546000# GND efet w=52500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4904 diff_83000_3098000# diff_1399000_598000# diff_1383000_625000# GND efet w=231000 l=8000
+ ad=0 pd=0 as=-3.56967e+08 ps=640000 
M4905 diff_95000_5192000# diff_1383000_625000# diff_1383000_625000# GND efet w=16000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4906 diff_83000_3098000# diff_1204000_546000# diff_1430000_565000# GND efet w=275000 l=9000
+ ad=0 pd=0 as=2.00707e+09 ps=1.486e+06 
M4907 diff_1383000_625000# diff_680000_1019000# diff_1277000_568000# GND efet w=35000 l=11000
+ ad=0 pd=0 as=5.93e+08 ps=176000 
M4908 diff_83000_3098000# diff_553000_1211000# diff_1430000_565000# GND efet w=298000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4909 diff_1430000_565000# diff_1204000_546000# diff_83000_3098000# GND efet w=46000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4910 diff_95000_5192000# diff_969000_456000# diff_801000_364000# GND efet w=171000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4911 diff_95000_5192000# diff_969000_456000# diff_801000_364000# GND efet w=172000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4912 diff_83000_3098000# diff_553000_1211000# diff_126000_347000# GND efet w=120500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4913 diff_95000_5192000# diff_126000_347000# diff_135000_355000# GND efet w=244000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4914 diff_83000_3098000# diff_174000_153000# diff_126000_347000# GND efet w=499500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4915 diff_801000_364000# diff_792000_356000# diff_83000_3098000# GND efet w=512500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4916 diff_95000_5192000# diff_126000_347000# diff_135000_355000# GND efet w=488000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4917 diff_126000_347000# diff_126000_347000# diff_95000_5192000# GND efet w=42000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4918 diff_174000_153000# diff_174000_153000# diff_95000_5192000# GND efet w=34000 l=9000
+ ad=2.07507e+09 pd=1.452e+06 as=0 ps=0 
M4919 diff_83000_3098000# diff_174000_153000# diff_135000_355000# GND efet w=604000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4920 diff_135000_355000# diff_174000_153000# diff_83000_3098000# GND efet w=830000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4921 diff_83000_3098000# diff_553000_1211000# diff_174000_153000# GND efet w=377500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4922 diff_709000_308000# diff_680000_1019000# diff_692000_115000# GND efet w=34000 l=11000
+ ad=0 pd=0 as=5.25e+08 ps=130000 
M4923 diff_83000_3098000# diff_692000_115000# diff_174000_153000# GND efet w=395500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4924 diff_801000_364000# diff_792000_356000# diff_83000_3098000# GND efet w=276000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4925 diff_95000_5192000# diff_969000_456000# diff_801000_364000# GND efet w=120500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4926 diff_1218000_195000# diff_1204000_546000# diff_95000_5192000# GND efet w=189000 l=8000
+ ad=-1.98706e+08 pd=4.556e+06 as=0 ps=0 
M4927 diff_95000_5192000# diff_1204000_546000# diff_1218000_195000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4928 diff_1218000_195000# diff_1204000_546000# diff_95000_5192000# GND efet w=650000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4929 diff_95000_5192000# diff_1204000_546000# diff_1218000_195000# GND efet w=203000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4930 diff_95000_5192000# diff_1204000_546000# diff_1218000_195000# GND efet w=206500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4931 diff_1430000_565000# diff_1430000_565000# diff_95000_5192000# GND efet w=35000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4932 diff_1430000_565000# diff_553000_1211000# diff_83000_3098000# GND efet w=54000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4933 diff_83000_3098000# diff_1430000_565000# diff_1218000_195000# GND efet w=191500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4934 diff_83000_3098000# diff_553000_1211000# diff_1620000_123000# GND efet w=55000 l=9000
+ ad=0 pd=0 as=1.87907e+09 ps=1.488e+06 
M4935 diff_83000_3098000# diff_553000_1211000# diff_1620000_123000# GND efet w=301000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4936 diff_83000_3098000# diff_1694000_585000# diff_1620000_123000# GND efet w=274000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4937 diff_83000_3098000# diff_72000_4515000# diff_3120000_2492000# GND efet w=71000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4938 diff_2893000_2725000# diff_72000_4515000# diff_83000_3098000# GND efet w=71000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4939 diff_95000_5192000# diff_95000_5192000# diff_1851000_1079000# GND efet w=12000 l=103000
+ ad=0 pd=0 as=0 ps=0 
M4940 diff_3428000_1309000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=32000
+ ad=0 pd=0 as=0 ps=0 
M4941 diff_3436000_1405000# diff_95000_5192000# diff_3374000_1306000# GND efet w=12500 l=79500
+ ad=0 pd=0 as=0 ps=0 
M4942 diff_3436000_1405000# diff_95000_5192000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4943 diff_95000_5192000# diff_95000_5192000# diff_3427000_1189000# GND efet w=12000 l=33000
+ ad=0 pd=0 as=9.25e+08 ps=190000 
M4944 diff_3436000_1099000# diff_95000_5192000# diff_3374000_1153000# GND efet w=12000 l=74000
+ ad=2.80327e+07 pd=728000 as=1.524e+09 ps=370000 
M4945 diff_95000_5192000# diff_95000_5192000# diff_3436000_1099000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4946 diff_817000_1211000# diff_3171000_2725000# diff_3374000_1153000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4947 diff_3436000_1405000# diff_3439000_2492000# diff_817000_1286000# GND efet w=104500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4948 diff_3577000_1368000# diff_3567000_785000# diff_3436000_1405000# GND efet w=108000 l=10000
+ ad=-2.06493e+09 pd=1.358e+06 as=0 ps=0 
M4949 diff_848000_1262000# diff_3596000_2395000# diff_3577000_1368000# GND efet w=120000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4950 diff_3632000_1324000# diff_3354000_2409000# diff_848000_1262000# GND efet w=19000 l=10000
+ ad=1.011e+09 pd=246000 as=0 ps=0 
M4951 diff_3436000_1099000# diff_3439000_2492000# diff_817000_1211000# GND efet w=105500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4952 diff_3577000_1134000# diff_3567000_785000# diff_3436000_1099000# GND efet w=109000 l=10000
+ ad=-2.09093e+09 pd=1.362e+06 as=0 ps=0 
M4953 diff_3374000_1153000# diff_3354000_2409000# diff_1851000_1079000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4954 diff_3374000_929000# diff_3354000_2409000# diff_1851000_999000# GND efet w=20000 l=9000
+ ad=1.534e+09 pd=388000 as=0 ps=0 
M4955 diff_1851000_999000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=103000
+ ad=0 pd=0 as=0 ps=0 
M4956 diff_3427000_1189000# diff_3374000_1153000# diff_83000_3098000# GND efet w=64000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4957 diff_3436000_1099000# diff_3427000_1189000# diff_83000_3098000# GND efet w=204500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4958 diff_1851000_1079000# diff_3474000_792000# diff_3436000_1099000# GND efet w=86000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4959 diff_3436000_1028000# diff_3428000_935000# diff_83000_3098000# GND efet w=205500 l=7500
+ ad=-3.99673e+07 pd=710000 as=0 ps=0 
M4960 diff_3428000_935000# diff_3374000_929000# diff_83000_3098000# GND efet w=72000 l=8000
+ ad=9.26e+08 pd=190000 as=0 ps=0 
M4961 diff_1851000_999000# diff_3474000_792000# diff_3436000_1028000# GND efet w=86000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4962 diff_848000_1211000# diff_3596000_2395000# diff_3577000_1134000# GND efet w=120000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4963 diff_817000_1663000# diff_3800000_830000# diff_3696000_1783000# GND efet w=102500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M4964 diff_3846000_1700000# diff_3830000_787000# diff_817000_1663000# GND efet w=102500 l=9500
+ ad=-1.71967e+08 pd=720000 as=0 ps=0 
M4965 diff_3846000_1700000# diff_3695000_2725000# diff_3577000_1746000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4966 diff_83000_3098000# diff_3902000_1795000# diff_3846000_1700000# GND efet w=204000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4967 diff_3902000_1795000# diff_3939000_1680000# diff_83000_3098000# GND efet w=63000 l=8000
+ ad=1.048e+09 pd=194000 as=0 ps=0 
M4968 diff_817000_1588000# diff_3800000_830000# diff_3696000_1475000# GND efet w=102000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4969 diff_3846000_1504000# diff_3830000_787000# diff_817000_1588000# GND efet w=102500 l=9500
+ ad=-1.40967e+08 pd=716000 as=0 ps=0 
M4970 diff_3686000_1562000# diff_3632000_1546000# diff_83000_3098000# GND efet w=65500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4971 diff_3696000_1475000# diff_3686000_1562000# diff_83000_3098000# GND efet w=203000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4972 diff_3577000_1511000# diff_3739000_826000# diff_3696000_1475000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4973 diff_4057000_1845000# diff_4036000_1950000# diff_83000_3098000# GND efet w=60500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4974 diff_4066000_1853000# diff_4057000_1845000# diff_83000_3098000# GND efet w=203500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M4975 diff_817000_1965000# diff_4108000_2725000# diff_4066000_1853000# GND efet w=86000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4976 diff_3577000_1888000# diff_3749000_2434000# diff_4066000_1853000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M4977 diff_4462000_2971000# diff_4462000_2971000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M4978 diff_83000_3098000# diff_4495000_3314000# diff_4517000_3010000# GND efet w=72000 l=8000
+ ad=0 pd=0 as=1.154e+09 ps=266000 
M4979 diff_4591000_3170000# diff_4517000_3010000# diff_83000_3098000# GND efet w=64000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M4980 diff_83000_3098000# diff_4591000_3170000# diff_4656000_3020000# GND efet w=104000 l=8000
+ ad=0 pd=0 as=4.59033e+08 ps=934000 
M4981 diff_4656000_3020000# diff_860000_2987000# diff_83000_3098000# GND efet w=114000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4982 diff_83000_3098000# diff_906000_3226000# diff_4656000_3020000# GND efet w=113500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M4983 diff_95000_5192000# diff_4591000_3170000# diff_4591000_3170000# GND efet w=11000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M4984 diff_4517000_3010000# diff_4517000_3010000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M4985 diff_4656000_3020000# diff_4656000_3020000# diff_95000_5192000# GND efet w=13000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M4986 diff_4716000_3243000# diff_72000_4515000# diff_4843000_3181000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=5.24e+08 ps=140000 
M4987 diff_4814000_3335000# diff_72000_4515000# diff_4865000_3205000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=3.98e+08 ps=120000 
M4988 diff_83000_3098000# diff_4779000_3198000# diff_4777000_2951000# GND efet w=72500 l=8500
+ ad=0 pd=0 as=-1.14497e+09 ps=660000 
M4989 diff_4777000_2951000# diff_3569000_3530000# diff_83000_3098000# GND efet w=62000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4990 diff_83000_3098000# diff_4843000_3181000# diff_4843000_3067000# GND efet w=63000 l=8000
+ ad=0 pd=0 as=3.31033e+08 ps=874000 
M4991 diff_4843000_3067000# diff_4865000_3205000# diff_83000_3098000# GND efet w=63000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M4992 diff_4806000_4501000# diff_72000_4515000# diff_4923000_2911000# GND efet w=11000 l=11000
+ ad=0 pd=0 as=3.33e+08 ps=110000 
M4993 diff_95000_5192000# diff_4777000_2951000# diff_4777000_2951000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M4994 diff_4904000_3051000# diff_68000_5288000# diff_817000_1286000# GND efet w=12000 l=11000
+ ad=6.19e+08 pd=128000 as=0 ps=0 
M4995 diff_4966000_3079000# diff_4904000_3051000# diff_83000_3098000# GND efet w=131000 l=9000
+ ad=1.179e+09 pd=280000 as=0 ps=0 
M4996 diff_4983000_2920000# diff_4927000_3400000# diff_4966000_3079000# GND efet w=131000 l=8000
+ ad=9.08033e+08 pd=882000 as=0 ps=0 
M4997 diff_5439000_3442000# diff_5357000_3322000# diff_83000_3098000# GND efet w=97000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M4998 diff_5920000_3449000# diff_5920000_3449000# diff_95000_5192000# GND efet w=12000 l=37000
+ ad=1.876e+09 pd=492000 as=0 ps=0 
M4999 diff_3254000_2509000# diff_72000_4515000# diff_5432000_3451000# GND efet w=13000 l=11000
+ ad=1.445e+09 pd=300000 as=3.18e+08 ps=82000 
M5000 diff_5920000_3449000# diff_5068000_4962000# diff_6006000_3447000# GND efet w=85000 l=9000
+ ad=0 pd=0 as=7.65e+08 ps=188000 
M5001 diff_6160000_3457000# diff_5920000_3449000# diff_6112000_3388000# GND efet w=90500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5002 diff_95000_5192000# diff_3254000_2509000# diff_3254000_2509000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5003 diff_3254000_2509000# diff_5578000_3393000# diff_83000_3098000# GND efet w=72000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5004 diff_6006000_3447000# diff_5098000_4894000# diff_83000_3098000# GND efet w=85000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5005 diff_4883000_4962000# diff_72000_4515000# diff_5407000_3340000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=5.34e+08 ps=134000 
M5006 diff_5531000_3344000# diff_4265000_3070000# diff_83000_3098000# GND efet w=93000 l=8000
+ ad=9.65e+08 pd=224000 as=0 ps=0 
M5007 diff_83000_3098000# diff_5039000_4962000# diff_6076000_3942000# GND efet w=42000 l=9000
+ ad=0 pd=0 as=-1.69697e+09 ps=554000 
M5008 diff_6120000_3397000# diff_6112000_3388000# diff_83000_3098000# GND efet w=103500 l=8500
+ ad=2.012e+09 pd=382000 as=0 ps=0 
M5009 diff_83000_3098000# diff_5696000_3194000# diff_6120000_3397000# GND efet w=90000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5010 diff_95000_5192000# diff_6076000_3942000# diff_6076000_3942000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M5011 diff_6076000_3942000# diff_6180000_3356000# diff_6120000_3397000# GND efet w=88000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5012 diff_5531000_3344000# diff_5407000_3340000# diff_5048000_3693000# GND efet w=103000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5013 diff_83000_3098000# diff_5407000_3340000# diff_5357000_3322000# GND efet w=48000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5014 diff_83000_3098000# diff_5009000_4962000# diff_5696000_3194000# GND efet w=66000 l=9000
+ ad=0 pd=0 as=1.725e+09 ps=386000 
M5015 diff_95000_5192000# diff_6180000_3356000# diff_6180000_3356000# GND efet w=11000 l=35000
+ ad=0 pd=0 as=1.657e+09 ps=346000 
M5016 diff_83000_3098000# diff_5469000_3309000# diff_5357000_3322000# GND efet w=44000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5017 diff_5357000_3322000# diff_5357000_3322000# diff_95000_5192000# GND efet w=12000 l=34000
+ ad=0 pd=0 as=0 ps=0 
M5018 diff_5048000_3693000# diff_5469000_3309000# diff_83000_3098000# GND efet w=42000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5019 diff_5469000_3309000# diff_72000_4515000# diff_65000_4220000# GND efet w=12000 l=12000
+ ad=2.43e+08 pd=70000 as=0 ps=0 
M5020 diff_5084000_3006000# diff_68000_5288000# diff_4983000_2920000# GND efet w=12000 l=12000
+ ad=5.6e+08 pd=136000 as=0 ps=0 
M5021 diff_95000_5192000# diff_4265000_3070000# diff_4265000_3070000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=1.658e+09 ps=358000 
M5022 diff_4265000_3070000# diff_5576000_3241000# diff_83000_3098000# GND efet w=78500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5023 diff_95000_5192000# diff_4843000_3067000# diff_4843000_3067000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M5024 diff_83000_3098000# diff_4923000_2911000# diff_4912000_2900000# GND efet w=142000 l=7000
+ ad=0 pd=0 as=-1.61897e+09 ps=508000 
M5025 diff_4983000_2920000# diff_4975000_2910000# diff_4912000_2900000# GND efet w=142000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5026 diff_5010000_3006000# diff_4871000_3351000# diff_4983000_2920000# GND efet w=129000 l=8000
+ ad=1.161e+09 pd=276000 as=0 ps=0 
M5027 diff_83000_3098000# diff_5019000_2993000# diff_5010000_3006000# GND efet w=129000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5028 diff_3321000_2527000# diff_72000_4515000# diff_5019000_2993000# GND efet w=12000 l=10000
+ ad=1.964e+09 pd=392000 as=3.39e+08 ps=118000 
M5029 diff_83000_3098000# diff_5084000_3006000# diff_3321000_2527000# GND efet w=92500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5030 diff_95000_5192000# diff_4983000_2920000# diff_4983000_2920000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M5031 diff_95000_5192000# diff_3321000_2527000# diff_3321000_2527000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M5032 diff_4954000_639000# diff_72000_4515000# diff_83000_3098000# GND efet w=272000 l=9000
+ ad=1.60803e+09 pd=848000 as=0 ps=0 
M5033 diff_83000_3098000# diff_5214000_3050000# diff_4954000_639000# GND efet w=270000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5034 diff_83000_3098000# diff_5087000_472000# diff_5214000_3050000# GND efet w=125500 l=8500
+ ad=0 pd=0 as=-2.08297e+09 ps=334000 
M5035 diff_5696000_3194000# diff_72000_4515000# diff_5576000_3241000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=2.32e+08 ps=68000 
M5036 diff_5696000_3194000# diff_5696000_3194000# diff_95000_5192000# GND efet w=11000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M5037 diff_6180000_3356000# diff_5696000_3194000# diff_6269000_3300000# GND efet w=131000 l=9000
+ ad=0 pd=0 as=1.179e+09 ps=280000 
M5038 diff_6269000_3300000# diff_5068000_4962000# diff_6269000_3282000# GND efet w=131000 l=8000
+ ad=0 pd=0 as=1.31e+09 ps=282000 
M5039 diff_6269000_3282000# diff_6252000_3157000# diff_83000_3098000# GND efet w=131000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5040 diff_5214000_3050000# diff_5214000_3050000# diff_95000_5192000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5041 diff_4358000_3758000# diff_72000_4515000# diff_4391000_2778000# GND efet w=19000 l=14000
+ ad=0 pd=0 as=9.09e+08 ps=148000 
M5042 diff_4415000_3774000# diff_72000_4515000# diff_4443000_2778000# GND efet w=20000 l=13000
+ ad=0 pd=0 as=9.36e+08 ps=150000 
M5043 diff_4462000_2971000# diff_72000_4515000# diff_4494000_2778000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=9.09e+08 ps=148000 
M5044 diff_4462000_3008000# diff_72000_4515000# diff_4546000_2778000# GND efet w=19000 l=13000
+ ad=0 pd=0 as=9.01e+08 ps=148000 
M5045 diff_4697000_3226000# diff_72000_4515000# diff_4689000_2592000# GND efet w=12000 l=8000
+ ad=0 pd=0 as=9.75e+08 ps=148000 
M5046 diff_4716000_3243000# diff_72000_4515000# diff_4785000_2783000# GND efet w=13000 l=9000
+ ad=0 pd=0 as=1.057e+09 ps=178000 
M5047 diff_95000_5192000# diff_4602000_2752000# diff_4602000_2752000# GND efet w=18000 l=8000
+ ad=0 pd=0 as=3.01033e+08 ps=964000 
M5048 diff_4374000_833000# diff_4391000_2778000# diff_83000_3098000# GND efet w=245000 l=8000
+ ad=6.75033e+08 pd=942000 as=0 ps=0 
M5049 diff_95000_5192000# diff_4374000_833000# diff_4374000_833000# GND efet w=18000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M5050 diff_4417000_952000# diff_4417000_952000# diff_95000_5192000# GND efet w=18000 l=7000
+ ad=3.58033e+08 pd=886000 as=0 ps=0 
M5051 diff_83000_3098000# diff_72000_4515000# diff_4374000_833000# GND efet w=203000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5052 diff_4417000_952000# diff_72000_4515000# diff_83000_3098000# GND efet w=203000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5053 diff_83000_3098000# diff_4443000_2778000# diff_4417000_952000# GND efet w=244000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5054 diff_4498000_2492000# diff_4494000_2778000# diff_83000_3098000# GND efet w=245000 l=8000
+ ad=2.63033e+08 pd=886000 as=0 ps=0 
M5055 diff_95000_5192000# diff_4498000_2492000# diff_4498000_2492000# GND efet w=18000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5056 diff_4548000_2725000# diff_4548000_2725000# diff_95000_5192000# GND efet w=18000 l=8000
+ ad=4.64033e+08 pd=886000 as=0 ps=0 
M5057 diff_83000_3098000# diff_72000_4515000# diff_4498000_2492000# GND efet w=204000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5058 diff_4548000_2725000# diff_72000_4515000# diff_83000_3098000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5059 diff_83000_3098000# diff_4546000_2778000# diff_4548000_2725000# GND efet w=244500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5060 diff_4328000_910000# diff_4328000_910000# diff_95000_5192000# GND efet w=24000 l=8000
+ ad=-4.66935e+08 pd=1.438e+06 as=0 ps=0 
M5061 diff_4777000_2951000# diff_68000_5288000# diff_4883000_2653000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=9.28e+08 ps=162000 
M5062 diff_83000_3098000# diff_72000_4515000# diff_4602000_2752000# GND efet w=200500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5063 diff_83000_3098000# diff_4224000_2739000# diff_817000_1965000# GND efet w=87000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5064 diff_4066000_1783000# diff_4057000_1774000# diff_83000_3098000# GND efet w=203500 l=7500
+ ad=-3.66967e+08 pd=696000 as=0 ps=0 
M5065 diff_83000_3098000# diff_4037000_1674000# diff_4057000_1774000# GND efet w=60500 l=8500
+ ad=0 pd=0 as=9.51e+08 ps=186000 
M5066 diff_817000_1663000# diff_4108000_2725000# diff_4066000_1783000# GND efet w=86000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5067 diff_83000_3098000# diff_3901000_2725000# diff_3577000_1888000# GND efet w=105000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5068 diff_4235000_1886000# diff_4066000_2160000# diff_83000_3098000# GND efet w=75000 l=8000
+ ad=-1.67297e+09 pd=410000 as=0 ps=0 
M5069 diff_83000_3098000# diff_4066000_1853000# diff_4235000_1886000# GND efet w=72000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5070 diff_83000_3098000# diff_3901000_2725000# diff_3577000_1746000# GND efet w=105500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5071 diff_3846000_1700000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5072 diff_3939000_1680000# diff_95000_5192000# diff_3846000_1700000# GND efet w=12500 l=77500
+ ad=8.1e+08 pd=232000 as=0 ps=0 
M5073 diff_3902000_1795000# diff_95000_5192000# diff_95000_5192000# GND efet w=13000 l=31000
+ ad=0 pd=0 as=0 ps=0 
M5074 diff_817000_1663000# diff_3922000_786000# diff_3939000_1680000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5075 diff_4037000_1674000# diff_4004000_2725000# diff_817000_1663000# GND efet w=20000 l=11000
+ ad=8.47e+08 pd=220000 as=0 ps=0 
M5076 diff_3938000_1563000# diff_95000_5192000# diff_3846000_1504000# GND efet w=12000 l=75000
+ ad=7.84e+08 pd=248000 as=0 ps=0 
M5077 diff_95000_5192000# diff_95000_5192000# diff_3846000_1504000# GND efet w=11000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5078 diff_95000_5192000# diff_95000_5192000# diff_3902000_1451000# GND efet w=13000 l=32000
+ ad=0 pd=0 as=1.022e+09 ps=192000 
M5079 diff_4057000_1774000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=31000
+ ad=0 pd=0 as=0 ps=0 
M5080 diff_4066000_1783000# diff_95000_5192000# diff_4037000_1674000# GND efet w=12000 l=78000
+ ad=0 pd=0 as=0 ps=0 
M5081 diff_4066000_1783000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5082 diff_4066000_1475000# diff_95000_5192000# diff_4037000_1573000# GND efet w=12000 l=75000
+ ad=-3.29967e+08 pd=692000 as=8.29e+08 ps=232000 
M5083 diff_817000_1588000# diff_3922000_786000# diff_3938000_1563000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5084 diff_4037000_1573000# diff_4004000_2725000# diff_817000_1588000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5085 diff_95000_5192000# diff_95000_5192000# diff_4057000_1467000# GND efet w=13000 l=32000
+ ad=0 pd=0 as=9.65e+08 ps=188000 
M5086 diff_3577000_1746000# diff_3749000_2434000# diff_4066000_1783000# GND efet w=87000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5087 diff_4226000_1649000# diff_4066000_1783000# diff_4235000_1886000# GND efet w=71000 l=8000
+ ad=-2.04797e+09 pd=402000 as=0 ps=0 
M5088 diff_95000_5192000# diff_95000_5192000# diff_4066000_1475000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5089 diff_3696000_1405000# diff_3687000_1311000# diff_83000_3098000# GND efet w=204000 l=8000
+ ad=-3.81967e+08 pd=714000 as=0 ps=0 
M5090 diff_3687000_1311000# diff_3632000_1324000# diff_83000_3098000# GND efet w=70500 l=8500
+ ad=1.029e+09 pd=202000 as=0 ps=0 
M5091 diff_3577000_1368000# diff_3739000_826000# diff_3696000_1405000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5092 diff_3846000_1504000# diff_3695000_2725000# diff_3577000_1511000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5093 diff_83000_3098000# diff_3902000_1451000# diff_3846000_1504000# GND efet w=204000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5094 diff_3902000_1451000# diff_3938000_1563000# diff_83000_3098000# GND efet w=62000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5095 diff_817000_1286000# diff_3489000_2725000# diff_3632000_1324000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5096 diff_3687000_1311000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=32000
+ ad=0 pd=0 as=0 ps=0 
M5097 diff_3696000_1405000# diff_95000_5192000# diff_3632000_1324000# GND efet w=12500 l=78500
+ ad=0 pd=0 as=0 ps=0 
M5098 diff_3696000_1405000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5099 diff_817000_1211000# diff_3489000_2725000# diff_3632000_1169000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=9.87e+08 ps=234000 
M5100 diff_95000_5192000# diff_95000_5192000# diff_3686000_1185000# GND efet w=13000 l=33000
+ ad=0 pd=0 as=1.046e+09 ps=200000 
M5101 diff_3696000_1098000# diff_95000_5192000# diff_3632000_1169000# GND efet w=12000 l=74000
+ ad=-1.94967e+08 pd=718000 as=0 ps=0 
M5102 diff_95000_5192000# diff_95000_5192000# diff_3696000_1098000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5103 diff_3632000_1169000# diff_3354000_2409000# diff_848000_1211000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5104 diff_817000_909000# diff_3171000_2725000# diff_3374000_929000# GND efet w=19000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5105 diff_3428000_935000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=33000
+ ad=0 pd=0 as=0 ps=0 
M5106 diff_3436000_1028000# diff_95000_5192000# diff_3374000_929000# GND efet w=12500 l=81500
+ ad=0 pd=0 as=0 ps=0 
M5107 diff_3436000_1028000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5108 diff_3436000_1028000# diff_3439000_2492000# diff_817000_909000# GND efet w=104500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5109 diff_3577000_991000# diff_3567000_785000# diff_3436000_1028000# GND efet w=107500 l=9500
+ ad=-1.95493e+09 pd=1.346e+06 as=0 ps=0 
M5110 diff_848000_885000# diff_3596000_2395000# diff_3577000_991000# GND efet w=120000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5111 diff_3631000_947000# diff_3354000_2409000# diff_848000_885000# GND efet w=19000 l=10000
+ ad=1.027e+09 pd=254000 as=0 ps=0 
M5112 diff_3354000_2409000# diff_72000_4515000# diff_83000_3098000# GND efet w=81000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5113 diff_3171000_2725000# diff_72000_4515000# diff_83000_3098000# GND efet w=84000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5114 diff_817000_1286000# diff_3800000_830000# diff_3696000_1405000# GND efet w=102000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5115 diff_3846000_1323000# diff_3830000_787000# diff_817000_1286000# GND efet w=102000 l=10000
+ ad=-1.78967e+08 pd=718000 as=0 ps=0 
M5116 diff_3846000_1323000# diff_3695000_2725000# diff_3577000_1368000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5117 diff_83000_3098000# diff_3902000_1418000# diff_3846000_1323000# GND efet w=205000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5118 diff_3902000_1418000# diff_3939000_1303000# diff_83000_3098000# GND efet w=63500 l=7500
+ ad=1.06e+09 pd=194000 as=0 ps=0 
M5119 diff_817000_1211000# diff_3800000_830000# diff_3696000_1098000# GND efet w=101500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5120 diff_3846000_1128000# diff_3830000_787000# diff_817000_1211000# GND efet w=101000 l=10000
+ ad=-7.49673e+07 pd=714000 as=0 ps=0 
M5121 diff_3686000_1185000# diff_3632000_1169000# diff_83000_3098000# GND efet w=64500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5122 diff_3696000_1098000# diff_3686000_1185000# diff_83000_3098000# GND efet w=202000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5123 diff_3577000_1134000# diff_3739000_826000# diff_3696000_1098000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5124 diff_4057000_1467000# diff_4037000_1573000# diff_83000_3098000# GND efet w=60000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5125 diff_4066000_1475000# diff_4057000_1467000# diff_83000_3098000# GND efet w=203500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5126 diff_817000_1588000# diff_4108000_2725000# diff_4066000_1475000# GND efet w=86000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5127 diff_3577000_1511000# diff_3749000_2434000# diff_4066000_1475000# GND efet w=85000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5128 diff_817000_1663000# diff_4277000_2781000# diff_83000_3098000# GND efet w=84000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5129 diff_83000_3098000# diff_3321000_2527000# diff_4275000_1613000# GND efet w=43000 l=9000
+ ad=0 pd=0 as=8.36e+08 ps=168000 
M5130 diff_4226000_1649000# diff_4226000_1649000# diff_95000_5192000# GND efet w=11000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M5131 diff_4275000_1613000# diff_4275000_1613000# diff_95000_5192000# GND efet w=13000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M5132 diff_95000_5192000# diff_4285000_1501000# diff_4285000_1501000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=-2.16967e+08 ps=832000 
M5133 diff_4066000_1405000# diff_4057000_1397000# diff_83000_3098000# GND efet w=204500 l=7500
+ ad=-3.71967e+08 pd=694000 as=0 ps=0 
M5134 diff_83000_3098000# diff_4036000_1297000# diff_4057000_1397000# GND efet w=61000 l=8000
+ ad=0 pd=0 as=9.6e+08 ps=186000 
M5135 diff_817000_1286000# diff_4108000_2725000# diff_4066000_1405000# GND efet w=86000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5136 diff_83000_3098000# diff_3901000_2725000# diff_3577000_1511000# GND efet w=106500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5137 diff_83000_3098000# diff_3901000_2725000# diff_3577000_1368000# GND efet w=105000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5138 diff_4266000_1501000# diff_4226000_1649000# diff_83000_3098000# GND efet w=101000 l=9000
+ ad=1.01e+09 pd=222000 as=0 ps=0 
M5139 diff_4285000_1501000# diff_4275000_1613000# diff_4266000_1501000# GND efet w=101000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5140 diff_95000_5192000# diff_4253000_1284000# diff_4253000_1284000# GND efet w=12000 l=38000
+ ad=0 pd=0 as=9.34e+08 ps=206000 
M5141 diff_3577000_2265000# diff_4328000_910000# diff_95000_5192000# GND efet w=99500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5142 diff_3577000_2123000# diff_4328000_910000# diff_95000_5192000# GND efet w=100000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5143 diff_83000_3098000# diff_4602000_2752000# diff_4328000_910000# GND efet w=449000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5144 diff_4760000_2748000# diff_68000_5288000# diff_4705000_2611000# GND efet w=14000 l=12000
+ ad=9.4e+08 pd=160000 as=1.931e+09 ps=386000 
M5145 diff_4740000_2641000# diff_4740000_2641000# diff_95000_5192000# GND efet w=12000 l=8000
+ ad=-1.64797e+09 pd=608000 as=0 ps=0 
M5146 diff_95000_5192000# diff_4705000_2611000# diff_4705000_2611000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M5147 diff_4705000_2611000# diff_4689000_2592000# diff_83000_3098000# GND efet w=66500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5148 diff_83000_3098000# diff_4760000_2748000# diff_4740000_2641000# GND efet w=161500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5149 diff_4837000_2758000# diff_68000_5288000# diff_4805000_2759000# GND efet w=15000 l=11000
+ ad=1.002e+09 pd=168000 as=1.74e+09 ps=368000 
M5150 diff_4839000_2618000# diff_4839000_2618000# diff_95000_5192000# GND efet w=12000 l=8000
+ ad=-1.72097e+09 pd=570000 as=0 ps=0 
M5151 diff_4768000_996000# diff_4768000_996000# diff_95000_5192000# GND efet w=12000 l=8000
+ ad=-1.34197e+09 pd=638000 as=0 ps=0 
M5152 diff_4768000_996000# diff_4883000_2653000# diff_83000_3098000# GND efet w=167500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5153 diff_95000_5192000# diff_4805000_2759000# diff_4805000_2759000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5154 diff_4805000_2759000# diff_4785000_2783000# diff_83000_3098000# GND efet w=76000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5155 diff_4433000_2246000# diff_4374000_833000# diff_83000_3098000# GND efet w=20000 l=10000
+ ad=1.675e+09 pd=328000 as=0 ps=0 
M5156 diff_4459000_2246000# diff_4417000_952000# diff_4433000_2246000# GND efet w=20000 l=10000
+ ad=-9.77967e+08 pd=722000 as=0 ps=0 
M5157 diff_95000_5192000# diff_95000_5192000# diff_3577000_2265000# GND efet w=13000 l=103000
+ ad=0 pd=0 as=0 ps=0 
M5158 diff_95000_5192000# diff_4518000_2327000# diff_4518000_2327000# GND efet w=12000 l=19000
+ ad=0 pd=0 as=2.035e+09 ps=412000 
M5159 diff_4518000_2327000# diff_3577000_2265000# diff_83000_3098000# GND efet w=49000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5160 diff_95000_5192000# diff_4575000_2328000# diff_4575000_2328000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=1.582e+09 ps=308000 
M5161 diff_95000_5192000# diff_4608000_2224000# diff_4608000_2224000# GND efet w=13000 l=20000
+ ad=0 pd=0 as=1.819e+09 ps=406000 
M5162 diff_4575000_2328000# diff_4498000_2492000# diff_4433000_2246000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5163 diff_83000_3098000# diff_4837000_2758000# diff_4839000_2618000# GND efet w=160000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5164 diff_95000_5192000# diff_4945000_2494000# diff_4945000_2494000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=1.27033e+08 ps=724000 
M5165 diff_5170000_2830000# diff_72000_4515000# diff_4975000_2910000# GND efet w=13000 l=11000
+ ad=2.043e+09 pd=430000 as=7.86e+08 ps=206000 
M5166 diff_4762000_3821000# diff_72000_4515000# diff_4932000_2482000# GND efet w=15000 l=11000
+ ad=0 pd=0 as=1.101e+09 ps=158000 
M5167 diff_4843000_3067000# diff_68000_5288000# diff_5114000_2490000# GND efet w=20000 l=12000
+ ad=0 pd=0 as=5.28e+08 ps=118000 
M5168 diff_4954000_639000# diff_4954000_639000# diff_95000_5192000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5169 diff_4495000_3314000# diff_72000_4515000# diff_5265000_2778000# GND efet w=20000 l=12000
+ ad=0 pd=0 as=8.98e+08 ps=152000 
M5170 diff_4656000_3020000# diff_72000_4515000# diff_5318000_2778000# GND efet w=20000 l=12000
+ ad=0 pd=0 as=9.1e+08 ps=136000 
M5171 diff_5012000_2755000# diff_68000_5288000# diff_4959000_2608000# GND efet w=14000 l=11000
+ ad=1.008e+09 pd=170000 as=1.541e+09 ps=324000 
M5172 diff_95000_5192000# diff_4932000_827000# diff_4932000_827000# GND efet w=17000 l=9000
+ ad=0 pd=0 as=7.37033e+08 ps=924000 
M5173 diff_4994000_2634000# diff_4994000_2634000# diff_95000_5192000# GND efet w=13000 l=8000
+ ad=2.092e+09 pd=484000 as=0 ps=0 
M5174 diff_83000_3098000# diff_5012000_2755000# diff_4994000_2634000# GND efet w=176500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5175 diff_4932000_827000# diff_4328000_910000# diff_83000_3098000# GND efet w=233000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5176 diff_83000_3098000# diff_72000_4515000# diff_4932000_827000# GND efet w=212500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5177 diff_5187000_2412000# diff_5187000_2412000# diff_95000_5192000# GND efet w=11000 l=15000
+ ad=-8.34967e+08 pd=662000 as=0 ps=0 
M5178 diff_95000_5192000# diff_4959000_2608000# diff_4959000_2608000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5179 diff_4959000_2608000# diff_4945000_2494000# diff_83000_3098000# GND efet w=74000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5180 diff_83000_3098000# diff_4932000_2482000# diff_4945000_2494000# GND efet w=63000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5181 diff_95000_5192000# diff_4694000_2317000# diff_4694000_2317000# GND efet w=13000 l=25000
+ ad=0 pd=0 as=-1.19197e+09 ps=546000 
M5182 diff_95000_5192000# diff_4727000_2238000# diff_4727000_2238000# GND efet w=13000 l=25000
+ ad=0 pd=0 as=1.506e+09 ps=296000 
M5183 diff_3577000_2123000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=103000
+ ad=0 pd=0 as=0 ps=0 
M5184 diff_4518000_2032000# diff_3577000_2123000# diff_83000_3098000# GND efet w=49000 l=8000
+ ad=1.967e+09 pd=410000 as=0 ps=0 
M5185 diff_83000_3098000# diff_4608000_2224000# diff_4575000_2328000# GND efet w=48000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5186 diff_4608000_2224000# diff_817000_2342000# diff_83000_3098000# GND efet w=67000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5187 diff_4433000_2246000# diff_4548000_2725000# diff_4608000_2224000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5188 diff_4705000_2274000# diff_4602000_2752000# diff_4433000_2246000# GND efet w=21000 l=12000
+ ad=3.99e+08 pd=80000 as=0 ps=0 
M5189 diff_4459000_2246000# diff_4498000_2492000# diff_4433000_2037000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=-1.84497e+09 ps=524000 
M5190 diff_83000_3098000# diff_4608000_2077000# diff_4459000_2246000# GND efet w=50000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5191 diff_4608000_2077000# diff_817000_2040000# diff_83000_3098000# GND efet w=67000 l=8000
+ ad=1.808e+09 pd=404000 as=0 ps=0 
M5192 diff_4705000_2229000# diff_4602000_2752000# diff_4518000_2327000# GND efet w=20000 l=12000
+ ad=4.42e+08 pd=136000 as=0 ps=0 
M5193 diff_83000_3098000# diff_4705000_2229000# diff_4727000_2238000# GND efet w=49000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5194 diff_4786000_2230000# diff_4740000_2641000# diff_83000_3098000# GND efet w=148500 l=8500
+ ad=1.868e+09 pd=370000 as=0 ps=0 
M5195 diff_4808000_2269000# diff_4727000_2238000# diff_4786000_2230000# GND efet w=126000 l=9000
+ ad=-2.03897e+09 pd=420000 as=0 ps=0 
M5196 diff_4694000_2317000# diff_4705000_2274000# diff_4808000_2269000# GND efet w=69000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5197 diff_95000_5192000# diff_4871000_2311000# diff_4871000_2311000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=-1.44797e+09 ps=464000 
M5198 diff_83000_3098000# diff_3408000_4288000# diff_5187000_2412000# GND efet w=103000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5199 diff_95000_5192000# diff_5122000_2495000# diff_5122000_2495000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=-1.22297e+09 ps=570000 
M5200 diff_95000_5192000# diff_4932000_827000# diff_5142000_2400000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=1.09603e+09 ps=1.018e+06 
M5201 diff_83000_3098000# diff_5122000_2495000# diff_5142000_2400000# GND efet w=163500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5202 diff_5122000_2495000# diff_5114000_2490000# diff_83000_3098000# GND efet w=65000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5203 diff_83000_3098000# diff_4932000_827000# diff_5122000_2495000# GND efet w=91500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5204 diff_83000_3098000# diff_4705000_2274000# diff_4871000_2311000# GND efet w=51000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5205 diff_4871000_2311000# diff_4839000_2618000# diff_83000_3098000# GND efet w=61000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5206 diff_4694000_2317000# diff_4705000_2274000# diff_4808000_2269000# GND efet w=68500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5207 diff_4705000_2151000# diff_4602000_2752000# diff_4518000_2032000# GND efet w=20000 l=12000
+ ad=4.65e+08 pd=136000 as=0 ps=0 
M5208 diff_4808000_2269000# diff_4727000_2238000# diff_4786000_2230000# GND efet w=12000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5209 diff_83000_3098000# diff_4839000_2618000# diff_4694000_2317000# GND efet w=51000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5210 diff_4808000_2024000# diff_4727000_2138000# diff_4786000_2160000# GND efet w=10000 l=8000
+ ad=-2.06697e+09 pd=420000 as=1.943e+09 ps=370000 
M5211 diff_3577000_1888000# diff_4328000_910000# diff_95000_5192000# GND efet w=102000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M5212 diff_4459000_2026000# diff_4417000_952000# diff_4433000_2037000# GND efet w=19000 l=10000
+ ad=-1.63897e+09 pd=560000 as=0 ps=0 
M5213 diff_4433000_2037000# diff_4374000_833000# diff_4285000_1501000# GND efet w=19000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5214 diff_4518000_2032000# diff_4518000_2032000# diff_95000_5192000# GND efet w=12000 l=19000
+ ad=0 pd=0 as=0 ps=0 
M5215 diff_4434000_1906000# diff_4374000_833000# diff_4285000_1501000# GND efet w=19000 l=10000
+ ad=1.541e+09 pd=332000 as=0 ps=0 
M5216 diff_3577000_1746000# diff_4328000_910000# diff_95000_5192000# GND efet w=100000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5217 diff_4459000_1862000# diff_4417000_952000# diff_4434000_1906000# GND efet w=21000 l=9000
+ ad=-7.75967e+08 pd=730000 as=0 ps=0 
M5218 diff_95000_5192000# diff_95000_5192000# diff_3577000_1888000# GND efet w=12000 l=104000
+ ad=0 pd=0 as=0 ps=0 
M5219 diff_95000_5192000# diff_4518000_1950000# diff_4518000_1950000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=2.056e+09 ps=412000 
M5220 diff_4518000_1950000# diff_3577000_1888000# diff_83000_3098000# GND efet w=49000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5221 diff_4433000_2037000# diff_4548000_2725000# diff_4608000_2077000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5222 diff_4705000_2105000# diff_4602000_2752000# diff_4433000_2037000# GND efet w=20000 l=12000
+ ad=3.99e+08 pd=80000 as=0 ps=0 
M5223 diff_83000_3098000# diff_4705000_2151000# diff_4727000_2138000# GND efet w=50000 l=8000
+ ad=0 pd=0 as=1.513e+09 ps=300000 
M5224 diff_4786000_2160000# diff_4740000_2641000# diff_83000_3098000# GND efet w=147500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5225 diff_4459000_2246000# diff_4459000_2246000# diff_95000_5192000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M5226 diff_4608000_2077000# diff_4608000_2077000# diff_95000_5192000# GND efet w=13000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M5227 diff_95000_5192000# diff_4459000_2026000# diff_4459000_2026000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M5228 diff_95000_5192000# diff_4608000_1847000# diff_4608000_1847000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=1.792e+09 ps=402000 
M5229 diff_4459000_2026000# diff_4498000_2492000# diff_4434000_1906000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5230 diff_4693000_2058000# diff_4693000_2058000# diff_95000_5192000# GND efet w=13000 l=25000
+ ad=-1.27797e+09 pd=540000 as=0 ps=0 
M5231 diff_4727000_2138000# diff_4727000_2138000# diff_95000_5192000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M5232 diff_4808000_2024000# diff_4727000_2138000# diff_4786000_2160000# GND efet w=125000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5233 diff_4693000_2058000# diff_4705000_2105000# diff_4808000_2024000# GND efet w=66500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5234 diff_83000_3098000# diff_4727000_2238000# diff_4871000_2311000# GND efet w=58000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5235 diff_4950000_2236000# diff_4705000_2274000# diff_83000_3098000# GND efet w=134000 l=8000
+ ad=1.474e+09 pd=290000 as=0 ps=0 
M5236 diff_4970000_2236000# diff_4768000_996000# diff_4950000_2236000# GND efet w=134000 l=9000
+ ad=1.818e+09 pd=352000 as=0 ps=0 
M5237 diff_4990000_2211000# diff_4727000_2238000# diff_4970000_2236000# GND efet w=95000 l=7000
+ ad=-2.80967e+08 pd=692000 as=0 ps=0 
M5238 diff_5271000_2493000# diff_5265000_2778000# diff_83000_3098000# GND efet w=245500 l=8500
+ ad=2.59033e+08 pd=874000 as=0 ps=0 
M5239 diff_95000_5192000# diff_5271000_2493000# diff_5271000_2493000# GND efet w=17000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5240 diff_5011000_576000# diff_5011000_576000# diff_95000_5192000# GND efet w=22000 l=7000
+ ad=4.54065e+08 pd=1.334e+06 as=0 ps=0 
M5241 diff_83000_3098000# diff_72000_4515000# diff_5271000_2493000# GND efet w=202500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5242 diff_83000_3098000# diff_3043000_2723000# diff_5187000_2412000# GND efet w=104000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5243 diff_5011000_576000# diff_72000_4515000# diff_83000_3098000# GND efet w=256000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5244 diff_83000_3098000# diff_5318000_2778000# diff_5011000_576000# GND efet w=125000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5245 diff_5011000_576000# diff_5318000_2778000# diff_83000_3098000# GND efet w=153000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M5246 diff_83000_3098000# diff_5187000_2412000# diff_817000_2342000# GND efet w=89500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5247 diff_6213000_3183000# diff_3569000_3530000# diff_83000_3098000# GND efet w=92500 l=8500
+ ad=-1.44697e+09 pd=502000 as=0 ps=0 
M5248 diff_83000_3098000# diff_4241000_2640000# diff_6213000_3183000# GND efet w=92000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5249 diff_6252000_3157000# diff_5098000_4894000# diff_6213000_3183000# GND efet w=91500 l=8500
+ ad=-1.03797e+09 pd=600000 as=0 ps=0 
M5250 diff_83000_3098000# diff_5009000_4962000# diff_5988000_3969000# GND efet w=41000 l=9000
+ ad=0 pd=0 as=-2.13297e+09 ps=440000 
M5251 diff_6213000_3183000# diff_3408000_4288000# diff_6252000_3157000# GND efet w=86000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5252 diff_5988000_3969000# diff_5068000_4962000# diff_83000_3098000# GND efet w=41000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5253 diff_83000_3098000# diff_5039000_4962000# diff_5988000_3969000# GND efet w=41000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5254 diff_95000_5192000# diff_6252000_3157000# diff_6252000_3157000# GND efet w=13000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M5255 diff_5988000_3969000# diff_5988000_3969000# diff_95000_5192000# GND efet w=13000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M5256 diff_5626000_2884000# diff_5619000_2893000# diff_83000_3098000# GND efet w=156000 l=10000
+ ad=-2.03797e+09 pd=400000 as=0 ps=0 
M5257 diff_5626000_2884000# diff_72000_4515000# diff_5618000_2718000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=1.045e+09 ps=234000 
M5258 diff_5769000_2821000# diff_5087000_472000# diff_83000_3098000# GND efet w=484000 l=9000
+ ad=1.27107e+09 pd=1.608e+06 as=0 ps=0 
M5259 diff_95000_5192000# diff_5626000_2884000# diff_5626000_2884000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5260 diff_95000_5192000# diff_5769000_2821000# diff_5619000_2893000# GND efet w=731000 l=8000
+ ad=0 pd=0 as=-2.64026e+06 ps=6.908e+06 
M5261 diff_95000_5192000# diff_5651000_2807000# diff_5618000_2718000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5262 diff_5651000_2807000# diff_5632000_2727000# diff_83000_3098000# GND efet w=46500 l=7500
+ ad=1.134e+09 pd=212000 as=0 ps=0 
M5263 diff_95000_5192000# diff_5769000_2821000# diff_5619000_2893000# GND efet w=287000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5264 diff_83000_3098000# diff_83000_3098000# diff_5619000_2893000# GND efet w=80000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M5265 diff_5619000_2172000# diff_83000_3098000# diff_83000_3098000# GND efet w=80000 l=12000
+ ad=-1.27161e+09 pd=7.502e+06 as=0 ps=0 
M5266 diff_5769000_2821000# diff_5697000_2542000# diff_83000_3098000# GND efet w=478000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5267 diff_95000_5192000# diff_5651000_2807000# diff_5651000_2807000# GND efet w=11000 l=35000
+ ad=0 pd=0 as=0 ps=0 
M5268 diff_95000_5192000# diff_5769000_2821000# diff_5619000_2893000# GND efet w=285500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5269 diff_5651000_2807000# diff_72000_4515000# diff_83000_3098000# GND efet w=27000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5270 diff_5632000_2727000# diff_5618000_2718000# diff_83000_3098000# GND efet w=222500 l=8500
+ ad=-5.59967e+08 pd=726000 as=0 ps=0 
M5271 diff_95000_5192000# diff_5632000_2727000# diff_5632000_2727000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M5272 diff_5619000_2893000# diff_5769000_2821000# diff_95000_5192000# GND efet w=287500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5273 diff_5769000_2821000# diff_5769000_2821000# diff_95000_5192000# GND efet w=44000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5274 diff_95000_5192000# diff_5697000_2542000# diff_5697000_2542000# GND efet w=33000 l=8000
+ ad=0 pd=0 as=2.02107e+09 ps=1.772e+06 
M5275 diff_83000_3098000# diff_5697000_2542000# diff_5619000_2893000# GND efet w=238500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5276 diff_5697000_2542000# diff_5087000_472000# diff_83000_3098000# GND efet w=476500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5277 diff_5632000_2727000# diff_5011000_576000# diff_817000_2342000# GND efet w=87000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5278 diff_83000_3098000# diff_5651000_2541000# diff_5697000_2542000# GND efet w=513500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5279 diff_95000_5192000# diff_4990000_2211000# diff_4990000_2211000# GND efet w=13000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M5280 diff_5123000_2369000# diff_4932000_827000# diff_95000_5192000# GND efet w=12000 l=8000
+ ad=-3.79673e+07 pd=890000 as=0 ps=0 
M5281 diff_5142000_2400000# diff_4990000_2211000# diff_5123000_2369000# GND efet w=129000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5282 diff_95000_5192000# diff_5069000_2349000# diff_5069000_2349000# GND efet w=13000 l=20000
+ ad=0 pd=0 as=1.675e+09 ps=364000 
M5283 diff_83000_3098000# diff_4727000_2138000# diff_4870000_2082000# GND efet w=59000 l=8000
+ ad=0 pd=0 as=-1.34397e+09 ps=476000 
M5284 diff_83000_3098000# diff_4839000_2618000# diff_4693000_2058000# GND efet w=49000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5285 diff_4990000_2211000# diff_4727000_2238000# diff_4970000_2236000# GND efet w=33000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M5286 diff_83000_3098000# diff_4994000_2634000# diff_4990000_2211000# GND efet w=55000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5287 diff_4990000_2211000# diff_4871000_2311000# diff_83000_3098000# GND efet w=44000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M5288 diff_5123000_2369000# diff_5069000_2349000# diff_83000_3098000# GND efet w=90000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5289 diff_5069000_2349000# diff_4694000_2317000# diff_83000_3098000# GND efet w=65500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5290 diff_83000_3098000# diff_4932000_827000# diff_5069000_2349000# GND efet w=65000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5291 diff_5243000_2360000# diff_5243000_2360000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=2.14e+09 pd=498000 as=0 ps=0 
M5292 diff_5288000_2302000# diff_4990000_2211000# diff_5243000_2360000# GND efet w=77500 l=8500
+ ad=1.377e+09 pd=336000 as=0 ps=0 
M5293 diff_95000_5192000# diff_5202000_2342000# diff_5202000_2342000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=1.634e+09 ps=352000 
M5294 diff_4693000_2058000# diff_4705000_2105000# diff_4808000_2024000# GND efet w=68000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5295 diff_4870000_2082000# diff_4839000_2618000# diff_83000_3098000# GND efet w=57500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5296 diff_95000_5192000# diff_4694000_1940000# diff_4694000_1940000# GND efet w=13000 l=25000
+ ad=0 pd=0 as=-1.18997e+09 ps=546000 
M5297 diff_95000_5192000# diff_4727000_1861000# diff_4727000_1861000# GND efet w=13000 l=24000
+ ad=0 pd=0 as=1.497e+09 ps=296000 
M5298 diff_4253000_1284000# diff_4226000_1649000# diff_83000_3098000# GND efet w=51500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5299 diff_3846000_1323000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5300 diff_3939000_1303000# diff_95000_5192000# diff_3846000_1323000# GND efet w=12500 l=78500
+ ad=8.14e+08 pd=238000 as=0 ps=0 
M5301 diff_3902000_1418000# diff_95000_5192000# diff_95000_5192000# GND efet w=13000 l=31000
+ ad=0 pd=0 as=0 ps=0 
M5302 diff_817000_1286000# diff_3922000_786000# diff_3939000_1303000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5303 diff_4036000_1297000# diff_4004000_2725000# diff_817000_1286000# GND efet w=20000 l=10000
+ ad=8.53e+08 pd=226000 as=0 ps=0 
M5304 diff_95000_5192000# diff_95000_5192000# diff_3846000_1128000# GND efet w=11000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5305 diff_3938000_1186000# diff_95000_5192000# diff_3846000_1128000# GND efet w=12000 l=74000
+ ad=8.01e+08 pd=252000 as=0 ps=0 
M5306 diff_95000_5192000# diff_95000_5192000# diff_3902000_1074000# GND efet w=13000 l=33000
+ ad=0 pd=0 as=1.025e+09 ps=192000 
M5307 diff_4057000_1397000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=31000
+ ad=0 pd=0 as=0 ps=0 
M5308 diff_4066000_1405000# diff_95000_5192000# diff_4036000_1297000# GND efet w=12000 l=79000
+ ad=0 pd=0 as=0 ps=0 
M5309 diff_4066000_1405000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5310 diff_3696000_1028000# diff_3687000_935000# diff_83000_3098000# GND efet w=204000 l=8000
+ ad=-2.73967e+08 pd=706000 as=0 ps=0 
M5311 diff_3687000_935000# diff_3631000_947000# diff_83000_3098000# GND efet w=70500 l=8500
+ ad=9.78e+08 pd=200000 as=0 ps=0 
M5312 diff_3577000_991000# diff_3739000_826000# diff_3696000_1028000# GND efet w=87000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5313 diff_3846000_1128000# diff_3695000_2725000# diff_3577000_1134000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5314 diff_817000_1211000# diff_3922000_786000# diff_3938000_1186000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5315 diff_4036000_1196000# diff_4004000_2725000# diff_817000_1211000# GND efet w=20000 l=10000
+ ad=8.45e+08 pd=234000 as=0 ps=0 
M5316 diff_95000_5192000# diff_95000_5192000# diff_4057000_1091000# GND efet w=13000 l=33000
+ ad=0 pd=0 as=9.68e+08 ps=188000 
M5317 diff_4066000_1098000# diff_95000_5192000# diff_4036000_1196000# GND efet w=12000 l=74000
+ ad=-2.65967e+08 pd=692000 as=0 ps=0 
M5318 diff_3577000_1368000# diff_3749000_2434000# diff_4066000_1405000# GND efet w=87000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5319 diff_95000_5192000# diff_95000_5192000# diff_4066000_1098000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5320 diff_83000_3098000# diff_3902000_1074000# diff_3846000_1128000# GND efet w=203000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5321 diff_3902000_1074000# diff_3938000_1186000# diff_83000_3098000# GND efet w=62000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5322 diff_817000_909000# diff_3489000_2725000# diff_3631000_947000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5323 diff_3687000_935000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=33000
+ ad=0 pd=0 as=0 ps=0 
M5324 diff_3696000_1028000# diff_95000_5192000# diff_3631000_947000# GND efet w=12500 l=80500
+ ad=0 pd=0 as=0 ps=0 
M5325 diff_3696000_1028000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5326 diff_3474000_792000# diff_72000_4515000# diff_83000_3098000# GND efet w=78000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5327 diff_3439000_2492000# diff_72000_4515000# diff_83000_3098000# GND efet w=74000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5328 diff_817000_909000# diff_3800000_830000# diff_3696000_1028000# GND efet w=101500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5329 diff_3846000_946000# diff_3830000_787000# diff_817000_909000# GND efet w=101000 l=10000
+ ad=-2.12967e+08 pd=710000 as=0 ps=0 
M5330 diff_3846000_946000# diff_3695000_2725000# diff_3577000_991000# GND efet w=87000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5331 diff_83000_3098000# diff_3902000_1041000# diff_3846000_946000# GND efet w=205000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5332 diff_3902000_1041000# diff_3939000_927000# diff_83000_3098000# GND efet w=63500 l=7500
+ ad=1.015e+09 pd=192000 as=0 ps=0 
M5333 diff_4057000_1091000# diff_4036000_1196000# diff_83000_3098000# GND efet w=60000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5334 diff_4066000_1098000# diff_4057000_1091000# diff_83000_3098000# GND efet w=202500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5335 diff_817000_1211000# diff_4108000_2725000# diff_4066000_1098000# GND efet w=86000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5336 diff_3577000_1134000# diff_3749000_2434000# diff_4066000_1098000# GND efet w=85000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5337 diff_4241000_1304000# diff_4066000_1475000# diff_83000_3098000# GND efet w=108000 l=9000
+ ad=1.406e+09 pd=304000 as=0 ps=0 
M5338 diff_4261000_1288000# diff_4253000_1284000# diff_4241000_1304000# GND efet w=28000 l=9000
+ ad=1.48203e+09 pd=876000 as=0 ps=0 
M5339 diff_4261000_1288000# diff_4253000_1284000# diff_4241000_1304000# GND efet w=78000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5340 diff_83000_3098000# diff_4066000_1405000# diff_4261000_1288000# GND efet w=72000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5341 diff_3577000_1511000# diff_4328000_910000# diff_95000_5192000# GND efet w=99000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5342 diff_3577000_1746000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=103000
+ ad=0 pd=0 as=0 ps=0 
M5343 diff_4518000_1655000# diff_3577000_1746000# diff_83000_3098000# GND efet w=49000 l=8000
+ ad=1.977e+09 pd=410000 as=0 ps=0 
M5344 diff_83000_3098000# diff_4608000_1847000# diff_4459000_2026000# GND efet w=48000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5345 diff_4608000_1847000# diff_817000_1965000# diff_83000_3098000# GND efet w=66000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5346 diff_4434000_1906000# diff_4548000_2725000# diff_4608000_1847000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5347 diff_4705000_1896000# diff_4602000_2752000# diff_4434000_1906000# GND efet w=21000 l=12000
+ ad=3.99e+08 pd=80000 as=0 ps=0 
M5348 diff_4459000_1862000# diff_4498000_2492000# diff_4430000_1714000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=2.059e+09 ps=440000 
M5349 diff_83000_3098000# diff_4608000_1700000# diff_4459000_1862000# GND efet w=49000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5350 diff_4608000_1700000# diff_817000_1663000# diff_83000_3098000# GND efet w=67000 l=8000
+ ad=1.775e+09 pd=404000 as=0 ps=0 
M5351 diff_4705000_1851000# diff_4602000_2752000# diff_4518000_1950000# GND efet w=21000 l=12000
+ ad=4.67e+08 pd=138000 as=0 ps=0 
M5352 diff_83000_3098000# diff_4705000_1851000# diff_4727000_1861000# GND efet w=49000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5353 diff_4786000_1853000# diff_4740000_2641000# diff_83000_3098000# GND efet w=148500 l=8500
+ ad=1.87e+09 pd=370000 as=0 ps=0 
M5354 diff_4808000_1891000# diff_4727000_1861000# diff_4786000_1853000# GND efet w=126000 l=9000
+ ad=-2.03797e+09 pd=420000 as=0 ps=0 
M5355 diff_4694000_1940000# diff_4705000_1896000# diff_4808000_1891000# GND efet w=69000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5356 diff_83000_3098000# diff_4705000_2105000# diff_4870000_2082000# GND efet w=53000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5357 diff_4870000_2082000# diff_4870000_2082000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M5358 diff_4951000_2028000# diff_4705000_2105000# diff_83000_3098000# GND efet w=135000 l=9000
+ ad=1.35e+09 pd=290000 as=0 ps=0 
M5359 diff_4970000_2028000# diff_4768000_996000# diff_4951000_2028000# GND efet w=135000 l=9000
+ ad=1.831e+09 pd=354000 as=0 ps=0 
M5360 diff_4990000_2028000# diff_4727000_2138000# diff_4970000_2028000# GND efet w=32000 l=7000
+ ad=-4.20967e+08 pd=692000 as=0 ps=0 
M5361 diff_5333000_2356000# diff_72000_4515000# diff_5243000_2360000# GND efet w=20000 l=11000
+ ad=2e+08 pd=60000 as=0 ps=0 
M5362 diff_5354000_2356000# diff_4328000_910000# diff_5333000_2356000# GND efet w=20000 l=11000
+ ad=3.26e+08 pd=100000 as=0 ps=0 
M5363 diff_5202000_2342000# diff_5142000_2400000# diff_83000_3098000# GND efet w=77000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5364 diff_5123000_2369000# diff_5069000_2349000# diff_83000_3098000# GND efet w=48000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5365 diff_5123000_2018000# diff_5069000_2032000# diff_83000_3098000# GND efet w=122000 l=9000
+ ad=1.06033e+08 pd=852000 as=0 ps=0 
M5366 diff_4990000_2028000# diff_4727000_2138000# diff_4970000_2028000# GND efet w=97000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M5367 diff_83000_3098000# diff_4994000_2634000# diff_4990000_2028000# GND efet w=53000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5368 diff_4990000_2028000# diff_4870000_2082000# diff_83000_3098000# GND efet w=44000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M5369 diff_5069000_2032000# diff_4693000_2058000# diff_83000_3098000# GND efet w=64500 l=8500
+ ad=1.771e+09 pd=360000 as=0 ps=0 
M5370 diff_83000_3098000# diff_4932000_827000# diff_5069000_2032000# GND efet w=65000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5371 diff_95000_5192000# diff_4871000_1932000# diff_4871000_1932000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=-1.41297e+09 ps=468000 
M5372 diff_83000_3098000# diff_4705000_1896000# diff_4871000_1932000# GND efet w=52000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5373 diff_4871000_1932000# diff_4839000_2618000# diff_83000_3098000# GND efet w=60000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M5374 diff_4694000_1940000# diff_4705000_1896000# diff_4808000_1891000# GND efet w=68500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5375 diff_4705000_1773000# diff_4602000_2752000# diff_4518000_1655000# GND efet w=20000 l=12000
+ ad=4.63e+08 pd=138000 as=0 ps=0 
M5376 diff_4808000_1891000# diff_4727000_1861000# diff_4786000_1853000# GND efet w=12000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5377 diff_83000_3098000# diff_4839000_2618000# diff_4694000_1940000# GND efet w=51000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5378 diff_4808000_1647000# diff_4727000_1761000# diff_4786000_1782000# GND efet w=10000 l=8000
+ ad=-2.04997e+09 pd=420000 as=1.952e+09 ps=370000 
M5379 diff_4459000_1639000# diff_4417000_952000# diff_4430000_1714000# GND efet w=20000 l=10000
+ ad=-1.71097e+09 pd=544000 as=0 ps=0 
M5380 diff_4430000_1714000# diff_4374000_833000# diff_83000_3098000# GND efet w=19000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5381 diff_4518000_1655000# diff_4518000_1655000# diff_95000_5192000# GND efet w=12000 l=19000
+ ad=0 pd=0 as=0 ps=0 
M5382 diff_4434000_1491000# diff_4374000_833000# diff_83000_3098000# GND efet w=19000 l=10000
+ ad=1.463e+09 pd=314000 as=0 ps=0 
M5383 diff_4458000_1491000# diff_4417000_952000# diff_4434000_1491000# GND efet w=19000 l=10000
+ ad=-9.04967e+08 pd=740000 as=0 ps=0 
M5384 diff_95000_5192000# diff_95000_5192000# diff_3577000_1511000# GND efet w=12000 l=105000
+ ad=0 pd=0 as=0 ps=0 
M5385 diff_95000_5192000# diff_4518000_1573000# diff_4518000_1573000# GND efet w=12000 l=19000
+ ad=0 pd=0 as=2.014e+09 ps=412000 
M5386 diff_4518000_1573000# diff_3577000_1511000# diff_83000_3098000# GND efet w=49000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5387 diff_4430000_1714000# diff_4548000_2725000# diff_4608000_1700000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5388 diff_4705000_1728000# diff_4602000_2752000# diff_4430000_1714000# GND efet w=20000 l=12000
+ ad=4e+08 pd=80000 as=0 ps=0 
M5389 diff_83000_3098000# diff_4705000_1773000# diff_4727000_1761000# GND efet w=50000 l=8000
+ ad=0 pd=0 as=1.511e+09 ps=300000 
M5390 diff_4786000_1782000# diff_4740000_2641000# diff_83000_3098000# GND efet w=147500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5391 diff_4459000_1862000# diff_4459000_1862000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M5392 diff_4608000_1700000# diff_4608000_1700000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M5393 diff_95000_5192000# diff_4459000_1639000# diff_4459000_1639000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M5394 diff_95000_5192000# diff_4608000_1471000# diff_4608000_1471000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=1.79e+09 ps=404000 
M5395 diff_4459000_1639000# diff_4498000_2492000# diff_4434000_1491000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5396 diff_4693000_1681000# diff_4693000_1681000# diff_95000_5192000# GND efet w=13000 l=25000
+ ad=-1.27397e+09 pd=540000 as=0 ps=0 
M5397 diff_4727000_1761000# diff_4727000_1761000# diff_95000_5192000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M5398 diff_4808000_1647000# diff_4727000_1761000# diff_4786000_1782000# GND efet w=126000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5399 diff_4693000_1681000# diff_4705000_1728000# diff_4808000_1647000# GND efet w=66500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5400 diff_83000_3098000# diff_4727000_1861000# diff_4871000_1932000# GND efet w=58000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5401 diff_4950000_1859000# diff_4705000_1896000# diff_83000_3098000# GND efet w=135000 l=8000
+ ad=1.485e+09 pd=292000 as=0 ps=0 
M5402 diff_4970000_1859000# diff_4768000_996000# diff_4950000_1859000# GND efet w=135000 l=9000
+ ad=1.831e+09 pd=354000 as=0 ps=0 
M5403 diff_4990000_1834000# diff_4727000_1861000# diff_4970000_1859000# GND efet w=96000 l=7000
+ ad=-2.72967e+08 pd=692000 as=0 ps=0 
M5404 diff_4990000_2028000# diff_4990000_2028000# diff_95000_5192000# GND efet w=13000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M5405 diff_5069000_2032000# diff_5069000_2032000# diff_95000_5192000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M5406 diff_5123000_2369000# diff_4990000_2028000# diff_5123000_2018000# GND efet w=40000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5407 diff_5123000_2018000# diff_5069000_2032000# diff_83000_3098000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5408 diff_5123000_2369000# diff_4990000_2028000# diff_5123000_2018000# GND efet w=70000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5409 diff_83000_3098000# diff_4990000_2211000# diff_5202000_2342000# GND efet w=70500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5410 diff_5243000_2360000# diff_5202000_2342000# diff_83000_3098000# GND efet w=63500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5411 diff_5288000_2302000# diff_4990000_2211000# diff_5243000_2360000# GND efet w=32000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5412 diff_83000_3098000# diff_5142000_2400000# diff_5288000_2302000# GND efet w=115500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5413 diff_5201000_2038000# diff_5123000_2369000# diff_83000_3098000# GND efet w=78000 l=8000
+ ad=1.566e+09 pd=344000 as=0 ps=0 
M5414 diff_83000_3098000# diff_4990000_2028000# diff_5201000_2038000# GND efet w=70500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5415 diff_83000_3098000# diff_5123000_2369000# diff_5288000_2043000# GND efet w=119000 l=8000
+ ad=0 pd=0 as=1.396e+09 ps=338000 
M5416 diff_5243000_2018000# diff_5201000_2038000# diff_83000_3098000# GND efet w=63500 l=8500
+ ad=-1.99497e+09 pd=502000 as=0 ps=0 
M5417 diff_5288000_2043000# diff_4990000_2028000# diff_5243000_2018000# GND efet w=33000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5418 diff_5201000_2038000# diff_5201000_2038000# diff_95000_5192000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M5419 diff_5123000_2018000# diff_4932000_827000# diff_95000_5192000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5420 diff_5288000_2043000# diff_4990000_2028000# diff_5243000_2018000# GND efet w=74000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5421 diff_95000_5192000# diff_5375000_2327000# diff_5375000_2327000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=-1.54797e+09 ps=536000 
M5422 diff_5375000_2327000# diff_5354000_2356000# diff_83000_3098000# GND efet w=190000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5423 diff_5331000_4062000# diff_5375000_2327000# diff_83000_3098000# GND efet w=155500 l=7500
+ ad=-2.14284e+09 pd=3.714e+06 as=0 ps=0 
M5424 diff_817000_2342000# diff_5271000_2493000# diff_5375000_2327000# GND efet w=86500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5425 diff_5375000_2058000# diff_5354000_2022000# diff_83000_3098000# GND efet w=199500 l=8500
+ ad=-1.50297e+09 pd=518000 as=0 ps=0 
M5426 diff_5331000_4062000# diff_5375000_2058000# diff_83000_3098000# GND efet w=154500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5427 diff_5243000_2018000# diff_5243000_2018000# diff_95000_5192000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M5428 diff_5334000_2022000# diff_72000_4515000# diff_5243000_2018000# GND efet w=19000 l=12000
+ ad=1.52e+08 pd=54000 as=0 ps=0 
M5429 diff_5354000_2022000# diff_4328000_910000# diff_5334000_2022000# GND efet w=19000 l=12000
+ ad=3.38e+08 pd=90000 as=0 ps=0 
M5430 diff_5375000_2058000# diff_5375000_2058000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M5431 diff_817000_2040000# diff_5271000_2493000# diff_5375000_2058000# GND efet w=86500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5432 diff_817000_2342000# diff_4954000_639000# diff_5651000_2541000# GND efet w=35000 l=12000
+ ad=0 pd=0 as=-1.58597e+09 ps=322000 
M5433 diff_83000_3098000# diff_5697000_2542000# diff_5619000_2893000# GND efet w=289000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5434 diff_83000_3098000# diff_5697000_2542000# diff_5619000_2893000# GND efet w=289500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5435 diff_5619000_2893000# diff_5697000_2542000# diff_83000_3098000# GND efet w=800500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5436 diff_5696000_2524000# diff_5651000_2472000# diff_83000_3098000# GND efet w=516000 l=9000
+ ad=1.58607e+09 pd=1.788e+06 as=0 ps=0 
M5437 diff_83000_3098000# diff_5696000_2524000# diff_5619000_2172000# GND efet w=795500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5438 diff_83000_3098000# diff_5087000_472000# diff_5696000_2524000# GND efet w=474000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5439 diff_5651000_2472000# diff_4954000_639000# diff_817000_2040000# GND efet w=35000 l=11000
+ ad=-1.70097e+09 pd=296000 as=0 ps=0 
M5440 diff_817000_2040000# diff_5011000_576000# diff_5632000_2276000# GND efet w=87000 l=10000
+ ad=0 pd=0 as=-2.52967e+08 ps=744000 
M5441 diff_5632000_2276000# diff_5618000_2219000# diff_83000_3098000# GND efet w=221000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5442 diff_83000_3098000# diff_5696000_2524000# diff_5619000_2172000# GND efet w=289500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5443 diff_83000_3098000# diff_5696000_2524000# diff_5619000_2172000# GND efet w=289000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5444 diff_5619000_2172000# diff_5696000_2524000# diff_83000_3098000# GND efet w=238500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5445 diff_5696000_2524000# diff_5696000_2524000# diff_5696000_2524000# GND efet w=2000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M5446 diff_5696000_2524000# diff_5696000_2524000# diff_95000_5192000# GND efet w=36000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5447 diff_95000_5192000# diff_4990000_1834000# diff_4990000_1834000# GND efet w=13000 l=26000
+ ad=0 pd=0 as=0 ps=0 
M5448 diff_5123000_1992000# diff_4932000_827000# diff_95000_5192000# GND efet w=12000 l=8000
+ ad=-1.59673e+07 pd=892000 as=0 ps=0 
M5449 diff_5123000_2018000# diff_4990000_1834000# diff_5123000_1992000# GND efet w=128500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5450 diff_95000_5192000# diff_5069000_1972000# diff_5069000_1972000# GND efet w=13000 l=20000
+ ad=0 pd=0 as=1.612e+09 ps=362000 
M5451 diff_83000_3098000# diff_4727000_1761000# diff_4870000_1705000# GND efet w=59000 l=8000
+ ad=0 pd=0 as=-1.29097e+09 ps=476000 
M5452 diff_83000_3098000# diff_4839000_2618000# diff_4693000_1681000# GND efet w=50000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5453 diff_4990000_1834000# diff_4727000_1861000# diff_4970000_1859000# GND efet w=33000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M5454 diff_83000_3098000# diff_4994000_2634000# diff_4990000_1834000# GND efet w=55000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5455 diff_4990000_1834000# diff_4871000_1932000# diff_83000_3098000# GND efet w=44000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M5456 diff_5123000_1992000# diff_5069000_1972000# diff_83000_3098000# GND efet w=89500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5457 diff_5069000_1972000# diff_4694000_1940000# diff_83000_3098000# GND efet w=65500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5458 diff_83000_3098000# diff_4932000_827000# diff_5069000_1972000# GND efet w=66000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5459 diff_5243000_1983000# diff_5243000_1983000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=-2.12097e+09 pd=500000 as=0 ps=0 
M5460 diff_95000_5192000# diff_5202000_1964000# diff_5202000_1964000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=1.62e+09 ps=350000 
M5461 diff_5288000_1925000# diff_4990000_1834000# diff_5243000_1983000# GND efet w=76500 l=8500
+ ad=1.367e+09 pd=334000 as=0 ps=0 
M5462 diff_4693000_1681000# diff_4705000_1728000# diff_4808000_1647000# GND efet w=68000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5463 diff_4870000_1705000# diff_4839000_2618000# diff_83000_3098000# GND efet w=58500 l=6500
+ ad=0 pd=0 as=0 ps=0 
M5464 diff_95000_5192000# diff_4694000_1563000# diff_4694000_1563000# GND efet w=13000 l=24000
+ ad=0 pd=0 as=-1.19997e+09 ps=548000 
M5465 diff_95000_5192000# diff_4727000_1483000# diff_4727000_1483000# GND efet w=13000 l=24000
+ ad=0 pd=0 as=1.539e+09 ps=300000 
M5466 diff_3577000_1368000# diff_4328000_910000# diff_95000_5192000# GND efet w=102000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5467 diff_4318000_999000# diff_3408000_4288000# diff_83000_3098000# GND efet w=52500 l=8500
+ ad=6.95e+08 pd=148000 as=0 ps=0 
M5468 diff_83000_3098000# diff_4066000_1098000# diff_4261000_1288000# GND efet w=83000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5469 diff_95000_5192000# diff_4225000_1221000# diff_4225000_1221000# GND efet w=12000 l=35000
+ ad=0 pd=0 as=-1.60197e+09 ps=390000 
M5470 diff_4318000_999000# diff_4318000_999000# diff_95000_5192000# GND efet w=12000 l=37000
+ ad=0 pd=0 as=0 ps=0 
M5471 diff_95000_5192000# diff_4307000_1187000# diff_4307000_1187000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=-6.24967e+08 ps=698000 
M5472 diff_4066000_1028000# diff_4057000_1020000# diff_83000_3098000# GND efet w=204500 l=7500
+ ad=-4.87967e+08 pd=686000 as=0 ps=0 
M5473 diff_83000_3098000# diff_4036000_920000# diff_4057000_1020000# GND efet w=61000 l=8000
+ ad=0 pd=0 as=9.53e+08 ps=184000 
M5474 diff_817000_909000# diff_4108000_2725000# diff_4066000_1028000# GND efet w=87000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5475 diff_83000_3098000# diff_3901000_2725000# diff_3577000_1134000# GND efet w=105000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5476 diff_83000_3098000# diff_3901000_2725000# diff_3577000_991000# GND efet w=104500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5477 diff_4261000_1288000# diff_4066000_1028000# diff_4225000_1221000# GND efet w=109000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5478 diff_3846000_946000# diff_95000_5192000# diff_95000_5192000# GND efet w=11000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5479 diff_3939000_927000# diff_95000_5192000# diff_3846000_946000# GND efet w=11500 l=80500
+ ad=7.78e+08 pd=238000 as=0 ps=0 
M5480 diff_83000_3098000# diff_72000_4515000# diff_3567000_785000# GND efet w=70000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5481 diff_3596000_2395000# diff_72000_4515000# diff_83000_3098000# GND efet w=93500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5482 diff_83000_3098000# diff_72000_4515000# diff_3354000_2409000# GND efet w=70000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5483 diff_3489000_2725000# diff_72000_4515000# diff_83000_3098000# GND efet w=70000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5484 diff_83000_3098000# diff_72000_4515000# diff_3739000_826000# GND efet w=77000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5485 diff_3800000_830000# diff_72000_4515000# diff_83000_3098000# GND efet w=74000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5486 diff_3902000_1041000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=33000
+ ad=0 pd=0 as=0 ps=0 
M5487 diff_817000_909000# diff_3922000_786000# diff_3939000_927000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5488 diff_4036000_920000# diff_4004000_2725000# diff_817000_909000# GND efet w=20000 l=10000
+ ad=8.45e+08 pd=228000 as=0 ps=0 
M5489 diff_4057000_1020000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=33000
+ ad=0 pd=0 as=0 ps=0 
M5490 diff_4066000_1028000# diff_95000_5192000# diff_4036000_920000# GND efet w=12000 l=81000
+ ad=0 pd=0 as=0 ps=0 
M5491 diff_4066000_1028000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5492 diff_83000_3098000# diff_72000_4515000# diff_3830000_787000# GND efet w=70000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5493 diff_3695000_2725000# diff_72000_4515000# diff_83000_3098000# GND efet w=96500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5494 diff_3577000_991000# diff_3749000_2434000# diff_4066000_1028000# GND efet w=86000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5495 diff_4307000_1010000# diff_4225000_1221000# diff_83000_3098000# GND efet w=101000 l=8000
+ ad=1.111e+09 pd=224000 as=0 ps=0 
M5496 diff_4307000_1187000# diff_4318000_999000# diff_4307000_1010000# GND efet w=101000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5497 diff_3577000_1368000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=104000
+ ad=0 pd=0 as=0 ps=0 
M5498 diff_4518000_1278000# diff_3577000_1368000# diff_83000_3098000# GND efet w=49000 l=8000
+ ad=1.99e+09 pd=410000 as=0 ps=0 
M5499 diff_83000_3098000# diff_4608000_1471000# diff_4459000_1639000# GND efet w=48000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5500 diff_4608000_1471000# diff_817000_1588000# diff_83000_3098000# GND efet w=66000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5501 diff_4434000_1491000# diff_4548000_2725000# diff_4608000_1471000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5502 diff_4705000_1519000# diff_4602000_2752000# diff_4434000_1491000# GND efet w=21000 l=12000
+ ad=3.99e+08 pd=80000 as=0 ps=0 
M5503 diff_4458000_1491000# diff_4498000_2492000# diff_4432000_1237000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=-2.13097e+09 ps=466000 
M5504 diff_83000_3098000# diff_4608000_1323000# diff_4458000_1491000# GND efet w=50000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5505 diff_4608000_1323000# diff_817000_1286000# diff_83000_3098000# GND efet w=67000 l=8000
+ ad=1.768e+09 pd=402000 as=0 ps=0 
M5506 diff_4705000_1475000# diff_4602000_2752000# diff_4518000_1573000# GND efet w=20000 l=12000
+ ad=4.73e+08 pd=138000 as=0 ps=0 
M5507 diff_83000_3098000# diff_4705000_1475000# diff_4727000_1483000# GND efet w=50000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5508 diff_4786000_1476000# diff_4740000_2641000# diff_83000_3098000# GND efet w=148500 l=8500
+ ad=1.868e+09 pd=370000 as=0 ps=0 
M5509 diff_4808000_1515000# diff_4727000_1483000# diff_4786000_1476000# GND efet w=126000 l=9000
+ ad=-2.03897e+09 pd=420000 as=0 ps=0 
M5510 diff_4694000_1563000# diff_4705000_1519000# diff_4808000_1515000# GND efet w=69000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5511 diff_83000_3098000# diff_4705000_1728000# diff_4870000_1705000# GND efet w=53000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5512 diff_4870000_1705000# diff_4870000_1705000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M5513 diff_4951000_1651000# diff_4705000_1728000# diff_83000_3098000# GND efet w=135000 l=9000
+ ad=1.35e+09 pd=290000 as=0 ps=0 
M5514 diff_4970000_1651000# diff_4768000_996000# diff_4951000_1651000# GND efet w=135000 l=9000
+ ad=1.831e+09 pd=354000 as=0 ps=0 
M5515 diff_4990000_1651000# diff_4727000_1761000# diff_4970000_1651000# GND efet w=32000 l=7000
+ ad=-4.25967e+08 pd=692000 as=0 ps=0 
M5516 diff_5334000_1978000# diff_72000_4515000# diff_5243000_1983000# GND efet w=21000 l=12000
+ ad=1.68e+08 pd=58000 as=0 ps=0 
M5517 diff_5354000_1978000# diff_4328000_910000# diff_5334000_1978000# GND efet w=21000 l=12000
+ ad=3.38e+08 pd=104000 as=0 ps=0 
M5518 diff_5123000_1992000# diff_5069000_1972000# diff_83000_3098000# GND efet w=48000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5519 diff_5202000_1964000# diff_5123000_2018000# diff_83000_3098000# GND efet w=77000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5520 diff_4990000_1651000# diff_4727000_1761000# diff_4970000_1651000# GND efet w=97000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M5521 diff_83000_3098000# diff_4994000_2634000# diff_4990000_1651000# GND efet w=54000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5522 diff_4990000_1651000# diff_4870000_1705000# diff_83000_3098000# GND efet w=45000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M5523 diff_5069000_1655000# diff_4693000_1681000# diff_83000_3098000# GND efet w=64500 l=8500
+ ad=1.74e+09 pd=362000 as=0 ps=0 
M5524 diff_83000_3098000# diff_4932000_827000# diff_5069000_1655000# GND efet w=65500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5525 diff_5123000_1641000# diff_5069000_1655000# diff_83000_3098000# GND efet w=123000 l=9000
+ ad=-1.65797e+09 pd=512000 as=0 ps=0 
M5526 diff_95000_5192000# diff_4871000_1557000# diff_4871000_1557000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=-1.44597e+09 ps=462000 
M5527 diff_83000_3098000# diff_4705000_1519000# diff_4871000_1557000# GND efet w=51000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5528 diff_4871000_1557000# diff_4839000_2618000# diff_83000_3098000# GND efet w=61500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5529 diff_4694000_1563000# diff_4705000_1519000# diff_4808000_1515000# GND efet w=68500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5530 diff_4705000_1396000# diff_4602000_2752000# diff_4518000_1278000# GND efet w=21000 l=12000
+ ad=4.78e+08 pd=138000 as=0 ps=0 
M5531 diff_4808000_1515000# diff_4727000_1483000# diff_4786000_1476000# GND efet w=12000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5532 diff_83000_3098000# diff_4839000_2618000# diff_4694000_1563000# GND efet w=51000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5533 diff_4808000_1269000# diff_4727000_1383000# diff_4786000_1406000# GND efet w=10000 l=8000
+ ad=-2.12197e+09 pd=420000 as=1.815e+09 ps=372000 
M5534 diff_4432000_1237000# diff_4374000_833000# diff_4307000_1187000# GND efet w=20000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5535 diff_4459000_1183000# diff_4417000_952000# diff_4432000_1237000# GND efet w=20000 l=10000
+ ad=-1.86197e+09 pd=486000 as=0 ps=0 
M5536 diff_3577000_1134000# diff_4328000_910000# diff_95000_5192000# GND efet w=100500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5537 diff_4518000_1278000# diff_4518000_1278000# diff_95000_5192000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M5538 diff_4432000_1144000# diff_4374000_833000# diff_4307000_1187000# GND efet w=21000 l=9000
+ ad=1.614e+09 pd=326000 as=0 ps=0 
M5539 diff_3577000_991000# diff_4328000_910000# diff_95000_5192000# GND efet w=87000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5540 diff_1758000_613000# diff_1758000_613000# diff_95000_5192000# GND efet w=16000 l=8000
+ ad=-4.84967e+08 pd=636000 as=0 ps=0 
M5541 diff_83000_3098000# diff_1757000_739000# diff_1758000_613000# GND efet w=231000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5542 diff_1694000_585000# diff_1694000_585000# diff_95000_5192000# GND efet w=50500 l=7500
+ ad=-8.69019e+07 pd=1.982e+06 as=0 ps=0 
M5543 diff_83000_3098000# diff_1844000_568000# diff_1694000_585000# GND efet w=485500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5544 diff_1844000_568000# diff_680000_1019000# diff_1758000_613000# GND efet w=35000 l=11000
+ ad=7.6e+08 pd=180000 as=0 ps=0 
M5545 diff_95000_5192000# diff_1620000_123000# diff_1620000_123000# GND efet w=36000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5546 diff_83000_3098000# diff_553000_1211000# diff_1694000_585000# GND efet w=437000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5547 diff_1620000_123000# diff_1694000_585000# diff_83000_3098000# GND efet w=44000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5548 diff_83000_3098000# diff_2108000_568000# diff_2035000_545000# GND efet w=487500 l=8500
+ ad=0 pd=0 as=-1.92902e+08 ps=1.988e+06 
M5549 diff_83000_3098000# diff_553000_1211000# diff_2035000_545000# GND efet w=437000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5550 diff_95000_5192000# diff_2035000_545000# diff_2035000_545000# GND efet w=52500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5551 diff_83000_3098000# diff_1774000_760000# diff_2214000_625000# GND efet w=231500 l=8500
+ ad=0 pd=0 as=-4.26967e+08 ps=638000 
M5552 diff_95000_5192000# diff_2214000_625000# diff_2214000_625000# GND efet w=16000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5553 diff_2214000_625000# diff_680000_1019000# diff_2108000_568000# GND efet w=35000 l=11000
+ ad=0 pd=0 as=6.82e+08 ps=178000 
M5554 diff_83000_3098000# diff_2035000_545000# diff_2261000_565000# GND efet w=274000 l=8000
+ ad=0 pd=0 as=2.04607e+09 ps=1.492e+06 
M5555 diff_83000_3098000# diff_553000_1211000# diff_2261000_565000# GND efet w=299500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5556 diff_2261000_565000# diff_2035000_545000# diff_83000_3098000# GND efet w=45000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5557 diff_83000_3098000# diff_1430000_565000# diff_1218000_195000# GND efet w=183500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5558 diff_83000_3098000# diff_1430000_565000# diff_1218000_195000# GND efet w=182000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5559 diff_1627000_456000# diff_1620000_123000# diff_83000_3098000# GND efet w=182000 l=8000
+ ad=1.60294e+08 pd=4.552e+06 as=0 ps=0 
M5560 diff_83000_3098000# diff_1430000_565000# diff_1218000_195000# GND efet w=649500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5561 diff_95000_5192000# diff_969000_456000# diff_801000_364000# GND efet w=523000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5562 diff_801000_364000# diff_969000_456000# diff_95000_5192000# GND efet w=260000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5563 diff_1218000_195000# diff_1204000_546000# diff_95000_5192000# GND efet w=268500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5564 diff_83000_3098000# diff_1620000_123000# diff_1627000_456000# GND efet w=184000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5565 diff_1627000_456000# diff_1620000_123000# diff_83000_3098000# GND efet w=647500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5566 diff_83000_3098000# diff_1620000_123000# diff_1627000_456000# GND efet w=191500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5567 diff_95000_5192000# diff_1694000_585000# diff_1627000_456000# GND efet w=208000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5568 diff_95000_5192000# diff_1694000_585000# diff_1627000_456000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5569 diff_95000_5192000# diff_1694000_585000# diff_1627000_456000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5570 diff_95000_5192000# diff_1694000_585000# diff_1627000_456000# GND efet w=189500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5571 diff_2049000_194000# diff_2035000_545000# diff_95000_5192000# GND efet w=191000 l=8000
+ ad=-7.17057e+07 pd=4.558e+06 as=0 ps=0 
M5572 diff_95000_5192000# diff_1694000_585000# diff_1627000_456000# GND efet w=650000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5573 diff_1218000_195000# diff_1430000_565000# diff_83000_3098000# GND efet w=280000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5574 diff_1627000_456000# diff_1620000_123000# diff_83000_3098000# GND efet w=280000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5575 diff_95000_5192000# diff_2035000_545000# diff_2049000_194000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5576 diff_2049000_194000# diff_2035000_545000# diff_95000_5192000# GND efet w=650000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5577 diff_95000_5192000# diff_2035000_545000# diff_2049000_194000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5578 diff_95000_5192000# diff_2035000_545000# diff_2049000_194000# GND efet w=208000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5579 diff_2261000_565000# diff_2261000_565000# diff_95000_5192000# GND efet w=35000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5580 diff_2261000_565000# diff_553000_1211000# diff_83000_3098000# GND efet w=56000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5581 diff_83000_3098000# diff_2261000_565000# diff_2049000_194000# GND efet w=191500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5582 diff_83000_3098000# diff_553000_1211000# diff_2450000_123000# GND efet w=56000 l=8000
+ ad=0 pd=0 as=2.02607e+09 ps=1.488e+06 
M5583 diff_83000_3098000# diff_553000_1211000# diff_2450000_123000# GND efet w=299500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5584 diff_83000_3098000# diff_2524000_585000# diff_2450000_123000# GND efet w=274000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5585 diff_2589000_613000# diff_2589000_613000# diff_95000_5192000# GND efet w=16000 l=8000
+ ad=-6.16967e+08 pd=636000 as=0 ps=0 
M5586 diff_83000_3098000# diff_1791000_798000# diff_2589000_613000# GND efet w=231500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5587 diff_2524000_585000# diff_2524000_585000# diff_95000_5192000# GND efet w=50000 l=8000
+ ad=-1.94902e+08 pd=1.982e+06 as=0 ps=0 
M5588 diff_83000_3098000# diff_2674000_568000# diff_2524000_585000# GND efet w=483500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5589 diff_2674000_568000# diff_680000_1019000# diff_2589000_613000# GND efet w=35000 l=12000
+ ad=6.92e+08 pd=178000 as=0 ps=0 
M5590 diff_95000_5192000# diff_2450000_123000# diff_2450000_123000# GND efet w=34000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5591 diff_83000_3098000# diff_553000_1211000# diff_2524000_585000# GND efet w=439000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5592 diff_2450000_123000# diff_2524000_585000# diff_83000_3098000# GND efet w=45000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5593 diff_83000_3098000# diff_553000_1211000# diff_3258000_123000# GND efet w=56000 l=9000
+ ad=0 pd=0 as=1.79907e+09 ps=1.484e+06 
M5594 diff_83000_3098000# diff_553000_1211000# diff_3258000_123000# GND efet w=302000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5595 diff_83000_3098000# diff_3332000_585000# diff_3258000_123000# GND efet w=272000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5596 diff_83000_3098000# diff_2261000_565000# diff_2049000_194000# GND efet w=184500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5597 diff_83000_3098000# diff_2261000_565000# diff_2049000_194000# GND efet w=181000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5598 diff_2458000_131000# diff_2450000_123000# diff_83000_3098000# GND efet w=183000 l=8000
+ ad=3.58294e+08 pd=4.556e+06 as=0 ps=0 
M5599 diff_83000_3098000# diff_2261000_565000# diff_2049000_194000# GND efet w=646500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5600 diff_83000_3098000# diff_2450000_123000# diff_2458000_131000# GND efet w=184500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5601 diff_2458000_131000# diff_2450000_123000# diff_83000_3098000# GND efet w=648500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5602 diff_83000_3098000# diff_2450000_123000# diff_2458000_131000# GND efet w=191000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5603 diff_95000_5192000# diff_2524000_585000# diff_2458000_131000# GND efet w=208000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5604 diff_95000_5192000# diff_2524000_585000# diff_2458000_131000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5605 diff_95000_5192000# diff_2524000_585000# diff_2458000_131000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5606 diff_95000_5192000# diff_2524000_585000# diff_2458000_131000# GND efet w=189000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5607 diff_95000_5192000# diff_2524000_585000# diff_2458000_131000# GND efet w=646000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5608 diff_1627000_456000# diff_1694000_585000# diff_95000_5192000# GND efet w=269000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5609 diff_2049000_194000# diff_2035000_545000# diff_95000_5192000# GND efet w=270000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5610 diff_2049000_194000# diff_2261000_565000# diff_83000_3098000# GND efet w=280000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5611 diff_2458000_131000# diff_2450000_123000# diff_83000_3098000# GND efet w=281000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5612 diff_83000_3098000# diff_72000_4515000# diff_3922000_786000# GND efet w=102500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5613 diff_4004000_2725000# diff_72000_4515000# diff_83000_3098000# GND efet w=69000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5614 diff_83000_3098000# diff_72000_4515000# diff_4045000_823000# GND efet w=111000 l=8000
+ ad=0 pd=0 as=1.932e+09 ps=304000 
M5615 diff_95000_5192000# diff_4045000_823000# diff_4045000_823000# GND efet w=13000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M5616 diff_4108000_2725000# diff_72000_4515000# diff_83000_3098000# GND efet w=74500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5617 diff_83000_3098000# diff_72000_4515000# diff_3749000_2434000# GND efet w=74000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5618 diff_3901000_2725000# diff_72000_4515000# diff_83000_3098000# GND efet w=75000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5619 diff_4328000_910000# diff_4045000_823000# diff_83000_3098000# GND efet w=72000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5620 diff_4459000_1108000# diff_4417000_952000# diff_4432000_1144000# GND efet w=21000 l=8000
+ ad=-9.55967e+08 pd=728000 as=0 ps=0 
M5621 diff_95000_5192000# diff_95000_5192000# diff_3577000_1134000# GND efet w=12000 l=104000
+ ad=0 pd=0 as=0 ps=0 
M5622 diff_95000_5192000# diff_4518000_1196000# diff_4518000_1196000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=2.049e+09 ps=412000 
M5623 diff_4518000_1196000# diff_3577000_1134000# diff_83000_3098000# GND efet w=49000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5624 diff_4432000_1237000# diff_4548000_2725000# diff_4608000_1323000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5625 diff_4705000_1351000# diff_4602000_2752000# diff_4432000_1237000# GND efet w=20000 l=12000
+ ad=4e+08 pd=80000 as=0 ps=0 
M5626 diff_83000_3098000# diff_4705000_1396000# diff_4727000_1383000# GND efet w=50000 l=8000
+ ad=0 pd=0 as=1.51e+09 ps=300000 
M5627 diff_4786000_1406000# diff_4740000_2641000# diff_83000_3098000# GND efet w=148000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5628 diff_4458000_1491000# diff_4458000_1491000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M5629 diff_4608000_1323000# diff_4608000_1323000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M5630 diff_95000_5192000# diff_4459000_1183000# diff_4459000_1183000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M5631 diff_95000_5192000# diff_4608000_1093000# diff_4608000_1093000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=1.777e+09 ps=400000 
M5632 diff_4459000_1183000# diff_4498000_2492000# diff_4432000_1144000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5633 diff_4693000_1304000# diff_4693000_1304000# diff_95000_5192000# GND efet w=13000 l=25000
+ ad=-1.29497e+09 pd=540000 as=0 ps=0 
M5634 diff_4727000_1383000# diff_4727000_1383000# diff_95000_5192000# GND efet w=14000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M5635 diff_4808000_1269000# diff_4727000_1383000# diff_4786000_1406000# GND efet w=126000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5636 diff_4693000_1304000# diff_4705000_1351000# diff_4808000_1269000# GND efet w=66500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5637 diff_83000_3098000# diff_4727000_1483000# diff_4871000_1557000# GND efet w=58000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5638 diff_4950000_1482000# diff_4705000_1519000# diff_83000_3098000# GND efet w=134000 l=8000
+ ad=1.474e+09 pd=290000 as=0 ps=0 
M5639 diff_4970000_1482000# diff_4768000_996000# diff_4950000_1482000# GND efet w=134000 l=9000
+ ad=1.819e+09 pd=352000 as=0 ps=0 
M5640 diff_4990000_1457000# diff_4727000_1483000# diff_4970000_1482000# GND efet w=95000 l=7000
+ ad=-2.82967e+08 pd=692000 as=0 ps=0 
M5641 diff_4990000_1651000# diff_4990000_1651000# diff_95000_5192000# GND efet w=13000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M5642 diff_5069000_1655000# diff_5069000_1655000# diff_95000_5192000# GND efet w=12000 l=19000
+ ad=0 pd=0 as=0 ps=0 
M5643 diff_5123000_1992000# diff_4990000_1651000# diff_5123000_1641000# GND efet w=41000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5644 diff_5123000_1641000# diff_5069000_1655000# diff_83000_3098000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5645 diff_5123000_1992000# diff_4990000_1651000# diff_5123000_1641000# GND efet w=71000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5646 diff_83000_3098000# diff_4990000_1834000# diff_5202000_1964000# GND efet w=70500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5647 diff_5243000_1983000# diff_5202000_1964000# diff_83000_3098000# GND efet w=63500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5648 diff_5288000_1925000# diff_4990000_1834000# diff_5243000_1983000# GND efet w=32000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5649 diff_83000_3098000# diff_5123000_2018000# diff_5288000_1925000# GND efet w=115500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5650 diff_5201000_1660000# diff_5123000_1992000# diff_83000_3098000# GND efet w=78000 l=8000
+ ad=1.576e+09 pd=346000 as=0 ps=0 
M5651 diff_83000_3098000# diff_4990000_1651000# diff_5201000_1660000# GND efet w=71500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5652 diff_83000_3098000# diff_5123000_1992000# diff_5288000_1666000# GND efet w=118500 l=8500
+ ad=0 pd=0 as=1.383e+09 ps=336000 
M5653 diff_5243000_1641000# diff_5201000_1660000# diff_83000_3098000# GND efet w=63500 l=8500
+ ad=-2.02297e+09 pd=502000 as=0 ps=0 
M5654 diff_5288000_1666000# diff_4990000_1651000# diff_5243000_1641000# GND efet w=33000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5655 diff_5201000_1660000# diff_5201000_1660000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5656 diff_5123000_1641000# diff_4932000_827000# diff_95000_5192000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5657 diff_5288000_1666000# diff_4990000_1651000# diff_5243000_1641000# GND efet w=74500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5658 diff_95000_5192000# diff_5375000_1950000# diff_5375000_1950000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=-1.53997e+09 ps=540000 
M5659 diff_5375000_1950000# diff_5354000_1978000# diff_83000_3098000# GND efet w=191000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5660 diff_5331000_4062000# diff_5375000_1950000# diff_83000_3098000# GND efet w=155500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5661 diff_83000_3098000# diff_5159000_1628000# diff_5170000_2830000# GND efet w=103500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5662 diff_5170000_2830000# diff_5170000_2830000# diff_95000_5192000# GND efet w=12000 l=15000
+ ad=0 pd=0 as=0 ps=0 
M5663 diff_817000_1965000# diff_5271000_2493000# diff_5375000_1950000# GND efet w=88000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5664 diff_95000_5192000# diff_5473000_1600000# diff_5473000_1600000# GND efet w=12000 l=14000
+ ad=0 pd=0 as=1.792e+09 ps=364000 
M5665 diff_5473000_1600000# diff_5473000_1600000# diff_5473000_1600000# GND efet w=1000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5666 diff_5375000_1681000# diff_5354000_1645000# diff_83000_3098000# GND efet w=198000 l=8000
+ ad=-1.49897e+09 pd=520000 as=0 ps=0 
M5667 diff_5331000_4062000# diff_5375000_1681000# diff_83000_3098000# GND efet w=154500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5668 diff_5473000_1600000# diff_5123000_1641000# diff_83000_3098000# GND efet w=96000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5669 diff_95000_5192000# diff_5632000_2276000# diff_5632000_2276000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M5670 diff_83000_3098000# diff_72000_4515000# diff_5651000_2257000# GND efet w=28000 l=9000
+ ad=0 pd=0 as=1.184e+09 ps=216000 
M5671 diff_95000_5192000# diff_5769000_2161000# diff_5769000_2161000# GND efet w=44000 l=9000
+ ad=0 pd=0 as=1.33207e+09 ps=1.612e+06 
M5672 diff_83000_3098000# diff_5696000_2524000# diff_5769000_2161000# GND efet w=478000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5673 diff_5619000_2172000# diff_5769000_2161000# diff_95000_5192000# GND efet w=286000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5674 diff_5632000_2276000# diff_5632000_2276000# diff_5632000_2276000# GND efet w=1000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M5675 diff_95000_5192000# diff_5769000_2161000# diff_5619000_2172000# GND efet w=285500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5676 diff_95000_5192000# diff_5651000_2257000# diff_5651000_2257000# GND efet w=12000 l=35000
+ ad=0 pd=0 as=0 ps=0 
M5677 diff_5651000_2257000# diff_5632000_2276000# diff_83000_3098000# GND efet w=43500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5678 diff_95000_5192000# diff_5651000_2257000# diff_5618000_2219000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=9.4e+08 ps=230000 
M5679 diff_83000_3098000# diff_5087000_472000# diff_5769000_2161000# GND efet w=486000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5680 diff_95000_5192000# diff_5769000_2161000# diff_5619000_2172000# GND efet w=285500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5681 diff_5618000_2219000# diff_72000_4515000# diff_5626000_2182000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=2.098e+09 ps=394000 
M5682 diff_95000_5192000# diff_5626000_2182000# diff_5626000_2182000# GND efet w=13000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5683 diff_5626000_2182000# diff_5619000_2172000# diff_83000_3098000# GND efet w=154500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5684 diff_5619000_2172000# diff_5769000_2161000# diff_95000_5192000# GND efet w=775000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5685 diff_5626000_2091000# diff_5619000_2102000# diff_83000_3098000# GND efet w=155000 l=9000
+ ad=-1.96197e+09 pd=400000 as=0 ps=0 
M5686 diff_5769000_2028000# diff_5087000_472000# diff_83000_3098000# GND efet w=485000 l=9000
+ ad=1.45407e+09 pd=1.61e+06 as=0 ps=0 
M5687 diff_5626000_2091000# diff_72000_4515000# diff_5618000_1925000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=1.023e+09 ps=234000 
M5688 diff_95000_5192000# diff_5626000_2091000# diff_5626000_2091000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5689 diff_95000_5192000# diff_5769000_2028000# diff_5619000_2102000# GND efet w=778000 l=8000
+ ad=0 pd=0 as=-2.05864e+09 ps=6.806e+06 
M5690 diff_95000_5192000# diff_5651000_2014000# diff_5618000_1925000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5691 diff_5651000_2014000# diff_5632000_1934000# diff_83000_3098000# GND efet w=47000 l=8000
+ ad=1.164e+09 pd=214000 as=0 ps=0 
M5692 diff_95000_5192000# diff_5769000_2028000# diff_5619000_2102000# GND efet w=286000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5693 diff_5769000_2028000# diff_5697000_1749000# diff_83000_3098000# GND efet w=478000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5694 diff_95000_5192000# diff_5651000_2014000# diff_5651000_2014000# GND efet w=12000 l=35000
+ ad=0 pd=0 as=0 ps=0 
M5695 diff_95000_5192000# diff_5769000_2028000# diff_5619000_2102000# GND efet w=285500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5696 diff_5651000_2014000# diff_72000_4515000# diff_83000_3098000# GND efet w=28000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5697 diff_5632000_1934000# diff_5618000_1925000# diff_83000_3098000# GND efet w=222500 l=8500
+ ad=-5.04967e+08 pd=730000 as=0 ps=0 
M5698 diff_5243000_1641000# diff_5243000_1641000# diff_95000_5192000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M5699 diff_5333000_1645000# diff_72000_4515000# diff_5243000_1641000# GND efet w=19000 l=11000
+ ad=1.71e+08 pd=56000 as=0 ps=0 
M5700 diff_5354000_1645000# diff_4328000_910000# diff_5333000_1645000# GND efet w=19000 l=12000
+ ad=3.38e+08 pd=90000 as=0 ps=0 
M5701 diff_5375000_1681000# diff_5375000_1681000# diff_95000_5192000# GND efet w=13000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M5702 diff_817000_1663000# diff_5271000_2493000# diff_5375000_1681000# GND efet w=87500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5703 diff_95000_5192000# diff_4990000_1457000# diff_4990000_1457000# GND efet w=13000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M5704 diff_95000_5192000# diff_5069000_1595000# diff_5069000_1595000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=1.669e+09 ps=364000 
M5705 diff_5123000_1614000# diff_4932000_827000# diff_95000_5192000# GND efet w=13000 l=8000
+ ad=-8.9673e+06 pd=892000 as=0 ps=0 
M5706 diff_5159000_1628000# diff_4990000_1457000# diff_5123000_1614000# GND efet w=129500 l=9500
+ ad=-7.99967e+08 pd=692000 as=0 ps=0 
M5707 diff_83000_3098000# diff_4727000_1383000# diff_4870000_1328000# GND efet w=59000 l=8000
+ ad=0 pd=0 as=-1.30597e+09 ps=476000 
M5708 diff_83000_3098000# diff_4839000_2618000# diff_4693000_1304000# GND efet w=50000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5709 diff_4990000_1457000# diff_4727000_1483000# diff_4970000_1482000# GND efet w=33000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M5710 diff_83000_3098000# diff_4994000_2634000# diff_4990000_1457000# GND efet w=55000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5711 diff_4990000_1457000# diff_4871000_1557000# diff_83000_3098000# GND efet w=44000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M5712 diff_5123000_1614000# diff_5069000_1595000# diff_83000_3098000# GND efet w=90000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5713 diff_5069000_1595000# diff_4694000_1563000# diff_83000_3098000# GND efet w=65500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5714 diff_83000_3098000# diff_4932000_827000# diff_5069000_1595000# GND efet w=65000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5715 diff_5243000_1607000# diff_5243000_1607000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=2.139e+09 pd=498000 as=0 ps=0 
M5716 diff_95000_5192000# diff_5202000_1588000# diff_5202000_1588000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=1.631e+09 ps=352000 
M5717 diff_5288000_1548000# diff_4990000_1457000# diff_5243000_1607000# GND efet w=77500 l=8500
+ ad=1.376e+09 pd=336000 as=0 ps=0 
M5718 diff_4693000_1304000# diff_4705000_1351000# diff_4808000_1269000# GND efet w=69000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5719 diff_4870000_1328000# diff_4839000_2618000# diff_83000_3098000# GND efet w=58000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M5720 diff_95000_5192000# diff_4694000_1185000# diff_4694000_1185000# GND efet w=13000 l=25000
+ ad=0 pd=0 as=-1.17697e+09 ps=544000 
M5721 diff_95000_5192000# diff_4727000_1106000# diff_4727000_1106000# GND efet w=13000 l=24000
+ ad=0 pd=0 as=1.519e+09 ps=298000 
M5722 diff_4424000_962000# diff_4374000_833000# diff_83000_3098000# GND efet w=20000 l=9000
+ ad=1.794e+09 pd=386000 as=0 ps=0 
M5723 diff_4424000_962000# diff_4417000_952000# diff_4363000_2478000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5724 diff_3577000_991000# diff_95000_5192000# diff_95000_5192000# GND efet w=13000 l=104000
+ ad=0 pd=0 as=0 ps=0 
M5725 diff_4518000_901000# diff_3577000_991000# diff_83000_3098000# GND efet w=49000 l=8000
+ ad=1.962e+09 pd=392000 as=0 ps=0 
M5726 diff_83000_3098000# diff_4608000_1093000# diff_4459000_1183000# GND efet w=48000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5727 diff_4608000_1093000# diff_817000_1211000# diff_83000_3098000# GND efet w=66000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5728 diff_4432000_1144000# diff_4548000_2725000# diff_4608000_1093000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5729 diff_4705000_1142000# diff_4602000_2752000# diff_4432000_1144000# GND efet w=21000 l=12000
+ ad=3.99e+08 pd=80000 as=0 ps=0 
M5730 diff_4459000_1108000# diff_4498000_2492000# diff_4424000_962000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5731 diff_83000_3098000# diff_4608000_946000# diff_4459000_1108000# GND efet w=49000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5732 diff_4608000_946000# diff_817000_909000# diff_83000_3098000# GND efet w=67000 l=8000
+ ad=1.778e+09 pd=402000 as=0 ps=0 
M5733 diff_4705000_1097000# diff_4602000_2752000# diff_4518000_1196000# GND efet w=21000 l=12000
+ ad=4.68e+08 pd=138000 as=0 ps=0 
M5734 diff_83000_3098000# diff_4705000_1097000# diff_4727000_1106000# GND efet w=49000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5735 diff_4785000_1099000# diff_4740000_2641000# diff_83000_3098000# GND efet w=148500 l=8500
+ ad=1.748e+09 pd=370000 as=0 ps=0 
M5736 diff_4808000_1138000# diff_4727000_1106000# diff_4785000_1099000# GND efet w=126000 l=9000
+ ad=-2.05097e+09 pd=418000 as=0 ps=0 
M5737 diff_4694000_1185000# diff_4705000_1142000# diff_4808000_1138000# GND efet w=69000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5738 diff_83000_3098000# diff_4705000_1351000# diff_4870000_1328000# GND efet w=54000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5739 diff_4870000_1328000# diff_4870000_1328000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5740 diff_4951000_1273000# diff_4705000_1351000# diff_83000_3098000# GND efet w=135000 l=9000
+ ad=1.35e+09 pd=290000 as=0 ps=0 
M5741 diff_4970000_1273000# diff_4768000_996000# diff_4951000_1273000# GND efet w=135000 l=9000
+ ad=1.827e+09 pd=354000 as=0 ps=0 
M5742 diff_4990000_1273000# diff_4727000_1383000# diff_4970000_1273000# GND efet w=31000 l=7000
+ ad=-4.38967e+08 pd=692000 as=0 ps=0 
M5743 diff_5333000_1602000# diff_72000_4515000# diff_5243000_1607000# GND efet w=20000 l=11000
+ ad=1.8e+08 pd=58000 as=0 ps=0 
M5744 diff_5354000_1602000# diff_4328000_910000# diff_5333000_1602000# GND efet w=20000 l=12000
+ ad=3.19e+08 pd=102000 as=0 ps=0 
M5745 diff_5202000_1588000# diff_5159000_1628000# diff_83000_3098000# GND efet w=77000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5746 diff_5123000_1614000# diff_5069000_1595000# diff_83000_3098000# GND efet w=47500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5747 diff_5123000_1263000# diff_5069000_1278000# diff_83000_3098000# GND efet w=122000 l=9000
+ ad=1.00033e+08 pd=854000 as=0 ps=0 
M5748 diff_4990000_1273000# diff_4727000_1383000# diff_4970000_1273000# GND efet w=97000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M5749 diff_83000_3098000# diff_4994000_2634000# diff_4990000_1273000# GND efet w=54000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5750 diff_4990000_1273000# diff_4870000_1328000# diff_83000_3098000# GND efet w=45000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M5751 diff_5069000_1278000# diff_4693000_1304000# diff_83000_3098000# GND efet w=63500 l=8500
+ ad=1.762e+09 pd=358000 as=0 ps=0 
M5752 diff_83000_3098000# diff_4932000_827000# diff_5069000_1278000# GND efet w=64000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5753 diff_95000_5192000# diff_4871000_1180000# diff_4871000_1180000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=-1.49297e+09 ps=464000 
M5754 diff_83000_3098000# diff_4705000_1142000# diff_4871000_1180000# GND efet w=51000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5755 diff_4871000_1180000# diff_4839000_2618000# diff_83000_3098000# GND efet w=63000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5756 diff_4694000_1185000# diff_4705000_1142000# diff_4808000_1138000# GND efet w=68500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5757 diff_4808000_1138000# diff_4727000_1106000# diff_4785000_1099000# GND efet w=11000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5758 diff_83000_3098000# diff_4839000_2618000# diff_4694000_1185000# GND efet w=51000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5759 diff_4705000_1019000# diff_4602000_2752000# diff_4518000_901000# GND efet w=20000 l=12000
+ ad=4.63e+08 pd=118000 as=0 ps=0 
M5760 diff_4518000_901000# diff_4518000_901000# diff_95000_5192000# GND efet w=13000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M5761 diff_83000_3098000# diff_72000_4515000# diff_4374000_833000# GND efet w=82000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5762 diff_4417000_952000# diff_72000_4515000# diff_83000_3098000# GND efet w=70000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5763 diff_4424000_962000# diff_4548000_2725000# diff_4608000_946000# GND efet w=20000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5764 diff_4705000_974000# diff_4602000_2752000# diff_4424000_962000# GND efet w=20000 l=12000
+ ad=4e+08 pd=80000 as=0 ps=0 
M5765 diff_83000_3098000# diff_4705000_1019000# diff_4727000_1006000# GND efet w=50000 l=8000
+ ad=0 pd=0 as=1.497e+09 ps=298000 
M5766 diff_4786000_981000# diff_4768000_996000# diff_83000_3098000# GND efet w=26000 l=9000
+ ad=1.883e+09 pd=400000 as=0 ps=0 
M5767 diff_4808000_919000# diff_4727000_1006000# diff_4786000_981000# GND efet w=10000 l=9000
+ ad=-2.10897e+09 pd=436000 as=0 ps=0 
M5768 diff_4808000_919000# diff_4727000_1006000# diff_4786000_981000# GND efet w=137000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5769 diff_4693000_927000# diff_4705000_974000# diff_4808000_919000# GND efet w=67500 l=8500
+ ad=-1.35097e+09 pd=550000 as=0 ps=0 
M5770 diff_4786000_981000# diff_4768000_996000# diff_83000_3098000# GND efet w=108000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5771 diff_4459000_1108000# diff_4459000_1108000# diff_95000_5192000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M5772 diff_4608000_946000# diff_4608000_946000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M5773 diff_83000_3098000# diff_72000_4515000# diff_4498000_2492000# GND efet w=75000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5774 diff_4548000_2725000# diff_72000_4515000# diff_83000_3098000# GND efet w=75000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5775 diff_4602000_2752000# diff_72000_4515000# diff_83000_3098000# GND efet w=74500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5776 diff_4693000_927000# diff_4693000_927000# diff_95000_5192000# GND efet w=12000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M5777 diff_4727000_1006000# diff_4727000_1006000# diff_95000_5192000# GND efet w=14000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M5778 diff_83000_3098000# diff_4727000_1106000# diff_4871000_1180000# GND efet w=58000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5779 diff_4950000_1104000# diff_4705000_1142000# diff_83000_3098000# GND efet w=135000 l=8000
+ ad=1.485e+09 pd=292000 as=0 ps=0 
M5780 diff_4970000_1104000# diff_4768000_996000# diff_4950000_1104000# GND efet w=135000 l=9000
+ ad=1.831e+09 pd=354000 as=0 ps=0 
M5781 diff_4990000_1079000# diff_4727000_1106000# diff_4970000_1104000# GND efet w=96000 l=7000
+ ad=-1.88967e+08 pd=696000 as=0 ps=0 
M5782 diff_4990000_1273000# diff_4990000_1273000# diff_95000_5192000# GND efet w=13000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M5783 diff_5069000_1278000# diff_5069000_1278000# diff_95000_5192000# GND efet w=12000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M5784 diff_5123000_1614000# diff_4990000_1273000# diff_5123000_1263000# GND efet w=41000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5785 diff_83000_3098000# diff_4990000_1457000# diff_5202000_1588000# GND efet w=70500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5786 diff_5243000_1607000# diff_5202000_1588000# diff_83000_3098000# GND efet w=63500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5787 diff_5288000_1548000# diff_4990000_1457000# diff_5243000_1607000# GND efet w=32000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5788 diff_83000_3098000# diff_5159000_1628000# diff_5288000_1548000# GND efet w=115500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5789 diff_5201000_1284000# diff_5123000_1614000# diff_83000_3098000# GND efet w=77000 l=8000
+ ad=1.57e+09 pd=344000 as=0 ps=0 
M5790 diff_83000_3098000# diff_4990000_1273000# diff_5201000_1284000# GND efet w=70500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5791 diff_83000_3098000# diff_5123000_1614000# diff_5288000_1289000# GND efet w=119500 l=8500
+ ad=0 pd=0 as=1.4e+09 ps=338000 
M5792 diff_5243000_1264000# diff_5201000_1284000# diff_83000_3098000# GND efet w=64500 l=8500
+ ad=-2.04297e+09 pd=502000 as=0 ps=0 
M5793 diff_5123000_1263000# diff_5069000_1278000# diff_83000_3098000# GND efet w=22000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5794 diff_5123000_1614000# diff_4990000_1273000# diff_5123000_1263000# GND efet w=71000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5795 diff_5288000_1289000# diff_4990000_1273000# diff_5243000_1264000# GND efet w=34000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5796 diff_5201000_1284000# diff_5201000_1284000# diff_95000_5192000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5797 diff_5123000_1263000# diff_4932000_827000# diff_95000_5192000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5798 diff_5288000_1289000# diff_4990000_1273000# diff_5243000_1264000# GND efet w=74000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5799 diff_95000_5192000# diff_5375000_1574000# diff_5375000_1574000# GND efet w=13000 l=22000
+ ad=0 pd=0 as=-1.55597e+09 ps=536000 
M5800 diff_5375000_1574000# diff_5354000_1602000# diff_83000_3098000# GND efet w=190000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5801 diff_5331000_4062000# diff_5375000_1574000# diff_83000_3098000# GND efet w=155500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5802 diff_817000_1588000# diff_5271000_2493000# diff_5375000_1574000# GND efet w=87500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5803 diff_95000_5192000# diff_5632000_1934000# diff_5632000_1934000# GND efet w=12000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M5804 diff_83000_3098000# diff_83000_3098000# diff_5619000_2102000# GND efet w=92500 l=12500
+ ad=0 pd=0 as=0 ps=0 
M5805 diff_5619000_2102000# diff_5769000_2028000# diff_95000_5192000# GND efet w=287000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5806 diff_5769000_2028000# diff_5769000_2028000# diff_95000_5192000# GND efet w=44000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5807 diff_83000_3098000# diff_5697000_1749000# diff_5619000_2102000# GND efet w=239000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5808 diff_95000_5192000# diff_5697000_1749000# diff_5697000_1749000# GND efet w=33000 l=8000
+ ad=0 pd=0 as=2.09107e+09 ps=1.774e+06 
M5809 diff_5697000_1749000# diff_5087000_472000# diff_83000_3098000# GND efet w=475000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5810 diff_5632000_1934000# diff_5011000_576000# diff_817000_1965000# GND efet w=87000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5811 diff_83000_3098000# diff_5650000_1749000# diff_5697000_1749000# GND efet w=513000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5812 diff_817000_1965000# diff_4954000_639000# diff_5650000_1749000# GND efet w=35000 l=12000
+ ad=0 pd=0 as=-1.50297e+09 ps=322000 
M5813 diff_83000_3098000# diff_5697000_1749000# diff_5619000_2102000# GND efet w=289000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5814 diff_83000_3098000# diff_5697000_1749000# diff_5619000_2102000# GND efet w=290000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5815 diff_5619000_2102000# diff_5697000_1749000# diff_83000_3098000# GND efet w=801500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5816 diff_5696000_1731000# diff_5650000_1678000# diff_83000_3098000# GND efet w=514000 l=9000
+ ad=1.81607e+09 pd=1.792e+06 as=0 ps=0 
M5817 diff_83000_3098000# diff_5696000_1731000# diff_5619000_1381000# GND efet w=803000 l=10000
+ ad=0 pd=0 as=1.29633e+09 ps=6.762e+06 
M5818 diff_83000_3098000# diff_5087000_472000# diff_5696000_1731000# GND efet w=475500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5819 diff_5650000_1678000# diff_4954000_639000# diff_817000_1663000# GND efet w=35000 l=11000
+ ad=-1.53797e+09 pd=300000 as=0 ps=0 
M5820 diff_817000_1663000# diff_5011000_576000# diff_5632000_1485000# GND efet w=87000 l=11000
+ ad=0 pd=0 as=-2.60967e+08 ps=734000 
M5821 diff_95000_5192000# diff_95000_5192000# diff_5159000_1628000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M5822 diff_5159000_1628000# diff_5473000_1600000# diff_83000_3098000# GND efet w=126000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5823 diff_5375000_1305000# diff_5354000_1269000# diff_83000_3098000# GND efet w=198000 l=8000
+ ad=-1.50697e+09 pd=518000 as=0 ps=0 
M5824 diff_5331000_4062000# diff_5375000_1305000# diff_83000_3098000# GND efet w=153500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5825 diff_5243000_1264000# diff_5243000_1264000# diff_95000_5192000# GND efet w=11000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M5826 diff_5334000_1269000# diff_72000_4515000# diff_5243000_1264000# GND efet w=19000 l=12000
+ ad=1.52e+08 pd=54000 as=0 ps=0 
M5827 diff_5354000_1269000# diff_4328000_910000# diff_5334000_1269000# GND efet w=19000 l=12000
+ ad=3.34e+08 pd=92000 as=0 ps=0 
M5828 diff_5375000_1305000# diff_5375000_1305000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M5829 diff_817000_1286000# diff_5271000_2493000# diff_5375000_1305000# GND efet w=87500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5830 diff_95000_5192000# diff_4990000_1079000# diff_4990000_1079000# GND efet w=13000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M5831 diff_95000_5192000# diff_5069000_1218000# diff_5069000_1218000# GND efet w=13000 l=20000
+ ad=0 pd=0 as=1.684e+09 ps=366000 
M5832 diff_5123000_1237000# diff_4932000_827000# diff_95000_5192000# GND efet w=13000 l=8000
+ ad=2.69033e+08 pd=962000 as=0 ps=0 
M5833 diff_5123000_1263000# diff_4990000_1079000# diff_5123000_1237000# GND efet w=129500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5834 diff_83000_3098000# diff_4727000_1006000# diff_4870000_939000# GND efet w=60000 l=8000
+ ad=0 pd=0 as=-9.88967e+08 ps=606000 
M5835 diff_4990000_1079000# diff_4727000_1106000# diff_4970000_1104000# GND efet w=33000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M5836 diff_83000_3098000# diff_4994000_2634000# diff_4990000_1079000# GND efet w=55000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5837 diff_4990000_1079000# diff_4871000_1180000# diff_83000_3098000# GND efet w=45000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M5838 diff_5123000_1237000# diff_5069000_1218000# diff_83000_3098000# GND efet w=90000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5839 diff_5069000_1218000# diff_4694000_1185000# diff_83000_3098000# GND efet w=65500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5840 diff_83000_3098000# diff_4932000_827000# diff_5069000_1218000# GND efet w=66000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5841 diff_5243000_1229000# diff_5243000_1229000# diff_95000_5192000# GND efet w=13000 l=21000
+ ad=-2.09097e+09 pd=502000 as=0 ps=0 
M5842 diff_5288000_1171000# diff_4990000_1079000# diff_5243000_1229000# GND efet w=77500 l=8500
+ ad=1.38e+09 pd=336000 as=0 ps=0 
M5843 diff_95000_5192000# diff_5202000_1210000# diff_5202000_1210000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=1.609e+09 ps=350000 
M5844 diff_83000_3098000# diff_4839000_2618000# diff_4870000_939000# GND efet w=58000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5845 diff_4693000_927000# diff_4705000_974000# diff_4808000_919000# GND efet w=76000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5846 diff_4870000_939000# diff_4870000_939000# diff_95000_5192000# GND efet w=12000 l=22000
+ ad=0 pd=0 as=0 ps=0 
M5847 diff_83000_3098000# diff_4705000_974000# diff_4870000_939000# GND efet w=52500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5848 diff_4707000_840000# diff_4707000_840000# diff_95000_5192000# GND efet w=13000 l=36000
+ ad=1.332e+09 pd=254000 as=0 ps=0 
M5849 diff_4948000_897000# diff_4705000_974000# diff_83000_3098000# GND efet w=133000 l=9000
+ ad=1.832e+09 pd=352000 as=0 ps=0 
M5850 diff_4969000_890000# diff_4768000_996000# diff_4948000_897000# GND efet w=64000 l=9000
+ ad=1.895e+09 pd=416000 as=0 ps=0 
M5851 diff_4990000_890000# diff_4727000_1006000# diff_4969000_890000# GND efet w=32000 l=7000
+ ad=-2.75967e+08 pd=710000 as=0 ps=0 
M5852 diff_5334000_1225000# diff_72000_4515000# diff_5243000_1229000# GND efet w=21000 l=12000
+ ad=1.68e+08 pd=58000 as=0 ps=0 
M5853 diff_5354000_1225000# diff_4328000_910000# diff_5334000_1225000# GND efet w=21000 l=12000
+ ad=3.36e+08 pd=102000 as=0 ps=0 
M5854 diff_5202000_1210000# diff_5123000_1263000# diff_83000_3098000# GND efet w=77000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5855 diff_5123000_1237000# diff_5069000_1218000# diff_83000_3098000# GND efet w=47000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5856 diff_5123000_886000# diff_5069000_901000# diff_83000_3098000# GND efet w=122000 l=9000
+ ad=-1.60897e+09 pd=550000 as=0 ps=0 
M5857 diff_95000_5192000# diff_4838000_814000# diff_4838000_814000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=1.06e+09 ps=206000 
M5858 diff_4969000_890000# diff_4768000_996000# diff_4948000_897000# GND efet w=65000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5859 diff_4990000_890000# diff_4727000_1006000# diff_4969000_890000# GND efet w=113500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5860 diff_83000_3098000# diff_4994000_2634000# diff_4990000_890000# GND efet w=50000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5861 diff_4990000_890000# diff_4870000_939000# diff_83000_3098000# GND efet w=45000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M5862 diff_5069000_901000# diff_4693000_927000# diff_83000_3098000# GND efet w=64500 l=8500
+ ad=1.795e+09 pd=360000 as=0 ps=0 
M5863 diff_83000_3098000# diff_4932000_827000# diff_5069000_901000# GND efet w=65000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5864 diff_4990000_890000# diff_4990000_890000# diff_95000_5192000# GND efet w=12000 l=25000
+ ad=0 pd=0 as=0 ps=0 
M5865 diff_5069000_901000# diff_5069000_901000# diff_95000_5192000# GND efet w=12000 l=19000
+ ad=0 pd=0 as=0 ps=0 
M5866 diff_5123000_1237000# diff_4990000_890000# diff_5123000_886000# GND efet w=41000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5867 diff_83000_3098000# diff_4990000_1079000# diff_5202000_1210000# GND efet w=71500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5868 diff_5243000_1229000# diff_5202000_1210000# diff_83000_3098000# GND efet w=63500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5869 diff_5288000_1171000# diff_4990000_1079000# diff_5243000_1229000# GND efet w=33000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5870 diff_83000_3098000# diff_5123000_1263000# diff_5288000_1171000# GND efet w=115500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5871 diff_5201000_907000# diff_5123000_1237000# diff_83000_3098000# GND efet w=77000 l=8000
+ ad=1.577e+09 pd=344000 as=0 ps=0 
M5872 diff_83000_3098000# diff_4990000_890000# diff_5201000_907000# GND efet w=70500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5873 diff_83000_3098000# diff_5123000_1237000# diff_5288000_912000# GND efet w=118500 l=8500
+ ad=0 pd=0 as=1.388e+09 ps=338000 
M5874 diff_5243000_887000# diff_5201000_907000# diff_83000_3098000# GND efet w=64500 l=8500
+ ad=-2.04097e+09 pd=502000 as=0 ps=0 
M5875 diff_5123000_886000# diff_5069000_901000# diff_83000_3098000# GND efet w=21000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5876 diff_5123000_1237000# diff_4990000_890000# diff_5123000_886000# GND efet w=71000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5877 diff_5288000_912000# diff_4990000_890000# diff_5243000_887000# GND efet w=34000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5878 diff_5123000_886000# diff_4932000_827000# diff_95000_5192000# GND efet w=13000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5879 diff_5201000_907000# diff_5201000_907000# diff_95000_5192000# GND efet w=13000 l=23000
+ ad=0 pd=0 as=0 ps=0 
M5880 diff_5288000_912000# diff_4990000_890000# diff_5243000_887000# GND efet w=74000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5881 diff_95000_5192000# diff_5375000_1196000# diff_5375000_1196000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=-1.51397e+09 ps=538000 
M5882 diff_5375000_1196000# diff_5354000_1225000# diff_83000_3098000# GND efet w=193000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5883 diff_5331000_4062000# diff_5375000_1196000# diff_83000_3098000# GND efet w=155500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5884 diff_817000_1211000# diff_5271000_2493000# diff_5375000_1196000# GND efet w=87500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5885 diff_5371000_3654000# diff_5354000_892000# diff_83000_3098000# GND efet w=197000 l=8000
+ ad=1.32707e+09 pd=1.962e+06 as=0 ps=0 
M5886 diff_5331000_4062000# diff_5371000_3654000# diff_83000_3098000# GND efet w=154500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5887 diff_5243000_887000# diff_5243000_887000# diff_95000_5192000# GND efet w=11000 l=20000
+ ad=0 pd=0 as=0 ps=0 
M5888 diff_5333000_892000# diff_72000_4515000# diff_5243000_887000# GND efet w=19000 l=11000
+ ad=1.9e+08 pd=58000 as=0 ps=0 
M5889 diff_5354000_892000# diff_4328000_910000# diff_5333000_892000# GND efet w=19000 l=11000
+ ad=3.28e+08 pd=90000 as=0 ps=0 
M5890 diff_5371000_3654000# diff_5371000_3654000# diff_95000_5192000# GND efet w=13000 l=14000
+ ad=0 pd=0 as=0 ps=0 
M5891 diff_817000_909000# diff_5271000_2493000# diff_5371000_3654000# GND efet w=88500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5892 diff_5632000_1485000# diff_5618000_1427000# diff_83000_3098000# GND efet w=220500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5893 diff_83000_3098000# diff_5696000_1731000# diff_5619000_1381000# GND efet w=289500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M5894 diff_83000_3098000# diff_5696000_1731000# diff_5619000_1381000# GND efet w=288500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5895 diff_5696000_1731000# diff_5696000_1731000# diff_5696000_1731000# GND efet w=2000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M5896 diff_5619000_1381000# diff_5696000_1731000# diff_83000_3098000# GND efet w=238500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M5897 diff_5696000_1731000# diff_5696000_1731000# diff_95000_5192000# GND efet w=36000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M5898 diff_95000_5192000# diff_5632000_1485000# diff_5632000_1485000# GND efet w=11000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M5899 diff_83000_3098000# diff_72000_4515000# diff_5651000_1464000# GND efet w=28000 l=9000
+ ad=0 pd=0 as=1.145e+09 ps=214000 
M5900 diff_95000_5192000# diff_5769000_1368000# diff_5769000_1368000# GND efet w=44000 l=8000
+ ad=0 pd=0 as=1.18607e+09 ps=1.612e+06 
M5901 diff_83000_3098000# diff_5696000_1731000# diff_5769000_1368000# GND efet w=478000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5902 diff_5619000_1381000# diff_5769000_1368000# diff_95000_5192000# GND efet w=285000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5903 diff_95000_5192000# diff_5769000_1368000# diff_5619000_1381000# GND efet w=285500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5904 diff_95000_5192000# diff_5651000_1464000# diff_5651000_1464000# GND efet w=11000 l=35000
+ ad=0 pd=0 as=0 ps=0 
M5905 diff_5651000_1464000# diff_5632000_1485000# diff_83000_3098000# GND efet w=43500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5906 diff_95000_5192000# diff_5651000_1464000# diff_5618000_1427000# GND efet w=14000 l=12000
+ ad=0 pd=0 as=1.025e+09 ps=232000 
M5907 diff_83000_3098000# diff_5087000_472000# diff_5769000_1368000# GND efet w=485500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5908 diff_95000_5192000# diff_5769000_1368000# diff_5619000_1381000# GND efet w=286000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5909 diff_5618000_1427000# diff_72000_4515000# diff_5626000_1390000# GND efet w=19000 l=10000
+ ad=0 pd=0 as=1.991e+09 ps=396000 
M5910 diff_95000_5192000# diff_5626000_1390000# diff_5626000_1390000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M5911 diff_5619000_1381000# diff_5769000_1368000# diff_95000_5192000# GND efet w=786000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5912 diff_5626000_1390000# diff_5619000_1381000# diff_83000_3098000# GND efet w=155000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5913 diff_83000_3098000# diff_83000_3098000# diff_5619000_1381000# GND efet w=97000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M5914 diff_5626000_1299000# diff_5619000_1309000# diff_83000_3098000# GND efet w=155500 l=9500
+ ad=-1.96397e+09 pd=400000 as=0 ps=0 
M5915 diff_5769000_1236000# diff_5087000_472000# diff_83000_3098000# GND efet w=485000 l=9000
+ ad=1.28307e+09 pd=1.608e+06 as=0 ps=0 
M5916 diff_83000_3098000# diff_4727000_1006000# diff_4707000_840000# GND efet w=42000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M5917 diff_4776000_738000# diff_4705000_974000# diff_83000_3098000# GND efet w=42000 l=8000
+ ad=1.176e+09 pd=258000 as=0 ps=0 
M5918 diff_83000_3098000# diff_4870000_939000# diff_4838000_814000# GND efet w=43000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5919 diff_83000_3098000# diff_72000_4515000# diff_4932000_827000# GND efet w=71000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M5920 diff_83000_3098000# diff_4707000_840000# diff_5009000_805000# GND efet w=137500 l=7500
+ ad=0 pd=0 as=-7.66967e+08 ps=628000 
M5921 diff_4776000_738000# diff_4776000_738000# diff_95000_5192000# GND efet w=12000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M5922 diff_3396000_614000# diff_3396000_614000# diff_95000_5192000# GND efet w=16000 l=8000
+ ad=-5.07967e+08 pd=636000 as=0 ps=0 
M5923 diff_83000_3098000# diff_1851000_1456000# diff_3396000_614000# GND efet w=231000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5924 diff_3332000_585000# diff_3332000_585000# diff_95000_5192000# GND efet w=50500 l=7500
+ ad=-7.99019e+07 pd=1.982e+06 as=0 ps=0 
M5925 diff_83000_3098000# diff_3482000_568000# diff_3332000_585000# GND efet w=483500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5926 diff_3482000_568000# diff_680000_1019000# diff_3396000_614000# GND efet w=35000 l=11000
+ ad=7.5e+08 pd=182000 as=0 ps=0 
M5927 diff_95000_5192000# diff_3258000_123000# diff_3258000_123000# GND efet w=34000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5928 diff_83000_3098000# diff_553000_1211000# diff_3332000_585000# GND efet w=437000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5929 diff_3258000_123000# diff_3332000_585000# diff_83000_3098000# GND efet w=44000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5930 diff_83000_3098000# diff_3746000_568000# diff_3673000_545000# GND efet w=489500 l=8500
+ ad=0 pd=0 as=-1.76902e+08 ps=1.99e+06 
M5931 diff_83000_3098000# diff_553000_1211000# diff_3673000_545000# GND efet w=437000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5932 diff_95000_5192000# diff_3673000_545000# diff_3673000_545000# GND efet w=52500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M5933 diff_83000_3098000# diff_1851000_1376000# diff_3852000_625000# GND efet w=231500 l=8500
+ ad=0 pd=0 as=-3.52967e+08 ps=640000 
M5934 diff_95000_5192000# diff_3852000_625000# diff_3852000_625000# GND efet w=16000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5935 diff_3852000_625000# diff_680000_1019000# diff_3746000_568000# GND efet w=35000 l=11000
+ ad=0 pd=0 as=6.62e+08 ps=176000 
M5936 diff_83000_3098000# diff_3673000_545000# diff_3899000_565000# GND efet w=273000 l=8000
+ ad=0 pd=0 as=2.07007e+09 ps=1.494e+06 
M5937 diff_83000_3098000# diff_553000_1211000# diff_3899000_565000# GND efet w=301500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5938 diff_3899000_565000# diff_3673000_545000# diff_83000_3098000# GND efet w=45000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5939 diff_3265000_456000# diff_3258000_123000# diff_83000_3098000# GND efet w=183000 l=8000
+ ad=1.00294e+08 pd=4.558e+06 as=0 ps=0 
M5940 diff_83000_3098000# diff_3258000_123000# diff_3265000_456000# GND efet w=184000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5941 diff_2458000_131000# diff_2524000_585000# diff_95000_5192000# GND efet w=269000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5942 diff_3265000_456000# diff_3258000_123000# diff_83000_3098000# GND efet w=646500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5943 diff_83000_3098000# diff_3258000_123000# diff_3265000_456000# GND efet w=191000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5944 diff_95000_5192000# diff_3332000_585000# diff_3265000_456000# GND efet w=208000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5945 diff_95000_5192000# diff_3332000_585000# diff_3265000_456000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5946 diff_95000_5192000# diff_3332000_585000# diff_3265000_456000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5947 diff_95000_5192000# diff_3332000_585000# diff_3265000_456000# GND efet w=190000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5948 diff_3687000_194000# diff_3673000_545000# diff_95000_5192000# GND efet w=191000 l=8000
+ ad=5.62943e+07 pd=4.556e+06 as=0 ps=0 
M5949 diff_95000_5192000# diff_3332000_585000# diff_3265000_456000# GND efet w=651000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5950 diff_3265000_456000# diff_3258000_123000# diff_83000_3098000# GND efet w=280000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5951 diff_95000_5192000# diff_3673000_545000# diff_3687000_194000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5952 diff_3687000_194000# diff_3673000_545000# diff_95000_5192000# GND efet w=651000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5953 diff_95000_5192000# diff_3673000_545000# diff_3687000_194000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5954 diff_95000_5192000# diff_3673000_545000# diff_3687000_194000# GND efet w=208000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5955 diff_3899000_565000# diff_3899000_565000# diff_95000_5192000# GND efet w=34000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5956 diff_3899000_565000# diff_553000_1211000# diff_83000_3098000# GND efet w=56000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5957 diff_83000_3098000# diff_3899000_565000# diff_3687000_194000# GND efet w=191000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5958 diff_83000_3098000# diff_553000_1211000# diff_4088000_123000# GND efet w=56000 l=8000
+ ad=0 pd=0 as=2.01407e+09 ps=1.486e+06 
M5959 diff_83000_3098000# diff_553000_1211000# diff_4088000_123000# GND efet w=300000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5960 diff_83000_3098000# diff_4162000_585000# diff_4088000_123000# GND efet w=272000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5961 diff_4227000_613000# diff_4227000_613000# diff_95000_5192000# GND efet w=16000 l=8000
+ ad=-5.87967e+08 pd=636000 as=0 ps=0 
M5962 diff_83000_3098000# diff_1851000_1079000# diff_4227000_613000# GND efet w=232000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5963 diff_4162000_585000# diff_4162000_585000# diff_95000_5192000# GND efet w=51000 l=8000
+ ad=-2.35902e+08 pd=1.986e+06 as=0 ps=0 
M5964 diff_83000_3098000# diff_4312000_568000# diff_4162000_585000# GND efet w=483500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5965 diff_4312000_568000# diff_680000_1019000# diff_4227000_613000# GND efet w=35000 l=12000
+ ad=6.92e+08 pd=178000 as=0 ps=0 
M5966 diff_95000_5192000# diff_4088000_123000# diff_4088000_123000# GND efet w=34000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5967 diff_83000_3098000# diff_553000_1211000# diff_4162000_585000# GND efet w=439000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5968 diff_4088000_123000# diff_4162000_585000# diff_83000_3098000# GND efet w=44000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5969 diff_83000_3098000# diff_3899000_565000# diff_3687000_194000# GND efet w=184500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5970 diff_83000_3098000# diff_3899000_565000# diff_3687000_194000# GND efet w=181000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5971 diff_4096000_194000# diff_4088000_123000# diff_83000_3098000# GND efet w=182000 l=8000
+ ad=3.25294e+08 pd=4.544e+06 as=0 ps=0 
M5972 diff_83000_3098000# diff_3899000_565000# diff_3687000_194000# GND efet w=644500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5973 diff_83000_3098000# diff_4088000_123000# diff_4096000_194000# GND efet w=181500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5974 diff_83000_3098000# diff_4576000_568000# diff_4503000_546000# GND efet w=487500 l=8500
+ ad=0 pd=0 as=-2.53902e+08 ps=1.99e+06 
M5975 diff_83000_3098000# diff_553000_1211000# diff_4503000_546000# GND efet w=439000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5976 diff_95000_5192000# diff_4503000_546000# diff_4503000_546000# GND efet w=52000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5977 diff_83000_3098000# diff_1851000_999000# diff_4683000_625000# GND efet w=230000 l=8000
+ ad=0 pd=0 as=-3.47967e+08 ps=638000 
M5978 diff_95000_5192000# diff_4683000_625000# diff_4683000_625000# GND efet w=16000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5979 diff_83000_3098000# diff_4503000_546000# diff_4729000_565000# GND efet w=273000 l=9000
+ ad=0 pd=0 as=-2.1379e+09 ps=1.494e+06 
M5980 diff_4683000_625000# diff_680000_1019000# diff_4576000_568000# GND efet w=35000 l=12000
+ ad=0 pd=0 as=6.84e+08 ps=176000 
M5981 diff_83000_3098000# diff_553000_1211000# diff_4729000_565000# GND efet w=300000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5982 diff_4729000_565000# diff_4503000_546000# diff_83000_3098000# GND efet w=45000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5983 diff_4096000_194000# diff_4088000_123000# diff_83000_3098000# GND efet w=648500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5984 diff_83000_3098000# diff_4088000_123000# diff_4096000_194000# GND efet w=188500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5985 diff_95000_5192000# diff_4162000_585000# diff_4096000_194000# GND efet w=206500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5986 diff_95000_5192000# diff_4162000_585000# diff_4096000_194000# GND efet w=203000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5987 diff_95000_5192000# diff_4162000_585000# diff_4096000_194000# GND efet w=203500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5988 diff_95000_5192000# diff_4162000_585000# diff_4096000_194000# GND efet w=188000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5989 diff_4518000_194000# diff_4503000_546000# diff_95000_5192000# GND efet w=190000 l=8000
+ ad=1.56294e+08 pd=4.562e+06 as=0 ps=0 
M5990 diff_95000_5192000# diff_4503000_546000# diff_4518000_194000# GND efet w=205500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5991 diff_95000_5192000# diff_4162000_585000# diff_4096000_194000# GND efet w=646000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5992 diff_3265000_456000# diff_3332000_585000# diff_95000_5192000# GND efet w=270000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5993 diff_3687000_194000# diff_3673000_545000# diff_95000_5192000# GND efet w=270000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5994 diff_3687000_194000# diff_3899000_565000# diff_83000_3098000# GND efet w=279500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M5995 diff_4096000_194000# diff_4088000_123000# diff_83000_3098000# GND efet w=281000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5996 diff_4518000_194000# diff_4503000_546000# diff_95000_5192000# GND efet w=648000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M5997 diff_95000_5192000# diff_4503000_546000# diff_4518000_194000# GND efet w=205000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5998 diff_95000_5192000# diff_4503000_546000# diff_4518000_194000# GND efet w=210000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M5999 diff_4729000_565000# diff_4729000_565000# diff_95000_5192000# GND efet w=35000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6000 diff_4729000_565000# diff_553000_1211000# diff_83000_3098000# GND efet w=56000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M6001 diff_5009000_805000# diff_4776000_738000# diff_83000_3098000# GND efet w=130500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M6002 diff_83000_3098000# diff_5070000_815000# diff_5009000_805000# GND efet w=136500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M6003 diff_2351000_3074000# diff_2351000_3074000# diff_95000_5192000# GND efet w=18000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M6004 diff_83000_3098000# diff_5123000_886000# diff_2351000_3074000# GND efet w=256500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M6005 diff_5331000_4062000# diff_5331000_4062000# diff_95000_5192000# GND efet w=13000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M6006 diff_4328000_910000# diff_4045000_823000# diff_83000_3098000# GND efet w=71000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M6007 diff_5626000_1299000# diff_72000_4515000# diff_5618000_1133000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=1.04e+09 ps=234000 
M6008 diff_95000_5192000# diff_5626000_1299000# diff_5626000_1299000# GND efet w=13000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M6009 diff_95000_5192000# diff_5769000_1236000# diff_5619000_1309000# GND efet w=779000 l=8000
+ ad=0 pd=0 as=-1.68964e+09 ps=6.926e+06 
M6010 diff_95000_5192000# diff_5651000_1222000# diff_5618000_1133000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M6011 diff_5651000_1222000# diff_5632000_1142000# diff_83000_3098000# GND efet w=47000 l=8000
+ ad=1.163e+09 pd=214000 as=0 ps=0 
M6012 diff_95000_5192000# diff_5769000_1236000# diff_5619000_1309000# GND efet w=286000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6013 diff_5769000_1236000# diff_5697000_957000# diff_83000_3098000# GND efet w=478000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6014 diff_95000_5192000# diff_5651000_1222000# diff_5651000_1222000# GND efet w=12000 l=35000
+ ad=0 pd=0 as=0 ps=0 
M6015 diff_95000_5192000# diff_5769000_1236000# diff_5619000_1309000# GND efet w=285500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M6016 diff_5651000_1222000# diff_72000_4515000# diff_83000_3098000# GND efet w=28000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M6017 diff_5632000_1142000# diff_5618000_1133000# diff_83000_3098000# GND efet w=223500 l=8500
+ ad=-5.06967e+08 pd=730000 as=0 ps=0 
M6018 diff_95000_5192000# diff_5632000_1142000# diff_5632000_1142000# GND efet w=14000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M6019 diff_5619000_1309000# diff_5769000_1236000# diff_95000_5192000# GND efet w=287000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6020 diff_83000_3098000# diff_83000_3098000# diff_5619000_1309000# GND efet w=93500 l=12500
+ ad=0 pd=0 as=0 ps=0 
M6021 diff_5769000_1236000# diff_5769000_1236000# diff_95000_5192000# GND efet w=44000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6022 diff_83000_3098000# diff_5697000_957000# diff_5619000_1309000# GND efet w=239000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6023 diff_95000_5192000# diff_5697000_957000# diff_5697000_957000# GND efet w=33000 l=8000
+ ad=0 pd=0 as=1.97607e+09 ps=1.77e+06 
M6024 diff_5697000_957000# diff_5087000_472000# diff_83000_3098000# GND efet w=475000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6025 diff_5632000_1142000# diff_5011000_576000# diff_817000_1588000# GND efet w=87000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M6026 diff_83000_3098000# diff_5651000_957000# diff_5697000_957000# GND efet w=513000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M6027 diff_817000_1588000# diff_4954000_639000# diff_5651000_957000# GND efet w=35000 l=12000
+ ad=0 pd=0 as=-1.62097e+09 ps=320000 
M6028 diff_83000_3098000# diff_5697000_957000# diff_5619000_1309000# GND efet w=289000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6029 diff_83000_3098000# diff_5697000_957000# diff_5619000_1309000# GND efet w=290000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M6030 diff_5619000_1309000# diff_5697000_957000# diff_83000_3098000# GND efet w=800500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M6031 diff_5696000_939000# diff_5651000_888000# diff_83000_3098000# GND efet w=514000 l=9000
+ ad=1.62107e+09 pd=1.786e+06 as=0 ps=0 
M6032 diff_83000_3098000# diff_5696000_939000# diff_5600000_575000# GND efet w=804000 l=10000
+ ad=0 pd=0 as=-6.2264e+08 ps=7.076e+06 
M6033 diff_83000_3098000# diff_5087000_472000# diff_5696000_939000# GND efet w=475500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M6034 diff_5009000_805000# diff_95000_5192000# diff_95000_5192000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M6035 diff_83000_3098000# diff_5123000_1237000# diff_5070000_815000# GND efet w=55000 l=8000
+ ad=0 pd=0 as=9.19e+08 ps=210000 
M6036 diff_5070000_815000# diff_5070000_815000# diff_95000_5192000# GND efet w=10000 l=36000
+ ad=0 pd=0 as=0 ps=0 
M6037 diff_5387000_800000# diff_5277000_710000# diff_83000_3098000# GND efet w=172500 l=8500
+ ad=-6.61935e+08 pd=1.472e+06 as=0 ps=0 
M6038 diff_5651000_888000# diff_4954000_639000# diff_817000_1286000# GND efet w=35000 l=11000
+ ad=-1.75597e+09 pd=296000 as=0 ps=0 
M6039 diff_83000_3098000# diff_5009000_805000# diff_5387000_800000# GND efet w=164000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M6040 diff_5277000_710000# diff_5123000_1237000# diff_83000_3098000# GND efet w=130500 l=8500
+ ad=-9.16967e+08 pd=632000 as=0 ps=0 
M6041 diff_83000_3098000# diff_4838000_814000# diff_5277000_710000# GND efet w=125500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M6042 diff_817000_909000# diff_4954000_639000# diff_4944000_580000# GND efet w=46000 l=11000
+ ad=0 pd=0 as=2.115e+09 ps=226000 
M6043 diff_5026000_597000# diff_5011000_576000# diff_817000_909000# GND efet w=84000 l=11000
+ ad=-1.59967e+08 pd=570000 as=0 ps=0 
M6044 diff_95000_5192000# diff_5026000_597000# diff_5026000_597000# GND efet w=11000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M6045 diff_5115000_587000# diff_5115000_587000# diff_95000_5192000# GND efet w=14000 l=36000
+ ad=2.142e+09 pd=480000 as=0 ps=0 
M6046 diff_83000_3098000# diff_5039000_607000# diff_5026000_597000# GND efet w=228000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6047 diff_5115000_587000# diff_5026000_597000# diff_83000_3098000# GND efet w=34000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M6048 diff_83000_3098000# diff_72000_4515000# diff_5115000_587000# GND efet w=26000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M6049 diff_95000_5192000# diff_5115000_587000# diff_5039000_607000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=9.86e+08 ps=270000 
M6050 diff_95000_5192000# diff_5213000_615000# diff_5213000_615000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=2.14e+09 ps=434000 
M6051 diff_5213000_615000# diff_72000_4515000# diff_5039000_607000# GND efet w=19000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M6052 diff_5271000_2493000# diff_72000_4515000# diff_83000_3098000# GND efet w=73500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M6053 diff_817000_1286000# diff_5011000_576000# diff_5632000_693000# GND efet w=87000 l=11000
+ ad=0 pd=0 as=-2.99967e+08 ps=736000 
M6054 diff_5632000_693000# diff_5618000_625000# diff_83000_3098000# GND efet w=219500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M6055 diff_83000_3098000# diff_5696000_939000# diff_5600000_575000# GND efet w=289500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M6056 diff_83000_3098000# diff_5696000_939000# diff_5600000_575000# GND efet w=288500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M6057 diff_5696000_939000# diff_5696000_939000# diff_5696000_939000# GND efet w=2000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M6058 diff_5600000_575000# diff_5696000_939000# diff_83000_3098000# GND efet w=238500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M6059 diff_5696000_939000# diff_5696000_939000# diff_95000_5192000# GND efet w=36000 l=7000
+ ad=0 pd=0 as=0 ps=0 
M6060 diff_95000_5192000# diff_95000_5192000# diff_5277000_710000# GND efet w=13000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6061 diff_95000_5192000# diff_5387000_800000# diff_5387000_800000# GND efet w=15000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M6062 diff_95000_5192000# diff_5632000_693000# diff_5632000_693000# GND efet w=13000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M6063 diff_83000_3098000# diff_72000_4515000# diff_5651000_672000# GND efet w=28000 l=9000
+ ad=0 pd=0 as=1.153e+09 ps=214000 
M6064 diff_95000_5192000# diff_5769000_579000# diff_5769000_579000# GND efet w=44000 l=8000
+ ad=0 pd=0 as=1.79107e+09 ps=1.616e+06 
M6065 diff_83000_3098000# diff_5696000_939000# diff_5769000_579000# GND efet w=478000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M6066 diff_5600000_575000# diff_5769000_579000# diff_95000_5192000# GND efet w=285000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6067 diff_95000_5192000# diff_5769000_579000# diff_5600000_575000# GND efet w=285500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M6068 diff_95000_5192000# diff_5651000_672000# diff_5651000_672000# GND efet w=12000 l=35000
+ ad=0 pd=0 as=0 ps=0 
M6069 diff_5651000_672000# diff_5632000_693000# diff_83000_3098000# GND efet w=42500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M6070 diff_95000_5192000# diff_5651000_672000# diff_5618000_625000# GND efet w=12000 l=12000
+ ad=0 pd=0 as=1.099e+09 ps=246000 
M6071 diff_83000_3098000# diff_5087000_472000# diff_5769000_579000# GND efet w=485500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M6072 diff_95000_5192000# diff_5769000_579000# diff_5600000_575000# GND efet w=286000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6073 diff_5618000_625000# diff_72000_4515000# diff_5610000_585000# GND efet w=19000 l=12000
+ ad=0 pd=0 as=-1.98797e+09 ps=396000 
M6074 diff_5213000_615000# diff_4952000_396000# diff_83000_3098000# GND efet w=127000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M6075 diff_83000_3098000# diff_4729000_565000# diff_4518000_194000# GND efet w=192500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M6076 diff_83000_3098000# diff_4729000_565000# diff_4518000_194000# GND efet w=184000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6077 diff_83000_3098000# diff_4729000_565000# diff_4518000_194000# GND efet w=181000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6078 diff_83000_3098000# diff_4729000_565000# diff_4518000_194000# GND efet w=649500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M6079 diff_83000_3098000# diff_4944000_580000# diff_4942000_386000# GND efet w=558500 l=7500
+ ad=0 pd=0 as=-2.79019e+07 ps=1.754e+06 
M6080 diff_95000_5192000# diff_5610000_585000# diff_5610000_585000# GND efet w=12000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M6081 diff_5600000_575000# diff_5769000_579000# diff_95000_5192000# GND efet w=785000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6082 diff_4942000_386000# diff_5087000_472000# diff_83000_3098000# GND efet w=542000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6083 diff_83000_3098000# diff_4942000_386000# diff_5240000_452000# GND efet w=572500 l=8500
+ ad=0 pd=0 as=-4.36902e+08 ps=1.72e+06 
M6084 diff_95000_5192000# diff_4942000_386000# diff_4942000_386000# GND efet w=35000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M6085 diff_5240000_452000# diff_5240000_452000# diff_95000_5192000# GND efet w=45000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6086 diff_83000_3098000# diff_5087000_472000# diff_5240000_452000# GND efet w=532500 l=7500
+ ad=0 pd=0 as=0 ps=0 
M6087 diff_5610000_585000# diff_5600000_575000# diff_83000_3098000# GND efet w=147500 l=10500
+ ad=0 pd=0 as=0 ps=0 
M6088 diff_83000_3098000# diff_83000_3098000# diff_5600000_575000# GND efet w=97000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M6089 diff_4952000_396000# diff_4942000_386000# diff_83000_3098000# GND efet w=241500 l=10500
+ ad=-1.62257e+09 pd=7.482e+06 as=0 ps=0 
M6090 diff_4952000_396000# diff_4942000_386000# diff_83000_3098000# GND efet w=932500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M6091 diff_4096000_194000# diff_4162000_585000# diff_95000_5192000# GND efet w=269000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6092 diff_4518000_194000# diff_4503000_546000# diff_95000_5192000# GND efet w=270000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6093 diff_4518000_194000# diff_4729000_565000# diff_83000_3098000# GND efet w=281000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6094 diff_4952000_396000# diff_4942000_386000# diff_83000_3098000# GND efet w=416000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6095 diff_95000_5192000# diff_5240000_452000# diff_4952000_396000# GND efet w=215000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6096 diff_95000_5192000# diff_5240000_452000# diff_4952000_396000# GND efet w=941000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6097 diff_95000_5192000# diff_5240000_452000# diff_4952000_396000# GND efet w=421500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M6098 diff_5606000_421000# diff_5596000_414000# diff_83000_3098000# GND efet w=143000 l=10000
+ ad=-1.69497e+09 pd=532000 as=0 ps=0 
M6099 diff_5769000_414000# diff_5087000_472000# diff_83000_3098000# GND efet w=485000 l=9000
+ ad=1.36207e+09 pd=1.61e+06 as=0 ps=0 
M6100 diff_5606000_421000# diff_72000_4515000# diff_5618000_311000# GND efet w=20000 l=11000
+ ad=0 pd=0 as=1.076e+09 ps=236000 
M6101 diff_95000_5192000# diff_5606000_421000# diff_5606000_421000# GND efet w=13000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M6102 diff_95000_5192000# diff_5769000_414000# diff_5596000_414000# GND efet w=779000 l=8000
+ ad=0 pd=0 as=6.1236e+08 ps=6.982e+06 
M6103 diff_95000_5192000# diff_5651000_400000# diff_5618000_311000# GND efet w=13000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M6104 diff_5651000_400000# diff_5632000_320000# diff_83000_3098000# GND efet w=47000 l=8000
+ ad=1.14e+09 pd=214000 as=0 ps=0 
M6105 diff_95000_5192000# diff_5769000_414000# diff_5596000_414000# GND efet w=286000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6106 diff_5769000_414000# diff_5697000_135000# diff_83000_3098000# GND efet w=478000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6107 diff_95000_5192000# diff_5651000_400000# diff_5651000_400000# GND efet w=11000 l=35000
+ ad=0 pd=0 as=0 ps=0 
M6108 diff_95000_5192000# diff_5769000_414000# diff_5596000_414000# GND efet w=285500 l=8500
+ ad=0 pd=0 as=0 ps=0 
M6109 diff_5651000_400000# diff_72000_4515000# diff_83000_3098000# GND efet w=28000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M6110 diff_5632000_320000# diff_5618000_311000# diff_83000_3098000# GND efet w=223500 l=8500
+ ad=-5.62967e+08 pd=730000 as=0 ps=0 
M6111 diff_95000_5192000# diff_5632000_320000# diff_5632000_320000# GND efet w=11000 l=21000
+ ad=0 pd=0 as=0 ps=0 
M6112 diff_5596000_414000# diff_5769000_414000# diff_95000_5192000# GND efet w=287000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6113 diff_83000_3098000# diff_83000_3098000# diff_5596000_414000# GND efet w=93000 l=13000
+ ad=0 pd=0 as=0 ps=0 
M6114 diff_5769000_414000# diff_5769000_414000# diff_95000_5192000# GND efet w=44000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6115 diff_83000_3098000# diff_5697000_135000# diff_5596000_414000# GND efet w=239000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6116 diff_95000_5192000# diff_5697000_135000# diff_5697000_135000# GND efet w=33000 l=8000
+ ad=0 pd=0 as=1.97107e+09 ps=1.77e+06 
M6117 diff_5697000_135000# diff_5087000_472000# diff_83000_3098000# GND efet w=475000 l=8000
+ ad=0 pd=0 as=0 ps=0 
M6118 diff_5632000_320000# diff_5011000_576000# diff_817000_1211000# GND efet w=87000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M6119 diff_83000_3098000# diff_5651000_135000# diff_5697000_135000# GND efet w=513000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M6120 diff_817000_1211000# diff_4954000_639000# diff_5651000_135000# GND efet w=34000 l=12000
+ ad=0 pd=0 as=-1.62997e+09 ps=318000 
M6121 diff_83000_3098000# diff_5697000_135000# diff_5596000_414000# GND efet w=289000 l=10000
+ ad=0 pd=0 as=0 ps=0 
M6122 diff_83000_3098000# diff_5697000_135000# diff_5596000_414000# GND efet w=290000 l=11000
+ ad=0 pd=0 as=0 ps=0 
M6123 diff_5596000_414000# diff_5697000_135000# diff_83000_3098000# GND efet w=770500 l=9500
+ ad=0 pd=0 as=0 ps=0 
M6124 diff_83000_3098000# diff_83000_3098000# diff_4952000_396000# GND efet w=98500 l=11500
+ ad=0 pd=0 as=0 ps=0 
C0 diff_5651000_135000# gnd! 550.8fF
C1 diff_5697000_135000# gnd! 2413.8fF
C2 diff_5632000_320000# gnd! 525.4fF
C3 diff_5651000_400000# gnd! 232.7fF
C4 diff_5618000_311000# gnd! 302.1fF
C5 diff_5769000_414000# gnd! 2007.7fF
C6 diff_5606000_421000# gnd! 341.6fF
C7 diff_5240000_452000# gnd! 2353.8fF
C8 diff_4942000_386000# gnd! 2769.2fF
C9 diff_5610000_585000# gnd! 295.1fF
C10 diff_5651000_672000# gnd! 230.9fF
C11 diff_5769000_579000# gnd! 2070.1fF
C12 diff_5632000_693000# gnd! 551.1fF
C13 diff_5618000_625000# gnd! 300.7fF
C14 diff_5213000_615000# gnd! 295.9fF
C15 diff_5039000_607000# gnd! 270.3fF
C16 diff_5115000_587000# gnd! 350.9fF
C17 diff_4944000_580000# gnd! 478.7fF
C18 diff_5026000_597000# gnd! 546.1fF
C19 diff_5277000_710000# gnd! 560.5fF
C20 diff_5696000_939000# gnd! 2434.5fF
C21 diff_5651000_888000# gnd! 536.1fF
C22 diff_5651000_957000# gnd! 551.9fF
C23 diff_5697000_957000# gnd! 2449.8fF
C24 diff_5632000_1142000# gnd! 531.4fF
C25 diff_5651000_1222000# gnd! 235.0fF
C26 diff_5618000_1133000# gnd! 298.2fF
C27 diff_4518000_194000# gnd! 4707.7fF
C28 diff_4729000_565000# gnd! 1948.1fF
C29 diff_4683000_625000# gnd! 476.3fF
C30 diff_4576000_568000# gnd! 314.2fF
C31 diff_4503000_546000# gnd! 2489.2fF
C32 diff_4096000_194000# gnd! 4851.7fF
C33 diff_4312000_568000# gnd! 309.2fF
C34 diff_4227000_613000# gnd! 452.1fF
C35 diff_4162000_585000# gnd! 2484.5fF
C36 diff_3687000_194000# gnd! 4688.1fF
C37 diff_3265000_456000# gnd! 4692.7fF
C38 diff_4088000_123000# gnd! 1936.3fF
C39 diff_3852000_625000# gnd! 476.0fF
C40 diff_3899000_565000# gnd! 2058.2fF
C41 diff_3746000_568000# gnd! 307.4fF
C42 diff_3673000_545000# gnd! 2477.9fF
C43 diff_3482000_568000# gnd! 312.2fF
C44 diff_5009000_805000# gnd! 694.3fF
C45 diff_5070000_815000# gnd! 298.8fF
C46 diff_4776000_738000# gnd! 410.2fF
C47 diff_5769000_1236000# gnd! 1999.2fF
C48 diff_5626000_1299000# gnd! 301.6fF
C49 diff_5626000_1390000# gnd! 264.4fF
C50 diff_5651000_1464000# gnd! 233.2fF
C51 diff_5769000_1368000# gnd! 2012.8fF
C52 diff_5333000_892000# gnd! 24.8fF
C53 diff_5354000_892000# gnd! 134.4fF
C54 diff_5375000_1196000# gnd! 518.3fF
C55 diff_5243000_887000# gnd! 305.4fF
C56 diff_5288000_912000# gnd! 172.6fF
C57 diff_5201000_907000# gnd! 299.6fF
C58 diff_5123000_886000# gnd! 457.1fF
C59 diff_4838000_814000# gnd! 485.4fF
C60 diff_5069000_901000# gnd! 388.1fF
C61 diff_5354000_1225000# gnd! 137.9fF
C62 diff_5334000_1225000# gnd! 22.6fF
C63 diff_4990000_890000# gnd! 861.9fF
C64 diff_4707000_840000# gnd! 376.7fF
C65 diff_4948000_897000# gnd! 218.4fF
C66 diff_4969000_890000# gnd! 231.1fF
C67 diff_5288000_1171000# gnd! 171.6fF
C68 diff_5202000_1210000# gnd! 300.1fF
C69 diff_5243000_1229000# gnd! 301.9fF
C70 diff_4870000_939000# gnd! 575.8fF
C71 diff_5123000_1237000# gnd! 939.8fF
C72 diff_5069000_1218000# gnd! 402.8fF
C73 diff_5334000_1269000# gnd! 20.6fF
C74 diff_5354000_1269000# gnd! 136.4fF
C75 diff_5375000_1305000# gnd! 516.5fF
C76 diff_5632000_1485000# gnd! 554.3fF
C77 diff_5618000_1427000# gnd! 296.6fF
C78 diff_5696000_1731000# gnd! 2454.6fF
C79 diff_5650000_1678000# gnd! 560.2fF
C80 diff_5650000_1749000# gnd! 563.9fF
C81 diff_5375000_1574000# gnd! 517.5fF
C82 diff_5243000_1264000# gnd! 305.2fF
C83 diff_5288000_1289000# gnd! 173.8fF
C84 diff_5201000_1284000# gnd! 296.6fF
C85 diff_4990000_1079000# gnd! 892.7fF
C86 diff_4970000_1104000# gnd! 218.5fF
C87 diff_4950000_1104000# gnd! 177.7fF
C88 diff_4693000_927000# gnd! 595.1fF
C89 diff_4808000_919000# gnd! 262.2fF
C90 diff_4786000_981000# gnd! 228.3fF
C91 diff_4705000_974000# gnd! 397.1fF
C92 diff_4705000_1019000# gnd! 104.9fF
C93 diff_4727000_1006000# gnd! 631.6fF
C94 diff_4871000_1180000# gnd! 457.3fF
C95 diff_5123000_1263000# gnd! 699.7fF
C96 diff_5069000_1278000# gnd! 385.2fF
C97 diff_5354000_1602000# gnd! 137.9fF
C98 diff_5333000_1602000# gnd! 23.8fF
C99 diff_4990000_1273000# gnd! 846.8fF
C100 diff_4951000_1273000# gnd! 164.0fF
C101 diff_4808000_1138000# gnd! 266.2fF
C102 diff_4785000_1099000# gnd! 211.8fF
C103 diff_4608000_946000# gnd! 310.6fF
C104 diff_4705000_1097000# gnd! 105.4fF
C105 diff_4518000_901000# gnd! 328.4fF
C106 diff_4424000_962000# gnd! 312.8fF
C107 diff_4694000_1185000# gnd! 607.6fF
C108 diff_4705000_1142000# gnd! 332.6fF
C109 diff_4727000_1106000# gnd! 561.0fF
C110 diff_4970000_1273000# gnd! 218.1fF
C111 diff_5288000_1548000# gnd! 171.2fF
C112 diff_5202000_1588000# gnd! 299.6fF
C113 diff_5243000_1607000# gnd! 293.6fF
C114 diff_4870000_1328000# gnd! 482.8fF
C115 diff_5123000_1614000# gnd! 691.5fF
C116 diff_5069000_1595000# gnd! 403.5fF
C117 diff_5333000_1645000# gnd! 22.7fF
C118 diff_5697000_1749000# gnd! 2462.2fF
C119 diff_5632000_1934000# gnd! 532.2fF
C120 diff_5651000_2014000# gnd! 235.1fF
C121 diff_5618000_1925000# gnd! 296.6fF
C122 diff_5769000_2028000# gnd! 2016.5fF
C123 diff_5626000_2091000# gnd! 300.9fF
C124 diff_5626000_2182000# gnd! 274.4fF
C125 diff_5651000_2257000# gnd! 237.3fF
C126 diff_5769000_2161000# gnd! 2032.0fF
C127 diff_5354000_1645000# gnd! 134.9fF
C128 diff_5375000_1681000# gnd! 519.5fF
C129 diff_5473000_1600000# gnd! 474.1fF
C130 diff_5375000_1950000# gnd! 518.6fF
C131 diff_5243000_1641000# gnd! 306.2fF
C132 diff_5288000_1666000# gnd! 171.9fF
C133 diff_5201000_1660000# gnd! 298.9fF
C134 diff_4990000_1457000# gnd! 883.1fF
C135 diff_4970000_1482000# gnd! 217.1fF
C136 diff_4950000_1482000# gnd! 176.4fF
C137 diff_4693000_1304000# gnd! 599.2fF
C138 diff_4608000_1093000# gnd! 311.9fF
C139 diff_4518000_1196000# gnd! 340.6fF
C140 diff_4459000_1108000# gnd! 500.1fF
C141 diff_3396000_614000# gnd! 460.1fF
C142 diff_2458000_131000# gnd! 4727.3fF
C143 diff_3332000_585000# gnd! 2488.9fF
C144 diff_3258000_123000# gnd! 1906.4fF
C145 diff_2674000_568000# gnd! 315.1fF
C146 diff_2589000_613000# gnd! 449.2fF
C147 diff_2524000_585000# gnd! 2490.8fF
C148 diff_2049000_194000# gnd! 4678.1fF
C149 diff_1627000_456000# gnd! 4698.1fF
C150 diff_2450000_123000# gnd! 1933.2fF
C151 diff_2261000_565000# gnd! 1935.8fF
C152 diff_2214000_625000# gnd! 468.4fF
C153 diff_2108000_568000# gnd! 305.0fF
C154 diff_2035000_545000# gnd! 2481.0fF
C155 diff_1844000_568000# gnd! 317.4fF
C156 diff_4045000_823000# gnd! 668.5fF
C157 diff_4432000_1144000# gnd! 287.9fF
C158 diff_4459000_1183000# gnd! 392.5fF
C159 diff_4808000_1269000# gnd! 259.3fF
C160 diff_4786000_1406000# gnd! 218.7fF
C161 diff_4705000_1351000# gnd! 342.3fF
C162 diff_4727000_1383000# gnd! 548.5fF
C163 diff_4705000_1396000# gnd! 104.0fF
C164 diff_4871000_1557000# gnd! 463.9fF
C165 diff_5123000_1641000# gnd! 491.5fF
C166 diff_5069000_1655000# gnd! 381.9fF
C167 diff_5354000_1978000# gnd! 138.8fF
C168 diff_5334000_1978000# gnd! 22.6fF
C169 diff_5288000_1925000# gnd! 170.1fF
C170 diff_4990000_1651000# gnd! 850.2fF
C171 diff_4951000_1651000# gnd! 164.0fF
C172 diff_4808000_1515000# gnd! 267.6fF
C173 diff_4786000_1476000# gnd! 223.8fF
C174 diff_4608000_1323000# gnd! 309.6fF
C175 diff_4705000_1475000# gnd! 103.5fF
C176 diff_4518000_1278000# gnd! 330.3fF
C177 diff_4432000_1237000# gnd! 357.8fF
C178 diff_4307000_1010000# gnd! 133.5fF
C179 diff_4036000_920000# gnd! 166.8fF
C180 diff_4057000_1020000# gnd! 254.9fF
C181 diff_4307000_1187000# gnd! 539.9fF
C182 diff_4066000_1028000# gnd! 636.7fF
C183 diff_4225000_1221000# gnd! 477.2fF
C184 diff_4318000_999000# gnd! 336.5fF
C185 diff_4694000_1563000# gnd! 606.0fF
C186 diff_4705000_1519000# gnd! 332.3fF
C187 diff_4727000_1483000# gnd! 564.4fF
C188 diff_4970000_1651000# gnd! 218.5fF
C189 diff_5202000_1964000# gnd! 301.2fF
C190 diff_5243000_1983000# gnd! 298.2fF
C191 diff_4870000_1705000# gnd! 482.8fF
C192 diff_5069000_1972000# gnd! 392.9fF
C193 diff_5123000_1992000# gnd! 695.8fF
C194 diff_5159000_1628000# gnd! 1041.2fF
C195 diff_5632000_2276000# gnd! 559.2fF
C196 diff_5618000_2219000# gnd! 287.8fF
C197 diff_5696000_2524000# gnd! 2414.8fF
C198 diff_5651000_2472000# gnd! 542.0fF
C199 diff_5334000_2022000# gnd! 20.6fF
C200 diff_5354000_2022000# gnd! 136.1fF
C201 diff_5375000_2058000# gnd! 519.1fF
C202 diff_5375000_2327000# gnd! 519.5fF
C203 diff_5243000_2018000# gnd! 310.4fF
C204 diff_5288000_2043000# gnd! 173.4fF
C205 diff_5201000_2038000# gnd! 298.6fF
C206 diff_4990000_1834000# gnd! 887.7fF
C207 diff_4970000_1859000# gnd! 218.5fF
C208 diff_4950000_1859000# gnd! 177.7fF
C209 diff_4693000_1681000# gnd! 593.1fF
C210 diff_4608000_1471000# gnd! 315.5fF
C211 diff_4518000_1573000# gnd! 335.7fF
C212 diff_4458000_1491000# gnd! 506.4fF
C213 diff_4434000_1491000# gnd! 271.2fF
C214 diff_4459000_1639000# gnd! 412.4fF
C215 diff_4808000_1647000# gnd! 266.5fF
C216 diff_4786000_1782000# gnd! 232.2fF
C217 diff_4727000_1761000# gnd! 555.9fF
C218 diff_4705000_1728000# gnd! 340.3fF
C219 diff_4705000_1773000# gnd! 104.9fF
C220 diff_4871000_1932000# gnd! 466.7fF
C221 diff_5123000_2018000# gnd! 700.1fF
C222 diff_5069000_2032000# gnd! 386.8fF
C223 diff_5354000_2356000# gnd! 137.5fF
C224 diff_5333000_2356000# gnd! 26.0fF
C225 diff_4990000_2028000# gnd! 850.0fF
C226 diff_4951000_2028000# gnd! 164.0fF
C227 diff_4808000_1891000# gnd! 267.7fF
C228 diff_4786000_1853000# gnd! 224.0fF
C229 diff_4608000_1700000# gnd! 311.8fF
C230 diff_4705000_1851000# gnd! 105.3fF
C231 diff_4518000_1655000# gnd! 332.2fF
C232 diff_4430000_1714000# gnd! 349.2fF
C233 diff_4261000_1288000# gnd! 665.3fF
C234 diff_4066000_1098000# gnd! 632.0fF
C235 diff_3939000_927000# gnd! 157.1fF
C236 diff_3846000_946000# gnd! 521.5fF
C237 diff_3902000_1041000# gnd! 251.1fF
C238 diff_4057000_1091000# gnd! 256.8fF
C239 diff_4036000_1196000# gnd! 169.2fF
C240 diff_3902000_1074000# gnd! 252.1fF
C241 diff_3696000_1028000# gnd! 514.0fF
C242 diff_3687000_935000# gnd! 252.7fF
C243 diff_3938000_1186000# gnd! 164.8fF
C244 diff_4241000_1304000# gnd! 171.0fF
C245 diff_4694000_1940000# gnd! 595.7fF
C246 diff_4727000_1861000# gnd! 558.5fF
C247 diff_4705000_1896000# gnd! 331.6fF
C248 diff_4970000_2028000# gnd! 218.5fF
C249 diff_5288000_2302000# gnd! 171.3fF
C250 diff_5202000_2342000# gnd! 302.1fF
C251 diff_5243000_2360000# gnd! 294.5fF
C252 diff_4870000_2082000# gnd! 477.5fF
C253 diff_5069000_2349000# gnd! 400.5fF
C254 diff_5123000_2369000# gnd! 686.5fF
C255 diff_5651000_2541000# gnd! 553.9fF
C256 diff_5697000_2542000# gnd! 2458.7fF
C257 diff_5632000_2727000# gnd! 524.4fF
C258 diff_5651000_2807000# gnd! 231.4fF
C259 diff_5618000_2718000# gnd! 301.1fF
C260 diff_5626000_2884000# gnd! 294.7fF
C261 diff_5769000_2821000# gnd! 1985.8fF
C262 diff_6213000_3183000# gnd! 335.0fF
C263 diff_4990000_2211000# gnd! 884.4fF
C264 diff_4970000_2236000# gnd! 217.0fF
C265 diff_4950000_2236000# gnd! 176.4fF
C266 diff_4693000_2058000# gnd! 600.0fF
C267 diff_4608000_1847000# gnd! 314.2fF
C268 diff_4518000_1950000# gnd! 337.1fF
C269 diff_4459000_1862000# gnd! 522.4fF
C270 diff_4434000_1906000# gnd! 281.9fF
C271 diff_4459000_2026000# gnd! 418.4fF
C272 diff_4808000_2024000# gnd! 264.8fF
C273 diff_4786000_2160000# gnd! 231.3fF
C274 diff_4705000_2105000# gnd! 337.1fF
C275 diff_4727000_2138000# gnd! 552.5fF
C276 diff_4705000_2151000# gnd! 102.5fF
C277 diff_5142000_2400000# gnd! 814.5fF
C278 diff_5122000_2495000# gnd! 528.7fF
C279 diff_4871000_2311000# gnd! 463.5fF
C280 diff_4808000_2269000# gnd! 267.6fF
C281 diff_4786000_2230000# gnd! 223.8fF
C282 diff_4608000_2077000# gnd! 313.5fF
C283 diff_4705000_2229000# gnd! 102.6fF
C284 diff_4518000_2032000# gnd! 330.8fF
C285 diff_4433000_2037000# gnd! 393.7fF
C286 diff_4694000_2317000# gnd! 607.1fF
C287 diff_4705000_2274000# gnd! 336.3fF
C288 diff_4727000_2238000# gnd! 560.3fF
C289 diff_5187000_2412000# gnd! 537.2fF
C290 diff_5011000_576000# gnd! 2089.9fF
C291 diff_5271000_2493000# gnd! 1549.2fF
C292 diff_5114000_2490000# gnd! 179.6fF
C293 diff_4994000_2634000# gnd! 969.8fF
C294 diff_4932000_827000# gnd! 1560.5fF
C295 diff_5012000_2755000# gnd! 220.1fF
C296 diff_4959000_2608000# gnd! 307.2fF
C297 diff_5318000_2778000# gnd! 255.8fF
C298 diff_5265000_2778000# gnd! 224.2fF
C299 diff_5170000_2830000# gnd! 211.2fF
C300 diff_4945000_2494000# gnd! 598.9fF
C301 diff_4608000_2224000# gnd! 316.8fF
C302 diff_4575000_2328000# gnd! 265.9fF
C303 diff_4518000_2327000# gnd! 334.8fF
C304 diff_4459000_2246000# gnd! 502.0fF
C305 diff_4768000_996000# gnd! 1275.6fF
C306 diff_4839000_2618000# gnd! 1168.8fF
C307 diff_4883000_2653000# gnd! 256.5fF
C308 diff_4805000_2759000# gnd! 332.6fF
C309 diff_4837000_2758000# gnd! 273.8fF
C310 diff_4740000_2641000# gnd! 940.0fF
C311 diff_4760000_2748000# gnd! 226.6fF
C312 diff_4705000_2611000# gnd! 353.0fF
C313 diff_4433000_2246000# gnd! 292.0fF
C314 diff_4253000_1284000# gnd! 366.1fF
C315 diff_4266000_1501000# gnd! 123.2fF
C316 diff_4036000_1297000# gnd! 166.8fF
C317 diff_4066000_1405000# gnd! 587.9fF
C318 diff_4057000_1397000# gnd! 256.3fF
C319 diff_4285000_1501000# gnd! 638.5fF
C320 diff_4275000_1613000# gnd! 240.1fF
C321 diff_4066000_1475000# gnd! 661.0fF
C322 diff_3846000_1128000# gnd! 535.7fF
C323 diff_3939000_1303000# gnd! 160.2fF
C324 diff_3846000_1323000# gnd! 525.7fF
C325 diff_3696000_1098000# gnd! 523.1fF
C326 diff_3631000_947000# gnd! 217.8fF
C327 diff_3577000_991000# gnd! 1156.4fF
C328 diff_3686000_1185000# gnd! 258.0fF
C329 diff_3632000_1169000# gnd! 214.3fF
C330 diff_3902000_1418000# gnd! 255.8fF
C331 diff_3696000_1405000# gnd! 504.0fF
C332 diff_3687000_1311000# gnd! 258.0fF
C333 diff_4057000_1467000# gnd! 258.4fF
C334 diff_4226000_1649000# gnd! 425.3fF
C335 diff_4037000_1573000# gnd! 166.3fF
C336 diff_3902000_1451000# gnd! 253.7fF
C337 diff_3938000_1563000# gnd! 162.0fF
C338 diff_4235000_1886000# gnd! 303.2fF
C339 diff_4037000_1674000# gnd! 166.1fF
C340 diff_4066000_1783000# gnd! 576.9fF
C341 diff_4057000_1774000# gnd! 255.6fF
C342 diff_4328000_910000# gnd! 1555.4fF
C343 diff_4548000_2725000# gnd! 1343.9fF
C344 diff_4498000_2492000# gnd! 1418.1fF
C345 diff_4417000_952000# gnd! 1320.7fF
C346 diff_4374000_833000# gnd! 1437.5fF
C347 diff_4602000_2752000# gnd! 1731.1fF
C348 diff_4546000_2778000# gnd! 229.8fF
C349 diff_4494000_2778000# gnd! 218.2fF
C350 diff_4443000_2778000# gnd! 227.8fF
C351 diff_4391000_2778000# gnd! 224.8fF
C352 diff_4785000_2783000# gnd! 270.8fF
C353 diff_4689000_2592000# gnd! 259.9fF
C354 diff_4932000_2482000# gnd! 135.4fF
C355 diff_6252000_3157000# gnd! 620.1fF
C356 diff_6269000_3282000# gnd! 159.2fF
C357 diff_6269000_3300000# gnd! 145.9fF
C358 diff_4954000_639000# gnd! 1329.5fF
C359 diff_5214000_3050000# gnd! 410.5fF
C360 diff_5010000_3006000# gnd! 143.7fF
C361 diff_4912000_2900000# gnd! 318.4fF
C362 diff_4975000_2910000# gnd! 237.8fF
C363 diff_5019000_2993000# gnd! 132.3fF
C364 diff_5576000_3241000# gnd! 95.7fF
C365 diff_5084000_3006000# gnd! 159.2fF
C366 diff_5469000_3309000# gnd! 100.8fF
C367 diff_6180000_3356000# gnd! 371.9fF
C368 diff_6120000_3397000# gnd! 239.4fF
C369 diff_5531000_3344000# gnd! 118.9fF
C370 diff_5407000_3340000# gnd! 164.7fF
C371 diff_6006000_3447000# gnd! 95.3fF
C372 diff_6160000_3457000# gnd! 102.8fF
C373 diff_4966000_3079000# gnd! 145.9fF
C374 diff_4983000_2920000# gnd! 772.0fF
C375 diff_4904000_3051000# gnd! 200.0fF
C376 diff_4923000_2911000# gnd! 206.9fF
C377 diff_4843000_3067000# gnd! 759.8fF
C378 diff_4865000_3205000# gnd! 91.7fF
C379 diff_4843000_3181000# gnd! 108.2fF
C380 diff_4777000_2951000# gnd! 500.7fF
C381 diff_4066000_1853000# gnd! 587.1fF
C382 diff_3846000_1504000# gnd! 529.8fF
C383 diff_3939000_1680000# gnd! 159.7fF
C384 diff_3846000_1700000# gnd! 527.1fF
C385 diff_3696000_1475000# gnd! 514.6fF
C386 diff_3436000_1028000# gnd! 533.1fF
C387 diff_3428000_935000# gnd! 249.0fF
C388 diff_3374000_929000# gnd! 277.9fF
C389 diff_3577000_1134000# gnd! 1139.0fF
C390 diff_3632000_1324000# gnd! 214.2fF
C391 diff_3436000_1099000# gnd! 541.7fF
C392 diff_3427000_1189000# gnd! 248.9fF
C393 diff_3374000_1153000# gnd! 278.2fF
C394 diff_1758000_613000# gnd! 462.4fF
C395 diff_1694000_585000# gnd! 2492.9fF
C396 diff_692000_115000# gnd! 232.7fF
C397 diff_174000_153000# gnd! 2258.7fF
C398 diff_1218000_195000# gnd! 4670.2fF
C399 diff_1620000_123000# gnd! 1919.0fF
C400 diff_1430000_565000# gnd! 1937.6fF
C401 diff_1383000_625000# gnd! 475.6fF
C402 diff_1277000_568000# gnd! 300.1fF
C403 diff_1204000_546000# gnd! 2467.2fF
C404 diff_801000_364000# gnd! 4474.8fF
C405 diff_135000_355000# gnd! 3173.7fF
C406 diff_126000_347000# gnd! 2147.8fF
C407 diff_969000_456000# gnd! 2187.2fF
C408 diff_3117000_1023000# gnd! 491.6fF
C409 diff_3099000_927000# gnd! 266.3fF
C410 diff_3577000_1368000# gnd! 1147.5fF
C411 diff_3686000_1562000# gnd! 261.8fF
C412 diff_3632000_1546000# gnd! 214.1fF
C413 diff_3902000_1795000# gnd! 256.5fF
C414 diff_3696000_1783000# gnd! 510.9fF
C415 diff_3687000_1689000# gnd! 259.5fF
C416 diff_4057000_1845000# gnd! 259.9fF
C417 diff_4036000_1950000# gnd! 168.4fF
C418 diff_3902000_1829000# gnd! 256.1fF
C419 diff_3938000_1940000# gnd! 164.1fF
C420 diff_4036000_2051000# gnd! 166.9fF
C421 diff_4066000_2160000# gnd! 649.6fF
C422 diff_4057000_2151000# gnd! 255.2fF
C423 diff_4066000_2230000# gnd! 511.7fF
C424 diff_3846000_1881000# gnd! 531.4fF
C425 diff_3939000_2058000# gnd! 160.3fF
C426 diff_3846000_2078000# gnd! 525.2fF
C427 diff_3696000_1853000# gnd! 521.5fF
C428 diff_3436000_1405000# gnd! 525.1fF
C429 diff_3428000_1309000# gnd! 251.1fF
C430 diff_3374000_1306000# gnd! 277.1fF
C431 diff_3117000_1087000# gnd! 506.6fF
C432 diff_3099000_1189000# gnd! 263.6fF
C433 diff_3029000_910000# gnd! 303.1fF
C434 diff_3577000_1511000# gnd! 1128.3fF
C435 diff_3632000_1701000# gnd! 213.8fF
C436 diff_3436000_1476000# gnd! 527.5fF
C437 diff_3427000_1566000# gnd! 250.7fF
C438 diff_3374000_1530000# gnd! 279.5fF
C439 diff_3029000_1168000# gnd! 303.4fF
C440 diff_3117000_1400000# gnd! 488.3fF
C441 diff_3099000_1304000# gnd! 259.1fF
C442 diff_3577000_1746000# gnd! 1137.5fF
C443 diff_3686000_1940000# gnd! 262.6fF
C444 diff_3632000_1923000# gnd! 214.4fF
C445 diff_3902000_2172000# gnd! 254.8fF
C446 diff_4057000_2222000# gnd! 259.6fF
C447 diff_4037000_2327000# gnd! 169.1fF
C448 diff_3902000_2206000# gnd! 257.2fF
C449 diff_3696000_2160000# gnd! 500.6fF
C450 diff_3687000_2066000# gnd! 258.1fF
C451 diff_3938000_2317000# gnd! 162.2fF
C452 diff_3846000_2258000# gnd! 528.2fF
C453 diff_3696000_2230000# gnd! 515.5fF
C454 diff_3436000_1783000# gnd! 521.7fF
C455 diff_3428000_1687000# gnd! 252.0fF
C456 diff_3374000_1683000# gnd! 279.6fF
C457 diff_3577000_1888000# gnd! 1137.7fF
C458 diff_3632000_2078000# gnd! 210.0fF
C459 diff_3436000_1854000# gnd! 533.0fF
C460 diff_3427000_1944000# gnd! 252.6fF
C461 diff_3374000_1907000# gnd! 279.1fF
C462 diff_3577000_2123000# gnd! 1126.4fF
C463 diff_3686000_2317000# gnd! 264.1fF
C464 diff_3632000_2301000# gnd! 213.9fF
C465 diff_4155000_2676000# gnd! 620.0fF
C466 diff_4277000_2781000# gnd! 591.0fF
C467 diff_4224000_2739000# gnd! 606.3fF
C468 diff_3436000_2160000# gnd! 534.3fF
C469 diff_3428000_2064000# gnd! 250.6fF
C470 diff_3374000_2060000# gnd! 277.7fF
C471 diff_3577000_2265000# gnd! 1160.7fF
C472 diff_3436000_2231000# gnd! 538.0fF
C473 diff_3374000_2284000# gnd! 278.8fF
C474 diff_3427000_2321000# gnd! 253.1fF
C475 diff_3117000_1464000# gnd! 500.2fF
C476 diff_3099000_1566000# gnd! 265.1fF
C477 diff_2915000_927000# gnd! 240.7fF
C478 diff_2876000_1039000# gnd! 260.1fF
C479 diff_2829000_939000# gnd! 516.0fF
C480 diff_2650000_947000# gnd! 132.0fF
C481 diff_2683000_1022000# gnd! 516.7fF
C482 diff_2674000_1013000# gnd! 263.9fF
C483 diff_2876000_1074000# gnd! 257.7fF
C484 diff_2915000_1188000# gnd! 241.5fF
C485 diff_2102000_884000# gnd! 19.4fF
C486 diff_2531000_969000# gnd! 241.0fF
C487 diff_2829000_1111000# gnd! 525.5fF
C488 diff_3029000_1287000# gnd! 295.6fF
C489 diff_3029000_1546000# gnd! 305.8fF
C490 diff_3117000_1777000# gnd! 489.9fF
C491 diff_3099000_1681000# gnd! 258.8fF
C492 diff_3117000_1841000# gnd! 505.1fF
C493 diff_3099000_1943000# gnd! 262.8fF
C494 diff_2914000_1304000# gnd! 242.7fF
C495 diff_2876000_1416000# gnd! 259.0fF
C496 diff_2829000_1316000# gnd! 513.8fF
C497 diff_2409000_958000# gnd! 143.0fF
C498 diff_2683000_1084000# gnd! 519.6fF
C499 diff_2651000_1168000# gnd! 134.6fF
C500 diff_2674000_1077000# gnd! 263.6fF
C501 diff_2531000_1102000# gnd! 230.8fF
C502 diff_2471000_1074000# gnd! 141.8fF
C503 diff_2460000_1079000# gnd! 199.9fF
C504 diff_2406000_1192000# gnd! 183.1fF
C505 diff_2335000_1127000# gnd! 393.2fF
C506 diff_2650000_1323000# gnd! 135.2fF
C507 diff_2683000_1400000# gnd! 496.4fF
C508 diff_2674000_1391000# gnd! 266.8fF
C509 diff_2876000_1451000# gnd! 257.7fF
C510 diff_2915000_1565000# gnd! 244.2fF
C511 diff_2290000_1091000# gnd! 277.1fF
C512 diff_2531000_1389000# gnd! 227.7fF
C513 diff_2459000_1348000# gnd! 208.6fF
C514 diff_2406000_1315000# gnd! 182.5fF
C515 diff_2335000_1372000# gnd! 410.4fF
C516 diff_2184000_926000# gnd! 268.2fF
C517 diff_2121000_884000# gnd! 402.9fF
C518 diff_2130000_913000# gnd! 453.7fF
C519 diff_2137000_920000# gnd! 225.7fF
C520 diff_2127000_952000# gnd! 551.6fF
C521 diff_2184000_1118000# gnd! 270.1fF
C522 diff_2137000_1204000# gnd! 218.7fF
C523 diff_2130000_1219000# gnd! 421.0fF
C524 diff_2050000_1017000# gnd! 142.8fF
C525 diff_1997000_985000# gnd! 462.1fF
C526 diff_1931000_949000# gnd! 167.4fF
C527 diff_1850000_941000# gnd! 507.5fF
C528 diff_1851000_999000# gnd! 1694.0fF
C529 diff_1881000_1041000# gnd! 273.1fF
C530 diff_2102000_1230000# gnd! 20.3fF
C531 diff_2050000_1081000# gnd! 140.7fF
C532 diff_2121000_1230000# gnd! 387.7fF
C533 diff_2127000_1169000# gnd! 639.4fF
C534 diff_2290000_1294000# gnd! 295.9fF
C535 diff_2471000_1358000# gnd! 142.1fF
C536 diff_2829000_1488000# gnd! 525.7fF
C537 diff_3029000_1664000# gnd! 296.4fF
C538 diff_3029000_1923000# gnd! 305.6fF
C539 diff_3117000_2154000# gnd! 482.1fF
C540 diff_3099000_2059000# gnd! 258.6fF
C541 diff_3117000_2217000# gnd! 503.0fF
C542 diff_3099000_2319000# gnd! 261.2fF
C543 diff_2914000_1681000# gnd! 243.9fF
C544 diff_2829000_1693000# gnd! 516.8fF
C545 diff_2683000_1461000# gnd! 506.2fF
C546 diff_2651000_1545000# gnd! 133.1fF
C547 diff_2674000_1454000# gnd! 263.2fF
C548 diff_2531000_1479000# gnd! 227.4fF
C549 diff_2876000_1793000# gnd! 261.6fF
C550 diff_2471000_1451000# gnd! 135.4fF
C551 diff_2459000_1456000# gnd! 209.4fF
C552 diff_2407000_1569000# gnd! 182.4fF
C553 diff_2335000_1514000# gnd! 409.2fF
C554 diff_2651000_1700000# gnd! 131.4fF
C555 diff_2683000_1777000# gnd! 505.3fF
C556 diff_2674000_1768000# gnd! 264.1fF
C557 diff_2876000_1829000# gnd! 256.3fF
C558 diff_2915000_1942000# gnd! 245.8fF
C559 diff_2291000_1482000# gnd! 245.1fF
C560 diff_2531000_1766000# gnd! 224.3fF
C561 diff_2460000_1725000# gnd! 198.5fF
C562 diff_2407000_1692000# gnd! 181.1fF
C563 diff_2471000_1736000# gnd! 138.9fF
C564 diff_2829000_1865000# gnd! 531.0fF
C565 diff_3029000_2041000# gnd! 297.8fF
C566 diff_3029000_2300000# gnd! 304.6fF
C567 diff_2914000_2058000# gnd! 244.2fF
C568 diff_2876000_2170000# gnd! 254.4fF
C569 diff_2829000_2070000# gnd! 516.8fF
C570 diff_2683000_1839000# gnd! 516.4fF
C571 diff_2650000_1921000# gnd! 137.9fF
C572 diff_2674000_1831000# gnd! 266.4fF
C573 diff_2531000_1855000# gnd! 227.9fF
C574 diff_2471000_1828000# gnd! 139.8fF
C575 diff_2460000_1833000# gnd! 201.3fF
C576 diff_2102000_1261000# gnd! 19.4fF
C577 diff_2184000_1302000# gnd! 267.4fF
C578 diff_2121000_1261000# gnd! 398.8fF
C579 diff_2130000_1289000# gnd! 407.0fF
C580 diff_2137000_1296000# gnd! 231.2fF
C581 diff_2127000_1328000# gnd! 698.9fF
C582 diff_2184000_1494000# gnd! 267.9fF
C583 diff_2137000_1580000# gnd! 222.5fF
C584 diff_2130000_1595000# gnd! 420.5fF
C585 diff_1997000_1091000# gnd! 445.9fF
C586 diff_1881000_1073000# gnd! 265.6fF
C587 diff_1851000_1079000# gnd! 1913.7fF
C588 diff_1932000_1177000# gnd! 176.1fF
C589 diff_1850000_1158000# gnd! 520.5fF
C590 diff_2050000_1393000# gnd! 139.6fF
C591 diff_1997000_1362000# gnd! 460.6fF
C592 diff_1932000_1328000# gnd! 169.8fF
C593 diff_1851000_1317000# gnd! 517.0fF
C594 diff_1851000_1376000# gnd! 1860.2fF
C595 diff_1881000_1418000# gnd! 275.1fF
C596 diff_2102000_1607000# gnd! 20.3fF
C597 diff_2050000_1457000# gnd! 141.7fF
C598 diff_2122000_1607000# gnd! 385.6fF
C599 diff_2102000_1637000# gnd! 20.3fF
C600 diff_2127000_1545000# gnd! 699.9fF
C601 diff_2330000_1775000# gnd! 438.6fF
C602 diff_2406000_1946000# gnd! 183.1fF
C603 diff_2651000_2077000# gnd! 131.3fF
C604 diff_2683000_2153000# gnd! 511.5fF
C605 diff_2674000_2144000# gnd! 259.9fF
C606 diff_2876000_2205000# gnd! 258.7fF
C607 diff_2915000_2318000# gnd! 245.0fF
C608 diff_2532000_2143000# gnd! 223.0fF
C609 diff_2829000_2242000# gnd! 531.9fF
C610 diff_4108000_2725000# gnd! 1386.8fF
C611 diff_3800000_830000# gnd! 1564.8fF
C612 diff_4004000_2725000# gnd! 560.8fF
C613 diff_3922000_786000# gnd! 578.3fF
C614 diff_3901000_2725000# gnd! 1463.3fF
C615 diff_3830000_787000# gnd! 1451.3fF
C616 diff_3739000_826000# gnd! 1549.5fF
C617 diff_3749000_2434000# gnd! 1470.4fF
C618 diff_3695000_2725000# gnd! 1650.7fF
C619 diff_3596000_2395000# gnd! 1470.8fF
C620 diff_3567000_785000# gnd! 1464.8fF
C621 diff_3474000_792000# gnd! 1498.5fF
C622 diff_3489000_2725000# gnd! 859.3fF
C623 diff_3439000_2492000# gnd! 1550.4fF
C624 diff_3354000_2409000# gnd! 2287.9fF
C625 diff_4104000_2778000# gnd! 232.3fF
C626 diff_4052000_2778000# gnd! 232.3fF
C627 diff_4001000_2778000# gnd! 232.4fF
C628 diff_3949000_2778000# gnd! 232.1fF
C629 diff_3898000_2778000# gnd! 227.8fF
C630 diff_3846000_2778000# gnd! 229.7fF
C631 diff_3794000_2778000# gnd! 227.2fF
C632 diff_3742000_2778000# gnd! 233.5fF
C633 diff_3692000_2778000# gnd! 229.9fF
C634 diff_3639000_2778000# gnd! 232.2fF
C635 diff_3589000_2778000# gnd! 218.3fF
C636 diff_3536000_2778000# gnd! 225.8fF
C637 diff_3486000_2778000# gnd! 229.7fF
C638 diff_3433000_2778000# gnd! 227.8fF
C639 diff_3383000_2778000# gnd! 229.7fF
C640 diff_4517000_3010000# gnd! 225.0fF
C641 diff_4656000_3020000# gnd! 932.0fF
C642 diff_4779000_3198000# gnd! 156.6fF
C643 diff_5439000_3442000# gnd! 108.5fF
C644 diff_5920000_3449000# gnd! 358.9fF
C645 diff_5432000_3451000# gnd! 144.2fF
C646 diff_5578000_3393000# gnd! 139.3fF
C647 diff_6160000_3507000# gnd! 88.6fF
C648 diff_5294000_3449000# gnd! 177.2fF
C649 diff_5472000_3486000# gnd! 95.6fF
C650 diff_5357000_3322000# gnd! 620.9fF
C651 diff_6112000_3388000# gnd! 535.8fF
C652 diff_6185000_3575000# gnd! 296.4fF
C653 diff_6185000_3600000# gnd! 159.1fF
C654 diff_6017000_3581000# gnd! 318.6fF
C655 diff_5660000_3640000# gnd! 87.2fF
C656 diff_5504000_3630000# gnd! 107.6fF
C657 diff_5513000_3639000# gnd! 156.1fF
C658 diff_5397000_3644000# gnd! 107.9fF
C659 diff_5228000_3587000# gnd! 746.2fF
C660 diff_4871000_3351000# gnd! 883.5fF
C661 diff_5022000_3615000# gnd! 95.8fF
C662 diff_5397000_3662000# gnd! 596.6fF
C663 diff_6146000_3754000# gnd! 346.2fF
C664 diff_6155000_3780000# gnd! 96.4fF
C665 diff_5397000_3688000# gnd! 110.4fF
C666 diff_5293000_3706000# gnd! 124.5fF
C667 diff_5491000_3760000# gnd! 97.5fF
C668 diff_5043000_3671000# gnd! 260.9fF
C669 diff_6155000_3762000# gnd! 367.1fF
C670 diff_6161000_3828000# gnd! 250.2fF
C671 diff_6151000_3839000# gnd! 354.6fF
C672 diff_5501000_3768000# gnd! 116.9fF
C673 diff_5678000_3740000# gnd! 114.5fF
C674 diff_5501000_3807000# gnd! 114.0fF
C675 diff_5039000_3682000# gnd! 241.5fF
C676 diff_5048000_3693000# gnd! 1144.3fF
C677 diff_4591000_3170000# gnd! 682.2fF
C678 diff_4462000_2971000# gnd! 146.1fF
C679 diff_4453000_3015000# gnd! 217.4fF
C680 diff_4435000_3015000# gnd! 237.2fF
C681 diff_4363000_2478000# gnd! 923.4fF
C682 diff_4278000_3058000# gnd! 151.0fF
C683 diff_4627000_3380000# gnd! 236.4fF
C684 diff_4994000_3787000# gnd! 80.5fF
C685 diff_6076000_3942000# gnd! 601.3fF
C686 diff_5983000_3917000# gnd! 484.6fF
C687 diff_5625000_3936000# gnd! 144.8fF
C688 diff_5988000_3969000# gnd! 403.1fF
C689 diff_5696000_3194000# gnd! 791.2fF
C690 diff_6196000_3985000# gnd! 354.9fF
C691 diff_5996000_3977000# gnd! 526.9fF
C692 diff_4997000_3824000# gnd! 201.6fF
C693 diff_4973000_3834000# gnd! 69.3fF
C694 diff_5321000_3744000# gnd! 243.8fF
C695 diff_5228000_3879000# gnd! 756.3fF
C696 diff_4973000_3872000# gnd! 216.8fF
C697 diff_5263000_3933000# gnd! 154.4fF
C698 diff_5067000_3914000# gnd! 195.2fF
C699 diff_4975000_3889000# gnd! 86.5fF
C700 diff_5264000_3945000# gnd! 246.3fF
C701 diff_5274000_3953000# gnd! 386.5fF
C702 diff_5080000_3926000# gnd! 104.9fF
C703 diff_4814000_3335000# gnd! 405.7fF
C704 diff_4716000_3243000# gnd! 406.5fF
C705 diff_5061000_3959000# gnd! 589.4fF
C706 diff_5625000_3954000# gnd! 406.6fF
C707 diff_5612000_4010000# gnd! 408.0fF
C708 diff_5850000_3991000# gnd! 508.1fF
C709 diff_5008000_3739000# gnd! 558.9fF
C710 diff_5356000_4035000# gnd! 154.4fF
C711 diff_5356000_4053000# gnd! 159.1fF
C712 diff_5356000_4071000# gnd! 1176.2fF
C713 diff_5331000_4062000# gnd! 2715.0fF
C714 diff_5371000_3654000# gnd! 1960.5fF
C715 diff_5055000_4064000# gnd! 76.5fF
C716 diff_5029000_4064000# gnd! 230.8fF
C717 diff_5918000_4120000# gnd! 747.5fF
C718 diff_5763000_4184000# gnd! 697.0fF
C719 diff_6179000_4193000# gnd! 337.2fF
C720 diff_6158000_4243000# gnd! 87.6fF
C721 diff_5674000_4156000# gnd! 364.8fF
C722 diff_5019000_4116000# gnd! 95.9fF
C723 diff_4778000_3875000# gnd! 167.8fF
C724 diff_4762000_3821000# gnd! 709.8fF
C725 diff_5114000_4071000# gnd! 498.5fF
C726 diff_5028000_4156000# gnd! 216.4fF
C727 diff_5004000_4150000# gnd! 64.8fF
C728 diff_4715000_3889000# gnd! 160.0fF
C729 diff_5387000_800000# gnd! 1026.2fF
C730 diff_6158000_4260000# gnd! 548.8fF
C731 diff_5164000_4226000# gnd! 334.1fF
C732 diff_5567000_4243000# gnd! 102.0fF
C733 diff_5575000_4252000# gnd! 156.5fF
C734 diff_6145000_4251000# gnd! 408.4fF
C735 diff_5956000_4224000# gnd! 440.6fF
C736 diff_6031000_4330000# gnd! 105.2fF
C737 diff_5603000_4298000# gnd! 157.9fF
C738 diff_5055000_4275000# gnd! 80.6fF
C739 diff_4697000_3226000# gnd! 858.7fF
C740 diff_5091000_4257000# gnd! 235.5fF
C741 diff_5376000_4257000# gnd! 269.9fF
C742 diff_5603000_4344000# gnd! 156.8fF
C743 diff_4241000_2640000# gnd! 1796.0fF
C744 diff_6146000_4381000# gnd! 289.8fF
C745 diff_6187000_3965000# gnd! 404.6fF
C746 diff_4981000_4331000# gnd! 92.5fF
C747 diff_5569000_4409000# gnd! 143.7fF
C748 diff_5389000_4389000# gnd! 158.0fF
C749 diff_5169000_4319000# gnd! 451.8fF
C750 diff_5346000_4399000# gnd! 644.6fF
C751 diff_5056000_4359000# gnd! 185.4fF
C752 diff_5561000_4418000# gnd! 106.5fF
C753 diff_5826000_4381000# gnd! 394.3fF
C754 diff_5949000_4452000# gnd! 282.5fF
C755 diff_6223000_4302000# gnd! 491.3fF
C756 diff_4303000_2657000# gnd! 1329.4fF
C757 diff_5258000_4376000# gnd! 650.5fF
C758 diff_4984000_4430000# gnd! 77.8fF
C759 diff_5389000_4406000# gnd! 1396.0fF
C760 diff_4182000_2528000# gnd! 1162.8fF
C761 diff_4995000_4438000# gnd! 209.3fF
C762 diff_5740000_4460000# gnd! 88.2fF
C763 diff_5980000_4397000# gnd! 417.8fF
C764 diff_5391000_4498000# gnd! 172.9fF
C765 diff_6153000_4534000# gnd! 435.7fF
C766 diff_5397000_4487000# gnd! 137.3fF
C767 diff_5022000_4457000# gnd! 226.4fF
C768 diff_4511000_3502000# gnd! 269.5fF
C769 diff_4495000_3314000# gnd! 923.8fF
C770 diff_4262000_2987000# gnd! 670.9fF
C771 diff_4306000_3185000# gnd! 127.2fF
C772 diff_4225000_2934000# gnd! 449.4fF
C773 diff_4052000_2818000# gnd! 436.4fF
C774 diff_4154000_3010000# gnd! 183.0fF
C775 diff_4297000_3178000# gnd! 363.1fF
C776 diff_4087000_3165000# gnd! 148.8fF
C777 diff_4068000_3124000# gnd! 320.6fF
C778 diff_4095000_3085000# gnd! 123.8fF
C779 diff_3949000_2818000# gnd! 389.6fF
C780 diff_3846000_2818000# gnd! 474.1fF
C781 diff_3904000_3049000# gnd! 86.2fF
C782 diff_4304000_3505000# gnd! 145.9fF
C783 diff_4022000_2818000# gnd! 710.3fF
C784 diff_4462000_3008000# gnd! 786.5fF
C785 diff_4415000_3774000# gnd! 1008.7fF
C786 diff_4419000_3822000# gnd! 147.3fF
C787 diff_4374000_3894000# gnd! 149.2fF
C788 diff_4358000_3758000# gnd! 573.3fF
C789 diff_4458000_3837000# gnd! 427.6fF
C790 diff_4516000_3837000# gnd! 561.1fF
C791 diff_5457000_4544000# gnd! 70.2fF
C792 diff_5229000_4554000# gnd! 275.9fF
C793 diff_5074000_4506000# gnd! 258.0fF
C794 diff_5096000_4554000# gnd! 264.1fF
C795 diff_5711000_4528000# gnd! 306.4fF
C796 diff_6079000_4659000# gnd! 144.8fF
C797 diff_6049000_4641000# gnd! 109.1fF
C798 diff_5337000_4569000# gnd! 286.5fF
C799 diff_5160000_4311000# gnd! 193.3fF
C800 diff_5476000_4643000# gnd! 68.3fF
C801 diff_5127000_4617000# gnd! 300.7fF
C802 diff_4806000_4501000# gnd! 780.7fF
C803 diff_5296000_4530000# gnd! 420.7fF
C804 diff_5127000_4637000# gnd! 81.6fF
C805 diff_5337000_4602000# gnd! 492.6fF
C806 diff_4920000_4669000# gnd! 159.7fF
C807 diff_5991000_4719000# gnd! 133.7fF
C808 diff_6078000_4738000# gnd! 159.2fF
C809 diff_6078000_4787000# gnd! 145.9fF
C810 diff_5641000_4717000# gnd! 330.6fF
C811 diff_4927000_3400000# gnd! 2509.9fF
C812 diff_5489000_4718000# gnd! 151.4fF
C813 diff_5488000_4745000# gnd! 117.9fF
C814 diff_6078000_4836000# gnd! 145.9fF
C815 diff_6029000_4851000# gnd! 113.8fF
C816 diff_5413000_4658000# gnd! 964.1fF
C817 diff_5601000_3945000# gnd! 1652.5fF
C818 diff_6078000_4885000# gnd! 145.9fF
C819 diff_6029000_4890000# gnd! 138.4fF
C820 diff_6029000_4913000# gnd! 169.8fF
C821 diff_5296000_4764000# gnd! 301.5fF
C822 diff_5220000_4035000# gnd! 913.9fF
C823 diff_5098000_4894000# gnd! 1489.8fF
C824 diff_5068000_4962000# gnd! 934.6fF
C825 diff_5039000_4962000# gnd! 786.2fF
C826 diff_5009000_4962000# gnd! 1712.5fF
C827 diff_4751000_4352000# gnd! 512.8fF
C828 diff_4788000_4476000# gnd! 428.1fF
C829 diff_4374000_4012000# gnd! 131.6fF
C830 diff_4265000_3070000# gnd! 1540.5fF
C831 diff_4527000_4142000# gnd! 507.9fF
C832 diff_4028000_3054000# gnd! 678.0fF
C833 diff_4003000_3074000# gnd! 435.3fF
C834 diff_3815000_2818000# gnd! 537.1fF
C835 diff_3917000_3246000# gnd! 88.7fF
C836 diff_3867000_2981000# gnd! 274.7fF
C837 diff_3742000_2818000# gnd! 435.8fF
C838 diff_3867000_3072000# gnd! 119.1fF
C839 diff_3712000_2818000# gnd! 369.2fF
C840 diff_3536000_2818000# gnd! 372.0fF
C841 diff_3639000_2818000# gnd! 586.4fF
C842 diff_4044000_3493000# gnd! 156.7fF
C843 diff_3609000_2818000# gnd! 622.1fF
C844 diff_3819000_3049000# gnd! 479.4fF
C845 diff_3506000_2818000# gnd! 475.1fF
C846 diff_3604000_3007000# gnd! 287.6fF
C847 diff_3579000_3164000# gnd! 81.0fF
C848 diff_3621000_3188000# gnd! 136.6fF
C849 diff_4218000_3818000# gnd! 119.9fF
C850 diff_4187000_3788000# gnd! 91.5fF
C851 diff_4163000_3767000# gnd! 287.4fF
C852 diff_4214000_3933000# gnd! 539.8fF
C853 diff_4169000_3959000# gnd! 90.2fF
C854 diff_4143000_3861000# gnd! 437.4fF
C855 diff_4423000_4318000# gnd! 809.8fF
C856 diff_4524000_4435000# gnd! 102.9fF
C857 diff_4469000_4450000# gnd! 1162.1fF
C858 diff_4694000_4601000# gnd! 728.8fF
C859 diff_4647000_4721000# gnd! 758.6fF
C860 diff_4318000_4212000# gnd! 2026.4fF
C861 diff_4247000_4333000# gnd! 145.9fF
C862 diff_4136000_4237000# gnd! 477.5fF
C863 diff_3791000_3500000# gnd! 190.4fF
C864 diff_3517000_3070000# gnd! 286.4fF
C865 diff_3433000_2818000# gnd! 541.3fF
C866 diff_3487000_3126000# gnd! 143.7fF
C867 diff_3283000_1426000# gnd! 415.8fF
C868 diff_3256000_1459000# gnd! 446.7fF
C869 diff_3321000_2527000# gnd! 872.5fF
C870 diff_3079000_2441000# gnd! 278.9fF
C871 diff_2460000_2101000# gnd! 199.4fF
C872 diff_2407000_2069000# gnd! 181.0fF
C873 diff_2320000_1883000# gnd! 469.3fF
C874 diff_2281000_1866000# gnd! 296.0fF
C875 diff_2184000_1679000# gnd! 268.7fF
C876 diff_2122000_1637000# gnd! 400.7fF
C877 diff_2130000_1666000# gnd! 414.8fF
C878 diff_2137000_1673000# gnd! 231.8fF
C879 diff_2127000_1705000# gnd! 592.3fF
C880 diff_2184000_1871000# gnd! 271.6fF
C881 diff_2137000_1957000# gnd! 222.3fF
C882 diff_2130000_1972000# gnd! 420.5fF
C883 diff_2471000_2112000# gnd! 138.9fF
C884 diff_2683000_2215000# gnd! 521.7fF
C885 diff_2651000_2299000# gnd! 134.2fF
C886 diff_2674000_2207000# gnd! 263.4fF
C887 diff_2532000_2233000# gnd! 222.6fF
C888 diff_2471000_2205000# gnd! 135.8fF
C889 diff_2460000_2210000# gnd! 200.0fF
C890 diff_1997000_1468000# gnd! 450.4fF
C891 diff_1881000_1450000# gnd! 261.5fF
C892 diff_1851000_1456000# gnd! 1625.6fF
C893 diff_1932000_1554000# gnd! 170.8fF
C894 diff_1850000_1535000# gnd! 525.3fF
C895 diff_1997000_1739000# gnd! 459.9fF
C896 diff_2050000_1770000# gnd! 141.7fF
C897 diff_1932000_1705000# gnd! 165.7fF
C898 diff_1851000_1695000# gnd! 503.0fF
C899 diff_1881000_1794000# gnd! 272.4fF
C900 diff_2102000_1984000# gnd! 19.4fF
C901 diff_2050000_1834000# gnd! 137.3fF
C902 diff_2122000_1984000# gnd! 383.5fF
C903 diff_2320000_2130000# gnd! 465.8fF
C904 diff_2127000_1922000# gnd! 610.7fF
C905 diff_2281000_2086000# gnd! 288.6fF
C906 diff_2406000_2323000# gnd! 184.1fF
C907 diff_2320000_2261000# gnd! 473.9fF
C908 diff_2102000_2014000# gnd! 20.3fF
C909 diff_2184000_2056000# gnd! 267.6fF
C910 diff_2122000_2014000# gnd! 402.3fF
C911 diff_2130000_2043000# gnd! 415.1fF
C912 diff_2137000_2050000# gnd! 231.4fF
C913 diff_2127000_2082000# gnd! 515.5fF
C914 diff_2281000_2195000# gnd! 293.2fF
C915 diff_3171000_2725000# gnd! 1500.5fF
C916 diff_3120000_2492000# gnd! 1463.2fF
C917 diff_3043000_2723000# gnd! 1029.9fF
C918 diff_2184000_2248000# gnd! 269.4fF
C919 diff_2137000_2334000# gnd! 223.8fF
C920 diff_2130000_2350000# gnd! 416.1fF
C921 diff_1997000_1845000# gnd! 449.4fF
C922 diff_1881000_1826000# gnd! 266.5fF
C923 diff_1932000_1931000# gnd! 171.9fF
C924 diff_2050000_2147000# gnd! 138.3fF
C925 diff_1997000_2116000# gnd! 458.0fF
C926 diff_1850000_1913000# gnd! 523.2fF
C927 diff_1932000_2082000# gnd! 168.3fF
C928 diff_1850000_2072000# gnd! 510.6fF
C929 diff_1881000_2171000# gnd! 271.7fF
C930 diff_2102000_2360000# gnd! 21.2fF
C931 diff_2050000_2211000# gnd! 143.0fF
C932 diff_2122000_2360000# gnd! 387.7fF
C933 diff_1997000_2222000# gnd! 449.2fF
C934 diff_1881000_2203000# gnd! 270.6fF
C935 diff_1932000_2308000# gnd! 175.6fF
C936 diff_1850000_2290000# gnd! 510.6fF
C937 diff_2996000_2725000# gnd! 1450.3fF
C938 diff_2939000_824000# gnd! 1157.6fF
C939 diff_2893000_2725000# gnd! 1568.0fF
C940 diff_2843000_1950000# gnd! 1469.5fF
C941 diff_2775000_765000# gnd! 1542.0fF
C942 diff_2713000_822000# gnd! 1483.0fF
C943 diff_2641000_934000# gnd! 1389.5fF
C944 diff_2638000_2492000# gnd! 1481.5fF
C945 diff_2583000_2725000# gnd! 1530.4fF
C946 diff_2534000_2492000# gnd! 1526.7fF
C947 diff_3168000_2777000# gnd! 231.8fF
C948 diff_3115000_2777000# gnd! 229.4fF
C949 diff_3047000_2783000# gnd! 280.5fF
C950 diff_2994000_2777000# gnd! 225.1fF
C951 diff_2941000_2777000# gnd! 223.4fF
C952 diff_2891000_2777000# gnd! 220.4fF
C953 diff_2838000_2777000# gnd! 235.0fF
C954 diff_2788000_2777000# gnd! 229.0fF
C955 diff_2735000_2777000# gnd! 234.2fF
C956 diff_2684000_2777000# gnd! 234.4fF
C957 diff_2632000_2777000# gnd! 228.0fF
C958 diff_2581000_2777000# gnd! 229.6fF
C959 diff_2529000_2777000# gnd! 229.4fF
C960 diff_2448000_2717000# gnd! 1570.6fF
C961 diff_3254000_2509000# gnd! 1030.9fF
C962 diff_3355000_3022000# gnd! 155.2fF
C963 diff_3365000_3033000# gnd! 358.9fF
C964 diff_3517000_3179000# gnd! 83.1fF
C965 diff_3551000_3277000# gnd! 826.3fF
C966 diff_2838000_2818000# gnd! 653.5fF
C967 diff_3187000_3099000# gnd! 228.0fF
C968 diff_3282000_3144000# gnd! 156.8fF
C969 diff_3231000_3142000# gnd! 145.9fF
C970 diff_3014000_2818000# gnd! 1354.0fF
C971 diff_3050000_2818000# gnd! 405.3fF
C972 diff_2941000_2818000# gnd! 389.8fF
C973 diff_3188000_2818000# gnd! 994.5fF
C974 diff_3944000_3772000# gnd! 121.8fF
C975 diff_3939000_3886000# gnd! 144.8fF
C976 diff_4066000_4315000# gnd! 131.7fF
C977 diff_4467000_4516000# gnd! 218.2fF
C978 diff_4920000_4772000# gnd! 535.3fF
C979 diff_4902000_4754000# gnd! 340.9fF
C980 diff_4883000_4962000# gnd! 817.1fF
C981 diff_4843000_4668000# gnd! 201.6fF
C982 diff_4824000_4962000# gnd! 135.1fF
C983 diff_4770000_4458000# gnd! 81.3fF
C984 diff_4428000_3813000# gnd! 446.8fF
C985 diff_4735000_4962000# gnd! 169.3fF
C986 diff_4382000_4593000# gnd! 380.0fF
C987 diff_4125000_2818000# gnd! 1101.6fF
C988 diff_4175000_4495000# gnd! 458.7fF
C989 diff_4126000_4460000# gnd! 401.7fF
C990 diff_3909000_4369000# gnd! 500.2fF
C991 diff_3702000_3518000# gnd! 88.7fF
C992 diff_3645000_3521000# gnd! 162.4fF
C993 diff_3444000_3167000# gnd! 793.2fF
C994 diff_3569000_3530000# gnd! 1342.1fF
C995 diff_3981000_4517000# gnd! 948.8fF
C996 diff_4020000_4533000# gnd! 296.8fF
C997 diff_3668000_3852000# gnd! 169.1fF
C998 diff_3122000_3080000# gnd! 118.7fF
C999 diff_3061000_3052000# gnd! 332.8fF
C1000 diff_3072000_3193000# gnd! 80.7fF
C1001 diff_3024000_3075000# gnd! 141.1fF
C1002 diff_2978000_3080000# gnd! 189.0fF
C1003 diff_2911000_2818000# gnd! 464.5fF
C1004 diff_2907000_3149000# gnd! 268.5fF
C1005 diff_2874000_3145000# gnd! 78.5fF
C1006 diff_2922000_3078000# gnd! 78.7fF
C1007 diff_2808000_2818000# gnd! 450.3fF
C1008 diff_2819000_3094000# gnd! 133.6fF
C1009 diff_2735000_2818000# gnd! 390.3fF
C1010 diff_2744000_3026000# gnd! 92.8fF
C1011 diff_3619000_3826000# gnd! 295.5fF
C1012 diff_3532000_3485000# gnd! 494.1fF
C1013 diff_3677000_3847000# gnd! 106.9fF
C1014 diff_3623000_3886000# gnd! 94.3fF
C1015 diff_3448000_3517000# gnd! 607.6fF
C1016 diff_3583000_4085000# gnd! 89.3fF
C1017 diff_3666000_4069000# gnd! 932.2fF
C1018 diff_3666000_4149000# gnd! 160.4fF
C1019 diff_3535000_3825000# gnd! 464.4fF
C1020 diff_3658000_4142000# gnd! 275.4fF
C1021 diff_3887000_4604000# gnd! 240.2fF
C1022 diff_3607000_4424000# gnd! 443.3fF
C1023 diff_3664000_4488000# gnd! 594.4fF
C1024 diff_3113000_3386000# gnd! 351.1fF
C1025 diff_2988000_3091000# gnd! 458.2fF
C1026 diff_3413000_3852000# gnd! 225.1fF
C1027 diff_3212000_3556000# gnd! 272.9fF
C1028 diff_2986000_3296000# gnd! 415.1fF
C1029 diff_2127000_2299000# gnd! 826.0fF
C1030 diff_2288000_2488000# gnd! 422.6fF
C1031 diff_2304000_1746000# gnd! 2125.3fF
C1032 diff_1791000_798000# gnd! 1596.3fF
C1033 diff_1774000_760000# gnd! 1815.0fF
C1034 diff_1386000_841000# gnd! 750.9fF
C1035 diff_1437000_884000# gnd! 30.4fF
C1036 diff_1556000_944000# gnd! 131.0fF
C1037 diff_1583000_1024000# gnd! 514.4fF
C1038 diff_1576000_1014000# gnd! 256.6fF
C1039 diff_1583000_1098000# gnd! 504.6fF
C1040 diff_1477000_942000# gnd! 485.9fF
C1041 diff_1460000_884000# gnd! 144.4fF
C1042 diff_1556000_1173000# gnd! 137.2fF
C1043 diff_1576000_1089000# gnd! 254.8fF
C1044 diff_1477000_1091000# gnd! 476.8fF
C1045 diff_1390000_920000# gnd! 162.0fF
C1046 diff_1345000_885000# gnd! 336.4fF
C1047 diff_1305000_907000# gnd! 270.1fF
C1048 diff_1390000_1180000# gnd! 163.2fF
C1049 diff_792000_356000# gnd! 2190.9fF
C1050 diff_906000_615000# gnd! 255.9fF
C1051 diff_123000_488000# gnd! 2288.8fF
C1052 diff_582000_709000# gnd! 264.2fF
C1053 diff_1460000_1230000# gnd! 148.9fF
C1054 diff_1437000_1230000# gnd! 31.8fF
C1055 diff_1305000_1208000# gnd! 269.6fF
C1056 diff_1238000_975000# gnd! 493.0fF
C1057 diff_1188000_1219000# gnd! 279.5fF
C1058 diff_1345000_1229000# gnd! 340.4fF
C1059 diff_1437000_1261000# gnd! 31.8fF
C1060 diff_1557000_1321000# gnd! 130.2fF
C1061 diff_1583000_1401000# gnd! 512.3fF
C1062 diff_1576000_1391000# gnd! 253.2fF
C1063 diff_1583000_1475000# gnd! 506.7fF
C1064 diff_1477000_1320000# gnd! 485.7fF
C1065 diff_1460000_1261000# gnd! 147.6fF
C1066 diff_1557000_1550000# gnd! 133.7fF
C1067 diff_1576000_1466000# gnd! 251.7fF
C1068 diff_1757000_739000# gnd! 1674.0fF
C1069 diff_1477000_1468000# gnd! 477.0fF
C1070 diff_1390000_1297000# gnd! 163.1fF
C1071 diff_1345000_1262000# gnd! 340.8fF
C1072 diff_1305000_1284000# gnd! 269.6fF
C1073 diff_1390000_1558000# gnd! 161.7fF
C1074 diff_1460000_1607000# gnd! 149.4fF
C1075 diff_1437000_1607000# gnd! 31.8fF
C1076 diff_1305000_1585000# gnd! 271.0fF
C1077 diff_1236000_1245000# gnd! 669.6fF
C1078 diff_1085000_969000# gnd! 184.7fF
C1079 diff_1064000_933000# gnd! 472.6fF
C1080 diff_132000_496000# gnd! 3747.3fF
C1081 diff_123000_700000# gnd! 2282.4fF
C1082 diff_1010000_1054000# gnd! 189.6fF
C1083 diff_970000_884000# gnd! 938.3fF
C1084 diff_889000_963000# gnd! 270.9fF
C1085 diff_914000_1003000# gnd! 270.2fF
C1086 diff_1085000_1080000# gnd! 183.8fF
C1087 diff_1010000_1073000# gnd! 198.1fF
C1088 diff_856000_890000# gnd! 230.2fF
C1089 diff_848000_885000# gnd! 1233.7fF
C1090 diff_582000_964000# gnd! 270.2fF
C1091 diff_1064000_1080000# gnd! 527.0fF
C1092 diff_889000_1153000# gnd! 273.6fF
C1093 diff_709000_308000# gnd! 1226.8fF
C1094 diff_914000_1079000# gnd! 265.9fF
C1095 diff_1188000_1277000# gnd! 315.0fF
C1096 diff_1236000_1424000# gnd! 647.1fF
C1097 diff_1085000_1346000# gnd! 184.8fF
C1098 diff_1063000_1310000# gnd! 547.0fF
C1099 diff_856000_1218000# gnd! 225.5fF
C1100 diff_817000_1211000# gnd! 2991.1fF
C1101 diff_848000_1211000# gnd! 1242.5fF
C1102 diff_123000_866000# gnd! 2268.9fF
C1103 diff_132000_874000# gnd! 3785.1fF
C1104 diff_123000_1087000# gnd! 2289.6fF
C1105 diff_1010000_1431000# gnd! 189.6fF
C1106 diff_752000_680000# gnd! 1039.3fF
C1107 diff_889000_1340000# gnd! 271.9fF
C1108 diff_914000_1380000# gnd! 265.9fF
C1109 diff_1345000_1606000# gnd! 343.1fF
C1110 diff_1437000_1638000# gnd! 31.8fF
C1111 diff_1556000_1698000# gnd! 131.9fF
C1112 diff_1583000_1778000# gnd! 506.4fF
C1113 diff_1576000_1768000# gnd! 254.9fF
C1114 diff_1399000_598000# gnd! 2021.4fF
C1115 diff_1583000_1852000# gnd! 504.0fF
C1116 diff_1477000_1697000# gnd! 496.6fF
C1117 diff_1460000_1638000# gnd! 146.8fF
C1118 diff_1556000_1927000# gnd! 135.8fF
C1119 diff_1576000_1843000# gnd! 249.8fF
C1120 diff_1477000_1846000# gnd! 485.4fF
C1121 diff_1196000_1522000# gnd! 250.3fF
C1122 diff_1085000_1457000# gnd! 183.9fF
C1123 diff_817000_1286000# gnd! 3615.2fF
C1124 diff_1010000_1450000# gnd! 200.8fF
C1125 diff_856000_1267000# gnd! 228.0fF
C1126 diff_848000_1262000# gnd! 1240.9fF
C1127 diff_123000_1243000# gnd! 2306.2fF
C1128 diff_1390000_1674000# gnd! 163.0fF
C1129 diff_1345000_1639000# gnd! 342.4fF
C1130 diff_1305000_1661000# gnd! 269.6fF
C1131 diff_1202000_1633000# gnd! 725.4fF
C1132 diff_1390000_1935000# gnd! 161.7fF
C1133 diff_1460000_1984000# gnd! 150.7fF
C1134 diff_1437000_1984000# gnd! 31.8fF
C1135 diff_1305000_1962000# gnd! 270.4fF
C1136 diff_1265000_1694000# gnd! 631.7fF
C1137 diff_1345000_1983000# gnd! 340.2fF
C1138 diff_1437000_2015000# gnd! 31.8fF
C1139 diff_1556000_2076000# gnd! 131.8fF
C1140 diff_1583000_2155000# gnd! 498.4fF
C1141 diff_1576000_2146000# gnd! 254.5fF
C1142 diff_1583000_2229000# gnd! 498.5fF
C1143 diff_1477000_2074000# gnd! 485.9fF
C1144 diff_1460000_2015000# gnd! 147.4fF
C1145 diff_1556000_2304000# gnd! 134.6fF
C1146 diff_1576000_2220000# gnd! 254.0fF
C1147 diff_1477000_2222000# gnd! 481.8fF
C1148 diff_1189000_1979000# gnd! 329.6fF
C1149 diff_1390000_2052000# gnd! 162.0fF
C1150 diff_1345000_2016000# gnd! 339.6fF
C1151 diff_1305000_2038000# gnd! 268.5fF
C1152 diff_1245000_1992000# gnd! 736.5fF
C1153 diff_1189000_2023000# gnd! 331.7fF
C1154 diff_1390000_2312000# gnd! 163.0fF
C1155 diff_1460000_2361000# gnd! 149.8fF
C1156 diff_1437000_2361000# gnd! 31.8fF
C1157 diff_1305000_2339000# gnd! 269.9fF
C1158 diff_1245000_2015000# gnd! 723.5fF
C1159 diff_1345000_2360000# gnd! 342.2fF
C1160 diff_2208000_2717000# gnd! 230.8fF
C1161 diff_1858000_1019000# gnd! 1618.5fF
C1162 diff_1837000_1364000# gnd! 1546.8fF
C1163 diff_2113000_2778000# gnd! 237.8fF
C1164 diff_2060000_2777000# gnd! 223.9fF
C1165 diff_2602000_2818000# gnd! 372.5fF
C1166 diff_2632000_2818000# gnd! 581.5fF
C1167 diff_2678000_3055000# gnd! 371.8fF
C1168 diff_2962000_3296000# gnd! 164.2fF
C1169 diff_3348000_3929000# gnd! 174.8fF
C1170 diff_3325000_3886000# gnd! 315.0fF
C1171 diff_3339000_4042000# gnd! 103.4fF
C1172 diff_3272000_3283000# gnd! 535.3fF
C1173 diff_3535000_4387000# gnd! 198.3fF
C1174 diff_3401000_3461000# gnd! 788.6fF
C1175 diff_3494000_4370000# gnd! 211.0fF
C1176 diff_3399000_4294000# gnd! 228.3fF
C1177 diff_3380000_4294000# gnd! 252.2fF
C1178 diff_3408000_4288000# gnd! 3608.6fF
C1179 diff_2790000_3479000# gnd! 99.8fF
C1180 diff_2810000_3352000# gnd! 414.9fF
C1181 diff_3017000_3539000# gnd! 191.7fF
C1182 diff_2573000_3039000# gnd! 102.7fF
C1183 diff_2561000_3213000# gnd! 531.0fF
C1184 diff_2521000_3105000# gnd! 88.8fF
C1185 diff_1729000_1868000# gnd! 667.5fF
C1186 diff_1729000_2091000# gnd! 516.7fF
C1187 diff_1931000_2739000# gnd! 332.9fF
C1188 diff_1728000_2245000# gnd! 505.3fF
C1189 diff_1874000_2769000# gnd! 232.2fF
C1190 diff_1189000_2359000# gnd! 321.0fF
C1191 diff_1063000_1457000# gnd! 538.3fF
C1192 diff_889000_1530000# gnd! 271.8fF
C1193 diff_719000_1030000# gnd! 992.6fF
C1194 diff_914000_1456000# gnd! 264.5fF
C1195 diff_1085000_1723000# gnd! 186.1fF
C1196 diff_1064000_1687000# gnd! 581.8fF
C1197 diff_856000_1595000# gnd! 228.6fF
C1198 diff_817000_1588000# gnd! 3392.7fF
C1199 diff_848000_1588000# gnd! 1370.6fF
C1200 diff_582000_1463000# gnd! 260.0fF
C1201 diff_132000_1251000# gnd! 3788.3fF
C1202 diff_123000_1453000# gnd! 2295.9fF
C1203 diff_1010000_1808000# gnd! 189.6fF
C1204 diff_719000_1426000# gnd! 964.1fF
C1205 diff_888000_1717000# gnd! 269.5fF
C1206 diff_914000_1757000# gnd! 262.4fF
C1207 diff_817000_1663000# gnd! 3446.2fF
C1208 diff_1085000_1834000# gnd! 183.7fF
C1209 diff_1010000_1827000# gnd! 200.8fF
C1210 diff_856000_1645000# gnd! 225.2fF
C1211 diff_848000_1639000# gnd! 1246.5fF
C1212 diff_582000_1718000# gnd! 270.1fF
C1213 diff_1064000_1834000# gnd! 606.9fF
C1214 diff_889000_1907000# gnd! 269.4fF
C1215 diff_719000_1784000# gnd! 881.3fF
C1216 diff_914000_1833000# gnd! 264.5fF
C1217 diff_1085000_2099000# gnd! 187.4fF
C1218 diff_1064000_2064000# gnd! 609.7fF
C1219 diff_856000_1972000# gnd! 230.7fF
C1220 diff_817000_1965000# gnd! 3416.1fF
C1221 diff_848000_1965000# gnd! 1357.3fF
C1222 diff_1010000_2185000# gnd! 189.7fF
C1223 diff_889000_2094000# gnd! 266.1fF
C1224 diff_914000_2134000# gnd! 262.4fF
C1225 diff_1085000_2211000# gnd! 184.6fF
C1226 diff_817000_2040000# gnd! 3727.5fF
C1227 diff_1010000_2204000# gnd! 196.5fF
C1228 diff_856000_2022000# gnd! 227.0fF
C1229 diff_848000_2016000# gnd! 1251.3fF
C1230 diff_123000_1620000# gnd! 2271.5fF
C1231 diff_132000_1628000# gnd! 3795.4fF
C1232 diff_123000_1841000# gnd! 2313.1fF
C1233 diff_719000_2180000# gnd! 866.3fF
C1234 diff_123000_1997000# gnd! 2291.8fF
C1235 diff_1064000_2211000# gnd! 606.1fF
C1236 diff_889000_2284000# gnd! 270.8fF
C1237 diff_914000_2210000# gnd! 262.3fF
C1238 diff_1094000_1020000# gnd! 2006.0fF
C1239 diff_1037000_877000# gnd! 2036.4fF
C1240 diff_856000_2349000# gnd! 226.1fF
C1241 diff_817000_2342000# gnd! 3158.0fF
C1242 diff_582000_2217000# gnd! 260.0fF
C1243 diff_848000_2342000# gnd! 1367.9fF
C1244 diff_1696000_986000# gnd! 1519.2fF
C1245 diff_1643000_833000# gnd! 1475.2fF
C1246 diff_1816000_2509000# gnd! 246.1fF
C1247 diff_1776000_2770000# gnd! 250.8fF
C1248 diff_1547000_932000# gnd! 2438.0fF
C1249 diff_1487000_841000# gnd! 2892.4fF
C1250 diff_1712000_2778000# gnd! 217.9fF
C1251 diff_1659000_2777000# gnd! 236.1fF
C1252 diff_1252000_2261000# gnd! 1037.0fF
C1253 diff_1237000_1921000# gnd! 2348.3fF
C1254 diff_1176000_1643000# gnd! 1827.9fF
C1255 diff_1393000_2558000# gnd! 502.1fF
C1256 diff_132000_2005000# gnd! 3407.9fF
C1257 diff_123000_2207000# gnd! 2286.9fF
C1258 diff_1281000_2492000# gnd! 296.0fF
C1259 diff_1150000_1007000# gnd! 2665.7fF
C1260 diff_1318000_2487000# gnd! 311.1fF
C1261 diff_1276000_2574000# gnd! 899.4fF
C1262 diff_1610000_2779000# gnd! 232.7fF
C1263 diff_1554000_2586000# gnd! 254.2fF
C1264 diff_2400000_2876000# gnd! 508.1fF
C1265 diff_2464000_2895000# gnd! 435.6fF
C1266 diff_2420000_3102000# gnd! 95.2fF
C1267 diff_2390000_3201000# gnd! 101.6fF
C1268 diff_2356000_3007000# gnd! 370.3fF
C1269 diff_2182000_3046000# gnd! 528.3fF
C1270 diff_2248000_3126000# gnd! 195.1fF
C1271 diff_2293000_3174000# gnd! 442.5fF
C1272 diff_2066000_3013000# gnd! 457.3fF
C1273 diff_2134000_3060000# gnd! 642.7fF
C1274 diff_2110000_2945000# gnd! 554.8fF
C1275 diff_2082000_3201000# gnd! 134.3fF
C1276 diff_1963000_2987000# gnd! 383.9fF
C1277 diff_1998000_3198000# gnd! 98.6fF
C1278 diff_2004000_3055000# gnd! 501.2fF
C1279 diff_1935000_3038000# gnd! 491.7fF
C1280 diff_817000_909000# gnd! 3582.8fF
C1281 diff_1808000_2942000# gnd! 194.3fF
C1282 diff_1751000_2974000# gnd! 442.8fF
C1283 diff_1840000_3083000# gnd! 341.1fF
C1284 diff_1826000_2942000# gnd! 538.1fF
C1285 diff_1962000_3117000# gnd! 185.1fF
C1286 diff_2351000_3074000# gnd! 2826.2fF
C1287 diff_3048000_3539000# gnd! 247.6fF
C1288 diff_2633000_3304000# gnd! 450.4fF
C1289 diff_2651000_3482000# gnd! 157.2fF
C1290 diff_2598000_3304000# gnd! 217.2fF
C1291 diff_2660000_3493000# gnd! 432.8fF
C1292 diff_2772000_3402000# gnd! 909.5fF
C1293 diff_3005000_3816000# gnd! 194.9fF
C1294 diff_3032000_3774000# gnd! 118.3fF
C1295 diff_1698000_2848000# gnd! 1129.7fF
C1296 diff_1817000_2934000# gnd! 722.9fF
C1297 diff_1733000_2883000# gnd! 856.0fF
C1298 diff_1438000_786000# gnd! 3152.0fF
C1299 diff_1586000_2912000# gnd! 138.3fF
C1300 diff_1259000_2736000# gnd! 185.2fF
C1301 diff_1259000_2792000# gnd! 559.9fF
C1302 diff_901000_991000# gnd! 1615.9fF
C1303 diff_877000_1128000# gnd! 2074.1fF
C1304 diff_1157000_2480000# gnd! 292.4fF
C1305 diff_955000_2507000# gnd! 271.9fF
C1306 diff_1716000_2866000# gnd! 763.7fF
C1307 diff_2219000_3479000# gnd! 258.7fF
C1308 diff_2882000_3711000# gnd! 212.1fF
C1309 diff_3024000_3904000# gnd! 89.3fF
C1310 diff_3009000_3950000# gnd! 151.8fF
C1311 diff_2821000_3543000# gnd! 584.8fF
C1312 diff_2909000_3804000# gnd! 391.1fF
C1313 diff_2904000_3862000# gnd! 265.9fF
C1314 diff_2868000_3892000# gnd! 151.3fF
C1315 diff_2965000_3936000# gnd! 107.3fF
C1316 diff_2697000_3827000# gnd! 137.3fF
C1317 diff_2270000_3390000# gnd! 622.2fF
C1318 diff_582000_2472000# gnd! 270.6fF
C1319 diff_680000_1019000# gnd! 1900.2fF
C1320 diff_719000_2538000# gnd! 1039.0fF
C1321 diff_123000_2374000# gnd! 2266.4fF
C1322 diff_132000_2382000# gnd! 3850.9fF
C1323 diff_123000_2595000# gnd! 2338.0fF
C1324 diff_553000_1211000# gnd! 9712.0fF
C1325 diff_938000_2548000# gnd! 637.2fF
C1326 diff_1405000_2969000# gnd! 149.1fF
C1327 diff_1459000_2943000# gnd! 385.6fF
C1328 diff_1482000_3103000# gnd! 109.1fF
C1329 diff_1411000_3066000# gnd! 102.4fF
C1330 diff_1334000_2958000# gnd! 699.4fF
C1331 diff_1340000_3008000# gnd! 606.5fF
C1332 diff_1604000_3123000# gnd! 1655.7fF
C1333 diff_1328000_3051000# gnd! 453.9fF
C1334 diff_1251000_3051000# gnd! 100.8fF
C1335 diff_2340000_3697000# gnd! 175.9fF
C1336 diff_2912000_3918000# gnd! 150.8fF
C1337 diff_2938000_3467000# gnd! 760.4fF
C1338 diff_2853000_4056000# gnd! 96.4fF
C1339 diff_2799000_4040000# gnd! 469.6fF
C1340 diff_3667000_4701000# gnd! 1056.7fF
C1341 diff_3754000_4644000# gnd! 286.5fF
C1342 diff_3700000_4748000# gnd! 855.0fF
C1343 diff_3539000_4683000# gnd! 106.4fF
C1344 diff_3272000_4383000# gnd! 189.7fF
C1345 diff_3430000_4645000# gnd! 169.5fF
C1346 diff_3421000_4638000# gnd! 375.7fF
C1347 diff_3488000_4662000# gnd! 805.1fF
C1348 diff_3359000_4501000# gnd! 1606.6fF
C1349 diff_3184000_4336000# gnd! 455.1fF
C1350 diff_3033000_4154000# gnd! 802.1fF
C1351 diff_3014000_3475000# gnd! 1100.0fF
C1352 diff_3012000_4154000# gnd! 394.5fF
C1353 diff_2559000_3889000# gnd! 929.0fF
C1354 diff_2895000_4350000# gnd! 126.5fF
C1355 diff_2913000_4304000# gnd! 334.1fF
C1356 diff_3062000_4310000# gnd! 401.6fF
C1357 diff_2877000_4437000# gnd! 93.0fF
C1358 diff_3009000_4523000# gnd! 648.7fF
C1359 diff_2971000_4656000# gnd! 856.6fF
C1360 diff_2931000_4557000# gnd! 1063.1fF
C1361 diff_2915000_4682000# gnd! 87.6fF
C1362 diff_2878000_4622000# gnd! 623.6fF
C1363 diff_2906000_4658000# gnd! 374.6fF
C1364 diff_2860000_4570000# gnd! 663.0fF
C1365 diff_2509000_3809000# gnd! 433.4fF
C1366 diff_2490000_3879000# gnd! 115.5fF
C1367 diff_2471000_3862000# gnd! 95.0fF
C1368 diff_2687000_4368000# gnd! 147.2fF
C1369 diff_2642000_3475000# gnd! 815.6fF
C1370 diff_2647000_4397000# gnd! 159.2fF
C1371 diff_2182000_3681000# gnd! 562.6fF
C1372 diff_2174000_3677000# gnd! 414.8fF
C1373 diff_2028000_3555000# gnd! 381.0fF
C1374 diff_1556000_2817000# gnd! 635.3fF
C1375 diff_1502000_2925000# gnd! 1665.6fF
C1376 diff_1276000_3249000# gnd! 73.6fF
C1377 diff_1188000_3107000# gnd! 711.7fF
C1378 diff_1281000_3071000# gnd! 591.2fF
C1379 diff_1148000_3109000# gnd! 114.0fF
C1380 diff_1028000_3008000# gnd! 446.6fF
C1381 diff_1048000_3119000# gnd! 1212.2fF
C1382 diff_967000_2989000# gnd! 659.6fF
C1383 diff_962000_3082000# gnd! 159.2fF
C1384 diff_917000_3186000# gnd! 98.6fF
C1385 diff_875000_3125000# gnd! 105.0fF
C1386 diff_912000_3048000# gnd! 360.6fF
C1387 diff_1979000_3617000# gnd! 254.9fF
C1388 diff_1659000_2818000# gnd! 949.8fF
C1389 diff_1834000_3561000# gnd! 144.8fF
C1390 diff_946000_3225000# gnd! 114.5fF
C1391 diff_2073000_3806000# gnd! 250.6fF
C1392 diff_2050000_3807000# gnd! 433.6fF
C1393 diff_2324000_3768000# gnd! 339.3fF
C1394 diff_2337000_4018000# gnd! 89.0fF
C1395 diff_2256000_3932000# gnd! 78.0fF
C1396 diff_2568000_4388000# gnd! 145.9fF
C1397 diff_2154000_3995000# gnd! 558.9fF
C1398 diff_2222000_4172000# gnd! 414.1fF
C1399 diff_2129000_4009000# gnd! 918.4fF
C1400 diff_2111000_3992000# gnd! 242.0fF
C1401 diff_2093000_3973000# gnd! 247.8fF
C1402 diff_2120000_4001000# gnd! 1526.2fF
C1403 diff_1944000_3756000# gnd! 160.2fF
C1404 diff_1465000_3204000# gnd! 573.4fF
C1405 diff_1993000_3921000# gnd! 217.4fF
C1406 diff_1976000_3921000# gnd! 217.4fF
C1407 diff_2198000_3000000# gnd! 1258.1fF
C1408 diff_2566000_3500000# gnd! 1094.4fF
C1409 diff_2405000_4387000# gnd! 493.9fF
C1410 diff_2570000_3912000# gnd! 1450.7fF
C1411 diff_2173000_3038000# gnd! 1431.9fF
C1412 diff_1953000_3750000# gnd! 550.4fF
C1413 diff_1902000_3917000# gnd! 159.2fF
C1414 diff_2194000_4240000# gnd! 178.3fF
C1415 diff_2187000_4495000# gnd! 921.1fF
C1416 diff_2063000_4304000# gnd! 696.6fF
C1417 diff_2060000_4467000# gnd! 96.4fF
C1418 diff_1475000_3480000# gnd! 88.3fF
C1419 diff_1622000_3414000# gnd! 204.8fF
C1420 diff_1539000_3467000# gnd! 192.2fF
C1421 diff_1561000_3639000# gnd! 264.1fF
C1422 diff_1459000_3632000# gnd! 89.3fF
C1423 diff_1646000_3414000# gnd! 723.9fF
C1424 diff_1713000_3885000# gnd! 291.3fF
C1425 diff_1741000_4000000# gnd! 84.3fF
C1426 diff_1589000_4012000# gnd! 105.5fF
C1427 diff_2005000_4584000# gnd! 218.1fF
C1428 diff_2135000_4721000# gnd! 648.4fF
C1429 diff_1966000_4584000# gnd! 529.1fF
C1430 diff_1276000_3285000# gnd! 1980.0fF
C1431 diff_743000_2974000# gnd! 1187.6fF
C1432 diff_1097000_3119000# gnd! 1634.7fF
C1433 diff_823000_3289000# gnd! 207.7fF
C1434 diff_1272000_3500000# gnd! 70.5fF
C1435 diff_1339000_3691000# gnd! 134.1fF
C1436 diff_1508000_3890000# gnd! 107.5fF
C1437 diff_1516000_3900000# gnd! 690.7fF
C1438 diff_1691000_4259000# gnd! 293.0fF
C1439 diff_1483000_3488000# gnd! 981.9fF
C1440 diff_1436000_3778000# gnd! 343.4fF
C1441 diff_1419000_3778000# gnd! 174.5fF
C1442 diff_1406000_3519000# gnd! 346.8fF
C1443 diff_1477000_3932000# gnd! 526.5fF
C1444 diff_640000_3020000# gnd! 89.6fF
C1445 diff_669000_2930000# gnd! 638.0fF
C1446 diff_687000_3101000# gnd! 817.3fF
C1447 diff_1740000_4513000# gnd! 247.4fF
C1448 diff_1549000_4377000# gnd! 115.5fF
C1449 diff_1595000_4502000# gnd! 367.1fF
C1450 diff_1523000_4349000# gnd! 103.8fF
C1451 diff_557000_2988000# gnd! 409.5fF
C1452 diff_534000_2989000# gnd! 136.2fF
C1453 diff_83000_3131000# gnd! 219.6fF
C1454 diff_83000_3148000# gnd! 285.1fF
C1455 diff_102000_3167000# gnd! 422.1fF
C1456 diff_111000_3254000# gnd! 83.1fF
C1457 diff_90000_3265000# gnd! 293.1fF
C1458 diff_1237000_3461000# gnd! 565.4fF
C1459 diff_906000_3226000# gnd! 2005.2fF
C1460 diff_1692000_4497000# gnd! 134.5fF
C1461 diff_1541000_4610000# gnd! 456.6fF
C1462 diff_1674000_4606000# gnd! 566.6fF
C1463 diff_860000_2987000# gnd! 1553.4fF
C1464 diff_128000_3343000# gnd! 246.7fF
C1465 diff_206000_3372000# gnd! 82.4fF
C1466 diff_111000_3358000# gnd! 523.5fF
C1467 diff_906000_3511000# gnd! 165.5fF
C1468 diff_946000_3261000# gnd! 1428.9fF
C1469 diff_1142000_3814000# gnd! 160.4fF
C1470 diff_1152000_3809000# gnd! 125.7fF
C1471 diff_1134000_3807000# gnd! 117.9fF
C1472 diff_1048000_3792000# gnd! 159.2fF
C1473 diff_784000_3633000# gnd! 1203.5fF
C1474 diff_731000_3544000# gnd! 136.6fF
C1475 diff_1079000_3958000# gnd! 86.8fF
C1476 diff_1029000_3949000# gnd! 117.7fF
C1477 diff_987000_3874000# gnd! 210.0fF
C1478 diff_1055000_3959000# gnd! 103.7fF
C1479 diff_856000_3301000# gnd! 911.5fF
C1480 diff_787000_3667000# gnd! 76.2fF
C1481 diff_111000_3412000# gnd! 107.8fF
C1482 diff_104000_3450000# gnd! 471.3fF
C1483 diff_104000_3496000# gnd! 99.4fF
C1484 diff_88000_3357000# gnd! 232.3fF
C1485 diff_124000_3549000# gnd! 104.0fF
C1486 diff_101000_3535000# gnd! 499.8fF
C1487 diff_929000_3956000# gnd! 85.9fF
C1488 diff_997000_3891000# gnd! 101.6fF
C1489 diff_1180000_3099000# gnd! 680.5fF
C1490 diff_1448000_4598000# gnd! 362.9fF
C1491 diff_1000000_2990000# gnd! 2097.2fF
C1492 diff_1262000_4413000# gnd! 132.6fF
C1493 diff_1195000_4346000# gnd! 165.1fF
C1494 diff_1149000_4301000# gnd! 206.7fF
C1495 diff_1200000_4480000# gnd! 104.8fF
C1496 diff_1235000_4461000# gnd! 834.1fF
C1497 diff_3227000_4780000# gnd! 1363.3fF
C1498 diff_991000_3076000# gnd! 1549.9fF
C1499 diff_807000_3040000# gnd! 991.3fF
C1500 diff_94000_3158000# gnd! 1915.2fF
C1501 diff_4617000_4962000# gnd! 200.1fF
C1502 diff_4587000_4962000# gnd! 180.1fF
C1503 diff_4559000_4962000# gnd! 183.8fF
C1504 diff_4529000_4962000# gnd! 679.2fF
C1505 diff_4499000_4962000# gnd! 641.1fF
C1506 diff_4469000_4962000# gnd! 501.1fF
C1507 diff_4319000_4839000# gnd! 923.2fF
C1508 diff_4411000_4962000# gnd! 318.9fF
C1509 diff_4381000_4962000# gnd! 252.3fF
C1510 diff_4351000_4962000# gnd! 430.8fF
C1511 diff_4323000_4962000# gnd! 203.8fF
C1512 diff_4293000_4962000# gnd! 234.2fF
C1513 diff_4223000_4962000# gnd! 647.0fF
C1514 diff_4193000_4962000# gnd! 638.4fF
C1515 diff_4165000_4929000# gnd! 649.4fF
C1516 diff_4135000_4962000# gnd! 538.5fF
C1517 diff_4105000_4962000# gnd! 385.3fF
C1518 diff_4075000_4962000# gnd! 292.8fF
C1519 diff_4047000_4930000# gnd! 278.9fF
C1520 diff_4017000_4962000# gnd! 274.6fF
C1521 diff_3987000_4962000# gnd! 224.3fF
C1522 diff_3957000_4962000# gnd! 133.3fF
C1523 diff_3929000_4962000# gnd! 690.9fF
C1524 diff_3899000_4962000# gnd! 410.9fF
C1525 diff_3870000_4934000# gnd! 219.4fF
C1526 diff_3840000_4962000# gnd! 584.1fF
C1527 diff_3811000_4962000# gnd! 609.0fF
C1528 diff_3781000_4962000# gnd! 377.6fF
C1529 diff_3713000_4962000# gnd! 616.0fF
C1530 diff_3683000_4962000# gnd! 862.0fF
C1531 diff_3654000_3515000# gnd! 777.4fF
C1532 diff_3625000_4962000# gnd! 197.8fF
C1533 diff_3595000_4962000# gnd! 172.4fF
C1534 diff_3565000_4962000# gnd! 170.6fF
C1535 diff_3537000_4962000# gnd! 348.8fF
C1536 diff_3507000_4962000# gnd! 303.6fF
C1537 diff_3477000_4962000# gnd! 360.8fF
C1538 diff_3447000_4962000# gnd! 353.4fF
C1539 diff_3419000_4962000# gnd! 362.6fF
C1540 diff_3389000_4962000# gnd! 315.5fF
C1541 diff_3360000_4962000# gnd! 357.8fF
C1542 diff_3330000_4962000# gnd! 252.7fF
C1543 diff_3301000_4962000# gnd! 166.9fF
C1544 diff_3271000_4962000# gnd! 347.9fF
C1545 diff_3204000_4962000# gnd! 195.3fF
C1546 diff_3174000_4962000# gnd! 1132.4fF
C1547 diff_3106000_3438000# gnd! 601.0fF
C1548 diff_3116000_4962000# gnd! 220.4fF
C1549 diff_3086000_4962000# gnd! 332.1fF
C1550 diff_3056000_4962000# gnd! 166.5fF
C1551 diff_3028000_4947000# gnd! 350.1fF
C1552 diff_2998000_4962000# gnd! 329.2fF
C1553 diff_2968000_4962000# gnd! 503.0fF
C1554 diff_2849000_2986000# gnd! 631.6fF
C1555 diff_2910000_4962000# gnd! 281.2fF
C1556 diff_2880000_4962000# gnd! 216.9fF
C1557 diff_2851000_4962000# gnd! 458.1fF
C1558 diff_2821000_4962000# gnd! 171.7fF
C1559 diff_2792000_4962000# gnd! 176.7fF
C1560 diff_2762000_4962000# gnd! 191.4fF
C1561 diff_2694000_4962000# gnd! 405.8fF
C1562 diff_2664000_4962000# gnd! 563.9fF
C1563 diff_2636000_4962000# gnd! 201.1fF
C1564 diff_2606000_4947000# gnd! 696.9fF
C1565 diff_2577000_4949000# gnd! 641.9fF
C1566 diff_2547000_4962000# gnd! 342.2fF
C1567 diff_2518000_4962000# gnd! 240.9fF
C1568 diff_2488000_4962000# gnd! 222.4fF
C1569 diff_2429000_4962000# gnd! 334.6fF
C1570 diff_2399000_4962000# gnd! 316.2fF
C1571 diff_2371000_4962000# gnd! 248.2fF
C1572 diff_2341000_4962000# gnd! 304.4fF
C1573 diff_2312000_4962000# gnd! 121.4fF
C1574 diff_2282000_4962000# gnd! 131.4fF
C1575 diff_2253000_4962000# gnd! 114.7fF
C1576 diff_2223000_4962000# gnd! 116.4fF
C1577 diff_2155000_4962000# gnd! 140.1fF
C1578 diff_2125000_4962000# gnd! 352.9fF
C1579 diff_2097000_4962000# gnd! 347.4fF
C1580 diff_2067000_4962000# gnd! 335.1fF
C1581 diff_2037000_4962000# gnd! 280.6fF
C1582 diff_2007000_4962000# gnd! 275.6fF
C1583 diff_1979000_4962000# gnd! 725.8fF
C1584 diff_1949000_4962000# gnd! 343.1fF
C1585 diff_1831000_4962000# gnd! 160.2fF
C1586 diff_1801000_4962000# gnd! 334.2fF
C1587 diff_1772000_4962000# gnd! 251.4fF
C1588 diff_1742000_4962000# gnd! 262.7fF
C1589 diff_1713000_4962000# gnd! 245.4fF
C1590 diff_1683000_4962000# gnd! 238.6fF
C1591 diff_1655000_4962000# gnd! 387.1fF
C1592 diff_1625000_4962000# gnd! 743.2fF
C1593 diff_873000_3938000# gnd! 610.0fF
C1594 diff_809000_3854000# gnd! 174.5fF
C1595 diff_792000_3825000# gnd! 491.6fF
C1596 diff_752000_3797000# gnd! 100.2fF
C1597 diff_732000_3738000# gnd! 415.4fF
C1598 diff_695000_3858000# gnd! 144.8fF
C1599 diff_635000_3800000# gnd! 755.8fF
C1600 diff_650000_3859000# gnd! 157.8fF
C1601 diff_182000_3691000# gnd! 87.8fF
C1602 diff_687000_3826000# gnd! 135.6fF
C1603 diff_608000_3765000# gnd! 296.1fF
C1604 diff_185000_3712000# gnd! 192.7fF
C1605 diff_118000_3658000# gnd! 121.5fF
C1606 diff_92000_3714000# gnd! 1435.9fF
C1607 diff_570000_3597000# gnd! 911.8fF
C1608 diff_660000_3853000# gnd! 355.8fF
C1609 diff_1126000_4459000# gnd! 108.5fF
C1610 diff_1163000_4605000# gnd! 852.1fF
C1611 diff_1053000_4267000# gnd! 506.9fF
C1612 diff_991000_4386000# gnd! 175.9fF
C1613 diff_975000_4364000# gnd! 501.7fF
C1614 diff_1001000_4394000# gnd! 2055.6fF
C1615 diff_1177000_4478000# gnd! 330.4fF
C1616 diff_1197000_3119000# gnd! 2071.4fF
C1617 diff_1253000_4407000# gnd! 1024.7fF
C1618 diff_1158000_4673000# gnd! 158.0fF
C1619 diff_1076000_4557000# gnd! 610.2fF
C1620 diff_1024000_4536000# gnd! 509.6fF
C1621 diff_691000_4135000# gnd! 578.5fF
C1622 diff_659000_4117000# gnd! 537.4fF
C1623 diff_637000_4100000# gnd! 423.9fF
C1624 diff_725000_4204000# gnd! 618.5fF
C1625 diff_94000_3753000# gnd! 562.3fF
C1626 diff_139000_3844000# gnd! 327.6fF
C1627 diff_132000_3835000# gnd! 120.8fF
C1628 diff_232000_3858000# gnd! 347.9fF
C1629 diff_130000_3949000# gnd! 362.6fF
C1630 diff_106000_3785000# gnd! 452.8fF
C1631 diff_282000_4044000# gnd! 397.9fF
C1632 diff_680000_4314000# gnd! 715.2fF
C1633 diff_128000_4097000# gnd! 916.4fF
C1634 diff_222000_4165000# gnd! 94.2fF
C1635 diff_773000_4078000# gnd! 785.4fF
C1636 diff_519000_3032000# gnd! 3064.9fF
C1637 diff_936000_4586000# gnd! 441.8fF
C1638 diff_853000_4510000# gnd! 238.0fF
C1639 diff_836000_4491000# gnd! 238.4fF
C1640 diff_793000_4433000# gnd! 147.3fF
C1641 diff_757000_4475000# gnd! 1036.0fF
C1642 diff_791000_4022000# gnd! 4981.0fF
C1643 diff_654000_4324000# gnd! 107.8fF
C1644 diff_597000_3013000# gnd! 2790.0fF
C1645 diff_1014000_4730000# gnd! 533.8fF
C1646 diff_1557000_4962000# gnd! 337.1fF
C1647 diff_1528000_4962000# gnd! 365.1fF
C1648 diff_1499000_4962000# gnd! 360.8fF
C1649 diff_1469000_4962000# gnd! 369.6fF
C1650 diff_1440000_4962000# gnd! 220.2fF
C1651 diff_1410000_4962000# gnd! 226.8fF
C1652 diff_1381000_4962000# gnd! 369.6fF
C1653 diff_1351000_4962000# gnd! 660.1fF
C1654 diff_1322000_4962000# gnd! 242.2fF
C1655 diff_1292000_4962000# gnd! 221.2fF
C1656 diff_1263000_4962000# gnd! 205.4fF
C1657 diff_1233000_4962000# gnd! 218.9fF
C1658 diff_1204000_4962000# gnd! 326.4fF
C1659 diff_1145000_4574000# gnd! 342.8fF
C1660 diff_1146000_4962000# gnd! 156.9fF
C1661 diff_1038000_4590000# gnd! 361.1fF
C1662 diff_861000_4692000# gnd! 345.1fF
C1663 diff_739000_4508000# gnd! 748.8fF
C1664 diff_583000_4388000# gnd! 85.4fF
C1665 diff_578000_4447000# gnd! 328.9fF
C1666 diff_686000_4521000# gnd! 1167.2fF
C1667 diff_725000_4490000# gnd! 756.0fF
C1668 diff_101000_4084000# gnd! 728.5fF
C1669 diff_354000_4247000# gnd! 152.7fF
C1670 diff_314000_4258000# gnd! 266.1fF
C1671 diff_96000_4258000# gnd! 276.3fF
C1672 diff_78000_4235000# gnd! 718.1fF
C1673 diff_106000_4268000# gnd! 145.3fF
C1674 diff_530000_4372000# gnd! 2867.5fF
C1675 diff_512000_4352000# gnd! 1413.5fF
C1676 diff_520000_4360000# gnd! 370.1fF
C1677 diff_480000_4480000# gnd! 492.7fF
C1678 diff_88000_4249000# gnd! 363.1fF
C1679 diff_109000_4359000# gnd! 226.7fF
C1680 diff_81000_4321000# gnd! 219.6fF
C1681 diff_83000_4448000# gnd! 320.6fF
C1682 diff_65000_4220000# gnd! 3119.1fF
C1683 diff_167000_4461000# gnd! 602.6fF
C1684 diff_782000_4737000# gnd! 317.9fF
C1685 diff_642000_4583000# gnd! 480.9fF
C1686 diff_531000_4622000# gnd! 3873.2fF
C1687 diff_559000_4358000# gnd! 1013.1fF
C1688 diff_74000_3122000# gnd! 1108.5fF
C1689 diff_337000_4528000# gnd! 1103.1fF
C1690 diff_153000_4530000# gnd! 246.8fF
C1691 diff_169000_4545000# gnd! 1988.7fF
C1692 diff_216000_4574000# gnd! 86.1fF
C1693 diff_106000_4536000# gnd! 97.8fF
C1694 diff_81000_4527000# gnd! 128.2fF
C1695 diff_230000_4601000# gnd! 1060.4fF
C1696 diff_121000_4669000# gnd! 254.7fF
C1697 diff_625000_4565000# gnd! 576.6fF
C1698 diff_231000_4715000# gnd! 204.8fF
C1699 diff_205000_4722000# gnd! 83.7fF
C1700 diff_85000_4683000# gnd! 590.2fF
C1701 diff_201000_4774000# gnd! 136.4fF
C1702 diff_409000_4783000# gnd! 279.5fF
C1703 diff_78000_4695000# gnd! 912.2fF
C1704 diff_984000_4377000# gnd! 376.3fF
C1705 diff_1018000_4962000# gnd! 146.9fF
C1706 diff_988000_4962000# gnd! 154.8fF
C1707 diff_886000_3953000# gnd! 341.0fF
C1708 diff_888000_4706000# gnd! 168.2fF
C1709 diff_861000_4716000# gnd! 155.4fF
C1710 diff_831000_4716000# gnd! 156.9fF
C1711 diff_764000_4721000# gnd! 304.6fF
C1712 diff_668000_4504000# gnd! 465.1fF
C1713 diff_700000_4694000# gnd! 197.9fF
C1714 diff_446000_4910000# gnd! 983.0fF
C1715 diff_667000_3269000# gnd! 1885.5fF
C1716 diff_4952000_396000# gnd! 5980.1fF
C1717 diff_5596000_414000# gnd! 5381.2fF
C1718 diff_778000_5046000# gnd! 2672.9fF
C1719 diff_376000_4961000# gnd! 4408.3fF
C1720 diff_6226000_5161000# gnd! 414.9fF
C1721 diff_5700000_5120000# gnd! 195.7fF
C1722 diff_5502000_5120000# gnd! 542.6fF
C1723 diff_5972000_5106000# gnd! 344.4fF
C1724 diff_6074000_5171000# gnd! 96.8fF
C1725 diff_5501000_5152000# gnd! 463.6fF
C1726 diff_775000_5076000# gnd! 2459.9fF
C1727 diff_6226000_5191000# gnd! 356.8fF
C1728 diff_6074000_5195000# gnd! 101.0fF
C1729 diff_5972000_5181000# gnd! 316.5fF
C1730 diff_775000_5103000# gnd! 1570.3fF
C1731 diff_5700000_5195000# gnd! 198.5fF
C1732 diff_5502000_5195000# gnd! 545.5fF
C1733 diff_5501000_5227000# gnd! 462.2fF
C1734 diff_775000_5134000# gnd! 2039.2fF
C1735 diff_6170000_5282000# gnd! 442.8fF
C1736 diff_6012000_5272000# gnd! 112.5fF
C1737 diff_5972000_5256000# gnd! 250.3fF
C1738 diff_5600000_575000# gnd! 5707.8fF
C1739 diff_775000_5160000# gnd! 2011.6fF
C1740 diff_5700000_5270000# gnd! 199.6fF
C1741 diff_5502000_5270000# gnd! 543.8fF
C1742 diff_5501000_5302000# gnd! 460.8fF
C1743 diff_465000_5069000# gnd! 472.1fF
C1744 diff_77000_4827000# gnd! 1176.7fF
C1745 diff_487000_5098000# gnd! 450.8fF
C1746 diff_514000_5204000# gnd! 244.3fF
C1747 diff_775000_5192000# gnd! 2032.0fF
C1748 diff_5619000_1309000# gnd! 5431.2fF
C1749 diff_6170000_5342000# gnd! 362.9fF
C1750 diff_5972000_5331000# gnd! 284.4fF
C1751 diff_6012000_5360000# gnd! 104.6fF
C1752 diff_5700000_5345000# gnd! 198.9fF
C1753 diff_775000_5218000# gnd! 1818.0fF
C1754 diff_5502000_5346000# gnd! 553.9fF
C1755 diff_5501000_5377000# gnd! 459.6fF
C1756 diff_775000_5249000# gnd! 2494.0fF
C1757 diff_95000_5160000# gnd! 3666.4fF
C1758 diff_100000_3992000# gnd! 2319.4fF
C1759 diff_465000_5280000# gnd! 370.5fF
C1760 diff_502000_5322000# gnd! 127.8fF
C1761 diff_64000_4639000# gnd! 592.5fF
C1762 diff_6017000_5422000# gnd! 100.8fF
C1763 diff_6170000_5416000# gnd! 365.9fF
C1764 diff_5619000_1381000# gnd! 5380.1fF
C1765 diff_5972000_5406000# gnd! 258.9fF
C1766 diff_5619000_2102000# gnd! 4716.2fF
C1767 diff_5700000_5421000# gnd! 199.8fF
C1768 diff_775000_5275000# gnd! 1623.1fF
C1769 diff_499000_5334000# gnd! 211.4fF
C1770 diff_493000_5343000# gnd! 145.3fF
C1771 diff_5502000_5421000# gnd! 544.9fF
C1772 diff_5501000_5453000# gnd! 486.6fF
C1773 diff_775000_5306000# gnd! 2543.1fF
C1774 diff_473000_5333000# gnd! 115.9fF
C1775 diff_75000_5299000# gnd! 260.1fF
C1776 diff_6194000_5481000# gnd! 329.3fF
C1777 diff_5972000_5482000# gnd! 276.1fF
C1778 diff_6017000_5510000# gnd! 119.4fF
C1779 diff_5700000_5496000# gnd! 190.9fF
C1780 diff_775000_5333000# gnd! 2060.6fF
C1781 diff_5502000_5496000# gnd! 557.8fF
C1782 diff_5501000_5528000# gnd! 474.3fF
C1783 diff_775000_5364000# gnd! 2731.8fF
C1784 diff_6016000_5535000# gnd! 123.2fF
C1785 diff_6194000_5553000# gnd! 329.6fF
C1786 diff_5619000_2172000# gnd! 4184.0fF
C1787 diff_5972000_5557000# gnd! 242.3fF
C1788 diff_5619000_2893000# gnd! 5513.7fF
C1789 diff_5700000_5571000# gnd! 188.7fF
C1790 diff_775000_5390000# gnd! 2063.2fF
C1791 diff_5502000_5571000# gnd! 538.0fF
C1792 diff_6022000_5610000# gnd! 101.6fF
C1793 diff_5501000_5603000# gnd! 464.4fF
C1794 diff_775000_5421000# gnd! 1901.1fF
C1795 diff_6174000_5604000# gnd! 357.9fF
C1796 diff_5972000_5632000# gnd! 336.9fF
C1797 diff_6062000_5632000# gnd! 963.4fF
C1798 diff_5700000_5646000# gnd! 190.2fF
C1799 diff_402000_4713000# gnd! 1946.1fF
C1800 diff_5082000_5587000# gnd! 762.2fF
C1801 diff_775000_5448000# gnd! 1436.2fF
C1802 diff_5024000_5587000# gnd! 775.6fF
C1803 diff_5502000_5646000# gnd! 538.1fF
C1804 diff_5252000_5062000# gnd! 2182.6fF
C1805 diff_5062000_5621000# gnd! 878.6fF
C1806 diff_5004000_5621000# gnd! 868.2fF
C1807 diff_4926000_5587000# gnd! 817.4fF
C1808 diff_4867000_5587000# gnd! 826.1fF
C1809 diff_4808000_5587000# gnd! 803.7fF
C1810 diff_4906000_5621000# gnd! 902.7fF
C1811 diff_4750000_5587000# gnd! 797.8fF
C1812 diff_4847000_5621000# gnd! 925.2fF
C1813 diff_4602000_5587000# gnd! 796.7fF
C1814 diff_4788000_5621000# gnd! 886.3fF
C1815 diff_4543000_5587000# gnd! 780.2fF
C1816 diff_4730000_5621000# gnd! 902.5fF
C1817 diff_5501000_5678000# gnd! 464.4fF
C1818 diff_775000_5479000# gnd! 2193.6fF
C1819 diff_5954000_5147000# gnd! 678.4fF
C1820 diff_6105000_5745000# gnd! 142.1fF
C1821 diff_5487000_5789000# gnd! 40.3fF
C1822 diff_5775000_5847000# gnd! 2234.1fF
C1823 diff_5928000_6128000# gnd! 3101.6fF
C1824 diff_5507000_5789000# gnd! 810.0fF
C1825 diff_5402000_5747000# gnd! 597.6fF
C1826 diff_5259000_5770000# gnd! 1049.0fF
C1827 diff_4484000_5587000# gnd! 806.2fF
C1828 diff_4582000_5621000# gnd! 880.8fF
C1829 diff_4425000_5587000# gnd! 800.4fF
C1830 diff_4523000_5621000# gnd! 921.8fF
C1831 diff_4366000_5587000# gnd! 778.0fF
C1832 diff_4464000_5621000# gnd! 868.8fF
C1833 diff_4307000_5587000# gnd! 787.8fF
C1834 diff_4405000_5621000# gnd! 894.5fF
C1835 diff_4346000_5621000# gnd! 874.7fF
C1836 diff_4288000_5621000# gnd! 911.2fF
C1837 diff_4208000_5587000# gnd! 818.3fF
C1838 diff_4149000_5587000# gnd! 828.7fF
C1839 diff_4090000_5587000# gnd! 769.0fF
C1840 diff_4188000_5621000# gnd! 859.2fF
C1841 diff_4031000_5587000# gnd! 814.8fF
C1842 diff_4129000_5621000# gnd! 911.6fF
C1843 diff_3972000_5587000# gnd! 799.8fF
C1844 diff_4070000_5621000# gnd! 923.2fF
C1845 diff_3913000_5587000# gnd! 793.0fF
C1846 diff_4011000_5621000# gnd! 912.5fF
C1847 diff_3854000_5587000# gnd! 798.9fF
C1848 diff_3952000_5621000# gnd! 907.7fF
C1849 diff_3796000_5587000# gnd! 815.7fF
C1850 diff_3893000_5621000# gnd! 905.7fF
C1851 diff_3834000_5621000# gnd! 940.4fF
C1852 diff_3776000_5621000# gnd! 877.4fF
C1853 diff_3698000_5587000# gnd! 780.7fF
C1854 diff_3639000_5587000# gnd! 829.2fF
C1855 diff_3580000_5587000# gnd! 824.9fF
C1856 diff_3678000_5621000# gnd! 918.8fF
C1857 diff_3521000_5587000# gnd! 787.8fF
C1858 diff_3619000_5621000# gnd! 893.4fF
C1859 diff_3462000_5587000# gnd! 804.5fF
C1860 diff_3560000_5621000# gnd! 932.0fF
C1861 diff_3403000_5587000# gnd! 780.2fF
C1862 diff_3501000_5621000# gnd! 882.3fF
C1863 diff_3344000_5587000# gnd! 803.5fF
C1864 diff_3442000_5621000# gnd! 881.6fF
C1865 diff_3286000_5587000# gnd! 790.7fF
C1866 diff_3383000_5621000# gnd! 923.0fF
C1867 diff_3324000_5621000# gnd! 907.5fF
C1868 diff_3266000_5621000# gnd! 900.4fF
C1869 diff_3189000_5587000# gnd! 805.5fF
C1870 diff_3130000_5587000# gnd! 847.8fF
C1871 diff_3071000_5587000# gnd! 804.7fF
C1872 diff_3169000_5621000# gnd! 873.5fF
C1873 diff_3012000_5587000# gnd! 820.9fF
C1874 diff_3110000_5621000# gnd! 883.5fF
C1875 diff_2953000_5587000# gnd! 800.9fF
C1876 diff_3051000_5621000# gnd! 913.5fF
C1877 diff_2894000_5587000# gnd! 834.1fF
C1878 diff_2992000_5621000# gnd! 881.8fF
C1879 diff_2835000_5587000# gnd! 815.7fF
C1880 diff_2933000_5621000# gnd! 883.4fF
C1881 diff_2777000_5587000# gnd! 786.5fF
C1882 diff_2874000_5621000# gnd! 927.8fF
C1883 diff_2815000_5621000# gnd! 910.3fF
C1884 diff_2757000_5621000# gnd! 874.0fF
C1885 diff_2679000_5587000# gnd! 810.3fF
C1886 diff_2620000_5587000# gnd! 827.5fF
C1887 diff_2561000_5587000# gnd! 799.4fF
C1888 diff_2659000_5621000# gnd! 887.4fF
C1889 diff_2503000_5587000# gnd! 841.0fF
C1890 diff_2600000_5621000# gnd! 881.7fF
C1891 diff_2414000_5587000# gnd! 788.2fF
C1892 diff_2541000_5621000# gnd! 884.4fF
C1893 diff_2355000_5587000# gnd! 840.5fF
C1894 diff_2483000_5621000# gnd! 913.6fF
C1895 diff_4478000_4817000# gnd! 1828.8fF
C1896 diff_5173000_5735000# gnd! 893.2fF
C1897 diff_5430000_5898000# gnd! 355.1fF
C1898 diff_5453000_5802000# gnd! 320.9fF
C1899 diff_5772000_6155000# gnd! 242.7fF
C1900 diff_5761000_6140000# gnd! 2269.4fF
C1901 diff_5087000_472000# gnd! 7670.0fF
C1902 diff_5406000_5992000# gnd! 624.7fF
C1903 diff_4427000_5701000# gnd! 393.7fF
C1904 diff_4356000_5717000# gnd! 607.9fF
C1905 diff_3962000_5824000# gnd! 264.9fF
C1906 diff_4198000_5803000# gnd! 296.4fF
C1907 diff_3903000_5737000# gnd! 447.1fF
C1908 diff_3872000_5819000# gnd! 715.4fF
C1909 diff_3884000_5844000# gnd! 476.9fF
C1910 diff_3757000_5782000# gnd! 264.9fF
C1911 diff_3677000_5839000# gnd! 620.5fF
C1912 diff_3695000_5841000# gnd! 593.1fF
C1913 diff_2296000_5587000# gnd! 785.0fF
C1914 diff_2394000_5621000# gnd! 874.0fF
C1915 diff_2238000_5587000# gnd! 802.0fF
C1916 diff_2335000_5621000# gnd! 913.7fF
C1917 diff_2276000_5621000# gnd! 951.2fF
C1918 diff_2218000_5621000# gnd! 888.7fF
C1919 diff_2139000_5587000# gnd! 820.9fF
C1920 diff_2081000_5587000# gnd! 792.2fF
C1921 diff_2022000_5587000# gnd! 798.0fF
C1922 diff_2119000_5621000# gnd! 930.3fF
C1923 diff_1964000_5587000# gnd! 793.6fF
C1924 diff_2061000_5621000# gnd! 891.7fF
C1925 diff_1815000_5587000# gnd! 792.0fF
C1926 diff_2002000_5621000# gnd! 874.1fF
C1927 diff_1757000_5587000# gnd! 828.7fF
C1928 diff_1944000_5621000# gnd! 873.2fF
C1929 diff_3505000_5809000# gnd! 578.8fF
C1930 diff_3099000_5787000# gnd! 262.6fF
C1931 diff_2983000_5746000# gnd! 162.0fF
C1932 diff_3583000_5810000# gnd! 499.0fF
C1933 diff_5067000_5900000# gnd! 608.1fF
C1934 diff_4398000_6171000# gnd! 557.7fF
C1935 diff_2748000_5772000# gnd! 195.8fF
C1936 diff_1581000_4325000# gnd! 1577.3fF
C1937 diff_2523000_5770000# gnd! 322.4fF
C1938 diff_2613000_5827000# gnd! 102.7fF
C1939 diff_2621000_5834000# gnd! 415.6fF
C1940 diff_2833000_5761000# gnd! 141.5fF
C1941 diff_2841000_5928000# gnd! 662.0fF
C1942 diff_2877000_5745000# gnd! 812.0fF
C1943 diff_2975000_5983000# gnd! 53.9fF ;**FLOATING
C1944 diff_2933000_6015000# gnd! 39.3fF ;**FLOATING
C1945 diff_2887000_5984000# gnd! 68.9fF ;**FLOATING
C1946 diff_2877000_6028000# gnd! 306.6fF ;**FLOATING
C1947 diff_2157000_5726000# gnd! 23.4fF
C1948 diff_2092000_5823000# gnd! 52.5fF
C1949 diff_2071000_5823000# gnd! 16.4fF
C1950 diff_1698000_5587000# gnd! 833.4fF
C1951 diff_1795000_5621000# gnd! 909.6fF
C1952 diff_1639000_5587000# gnd! 777.6fF
C1953 diff_1737000_5621000# gnd! 867.4fF
C1954 diff_1678000_5621000# gnd! 897.4fF
C1955 diff_1619000_5621000# gnd! 894.7fF
C1956 diff_1542000_5587000# gnd! 776.2fF
C1957 diff_1484000_5587000# gnd! 785.2fF
C1958 diff_1424000_5587000# gnd! 824.2fF
C1959 diff_1522000_5621000# gnd! 933.7fF
C1960 diff_1366000_5587000# gnd! 825.4fF
C1961 diff_1464000_5621000# gnd! 898.6fF
C1962 diff_1306000_5587000# gnd! 799.7fF
C1963 diff_1404000_5621000# gnd! 879.4fF
C1964 diff_1248000_5587000# gnd! 802.3fF
C1965 diff_1346000_5621000# gnd! 854.4fF
C1966 diff_1188000_5587000# gnd! 788.0fF
C1967 diff_1286000_5621000# gnd! 887.8fF
C1968 diff_1130000_5587000# gnd! 790.9fF
C1969 diff_1228000_5621000# gnd! 856.9fF
C1970 diff_1169000_5621000# gnd! 927.2fF
C1971 diff_1110000_5621000# gnd! 892.0fF
C1972 diff_1032000_5587000# gnd! 840.9fF
C1973 diff_973000_5587000# gnd! 798.3fF
C1974 diff_914000_5587000# gnd! 787.0fF
C1975 diff_1012000_5621000# gnd! 880.6fF
C1976 diff_855000_5587000# gnd! 769.0fF
C1977 diff_953000_5621000# gnd! 921.4fF
C1978 diff_797000_5587000# gnd! 806.3fF
C1979 diff_761000_5561000# gnd! 814.8fF
C1980 diff_894000_5621000# gnd! 899.4fF
C1981 diff_835000_5621000# gnd! 885.0fF
C1982 diff_135000_5507000# gnd! 1829.3fF
C1983 diff_91000_5337000# gnd! 2367.7fF
C1984 diff_506000_5537000# gnd! 2447.4fF
C1985 diff_474000_5143000# gnd! 4409.9fF
C1986 diff_571000_4610000# gnd! 814.6fF
C1987 diff_301000_4194000# gnd! 1312.0fF
C1988 diff_2049000_5823000# gnd! 237.6fF
C1989 diff_2194000_5726000# gnd! 314.3fF
C1990 diff_88000_5400000# gnd! 1478.1fF
C1991 diff_969000_5800000# gnd! 279.8fF
C1992 diff_235000_3317000# gnd! 897.0fF
C1993 diff_836000_5746000# gnd! 293.6fF
C1994 diff_509000_5593000# gnd! 111.0fF
C1995 diff_896000_5771000# gnd! 341.0fF
C1996 diff_774000_5785000# gnd! 171.1fF
C1997 diff_72000_4515000# gnd! 28959.8fF
C1998 diff_68000_5288000# gnd! 13568.1fF
C1999 diff_94000_3551000# gnd! 4917.9fF
C2000 diff_514000_5774000# gnd! 646.0fF
C2001 diff_1586000_5876000# gnd! 214.0fF
C2002 diff_1648000_5847000# gnd! 541.9fF
C2003 diff_197000_5470000# gnd! 3124.7fF
C2004 diff_95000_5192000# gnd! 217931.0fF
C2005 diff_1586000_6057000# gnd! 1405.8fF
C2006 diff_1120000_5760000# gnd! 1785.5fF
C2007 diff_1278000_5968000# gnd! 1760.4fF
C2008 diff_1128000_5767000# gnd! 4876.3fF
C2009 diff_744000_5834000# gnd! 565.6fF
C2010 diff_1748000_6170000# gnd! 967.5fF
C2011 diff_4056000_6171000# gnd! 365.7fF
C2012 diff_83000_3098000# gnd! 487066.0fF
C2013 diff_421000_6062000# gnd! 47.8fF ;**FLOATING
C2014 diff_379000_6062000# gnd! 52.2fF ;**FLOATING
C2015 diff_338000_6062000# gnd! 52.2fF ;**FLOATING
C2016 diff_297000_6062000# gnd! 57.7fF ;**FLOATING
C2017 diff_259000_6062000# gnd! 38.8fF ;**FLOATING
C2018 diff_221000_6061000# gnd! 36.5fF ;**FLOATING
C2019 diff_161000_6062000# gnd! 67.8fF ;**FLOATING
C2020 diff_617000_6170000# gnd! 1194.0fF
