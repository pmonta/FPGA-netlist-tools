* SPICE3 file created from 4004.ext - technology: nmos

.option scale=0.4u

M1000 GND diff_6584_29296# diff_5792_29180# GND efet w=736 l=88
+ ad=3.71736e+07 pd=951320 as=121984 ps=4048 
M1001 GND GND test GND efet w=986 l=114
+ ad=0 pd=0 as=506512 ps=15104 
M1002 reset GND GND GND efet w=974 l=114
+ ad=512192 pd=15960 as=0 ps=0 
M1003 GND diff_3668_29188# diff_4204_29396# GND efet w=208 l=100
+ ad=0 pd=0 as=228624 ps=7320 
M1004 GND diff_7588_29524# diff_7520_29516# GND efet w=240 l=98
+ ad=0 pd=0 as=11744 ps=552 
M1005 GND diff_2860_29380# diff_3668_29188# GND efet w=172 l=88
+ ad=0 pd=0 as=44464 ps=1168 
M1006 diff_4204_29396# diff_2860_29380# diff_4076_29024# GND efet w=640 l=88
+ ad=0 pd=0 as=74576 ps=2224 
M1007 diff_3668_29188# Vdd Vdd GND efet w=52 l=568
+ ad=0 pd=0 as=1.42129e+07 ps=432138 
M1008 diff_3668_29188# diff_3088_28840# GND GND efet w=190 l=106
+ ad=0 pd=0 as=0 ps=0 
M1009 Vdd Vdd diff_4204_29396# GND efet w=64 l=244
+ ad=0 pd=0 as=0 ps=0 
M1010 diff_4076_29024# diff_3088_28840# GND GND efet w=1124 l=156
+ ad=0 pd=0 as=0 ps=0 
M1011 diff_3808_28348# diff_5212_23848# diff_5404_29068# GND efet w=358 l=106
+ ad=1.07288e+06 pd=29168 as=126016 ps=3752 
M1012 diff_5792_29180# diff_5200_22772# diff_3808_28348# GND efet w=400 l=94
+ ad=0 pd=0 as=0 ps=0 
M1013 diff_7520_29516# diff_7348_23696# diff_6584_29296# GND efet w=208 l=100
+ ad=0 pd=0 as=92128 ps=3216 
M1014 diff_6584_29296# diff_6496_23704# diff_4204_29396# GND efet w=112 l=100
+ ad=0 pd=0 as=0 ps=0 
M1015 GND diff_3088_28840# diff_2764_28012# GND efet w=118 l=94
+ ad=0 pd=0 as=54432 ps=2080 
M1016 Vdd diff_2740_24880# diff_2860_29380# GND efet w=70 l=106
+ ad=0 pd=0 as=27872 ps=1256 
M1017 diff_3088_28840# diff_2656_22088# diff_3808_28348# GND efet w=166 l=94
+ ad=14288 pd=584 as=0 ps=0 
M1018 diff_5408_28300# diff_5020_23836# diff_3808_28348# GND efet w=364 l=82
+ ad=115936 pd=3712 as=0 ps=0 
M1019 diff_3436_29560# diff_2656_22088# diff_2728_27904# GND efet w=160 l=88
+ ad=1.1732e+06 pd=32960 as=21536 ps=704 
M1020 diff_2764_28012# diff_2728_27904# diff_2476_25724# GND efet w=112 l=94
+ ad=0 pd=0 as=62592 ps=2008 
M1021 diff_2860_29380# diff_2728_27904# diff_2680_25724# GND efet w=208 l=88
+ ad=0 pd=0 as=42672 ps=1336 
M1022 GND diff_2728_27904# diff_4084_27448# GND efet w=1012 l=88
+ ad=0 pd=0 as=71072 ps=2016 
M1023 GND diff_424_25960# sync GND efet w=10126 l=82
+ ad=0 pd=0 as=810608 ps=18840 
M1024 diff_5408_27856# diff_5020_23836# diff_3436_29560# GND efet w=340 l=88
+ ad=107968 pd=3664 as=0 ps=0 
M1025 Vdd diff_2740_24880# diff_2984_25724# GND efet w=100 l=112
+ ad=0 pd=0 as=28784 ps=1104 
M1026 diff_424_25960# diff_460_26224# diff_424_25960# GND efet w=566 l=104
+ ad=110464 pd=4200 as=0 ps=0 
M1027 Vdd Vdd diff_460_26224# GND efet w=40 l=100
+ ad=0 pd=0 as=2720 ps=216 
M1028 Vdd diff_460_26224# diff_424_25960# GND efet w=76 l=100
+ ad=0 pd=0 as=0 ps=0 
M1029 diff_424_25492# diff_472_25516# diff_424_25492# GND efet w=560 l=104
+ ad=105712 pd=4488 as=0 ps=0 
M1030 Vdd diff_472_25516# diff_424_25492# GND efet w=88 l=88
+ ad=0 pd=0 as=0 ps=0 
M1031 Vdd Vdd diff_472_25516# GND efet w=46 l=106
+ ad=0 pd=0 as=2720 ps=216 
M1032 sync diff_424_25492# Vdd GND efet w=5614 l=100
+ ad=0 pd=0 as=0 ps=0 
M1033 diff_4204_27092# diff_2984_25724# diff_4084_27448# GND efet w=556 l=88
+ ad=219840 pd=7416 as=0 ps=0 
M1034 GND diff_2728_27904# diff_3656_27268# GND efet w=184 l=76
+ ad=0 pd=0 as=48832 ps=1240 
M1035 diff_3656_27268# Vdd Vdd GND efet w=52 l=556
+ ad=0 pd=0 as=0 ps=0 
M1036 Vdd Vdd diff_4204_27092# GND efet w=52 l=220
+ ad=0 pd=0 as=0 ps=0 
M1037 diff_3656_27268# diff_2984_25724# GND GND efet w=190 l=94
+ ad=0 pd=0 as=0 ps=0 
M1038 diff_4204_27092# diff_3656_27268# GND GND efet w=208 l=88
+ ad=0 pd=0 as=0 ps=0 
M1039 GND diff_3656_26524# diff_4204_26720# GND efet w=208 l=88
+ ad=0 pd=0 as=213984 ps=7296 
M1040 GND diff_3136_26020# diff_3656_26524# GND efet w=190 l=88
+ ad=0 pd=0 as=49936 ps=1216 
M1041 diff_4204_26720# diff_3136_26020# diff_4072_26372# GND efet w=574 l=94
+ ad=0 pd=0 as=68240 ps=2064 
M1042 diff_3656_26524# Vdd Vdd GND efet w=58 l=550
+ ad=0 pd=0 as=0 ps=0 
M1043 diff_3656_26524# diff_2428_25648# GND GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M1044 Vdd Vdd diff_4204_26720# GND efet w=58 l=238
+ ad=0 pd=0 as=0 ps=0 
M1045 diff_4072_26372# diff_2428_25648# GND GND efet w=1030 l=94
+ ad=0 pd=0 as=0 ps=0 
M1046 diff_2984_25724# diff_2428_25648# diff_2980_25568# GND efet w=188 l=144
+ ad=0 pd=0 as=9248 ps=408 
M1047 diff_2476_25724# diff_2428_25648# diff_2476_25568# GND efet w=100 l=88
+ ad=0 pd=0 as=6800 ps=336 
M1048 diff_2680_25724# diff_2428_25648# diff_2680_25568# GND efet w=184 l=88
+ ad=0 pd=0 as=12512 ps=504 
M1049 Vdd diff_2740_24880# diff_3136_26020# GND efet w=66 l=106
+ ad=0 pd=0 as=51440 ps=1880 
M1050 diff_2428_25648# diff_2656_22088# diff_3244_29488# GND efet w=160 l=88
+ ad=14672 pd=584 as=1.25806e+06 ps=35352 
M1051 diff_4204_29396# diff_6020_23524# diff_6160_28852# GND efet w=112 l=102
+ ad=0 pd=0 as=99440 ps=3176 
M1052 diff_6176_28456# diff_5144_23548# diff_4204_29396# GND efet w=112 l=88
+ ad=97472 pd=3032 as=0 ps=0 
M1053 diff_6164_27928# diff_5144_23548# diff_4204_27092# GND efet w=136 l=76
+ ad=99872 pd=3200 as=0 ps=0 
M1054 diff_3436_29560# diff_5212_23848# diff_5428_27220# GND efet w=358 l=94
+ ad=0 pd=0 as=120592 ps=3808 
M1055 diff_4204_27092# diff_6020_23524# diff_6172_27580# GND efet w=124 l=100
+ ad=0 pd=0 as=98912 ps=3056 
M1056 diff_5792_27100# diff_5200_22772# diff_3436_29560# GND efet w=382 l=82
+ ad=106336 pd=3712 as=0 ps=0 
M1057 diff_3244_29488# diff_5212_23848# diff_5428_26392# GND efet w=358 l=112
+ ad=0 pd=0 as=124432 ps=3808 
M1058 diff_5780_26516# diff_5200_22772# diff_3244_29488# GND efet w=436 l=76
+ ad=110752 pd=3856 as=0 ps=0 
M1059 diff_5408_25636# diff_5020_23836# diff_3244_29488# GND efet w=352 l=88
+ ad=115840 pd=3664 as=0 ps=0 
M1060 diff_2476_25568# diff_2428_25492# diff_2476_25408# GND efet w=100 l=88
+ ad=0 pd=0 as=67568 ps=2504 
M1061 diff_2680_25568# diff_2428_25492# diff_2680_25420# GND efet w=184 l=88
+ ad=0 pd=0 as=88576 ps=2472 
M1062 diff_2980_25568# diff_2428_25492# diff_2680_25420# GND efet w=136 l=88
+ ad=0 pd=0 as=0 ps=0 
M1063 diff_3136_26020# diff_2428_25492# diff_2680_25420# GND efet w=64 l=88
+ ad=0 pd=0 as=0 ps=0 
M1064 diff_3040_29500# diff_2656_22088# diff_2428_25492# GND efet w=184 l=94
+ ad=1.2635e+06 pd=33656 as=13376 ps=528 
M1065 GND diff_2428_25492# diff_4072_24796# GND efet w=1030 l=94
+ ad=0 pd=0 as=70256 ps=2064 
M1066 diff_2476_25408# diff_2740_24880# Vdd GND efet w=58 l=94
+ ad=0 pd=0 as=0 ps=0 
M1067 diff_5396_25448# diff_5020_23836# diff_3040_29500# GND efet w=352 l=106
+ ad=109216 pd=3664 as=0 ps=0 
M1068 Vdd diff_2740_24880# diff_3608_24316# GND efet w=82 l=112
+ ad=0 pd=0 as=19696 ps=936 
M1069 diff_4204_24416# diff_3608_24316# diff_4072_24796# GND efet w=568 l=88
+ ad=219888 pd=7296 as=0 ps=0 
M1070 GND diff_2428_25492# diff_3656_24604# GND efet w=232 l=88
+ ad=0 pd=0 as=48592 ps=1312 
M1071 diff_3656_24604# Vdd Vdd GND efet w=58 l=550
+ ad=0 pd=0 as=0 ps=0 
M1072 Vdd Vdd diff_4204_24416# GND efet w=52 l=220
+ ad=0 pd=0 as=0 ps=0 
M1073 GND diff_2788_24040# diff_2680_25420# GND efet w=256 l=100
+ ad=0 pd=0 as=0 ps=0 
M1074 diff_3656_24604# diff_3608_24316# GND GND efet w=172 l=76
+ ad=0 pd=0 as=0 ps=0 
M1075 GND diff_424_25492# diff_424_25960# GND efet w=832 l=100
+ ad=0 pd=0 as=0 ps=0 
M1076 diff_3608_24316# diff_2788_24040# GND GND efet w=112 l=88
+ ad=0 pd=0 as=0 ps=0 
M1077 diff_4204_24416# diff_3656_24604# GND GND efet w=220 l=76
+ ad=0 pd=0 as=0 ps=0 
M1078 diff_2476_25408# diff_2788_24040# diff_2836_23896# GND efet w=112 l=88
+ ad=0 pd=0 as=28784 ps=1088 
M1079 GND diff_928_20116# diff_424_25492# GND efet w=922 l=106
+ ad=0 pd=0 as=0 ps=0 
M1080 GND diff_8704_29524# diff_8636_29492# GND efet w=204 l=116
+ ad=0 pd=0 as=10304 ps=552 
M1081 diff_8276_29332# diff_8096_29188# GND GND efet w=154 l=82
+ ad=12800 pd=552 as=0 ps=0 
M1082 diff_6584_29296# diff_8020_23696# diff_8276_29332# GND efet w=214 l=94
+ ad=0 pd=0 as=0 ps=0 
M1083 diff_8636_29492# diff_8548_23696# diff_6584_29296# GND efet w=208 l=94
+ ad=0 pd=0 as=0 ps=0 
M1084 diff_6584_29296# diff_9232_23696# diff_9392_29332# GND efet w=226 l=94
+ ad=0 pd=0 as=13184 ps=600 
M1085 diff_9392_29332# diff_9224_29188# GND GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M1086 diff_5404_29068# diff_6160_28852# GND GND efet w=596 l=126
+ ad=0 pd=0 as=0 ps=0 
M1087 diff_5792_29180# diff_7576_23716# diff_7588_29524# GND efet w=46 l=94
+ ad=0 pd=0 as=3344 ps=264 
M1088 diff_8096_29188# diff_7816_23824# diff_5792_29180# GND efet w=58 l=82
+ ad=3008 pd=264 as=0 ps=0 
M1089 diff_5404_29068# diff_7576_23716# diff_7588_28744# GND efet w=46 l=94
+ ad=0 pd=0 as=3200 ps=240 
M1090 diff_8096_29044# diff_7816_23824# diff_5404_29068# GND efet w=40 l=76
+ ad=3200 pd=240 as=0 ps=0 
M1091 diff_7508_28748# diff_7348_23696# diff_6160_28852# GND efet w=220 l=88
+ ad=12656 pd=576 as=0 ps=0 
M1092 GND diff_7588_28744# diff_7508_28748# GND efet w=198 l=122
+ ad=0 pd=0 as=0 ps=0 
M1093 diff_5792_29180# diff_8788_23696# diff_8704_29524# GND efet w=46 l=94
+ ad=0 pd=0 as=3344 ps=264 
M1094 diff_9224_29188# diff_9028_23696# diff_5792_29180# GND efet w=40 l=88
+ ad=2864 pd=240 as=0 ps=0 
M1095 diff_5404_29068# diff_8788_23696# diff_8704_28756# GND efet w=46 l=94
+ ad=0 pd=0 as=3200 ps=240 
M1096 diff_9224_29044# diff_9028_23696# diff_5404_29068# GND efet w=40 l=100
+ ad=3440 pd=288 as=0 ps=0 
M1097 GND diff_6176_28456# diff_5408_28300# GND efet w=592 l=106
+ ad=0 pd=0 as=0 ps=0 
M1098 diff_7520_28604# diff_7348_23696# diff_6176_28456# GND efet w=196 l=82
+ ad=11024 pd=552 as=0 ps=0 
M1099 GND diff_7588_28636# diff_7520_28604# GND efet w=192 l=122
+ ad=0 pd=0 as=0 ps=0 
M1100 diff_8276_28780# diff_8096_29044# GND GND efet w=174 l=110
+ ad=13616 pd=600 as=0 ps=0 
M1101 diff_6160_28852# diff_8020_23696# diff_8276_28780# GND efet w=220 l=88
+ ad=0 pd=0 as=0 ps=0 
M1102 diff_8636_28744# diff_8548_23696# diff_6160_28852# GND efet w=214 l=82
+ ad=14432 pd=576 as=0 ps=0 
M1103 GND diff_8704_28756# diff_8636_28744# GND efet w=186 l=94
+ ad=0 pd=0 as=0 ps=0 
M1104 diff_5408_27856# diff_6164_27928# GND GND efet w=580 l=106
+ ad=0 pd=0 as=0 ps=0 
M1105 diff_5408_28300# diff_7576_23716# diff_7588_28636# GND efet w=58 l=94
+ ad=0 pd=0 as=3728 ps=312 
M1106 diff_8276_28444# diff_8096_28300# GND GND efet w=186 l=122
+ ad=13520 pd=576 as=0 ps=0 
M1107 Vdd diff_8680_20596# diff_6584_29296# GND efet w=64 l=88
+ ad=0 pd=0 as=0 ps=0 
M1108 diff_10996_29140# diff_2656_22088# diff_3040_29500# GND efet w=112 l=100
+ ad=5744 pd=408 as=0 ps=0 
M1109 diff_11180_28768# diff_12328_25804# diff_12256_29344# GND efet w=136 l=100
+ ad=132064 pd=3816 as=134400 ps=4160 
M1110 GND diff_12256_29344# diff_11788_29092# GND efet w=520 l=88
+ ad=0 pd=0 as=139616 ps=4752 
M1111 Vdd Vdd diff_5792_29180# GND efet w=46 l=250
+ ad=0 pd=0 as=0 ps=0 
M1112 GND diff_10996_29140# diff_11180_28768# GND efet w=898 l=94
+ ad=0 pd=0 as=0 ps=0 
M1113 Vdd Vdd diff_5404_29068# GND efet w=50 l=254
+ ad=0 pd=0 as=0 ps=0 
M1114 GND diff_8716_28612# diff_8636_28604# GND efet w=198 l=98
+ ad=0 pd=0 as=13712 ps=576 
M1115 diff_6176_28456# diff_8020_23696# diff_8276_28444# GND efet w=202 l=88
+ ad=0 pd=0 as=0 ps=0 
M1116 diff_8636_28604# diff_8548_23696# diff_6176_28456# GND efet w=214 l=82
+ ad=0 pd=0 as=0 ps=0 
M1117 diff_9392_28796# diff_9224_29044# GND GND efet w=186 l=110
+ ad=13328 pd=552 as=0 ps=0 
M1118 diff_6160_28852# diff_9232_23696# diff_9392_28796# GND efet w=214 l=82
+ ad=0 pd=0 as=0 ps=0 
M1119 Vdd diff_8680_20596# diff_6160_28852# GND efet w=70 l=100
+ ad=0 pd=0 as=0 ps=0 
M1120 diff_3040_29500# diff_11872_25876# diff_11788_29092# GND efet w=376 l=88
+ ad=0 pd=0 as=0 ps=0 
M1121 diff_12236_28852# diff_12136_25792# diff_3040_29500# GND efet w=370 l=100
+ ad=129008 pd=4560 as=0 ps=0 
M1122 diff_11180_28768# Vdd Vdd GND efet w=58 l=178
+ ad=0 pd=0 as=0 ps=0 
M1123 diff_9392_28444# diff_9224_28300# GND GND efet w=186 l=110
+ ad=13664 pd=576 as=0 ps=0 
M1124 diff_6176_28456# diff_9232_23696# diff_9392_28444# GND efet w=226 l=82
+ ad=0 pd=0 as=0 ps=0 
M1125 diff_8096_28300# diff_7816_23824# diff_5408_28300# GND efet w=46 l=76
+ ad=3488 pd=264 as=0 ps=0 
M1126 diff_5408_27856# diff_7576_23716# diff_7588_27856# GND efet w=40 l=76
+ ad=0 pd=0 as=3200 ps=240 
M1127 diff_8096_28156# diff_7816_23824# diff_5408_27856# GND efet w=40 l=76
+ ad=3200 pd=240 as=0 ps=0 
M1128 diff_7508_27856# diff_7348_23696# diff_6164_27928# GND efet w=226 l=82
+ ad=12608 pd=600 as=0 ps=0 
M1129 GND diff_7588_27856# diff_7508_27856# GND efet w=192 l=104
+ ad=0 pd=0 as=0 ps=0 
M1130 diff_5408_28300# diff_8788_23696# diff_8716_28612# GND efet w=46 l=94
+ ad=0 pd=0 as=3392 ps=288 
M1131 Vdd diff_8680_20596# diff_6176_28456# GND efet w=70 l=106
+ ad=0 pd=0 as=0 ps=0 
M1132 diff_11180_28552# Vdd Vdd GND efet w=58 l=166
+ ad=122320 pd=3648 as=0 ps=0 
M1133 diff_9224_28300# diff_9028_23696# diff_5408_28300# GND efet w=40 l=88
+ ad=3200 pd=240 as=0 ps=0 
M1134 diff_5408_27856# diff_8788_23696# diff_8704_27856# GND efet w=46 l=76
+ ad=0 pd=0 as=3200 ps=240 
M1135 diff_9224_28156# diff_9028_23696# diff_5408_27856# GND efet w=40 l=88
+ ad=3392 pd=264 as=0 ps=0 
M1136 GND diff_6172_27580# diff_5428_27220# GND efet w=520 l=88
+ ad=0 pd=0 as=0 ps=0 
M1137 diff_7520_27716# diff_7348_23696# diff_6172_27580# GND efet w=196 l=82
+ ad=11216 pd=528 as=0 ps=0 
M1138 GND diff_7588_27736# diff_7520_27716# GND efet w=192 l=116
+ ad=0 pd=0 as=0 ps=0 
M1139 diff_8264_27920# diff_8096_28156# GND GND efet w=186 l=110
+ ad=12896 pd=576 as=0 ps=0 
M1140 diff_6164_27928# diff_8020_23696# diff_8264_27920# GND efet w=208 l=88
+ ad=0 pd=0 as=0 ps=0 
M1141 diff_8636_27856# diff_8548_23696# diff_6164_27928# GND efet w=214 l=82
+ ad=14240 pd=576 as=0 ps=0 
M1142 GND diff_8704_27856# diff_8636_27856# GND efet w=192 l=92
+ ad=0 pd=0 as=0 ps=0 
M1143 Vdd Vdd diff_5408_28300# GND efet w=52 l=256
+ ad=0 pd=0 as=0 ps=0 
M1144 GND diff_10996_28180# diff_11180_28552# GND efet w=940 l=88
+ ad=0 pd=0 as=0 ps=0 
M1145 Vdd Vdd diff_5408_27856# GND efet w=50 l=246
+ ad=0 pd=0 as=0 ps=0 
M1146 diff_9392_27908# diff_9224_28156# GND GND efet w=186 l=146
+ ad=13712 pd=576 as=0 ps=0 
M1147 diff_8276_27568# diff_8096_27412# GND GND efet w=174 l=122
+ ad=11936 pd=552 as=0 ps=0 
M1148 GND diff_8704_27736# diff_8636_27692# GND efet w=186 l=98
+ ad=0 pd=0 as=13328 ps=552 
M1149 diff_6172_27580# diff_8020_23696# diff_8276_27568# GND efet w=214 l=82
+ ad=0 pd=0 as=0 ps=0 
M1150 diff_8636_27692# diff_8548_23696# diff_6172_27580# GND efet w=202 l=82
+ ad=0 pd=0 as=0 ps=0 
M1151 diff_6164_27928# diff_9232_23696# diff_9392_27908# GND efet w=208 l=88
+ ad=0 pd=0 as=0 ps=0 
M1152 Vdd diff_8680_20596# diff_6164_27928# GND efet w=64 l=100
+ ad=0 pd=0 as=0 ps=0 
M1153 diff_3244_29488# diff_11872_25876# diff_11800_28096# GND efet w=364 l=88
+ ad=0 pd=0 as=134672 ps=4584 
M1154 diff_12236_28156# diff_12136_25792# diff_3244_29488# GND efet w=376 l=88
+ ad=129824 pd=4536 as=0 ps=0 
M1155 diff_12680_28816# diff_12544_25804# diff_11180_28768# GND efet w=106 l=100
+ ad=138992 pd=4200 as=0 ps=0 
M1156 diff_12236_28852# diff_12680_28816# GND GND efet w=484 l=88
+ ad=0 pd=0 as=0 ps=0 
M1157 diff_13844_29468# diff_13744_27736# diff_12256_29344# GND efet w=196 l=100
+ ad=10544 pd=528 as=0 ps=0 
M1158 GND diff_13912_29200# diff_13844_29468# GND efet w=204 l=116
+ ad=0 pd=0 as=0 ps=0 
M1159 diff_14600_29332# diff_14420_29176# GND GND efet w=192 l=116
+ ad=10016 pd=504 as=0 ps=0 
M1160 diff_12256_29344# diff_14416_25448# diff_14600_29332# GND efet w=196 l=100
+ ad=0 pd=0 as=0 ps=0 
M1161 diff_14960_29468# diff_14860_29452# diff_12256_29344# GND efet w=208 l=100
+ ad=12224 pd=528 as=0 ps=0 
M1162 GND diff_15028_29188# diff_14960_29468# GND efet w=186 l=110
+ ad=0 pd=0 as=0 ps=0 
M1163 diff_15716_29332# diff_15536_29176# GND GND efet w=198 l=134
+ ad=9728 pd=504 as=0 ps=0 
M1164 diff_12256_29344# diff_15592_25448# diff_15716_29332# GND efet w=196 l=106
+ ad=0 pd=0 as=0 ps=0 
M1165 diff_16076_29492# diff_15976_29452# diff_12256_29344# GND efet w=208 l=112
+ ad=10448 pd=552 as=0 ps=0 
M1166 GND diff_16132_29488# diff_16076_29492# GND efet w=210 l=158
+ ad=0 pd=0 as=0 ps=0 
M1167 diff_16832_29320# diff_16652_29176# GND GND efet w=198 l=110
+ ad=9632 pd=576 as=0 ps=0 
M1168 diff_12256_29344# diff_16768_25436# diff_16832_29320# GND efet w=244 l=100
+ ad=0 pd=0 as=0 ps=0 
M1169 diff_11788_29092# diff_13972_25448# diff_13912_29200# GND efet w=40 l=88
+ ad=0 pd=0 as=2816 ps=264 
M1170 diff_14420_29176# diff_14224_25448# diff_11788_29092# GND efet w=40 l=88
+ ad=2864 pd=240 as=0 ps=0 
M1171 diff_11788_29092# diff_15148_25448# diff_15028_29188# GND efet w=46 l=94
+ ad=0 pd=0 as=3008 ps=264 
M1172 diff_12236_28852# diff_13972_25448# diff_13900_28732# GND efet w=40 l=88
+ ad=0 pd=0 as=2720 ps=216 
M1173 diff_14420_29032# diff_14224_25448# diff_12236_28852# GND efet w=40 l=88
+ ad=3008 pd=264 as=0 ps=0 
M1174 diff_13832_28732# diff_13744_27736# diff_12680_28816# GND efet w=220 l=100
+ ad=12800 pd=576 as=0 ps=0 
M1175 GND diff_13900_28732# diff_13832_28732# GND efet w=192 l=98
+ ad=0 pd=0 as=0 ps=0 
M1176 diff_15536_29176# diff_15388_25448# diff_11788_29092# GND efet w=40 l=88
+ ad=3200 pd=240 as=0 ps=0 
M1177 GND diff_13900_28612# diff_13832_28604# GND efet w=186 l=110
+ ad=0 pd=0 as=12032 ps=552 
M1178 diff_10996_28180# diff_2656_22088# diff_3244_29488# GND efet w=100 l=88
+ ad=10400 pd=408 as=0 ps=0 
M1179 diff_9392_27568# diff_9212_27412# GND GND efet w=192 l=134
+ ad=12800 pd=552 as=0 ps=0 
M1180 diff_6172_27580# diff_9232_23696# diff_9392_27568# GND efet w=202 l=82
+ ad=0 pd=0 as=0 ps=0 
M1181 GND diff_6584_27052# diff_5792_27100# GND efet w=562 l=106
+ ad=0 pd=0 as=0 ps=0 
M1182 diff_6584_27052# diff_6496_23704# diff_4204_27092# GND efet w=100 l=88
+ ad=94432 pd=3000 as=0 ps=0 
M1183 diff_5428_27220# diff_7576_23716# diff_7588_27736# GND efet w=58 l=94
+ ad=0 pd=0 as=4448 ps=288 
M1184 diff_8096_27412# diff_7816_23824# diff_5428_27220# GND efet w=40 l=94
+ ad=3584 pd=312 as=0 ps=0 
M1185 diff_5792_27100# diff_7576_23716# diff_7588_26968# GND efet w=40 l=76
+ ad=0 pd=0 as=3680 ps=264 
M1186 diff_8096_27268# diff_7816_23824# diff_5792_27100# GND efet w=40 l=76
+ ad=3200 pd=240 as=0 ps=0 
M1187 diff_7508_26968# diff_7348_23696# diff_6584_27052# GND efet w=220 l=82
+ ad=12656 pd=576 as=0 ps=0 
M1188 GND diff_7588_26968# diff_7508_26968# GND efet w=186 l=98
+ ad=0 pd=0 as=0 ps=0 
M1189 diff_5428_27220# diff_8788_23696# diff_8704_27736# GND efet w=46 l=82
+ ad=0 pd=0 as=3488 ps=288 
M1190 diff_9212_27412# diff_9028_23696# diff_5428_27220# GND efet w=40 l=76
+ ad=3680 pd=264 as=0 ps=0 
M1191 diff_5792_27100# diff_8788_23696# diff_8704_26968# GND efet w=40 l=76
+ ad=0 pd=0 as=3200 ps=240 
M1192 diff_9212_27268# diff_9028_23696# diff_5792_27100# GND efet w=40 l=76
+ ad=3680 pd=264 as=0 ps=0 
M1193 GND diff_6572_26696# diff_5780_26516# GND efet w=598 l=94
+ ad=0 pd=0 as=0 ps=0 
M1194 diff_6572_26696# diff_6496_23704# diff_4204_26720# GND efet w=112 l=82
+ ad=93136 pd=3056 as=0 ps=0 
M1195 diff_4204_26720# diff_6020_23524# diff_6172_26164# GND efet w=112 l=100
+ ad=0 pd=0 as=99968 ps=3200 
M1196 diff_7508_26840# diff_7348_23696# diff_6572_26696# GND efet w=214 l=82
+ ad=11648 pd=552 as=0 ps=0 
M1197 GND diff_7588_26848# diff_7508_26840# GND efet w=192 l=104
+ ad=0 pd=0 as=0 ps=0 
M1198 diff_8276_27004# diff_8096_27268# GND GND efet w=180 l=116
+ ad=13328 pd=552 as=0 ps=0 
M1199 diff_6584_27052# diff_8020_23696# diff_8276_27004# GND efet w=220 l=88
+ ad=0 pd=0 as=0 ps=0 
M1200 diff_8636_26968# diff_8548_23696# diff_6584_27052# GND efet w=220 l=88
+ ad=14384 pd=576 as=0 ps=0 
M1201 GND diff_8704_26968# diff_8636_26968# GND efet w=192 l=92
+ ad=0 pd=0 as=0 ps=0 
M1202 Vdd diff_8680_20596# diff_6172_27580# GND efet w=64 l=88
+ ad=0 pd=0 as=0 ps=0 
M1203 diff_10996_27364# diff_2656_22088# diff_3436_29560# GND efet w=112 l=100
+ ad=11600 pd=432 as=0 ps=0 
M1204 diff_6152_25792# diff_5144_23548# diff_4204_26720# GND efet w=112 l=100
+ ad=96704 pd=3032 as=0 ps=0 
M1205 diff_6152_25264# diff_5144_23548# diff_4204_24416# GND efet w=118 l=94
+ ad=96800 pd=3128 as=0 ps=0 
M1206 diff_5428_26392# diff_6172_26164# GND GND efet w=538 l=82
+ ad=0 pd=0 as=0 ps=0 
M1207 diff_5780_26516# diff_7576_23716# diff_7588_26848# GND efet w=46 l=100
+ ad=0 pd=0 as=3632 ps=288 
M1208 diff_8264_26680# diff_8096_26524# GND GND efet w=180 l=116
+ ad=14096 pd=552 as=0 ps=0 
M1209 GND diff_8704_26848# diff_8624_26828# GND efet w=204 l=104
+ ad=0 pd=0 as=13424 ps=576 
M1210 diff_6572_26696# diff_8020_23696# diff_8264_26680# GND efet w=202 l=94
+ ad=0 pd=0 as=0 ps=0 
M1211 diff_8624_26828# diff_8548_23696# diff_6572_26696# GND efet w=208 l=88
+ ad=0 pd=0 as=0 ps=0 
M1212 diff_9392_27008# diff_9212_27268# GND GND efet w=192 l=104
+ ad=13280 pd=552 as=0 ps=0 
M1213 diff_6584_27052# diff_9232_23696# diff_9392_27008# GND efet w=208 l=88
+ ad=0 pd=0 as=0 ps=0 
M1214 Vdd Vdd diff_5428_27220# GND efet w=46 l=238
+ ad=0 pd=0 as=0 ps=0 
M1215 GND diff_10996_27364# diff_11180_26992# GND efet w=898 l=82
+ ad=0 pd=0 as=126544 ps=3600 
M1216 diff_3436_29560# diff_11872_25876# diff_11800_27280# GND efet w=358 l=94
+ ad=0 pd=0 as=133760 ps=4544 
M1217 Vdd Vdd diff_5792_27100# GND efet w=50 l=234
+ ad=0 pd=0 as=0 ps=0 
M1218 Vdd diff_8680_20596# diff_6584_27052# GND efet w=76 l=88
+ ad=0 pd=0 as=0 ps=0 
M1219 diff_12680_28456# diff_12544_25804# diff_11180_28552# GND efet w=100 l=100
+ ad=137120 pd=4200 as=0 ps=0 
M1220 diff_11180_28552# diff_12328_25804# diff_12256_27952# GND efet w=100 l=88
+ ad=0 pd=0 as=141744 ps=4352 
M1221 diff_11180_26992# diff_12328_25804# diff_12256_27580# GND efet w=100 l=88
+ ad=0 pd=0 as=140064 ps=4304 
M1222 diff_9392_26668# diff_9212_26524# GND GND efet w=198 l=110
+ ad=13040 pd=552 as=0 ps=0 
M1223 diff_8096_26524# diff_7816_23824# diff_5780_26516# GND efet w=40 l=88
+ ad=3344 pd=264 as=0 ps=0 
M1224 diff_8096_26380# diff_7816_23824# diff_5428_26392# GND efet w=40 l=100
+ ad=3200 pd=240 as=0 ps=0 
M1225 diff_5428_26392# diff_7576_23716# diff_7588_26080# GND efet w=40 l=88
+ ad=0 pd=0 as=3200 ps=240 
M1226 diff_7508_26080# diff_7348_23696# diff_6172_26164# GND efet w=226 l=82
+ ad=13088 pd=576 as=0 ps=0 
M1227 GND diff_7588_26080# diff_7508_26080# GND efet w=186 l=98
+ ad=0 pd=0 as=0 ps=0 
M1228 diff_6572_26696# diff_9232_23696# diff_9392_26668# GND efet w=202 l=94
+ ad=0 pd=0 as=0 ps=0 
M1229 diff_5780_26516# diff_8788_23696# diff_8704_26848# GND efet w=40 l=76
+ ad=0 pd=0 as=3344 ps=264 
M1230 diff_9212_26524# diff_9028_23696# diff_5780_26516# GND efet w=40 l=76
+ ad=3344 pd=264 as=0 ps=0 
M1231 diff_5428_26392# diff_8788_23696# diff_8704_26080# GND efet w=40 l=76
+ ad=0 pd=0 as=3200 ps=240 
M1232 diff_9212_26380# diff_9028_23696# diff_5428_26392# GND efet w=40 l=88
+ ad=3200 pd=240 as=0 ps=0 
M1233 diff_8264_26128# diff_8096_26380# GND GND efet w=186 l=98
+ ad=14672 pd=600 as=0 ps=0 
M1234 GND diff_7588_25948# diff_7508_25952# GND efet w=198 l=110
+ ad=0 pd=0 as=11792 ps=552 
M1235 GND diff_6152_25792# diff_5408_25636# GND efet w=568 l=88
+ ad=0 pd=0 as=0 ps=0 
M1236 diff_7508_25952# diff_7348_23696# diff_6152_25792# GND efet w=202 l=82
+ ad=0 pd=0 as=0 ps=0 
M1237 diff_6172_26164# diff_8020_23696# diff_8264_26128# GND efet w=214 l=82
+ ad=0 pd=0 as=0 ps=0 
M1238 diff_8636_26080# diff_8548_23696# diff_6172_26164# GND efet w=208 l=88
+ ad=13616 pd=600 as=0 ps=0 
M1239 GND diff_8704_26080# diff_8636_26080# GND efet w=204 l=92
+ ad=0 pd=0 as=0 ps=0 
M1240 diff_5396_25448# diff_6152_25264# GND GND efet w=556 l=100
+ ad=0 pd=0 as=0 ps=0 
M1241 diff_8264_25820# diff_8096_25636# GND GND efet w=192 l=104
+ ad=13904 pd=600 as=0 ps=0 
M1242 GND diff_8704_25960# diff_8636_25916# GND efet w=186 l=98
+ ad=0 pd=0 as=13472 ps=552 
M1243 diff_6152_25792# diff_8020_23696# diff_8264_25820# GND efet w=208 l=88
+ ad=0 pd=0 as=0 ps=0 
M1244 diff_8636_25916# diff_8548_23696# diff_6152_25792# GND efet w=208 l=88
+ ad=0 pd=0 as=0 ps=0 
M1245 diff_9392_26120# diff_9212_26380# GND GND efet w=186 l=110
+ ad=12320 pd=528 as=0 ps=0 
M1246 diff_6172_26164# diff_9232_23696# diff_9392_26120# GND efet w=196 l=88
+ ad=0 pd=0 as=0 ps=0 
M1247 diff_11180_26992# Vdd Vdd GND efet w=52 l=160
+ ad=0 pd=0 as=0 ps=0 
M1248 Vdd diff_8680_20596# diff_6572_26696# GND efet w=70 l=106
+ ad=0 pd=0 as=0 ps=0 
M1249 Vdd Vdd diff_5780_26516# GND efet w=44 l=240
+ ad=0 pd=0 as=0 ps=0 
M1250 diff_11180_26776# Vdd Vdd GND efet w=58 l=160
+ ad=120256 pd=3696 as=0 ps=0 
M1251 GND diff_10996_26404# diff_11180_26776# GND efet w=940 l=100
+ ad=0 pd=0 as=0 ps=0 
M1252 diff_12236_27076# diff_12136_25792# diff_3436_29560# GND efet w=364 l=88
+ ad=126128 pd=4584 as=0 ps=0 
M1253 GND diff_12680_28456# diff_12236_28156# GND efet w=484 l=88
+ ad=0 pd=0 as=0 ps=0 
M1254 diff_11800_28096# diff_12256_27952# GND GND efet w=490 l=82
+ ad=0 pd=0 as=0 ps=0 
M1255 diff_13832_28604# diff_13744_27736# diff_12680_28456# GND efet w=208 l=88
+ ad=0 pd=0 as=0 ps=0 
M1256 diff_14588_28784# diff_14420_29032# GND GND efet w=228 l=116
+ ad=12224 pd=600 as=0 ps=0 
M1257 diff_12680_28816# diff_14416_25448# diff_14588_28784# GND efet w=220 l=88
+ ad=0 pd=0 as=0 ps=0 
M1258 diff_14948_28736# diff_14860_29452# diff_12680_28816# GND efet w=208 l=100
+ ad=12224 pd=552 as=0 ps=0 
M1259 diff_12236_28852# diff_15148_25448# diff_15028_28720# GND efet w=40 l=88
+ ad=0 pd=0 as=2720 ps=216 
M1260 diff_15536_29032# diff_15388_25448# diff_12236_28852# GND efet w=40 l=88
+ ad=3200 pd=240 as=0 ps=0 
M1261 GND diff_15028_28720# diff_14948_28736# GND efet w=168 l=104
+ ad=0 pd=0 as=0 ps=0 
M1262 diff_15716_28780# diff_15536_29032# GND GND efet w=192 l=128
+ ad=9920 pd=528 as=0 ps=0 
M1263 diff_17192_29468# diff_17092_28684# diff_12256_29344# GND efet w=220 l=100
+ ad=10304 pd=552 as=0 ps=0 
M1264 GND diff_17248_29488# diff_17192_29468# GND efet w=210 l=156
+ ad=0 pd=0 as=0 ps=0 
M1265 diff_17948_29320# diff_17780_29176# GND GND efet w=216 l=104
+ ad=9200 pd=552 as=0 ps=0 
M1266 diff_12256_29344# diff_17932_25436# diff_17948_29320# GND efet w=232 l=106
+ ad=0 pd=0 as=0 ps=0 
M1267 diff_12680_28816# diff_15592_25448# diff_15716_28780# GND efet w=214 l=106
+ ad=0 pd=0 as=0 ps=0 
M1268 diff_11788_29092# diff_16312_25436# diff_16132_29488# GND efet w=40 l=100
+ ad=0 pd=0 as=2864 ps=240 
M1269 diff_16652_29176# diff_16516_26800# diff_11788_29092# GND efet w=58 l=94
+ ad=2672 pd=240 as=0 ps=0 
M1270 diff_12236_28852# diff_16312_25436# diff_16144_28720# GND efet w=52 l=100
+ ad=0 pd=0 as=2720 ps=216 
M1271 GND diff_16144_28720# diff_16076_28732# GND efet w=168 l=116
+ ad=0 pd=0 as=12224 ps=528 
M1272 diff_16652_29032# diff_16516_26800# diff_12236_28852# GND efet w=46 l=94
+ ad=3008 pd=240 as=0 ps=0 
M1273 diff_16076_28732# diff_15976_29452# diff_12680_28816# GND efet w=196 l=88
+ ad=0 pd=0 as=0 ps=0 
M1274 diff_14588_28444# diff_14420_28288# GND GND efet w=210 l=122
+ ad=12512 pd=624 as=0 ps=0 
M1275 diff_12236_28156# diff_13972_25448# diff_13900_28612# GND efet w=40 l=88
+ ad=0 pd=0 as=3056 ps=264 
M1276 GND diff_15028_28612# diff_14948_28604# GND efet w=180 l=122
+ ad=0 pd=0 as=12272 ps=576 
M1277 diff_12680_28456# diff_14416_25448# diff_14588_28444# GND efet w=226 l=82
+ ad=0 pd=0 as=0 ps=0 
M1278 diff_14948_28604# diff_14860_29452# diff_12680_28456# GND efet w=202 l=82
+ ad=0 pd=0 as=0 ps=0 
M1279 diff_11788_29092# diff_17440_26356# diff_17248_29488# GND efet w=40 l=100
+ ad=0 pd=0 as=2720 ps=216 
M1280 diff_17780_29176# diff_17632_26752# diff_11788_29092# GND efet w=40 l=112
+ ad=2240 pd=192 as=0 ps=0 
M1281 diff_12236_28852# diff_17440_26356# diff_17272_28708# GND efet w=52 l=106
+ ad=0 pd=0 as=2912 ps=240 
M1282 diff_17780_29020# diff_17632_26752# diff_12236_28852# GND efet w=58 l=118
+ ad=3056 pd=240 as=0 ps=0 
M1283 diff_15704_28432# diff_15536_28288# GND GND efet w=198 l=134
+ ad=12368 pd=624 as=0 ps=0 
M1284 diff_14420_28288# diff_14224_25448# diff_12236_28156# GND efet w=40 l=88
+ ad=3200 pd=240 as=0 ps=0 
M1285 diff_11800_28096# diff_13972_25448# diff_13912_27832# GND efet w=40 l=88
+ ad=0 pd=0 as=2720 ps=216 
M1286 diff_14420_28144# diff_14224_25448# diff_11800_28096# GND efet w=40 l=88
+ ad=3200 pd=240 as=0 ps=0 
M1287 diff_13832_27860# diff_13744_27736# diff_12256_27952# GND efet w=220 l=88
+ ad=12176 pd=552 as=0 ps=0 
M1288 GND diff_13912_27832# diff_13832_27860# GND efet w=180 l=104
+ ad=0 pd=0 as=0 ps=0 
M1289 diff_12236_28156# diff_15148_25448# diff_15028_28612# GND efet w=46 l=82
+ ad=0 pd=0 as=3152 ps=264 
M1290 diff_12680_28456# diff_15592_25448# diff_15704_28432# GND efet w=220 l=100
+ ad=0 pd=0 as=0 ps=0 
M1291 diff_16076_28580# diff_15976_29452# diff_12680_28456# GND efet w=202 l=100
+ ad=12656 pd=552 as=0 ps=0 
M1292 GND diff_16144_28612# diff_16076_28580# GND efet w=174 l=110
+ ad=0 pd=0 as=0 ps=0 
M1293 diff_16832_28768# diff_16652_29032# GND GND efet w=210 l=110
+ ad=9584 pd=528 as=0 ps=0 
M1294 diff_12680_28816# diff_16768_25436# diff_16832_28768# GND efet w=202 l=94
+ ad=0 pd=0 as=0 ps=0 
M1295 diff_17192_28732# diff_17092_28684# diff_12680_28816# GND efet w=202 l=94
+ ad=12896 pd=528 as=0 ps=0 
M1296 GND diff_17272_28708# diff_17192_28732# GND efet w=160 l=100
+ ad=0 pd=0 as=0 ps=0 
M1297 diff_16832_28432# diff_16652_28288# GND GND efet w=204 l=104
+ ad=10160 pd=552 as=0 ps=0 
M1298 diff_12680_28456# diff_16768_25436# diff_16832_28432# GND efet w=208 l=94
+ ad=0 pd=0 as=0 ps=0 
M1299 diff_17948_28768# diff_17780_29020# GND GND efet w=204 l=104
+ ad=9296 pd=528 as=0 ps=0 
M1300 diff_12680_28816# diff_17932_25436# diff_17948_28768# GND efet w=208 l=112
+ ad=0 pd=0 as=0 ps=0 
M1301 diff_15536_28288# diff_15388_25448# diff_12236_28156# GND efet w=40 l=88
+ ad=3200 pd=240 as=0 ps=0 
M1302 diff_11800_28096# diff_15148_25448# diff_15028_27832# GND efet w=40 l=82
+ ad=0 pd=0 as=2720 ps=216 
M1303 diff_15536_28144# diff_15388_25448# diff_11800_28096# GND efet w=40 l=88
+ ad=3200 pd=240 as=0 ps=0 
M1304 diff_14588_28028# diff_14420_28144# GND GND efet w=192 l=104
+ ad=11984 pd=600 as=0 ps=0 
M1305 GND diff_13912_27712# diff_13844_27692# GND efet w=186 l=110
+ ad=0 pd=0 as=11936 ps=528 
M1306 GND diff_12256_27580# diff_11800_27280# GND efet w=478 l=94
+ ad=0 pd=0 as=0 ps=0 
M1307 diff_13844_27692# diff_13744_27736# diff_12256_27580# GND efet w=202 l=94
+ ad=0 pd=0 as=0 ps=0 
M1308 diff_12256_27952# diff_14416_25448# diff_14588_28028# GND efet w=232 l=82
+ ad=0 pd=0 as=0 ps=0 
M1309 diff_14960_27844# diff_14860_29452# diff_12256_27952# GND efet w=208 l=88
+ ad=12800 pd=552 as=0 ps=0 
M1310 GND diff_15028_27832# diff_14960_27844# GND efet w=180 l=104
+ ad=0 pd=0 as=0 ps=0 
M1311 diff_17192_28580# diff_17092_28684# diff_12680_28456# GND efet w=196 l=88
+ ad=12560 pd=552 as=0 ps=0 
M1312 GND diff_17272_28288# diff_17192_28580# GND efet w=166 l=106
+ ad=0 pd=0 as=0 ps=0 
M1313 Vdd diff_17152_20864# diff_12256_29344# GND efet w=88 l=112
+ ad=0 pd=0 as=0 ps=0 
M1314 Vdd Vdd diff_11788_29092# GND efet w=64 l=268
+ ad=0 pd=0 as=0 ps=0 
M1315 Vdd Vdd diff_12236_28852# GND efet w=64 l=268
+ ad=0 pd=0 as=0 ps=0 
M1316 Vdd diff_17152_20864# diff_12680_28816# GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M1317 diff_17948_28432# diff_17780_28288# GND GND efet w=204 l=104
+ ad=9968 pd=528 as=0 ps=0 
M1318 diff_12236_28156# diff_16312_25436# diff_16144_28612# GND efet w=40 l=100
+ ad=0 pd=0 as=2864 ps=240 
M1319 diff_16652_28288# diff_16516_26800# diff_12236_28156# GND efet w=40 l=88
+ ad=3200 pd=240 as=0 ps=0 
M1320 diff_11800_28096# diff_16312_25436# diff_16144_27832# GND efet w=40 l=112
+ ad=0 pd=0 as=2720 ps=216 
M1321 diff_16652_28144# diff_16516_26800# diff_11800_28096# GND efet w=52 l=100
+ ad=3296 pd=264 as=0 ps=0 
M1322 diff_12236_27076# diff_12680_27040# GND GND efet w=508 l=88
+ ad=0 pd=0 as=0 ps=0 
M1323 diff_12680_27040# diff_12544_25804# diff_11180_26992# GND efet w=100 l=88
+ ad=139328 pd=4224 as=0 ps=0 
M1324 diff_14600_27556# diff_14420_27400# GND GND efet w=180 l=104
+ ad=12080 pd=528 as=0 ps=0 
M1325 diff_12256_27580# diff_14416_25448# diff_14600_27556# GND efet w=220 l=88
+ ad=0 pd=0 as=0 ps=0 
M1326 diff_14960_27692# diff_14860_29452# diff_12256_27580# GND efet w=196 l=88
+ ad=12080 pd=528 as=0 ps=0 
M1327 GND diff_15028_27712# diff_14960_27692# GND efet w=180 l=104
+ ad=0 pd=0 as=0 ps=0 
M1328 diff_15716_27892# diff_15536_28144# GND GND efet w=186 l=110
+ ad=11168 pd=576 as=0 ps=0 
M1329 diff_12256_27952# diff_15592_25448# diff_15716_27892# GND efet w=220 l=88
+ ad=0 pd=0 as=0 ps=0 
M1330 diff_16076_27844# diff_15976_29452# diff_12256_27952# GND efet w=208 l=88
+ ad=13328 pd=552 as=0 ps=0 
M1331 GND diff_16144_27832# diff_16076_27844# GND efet w=180 l=116
+ ad=0 pd=0 as=0 ps=0 
M1332 diff_12680_28456# diff_17932_25436# diff_17948_28432# GND efet w=208 l=112
+ ad=0 pd=0 as=0 ps=0 
M1333 diff_12236_28156# diff_17440_26356# diff_17272_28288# GND efet w=40 l=100
+ ad=0 pd=0 as=2720 ps=216 
M1334 diff_17780_28288# diff_17632_26752# diff_12236_28156# GND efet w=46 l=106
+ ad=2720 pd=216 as=0 ps=0 
M1335 diff_11800_28096# diff_17440_26356# diff_17272_27832# GND efet w=52 l=100
+ ad=0 pd=0 as=3536 ps=240 
M1336 diff_16832_27892# diff_16652_28144# GND GND efet w=180 l=110
+ ad=9968 pd=552 as=0 ps=0 
M1337 diff_12256_27952# diff_16768_25436# diff_16832_27892# GND efet w=202 l=106
+ ad=0 pd=0 as=0 ps=0 
M1338 diff_17192_27844# diff_17092_28684# diff_12256_27952# GND efet w=196 l=94
+ ad=12944 pd=552 as=0 ps=0 
M1339 GND diff_17272_27832# diff_17192_27844# GND efet w=156 l=88
+ ad=0 pd=0 as=0 ps=0 
M1340 diff_15716_27556# diff_15536_27428# GND GND efet w=180 l=116
+ ad=11792 pd=528 as=0 ps=0 
M1341 diff_11800_27280# diff_13972_25448# diff_13912_27712# GND efet w=40 l=94
+ ad=0 pd=0 as=2240 ps=240 
M1342 diff_14420_27400# diff_14224_25448# diff_11800_27280# GND efet w=46 l=94
+ ad=3392 pd=288 as=0 ps=0 
M1343 diff_12236_27076# diff_13972_25448# diff_13912_26956# GND efet w=58 l=82
+ ad=0 pd=0 as=3104 ps=264 
M1344 diff_14420_27256# diff_14224_25448# diff_12236_27076# GND efet w=40 l=88
+ ad=3200 pd=240 as=0 ps=0 
M1345 diff_13844_26968# diff_13744_27736# diff_12680_27040# GND efet w=196 l=88
+ ad=11936 pd=528 as=0 ps=0 
M1346 GND diff_13912_26956# diff_13844_26968# GND efet w=180 l=104
+ ad=0 pd=0 as=0 ps=0 
M1347 Vdd Vdd diff_5428_26392# GND efet w=44 l=240
+ ad=0 pd=0 as=0 ps=0 
M1348 Vdd diff_8680_20596# diff_6172_26164# GND efet w=82 l=88
+ ad=0 pd=0 as=0 ps=0 
M1349 diff_10996_26404# diff_2656_22088# diff_3808_28348# GND efet w=100 l=88
+ ad=10592 pd=456 as=0 ps=0 
M1350 diff_3808_28348# diff_11872_25876# diff_11800_26332# GND efet w=376 l=88
+ ad=0 pd=0 as=133904 ps=4592 
M1351 diff_12236_26380# diff_12136_25792# diff_3808_28348# GND efet w=364 l=88
+ ad=127952 pd=4536 as=0 ps=0 
M1352 diff_9392_25792# diff_9212_25636# GND GND efet w=186 l=122
+ ad=12512 pd=552 as=0 ps=0 
M1353 diff_5408_25636# diff_7576_23716# diff_7588_25948# GND efet w=40 l=88
+ ad=0 pd=0 as=3200 ps=240 
M1354 diff_8096_25636# diff_7816_23824# diff_5408_25636# GND efet w=40 l=88
+ ad=3344 pd=264 as=0 ps=0 
M1355 diff_6152_25792# diff_9232_23696# diff_9392_25792# GND efet w=202 l=88
+ ad=0 pd=0 as=0 ps=0 
M1356 diff_5408_25636# diff_8788_23696# diff_8704_25960# GND efet w=40 l=76
+ ad=0 pd=0 as=3488 ps=264 
M1357 diff_9212_25636# diff_9028_23696# diff_5408_25636# GND efet w=40 l=76
+ ad=3344 pd=264 as=0 ps=0 
M1358 diff_5396_25448# diff_7576_23716# diff_7588_25192# GND efet w=40 l=88
+ ad=0 pd=0 as=3200 ps=240 
M1359 diff_8096_25492# diff_7816_23824# diff_5396_25448# GND efet w=40 l=88
+ ad=3200 pd=240 as=0 ps=0 
M1360 diff_7508_25192# diff_7348_23696# diff_6152_25264# GND efet w=220 l=82
+ ad=13088 pd=576 as=0 ps=0 
M1361 GND diff_7588_25192# diff_7508_25192# GND efet w=186 l=98
+ ad=0 pd=0 as=0 ps=0 
M1362 diff_8264_25240# diff_8096_25492# GND GND efet w=186 l=110
+ ad=12944 pd=576 as=0 ps=0 
M1363 diff_5396_25448# diff_8788_23696# diff_8704_25192# GND efet w=40 l=76
+ ad=0 pd=0 as=3200 ps=240 
M1364 diff_9212_25492# diff_9028_23696# diff_5396_25448# GND efet w=40 l=82
+ ad=3200 pd=240 as=0 ps=0 
M1365 GND diff_6160_24964# diff_5428_24556# GND efet w=556 l=88
+ ad=0 pd=0 as=128032 ps=3904 
M1366 GND diff_7588_25072# diff_7508_25052# GND efet w=192 l=116
+ ad=0 pd=0 as=12224 ps=552 
M1367 diff_4204_24416# diff_6020_23524# diff_6160_24964# GND efet w=112 l=88
+ ad=0 pd=0 as=95408 ps=3104 
M1368 diff_3040_29500# diff_5212_23848# diff_5428_24556# GND efet w=352 l=88
+ ad=0 pd=0 as=0 ps=0 
M1369 diff_5792_24436# diff_5200_22772# diff_3040_29500# GND efet w=394 l=82
+ ad=105040 pd=3616 as=0 ps=0 
M1370 Vdd diff_2740_24880# diff_2836_23896# GND efet w=52 l=88
+ ad=0 pd=0 as=0 ps=0 
M1371 diff_4040_23804# diff_2836_23896# GND GND efet w=232 l=88
+ ad=37408 pd=1344 as=0 ps=0 
M1372 diff_7508_25052# diff_7348_23696# diff_6160_24964# GND efet w=208 l=88
+ ad=0 pd=0 as=0 ps=0 
M1373 diff_6152_25264# diff_8020_23696# diff_8264_25240# GND efet w=202 l=82
+ ad=0 pd=0 as=0 ps=0 
M1374 diff_8636_25192# diff_8548_23696# diff_6152_25264# GND efet w=208 l=88
+ ad=12560 pd=600 as=0 ps=0 
M1375 GND diff_8704_25192# diff_8636_25192# GND efet w=186 l=104
+ ad=0 pd=0 as=0 ps=0 
M1376 diff_9392_25228# diff_9212_25492# GND GND efet w=178 l=122
+ ad=12368 pd=528 as=0 ps=0 
M1377 diff_8276_24904# diff_8096_24748# GND GND efet w=168 l=116
+ ad=11840 pd=528 as=0 ps=0 
M1378 diff_6160_24964# diff_8020_23696# diff_8276_24904# GND efet w=202 l=82
+ ad=0 pd=0 as=0 ps=0 
M1379 GND diff_6584_24388# diff_5792_24436# GND efet w=562 l=106
+ ad=0 pd=0 as=0 ps=0 
M1380 diff_6584_24388# diff_6496_23704# diff_4204_24416# GND efet w=100 l=88
+ ad=92752 pd=3024 as=0 ps=0 
M1381 Vdd Vdd diff_4040_23804# GND efet w=52 l=532
+ ad=0 pd=0 as=0 ps=0 
M1382 GND diff_1132_21544# diff_3508_23020# GND efet w=196 l=88
+ ad=0 pd=0 as=47072 ps=1352 
M1383 diff_4040_23804# clk2 diff_3952_23632# GND efet w=96 l=116
+ ad=0 pd=0 as=5600 ps=392 
M1384 cm_rom diff_928_16456# Vdd GND efet w=3448 l=88
+ ad=399536 pd=10240 as=0 ps=0 
M1385 GND diff_1232_22576# cm_rom GND efet w=5020 l=82
+ ad=0 pd=0 as=0 ps=0 
M1386 GND diff_2140_5752# diff_3508_23020# GND efet w=214 l=94
+ ad=0 pd=0 as=0 ps=0 
M1387 diff_2740_24880# Vdd clk1 GND efet w=280 l=88
+ ad=21888 pd=776 as=1.10218e+06 ps=23528 
M1388 Vdd Vdd diff_6020_23524# GND efet w=40 l=220
+ ad=0 pd=0 as=38640 ps=1600 
M1389 GND diff_2140_4552# diff_3200_23188# GND efet w=100 l=94
+ ad=0 pd=0 as=45792 ps=1704 
M1390 diff_4052_23284# diff_3952_23632# GND GND efet w=160 l=88
+ ad=36016 pd=1024 as=0 ps=0 
M1391 diff_5144_23548# Vdd Vdd GND efet w=52 l=220
+ ad=64896 pd=2416 as=0 ps=0 
M1392 GND diff_4436_22444# diff_5144_23548# GND efet w=228 l=104
+ ad=0 pd=0 as=0 ps=0 
M1393 Vdd Vdd diff_4052_23284# GND efet w=46 l=418
+ ad=0 pd=0 as=0 ps=0 
M1394 diff_3200_23188# Vdd Vdd GND efet w=46 l=550
+ ad=0 pd=0 as=0 ps=0 
M1395 diff_4052_23284# clk1 diff_3952_23104# GND efet w=64 l=88
+ ad=0 pd=0 as=13280 ps=632 
M1396 diff_1232_22576# Vdd Vdd GND efet w=70 l=106
+ ad=63056 pd=2280 as=0 ps=0 
M1397 GND diff_3856_18340# diff_5144_23548# GND efet w=292 l=88
+ ad=0 pd=0 as=0 ps=0 
M1398 diff_8636_25028# diff_8548_23696# diff_6160_24964# GND efet w=196 l=88
+ ad=11696 pd=552 as=0 ps=0 
M1399 GND diff_8704_25072# diff_8636_25028# GND efet w=180 l=116
+ ad=0 pd=0 as=0 ps=0 
M1400 diff_6152_25264# diff_9232_23696# diff_9392_25228# GND efet w=196 l=88
+ ad=0 pd=0 as=0 ps=0 
M1401 Vdd diff_8680_20596# diff_6152_25792# GND efet w=64 l=100
+ ad=0 pd=0 as=0 ps=0 
M1402 diff_12680_26680# diff_12544_25804# diff_11180_26776# GND efet w=100 l=88
+ ad=135392 pd=4152 as=0 ps=0 
M1403 diff_12256_27580# diff_15592_25448# diff_15716_27556# GND efet w=196 l=88
+ ad=0 pd=0 as=0 ps=0 
M1404 diff_16076_27692# diff_15976_29452# diff_12256_27580# GND efet w=196 l=88
+ ad=12224 pd=528 as=0 ps=0 
M1405 GND diff_16144_27724# diff_16076_27692# GND efet w=186 l=134
+ ad=0 pd=0 as=0 ps=0 
M1406 diff_17780_28132# diff_17632_26752# diff_11800_28096# GND efet w=58 l=118
+ ad=3680 pd=264 as=0 ps=0 
M1407 diff_17948_27880# diff_17780_28132# GND GND efet w=216 l=116
+ ad=9440 pd=528 as=0 ps=0 
M1408 diff_16832_27556# diff_16664_27400# GND GND efet w=180 l=116
+ ad=11120 pd=528 as=0 ps=0 
M1409 diff_11800_27280# diff_15148_25448# diff_15028_27712# GND efet w=40 l=100
+ ad=0 pd=0 as=2864 ps=240 
M1410 diff_15536_27428# diff_15388_25448# diff_11800_27280# GND efet w=48 l=82
+ ad=2864 pd=240 as=0 ps=0 
M1411 diff_12236_27076# diff_15148_25448# diff_15040_26944# GND efet w=40 l=88
+ ad=0 pd=0 as=3200 ps=240 
M1412 diff_15548_27256# diff_15388_25448# diff_12236_27076# GND efet w=40 l=88
+ ad=2864 pd=240 as=0 ps=0 
M1413 GND diff_13912_26836# diff_13844_26816# GND efet w=186 l=110
+ ad=0 pd=0 as=11792 ps=528 
M1414 diff_11180_26776# diff_12328_25804# diff_12256_26224# GND efet w=118 l=76
+ ad=0 pd=0 as=142704 ps=4400 
M1415 GND diff_12680_26680# diff_12236_26380# GND efet w=484 l=88
+ ad=0 pd=0 as=0 ps=0 
M1416 diff_13844_26816# diff_13744_27736# diff_12680_26680# GND efet w=196 l=88
+ ad=0 pd=0 as=0 ps=0 
M1417 diff_14600_27004# diff_14420_27256# GND GND efet w=186 l=110
+ ad=12080 pd=528 as=0 ps=0 
M1418 diff_12680_27040# diff_14416_25448# diff_14600_27004# GND efet w=196 l=88
+ ad=0 pd=0 as=0 ps=0 
M1419 diff_14960_26968# diff_14860_29452# diff_12680_27040# GND efet w=196 l=100
+ ad=12848 pd=576 as=0 ps=0 
M1420 GND diff_15040_26944# diff_14960_26968# GND efet w=198 l=98
+ ad=0 pd=0 as=0 ps=0 
M1421 diff_14600_26668# diff_14420_26524# GND GND efet w=180 l=104
+ ad=12368 pd=528 as=0 ps=0 
M1422 diff_12256_27580# diff_16768_25436# diff_16832_27556# GND efet w=202 l=94
+ ad=0 pd=0 as=0 ps=0 
M1423 diff_17192_27692# diff_17092_28684# diff_12256_27580# GND efet w=220 l=88
+ ad=13040 pd=576 as=0 ps=0 
M1424 GND diff_17272_27400# diff_17192_27692# GND efet w=160 l=88
+ ad=0 pd=0 as=0 ps=0 
M1425 diff_11800_27280# diff_16312_25436# diff_16144_27724# GND efet w=40 l=88
+ ad=0 pd=0 as=3200 ps=240 
M1426 diff_16664_27400# diff_16516_26800# diff_11800_27280# GND efet w=46 l=100
+ ad=2720 pd=216 as=0 ps=0 
M1427 diff_12256_27952# diff_17932_25436# diff_17948_27880# GND efet w=202 l=94
+ ad=0 pd=0 as=0 ps=0 
M1428 diff_17948_27544# diff_17780_27400# GND GND efet w=216 l=116
+ ad=10160 pd=552 as=0 ps=0 
M1429 Vdd diff_17152_20864# diff_12680_28456# GND efet w=88 l=108
+ ad=0 pd=0 as=0 ps=0 
M1430 Vdd Vdd diff_12236_28156# GND efet w=52 l=304
+ ad=0 pd=0 as=0 ps=0 
M1431 Vdd Vdd diff_11800_28096# GND efet w=58 l=286
+ ad=0 pd=0 as=0 ps=0 
M1432 Vdd diff_17152_20864# diff_12256_27952# GND efet w=94 l=106
+ ad=0 pd=0 as=0 ps=0 
M1433 diff_12256_27580# diff_17932_25436# diff_17948_27544# GND efet w=208 l=94
+ ad=0 pd=0 as=0 ps=0 
M1434 diff_12236_27076# diff_16312_25436# diff_16144_26956# GND efet w=40 l=88
+ ad=0 pd=0 as=3200 ps=240 
M1435 diff_11800_26332# diff_12256_26224# GND GND efet w=484 l=88
+ ad=0 pd=0 as=0 ps=0 
M1436 diff_12680_26680# diff_14416_25448# diff_14600_26668# GND efet w=196 l=88
+ ad=0 pd=0 as=0 ps=0 
M1437 diff_14960_26816# diff_14860_29452# diff_12680_26680# GND efet w=196 l=88
+ ad=12320 pd=552 as=0 ps=0 
M1438 GND diff_15028_26836# diff_14960_26816# GND efet w=210 l=104
+ ad=0 pd=0 as=0 ps=0 
M1439 diff_15716_27004# diff_15548_27256# GND GND efet w=186 l=122
+ ad=12512 pd=576 as=0 ps=0 
M1440 diff_12680_27040# diff_15592_25448# diff_15716_27004# GND efet w=226 l=82
+ ad=0 pd=0 as=0 ps=0 
M1441 diff_16076_26956# diff_15976_29452# diff_12680_27040# GND efet w=238 l=82
+ ad=13136 pd=624 as=0 ps=0 
M1442 GND diff_16144_26956# diff_16076_26956# GND efet w=198 l=110
+ ad=0 pd=0 as=0 ps=0 
M1443 diff_16664_27256# diff_16516_26800# diff_12236_27076# GND efet w=40 l=88
+ ad=2864 pd=240 as=0 ps=0 
M1444 diff_11800_27280# diff_17440_26356# diff_17272_27400# GND efet w=40 l=94
+ ad=0 pd=0 as=2720 ps=216 
M1445 diff_17780_27400# diff_17632_26752# diff_11800_27280# GND efet w=46 l=106
+ ad=2720 pd=216 as=0 ps=0 
M1446 diff_12236_27076# diff_17440_26356# diff_17272_26944# GND efet w=46 l=106
+ ad=0 pd=0 as=3008 ps=240 
M1447 diff_17780_27256# diff_17632_26752# diff_12236_27076# GND efet w=46 l=118
+ ad=2864 pd=240 as=0 ps=0 
M1448 diff_16832_27004# diff_16664_27256# GND GND efet w=192 l=104
+ ad=11648 pd=552 as=0 ps=0 
M1449 diff_12680_27040# diff_16768_25436# diff_16832_27004# GND efet w=214 l=94
+ ad=0 pd=0 as=0 ps=0 
M1450 diff_17192_26956# diff_17092_28684# diff_12680_27040# GND efet w=232 l=88
+ ad=11840 pd=576 as=0 ps=0 
M1451 diff_15716_26668# diff_15548_26512# GND GND efet w=180 l=110
+ ad=12320 pd=552 as=0 ps=0 
M1452 diff_12236_26380# diff_13972_25448# diff_13912_26836# GND efet w=46 l=106
+ ad=0 pd=0 as=3248 ps=312 
M1453 diff_14420_26524# diff_14224_25448# diff_12236_26380# GND efet w=28 l=94
+ ad=2240 pd=216 as=0 ps=0 
M1454 diff_11800_26332# diff_13972_25448# diff_13912_26068# GND efet w=52 l=88
+ ad=0 pd=0 as=3008 ps=264 
M1455 diff_14420_26368# diff_14224_25448# diff_11800_26332# GND efet w=40 l=88
+ ad=3200 pd=240 as=0 ps=0 
M1456 diff_13844_26080# diff_13744_27736# diff_12256_26224# GND efet w=196 l=106
+ ad=11792 pd=528 as=0 ps=0 
M1457 GND diff_13912_26068# diff_13844_26080# GND efet w=180 l=104
+ ad=0 pd=0 as=0 ps=0 
M1458 diff_12680_26680# diff_15592_25448# diff_15716_26668# GND efet w=214 l=88
+ ad=0 pd=0 as=0 ps=0 
M1459 diff_16076_26804# diff_15976_29452# diff_12680_26680# GND efet w=214 l=94
+ ad=11504 pd=576 as=0 ps=0 
M1460 GND diff_16156_26512# diff_16076_26804# GND efet w=204 l=128
+ ad=0 pd=0 as=0 ps=0 
M1461 GND diff_17272_26944# diff_17192_26956# GND efet w=166 l=118
+ ad=0 pd=0 as=0 ps=0 
M1462 diff_16832_26656# diff_16664_26512# GND GND efet w=192 l=116
+ ad=11936 pd=552 as=0 ps=0 
M1463 diff_12236_26380# diff_15148_25448# diff_15028_26836# GND efet w=52 l=88
+ ad=0 pd=0 as=3920 ps=264 
M1464 diff_15548_26512# diff_15388_25448# diff_12236_26380# GND efet w=46 l=106
+ ad=2864 pd=240 as=0 ps=0 
M1465 diff_11800_26332# diff_15148_25448# diff_15040_26056# GND efet w=40 l=88
+ ad=0 pd=0 as=3200 ps=240 
M1466 diff_15548_26368# diff_15388_25448# diff_11800_26332# GND efet w=40 l=88
+ ad=2864 pd=240 as=0 ps=0 
M1467 Vdd Vdd diff_5408_25636# GND efet w=40 l=244
+ ad=0 pd=0 as=0 ps=0 
M1468 GND diff_11224_25648# diff_10976_25588# GND efet w=100 l=100
+ ad=0 pd=0 as=36544 ps=1456 
M1469 diff_10976_25588# Vdd Vdd GND efet w=64 l=532
+ ad=0 pd=0 as=0 ps=0 
M1470 diff_11224_25648# diff_10976_25588# GND GND efet w=88 l=88
+ ad=42656 pd=1520 as=0 ps=0 
M1471 diff_14600_26116# diff_14420_26368# GND GND efet w=186 l=110
+ ad=12896 pd=576 as=0 ps=0 
M1472 diff_12256_26224# diff_14416_25448# diff_14600_26116# GND efet w=220 l=88
+ ad=0 pd=0 as=0 ps=0 
M1473 diff_14960_26068# diff_14860_29452# diff_12256_26224# GND efet w=220 l=100
+ ad=13376 pd=576 as=0 ps=0 
M1474 GND diff_15040_26056# diff_14960_26068# GND efet w=216 l=104
+ ad=0 pd=0 as=0 ps=0 
M1475 diff_12680_26680# diff_16768_25436# diff_16832_26656# GND efet w=208 l=100
+ ad=0 pd=0 as=0 ps=0 
M1476 diff_17192_26816# diff_17092_28684# diff_12680_26680# GND efet w=250 l=106
+ ad=11552 pd=552 as=0 ps=0 
M1477 GND diff_17260_26836# diff_17192_26816# GND efet w=178 l=140
+ ad=0 pd=0 as=0 ps=0 
M1478 diff_17948_26996# diff_17780_27256# GND GND efet w=234 l=122
+ ad=9728 pd=576 as=0 ps=0 
M1479 diff_12680_27040# diff_17932_25436# diff_17948_26996# GND efet w=220 l=100
+ ad=0 pd=0 as=0 ps=0 
M1480 Vdd diff_17152_20864# diff_12256_27580# GND efet w=112 l=112
+ ad=0 pd=0 as=0 ps=0 
M1481 Vdd Vdd diff_11800_27280# GND efet w=64 l=278
+ ad=0 pd=0 as=0 ps=0 
M1482 Vdd Vdd diff_12236_27076# GND efet w=58 l=262
+ ad=0 pd=0 as=0 ps=0 
M1483 Vdd diff_17152_20864# diff_12680_27040# GND efet w=88 l=100
+ ad=0 pd=0 as=0 ps=0 
M1484 diff_17948_26656# diff_17780_26512# GND GND efet w=228 l=100
+ ad=11792 pd=624 as=0 ps=0 
M1485 diff_12680_26680# diff_17932_25436# diff_17948_26656# GND efet w=232 l=88
+ ad=0 pd=0 as=0 ps=0 
M1486 diff_16664_26512# diff_16516_26800# diff_12236_26380# GND efet w=40 l=106
+ ad=2720 pd=216 as=0 ps=0 
M1487 diff_12236_26380# diff_16312_25436# diff_16156_26512# GND efet w=40 l=88
+ ad=0 pd=0 as=3152 ps=240 
M1488 diff_11800_26332# diff_16312_25436# diff_16156_26056# GND efet w=40 l=88
+ ad=0 pd=0 as=3152 ps=240 
M1489 diff_15716_26116# diff_15548_26368# GND GND efet w=186 l=110
+ ad=12944 pd=576 as=0 ps=0 
M1490 diff_12256_26224# diff_15592_25448# diff_15716_26116# GND efet w=220 l=88
+ ad=0 pd=0 as=0 ps=0 
M1491 diff_16076_26068# diff_15976_29452# diff_12256_26224# GND efet w=220 l=88
+ ad=12992 pd=600 as=0 ps=0 
M1492 GND diff_16156_26056# diff_16076_26068# GND efet w=198 l=110
+ ad=0 pd=0 as=0 ps=0 
M1493 diff_16664_26368# diff_16516_26800# diff_11800_26332# GND efet w=40 l=88
+ ad=2864 pd=240 as=0 ps=0 
M1494 diff_16832_26180# diff_16664_26368# GND GND efet w=214 l=116
+ ad=10976 pd=592 as=0 ps=0 
M1495 Vdd diff_17152_20864# diff_12680_26680# GND efet w=88 l=100
+ ad=0 pd=0 as=0 ps=0 
M1496 diff_12236_26380# diff_17440_26356# diff_17260_26836# GND efet w=40 l=88
+ ad=0 pd=0 as=2864 ps=240 
M1497 diff_17780_26512# diff_17632_26752# diff_12236_26380# GND efet w=40 l=100
+ ad=2720 pd=216 as=0 ps=0 
M1498 diff_11800_26332# diff_17440_26356# diff_17272_26056# GND efet w=40 l=100
+ ad=0 pd=0 as=3056 ps=264 
M1499 diff_17780_26356# diff_17632_26752# diff_11800_26332# GND efet w=52 l=112
+ ad=3440 pd=264 as=0 ps=0 
M1500 diff_12256_26224# diff_16768_25436# diff_16832_26180# GND efet w=208 l=94
+ ad=0 pd=0 as=0 ps=0 
M1501 diff_17204_26068# diff_17092_28684# diff_12256_26224# GND efet w=208 l=100
+ ad=11936 pd=576 as=0 ps=0 
M1502 GND diff_17272_26056# diff_17204_26068# GND efet w=216 l=128
+ ad=0 pd=0 as=0 ps=0 
M1503 Vdd Vdd diff_12236_26380# GND efet w=64 l=274
+ ad=0 pd=0 as=0 ps=0 
M1504 GND GND clk2 GND efet w=970 l=106
+ ad=0 pd=0 as=1.11096e+06 ps=19008 
M1505 GND GND clk1 GND efet w=928 l=100
+ ad=0 pd=0 as=0 ps=0 
M1506 Vdd Vdd diff_11800_26332# GND efet w=60 l=274
+ ad=0 pd=0 as=0 ps=0 
M1507 diff_17948_26108# diff_17780_26356# GND GND efet w=204 l=128
+ ad=10400 pd=528 as=0 ps=0 
M1508 diff_12256_26224# diff_17932_25436# diff_17948_26108# GND efet w=214 l=94
+ ad=0 pd=0 as=0 ps=0 
M1509 Vdd diff_17152_20864# diff_12256_26224# GND efet w=88 l=112
+ ad=0 pd=0 as=0 ps=0 
M1510 Vdd Vdd diff_5396_25448# GND efet w=40 l=232
+ ad=0 pd=0 as=0 ps=0 
M1511 Vdd Vdd diff_11224_25648# GND efet w=40 l=532
+ ad=0 pd=0 as=0 ps=0 
M1512 diff_9412_21772# Vdd Vdd GND efet w=64 l=544
+ ad=103616 pd=4024 as=0 ps=0 
M1513 GND diff_11224_25648# diff_9412_21772# GND efet w=118 l=82
+ ad=0 pd=0 as=0 ps=0 
M1514 diff_11708_25456# diff_10976_25588# GND GND efet w=112 l=88
+ ad=33040 pd=1360 as=0 ps=0 
M1515 GND diff_13484_25336# diff_13744_27736# GND efet w=112 l=88
+ ad=0 pd=0 as=15680 ps=504 
M1516 GND diff_13484_25336# diff_13972_25448# GND efet w=88 l=88
+ ad=0 pd=0 as=12320 ps=456 
M1517 GND diff_14164_25600# diff_14224_25448# GND efet w=88 l=88
+ ad=0 pd=0 as=12320 ps=456 
M1518 GND diff_14164_25600# diff_14416_25448# GND efet w=112 l=88
+ ad=0 pd=0 as=15680 ps=504 
M1519 Vdd Vdd diff_11708_25456# GND efet w=70 l=538
+ ad=0 pd=0 as=0 ps=0 
M1520 Vdd diff_8680_20596# diff_6152_25264# GND efet w=70 l=82
+ ad=0 pd=0 as=0 ps=0 
M1521 diff_9392_24904# diff_9212_24748# GND GND efet w=174 l=146
+ ad=11840 pd=528 as=0 ps=0 
M1522 diff_5428_24556# diff_7576_23716# diff_7588_25072# GND efet w=46 l=106
+ ad=0 pd=0 as=3248 ps=264 
M1523 diff_8096_24748# diff_7816_23824# diff_5428_24556# GND efet w=46 l=94
+ ad=3200 pd=240 as=0 ps=0 
M1524 diff_5792_24436# diff_7576_23716# diff_7588_24304# GND efet w=40 l=88
+ ad=0 pd=0 as=3200 ps=240 
M1525 diff_8096_24604# diff_7816_23824# diff_5792_24436# GND efet w=40 l=88
+ ad=3200 pd=240 as=0 ps=0 
M1526 diff_7508_24316# diff_7348_23696# diff_6584_24388# GND efet w=220 l=100
+ ad=12224 pd=552 as=0 ps=0 
M1527 GND diff_7588_24304# diff_7508_24316# GND efet w=186 l=98
+ ad=0 pd=0 as=0 ps=0 
M1528 diff_13484_25336# Vdd Vdd GND efet w=46 l=502
+ ad=41536 pd=1848 as=0 ps=0 
M1529 diff_13744_27736# diff_13708_25372# diff_13720_25264# GND efet w=130 l=82
+ ad=0 pd=0 as=302800 ps=9360 
M1530 diff_13972_25448# diff_13708_25372# diff_13972_25108# GND efet w=106 l=100
+ ad=0 pd=0 as=414288 ps=11072 
M1531 diff_14224_25448# diff_14164_25384# diff_13972_25108# GND efet w=94 l=82
+ ad=0 pd=0 as=0 ps=0 
M1532 diff_14416_25448# diff_14164_25384# diff_13720_25264# GND efet w=130 l=94
+ ad=0 pd=0 as=0 ps=0 
M1533 diff_9412_21772# diff_11020_25156# diff_11068_25000# GND efet w=64 l=76
+ ad=0 pd=0 as=4784 ps=288 
M1534 diff_11708_25456# diff_11020_25156# diff_11512_24664# GND efet w=64 l=100
+ ad=0 pd=0 as=5120 ps=288 
M1535 diff_6160_24964# diff_9232_23696# diff_9392_24904# GND efet w=196 l=88
+ ad=0 pd=0 as=0 ps=0 
M1536 diff_5428_24556# diff_8788_23696# diff_8704_25072# GND efet w=46 l=82
+ ad=0 pd=0 as=3536 ps=288 
M1537 diff_9212_24748# diff_9028_23696# diff_5428_24556# GND efet w=40 l=76
+ ad=3200 pd=240 as=0 ps=0 
M1538 diff_5792_24436# diff_8788_23696# diff_8704_24304# GND efet w=40 l=76
+ ad=0 pd=0 as=3200 ps=240 
M1539 diff_9212_24604# diff_9028_23696# diff_5792_24436# GND efet w=40 l=76
+ ad=3200 pd=240 as=0 ps=0 
M1540 diff_8264_24380# diff_8096_24604# GND GND efet w=204 l=104
+ ad=13568 pd=624 as=0 ps=0 
M1541 diff_6584_24388# diff_8020_23696# diff_8264_24380# GND efet w=220 l=100
+ ad=0 pd=0 as=0 ps=0 
M1542 diff_8636_24304# diff_8548_23696# diff_6584_24388# GND efet w=202 l=94
+ ad=12608 pd=600 as=0 ps=0 
M1543 diff_6496_23704# Vdd Vdd GND efet w=58 l=250
+ ad=59184 pd=1512 as=0 ps=0 
M1544 GND diff_8704_24304# diff_8636_24304# GND efet w=198 l=104
+ ad=0 pd=0 as=0 ps=0 
M1545 diff_9392_24340# diff_9212_24604# GND GND efet w=186 l=122
+ ad=12656 pd=552 as=0 ps=0 
M1546 diff_6584_24388# diff_9232_23696# diff_9392_24340# GND efet w=214 l=106
+ ad=0 pd=0 as=0 ps=0 
M1547 Vdd diff_8680_20596# diff_6160_24964# GND efet w=64 l=88
+ ad=0 pd=0 as=0 ps=0 
M1548 diff_11216_24704# diff_11000_24316# diff_10976_25588# GND efet w=172 l=94
+ ad=16400 pd=672 as=0 ps=0 
M1549 Vdd Vdd diff_5428_24556# GND efet w=46 l=262
+ ad=0 pd=0 as=0 ps=0 
M1550 GND diff_11068_25000# diff_11216_24704# GND efet w=274 l=88
+ ad=0 pd=0 as=0 ps=0 
M1551 diff_11600_24700# diff_11512_24664# GND GND efet w=280 l=88
+ ad=16496 pd=696 as=0 ps=0 
M1552 diff_11224_25648# diff_11000_24316# diff_11600_24700# GND efet w=160 l=88
+ ad=0 pd=0 as=0 ps=0 
M1553 Vdd Vdd diff_5792_24436# GND efet w=46 l=250
+ ad=0 pd=0 as=0 ps=0 
M1554 GND diff_14752_24940# diff_14860_29452# GND efet w=112 l=76
+ ad=0 pd=0 as=15680 ps=504 
M1555 GND diff_14752_24940# diff_15148_25448# GND efet w=88 l=76
+ ad=0 pd=0 as=12320 ps=456 
M1556 GND diff_15328_25624# diff_15388_25448# GND efet w=100 l=76
+ ad=0 pd=0 as=14000 ps=480 
M1557 GND diff_15328_25624# diff_15592_25448# GND efet w=124 l=76
+ ad=0 pd=0 as=15632 ps=528 
M1558 GND diff_15928_24928# diff_15976_29452# GND efet w=106 l=82
+ ad=0 pd=0 as=13184 ps=504 
M1559 diff_14860_29452# diff_14740_23060# diff_13720_25264# GND efet w=112 l=88
+ ad=0 pd=0 as=0 ps=0 
M1560 diff_15148_25448# diff_14740_23060# diff_13972_25108# GND efet w=94 l=94
+ ad=0 pd=0 as=0 ps=0 
M1561 diff_15388_25448# diff_15124_23692# diff_13972_25108# GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M1562 diff_15592_25448# diff_15124_23692# diff_13720_25264# GND efet w=112 l=100
+ ad=0 pd=0 as=0 ps=0 
M1563 GND diff_13708_25372# diff_13484_25336# GND efet w=88 l=100
+ ad=0 pd=0 as=0 ps=0 
M1564 diff_14164_25600# diff_14164_25384# GND GND efet w=76 l=88
+ ad=27088 pd=1008 as=0 ps=0 
M1565 diff_11872_25876# diff_12848_24544# diff_11872_25876# GND efet w=630 l=50
+ ad=230448 pd=8792 as=0 ps=0 
M1566 diff_11872_25876# diff_12848_24544# Vdd GND efet w=76 l=184
+ ad=0 pd=0 as=0 ps=0 
M1567 diff_12848_24544# Vdd Vdd GND efet w=46 l=106
+ ad=2240 pd=192 as=0 ps=0 
M1568 Vdd diff_8680_20596# diff_6584_24388# GND efet w=76 l=88
+ ad=0 pd=0 as=0 ps=0 
M1569 diff_11000_24316# Vdd Vdd GND efet w=46 l=586
+ ad=43184 pd=1376 as=0 ps=0 
M1570 GND diff_11020_25156# diff_11000_24316# GND efet w=88 l=88
+ ad=0 pd=0 as=0 ps=0 
M1571 diff_11020_25156# diff_11000_24316# GND GND efet w=100 l=88
+ ad=43696 pd=1568 as=0 ps=0 
M1572 GND diff_14740_23060# diff_14752_24940# GND efet w=82 l=94
+ ad=0 pd=0 as=28288 ps=1008 
M1573 diff_15328_25624# diff_15124_23692# GND GND efet w=76 l=100
+ ad=26224 pd=936 as=0 ps=0 
M1574 GND diff_15928_24928# diff_16312_25436# GND efet w=100 l=82
+ ad=0 pd=0 as=14000 ps=480 
M1575 GND diff_16504_25588# diff_16516_26800# GND efet w=88 l=88
+ ad=0 pd=0 as=12320 ps=456 
M1576 GND diff_16504_25588# diff_16768_25436# GND efet w=100 l=94
+ ad=0 pd=0 as=14000 ps=480 
M1577 diff_15976_29452# diff_15676_23048# diff_13720_25264# GND efet w=112 l=82
+ ad=0 pd=0 as=0 ps=0 
M1578 diff_13972_25108# diff_15676_23048# diff_16312_25436# GND efet w=94 l=82
+ ad=0 pd=0 as=0 ps=0 
M1579 diff_16516_26800# diff_16120_23288# diff_13972_25108# GND efet w=94 l=82
+ ad=0 pd=0 as=0 ps=0 
M1580 diff_16768_25436# diff_16120_23288# diff_13720_25264# GND efet w=100 l=76
+ ad=0 pd=0 as=0 ps=0 
M1581 GND diff_15676_23048# diff_15928_24928# GND efet w=94 l=94
+ ad=0 pd=0 as=28048 ps=1008 
M1582 diff_14164_25600# Vdd Vdd GND efet w=46 l=370
+ ad=0 pd=0 as=0 ps=0 
M1583 Vdd Vdd diff_14752_24940# GND efet w=54 l=418
+ ad=0 pd=0 as=0 ps=0 
M1584 diff_16504_25588# diff_16120_23288# GND GND efet w=88 l=100
+ ad=26752 pd=984 as=0 ps=0 
M1585 GND diff_17092_24928# diff_17092_28684# GND efet w=112 l=88
+ ad=0 pd=0 as=15680 ps=504 
M1586 GND diff_17092_24928# diff_17440_26356# GND efet w=88 l=88
+ ad=0 pd=0 as=12320 ps=456 
M1587 GND diff_17668_25588# diff_17632_26752# GND efet w=88 l=88
+ ad=0 pd=0 as=12320 ps=456 
M1588 GND diff_17668_25588# diff_17932_25436# GND efet w=112 l=88
+ ad=0 pd=0 as=15152 ps=528 
M1589 diff_17092_28684# diff_16636_23048# diff_13720_25264# GND efet w=118 l=82
+ ad=0 pd=0 as=0 ps=0 
M1590 diff_17440_26356# diff_16636_23048# diff_13972_25108# GND efet w=94 l=82
+ ad=0 pd=0 as=0 ps=0 
M1591 diff_17632_26752# diff_17068_23276# diff_13972_25108# GND efet w=94 l=82
+ ad=0 pd=0 as=0 ps=0 
M1592 diff_17932_25436# diff_17068_23276# diff_13720_25264# GND efet w=112 l=88
+ ad=0 pd=0 as=0 ps=0 
M1593 diff_15328_25624# Vdd Vdd GND efet w=40 l=388
+ ad=0 pd=0 as=0 ps=0 
M1594 Vdd Vdd diff_15928_24928# GND efet w=46 l=430
+ ad=0 pd=0 as=0 ps=0 
M1595 GND diff_16636_23048# diff_17092_24928# GND efet w=76 l=100
+ ad=0 pd=0 as=26368 ps=936 
M1596 diff_17668_25588# diff_17068_23276# GND GND efet w=76 l=100
+ ad=25264 pd=960 as=0 ps=0 
M1597 Vdd Vdd diff_15472_24352# GND efet w=100 l=370
+ ad=0 pd=0 as=70336 ps=2432 
M1598 diff_16504_25588# Vdd Vdd GND efet w=46 l=394
+ ad=0 pd=0 as=0 ps=0 
M1599 Vdd Vdd diff_17092_24928# GND efet w=40 l=388
+ ad=0 pd=0 as=0 ps=0 
M1600 diff_17668_25588# Vdd Vdd GND efet w=40 l=388
+ ad=0 pd=0 as=0 ps=0 
M1601 GND diff_13816_24448# diff_13792_23696# GND efet w=220 l=100
+ ad=0 pd=0 as=99296 ps=2640 
M1602 Vdd Vdd diff_13816_24448# GND efet w=52 l=232
+ ad=0 pd=0 as=31504 ps=1296 
M1603 Vdd Vdd diff_11020_25156# GND efet w=46 l=562
+ ad=0 pd=0 as=0 ps=0 
M1604 diff_12848_24340# Vdd Vdd GND efet w=46 l=102
+ ad=2576 pd=264 as=0 ps=0 
M1605 diff_9412_21556# Vdd Vdd GND efet w=70 l=604
+ ad=100352 pd=3976 as=0 ps=0 
M1606 GND diff_11020_25156# diff_9412_21556# GND efet w=106 l=82
+ ad=0 pd=0 as=0 ps=0 
M1607 diff_11708_24184# diff_11000_24316# GND GND efet w=100 l=88
+ ad=32368 pd=1336 as=0 ps=0 
M1608 diff_12136_25792# diff_12848_24340# diff_12136_25792# GND efet w=466 l=122
+ ad=322432 pd=9928 as=0 ps=0 
M1609 Vdd Vdd diff_11708_24184# GND efet w=64 l=544
+ ad=0 pd=0 as=0 ps=0 
M1610 diff_12136_25792# diff_12848_24340# Vdd GND efet w=52 l=172
+ ad=0 pd=0 as=0 ps=0 
M1611 diff_6020_23524# diff_4700_19432# GND GND efet w=220 l=88
+ ad=0 pd=0 as=0 ps=0 
M1612 GND diff_4156_19880# diff_6496_23704# GND efet w=232 l=100
+ ad=0 pd=0 as=0 ps=0 
M1613 GND diff_4436_22444# diff_6020_23524# GND efet w=216 l=98
+ ad=0 pd=0 as=0 ps=0 
M1614 diff_6496_23704# diff_4436_22444# GND GND efet w=234 l=82
+ ad=0 pd=0 as=0 ps=0 
M1615 GND diff_7180_23308# diff_7348_23696# GND efet w=124 l=76
+ ad=0 pd=0 as=17360 ps=528 
M1616 GND diff_7180_23308# diff_7576_23716# GND efet w=88 l=76
+ ad=0 pd=0 as=12080 ps=456 
M1617 GND diff_7768_23848# diff_7816_23824# GND efet w=88 l=88
+ ad=0 pd=0 as=12368 ps=480 
M1618 GND diff_7768_23848# diff_8020_23696# GND efet w=124 l=76
+ ad=0 pd=0 as=17360 ps=528 
M1619 diff_7348_23696# diff_7288_23632# diff_6400_21080# GND efet w=124 l=88
+ ad=0 pd=0 as=142928 ps=4264 
M1620 diff_7576_23716# diff_7288_23632# diff_6952_20728# GND efet w=76 l=88
+ ad=0 pd=0 as=193008 ps=5184 
M1621 diff_7816_23824# diff_7768_23620# diff_6952_20728# GND efet w=94 l=94
+ ad=0 pd=0 as=0 ps=0 
M1622 diff_8020_23696# diff_7768_23620# diff_6400_21080# GND efet w=124 l=88
+ ad=0 pd=0 as=0 ps=0 
M1623 diff_3200_23188# diff_3460_23104# diff_3508_23020# GND efet w=184 l=76
+ ad=0 pd=0 as=0 ps=0 
M1624 GND diff_8380_23308# diff_8548_23696# GND efet w=124 l=76
+ ad=0 pd=0 as=17360 ps=528 
M1625 GND diff_8380_23308# diff_8788_23696# GND efet w=88 l=88
+ ad=0 pd=0 as=10784 ps=456 
M1626 GND diff_8968_23872# diff_9028_23696# GND efet w=88 l=88
+ ad=0 pd=0 as=11264 ps=432 
M1627 diff_9232_23696# diff_8968_23872# GND GND efet w=124 l=100
+ ad=14528 pd=528 as=0 ps=0 
M1628 diff_9412_21556# clk1 diff_11068_23716# GND efet w=52 l=88
+ ad=0 pd=0 as=3680 ps=264 
M1629 diff_14164_25384# diff_13816_24448# GND GND efet w=112 l=76
+ ad=88608 pd=3992 as=0 ps=0 
M1630 diff_14740_23060# diff_13816_24448# GND GND efet w=112 l=88
+ ad=85728 pd=2896 as=0 ps=0 
M1631 diff_15124_23692# diff_13816_24448# GND GND efet w=106 l=112
+ ad=85152 pd=3072 as=0 ps=0 
M1632 diff_15676_23048# diff_15472_24352# GND GND efet w=106 l=106
+ ad=88560 pd=3024 as=0 ps=0 
M1633 diff_13816_24448# diff_15472_24352# GND GND efet w=262 l=82
+ ad=0 pd=0 as=0 ps=0 
M1634 diff_16120_23288# diff_15472_24352# GND GND efet w=118 l=94
+ ad=84048 pd=2992 as=0 ps=0 
M1635 diff_16636_23048# diff_15472_24352# GND GND efet w=106 l=106
+ ad=94416 pd=3256 as=0 ps=0 
M1636 diff_17068_23276# diff_15472_24352# GND GND efet w=130 l=100
+ ad=100464 pd=3496 as=0 ps=0 
M1637 diff_15472_24352# diff_18340_24112# GND GND efet w=426 l=118
+ ad=0 pd=0 as=0 ps=0 
M1638 diff_13792_23696# diff_13816_24208# GND GND efet w=220 l=76
+ ad=0 pd=0 as=0 ps=0 
M1639 diff_14164_25384# diff_13816_24208# GND GND efet w=108 l=82
+ ad=0 pd=0 as=0 ps=0 
M1640 GND diff_13816_24208# diff_15676_23048# GND efet w=106 l=94
+ ad=0 pd=0 as=0 ps=0 
M1641 GND diff_13816_24208# diff_16120_23288# GND efet w=106 l=82
+ ad=0 pd=0 as=0 ps=0 
M1642 diff_14740_23060# diff_14812_24004# GND GND efet w=106 l=106
+ ad=0 pd=0 as=0 ps=0 
M1643 GND diff_13816_24004# diff_13792_23696# GND efet w=232 l=88
+ ad=0 pd=0 as=0 ps=0 
M1644 diff_15124_23692# diff_14812_24004# GND GND efet w=106 l=106
+ ad=0 pd=0 as=0 ps=0 
M1645 diff_11708_24184# clk1 diff_11512_23488# GND efet w=52 l=100
+ ad=0 pd=0 as=3680 ps=264 
M1646 diff_16636_23048# diff_14812_24004# GND GND efet w=100 l=76
+ ad=0 pd=0 as=0 ps=0 
M1647 diff_17068_23276# diff_14812_24004# GND GND efet w=124 l=124
+ ad=0 pd=0 as=0 ps=0 
M1648 Vdd Vdd diff_13816_24208# GND efet w=41 l=338
+ ad=0 pd=0 as=37840 ps=1352 
M1649 diff_14740_23060# diff_13816_24004# GND GND efet w=112 l=124
+ ad=0 pd=0 as=0 ps=0 
M1650 diff_8548_23696# diff_8320_21824# diff_6400_21080# GND efet w=124 l=88
+ ad=0 pd=0 as=0 ps=0 
M1651 diff_8788_23696# diff_8320_21824# diff_6952_20728# GND efet w=82 l=106
+ ad=0 pd=0 as=0 ps=0 
M1652 diff_9028_23696# diff_8740_22024# diff_6952_20728# GND efet w=88 l=88
+ ad=0 pd=0 as=0 ps=0 
M1653 diff_9232_23696# diff_8740_22024# diff_6400_21080# GND efet w=142 l=94
+ ad=0 pd=0 as=0 ps=0 
M1654 GND diff_11068_23716# diff_11216_23416# GND efet w=328 l=88
+ ad=0 pd=0 as=16112 ps=760 
M1655 GND diff_7288_23632# diff_7180_23308# GND efet w=94 l=94
+ ad=0 pd=0 as=32080 ps=1184 
M1656 diff_7768_23848# diff_7768_23620# GND GND efet w=88 l=88
+ ad=18400 pd=640 as=0 ps=0 
M1657 diff_11216_23416# diff_10516_20840# diff_11000_24316# GND efet w=172 l=100
+ ad=0 pd=0 as=0 ps=0 
M1658 diff_11600_23524# diff_11512_23488# GND GND efet w=310 l=94
+ ad=15776 pd=736 as=0 ps=0 
M1659 GND diff_13816_24004# diff_15676_23048# GND efet w=112 l=100
+ ad=0 pd=0 as=0 ps=0 
M1660 diff_11020_25156# diff_10516_20840# diff_11600_23524# GND efet w=154 l=100
+ ad=0 pd=0 as=0 ps=0 
M1661 diff_13792_23696# diff_12916_19724# diff_13708_25372# GND efet w=334 l=94
+ ad=0 pd=0 as=53296 ps=1592 
M1662 diff_13352_23512# Vdd Vdd GND efet w=64 l=328
+ ad=29200 pd=1096 as=0 ps=0 
M1663 GND diff_12916_19724# diff_13352_23512# GND efet w=232 l=88
+ ad=0 pd=0 as=0 ps=0 
M1664 Vdd Vdd diff_8968_23872# GND efet w=40 l=496
+ ad=0 pd=0 as=52960 ps=2032 
M1665 diff_3460_23104# diff_3952_23104# GND GND efet w=154 l=94
+ ad=22048 pd=768 as=0 ps=0 
M1666 Vdd Vdd diff_3460_23104# GND efet w=64 l=532
+ ad=0 pd=0 as=0 ps=0 
M1667 GND diff_3200_23188# diff_2788_24040# GND efet w=106 l=88
+ ad=0 pd=0 as=50032 ps=1624 
M1668 GND diff_5824_22268# diff_5020_23836# GND efet w=352 l=100
+ ad=0 pd=0 as=107984 ps=3536 
M1669 diff_5200_22772# Vdd Vdd GND efet w=58 l=184
+ ad=49952 pd=1832 as=0 ps=0 
M1670 diff_4436_22444# clk2 GND GND efet w=208 l=100
+ ad=116224 pd=4072 as=0 ps=0 
M1671 diff_2788_24040# Vdd Vdd GND efet w=76 l=412
+ ad=0 pd=0 as=0 ps=0 
M1672 diff_2788_24040# clk1 GND GND efet w=124 l=76
+ ad=0 pd=0 as=0 ps=0 
M1673 Vdd Vdd diff_4436_22444# GND efet w=46 l=238
+ ad=0 pd=0 as=0 ps=0 
M1674 GND diff_928_16456# diff_1232_22576# GND efet w=772 l=100
+ ad=0 pd=0 as=0 ps=0 
M1675 diff_2656_22088# diff_2284_21260# Vdd GND efet w=186 l=122
+ ad=111840 pd=3192 as=0 ps=0 
M1676 GND diff_2344_20804# diff_2656_22088# GND efet w=160 l=106
+ ad=0 pd=0 as=0 ps=0 
M1677 diff_2284_21260# diff_2072_21376# diff_2284_21260# GND efet w=462 l=116
+ ad=49728 pd=2536 as=0 ps=0 
M1678 diff_2072_21376# Vdd Vdd GND efet w=52 l=88
+ ad=3536 pd=240 as=0 ps=0 
M1679 GND diff_2344_20804# diff_2284_21260# GND efet w=112 l=88
+ ad=0 pd=0 as=0 ps=0 
M1680 diff_3872_22168# Vdd Vdd GND efet w=58 l=496
+ ad=44864 pd=1616 as=0 ps=0 
M1681 GND diff_2392_18688# diff_3872_22168# GND efet w=124 l=76
+ ad=0 pd=0 as=0 ps=0 
M1682 diff_5212_23848# Vdd Vdd GND efet w=58 l=214
+ ad=42848 pd=1376 as=0 ps=0 
M1683 diff_5020_23836# Vdd Vdd GND efet w=64 l=172
+ ad=0 pd=0 as=0 ps=0 
M1684 diff_5212_23848# clk2 GND GND efet w=412 l=88
+ ad=0 pd=0 as=0 ps=0 
M1685 GND diff_6208_22352# diff_5212_23848# GND efet w=346 l=106
+ ad=0 pd=0 as=0 ps=0 
M1686 diff_5200_22772# clk2 GND GND efet w=436 l=100
+ ad=0 pd=0 as=0 ps=0 
M1687 GND diff_6580_22360# diff_5200_22772# GND efet w=406 l=88
+ ad=0 pd=0 as=0 ps=0 
M1688 Vdd Vdd diff_7180_23308# GND efet w=40 l=508
+ ad=0 pd=0 as=0 ps=0 
M1689 GND diff_8320_21824# diff_8380_23308# GND efet w=88 l=82
+ ad=0 pd=0 as=14656 ps=616 
M1690 diff_8968_23872# diff_8740_22024# GND GND efet w=88 l=88
+ ad=0 pd=0 as=0 ps=0 
M1691 Vdd Vdd diff_7768_23848# GND efet w=46 l=406
+ ad=0 pd=0 as=0 ps=0 
M1692 diff_8380_23308# Vdd Vdd GND efet w=40 l=424
+ ad=0 pd=0 as=0 ps=0 
M1693 diff_7492_22408# diff_7840_22408# GND GND efet w=190 l=82
+ ad=26560 pd=792 as=0 ps=0 
M1694 GND diff_13816_24004# diff_16636_23048# GND efet w=100 l=76
+ ad=0 pd=0 as=0 ps=0 
M1695 GND diff_14320_23620# diff_14164_25384# GND efet w=118 l=82
+ ad=0 pd=0 as=0 ps=0 
M1696 diff_15124_23692# diff_14320_23620# GND GND efet w=112 l=88
+ ad=0 pd=0 as=0 ps=0 
M1697 diff_16120_23288# diff_14320_23620# GND GND efet w=112 l=76
+ ad=0 pd=0 as=0 ps=0 
M1698 diff_17068_23276# diff_14320_23620# GND GND efet w=112 l=94
+ ad=0 pd=0 as=0 ps=0 
M1699 diff_14164_25384# diff_13352_23512# GND GND efet w=112 l=106
+ ad=0 pd=0 as=0 ps=0 
M1700 diff_14740_23060# diff_13352_23512# GND GND efet w=118 l=106
+ ad=0 pd=0 as=0 ps=0 
M1701 diff_15124_23692# diff_13352_23512# GND GND efet w=118 l=94
+ ad=0 pd=0 as=0 ps=0 
M1702 diff_15676_23048# diff_13352_23512# GND GND efet w=130 l=88
+ ad=0 pd=0 as=0 ps=0 
M1703 diff_16120_23288# diff_13352_23512# GND GND efet w=118 l=82
+ ad=0 pd=0 as=0 ps=0 
M1704 GND diff_13352_23512# diff_16636_23048# GND efet w=112 l=88
+ ad=0 pd=0 as=0 ps=0 
M1705 GND diff_13352_23512# diff_17068_23276# GND efet w=112 l=100
+ ad=0 pd=0 as=0 ps=0 
M1706 diff_14164_25384# diff_14236_22696# diff_14164_25384# GND efet w=470 l=242
+ ad=0 pd=0 as=0 ps=0 
M1707 Vdd Vdd diff_7492_22408# GND efet w=64 l=532
+ ad=0 pd=0 as=0 ps=0 
M1708 diff_13708_25372# diff_13744_22612# diff_13708_25372# GND efet w=128 l=412
+ ad=0 pd=0 as=0 ps=0 
M1709 diff_11000_22924# Vdd Vdd GND efet w=52 l=532
+ ad=36496 pd=1336 as=0 ps=0 
M1710 GND diff_11224_22636# diff_11000_22924# GND efet w=112 l=100
+ ad=0 pd=0 as=0 ps=0 
M1711 diff_8320_21824# diff_7492_22408# GND GND efet w=88 l=100
+ ad=72384 pd=2208 as=0 ps=0 
M1712 diff_11224_22636# diff_11000_22924# GND GND efet w=100 l=88
+ ad=42944 pd=1448 as=0 ps=0 
M1713 Vdd Vdd diff_11224_22636# GND efet w=46 l=550
+ ad=0 pd=0 as=0 ps=0 
M1714 diff_9932_21748# Vdd Vdd GND efet w=64 l=556
+ ad=106528 pd=3720 as=0 ps=0 
M1715 GND diff_11224_22636# diff_9932_21748# GND efet w=118 l=100
+ ad=0 pd=0 as=0 ps=0 
M1716 diff_11708_22792# diff_11000_22924# GND GND efet w=112 l=100
+ ad=32320 pd=1360 as=0 ps=0 
M1717 Vdd Vdd diff_11708_22792# GND efet w=64 l=544
+ ad=0 pd=0 as=0 ps=0 
M1718 diff_8740_22024# diff_7840_22408# GND GND efet w=154 l=94
+ ad=69424 pd=3040 as=0 ps=0 
M1719 diff_9932_21748# diff_11020_22492# diff_11068_22336# GND efet w=64 l=88
+ ad=0 pd=0 as=4400 ps=288 
M1720 diff_11708_22792# diff_11020_22492# diff_11512_22108# GND efet w=70 l=94
+ ad=0 pd=0 as=4112 ps=336 
M1721 diff_3872_22168# clk2 diff_5824_22268# GND efet w=52 l=100
+ ad=0 pd=0 as=3824 ps=288 
M1722 diff_6208_22352# clk2 diff_3500_21460# GND efet w=52 l=88
+ ad=3680 pd=264 as=33296 ps=1232 
M1723 diff_6580_22360# clk2 diff_3052_21280# GND efet w=58 l=106
+ ad=3584 pd=264 as=56960 ps=1936 
M1724 diff_2284_21260# diff_2072_21376# Vdd GND efet w=54 l=304
+ ad=0 pd=0 as=0 ps=0 
M1725 diff_3500_21460# diff_2140_4552# GND GND efet w=112 l=88
+ ad=0 pd=0 as=0 ps=0 
M1726 GND diff_2140_5752# diff_3052_21280# GND efet w=124 l=76
+ ad=0 pd=0 as=0 ps=0 
M1727 diff_3052_21280# Vdd Vdd GND efet w=66 l=458
+ ad=0 pd=0 as=0 ps=0 
M1728 Vdd Vdd diff_2344_20804# GND efet w=60 l=284
+ ad=0 pd=0 as=67712 ps=3584 
M1729 diff_2344_20804# clk1 diff_2192_20392# GND efet w=390 l=122
+ ad=0 pd=0 as=24656 ps=864 
M1730 GND diff_1840_19936# diff_2344_20804# GND efet w=178 l=100
+ ad=0 pd=0 as=0 ps=0 
M1731 diff_2344_20804# diff_2068_14080# GND GND efet w=184 l=64
+ ad=0 pd=0 as=0 ps=0 
M1732 diff_2192_20392# diff_1912_20180# GND GND efet w=358 l=94
+ ad=0 pd=0 as=0 ps=0 
M1733 Vdd Vdd diff_1696_20020# GND efet w=46 l=334
+ ad=0 pd=0 as=50208 ps=2248 
M1734 diff_3500_21460# Vdd Vdd GND efet w=46 l=430
+ ad=0 pd=0 as=0 ps=0 
M1735 diff_1912_20180# clk2 diff_1696_20020# GND efet w=112 l=88
+ ad=15584 pd=624 as=0 ps=0 
M1736 GND diff_1840_19936# diff_1696_20020# GND efet w=162 l=98
+ ad=0 pd=0 as=0 ps=0 
M1737 diff_5020_23836# clk2 GND GND efet w=352 l=88
+ ad=0 pd=0 as=0 ps=0 
M1738 diff_7288_23632# diff_7492_22408# GND GND efet w=100 l=76
+ ad=88688 pd=2768 as=0 ps=0 
M1739 diff_7768_23620# diff_7840_22408# GND GND efet w=160 l=76
+ ad=69568 pd=3016 as=0 ps=0 
M1740 diff_7288_23632# diff_7492_22216# GND GND efet w=94 l=76
+ ad=0 pd=0 as=0 ps=0 
M1741 GND diff_7492_22216# diff_7768_23620# GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M1742 GND diff_8344_22228# diff_8320_21824# GND efet w=160 l=76
+ ad=0 pd=0 as=0 ps=0 
M1743 GND diff_8344_22228# diff_8740_22024# GND efet w=160 l=100
+ ad=0 pd=0 as=0 ps=0 
M1744 diff_7288_23632# diff_7324_21436# diff_7288_23632# GND efet w=244 l=290
+ ad=0 pd=0 as=0 ps=0 
M1745 GND diff_1132_21544# diff_1696_20020# GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M1746 Vdd Vdd diff_4156_19880# GND efet w=48 l=568
+ ad=0 pd=0 as=121696 ps=4536 
M1747 diff_7288_23632# diff_7324_21436# Vdd GND efet w=52 l=460
+ ad=0 pd=0 as=0 ps=0 
M1748 diff_7768_23620# diff_7816_21928# diff_7768_23620# GND efet w=492 l=248
+ ad=0 pd=0 as=0 ps=0 
M1749 diff_8320_21824# diff_8272_21388# diff_8320_21824# GND efet w=238 l=490
+ ad=0 pd=0 as=0 ps=0 
M1750 GND diff_11068_22336# diff_11216_22036# GND efet w=316 l=88
+ ad=0 pd=0 as=16160 ps=736 
M1751 diff_11216_22036# diff_11000_21736# diff_11000_22924# GND efet w=172 l=112
+ ad=0 pd=0 as=0 ps=0 
M1752 diff_8740_22024# diff_8764_21368# diff_8740_22024# GND efet w=504 l=260
+ ad=0 pd=0 as=0 ps=0 
M1753 Vdd Vdd diff_6404_20440# GND efet w=50 l=494
+ ad=0 pd=0 as=11440 ps=656 
M1754 diff_7768_23620# diff_7816_21928# Vdd GND efet w=52 l=448
+ ad=0 pd=0 as=0 ps=0 
M1755 diff_8320_21824# diff_8272_21388# Vdd GND efet w=52 l=460
+ ad=0 pd=0 as=0 ps=0 
M1756 diff_7492_22216# diff_8344_22228# GND GND efet w=196 l=88
+ ad=27904 pd=920 as=0 ps=0 
M1757 Vdd Vdd diff_7492_22216# GND efet w=64 l=544
+ ad=0 pd=0 as=0 ps=0 
M1758 diff_11600_22144# diff_11512_22108# GND GND efet w=316 l=100
+ ad=15824 pd=688 as=0 ps=0 
M1759 diff_11224_22636# diff_11000_21736# diff_11600_22144# GND efet w=154 l=106
+ ad=0 pd=0 as=0 ps=0 
M1760 diff_13708_25372# diff_13744_22612# Vdd GND efet w=76 l=454
+ ad=0 pd=0 as=0 ps=0 
M1761 diff_14740_23060# diff_14680_22624# diff_14740_23060# GND efet w=226 l=254
+ ad=0 pd=0 as=0 ps=0 
M1762 diff_14164_25384# diff_14236_22696# Vdd GND efet w=58 l=490
+ ad=0 pd=0 as=0 ps=0 
M1763 diff_14740_23060# diff_14680_22624# Vdd GND efet w=52 l=460
+ ad=0 pd=0 as=0 ps=0 
M1764 diff_15124_23692# diff_15172_22876# diff_15124_23692# GND efet w=234 l=448
+ ad=0 pd=0 as=0 ps=0 
M1765 diff_15676_23048# diff_15616_22684# diff_15676_23048# GND efet w=234 l=426
+ ad=0 pd=0 as=0 ps=0 
M1766 diff_16120_23288# diff_16108_22948# diff_16120_23288# GND efet w=238 l=430
+ ad=0 pd=0 as=0 ps=0 
M1767 diff_15124_23692# diff_15172_22876# Vdd GND efet w=52 l=460
+ ad=0 pd=0 as=0 ps=0 
M1768 diff_13744_22612# Vdd Vdd GND efet w=64 l=88
+ ad=6032 pd=360 as=0 ps=0 
M1769 diff_14236_22696# Vdd Vdd GND efet w=64 l=94
+ ad=5264 pd=312 as=0 ps=0 
M1770 diff_15676_23048# diff_15616_22684# Vdd GND efet w=64 l=484
+ ad=0 pd=0 as=0 ps=0 
M1771 diff_16636_23048# diff_16576_22612# diff_16636_23048# GND efet w=244 l=254
+ ad=0 pd=0 as=0 ps=0 
M1772 diff_16120_23288# diff_16108_22948# Vdd GND efet w=70 l=442
+ ad=0 pd=0 as=0 ps=0 
M1773 diff_14680_22624# Vdd Vdd GND efet w=76 l=76
+ ad=6368 pd=336 as=0 ps=0 
M1774 diff_15172_22876# Vdd Vdd GND efet w=76 l=76
+ ad=6224 pd=336 as=0 ps=0 
M1775 diff_16636_23048# diff_16576_22612# Vdd GND efet w=70 l=454
+ ad=0 pd=0 as=0 ps=0 
M1776 diff_13816_24208# diff_14812_24004# GND GND efet w=208 l=88
+ ad=0 pd=0 as=0 ps=0 
M1777 diff_14812_24004# diff_16420_22148# GND GND efet w=424 l=100
+ ad=44560 pd=1528 as=0 ps=0 
M1778 Vdd Vdd diff_14812_24004# GND efet w=64 l=304
+ ad=0 pd=0 as=0 ps=0 
M1779 Vdd Vdd diff_13816_24004# GND efet w=88 l=346
+ ad=0 pd=0 as=49264 ps=1576 
M1780 diff_17068_23276# diff_17068_22816# diff_17068_23276# GND efet w=244 l=258
+ ad=0 pd=0 as=0 ps=0 
M1781 diff_13816_24004# diff_14320_23620# GND GND efet w=208 l=76
+ ad=0 pd=0 as=0 ps=0 
M1782 diff_14320_23620# diff_13360_22252# GND GND efet w=394 l=82
+ ad=40240 pd=1488 as=0 ps=0 
M1783 Vdd Vdd diff_14320_23620# GND efet w=76 l=358
+ ad=0 pd=0 as=0 ps=0 
M1784 diff_15616_22684# Vdd Vdd GND efet w=64 l=76
+ ad=5264 pd=312 as=0 ps=0 
M1785 diff_16108_22948# Vdd Vdd GND efet w=70 l=82
+ ad=5120 pd=288 as=0 ps=0 
M1786 diff_17068_23276# diff_17068_22816# Vdd GND efet w=52 l=436
+ ad=0 pd=0 as=0 ps=0 
M1787 diff_3244_29488# diff_18892_22660# diff_13360_22252# GND efet w=64 l=100
+ ad=0 pd=0 as=87184 ps=3632 
M1788 diff_3436_29560# diff_18892_22660# diff_16420_22148# GND efet w=52 l=100
+ ad=0 pd=0 as=96768 ps=2752 
M1789 diff_16576_22612# Vdd Vdd GND efet w=82 l=112
+ ad=5456 pd=336 as=0 ps=0 
M1790 diff_17068_22816# Vdd Vdd GND efet w=76 l=88
+ ad=6080 pd=312 as=0 ps=0 
M1791 Vdd Vdd diff_13492_21712# GND efet w=40 l=562
+ ad=0 pd=0 as=73424 ps=1928 
M1792 Vdd Vdd diff_14068_21556# GND efet w=46 l=538
+ ad=0 pd=0 as=80848 ps=2344 
M1793 Vdd Vdd diff_14824_21716# GND efet w=40 l=544
+ ad=0 pd=0 as=23632 ps=1096 
M1794 Vdd Vdd diff_15892_21560# GND efet w=40 l=520
+ ad=0 pd=0 as=69248 ps=1712 
M1795 diff_13360_22252# diff_13816_22024# diff_14012_21652# GND efet w=64 l=88
+ ad=0 pd=0 as=65184 ps=1976 
M1796 Vdd Vdd diff_14012_21652# GND efet w=40 l=268
+ ad=0 pd=0 as=0 ps=0 
M1797 Vdd Vdd diff_16456_21556# GND efet w=40 l=592
+ ad=0 pd=0 as=83968 ps=2392 
M1798 Vdd Vdd diff_17212_21704# GND efet w=40 l=520
+ ad=0 pd=0 as=24928 ps=1048 
M1799 diff_16400_21640# Vdd Vdd GND efet w=50 l=334
+ ad=69504 pd=1952 as=0 ps=0 
M1800 diff_16420_22148# diff_13816_22024# diff_16400_21640# GND efet w=82 l=82
+ ad=0 pd=0 as=0 ps=0 
M1801 diff_5704_20956# diff_5656_20560# diff_5704_20956# GND efet w=596 l=240
+ ad=127008 pd=5144 as=0 ps=0 
M1802 diff_7324_21436# Vdd Vdd GND efet w=76 l=88
+ ad=6080 pd=312 as=0 ps=0 
M1803 diff_7816_21928# Vdd Vdd GND efet w=88 l=76
+ ad=5840 pd=312 as=0 ps=0 
M1804 diff_8740_22024# diff_8764_21368# Vdd GND efet w=52 l=436
+ ad=0 pd=0 as=0 ps=0 
M1805 diff_7840_22408# diff_2104_10732# diff_9412_21772# GND efet w=64 l=88
+ ad=18656 pd=648 as=0 ps=0 
M1806 diff_9932_21748# diff_2392_18688# diff_7840_22408# GND efet w=64 l=88
+ ad=0 pd=0 as=0 ps=0 
M1807 diff_8344_22228# diff_2104_10732# diff_9412_21556# GND efet w=64 l=88
+ ad=8800 pd=648 as=0 ps=0 
M1808 diff_9932_21580# diff_2392_18688# diff_8344_22228# GND efet w=58 l=100
+ ad=125328 pd=4184 as=0 ps=0 
M1809 diff_8272_21388# Vdd Vdd GND efet w=82 l=76
+ ad=6176 pd=336 as=0 ps=0 
M1810 diff_8764_21368# Vdd Vdd GND efet w=88 l=88
+ ad=5840 pd=336 as=0 ps=0 
M1811 diff_6400_21080# diff_5704_20956# Vdd GND efet w=330 l=170
+ ad=0 pd=0 as=0 ps=0 
M1812 Vdd Vdd diff_5656_20560# GND efet w=58 l=94
+ ad=0 pd=0 as=3248 ps=248 
M1813 Vdd diff_5656_20560# diff_5704_20956# GND efet w=40 l=352
+ ad=0 pd=0 as=0 ps=0 
M1814 GND diff_6404_20440# diff_6400_21080# GND efet w=238 l=94
+ ad=0 pd=0 as=0 ps=0 
M1815 Vdd Vdd diff_7084_20800# GND efet w=64 l=418
+ ad=0 pd=0 as=13936 ps=872 
M1816 GND diff_7084_20800# diff_6952_20728# GND efet w=160 l=76
+ ad=0 pd=0 as=0 ps=0 
M1817 Vdd diff_8068_20716# diff_7084_20632# GND efet w=52 l=328
+ ad=0 pd=0 as=88192 ps=4784 
M1818 GND diff_4996_19156# diff_4928_19924# GND efet w=270 l=110
+ ad=0 pd=0 as=16592 ps=624 
M1819 Vdd Vdd diff_4700_19432# GND efet w=46 l=562
+ ad=0 pd=0 as=94176 ps=3440 
M1820 diff_4700_19924# diff_2212_11356# diff_4156_19880# GND efet w=244 l=88
+ ad=34160 pd=768 as=0 ps=0 
M1821 diff_4928_19924# diff_4576_17684# diff_4700_19924# GND efet w=244 l=88
+ ad=0 pd=0 as=0 ps=0 
M1822 diff_5084_19444# diff_1840_19936# GND GND efet w=262 l=94
+ ad=45184 pd=1984 as=0 ps=0 
M1823 diff_4156_19880# diff_1132_21544# GND GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M1824 diff_5084_19444# diff_4996_19156# diff_4928_19444# GND efet w=298 l=160
+ ad=0 pd=0 as=15776 ps=600 
M1825 diff_4376_19432# diff_3868_15448# GND GND efet w=244 l=100
+ ad=18992 pd=648 as=0 ps=0 
M1826 diff_4544_19444# diff_4456_18616# diff_4376_19432# GND efet w=232 l=100
+ ad=16352 pd=624 as=0 ps=0 
M1827 diff_4700_19432# diff_2212_11356# diff_4544_19444# GND efet w=244 l=88
+ ad=0 pd=0 as=0 ps=0 
M1828 diff_4928_19444# diff_4576_17684# diff_4700_19432# GND efet w=232 l=88
+ ad=0 pd=0 as=0 ps=0 
M1829 diff_5240_19432# diff_5152_19192# diff_5084_19444# GND efet w=244 l=88
+ ad=16592 pd=624 as=0 ps=0 
M1830 diff_4700_19432# diff_5308_19396# diff_5240_19432# GND efet w=250 l=94
+ ad=0 pd=0 as=0 ps=0 
M1831 diff_6404_20440# diff_5704_20956# GND GND efet w=100 l=112
+ ad=0 pd=0 as=0 ps=0 
M1832 Vdd Vdd diff_8068_20716# GND efet w=40 l=76
+ ad=0 pd=0 as=3200 ps=240 
M1833 Vdd Vdd diff_8668_20836# GND efet w=40 l=88
+ ad=0 pd=0 as=3536 ps=288 
M1834 Vdd diff_8668_20836# diff_8680_20596# GND efet w=58 l=142
+ ad=0 pd=0 as=192656 ps=6240 
M1835 diff_7084_20632# diff_8068_20716# diff_7084_20632# GND efet w=390 l=188
+ ad=0 pd=0 as=0 ps=0 
M1836 Vdd diff_7084_20632# diff_6952_20728# GND efet w=166 l=94
+ ad=0 pd=0 as=0 ps=0 
M1837 GND diff_7084_20632# diff_7084_20800# GND efet w=106 l=106
+ ad=0 pd=0 as=0 ps=0 
M1838 diff_8680_20596# diff_8668_20836# diff_8680_20596# GND efet w=662 l=186
+ ad=0 pd=0 as=0 ps=0 
M1839 diff_8680_20596# diff_9280_20260# GND GND efet w=286 l=94
+ ad=0 pd=0 as=0 ps=0 
M1840 GND diff_6532_20236# diff_8680_20596# GND efet w=292 l=88
+ ad=0 pd=0 as=0 ps=0 
M1841 GND diff_9592_20488# diff_8680_20596# GND efet w=280 l=88
+ ad=0 pd=0 as=0 ps=0 
M1842 Vdd Vdd diff_6688_20020# GND efet w=40 l=412
+ ad=0 pd=0 as=12112 ps=752 
M1843 diff_5704_20956# diff_6532_20236# GND GND efet w=106 l=82
+ ad=0 pd=0 as=0 ps=0 
M1844 diff_7084_20632# diff_7744_20500# GND GND efet w=106 l=82
+ ad=0 pd=0 as=0 ps=0 
M1845 diff_7084_20632# diff_7516_20284# diff_7408_20204# GND efet w=238 l=82
+ ad=0 pd=0 as=24416 ps=936 
M1846 diff_5704_20956# diff_4192_12940# GND GND efet w=118 l=94
+ ad=0 pd=0 as=0 ps=0 
M1847 GND diff_6496_19828# diff_5704_20956# GND efet w=112 l=94
+ ad=0 pd=0 as=0 ps=0 
M1848 diff_5704_20956# diff_6688_20020# GND GND efet w=112 l=88
+ ad=0 pd=0 as=0 ps=0 
M1849 diff_7408_20204# diff_4456_18616# GND GND efet w=238 l=82
+ ad=0 pd=0 as=0 ps=0 
M1850 GND diff_7324_19300# diff_7084_20632# GND efet w=118 l=82
+ ad=0 pd=0 as=0 ps=0 
M1851 GND diff_2140_5752# diff_4700_19432# GND efet w=142 l=106
+ ad=0 pd=0 as=0 ps=0 
M1852 diff_6688_20020# clk2 GND GND efet w=112 l=76
+ ad=0 pd=0 as=0 ps=0 
M1853 GND diff_4456_14788# diff_5308_19396# GND efet w=270 l=110
+ ad=0 pd=0 as=76976 ps=3328 
M1854 diff_5308_19396# diff_3868_15448# GND GND efet w=214 l=106
+ ad=0 pd=0 as=0 ps=0 
M1855 diff_4556_18160# diff_3868_15448# diff_3856_18340# GND efet w=262 l=76
+ ad=19520 pd=648 as=214960 ps=9008 
M1856 diff_3856_18340# diff_2140_4552# GND GND efet w=94 l=82
+ ad=0 pd=0 as=0 ps=0 
M1857 diff_4712_18160# diff_4456_18616# diff_4556_18160# GND efet w=256 l=76
+ ad=18896 pd=672 as=0 ps=0 
M1858 GND diff_2392_18688# diff_4712_18160# GND efet w=244 l=76
+ ad=0 pd=0 as=0 ps=0 
M1859 Vdd Vdd diff_3856_18340# GND efet w=58 l=526
+ ad=0 pd=0 as=0 ps=0 
M1860 diff_5240_18248# diff_4576_17684# diff_5092_17944# GND efet w=292 l=88
+ ad=21584 pd=768 as=105872 ps=3152 
M1861 diff_3856_18340# diff_4996_19156# diff_5240_18248# GND efet w=310 l=82
+ ad=0 pd=0 as=0 ps=0 
M1862 diff_5624_18136# diff_5152_19192# diff_3856_18340# GND efet w=268 l=88
+ ad=18224 pd=672 as=0 ps=0 
M1863 diff_5092_17944# diff_5308_19396# diff_5624_18136# GND efet w=268 l=88
+ ad=0 pd=0 as=0 ps=0 
M1864 GND diff_2068_14080# diff_5092_17944# GND efet w=280 l=76
+ ad=0 pd=0 as=0 ps=0 
M1865 GND diff_3868_15448# diff_4576_17684# GND efet w=220 l=82
+ ad=0 pd=0 as=19648 ps=880 
M1866 diff_4576_17684# Vdd Vdd GND efet w=40 l=220
+ ad=0 pd=0 as=0 ps=0 
M1867 diff_5308_19396# Vdd Vdd GND efet w=46 l=226
+ ad=0 pd=0 as=0 ps=0 
M1868 diff_4408_17236# diff_4936_17224# Vdd GND efet w=46 l=226
+ ad=58656 pd=2984 as=0 ps=0 
M1869 Vdd diff_4408_17236# diff_3868_15448# GND efet w=304 l=88
+ ad=0 pd=0 as=105632 ps=2256 
M1870 Vdd Vdd diff_4936_17224# GND efet w=46 l=100
+ ad=0 pd=0 as=2912 ps=240 
M1871 GND diff_2104_10732# diff_6496_19828# GND efet w=118 l=94
+ ad=0 pd=0 as=56448 ps=2504 
M1872 GND diff_2392_18688# diff_6496_19828# GND efet w=94 l=94
+ ad=0 pd=0 as=0 ps=0 
M1873 Vdd Vdd diff_7744_20500# GND efet w=46 l=418
+ ad=0 pd=0 as=22384 ps=832 
M1874 diff_6496_19828# Vdd Vdd GND efet w=40 l=544
+ ad=0 pd=0 as=0 ps=0 
M1875 diff_7744_20500# clk1 GND GND efet w=112 l=76
+ ad=0 pd=0 as=0 ps=0 
M1876 Vdd Vdd diff_7228_18940# GND efet w=40 l=220
+ ad=0 pd=0 as=43712 ps=1848 
M1877 Vdd Vdd diff_6532_20236# GND efet w=40 l=232
+ ad=0 pd=0 as=72144 ps=2512 
M1878 diff_9080_19840# Vdd Vdd GND efet w=58 l=442
+ ad=87360 pd=2840 as=0 ps=0 
M1879 diff_9280_20260# clk2 diff_9080_19840# GND efet w=70 l=118
+ ad=9104 pd=552 as=0 ps=0 
M1880 diff_11000_21736# Vdd Vdd GND efet w=46 l=598
+ ad=35392 pd=1360 as=0 ps=0 
M1881 GND diff_11020_22492# diff_11000_21736# GND efet w=88 l=88
+ ad=0 pd=0 as=0 ps=0 
M1882 diff_11020_22492# diff_11000_21736# GND GND efet w=100 l=88
+ ad=45808 pd=1664 as=0 ps=0 
M1883 Vdd Vdd diff_11020_22492# GND efet w=46 l=532
+ ad=0 pd=0 as=0 ps=0 
M1884 GND diff_11020_22492# diff_9932_21580# GND efet w=148 l=76
+ ad=0 pd=0 as=0 ps=0 
M1885 diff_9932_21580# Vdd Vdd GND efet w=58 l=562
+ ad=0 pd=0 as=0 ps=0 
M1886 diff_11708_21568# diff_11000_21736# GND GND efet w=112 l=88
+ ad=31936 pd=1384 as=0 ps=0 
M1887 Vdd Vdd diff_11708_21568# GND efet w=70 l=622
+ ad=0 pd=0 as=0 ps=0 
M1888 diff_9932_21580# clk1 diff_11068_21100# GND efet w=64 l=82
+ ad=0 pd=0 as=4208 ps=288 
M1889 diff_11708_21568# clk1 diff_11512_20872# GND efet w=52 l=76
+ ad=0 pd=0 as=4160 ps=264 
M1890 diff_14012_21652# clk1 diff_13408_21340# GND efet w=58 l=118
+ ad=0 pd=0 as=3488 ps=240 
M1891 diff_13492_21712# diff_13336_21568# diff_13468_21416# GND efet w=196 l=94
+ ad=0 pd=0 as=17216 ps=720 
M1892 diff_13468_21416# diff_13408_21340# GND GND efet w=274 l=94
+ ad=0 pd=0 as=0 ps=0 
M1893 diff_14012_21652# diff_14068_21556# GND GND efet w=172 l=88
+ ad=0 pd=0 as=0 ps=0 
M1894 GND diff_14068_21556# diff_13492_21712# GND efet w=94 l=94
+ ad=0 pd=0 as=0 ps=0 
M1895 diff_15116_21748# clk1 diff_14824_21716# GND efet w=58 l=106
+ ad=3344 pd=264 as=0 ps=0 
M1896 diff_14824_21716# diff_13492_21712# GND GND efet w=94 l=94
+ ad=0 pd=0 as=0 ps=0 
M1897 diff_14068_21556# diff_13492_21712# GND GND efet w=94 l=94
+ ad=0 pd=0 as=0 ps=0 
M1898 diff_16400_21640# diff_13492_21712# diff_15796_21328# GND efet w=76 l=94
+ ad=0 pd=0 as=2960 ps=240 
M1899 GND diff_11068_21100# diff_11216_20812# GND efet w=316 l=100
+ ad=0 pd=0 as=15728 ps=712 
M1900 Vdd Vdd diff_10264_20224# GND efet w=52 l=532
+ ad=0 pd=0 as=26464 ps=1416 
M1901 diff_10516_20840# Vdd Vdd GND efet w=46 l=226
+ ad=44768 pd=1368 as=0 ps=0 
M1902 diff_11216_20812# diff_11060_20488# diff_11000_21736# GND efet w=154 l=112
+ ad=0 pd=0 as=0 ps=0 
M1903 diff_11600_20908# diff_11512_20872# GND GND efet w=316 l=88
+ ad=15824 pd=688 as=0 ps=0 
M1904 diff_11020_22492# diff_11060_20488# diff_11600_20908# GND efet w=160 l=100
+ ad=0 pd=0 as=0 ps=0 
M1905 diff_14068_21556# diff_13336_21568# diff_15232_21416# GND efet w=166 l=94
+ ad=0 pd=0 as=17696 ps=696 
M1906 diff_17516_21736# diff_13492_21712# diff_17212_21704# GND efet w=64 l=100
+ ad=4160 pd=288 as=0 ps=0 
M1907 GND diff_15892_21560# diff_17212_21704# GND efet w=100 l=94
+ ad=0 pd=0 as=0 ps=0 
M1908 diff_15892_21560# diff_14068_21556# diff_15856_21436# GND efet w=172 l=100
+ ad=0 pd=0 as=17744 ps=696 
M1909 diff_16400_21640# diff_16456_21556# GND GND efet w=172 l=76
+ ad=0 pd=0 as=0 ps=0 
M1910 diff_15892_21560# diff_16456_21556# GND GND efet w=88 l=76
+ ad=0 pd=0 as=0 ps=0 
M1911 diff_15232_21416# diff_15116_21748# GND GND efet w=286 l=100
+ ad=0 pd=0 as=0 ps=0 
M1912 diff_15856_21436# diff_15796_21328# GND GND efet w=268 l=88
+ ad=0 pd=0 as=0 ps=0 
M1913 GND diff_8908_18832# diff_11872_25876# GND efet w=250 l=118
+ ad=0 pd=0 as=0 ps=0 
M1914 GND diff_12416_19756# diff_11872_25876# GND efet w=328 l=94
+ ad=0 pd=0 as=0 ps=0 
M1915 GND diff_10264_20224# diff_10516_20840# GND efet w=208 l=88
+ ad=0 pd=0 as=0 ps=0 
M1916 Vdd Vdd diff_9592_20488# GND efet w=40 l=292
+ ad=0 pd=0 as=35104 ps=1528 
M1917 diff_11060_20488# diff_10972_20356# GND GND efet w=214 l=100
+ ad=116384 pd=5008 as=0 ps=0 
M1918 diff_11872_25876# clk2 GND GND efet w=232 l=100
+ ad=0 pd=0 as=0 ps=0 
M1919 Vdd Vdd diff_11060_20488# GND efet w=70 l=248
+ ad=0 pd=0 as=0 ps=0 
M1920 GND clk2 diff_10664_19996# GND efet w=238 l=118
+ ad=0 pd=0 as=21296 ps=744 
M1921 diff_10664_19996# diff_2392_18688# diff_10508_20008# GND efet w=250 l=94
+ ad=0 pd=0 as=16064 ps=624 
M1922 diff_7172_18664# diff_2104_10732# GND GND efet w=172 l=100
+ ad=11696 pd=480 as=0 ps=0 
M1923 diff_7324_19300# clk2 diff_7160_18400# GND efet w=58 l=94
+ ad=5120 pd=392 as=51744 ps=2304 
M1924 diff_7160_18400# diff_7228_18940# diff_7172_18664# GND efet w=172 l=88
+ ad=0 pd=0 as=0 ps=0 
M1925 GND diff_6532_20236# diff_7228_18940# GND efet w=208 l=106
+ ad=0 pd=0 as=0 ps=0 
M1926 GND diff_8476_18004# diff_6532_20236# GND efet w=208 l=88
+ ad=0 pd=0 as=0 ps=0 
M1927 GND diff_2068_14080# diff_9080_19840# GND efet w=148 l=88
+ ad=0 pd=0 as=0 ps=0 
M1928 diff_7516_20284# diff_3868_15448# GND GND efet w=112 l=82
+ ad=29488 pd=1384 as=0 ps=0 
M1929 Vdd Vdd diff_8308_18688# GND efet w=40 l=424
+ ad=0 pd=0 as=20368 ps=920 
M1930 diff_7160_18400# Vdd Vdd GND efet w=40 l=532
+ ad=0 pd=0 as=0 ps=0 
M1931 diff_7160_18400# diff_1132_21544# GND GND efet w=116 l=82
+ ad=0 pd=0 as=0 ps=0 
M1932 diff_7516_20284# Vdd Vdd GND efet w=52 l=388
+ ad=0 pd=0 as=0 ps=0 
M1933 GND diff_8908_18832# diff_8476_18344# GND efet w=238 l=94
+ ad=0 pd=0 as=98368 ps=3520 
M1934 diff_9592_20488# clk1 GND GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M1935 diff_10508_20008# diff_7228_18940# diff_10264_20224# GND efet w=232 l=88
+ ad=0 pd=0 as=0 ps=0 
M1936 GND diff_2212_11356# diff_9080_19840# GND efet w=118 l=94
+ ad=0 pd=0 as=0 ps=0 
M1937 GND diff_4456_14788# diff_8308_18688# GND efet w=130 l=88
+ ad=0 pd=0 as=0 ps=0 
M1938 GND diff_3868_15448# diff_9064_18608# GND efet w=172 l=88
+ ad=0 pd=0 as=11696 ps=480 
M1939 diff_9064_18608# diff_4456_18616# diff_8476_18004# GND efet w=202 l=82
+ ad=0 pd=0 as=105968 ps=3464 
M1940 diff_8476_18344# diff_8308_18688# diff_8476_18188# GND efet w=238 l=94
+ ad=0 pd=0 as=15776 ps=600 
M1941 diff_8476_18188# diff_5152_19192# diff_8476_18004# GND efet w=232 l=88
+ ad=0 pd=0 as=0 ps=0 
M1942 diff_8476_18344# diff_4996_19156# diff_8476_18004# GND efet w=172 l=88
+ ad=0 pd=0 as=0 ps=0 
M1943 diff_10972_20356# Vdd diff_10972_20356# GND efet w=20 l=548
+ ad=104656 pd=4944 as=0 ps=0 
M1944 diff_10904_19228# diff_10792_18352# GND GND efet w=244 l=88
+ ad=16592 pd=624 as=0 ps=0 
M1945 diff_11060_19228# diff_2068_14080# diff_10904_19228# GND efet w=256 l=88
+ ad=16544 pd=648 as=0 ps=0 
M1946 diff_10972_20356# diff_8908_18832# diff_11060_19228# GND efet w=244 l=88
+ ad=0 pd=0 as=0 ps=0 
M1947 Vdd Vdd diff_11524_19384# GND efet w=40 l=268
+ ad=0 pd=0 as=22816 ps=1064 
M1948 Vdd Vdd diff_11984_19228# GND efet w=40 l=574
+ ad=0 pd=0 as=63216 ps=2312 
M1949 diff_12416_19756# clk2 diff_11984_19228# GND efet w=100 l=100
+ ad=6128 pd=344 as=0 ps=0 
M1950 GND clk2 diff_11524_19384# GND efet w=172 l=88
+ ad=0 pd=0 as=0 ps=0 
M1951 diff_16456_21556# diff_15892_21560# GND GND efet w=94 l=82
+ ad=0 pd=0 as=0 ps=0 
M1952 diff_16456_21556# diff_14068_21556# diff_17668_21404# GND efet w=172 l=100
+ ad=0 pd=0 as=17648 ps=720 
M1953 diff_17668_21404# diff_17516_21736# GND GND efet w=292 l=88
+ ad=0 pd=0 as=0 ps=0 
M1954 diff_3808_28348# diff_18892_22660# diff_18340_24112# GND efet w=72 l=104
+ ad=0 pd=0 as=82448 ps=2696 
M1955 Vdd Vdd diff_18316_21548# GND efet w=40 l=532
+ ad=0 pd=0 as=71120 ps=1760 
M1956 Vdd Vdd diff_18880_21544# GND efet w=46 l=550
+ ad=0 pd=0 as=87424 ps=2368 
M1957 Vdd Vdd diff_19648_21692# GND efet w=52 l=568
+ ad=0 pd=0 as=25024 ps=1032 
M1958 diff_18340_24112# diff_13816_22024# diff_18824_21640# GND efet w=52 l=88
+ ad=0 pd=0 as=65472 ps=1880 
M1959 Vdd Vdd diff_18824_21640# GND efet w=34 l=274
+ ad=0 pd=0 as=0 ps=0 
M1960 diff_18824_21640# diff_15892_21560# diff_18220_21328# GND efet w=58 l=94
+ ad=0 pd=0 as=2768 ps=272 
M1961 diff_18316_21548# diff_16456_21556# diff_18292_21404# GND efet w=166 l=94
+ ad=0 pd=0 as=19952 ps=720 
M1962 diff_18824_21640# diff_18880_21544# GND GND efet w=172 l=88
+ ad=0 pd=0 as=0 ps=0 
M1963 diff_18316_21548# diff_18880_21544# GND GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M1964 diff_18292_21404# diff_18220_21328# GND GND efet w=292 l=88
+ ad=0 pd=0 as=0 ps=0 
M1965 diff_19928_21736# diff_15892_21560# diff_19648_21692# GND efet w=78 l=122
+ ad=4448 pd=296 as=0 ps=0 
M1966 diff_19648_21692# diff_18316_21548# GND GND efet w=88 l=76
+ ad=0 pd=0 as=0 ps=0 
M1967 diff_18880_21544# diff_18316_21548# GND GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M1968 diff_18880_21544# diff_16456_21556# diff_20092_21392# GND efet w=192 l=128
+ ad=0 pd=0 as=17984 ps=680 
M1969 diff_20092_21392# diff_19928_21736# GND GND efet w=268 l=88
+ ad=0 pd=0 as=0 ps=0 
M1970 Vdd Vdd diff_12916_19724# GND efet w=40 l=418
+ ad=0 pd=0 as=151392 ps=6568 
M1971 GND diff_16300_20812# diff_12328_25804# GND efet w=196 l=88
+ ad=0 pd=0 as=76944 ps=2224 
M1972 GND diff_16732_20032# diff_13336_21568# GND efet w=166 l=94
+ ad=0 pd=0 as=42320 ps=1712 
M1973 diff_17152_20864# diff_17080_20656# diff_17152_20864# GND efet w=450 l=224
+ ad=162608 pd=7200 as=0 ps=0 
M1974 diff_12136_25792# diff_8908_18832# GND GND efet w=316 l=112
+ ad=0 pd=0 as=0 ps=0 
M1975 Vdd Vdd diff_13744_19760# GND efet w=40 l=580
+ ad=0 pd=0 as=60544 ps=2176 
M1976 GND diff_14128_19912# diff_12136_25792# GND efet w=298 l=116
+ ad=0 pd=0 as=0 ps=0 
M1977 GND clk2 diff_12136_25792# GND efet w=280 l=124
+ ad=0 pd=0 as=0 ps=0 
M1978 GND diff_11524_19384# diff_11060_20488# GND efet w=238 l=94
+ ad=0 pd=0 as=0 ps=0 
M1979 diff_13744_19760# clk2 diff_14128_19912# GND efet w=130 l=82
+ ad=0 pd=0 as=7856 ps=456 
M1980 diff_11828_19228# diff_2212_11356# GND GND efet w=178 l=94
+ ad=11456 pd=480 as=0 ps=0 
M1981 diff_12164_19364# diff_12028_18580# diff_11984_19228# GND efet w=262 l=106
+ ad=16544 pd=648 as=0 ps=0 
M1982 diff_11984_19228# diff_11884_18124# diff_11828_19228# GND efet w=172 l=94
+ ad=0 pd=0 as=0 ps=0 
M1983 diff_12344_19228# diff_2104_10732# diff_12164_19364# GND efet w=238 l=106
+ ad=13664 pd=600 as=0 ps=0 
M1984 diff_10664_18676# diff_10564_18232# GND GND efet w=186 l=94
+ ad=54800 pd=1816 as=0 ps=0 
M1985 diff_10664_18676# diff_2068_14080# diff_10972_20356# GND efet w=202 l=106
+ ad=0 pd=0 as=0 ps=0 
M1986 diff_10972_20356# diff_2212_11356# diff_10664_18676# GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M1987 diff_10972_20356# diff_2104_10732# diff_10664_18676# GND efet w=172 l=100
+ ad=0 pd=0 as=0 ps=0 
M1988 GND diff_12100_17968# diff_12344_19228# GND efet w=244 l=100
+ ad=0 pd=0 as=0 ps=0 
M1989 diff_13744_19760# diff_2104_10732# diff_13564_19592# GND efet w=250 l=118
+ ad=0 pd=0 as=84592 ps=3184 
M1990 diff_12916_19724# diff_2104_10732# diff_12856_19024# GND efet w=346 l=106
+ ad=0 pd=0 as=49616 ps=2200 
M1991 Vdd Vdd diff_8908_18832# GND efet w=64 l=196
+ ad=0 pd=0 as=64720 ps=2840 
M1992 diff_12328_25804# Vdd Vdd GND efet w=40 l=268
+ ad=0 pd=0 as=0 ps=0 
M1993 diff_15664_19120# Vdd Vdd GND efet w=40 l=568
+ ad=44704 pd=2288 as=0 ps=0 
M1994 diff_12544_25804# Vdd Vdd GND efet w=52 l=232
+ ad=163872 pd=5608 as=0 ps=0 
M1995 diff_13336_21568# Vdd Vdd GND efet w=40 l=292
+ ad=0 pd=0 as=0 ps=0 
M1996 diff_17152_20864# diff_17080_20656# Vdd GND efet w=76 l=220
+ ad=0 pd=0 as=0 ps=0 
M1997 diff_17152_20864# diff_17452_19928# GND GND efet w=300 l=116
+ ad=0 pd=0 as=0 ps=0 
M1998 GND diff_18040_19532# diff_18220_20996# GND efet w=94 l=94
+ ad=0 pd=0 as=55680 ps=2456 
M1999 diff_18220_20996# diff_18148_20656# diff_18220_20996# GND efet w=426 l=236
+ ad=0 pd=0 as=0 ps=0 
M2000 Vdd diff_18148_20656# diff_18220_20996# GND efet w=46 l=442
+ ad=0 pd=0 as=0 ps=0 
M2001 GND diff_18040_19532# diff_13972_25108# GND efet w=160 l=88
+ ad=0 pd=0 as=0 ps=0 
M2002 GND diff_19228_20764# diff_19900_20720# GND efet w=88 l=88
+ ad=0 pd=0 as=21040 ps=1176 
M2003 diff_19228_20764# diff_19156_20272# diff_19228_20764# GND efet w=426 l=146
+ ad=150656 pd=5664 as=0 ps=0 
M2004 diff_13972_25108# diff_18220_20996# Vdd GND efet w=148 l=88
+ ad=0 pd=0 as=0 ps=0 
M2005 diff_13720_25264# diff_19900_20720# GND GND efet w=192 l=88
+ ad=0 pd=0 as=0 ps=0 
M2006 diff_17080_20656# Vdd Vdd GND efet w=46 l=82
+ ad=3536 pd=288 as=0 ps=0 
M2007 diff_12544_25804# diff_15664_19120# GND GND efet w=268 l=110
+ ad=0 pd=0 as=0 ps=0 
M2008 diff_13564_19592# diff_8944_12928# diff_13564_19468# GND efet w=430 l=94
+ ad=0 pd=0 as=26960 ps=984 
M2009 diff_13004_19000# diff_8944_12928# diff_12856_19024# GND efet w=654 l=104
+ ad=27056 pd=1120 as=0 ps=0 
M2010 GND diff_11548_16012# diff_13004_19000# GND efet w=346 l=106
+ ad=0 pd=0 as=0 ps=0 
M2011 diff_8476_18004# Vdd Vdd GND efet w=40 l=496
+ ad=0 pd=0 as=0 ps=0 
M2012 GND diff_7864_17452# diff_7912_17540# GND efet w=256 l=94
+ ad=0 pd=0 as=122080 ps=4792 
M2013 diff_8212_16444# diff_7864_17452# GND GND efet w=262 l=82
+ ad=121232 pd=5024 as=0 ps=0 
M2014 GND diff_12100_17968# diff_13564_19468# GND efet w=238 l=94
+ ad=0 pd=0 as=0 ps=0 
M2015 GND diff_3868_15448# diff_14344_18812# GND efet w=238 l=106
+ ad=0 pd=0 as=39920 ps=1576 
M2016 diff_8908_18832# diff_3868_15448# GND GND efet w=490 l=100
+ ad=0 pd=0 as=0 ps=0 
M2017 GND diff_11884_18124# diff_13564_19592# GND efet w=172 l=76
+ ad=0 pd=0 as=0 ps=0 
M2018 diff_12028_18580# diff_8944_12928# GND GND efet w=448 l=88
+ ad=62048 pd=2112 as=0 ps=0 
M2019 GND diff_8908_18832# diff_15316_19232# GND efet w=244 l=88
+ ad=0 pd=0 as=16592 ps=624 
M2020 diff_15316_19232# diff_11884_18124# diff_15316_19108# GND efet w=250 l=82
+ ad=0 pd=0 as=48080 ps=1704 
M2021 diff_16732_20032# Vdd Vdd GND efet w=40 l=580
+ ad=28000 pd=1096 as=0 ps=0 
M2022 Vdd Vdd diff_17452_19928# GND efet w=40 l=580
+ ad=0 pd=0 as=73600 ps=2872 
M2023 diff_18148_20656# Vdd Vdd GND efet w=52 l=88
+ ad=4160 pd=264 as=0 ps=0 
M2024 diff_17452_19928# clk2 diff_17452_19432# GND efet w=244 l=76
+ ad=0 pd=0 as=34160 ps=1352 
M2025 diff_16732_20032# clk2 diff_16936_19336# GND efet w=244 l=88
+ ad=0 pd=0 as=28688 ps=1328 
M2026 diff_14344_18812# diff_2392_18688# diff_14344_18676# GND efet w=298 l=94
+ ad=0 pd=0 as=45824 ps=2120 
M2027 diff_14992_18404# diff_14872_18520# GND GND efet w=238 l=116
+ ad=45440 pd=1464 as=0 ps=0 
M2028 diff_12028_18580# Vdd Vdd GND efet w=40 l=220
+ ad=0 pd=0 as=0 ps=0 
M2029 GND diff_8908_18832# diff_8920_12124# GND efet w=196 l=88
+ ad=0 pd=0 as=144656 ps=5784 
M2030 GND diff_14516_18124# diff_14176_18496# GND efet w=226 l=112
+ ad=0 pd=0 as=28272 ps=1288 
M2031 diff_15316_19108# diff_8944_12928# diff_14872_18520# GND efet w=442 l=94
+ ad=0 pd=0 as=36224 ps=1464 
M2032 diff_14176_18496# Vdd Vdd GND efet w=40 l=220
+ ad=0 pd=0 as=0 ps=0 
M2033 diff_15992_19108# diff_14992_18404# diff_15836_18652# GND efet w=274 l=128
+ ad=14144 pd=648 as=40960 ps=2160 
M2034 GND diff_1840_19936# diff_15992_19108# GND efet w=274 l=100
+ ad=0 pd=0 as=0 ps=0 
M2035 diff_16376_19108# diff_2068_14080# GND GND efet w=250 l=106
+ ad=13664 pd=600 as=0 ps=0 
M2036 diff_16532_18520# diff_14992_18404# diff_16376_19108# GND efet w=244 l=100
+ ad=44416 pd=1912 as=0 ps=0 
M2037 diff_15836_18652# clk2 diff_15664_19120# GND efet w=274 l=94
+ ad=0 pd=0 as=0 ps=0 
M2038 diff_15992_18424# diff_8944_12928# diff_15836_18652# GND efet w=432 l=110
+ ad=18848 pd=936 as=0 ps=0 
M2039 diff_14516_18124# diff_13672_16400# diff_14344_18676# GND efet w=250 l=94
+ ad=19792 pd=840 as=0 ps=0 
M2040 Vdd Vdd diff_14516_18124# GND efet w=46 l=526
+ ad=0 pd=0 as=0 ps=0 
M2041 diff_14992_18404# Vdd Vdd GND efet w=40 l=220
+ ad=0 pd=0 as=0 ps=0 
M2042 diff_9784_10948# diff_7864_17452# GND GND efet w=244 l=122
+ ad=149984 pd=6000 as=0 ps=0 
M2043 GND diff_7864_17452# diff_10564_18232# GND efet w=244 l=100
+ ad=0 pd=0 as=78736 ps=2800 
M2044 diff_16376_18520# diff_14176_18496# GND GND efet w=250 l=106
+ ad=13664 pd=600 as=0 ps=0 
M2045 diff_19228_20764# diff_19156_20272# Vdd GND efet w=40 l=424
+ ad=0 pd=0 as=0 ps=0 
M2046 diff_17600_19420# diff_3868_15448# diff_17452_19432# GND efet w=258 l=122
+ ad=42592 pd=1552 as=0 ps=0 
M2047 diff_17084_19288# diff_2140_4552# diff_16936_19336# GND efet w=258 l=110
+ ad=13664 pd=600 as=0 ps=0 
M2048 GND diff_3868_15448# diff_17084_19288# GND efet w=244 l=112
+ ad=0 pd=0 as=0 ps=0 
M2049 GND diff_2068_14080# diff_17600_19420# GND efet w=250 l=118
+ ad=0 pd=0 as=0 ps=0 
M2050 Vdd Vdd diff_18040_19532# GND efet w=52 l=556
+ ad=0 pd=0 as=98144 ps=4152 
M2051 diff_19156_20272# Vdd Vdd GND efet w=46 l=82
+ ad=3200 pd=240 as=0 ps=0 
M2052 Vdd Vdd diff_19900_20720# GND efet w=40 l=424
+ ad=0 pd=0 as=0 ps=0 
M2053 diff_18040_19532# clk2 diff_18040_19408# GND efet w=298 l=82
+ ad=0 pd=0 as=26000 ps=1424 
M2054 diff_18008_19060# diff_1840_19936# GND GND efet w=244 l=88
+ ad=105440 pd=2864 as=0 ps=0 
M2055 diff_18356_18196# diff_2104_10732# diff_17980_18148# GND efet w=690 l=134
+ ad=156352 pd=5616 as=155024 ps=5456 
M2056 diff_18008_19060# diff_2140_4552# GND GND efet w=292 l=122
+ ad=0 pd=0 as=0 ps=0 
M2057 GND diff_2140_5752# diff_17600_19420# GND efet w=238 l=106
+ ad=0 pd=0 as=0 ps=0 
M2058 GND diff_14176_18496# diff_15992_18424# GND efet w=244 l=100
+ ad=0 pd=0 as=0 ps=0 
M2059 diff_16532_18520# diff_12028_18580# diff_16376_18520# GND efet w=244 l=100
+ ad=0 pd=0 as=0 ps=0 
M2060 diff_16300_20812# clk2 diff_16532_18520# GND efet w=256 l=100
+ ad=29680 pd=1000 as=0 ps=0 
M2061 Vdd Vdd diff_16300_20812# GND efet w=58 l=550
+ ad=0 pd=0 as=0 ps=0 
M2062 diff_14872_18520# Vdd Vdd GND efet w=40 l=532
+ ad=0 pd=0 as=0 ps=0 
M2063 diff_18008_19060# diff_3868_15448# diff_18040_19408# GND efet w=270 l=122
+ ad=0 pd=0 as=0 ps=0 
M2064 GND diff_4192_12940# diff_17980_18148# GND efet w=706 l=94
+ ad=0 pd=0 as=0 ps=0 
M2065 Vdd Vdd diff_13816_22024# GND efet w=40 l=280
+ ad=0 pd=0 as=149280 ps=4920 
M2066 diff_13720_25264# diff_19228_20764# Vdd GND efet w=172 l=76
+ ad=0 pd=0 as=0 ps=0 
M2067 Vdd Vdd diff_20572_19796# GND efet w=70 l=538
+ ad=0 pd=0 as=22192 ps=856 
M2068 Vdd Vdd diff_18892_22660# GND efet w=58 l=202
+ ad=0 pd=0 as=53344 ps=1920 
M2069 diff_18892_22660# diff_20572_19796# GND GND efet w=304 l=112
+ ad=0 pd=0 as=0 ps=0 
M2070 GND diff_4192_12940# diff_19228_20764# GND efet w=126 l=98
+ ad=0 pd=0 as=0 ps=0 
M2071 diff_19228_20764# diff_19336_18748# GND GND efet w=106 l=82
+ ad=0 pd=0 as=0 ps=0 
M2072 diff_20572_19796# diff_2068_14080# diff_20572_19660# GND efet w=262 l=94
+ ad=0 pd=0 as=20048 ps=792 
M2073 GND diff_20116_18580# diff_13816_22024# GND efet w=198 l=122
+ ad=0 pd=0 as=0 ps=0 
M2074 diff_18976_18112# clk2 diff_18356_18196# GND efet w=112 l=100
+ ad=11504 pd=600 as=0 ps=0 
M2075 diff_20572_19660# clk2 diff_20656_19484# GND efet w=244 l=88
+ ad=0 pd=0 as=16592 ps=624 
M2076 diff_20656_19484# diff_3868_15448# GND GND efet w=244 l=88
+ ad=0 pd=0 as=0 ps=0 
M2077 diff_19688_18628# diff_2104_10732# GND GND efet w=250 l=94
+ ad=50288 pd=1808 as=0 ps=0 
M2078 diff_11848_16852# diff_7864_17452# GND GND efet w=436 l=88
+ ad=159952 pd=4184 as=0 ps=0 
M2079 diff_13672_16400# diff_7864_17452# diff_13252_16600# GND efet w=384 l=88
+ ad=172544 pd=4608 as=184416 ps=6456 
M2080 diff_14164_15040# diff_7864_17452# GND GND efet w=246 l=92
+ ad=174896 pd=6288 as=0 ps=0 
M2081 diff_14644_15824# diff_7864_17452# GND GND efet w=244 l=82
+ ad=155072 pd=6744 as=0 ps=0 
M2082 diff_14992_15292# diff_7864_17452# GND GND efet w=250 l=104
+ ad=149792 pd=6720 as=0 ps=0 
M2083 diff_5152_19192# diff_6676_17296# GND GND efet w=406 l=88
+ ad=200352 pd=6208 as=0 ps=0 
M2084 GND diff_6676_17296# diff_6904_14332# GND efet w=202 l=100
+ ad=0 pd=0 as=127168 ps=5368 
M2085 diff_5812_16768# diff_6676_17296# GND GND efet w=190 l=106
+ ad=64048 pd=1976 as=0 ps=0 
M2086 diff_5204_16384# Vdd Vdd GND efet w=46 l=286
+ ad=38320 pd=1872 as=0 ps=0 
M2087 diff_4408_17236# diff_4936_17224# diff_4408_17236# GND efet w=564 l=38
+ ad=0 pd=0 as=0 ps=0 
M2088 GND diff_4720_16588# diff_3868_15448# GND efet w=244 l=88
+ ad=0 pd=0 as=0 ps=0 
M2089 diff_4408_17236# diff_4720_16588# GND GND efet w=232 l=88
+ ad=0 pd=0 as=0 ps=0 
M2090 GND diff_6676_17296# diff_6556_14212# GND efet w=196 l=88
+ ad=0 pd=0 as=118768 ps=4720 
M2091 GND diff_6676_17296# diff_7384_14632# GND efet w=190 l=94
+ ad=0 pd=0 as=69840 ps=2280 
M2092 GND diff_6676_17296# diff_4456_18616# GND efet w=364 l=88
+ ad=0 pd=0 as=212880 ps=6184 
M2093 diff_4996_19156# diff_6676_17296# GND GND efet w=358 l=88
+ ad=228880 pd=6672 as=0 ps=0 
M2094 GND diff_6676_17296# diff_8920_12124# GND efet w=184 l=100
+ ad=0 pd=0 as=0 ps=0 
M2095 diff_6556_14212# diff_6976_17140# GND GND efet w=250 l=88
+ ad=0 pd=0 as=0 ps=0 
M2096 diff_7912_17540# diff_6976_17140# GND GND efet w=238 l=94
+ ad=0 pd=0 as=0 ps=0 
M2097 diff_8212_16444# diff_6976_17140# GND GND efet w=250 l=88
+ ad=0 pd=0 as=0 ps=0 
M2098 diff_4996_19156# diff_6976_17140# GND GND efet w=454 l=106
+ ad=0 pd=0 as=0 ps=0 
M2099 GND diff_6676_17296# diff_10792_18352# GND efet w=196 l=88
+ ad=0 pd=0 as=75088 ps=2536 
M2100 GND diff_6676_17296# diff_11548_16012# GND efet w=184 l=88
+ ad=0 pd=0 as=84464 ps=3008 
M2101 diff_15292_15896# diff_7864_17452# GND GND efet w=252 l=100
+ ad=151152 pd=6320 as=0 ps=0 
M2102 GND diff_1132_21544# diff_19688_18628# GND efet w=238 l=106
+ ad=0 pd=0 as=0 ps=0 
M2103 diff_19688_18628# diff_3868_15448# diff_19532_18580# GND efet w=278 l=106
+ ad=0 pd=0 as=17408 ps=736 
M2104 GND diff_16144_12496# diff_17980_18148# GND efet w=670 l=94
+ ad=0 pd=0 as=0 ps=0 
M2105 GND diff_1132_21544# diff_18356_18196# GND efet w=414 l=122
+ ad=0 pd=0 as=0 ps=0 
M2106 diff_18356_18196# diff_1840_19936# GND GND efet w=294 l=106
+ ad=0 pd=0 as=0 ps=0 
M2107 GND diff_18976_18112# diff_17896_9496# GND efet w=426 l=106
+ ad=0 pd=0 as=218160 ps=5816 
M2108 diff_17896_9496# diff_18976_18112# GND GND efet w=492 l=116
+ ad=0 pd=0 as=0 ps=0 
M2109 diff_19532_18580# clk2 diff_19336_18748# GND efet w=244 l=64
+ ad=0 pd=0 as=35216 ps=1536 
M2110 GND diff_1840_19936# diff_20740_18860# GND efet w=238 l=82
+ ad=0 pd=0 as=21920 ps=672 
M2111 diff_20740_18860# diff_3868_15448# diff_20740_18704# GND efet w=238 l=82
+ ad=0 pd=0 as=18992 ps=648 
M2112 diff_20348_18460# diff_2140_5752# diff_20116_18580# GND efet w=186 l=70
+ ad=12512 pd=504 as=23680 ps=1056 
M2113 GND diff_3868_15448# diff_20348_18460# GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M2114 diff_20740_18704# clk2 diff_20740_18548# GND efet w=244 l=76
+ ad=0 pd=0 as=22912 ps=960 
M2115 diff_18356_18196# Vdd Vdd GND efet w=56 l=300
+ ad=0 pd=0 as=0 ps=0 
M2116 Vdd Vdd diff_19336_18748# GND efet w=46 l=526
+ ad=0 pd=0 as=0 ps=0 
M2117 diff_12100_17968# diff_6676_17296# diff_11848_16852# GND efet w=388 l=100
+ ad=279456 pd=10344 as=0 ps=0 
M2118 diff_13252_16600# diff_6676_17296# GND GND efet w=322 l=106
+ ad=0 pd=0 as=0 ps=0 
M2119 GND diff_6976_17140# diff_9520_16492# GND efet w=754 l=82
+ ad=0 pd=0 as=156640 ps=3528 
M2120 diff_8920_12124# diff_6976_17140# GND GND efet w=244 l=98
+ ad=0 pd=0 as=0 ps=0 
M2121 diff_10564_18232# diff_6976_17140# GND GND efet w=244 l=94
+ ad=0 pd=0 as=0 ps=0 
M2122 diff_5816_16240# diff_5152_19192# diff_5600_16228# GND efet w=288 l=128
+ ad=99312 pd=3712 as=91584 ps=3032 
M2123 diff_5204_16384# clk1 diff_4720_16588# GND efet w=112 l=100
+ ad=0 pd=0 as=19712 ps=720 
M2124 diff_5600_16228# diff_5812_16768# diff_5816_16240# GND efet w=268 l=112
+ ad=0 pd=0 as=0 ps=0 
M2125 diff_10792_18352# diff_6976_17140# GND GND efet w=256 l=88
+ ad=0 pd=0 as=0 ps=0 
M2126 GND diff_6676_17296# diff_11884_18124# GND efet w=196 l=88
+ ad=0 pd=0 as=60704 ps=2320 
M2127 GND diff_6676_17296# diff_15592_16384# GND efet w=196 l=88
+ ad=0 pd=0 as=130256 ps=5424 
M2128 diff_11848_16852# diff_6976_17140# diff_12100_17968# GND efet w=460 l=88
+ ad=0 pd=0 as=0 ps=0 
M2129 diff_13252_16600# diff_6976_17140# GND GND efet w=376 l=110
+ ad=0 pd=0 as=0 ps=0 
M2130 diff_15292_15896# diff_6976_17140# GND GND efet w=262 l=94
+ ad=0 pd=0 as=0 ps=0 
M2131 diff_9520_16492# diff_6676_16900# diff_5152_19192# GND efet w=808 l=88
+ ad=0 pd=0 as=0 ps=0 
M2132 GND diff_6676_16900# diff_5812_16768# GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M2133 GND diff_6676_16900# diff_6904_14332# GND efet w=190 l=106
+ ad=0 pd=0 as=0 ps=0 
M2134 GND diff_6676_16900# diff_7384_14632# GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M2135 diff_15592_16384# diff_6976_17140# GND GND efet w=262 l=94
+ ad=0 pd=0 as=0 ps=0 
M2136 GND diff_6676_16900# diff_4456_18616# GND efet w=364 l=76
+ ad=0 pd=0 as=0 ps=0 
M2137 diff_5812_16768# diff_6676_16672# GND GND efet w=246 l=94
+ ad=0 pd=0 as=0 ps=0 
M2138 diff_6556_14212# diff_6676_16672# GND GND efet w=256 l=100
+ ad=0 pd=0 as=0 ps=0 
M2139 diff_7384_14632# diff_6676_16672# GND GND efet w=238 l=88
+ ad=0 pd=0 as=0 ps=0 
M2140 diff_7912_17540# diff_6676_16672# GND GND efet w=234 l=88
+ ad=0 pd=0 as=0 ps=0 
M2141 diff_8212_16444# diff_6676_16672# GND GND efet w=244 l=94
+ ad=0 pd=0 as=0 ps=0 
M2142 GND diff_6676_16900# diff_9784_10948# GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M2143 GND diff_6676_16900# diff_11548_16012# GND efet w=190 l=94
+ ad=0 pd=0 as=0 ps=0 
M2144 GND diff_6676_16900# diff_11848_16852# GND efet w=376 l=124
+ ad=0 pd=0 as=0 ps=0 
M2145 diff_6676_16900# diff_17332_16324# Vdd GND efet w=380 l=168
+ ad=89120 pd=2208 as=0 ps=0 
M2146 Vdd diff_17320_17404# diff_6976_17140# GND efet w=268 l=124
+ ad=0 pd=0 as=66992 ps=1776 
M2147 diff_13252_16600# diff_6676_16900# diff_13672_16400# GND efet w=328 l=100
+ ad=0 pd=0 as=0 ps=0 
M2148 diff_11884_18124# diff_6676_16900# GND GND efet w=202 l=94
+ ad=0 pd=0 as=0 ps=0 
M2149 diff_4456_18616# diff_6676_16672# GND GND efet w=436 l=88
+ ad=0 pd=0 as=0 ps=0 
M2150 diff_9784_10948# diff_6676_16672# GND GND efet w=244 l=98
+ ad=0 pd=0 as=0 ps=0 
M2151 diff_8920_12124# diff_6676_16672# GND GND efet w=234 l=82
+ ad=0 pd=0 as=0 ps=0 
M2152 diff_9520_16492# diff_6676_16672# GND GND efet w=730 l=100
+ ad=0 pd=0 as=0 ps=0 
M2153 GND diff_6676_16900# diff_14164_15040# GND efet w=196 l=88
+ ad=0 pd=0 as=0 ps=0 
M2154 GND diff_6676_16900# diff_14644_15824# GND efet w=184 l=94
+ ad=0 pd=0 as=0 ps=0 
M2155 GND diff_6676_16900# diff_14992_15292# GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M2156 diff_11848_16852# diff_6676_16672# diff_12100_17968# GND efet w=462 l=112
+ ad=0 pd=0 as=0 ps=0 
M2157 GND diff_6676_16672# diff_13252_16600# GND efet w=370 l=88
+ ad=0 pd=0 as=0 ps=0 
M2158 diff_5600_16228# diff_2392_18688# GND GND efet w=304 l=100
+ ad=0 pd=0 as=0 ps=0 
M2159 diff_4376_15940# Vdd Vdd GND efet w=58 l=526
+ ad=9280 pd=608 as=0 ps=0 
M2160 GND diff_5272_16192# diff_5204_16384# GND efet w=174 l=82
+ ad=0 pd=0 as=0 ps=0 
M2161 diff_5816_16240# diff_4996_19156# diff_5600_16228# GND efet w=256 l=100
+ ad=0 pd=0 as=0 ps=0 
M2162 diff_5132_15892# diff_3868_15448# diff_5816_16240# GND efet w=280 l=88
+ ad=89488 pd=3144 as=0 ps=0 
M2163 GND diff_7276_16504# diff_6904_14332# GND efet w=190 l=94
+ ad=0 pd=0 as=0 ps=0 
M2164 GND diff_7276_16504# diff_4996_19156# GND efet w=376 l=100
+ ad=0 pd=0 as=0 ps=0 
M2165 diff_11548_16012# diff_6676_16672# GND GND efet w=184 l=76
+ ad=0 pd=0 as=0 ps=0 
M2166 diff_9520_16492# diff_7276_16504# diff_5152_19192# GND efet w=790 l=112
+ ad=0 pd=0 as=0 ps=0 
M2167 diff_6556_14212# diff_6976_16348# GND GND efet w=252 l=100
+ ad=0 pd=0 as=0 ps=0 
M2168 GND diff_7276_16504# diff_10564_18232# GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M2169 GND diff_7276_16504# diff_10792_18352# GND efet w=208 l=88
+ ad=0 pd=0 as=0 ps=0 
M2170 diff_13672_16400# diff_6676_16672# diff_13252_16600# GND efet w=376 l=100
+ ad=0 pd=0 as=0 ps=0 
M2171 GND diff_6676_16672# diff_11884_18124# GND efet w=244 l=94
+ ad=0 pd=0 as=0 ps=0 
M2172 diff_14164_15040# diff_6676_16672# GND GND efet w=252 l=88
+ ad=0 pd=0 as=0 ps=0 
M2173 GND diff_17332_16324# diff_6976_17140# GND efet w=262 l=106
+ ad=0 pd=0 as=0 ps=0 
M2174 diff_6676_16900# diff_17320_17404# GND GND efet w=238 l=106
+ ad=0 pd=0 as=0 ps=0 
M2175 diff_17896_9496# Vdd Vdd GND efet w=76 l=112
+ ad=0 pd=0 as=0 ps=0 
M2176 diff_6676_17296# diff_18280_16804# Vdd GND efet w=312 l=116
+ ad=56864 pd=1696 as=0 ps=0 
M2177 Vdd diff_18220_17272# diff_7864_17452# GND efet w=160 l=112
+ ad=0 pd=0 as=76352 ps=1728 
M2178 diff_6676_17296# diff_18220_17272# GND GND efet w=238 l=118
+ ad=0 pd=0 as=0 ps=0 
M2179 GND diff_18280_16804# diff_7864_17452# GND efet w=160 l=88
+ ad=0 pd=0 as=0 ps=0 
M2180 Vdd Vdd diff_20116_18580# GND efet w=52 l=496
+ ad=0 pd=0 as=0 ps=0 
M2181 diff_20740_18548# Vdd Vdd GND efet w=46 l=514
+ ad=0 pd=0 as=0 ps=0 
M2182 GND diff_20740_18548# diff_20980_18032# GND efet w=298 l=70
+ ad=0 pd=0 as=23872 ps=1048 
M2183 diff_20980_18032# Vdd Vdd GND efet w=46 l=208
+ ad=0 pd=0 as=0 ps=0 
M2184 diff_3040_29500# diff_20980_18032# diff_19180_16528# GND efet w=88 l=94
+ ad=0 pd=0 as=17936 ps=656 
M2185 diff_3436_29560# diff_20980_18032# diff_19720_16504# GND efet w=82 l=88
+ ad=0 pd=0 as=17072 ps=680 
M2186 diff_16852_16108# Vdd Vdd GND efet w=64 l=244
+ ad=40288 pd=1624 as=0 ps=0 
M2187 diff_17320_17404# Vdd Vdd GND efet w=80 l=262
+ ad=32608 pd=1416 as=0 ps=0 
M2188 GND diff_19180_16528# diff_16852_16108# GND efet w=478 l=106
+ ad=0 pd=0 as=0 ps=0 
M2189 GND diff_20848_16804# diff_18220_17272# GND efet w=508 l=88
+ ad=0 pd=0 as=42256 ps=2072 
M2190 diff_3244_29488# diff_20980_18032# diff_20260_16504# GND efet w=82 l=94
+ ad=0 pd=0 as=17984 ps=672 
M2191 diff_17824_15484# Vdd Vdd GND efet w=94 l=232
+ ad=37840 pd=1680 as=0 ps=0 
M2192 GND diff_19720_16504# diff_17320_17404# GND efet w=502 l=94
+ ad=0 pd=0 as=0 ps=0 
M2193 GND diff_7276_16504# diff_14644_15824# GND efet w=190 l=82
+ ad=0 pd=0 as=0 ps=0 
M2194 GND diff_7276_16504# diff_14992_15292# GND efet w=190 l=82
+ ad=0 pd=0 as=0 ps=0 
M2195 diff_15292_15896# diff_7276_16504# GND GND efet w=190 l=94
+ ad=0 pd=0 as=0 ps=0 
M2196 diff_6904_14332# diff_6976_16348# GND GND efet w=246 l=94
+ ad=0 pd=0 as=0 ps=0 
M2197 diff_8212_16444# diff_6976_16348# GND GND efet w=244 l=94
+ ad=0 pd=0 as=0 ps=0 
M2198 diff_4456_18616# diff_6976_16348# GND GND efet w=424 l=82
+ ad=0 pd=0 as=0 ps=0 
M2199 GND diff_2392_18688# diff_4376_15940# GND efet w=94 l=94
+ ad=0 pd=0 as=0 ps=0 
M2200 diff_4976_15892# diff_4376_15940# GND GND efet w=172 l=88
+ ad=11696 pd=480 as=0 ps=0 
M2201 diff_5132_15892# diff_4720_16588# diff_4976_15892# GND efet w=172 l=88
+ ad=0 pd=0 as=0 ps=0 
M2202 diff_5272_16192# clk2 diff_5132_15892# GND efet w=64 l=88
+ ad=7424 pd=360 as=0 ps=0 
M2203 diff_5132_15892# Vdd diff_5132_15892# GND efet w=26 l=578
+ ad=0 pd=0 as=0 ps=0 
M2204 diff_9784_10948# diff_6976_16348# GND GND efet w=234 l=82
+ ad=0 pd=0 as=0 ps=0 
M2205 GND diff_6976_16348# diff_5152_19192# GND efet w=436 l=88
+ ad=0 pd=0 as=0 ps=0 
M2206 diff_10792_18352# diff_6976_16348# GND GND efet w=250 l=76
+ ad=0 pd=0 as=0 ps=0 
M2207 GND diff_7276_16504# diff_15592_16384# GND efet w=196 l=88
+ ad=0 pd=0 as=0 ps=0 
M2208 diff_13672_16400# diff_6976_16348# diff_13252_16600# GND efet w=420 l=100
+ ad=0 pd=0 as=0 ps=0 
M2209 diff_11548_16012# diff_6976_16348# GND GND efet w=190 l=94
+ ad=0 pd=0 as=0 ps=0 
M2210 diff_14644_15824# diff_6976_16348# GND GND efet w=246 l=94
+ ad=0 pd=0 as=0 ps=0 
M2211 diff_7576_16108# diff_16852_15544# Vdd GND efet w=156 l=140
+ ad=35168 pd=1584 as=0 ps=0 
M2212 Vdd diff_16852_16108# diff_6976_16348# GND efet w=318 l=176
+ ad=0 pd=0 as=46624 ps=1696 
M2213 GND diff_6604_14548# diff_5812_16768# GND efet w=172 l=112
+ ad=0 pd=0 as=0 ps=0 
M2214 GND diff_7576_16108# diff_7384_14632# GND efet w=202 l=118
+ ad=0 pd=0 as=0 ps=0 
M2215 GND diff_7576_16108# diff_7912_17540# GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M2216 Vdd Vdd diff_4360_13720# GND efet w=46 l=322
+ ad=0 pd=0 as=21216 ps=992 
M2217 Vdd Vdd diff_4192_12940# GND efet w=58 l=178
+ ad=0 pd=0 as=711584 ps=22680 
M2218 diff_4456_14788# Vdd Vdd GND efet w=76 l=226
+ ad=44752 pd=1512 as=0 ps=0 
M2219 diff_5812_16768# Vdd Vdd GND efet w=40 l=484
+ ad=0 pd=0 as=0 ps=0 
M2220 GND diff_7576_16108# diff_10564_18232# GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M2221 GND diff_7576_16108# diff_14164_15040# GND efet w=196 l=76
+ ad=0 pd=0 as=0 ps=0 
M2222 GND diff_7576_16108# diff_14992_15292# GND efet w=184 l=94
+ ad=0 pd=0 as=0 ps=0 
M2223 diff_6556_14212# Vdd Vdd GND efet w=52 l=520
+ ad=0 pd=0 as=0 ps=0 
M2224 diff_6904_14332# Vdd Vdd GND efet w=40 l=508
+ ad=0 pd=0 as=0 ps=0 
M2225 diff_7384_14632# Vdd Vdd GND efet w=40 l=514
+ ad=0 pd=0 as=0 ps=0 
M2226 diff_7912_17540# Vdd Vdd GND efet w=70 l=598
+ ad=0 pd=0 as=0 ps=0 
M2227 Vdd Vdd diff_8044_14476# GND efet w=52 l=592
+ ad=0 pd=0 as=12544 ps=576 
M2228 Vdd Vdd diff_8212_16444# GND efet w=52 l=460
+ ad=0 pd=0 as=0 ps=0 
M2229 diff_4456_18616# Vdd Vdd GND efet w=52 l=298
+ ad=0 pd=0 as=0 ps=0 
M2230 Vdd Vdd diff_8480_14848# GND efet w=52 l=412
+ ad=0 pd=0 as=14944 ps=744 
M2231 diff_4996_19156# Vdd Vdd GND efet w=64 l=316
+ ad=0 pd=0 as=0 ps=0 
M2232 diff_5152_19192# Vdd Vdd GND efet w=64 l=280
+ ad=0 pd=0 as=0 ps=0 
M2233 diff_8920_12124# Vdd Vdd GND efet w=52 l=448
+ ad=0 pd=0 as=0 ps=0 
M2234 Vdd Vdd diff_8896_12352# GND efet w=40 l=520
+ ad=0 pd=0 as=74224 ps=2464 
M2235 GND diff_6604_14548# diff_7472_14668# GND efet w=310 l=82
+ ad=0 pd=0 as=19040 ps=792 
M2236 diff_7472_14668# diff_7384_14632# diff_5704_12496# GND efet w=184 l=100
+ ad=0 pd=0 as=45680 ps=1928 
M2237 GND diff_3868_15448# diff_6136_14300# GND efet w=268 l=76
+ ad=0 pd=0 as=20240 ps=720 
M2238 diff_4360_13720# diff_2140_4552# GND GND efet w=142 l=94
+ ad=0 pd=0 as=0 ps=0 
M2239 GND reset diff_4120_13972# GND efet w=286 l=94
+ ad=0 pd=0 as=64240 ps=2088 
M2240 GND diff_5020_13900# diff_4456_14788# GND efet w=466 l=100
+ ad=0 pd=0 as=0 ps=0 
M2241 GND diff_4120_13972# diff_4360_13720# GND efet w=154 l=94
+ ad=0 pd=0 as=0 ps=0 
M2242 diff_4192_12940# diff_4120_13972# GND GND efet w=454 l=94
+ ad=0 pd=0 as=0 ps=0 
M2243 diff_5536_14200# diff_5020_13900# GND GND efet w=172 l=100
+ ad=16928 pd=744 as=0 ps=0 
M2244 diff_5584_14080# diff_2392_18688# GND GND efet w=106 l=94
+ ad=11872 pd=704 as=0 ps=0 
M2245 diff_6136_14300# diff_2392_18688# diff_6136_14144# GND efet w=274 l=82
+ ad=0 pd=0 as=19520 ps=648 
M2246 GND diff_7912_17540# diff_8044_14476# GND efet w=102 l=88
+ ad=0 pd=0 as=0 ps=0 
M2247 diff_8480_14848# diff_8212_16444# GND GND efet w=118 l=94
+ ad=0 pd=0 as=0 ps=0 
M2248 Vdd diff_8480_14848# diff_7744_12340# GND efet w=232 l=88
+ ad=0 pd=0 as=58384 ps=1776 
M2249 GND diff_7912_17540# diff_5512_12820# GND efet w=280 l=88
+ ad=0 pd=0 as=20768 ps=696 
M2250 diff_5512_12820# diff_8044_14476# Vdd GND efet w=106 l=94
+ ad=0 pd=0 as=0 ps=0 
M2251 GND diff_6556_14212# diff_6604_14020# GND efet w=100 l=88
+ ad=0 pd=0 as=25568 ps=792 
M2252 GND diff_6904_14332# diff_6844_13916# GND efet w=106 l=94
+ ad=0 pd=0 as=26032 ps=1240 
M2253 diff_7744_12340# diff_8212_16444# GND GND efet w=238 l=94
+ ad=0 pd=0 as=0 ps=0 
M2254 Vdd Vdd diff_7264_8080# GND efet w=52 l=436
+ ad=0 pd=0 as=173184 ps=6592 
M2255 Vdd Vdd diff_7504_8092# GND efet w=40 l=538
+ ad=0 pd=0 as=208688 ps=7072 
M2256 Vdd Vdd diff_7696_2656# GND efet w=64 l=352
+ ad=0 pd=0 as=142048 ps=4392 
M2257 Vdd Vdd diff_6712_8284# GND efet w=64 l=352
+ ad=0 pd=0 as=110800 ps=3040 
M2258 diff_9784_10948# Vdd Vdd GND efet w=40 l=466
+ ad=0 pd=0 as=0 ps=0 
M2259 diff_10564_18232# Vdd Vdd GND efet w=46 l=466
+ ad=0 pd=0 as=0 ps=0 
M2260 diff_10792_18352# Vdd Vdd GND efet w=52 l=448
+ ad=0 pd=0 as=0 ps=0 
M2261 diff_11548_16012# Vdd Vdd GND efet w=46 l=496
+ ad=0 pd=0 as=0 ps=0 
M2262 diff_12100_17968# Vdd Vdd GND efet w=76 l=532
+ ad=0 pd=0 as=0 ps=0 
M2263 Vdd Vdd diff_10648_11020# GND efet w=40 l=460
+ ad=0 pd=0 as=46880 ps=1544 
M2264 Vdd Vdd diff_11596_12508# GND efet w=52 l=448
+ ad=0 pd=0 as=86992 ps=3232 
M2265 diff_11380_10888# Vdd Vdd GND efet w=46 l=448
+ ad=71872 pd=2368 as=0 ps=0 
M2266 diff_12196_12148# Vdd Vdd GND efet w=46 l=454
+ ad=75952 pd=3088 as=0 ps=0 
M2267 Vdd Vdd diff_12496_12980# GND efet w=52 l=460
+ ad=0 pd=0 as=88400 ps=3176 
M2268 diff_12764_14728# Vdd Vdd GND efet w=40 l=502
+ ad=75696 pd=2848 as=0 ps=0 
M2269 diff_13672_16400# Vdd Vdd GND efet w=40 l=532
+ ad=0 pd=0 as=0 ps=0 
M2270 Vdd Vdd diff_14164_15040# GND efet w=46 l=550
+ ad=0 pd=0 as=0 ps=0 
M2271 diff_11884_18124# Vdd Vdd GND efet w=52 l=412
+ ad=0 pd=0 as=0 ps=0 
M2272 diff_10648_11020# diff_5512_12820# GND GND efet w=310 l=82
+ ad=0 pd=0 as=0 ps=0 
M2273 Vdd Vdd diff_13024_11248# GND efet w=52 l=436
+ ad=0 pd=0 as=82064 ps=2960 
M2274 Vdd Vdd diff_13372_12532# GND efet w=46 l=430
+ ad=0 pd=0 as=81184 ps=3088 
M2275 Vdd Vdd diff_13684_12616# GND efet w=40 l=460
+ ad=0 pd=0 as=76192 ps=2984 
M2276 Vdd Vdd diff_13960_12484# GND efet w=52 l=514
+ ad=0 pd=0 as=73376 ps=2912 
M2277 diff_14644_15824# Vdd Vdd GND efet w=52 l=496
+ ad=0 pd=0 as=0 ps=0 
M2278 diff_14992_15292# Vdd Vdd GND efet w=52 l=484
+ ad=0 pd=0 as=0 ps=0 
M2279 diff_15292_15896# Vdd Vdd GND efet w=58 l=478
+ ad=0 pd=0 as=0 ps=0 
M2280 diff_15592_16384# Vdd Vdd GND efet w=48 l=520
+ ad=0 pd=0 as=0 ps=0 
M2281 diff_14164_12076# Vdd Vdd GND efet w=58 l=532
+ ad=79904 pd=3480 as=0 ps=0 
M2282 Vdd Vdd diff_14572_12520# GND efet w=52 l=460
+ ad=0 pd=0 as=87424 ps=3328 
M2283 diff_14872_12968# Vdd Vdd GND efet w=40 l=460
+ ad=86896 pd=2728 as=0 ps=0 
M2284 diff_7576_16108# diff_16852_16108# GND GND efet w=162 l=98
+ ad=0 pd=0 as=0 ps=0 
M2285 GND diff_16852_15544# diff_6976_16348# GND efet w=234 l=94
+ ad=0 pd=0 as=0 ps=0 
M2286 diff_6676_16672# diff_17824_15484# Vdd GND efet w=306 l=128
+ ad=68624 pd=2376 as=0 ps=0 
M2287 Vdd diff_17824_16204# diff_7276_16504# GND efet w=196 l=100
+ ad=0 pd=0 as=49472 ps=1632 
M2288 diff_16852_15544# diff_16852_16108# GND GND efet w=220 l=88
+ ad=36544 pd=1560 as=0 ps=0 
M2289 diff_18220_17272# Vdd Vdd GND efet w=64 l=268
+ ad=0 pd=0 as=0 ps=0 
M2290 GND diff_20260_16504# diff_17824_15484# GND efet w=472 l=88
+ ad=0 pd=0 as=0 ps=0 
M2291 diff_17332_16324# diff_17320_17404# GND GND efet w=232 l=88
+ ad=61280 pd=2184 as=0 ps=0 
M2292 diff_17824_16204# diff_17824_15484# GND GND efet w=232 l=76
+ ad=42352 pd=1456 as=0 ps=0 
M2293 diff_3808_28348# diff_20980_18032# diff_20848_16804# GND efet w=76 l=94
+ ad=0 pd=0 as=17216 ps=632 
M2294 diff_18280_16804# diff_18220_17272# GND GND efet w=214 l=82
+ ad=38576 pd=1488 as=0 ps=0 
M2295 diff_16852_15544# diff_19000_15988# diff_16852_15544# GND efet w=26 l=422
+ ad=0 pd=0 as=0 ps=0 
M2296 diff_6676_16672# diff_17824_16204# GND GND efet w=270 l=104
+ ad=0 pd=0 as=0 ps=0 
M2297 GND diff_17824_15484# diff_7276_16504# GND efet w=196 l=88
+ ad=0 pd=0 as=0 ps=0 
M2298 diff_17332_16324# Vdd diff_17332_16324# GND efet w=32 l=432
+ ad=0 pd=0 as=0 ps=0 
M2299 diff_17824_16204# Vdd diff_17824_16204# GND efet w=26 l=350
+ ad=0 pd=0 as=0 ps=0 
M2300 diff_18280_16804# Vdd diff_18280_16804# GND efet w=20 l=414
+ ad=0 pd=0 as=0 ps=0 
M2301 diff_3808_28348# diff_16636_10928# diff_8212_13960# GND efet w=478 l=106
+ ad=0 pd=0 as=172064 ps=4792 
M2302 Vdd Vdd diff_16144_12496# GND efet w=82 l=334
+ ad=0 pd=0 as=132304 ps=3704 
M2303 diff_14572_12520# diff_5512_12820# GND GND efet w=256 l=100
+ ad=0 pd=0 as=0 ps=0 
M2304 diff_14872_12968# diff_5512_12820# GND GND efet w=256 l=98
+ ad=0 pd=0 as=0 ps=0 
M2305 Vdd Vdd diff_15940_9388# GND efet w=40 l=400
+ ad=0 pd=0 as=43568 ps=1544 
M2306 GND diff_7012_10588# diff_17852_14980# GND efet w=106 l=94
+ ad=0 pd=0 as=20032 ps=1008 
M2307 diff_17852_14980# Vdd Vdd GND efet w=52 l=554
+ ad=0 pd=0 as=0 ps=0 
M2308 diff_18364_14864# diff_17852_14980# diff_15940_9388# GND efet w=220 l=88
+ ad=13856 pd=576 as=0 ps=0 
M2309 diff_18032_14824# Vdd Vdd GND efet w=52 l=634
+ ad=13888 pd=744 as=0 ps=0 
M2310 diff_18364_14864# diff_18032_14824# GND GND efet w=214 l=82
+ ad=0 pd=0 as=0 ps=0 
M2311 diff_18032_14824# diff_16144_12496# GND GND efet w=94 l=76
+ ad=0 pd=0 as=0 ps=0 
M2312 diff_5536_14200# diff_5584_14080# diff_5644_14008# GND efet w=160 l=88
+ ad=0 pd=0 as=47056 ps=1560 
M2313 diff_6136_14144# diff_6076_14080# diff_5644_14008# GND efet w=244 l=76
+ ad=0 pd=0 as=0 ps=0 
M2314 diff_2996_13528# clk2 GND GND efet w=208 l=88
+ ad=89520 pd=3408 as=0 ps=0 
M2315 diff_2996_13528# diff_3076_13504# diff_2996_13528# GND efet w=606 l=38
+ ad=0 pd=0 as=0 ps=0 
M2316 Vdd diff_3076_13504# diff_2996_13528# GND efet w=58 l=262
+ ad=0 pd=0 as=0 ps=0 
M2317 diff_2212_11356# clk2 diff_2608_13384# GND efet w=106 l=94
+ ad=394704 pd=11624 as=8768 ps=480 
M2318 Vdd Vdd diff_3076_13504# GND efet w=40 l=100
+ ad=0 pd=0 as=3008 ps=240 
M2319 diff_928_20116# diff_2996_13528# diff_2752_13076# GND efet w=220 l=88
+ ad=280736 pd=10432 as=70080 ps=2368 
M2320 diff_2752_13076# diff_2608_13384# GND GND efet w=508 l=100
+ ad=0 pd=0 as=0 ps=0 
M2321 Vdd Vdd diff_2752_13076# GND efet w=58 l=166
+ ad=0 pd=0 as=0 ps=0 
M2322 diff_2752_13076# clk1 diff_2428_12196# GND efet w=88 l=88
+ ad=0 pd=0 as=8432 ps=440 
M2323 GND diff_4360_13720# diff_4120_13972# GND efet w=268 l=88
+ ad=0 pd=0 as=0 ps=0 
M2324 diff_5240_13720# clk1 diff_5020_13900# GND efet w=112 l=88
+ ad=26368 pd=960 as=13664 ps=576 
M2325 GND diff_5308_13696# diff_5240_13720# GND efet w=214 l=94
+ ad=0 pd=0 as=0 ps=0 
M2326 diff_5644_14008# clk2 diff_5308_13696# GND efet w=64 l=88
+ ad=0 pd=0 as=9056 ps=528 
M2327 Vdd Vdd diff_5584_14080# GND efet w=52 l=688
+ ad=0 pd=0 as=0 ps=0 
M2328 GND test diff_4300_13492# GND efet w=292 l=76
+ ad=0 pd=0 as=94944 ps=3448 
M2329 Vdd Vdd diff_4300_13492# GND efet w=35 l=464
+ ad=0 pd=0 as=0 ps=0 
M2330 diff_4120_13972# Vdd Vdd GND efet w=40 l=208
+ ad=0 pd=0 as=0 ps=0 
M2331 Vdd Vdd diff_5240_13720# GND efet w=52 l=292
+ ad=0 pd=0 as=0 ps=0 
M2332 Vdd Vdd diff_4636_12124# GND efet w=40 l=412
+ ad=0 pd=0 as=21376 ps=1048 
M2333 diff_2780_12500# diff_2428_12196# GND GND efet w=256 l=82
+ ad=79248 pd=2968 as=0 ps=0 
M2334 Vdd Vdd diff_5116_11728# GND efet w=64 l=160
+ ad=0 pd=0 as=124304 ps=3784 
M2335 diff_5644_14008# Vdd Vdd GND efet w=46 l=514
+ ad=0 pd=0 as=0 ps=0 
M2336 GND diff_5512_12820# diff_5116_11728# GND efet w=484 l=88
+ ad=0 pd=0 as=0 ps=0 
M2337 diff_6604_14020# Vdd Vdd GND efet w=82 l=538
+ ad=0 pd=0 as=0 ps=0 
M2338 GND diff_6844_13916# diff_7060_14084# GND efet w=184 l=88
+ ad=0 pd=0 as=140720 ps=5440 
M2339 GND diff_7744_12340# diff_8896_12352# GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M2340 diff_7264_8080# diff_7744_12340# GND GND efet w=184 l=94
+ ad=0 pd=0 as=0 ps=0 
M2341 GND diff_7744_12340# diff_7504_8092# GND efet w=190 l=94
+ ad=0 pd=0 as=0 ps=0 
M2342 GND diff_7744_12340# diff_7696_2656# GND efet w=310 l=82
+ ad=0 pd=0 as=0 ps=0 
M2343 GND diff_7744_12340# diff_6712_8284# GND efet w=274 l=94
+ ad=0 pd=0 as=0 ps=0 
M2344 diff_11596_12508# diff_7744_12340# GND GND efet w=190 l=82
+ ad=0 pd=0 as=0 ps=0 
M2345 GND diff_7744_12340# diff_11380_10888# GND efet w=190 l=82
+ ad=0 pd=0 as=0 ps=0 
M2346 GND diff_7744_12340# diff_12196_12148# GND efet w=202 l=82
+ ad=0 pd=0 as=0 ps=0 
M2347 diff_7744_14056# diff_7588_13816# diff_7060_14084# GND efet w=358 l=118
+ ad=77520 pd=2752 as=0 ps=0 
M2348 diff_7060_14084# diff_6604_14020# diff_6076_14080# GND efet w=334 l=106
+ ad=0 pd=0 as=56992 ps=1536 
M2349 diff_6844_13916# Vdd Vdd GND efet w=40 l=472
+ ad=0 pd=0 as=0 ps=0 
M2350 diff_7060_14084# diff_7216_13264# diff_6076_14080# GND efet w=382 l=100
+ ad=0 pd=0 as=0 ps=0 
M2351 diff_6076_14080# Vdd Vdd GND efet w=40 l=406
+ ad=0 pd=0 as=0 ps=0 
M2352 Vdd Vdd diff_5704_12496# GND efet w=40 l=562
+ ad=0 pd=0 as=0 ps=0 
M2353 Vdd Vdd diff_6472_12712# GND efet w=46 l=208
+ ad=0 pd=0 as=46912 ps=2064 
M2354 diff_7060_14084# diff_8212_14116# diff_7744_14056# GND efet w=520 l=100
+ ad=0 pd=0 as=0 ps=0 
M2355 diff_8896_12352# diff_8212_14116# GND GND efet w=244 l=82
+ ad=0 pd=0 as=0 ps=0 
M2356 diff_7504_8092# diff_8212_14116# GND GND efet w=240 l=88
+ ad=0 pd=0 as=0 ps=0 
M2357 diff_7696_2656# diff_8212_14116# GND GND efet w=328 l=88
+ ad=0 pd=0 as=0 ps=0 
M2358 diff_6712_8284# diff_8212_14116# GND GND efet w=328 l=106
+ ad=0 pd=0 as=0 ps=0 
M2359 diff_7744_14056# diff_7720_13960# GND GND efet w=408 l=112
+ ad=0 pd=0 as=0 ps=0 
M2360 GND diff_8212_13960# diff_7744_14056# GND efet w=616 l=100
+ ad=0 pd=0 as=0 ps=0 
M2361 GND diff_7744_12340# diff_12496_12980# GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M2362 diff_12764_14728# diff_7744_12340# GND GND efet w=190 l=94
+ ad=0 pd=0 as=0 ps=0 
M2363 GND diff_7744_12340# diff_13024_11248# GND efet w=190 l=94
+ ad=0 pd=0 as=0 ps=0 
M2364 GND diff_7744_12340# diff_13372_12532# GND efet w=184 l=100
+ ad=0 pd=0 as=0 ps=0 
M2365 GND diff_7744_12340# diff_13684_12616# GND efet w=190 l=94
+ ad=0 pd=0 as=0 ps=0 
M2366 GND diff_5512_12820# diff_16144_12496# GND efet w=322 l=82
+ ad=0 pd=0 as=0 ps=0 
M2367 diff_15940_9388# diff_2140_4552# diff_16900_14392# GND efet w=252 l=92
+ ad=0 pd=0 as=23744 ps=840 
M2368 diff_3436_29560# diff_16636_10928# diff_8512_13708# GND efet w=502 l=130
+ ad=0 pd=0 as=142400 ps=4672 
M2369 GND diff_7744_12340# diff_13960_12484# GND efet w=184 l=76
+ ad=0 pd=0 as=0 ps=0 
M2370 diff_14164_12076# diff_7744_12340# GND GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M2371 GND diff_16144_12496# diff_16900_14392# GND efet w=254 l=114
+ ad=0 pd=0 as=0 ps=0 
M2372 diff_12764_14728# diff_8212_14116# GND GND efet w=250 l=100
+ ad=0 pd=0 as=0 ps=0 
M2373 diff_13372_12532# diff_8212_14116# GND GND efet w=244 l=86
+ ad=0 pd=0 as=0 ps=0 
M2374 diff_14572_12520# diff_8212_14116# GND GND efet w=262 l=88
+ ad=0 pd=0 as=0 ps=0 
M2375 diff_14872_12968# diff_8212_14116# GND GND efet w=244 l=110
+ ad=0 pd=0 as=0 ps=0 
M2376 diff_16144_12496# diff_8212_14116# GND GND efet w=364 l=88
+ ad=0 pd=0 as=0 ps=0 
M2377 GND diff_17252_11776# diff_8212_14116# GND efet w=238 l=88
+ ad=0 pd=0 as=51664 ps=2016 
M2378 diff_8212_13960# diff_17140_11656# GND GND efet w=466 l=94
+ ad=0 pd=0 as=0 ps=0 
M2379 GND diff_8212_13960# diff_7264_8080# GND efet w=184 l=94
+ ad=0 pd=0 as=0 ps=0 
M2380 GND diff_8212_13960# diff_10648_11020# GND efet w=256 l=76
+ ad=0 pd=0 as=0 ps=0 
M2381 GND diff_8212_13960# diff_11596_12508# GND efet w=196 l=76
+ ad=0 pd=0 as=0 ps=0 
M2382 GND diff_8212_13960# diff_11380_10888# GND efet w=190 l=82
+ ad=0 pd=0 as=0 ps=0 
M2383 GND diff_8212_13960# diff_12196_12148# GND efet w=184 l=76
+ ad=0 pd=0 as=0 ps=0 
M2384 GND diff_8212_13960# diff_12496_12980# GND efet w=184 l=76
+ ad=0 pd=0 as=0 ps=0 
M2385 GND diff_8212_13960# diff_13024_11248# GND efet w=196 l=88
+ ad=0 pd=0 as=0 ps=0 
M2386 GND diff_8212_13960# diff_13684_12616# GND efet w=190 l=82
+ ad=0 pd=0 as=0 ps=0 
M2387 GND diff_7720_13960# diff_7588_13816# GND efet w=100 l=88
+ ad=0 pd=0 as=20128 ps=1056 
M2388 diff_8896_12352# diff_8944_13720# GND GND efet w=244 l=82
+ ad=0 pd=0 as=0 ps=0 
M2389 GND diff_8512_13708# diff_8408_13540# GND efet w=364 l=112
+ ad=0 pd=0 as=37808 ps=1240 
M2390 diff_8408_13540# diff_7660_12052# diff_7720_13960# GND efet w=232 l=82
+ ad=0 pd=0 as=92336 ps=3272 
M2391 diff_7588_13816# Vdd Vdd GND efet w=40 l=412
+ ad=0 pd=0 as=0 ps=0 
M2392 diff_7504_8092# diff_8944_13720# GND GND efet w=244 l=82
+ ad=0 pd=0 as=0 ps=0 
M2393 diff_11596_12508# diff_8944_13720# GND GND efet w=256 l=94
+ ad=0 pd=0 as=0 ps=0 
M2394 diff_11380_10888# diff_8944_13720# GND GND efet w=246 l=100
+ ad=0 pd=0 as=0 ps=0 
M2395 diff_12196_12148# diff_8944_13720# GND GND efet w=240 l=88
+ ad=0 pd=0 as=0 ps=0 
M2396 diff_12496_12980# diff_8944_13720# GND GND efet w=250 l=92
+ ad=0 pd=0 as=0 ps=0 
M2397 GND diff_8212_13960# diff_13960_12484# GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M2398 GND diff_8212_13960# diff_14164_12076# GND efet w=196 l=88
+ ad=0 pd=0 as=0 ps=0 
M2399 GND diff_18332_11776# diff_8944_13720# GND efet w=294 l=122
+ ad=0 pd=0 as=52448 ps=1856 
M2400 diff_8512_13708# diff_18232_11632# GND GND efet w=442 l=128
+ ad=0 pd=0 as=0 ps=0 
M2401 diff_7720_13960# Vdd Vdd GND efet w=40 l=388
+ ad=0 pd=0 as=0 ps=0 
M2402 GND diff_8512_13708# diff_7696_2656# GND efet w=274 l=106
+ ad=0 pd=0 as=0 ps=0 
M2403 GND diff_8512_13708# diff_6712_8284# GND efet w=280 l=88
+ ad=0 pd=0 as=0 ps=0 
M2404 Vdd diff_17140_11656# diff_8212_14116# GND efet w=178 l=82
+ ad=0 pd=0 as=0 ps=0 
M2405 diff_8212_13960# diff_17252_11776# Vdd GND efet w=202 l=70
+ ad=0 pd=0 as=0 ps=0 
M2406 GND diff_8512_13708# diff_12764_14728# GND efet w=184 l=76
+ ad=0 pd=0 as=0 ps=0 
M2407 GND diff_8512_13708# diff_13024_11248# GND efet w=196 l=76
+ ad=0 pd=0 as=0 ps=0 
M2408 GND diff_8512_13708# diff_13372_12532# GND efet w=190 l=88
+ ad=0 pd=0 as=0 ps=0 
M2409 GND diff_8512_13708# diff_13684_12616# GND efet w=220 l=76
+ ad=0 pd=0 as=0 ps=0 
M2410 GND diff_8512_13708# diff_13960_12484# GND efet w=220 l=76
+ ad=0 pd=0 as=0 ps=0 
M2411 GND diff_8512_13708# diff_14164_12076# GND efet w=184 l=100
+ ad=0 pd=0 as=0 ps=0 
M2412 GND clk2 diff_6472_12712# GND efet w=388 l=76
+ ad=0 pd=0 as=0 ps=0 
M2413 Vdd Vdd diff_5792_12544# GND efet w=46 l=550
+ ad=0 pd=0 as=22912 ps=1152 
M2414 diff_2780_12500# diff_2860_12400# diff_2780_12500# GND efet w=588 l=44
+ ad=0 pd=0 as=0 ps=0 
M2415 Vdd diff_2860_12400# diff_2780_12500# GND efet w=46 l=214
+ ad=0 pd=0 as=0 ps=0 
M2416 Vdd Vdd diff_2860_12400# GND efet w=40 l=100
+ ad=0 pd=0 as=3248 ps=288 
M2417 diff_2392_18688# diff_2428_12196# GND GND efet w=256 l=88
+ ad=412416 pd=10336 as=0 ps=0 
M2418 diff_4636_12124# diff_4120_12124# GND GND efet w=112 l=88
+ ad=0 pd=0 as=0 ps=0 
M2419 diff_7100_12928# clk2 diff_2140_5752# GND efet w=64 l=88
+ ad=4784 pd=288 as=869584 ps=24424 
M2420 diff_5792_12544# diff_5704_12496# GND GND efet w=100 l=100
+ ad=0 pd=0 as=0 ps=0 
M2421 Vdd diff_2780_12500# diff_2392_18688# GND efet w=292 l=94
+ ad=0 pd=0 as=0 ps=0 
M2422 diff_4096_2464# diff_4120_12124# Vdd GND efet w=160 l=88
+ ad=77008 pd=2904 as=0 ps=0 
M2423 diff_7004_12508# diff_7100_12928# GND GND efet w=112 l=88
+ ad=29296 pd=1312 as=0 ps=0 
M2424 diff_7004_12508# diff_6472_12712# diff_6712_12448# GND efet w=64 l=100
+ ad=0 pd=0 as=11072 ps=560 
M2425 Vdd Vdd diff_7420_13000# GND efet w=46 l=88
+ ad=0 pd=0 as=19376 ps=888 
M2426 Vdd diff_7420_13000# diff_7516_12484# GND efet w=40 l=130
+ ad=0 pd=0 as=364368 ps=11824 
M2427 diff_7516_12484# diff_7420_13000# diff_7516_12484# GND efet w=568 l=214
+ ad=0 pd=0 as=0 ps=0 
M2428 diff_8396_13108# diff_5524_8116# diff_7720_13960# GND efet w=220 l=88
+ ad=30560 pd=1312 as=0 ps=0 
M2429 diff_6712_8284# diff_10204_13336# GND GND efet w=352 l=82
+ ad=0 pd=0 as=0 ps=0 
M2430 diff_11596_12508# diff_10204_13336# GND GND efet w=250 l=76
+ ad=0 pd=0 as=0 ps=0 
M2431 diff_12496_12980# diff_10204_13336# GND GND efet w=240 l=88
+ ad=0 pd=0 as=0 ps=0 
M2432 GND diff_8500_13252# diff_8396_13108# GND efet w=370 l=100
+ ad=0 pd=0 as=0 ps=0 
M2433 diff_12764_14728# diff_10204_13336# GND GND efet w=256 l=88
+ ad=0 pd=0 as=0 ps=0 
M2434 diff_13024_11248# diff_10204_13336# GND GND efet w=250 l=94
+ ad=0 pd=0 as=0 ps=0 
M2435 diff_13684_12616# diff_10204_13336# GND GND efet w=252 l=88
+ ad=0 pd=0 as=0 ps=0 
M2436 GND diff_8512_13708# diff_14572_12520# GND efet w=226 l=82
+ ad=0 pd=0 as=0 ps=0 
M2437 GND diff_8512_13708# diff_14872_12968# GND efet w=208 l=88
+ ad=0 pd=0 as=0 ps=0 
M2438 diff_14872_12968# diff_10204_13336# GND GND efet w=238 l=94
+ ad=0 pd=0 as=0 ps=0 
M2439 GND diff_4636_12124# diff_4096_2464# GND efet w=160 l=88
+ ad=0 pd=0 as=0 ps=0 
M2440 diff_5216_12100# diff_4360_8920# diff_4120_12124# GND efet w=244 l=76
+ ad=14960 pd=576 as=81632 ps=2864 
M2441 GND diff_5116_11728# diff_5216_12100# GND efet w=220 l=88
+ ad=0 pd=0 as=0 ps=0 
M2442 diff_5600_12100# diff_4576_11152# GND GND efet w=220 l=88
+ ad=35360 pd=1296 as=0 ps=0 
M2443 diff_4120_12124# diff_5792_12544# diff_5600_12100# GND efet w=238 l=94
+ ad=0 pd=0 as=0 ps=0 
M2444 GND diff_6076_12268# diff_4120_12124# GND efet w=118 l=94
+ ad=0 pd=0 as=0 ps=0 
M2445 GND clk2 diff_6508_12124# GND efet w=130 l=94
+ ad=0 pd=0 as=54528 ps=2576 
M2446 diff_6076_12268# diff_6712_12448# GND GND efet w=160 l=94
+ ad=18800 pd=768 as=0 ps=0 
M2447 Vdd Vdd diff_6076_12268# GND efet w=58 l=448
+ ad=0 pd=0 as=0 ps=0 
M2448 Vdd diff_2780_11284# diff_2212_11356# GND efet w=316 l=100
+ ad=0 pd=0 as=0 ps=0 
M2449 diff_2212_11356# diff_2404_11752# GND GND efet w=298 l=94
+ ad=0 pd=0 as=0 ps=0 
M2450 GND diff_2212_11356# diff_2068_11368# GND efet w=202 l=106
+ ad=0 pd=0 as=147200 ps=5288 
M2451 diff_2780_11284# diff_2860_11344# diff_2780_11284# GND efet w=570 l=44
+ ad=81120 pd=2832 as=0 ps=0 
M2452 diff_2780_11284# diff_2404_11752# GND GND efet w=244 l=88
+ ad=0 pd=0 as=0 ps=0 
M2453 Vdd Vdd diff_2860_11344# GND efet w=46 l=106
+ ad=0 pd=0 as=2384 ps=216 
M2454 Vdd diff_2860_11344# diff_2780_11284# GND efet w=52 l=220
+ ad=0 pd=0 as=0 ps=0 
M2455 diff_3028_10888# diff_2792_10864# GND GND efet w=214 l=82
+ ad=44848 pd=1752 as=0 ps=0 
M2456 diff_2792_10864# clk2 diff_2104_10732# GND efet w=100 l=106
+ ad=10880 pd=488 as=653008 ps=19936 
M2457 diff_2404_11752# clk1 diff_3028_10888# GND efet w=112 l=88
+ ad=10064 pd=488 as=0 ps=0 
M2458 Vdd Vdd diff_3028_10888# GND efet w=64 l=304
+ ad=0 pd=0 as=0 ps=0 
M2459 diff_6344_12028# diff_2212_11356# GND GND efet w=112 l=88
+ ad=16480 pd=808 as=0 ps=0 
M2460 diff_4120_12124# diff_5476_11636# diff_4120_12124# GND efet w=132 l=476
+ ad=0 pd=0 as=0 ps=0 
M2461 diff_2068_11368# diff_2104_10732# GND GND efet w=172 l=106
+ ad=0 pd=0 as=0 ps=0 
M2462 Vdd diff_2780_10084# diff_2104_10732# GND efet w=286 l=94
+ ad=0 pd=0 as=0 ps=0 
M2463 diff_2104_10732# diff_2416_10540# GND GND efet w=298 l=94
+ ad=0 pd=0 as=0 ps=0 
M2464 diff_2780_10084# diff_2860_10156# diff_2780_10084# GND efet w=612 l=44
+ ad=78336 pd=3024 as=0 ps=0 
M2465 diff_2780_10084# diff_2416_10540# GND GND efet w=208 l=82
+ ad=0 pd=0 as=0 ps=0 
M2466 Vdd Vdd diff_2860_10156# GND efet w=40 l=88
+ ad=0 pd=0 as=3008 ps=240 
M2467 Vdd diff_2860_10156# diff_2780_10084# GND efet w=58 l=214
+ ad=0 pd=0 as=0 ps=0 
M2468 Vdd diff_5476_11636# diff_4120_12124# GND efet w=40 l=322
+ ad=0 pd=0 as=0 ps=0 
M2469 diff_6512_11944# clk2 diff_6344_12028# GND efet w=64 l=88
+ ad=3872 pd=264 as=0 ps=0 
M2470 diff_7004_12508# Vdd Vdd GND efet w=40 l=400
+ ad=0 pd=0 as=0 ps=0 
M2471 GND diff_8500_13252# diff_8896_12352# GND efet w=196 l=100
+ ad=0 pd=0 as=0 ps=0 
M2472 GND diff_8500_13252# diff_7504_8092# GND efet w=232 l=88
+ ad=0 pd=0 as=0 ps=0 
M2473 GND diff_8500_13252# diff_7696_2656# GND efet w=268 l=88
+ ad=0 pd=0 as=0 ps=0 
M2474 GND diff_8500_13252# diff_11380_10888# GND efet w=190 l=94
+ ad=0 pd=0 as=0 ps=0 
M2475 GND diff_8500_13252# diff_12196_12148# GND efet w=196 l=82
+ ad=0 pd=0 as=0 ps=0 
M2476 GND diff_8500_13252# diff_13372_12532# GND efet w=184 l=76
+ ad=0 pd=0 as=0 ps=0 
M2477 GND diff_8500_13252# diff_13960_12484# GND efet w=184 l=76
+ ad=0 pd=0 as=0 ps=0 
M2478 GND diff_8500_13252# diff_14164_12076# GND efet w=196 l=100
+ ad=0 pd=0 as=0 ps=0 
M2479 GND diff_8500_13252# diff_14572_12520# GND efet w=190 l=100
+ ad=0 pd=0 as=0 ps=0 
M2480 diff_8672_12820# diff_4300_13492# diff_7720_13960# GND efet w=220 l=88
+ ad=36224 pd=1376 as=0 ps=0 
M2481 GND diff_6604_14548# diff_8672_12820# GND efet w=400 l=112
+ ad=0 pd=0 as=0 ps=0 
M2482 diff_8896_12352# diff_8944_12928# GND GND efet w=240 l=88
+ ad=0 pd=0 as=0 ps=0 
M2483 diff_7696_2656# diff_8944_12928# GND GND efet w=340 l=82
+ ad=0 pd=0 as=0 ps=0 
M2484 diff_6712_8284# diff_8944_12928# GND GND efet w=334 l=88
+ ad=0 pd=0 as=0 ps=0 
M2485 diff_11380_10888# diff_8944_12928# GND GND efet w=246 l=106
+ ad=0 pd=0 as=0 ps=0 
M2486 diff_12496_12980# diff_8944_12928# GND GND efet w=244 l=88
+ ad=0 pd=0 as=0 ps=0 
M2487 diff_13024_11248# diff_8944_12928# GND GND efet w=256 l=88
+ ad=0 pd=0 as=0 ps=0 
M2488 diff_13960_12484# diff_8944_12928# GND GND efet w=250 l=76
+ ad=0 pd=0 as=0 ps=0 
M2489 diff_14872_12968# diff_8944_12928# GND GND efet w=238 l=88
+ ad=0 pd=0 as=0 ps=0 
M2490 GND diff_6604_14548# diff_7504_8092# GND efet w=196 l=76
+ ad=0 pd=0 as=0 ps=0 
M2491 GND diff_6604_14548# diff_11596_12508# GND efet w=196 l=88
+ ad=0 pd=0 as=0 ps=0 
M2492 GND diff_6604_14548# diff_13372_12532# GND efet w=208 l=100
+ ad=0 pd=0 as=0 ps=0 
M2493 GND diff_6604_14548# diff_12196_12148# GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M2494 GND diff_6604_14548# diff_12764_14728# GND efet w=184 l=82
+ ad=0 pd=0 as=0 ps=0 
M2495 GND diff_6604_14548# diff_13684_12616# GND efet w=184 l=76
+ ad=0 pd=0 as=0 ps=0 
M2496 GND diff_6604_14548# diff_14164_12076# GND efet w=196 l=88
+ ad=0 pd=0 as=0 ps=0 
M2497 GND diff_6604_14548# diff_14572_12520# GND efet w=196 l=76
+ ad=0 pd=0 as=0 ps=0 
M2498 GND diff_7744_12340# diff_7516_12484# GND efet w=358 l=82
+ ad=0 pd=0 as=0 ps=0 
M2499 GND diff_8416_12352# diff_4432_7336# GND efet w=178 l=82
+ ad=0 pd=0 as=232848 ps=6888 
M2500 diff_4432_7336# diff_5912_10948# GND GND efet w=160 l=88
+ ad=0 pd=0 as=0 ps=0 
M2501 diff_8416_12352# diff_8896_12352# GND GND efet w=112 l=76
+ ad=19120 pd=1056 as=0 ps=0 
M2502 diff_9884_12392# diff_7504_8092# GND GND efet w=112 l=76
+ ad=220080 pd=9376 as=0 ps=0 
M2503 GND diff_5912_10948# diff_7516_12484# GND efet w=358 l=82
+ ad=0 pd=0 as=0 ps=0 
M2504 diff_6508_12124# diff_6512_11944# GND GND efet w=172 l=106
+ ad=0 pd=0 as=0 ps=0 
M2505 Vdd Vdd diff_6344_12028# GND efet w=40 l=388
+ ad=0 pd=0 as=0 ps=0 
M2506 diff_5476_11636# Vdd Vdd GND efet w=40 l=88
+ ad=7184 pd=456 as=0 ps=0 
M2507 Vdd Vdd diff_7012_10588# GND efet w=40 l=124
+ ad=0 pd=0 as=115280 ps=4096 
M2508 diff_8416_12352# Vdd Vdd GND efet w=46 l=526
+ ad=0 pd=0 as=0 ps=0 
M2509 GND diff_7696_2656# diff_9884_12392# GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M2510 diff_9884_12392# diff_6712_8284# GND GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M2511 Vdd Vdd diff_5912_10948# GND efet w=46 l=148
+ ad=0 pd=0 as=93936 ps=2776 
M2512 diff_7012_10588# diff_6508_12124# GND GND efet w=532 l=88
+ ad=0 pd=0 as=0 ps=0 
M2513 diff_4952_10516# Vdd Vdd GND efet w=40 l=460
+ ad=28912 pd=1576 as=0 ps=0 
M2514 Vdd Vdd diff_5420_10876# GND efet w=40 l=232
+ ad=0 pd=0 as=58512 ps=2288 
M2515 diff_6508_12124# Vdd Vdd GND efet w=40 l=292
+ ad=0 pd=0 as=0 ps=0 
M2516 Vdd Vdd diff_6076_10456# GND efet w=46 l=526
+ ad=0 pd=0 as=56736 ps=2704 
M2517 diff_3028_9676# diff_2792_9668# GND GND efet w=214 l=82
+ ad=44752 pd=1680 as=0 ps=0 
M2518 diff_2792_9668# clk2 diff_2068_14080# GND efet w=124 l=88
+ ad=11936 pd=488 as=195664 ps=5320 
M2519 diff_2416_10540# clk1 diff_3028_9676# GND efet w=112 l=88
+ ad=11168 pd=488 as=0 ps=0 
M2520 Vdd Vdd diff_3028_9676# GND efet w=52 l=244
+ ad=0 pd=0 as=0 ps=0 
M2521 diff_5420_10876# diff_5108_10516# GND GND efet w=280 l=94
+ ad=0 pd=0 as=0 ps=0 
M2522 GND clk2 diff_5420_10876# GND efet w=226 l=94
+ ad=0 pd=0 as=0 ps=0 
M2523 diff_5912_10948# diff_5420_10876# GND GND efet w=436 l=88
+ ad=0 pd=0 as=0 ps=0 
M2524 GND diff_5116_11728# diff_6076_10456# GND efet w=106 l=94
+ ad=0 pd=0 as=0 ps=0 
M2525 diff_6076_10456# diff_4192_12940# GND GND efet w=88 l=88
+ ad=0 pd=0 as=0 ps=0 
M2526 diff_5516_10504# diff_2212_11356# diff_5320_10684# GND efet w=232 l=100
+ ad=15776 pd=600 as=46304 ps=1424 
M2527 GND clk2 diff_5516_10504# GND efet w=238 l=106
+ ad=0 pd=0 as=0 ps=0 
M2528 diff_5840_10504# clk1 GND GND efet w=250 l=94
+ ad=17552 pd=672 as=0 ps=0 
M2529 diff_4952_10516# diff_2104_10732# GND GND efet w=118 l=94
+ ad=0 pd=0 as=0 ps=0 
M2530 diff_5108_10516# clk2 diff_4952_10516# GND efet w=70 l=94
+ ad=7184 pd=432 as=0 ps=0 
M2531 diff_5996_10504# diff_5420_10876# diff_5840_10504# GND efet w=250 l=82
+ ad=18224 pd=624 as=0 ps=0 
M2532 diff_5884_9412# diff_6076_10456# diff_5996_10504# GND efet w=238 l=94
+ ad=126960 pd=6440 as=0 ps=0 
M2533 diff_5320_10684# diff_5116_11728# diff_5884_9412# GND efet w=244 l=82
+ ad=0 pd=0 as=0 ps=0 
M2534 diff_5884_9412# diff_4192_12940# diff_5320_10684# GND efet w=232 l=88
+ ad=0 pd=0 as=0 ps=0 
M2535 diff_4432_7336# Vdd Vdd GND efet w=52 l=352
+ ad=0 pd=0 as=0 ps=0 
M2536 GND diff_8920_12124# diff_8752_10972# GND efet w=124 l=76
+ ad=0 pd=0 as=16672 ps=624 
M2537 diff_8752_10972# Vdd Vdd GND efet w=46 l=478
+ ad=0 pd=0 as=0 ps=0 
M2538 GND diff_7696_2656# diff_9964_12124# GND efet w=88 l=88
+ ad=0 pd=0 as=142928 ps=5200 
M2539 GND diff_7696_2656# diff_9916_11896# GND efet w=94 l=94
+ ad=0 pd=0 as=63472 ps=2976 
M2540 diff_10484_11956# diff_6712_8284# GND GND efet w=100 l=88
+ ad=109440 pd=4888 as=0 ps=0 
M2541 GND diff_9448_11716# diff_9184_10600# GND efet w=622 l=82
+ ad=0 pd=0 as=149328 ps=4696 
M2542 GND clk2 diff_4672_9160# GND efet w=172 l=100
+ ad=0 pd=0 as=38992 ps=1368 
M2543 diff_6772_10208# diff_5884_9412# Vdd GND efet w=166 l=88
+ ad=145808 pd=4496 as=0 ps=0 
M2544 Vdd Vdd diff_4672_9160# GND efet w=46 l=250
+ ad=0 pd=0 as=0 ps=0 
M2545 GND diff_2068_14080# diff_2068_11368# GND efet w=178 l=106
+ ad=0 pd=0 as=0 ps=0 
M2546 Vdd diff_2788_9316# diff_2068_14080# GND efet w=328 l=88
+ ad=0 pd=0 as=0 ps=0 
M2547 diff_2068_14080# diff_2416_9340# GND GND efet w=280 l=88
+ ad=0 pd=0 as=0 ps=0 
M2548 diff_2788_9316# diff_2860_8956# diff_2788_9316# GND efet w=570 l=44
+ ad=77952 pd=2792 as=0 ps=0 
M2549 diff_2788_9316# diff_2416_9340# GND GND efet w=220 l=100
+ ad=0 pd=0 as=0 ps=0 
M2550 Vdd Vdd diff_2860_8956# GND efet w=40 l=88
+ ad=0 pd=0 as=4160 ps=288 
M2551 Vdd diff_2860_8956# diff_2788_9316# GND efet w=28 l=250
+ ad=0 pd=0 as=0 ps=0 
M2552 Vdd Vdd diff_4772_9184# GND efet w=40 l=400
+ ad=0 pd=0 as=38176 ps=1744 
M2553 diff_5872_10088# Vdd Vdd GND efet w=48 l=592
+ ad=25488 pd=1008 as=0 ps=0 
M2554 diff_4772_9184# diff_4672_9160# diff_4528_9016# GND efet w=76 l=82
+ ad=0 pd=0 as=4064 ps=336 
M2555 diff_3028_8476# diff_2804_8464# GND GND efet w=214 l=82
+ ad=43312 pd=1752 as=0 ps=0 
M2556 diff_2804_8464# clk2 diff_1840_19936# GND efet w=106 l=118
+ ad=10736 pd=464 as=805760 ps=22136 
M2557 diff_2416_9340# clk1 diff_3028_8476# GND efet w=112 l=88
+ ad=10880 pd=536 as=0 ps=0 
M2558 diff_4360_8920# Vdd Vdd GND efet w=46 l=418
+ ad=81760 pd=3360 as=0 ps=0 
M2559 Vdd Vdd diff_3028_8476# GND efet w=58 l=310
+ ad=0 pd=0 as=0 ps=0 
M2560 diff_1840_19936# clk2 diff_4828_8656# GND efet w=64 l=98
+ ad=0 pd=0 as=4160 ps=296 
M2561 diff_6772_10208# diff_5872_10088# GND GND efet w=160 l=100
+ ad=0 pd=0 as=0 ps=0 
M2562 GND diff_5884_9412# diff_5872_10088# GND efet w=88 l=88
+ ad=0 pd=0 as=0 ps=0 
M2563 Vdd diff_5908_9436# diff_5884_9412# GND efet w=46 l=430
+ ad=0 pd=0 as=0 ps=0 
M2564 diff_5908_9436# Vdd Vdd GND efet w=46 l=94
+ ad=8192 pd=528 as=0 ps=0 
M2565 diff_5884_9412# diff_5908_9436# diff_5884_9412# GND efet w=570 l=38
+ ad=0 pd=0 as=0 ps=0 
M2566 Vdd Vdd diff_4576_11152# GND efet w=80 l=450
+ ad=0 pd=0 as=237632 ps=8136 
M2567 diff_7316_9668# Vdd diff_7316_9668# GND efet w=32 l=584
+ ad=29216 pd=1176 as=0 ps=0 
M2568 diff_2104_10732# clk2 diff_6652_8776# GND efet w=58 l=100
+ ad=0 pd=0 as=8768 ps=456 
M2569 diff_6212_9136# Vdd Vdd GND efet w=40 l=460
+ ad=48160 pd=1744 as=0 ps=0 
M2570 diff_6212_9136# diff_4672_9160# diff_5944_8812# GND efet w=82 l=82
+ ad=0 pd=0 as=5504 ps=416 
M2571 GND diff_5944_8812# diff_4576_11152# GND efet w=250 l=76
+ ad=0 pd=0 as=0 ps=0 
M2572 diff_7316_9668# diff_2104_10732# GND GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M2573 GND diff_4828_8656# diff_4772_9184# GND efet w=118 l=94
+ ad=0 pd=0 as=0 ps=0 
M2574 GND diff_6652_8776# diff_6212_9136# GND efet w=118 l=82
+ ad=0 pd=0 as=0 ps=0 
M2575 GND diff_4528_9016# diff_4360_8920# GND efet w=190 l=106
+ ad=0 pd=0 as=0 ps=0 
M2576 diff_2068_11368# diff_1840_19936# GND GND efet w=172 l=100
+ ad=0 pd=0 as=0 ps=0 
M2577 Vdd diff_2792_7532# diff_1840_19936# GND efet w=312 l=176
+ ad=0 pd=0 as=0 ps=0 
M2578 GND diff_5644_7940# diff_5908_8188# GND efet w=196 l=76
+ ad=0 pd=0 as=119808 ps=4008 
M2579 diff_1840_19936# diff_2416_8008# GND GND efet w=310 l=94
+ ad=0 pd=0 as=0 ps=0 
M2580 diff_928_16456# diff_4100_7756# diff_928_16456# GND efet w=534 l=56
+ ad=447680 pd=14752 as=0 ps=0 
M2581 GND diff_4192_12940# diff_928_16456# GND efet w=574 l=94
+ ad=0 pd=0 as=0 ps=0 
M2582 diff_928_16456# diff_4100_7756# Vdd GND efet w=76 l=124
+ ad=0 pd=0 as=0 ps=0 
M2583 diff_2792_7532# diff_2860_7660# diff_2792_7532# GND efet w=632 l=68
+ ad=81888 pd=3080 as=0 ps=0 
M2584 Vdd Vdd diff_2860_7660# GND efet w=46 l=88
+ ad=0 pd=0 as=4160 ps=288 
M2585 diff_2792_7532# diff_2416_8008# GND GND efet w=232 l=100
+ ad=0 pd=0 as=0 ps=0 
M2586 diff_4100_7756# Vdd Vdd GND efet w=64 l=100
+ ad=4496 pd=288 as=0 ps=0 
M2587 diff_5908_8188# diff_6244_8068# GND GND efet w=172 l=88
+ ad=0 pd=0 as=0 ps=0 
M2588 GND diff_5912_10948# diff_9184_10600# GND efet w=604 l=88
+ ad=0 pd=0 as=0 ps=0 
M2589 GND diff_9784_10948# diff_9884_12392# GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M2590 diff_9884_12392# diff_4192_12940# GND GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M2591 diff_10796_11596# diff_8920_12124# GND GND efet w=88 l=94
+ ad=38288 pd=1576 as=0 ps=0 
M2592 diff_9964_12124# diff_4192_12940# GND GND efet w=124 l=100
+ ad=0 pd=0 as=0 ps=0 
M2593 GND diff_12196_12148# diff_9884_12392# GND efet w=100 l=84
+ ad=0 pd=0 as=0 ps=0 
M2594 diff_9884_12392# diff_12496_12980# GND GND efet w=106 l=82
+ ad=0 pd=0 as=0 ps=0 
M2595 GND diff_13372_12532# diff_9884_12392# GND efet w=88 l=76
+ ad=0 pd=0 as=0 ps=0 
M2596 diff_9884_12392# diff_13684_12616# GND GND efet w=88 l=76
+ ad=0 pd=0 as=0 ps=0 
M2597 Vdd diff_18232_11632# diff_8944_13720# GND efet w=112 l=88
+ ad=0 pd=0 as=0 ps=0 
M2598 diff_8500_13252# diff_17692_11632# GND GND efet w=558 l=98
+ ad=153296 pd=4504 as=0 ps=0 
M2599 GND diff_17792_11776# diff_10204_13336# GND efet w=270 l=122
+ ad=0 pd=0 as=43616 ps=1672 
M2600 diff_9884_12392# diff_14164_12076# GND GND efet w=94 l=82
+ ad=0 pd=0 as=0 ps=0 
M2601 GND diff_14164_15040# diff_9884_12392# GND efet w=112 l=88
+ ad=0 pd=0 as=0 ps=0 
M2602 diff_9884_12392# diff_14644_15824# GND GND efet w=118 l=82
+ ad=0 pd=0 as=0 ps=0 
M2603 GND diff_14992_15292# diff_9884_12392# GND efet w=106 l=82
+ ad=0 pd=0 as=0 ps=0 
M2604 diff_9884_12392# diff_15292_15896# GND GND efet w=106 l=82
+ ad=0 pd=0 as=0 ps=0 
M2605 diff_9964_12124# diff_14644_15824# GND GND efet w=130 l=106
+ ad=0 pd=0 as=0 ps=0 
M2606 diff_9964_12124# diff_12496_12980# GND GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M2607 GND diff_12764_14728# diff_9964_12124# GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M2608 diff_9964_12124# diff_13024_11248# GND GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M2609 GND diff_13372_12532# diff_9964_12124# GND efet w=106 l=88
+ ad=0 pd=0 as=0 ps=0 
M2610 diff_9964_12124# diff_13684_12616# GND GND efet w=118 l=82
+ ad=0 pd=0 as=0 ps=0 
M2611 GND diff_13960_12484# diff_9964_12124# GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M2612 diff_9964_12124# diff_14164_12076# GND GND efet w=106 l=94
+ ad=0 pd=0 as=0 ps=0 
M2613 GND diff_14572_12520# diff_9964_12124# GND efet w=100 l=76
+ ad=0 pd=0 as=0 ps=0 
M2614 diff_9964_12124# diff_14872_12968# GND GND efet w=106 l=76
+ ad=0 pd=0 as=0 ps=0 
M2615 GND diff_11596_12508# diff_10484_11956# GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M2616 diff_10484_11956# diff_11380_10888# GND GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M2617 diff_9184_10600# diff_9448_11188# diff_9004_4732# GND efet w=610 l=82
+ ad=0 pd=0 as=269712 ps=7872 
M2618 diff_9004_4732# diff_7012_10588# diff_9184_10600# GND efet w=622 l=82
+ ad=0 pd=0 as=0 ps=0 
M2619 GND diff_8752_10972# diff_8740_10168# GND efet w=316 l=94
+ ad=0 pd=0 as=186816 ps=6552 
M2620 GND diff_9784_10948# diff_9448_11188# GND efet w=172 l=88
+ ad=0 pd=0 as=18544 ps=960 
M2621 GND diff_9448_11716# diff_9748_9256# GND efet w=112 l=88
+ ad=0 pd=0 as=40368 ps=1448 
M2622 GND diff_10648_11020# diff_9448_11716# GND efet w=172 l=88
+ ad=0 pd=0 as=30064 ps=1344 
M2623 diff_9916_11896# diff_12496_12980# GND GND efet w=100 l=100
+ ad=0 pd=0 as=0 ps=0 
M2624 diff_10484_11956# diff_13684_12616# GND GND efet w=94 l=112
+ ad=0 pd=0 as=0 ps=0 
M2625 GND diff_13372_12532# diff_10484_11956# GND efet w=94 l=82
+ ad=0 pd=0 as=0 ps=0 
M2626 GND diff_14992_15292# diff_9964_12124# GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M2627 GND diff_14572_12520# diff_10484_11956# GND efet w=88 l=76
+ ad=0 pd=0 as=0 ps=0 
M2628 diff_10484_11956# diff_14872_12968# GND GND efet w=100 l=100
+ ad=0 pd=0 as=0 ps=0 
M2629 diff_13112_11284# diff_13180_11488# diff_13112_11284# GND efet w=524 l=120
+ ad=219440 pd=8272 as=0 ps=0 
M2630 GND diff_12764_14728# diff_10796_11596# GND efet w=88 l=88
+ ad=0 pd=0 as=0 ps=0 
M2631 diff_13112_11284# diff_13024_11248# GND GND efet w=190 l=118
+ ad=0 pd=0 as=0 ps=0 
M2632 diff_11176_10672# diff_11380_10888# GND GND efet w=118 l=82
+ ad=28096 pd=1248 as=0 ps=0 
M2633 diff_9748_9256# diff_7012_10588# GND GND efet w=124 l=94
+ ad=0 pd=0 as=0 ps=0 
M2634 GND diff_7012_10588# diff_8740_10168# GND efet w=310 l=82
+ ad=0 pd=0 as=0 ps=0 
M2635 diff_8740_10168# diff_8680_9460# diff_8740_10168# GND efet w=684 l=230
+ ad=0 pd=0 as=0 ps=0 
M2636 diff_8740_10168# diff_8680_9460# Vdd GND efet w=64 l=196
+ ad=0 pd=0 as=0 ps=0 
M2637 diff_9004_4732# diff_9220_9376# diff_9004_4732# GND efet w=606 l=410
+ ad=0 pd=0 as=0 ps=0 
M2638 diff_9448_11188# Vdd diff_9448_11188# GND efet w=26 l=380
+ ad=0 pd=0 as=0 ps=0 
M2639 GND diff_7012_10588# diff_11032_10744# GND efet w=136 l=82
+ ad=0 pd=0 as=43200 ps=1560 
M2640 diff_13112_11284# diff_13180_11488# Vdd GND efet w=40 l=328
+ ad=0 pd=0 as=0 ps=0 
M2641 diff_10796_11596# diff_13684_12616# GND GND efet w=112 l=100
+ ad=0 pd=0 as=0 ps=0 
M2642 diff_10796_11596# Vdd Vdd GND efet w=52 l=544
+ ad=0 pd=0 as=0 ps=0 
M2643 diff_10484_11956# Vdd Vdd GND efet w=52 l=568
+ ad=0 pd=0 as=0 ps=0 
M2644 GND diff_11596_12508# diff_11752_10888# GND efet w=118 l=118
+ ad=0 pd=0 as=33280 ps=1560 
M2645 GND diff_11176_10672# diff_11032_10744# GND efet w=100 l=100
+ ad=0 pd=0 as=0 ps=0 
M2646 diff_9748_9256# Vdd Vdd GND efet w=44 l=588
+ ad=0 pd=0 as=0 ps=0 
M2647 diff_9448_11716# Vdd Vdd GND efet w=64 l=352
+ ad=0 pd=0 as=0 ps=0 
M2648 GND diff_7012_10588# diff_12064_8704# GND efet w=112 l=88
+ ad=0 pd=0 as=26544 ps=1056 
M2649 diff_12064_8704# diff_11752_10888# GND GND efet w=124 l=112
+ ad=0 pd=0 as=0 ps=0 
M2650 GND diff_12196_12148# diff_12628_10672# GND efet w=88 l=88
+ ad=0 pd=0 as=10384 ps=648 
M2651 diff_9004_4732# diff_9220_9376# Vdd GND efet w=78 l=238
+ ad=0 pd=0 as=0 ps=0 
M2652 diff_8680_9460# Vdd Vdd GND efet w=40 l=88
+ ad=3680 pd=264 as=0 ps=0 
M2653 diff_9220_9376# Vdd diff_9220_9376# GND efet w=20 l=152
+ ad=3680 pd=264 as=0 ps=0 
M2654 diff_11032_10744# Vdd Vdd GND efet w=64 l=532
+ ad=0 pd=0 as=0 ps=0 
M2655 diff_11176_10672# Vdd Vdd GND efet w=40 l=496
+ ad=0 pd=0 as=0 ps=0 
M2656 Vdd Vdd diff_13180_11488# GND efet w=46 l=106
+ ad=0 pd=0 as=9440 ps=552 
M2657 Vdd Vdd diff_11752_10888# GND efet w=58 l=694
+ ad=0 pd=0 as=0 ps=0 
M2658 diff_12064_8704# Vdd Vdd GND efet w=52 l=532
+ ad=0 pd=0 as=0 ps=0 
M2659 diff_12808_6016# diff_12628_10672# GND GND efet w=106 l=88
+ ad=135792 pd=6160 as=0 ps=0 
M2660 GND diff_6772_10208# diff_12808_6016# GND efet w=100 l=100
+ ad=0 pd=0 as=0 ps=0 
M2661 diff_9964_12124# Vdd Vdd GND efet w=46 l=520
+ ad=0 pd=0 as=0 ps=0 
M2662 diff_12628_10672# Vdd diff_12628_10672# GND efet w=26 l=722
+ ad=0 pd=0 as=0 ps=0 
M2663 GND diff_7316_9668# diff_9916_2584# GND efet w=150 l=102
+ ad=0 pd=0 as=129440 ps=5712 
M2664 diff_9916_11896# diff_14872_12968# GND GND efet w=94 l=130
+ ad=0 pd=0 as=0 ps=0 
M2665 diff_10484_11956# diff_14644_15824# GND GND efet w=100 l=100
+ ad=0 pd=0 as=0 ps=0 
M2666 GND diff_14992_15292# diff_10484_11956# GND efet w=106 l=94
+ ad=0 pd=0 as=0 ps=0 
M2667 GND diff_16144_12496# diff_9884_12392# GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M2668 GND diff_14572_12520# diff_13112_11284# GND efet w=172 l=100
+ ad=0 pd=0 as=0 ps=0 
M2669 GND diff_14992_15292# diff_9916_11896# GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M2670 diff_13112_11284# diff_14644_15824# GND GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M2671 diff_9916_11896# Vdd diff_9916_11896# GND efet w=20 l=524
+ ad=0 pd=0 as=0 ps=0 
M2672 Vdd diff_17692_11632# diff_10204_13336# GND efet w=240 l=212
+ ad=0 pd=0 as=0 ps=0 
M2673 diff_8500_13252# diff_17792_11776# Vdd GND efet w=210 l=134
+ ad=0 pd=0 as=0 ps=0 
M2674 Vdd Vdd diff_17252_11776# GND efet w=62 l=342
+ ad=0 pd=0 as=37504 ps=1416 
M2675 diff_8512_13708# diff_18332_11776# Vdd GND efet w=262 l=202
+ ad=0 pd=0 as=0 ps=0 
M2676 diff_3244_29488# diff_16636_10928# diff_8500_13252# GND efet w=478 l=142
+ ad=0 pd=0 as=0 ps=0 
M2677 GND clk2 diff_13444_2608# GND efet w=442 l=94
+ ad=0 pd=0 as=171680 ps=6768 
M2678 diff_13444_2608# diff_21968_13804# diff_13444_2608# GND efet w=528 l=128
+ ad=0 pd=0 as=0 ps=0 
M2679 diff_21968_13804# Vdd Vdd GND efet w=64 l=124
+ ad=3872 pd=288 as=0 ps=0 
M2680 Vdd Vdd diff_21340_13480# GND efet w=100 l=272
+ ad=0 pd=0 as=97024 ps=2440 
M2681 diff_3040_29500# diff_16636_10928# diff_6604_14548# GND efet w=532 l=100
+ ad=0 pd=0 as=187616 ps=5288 
M2682 GND diff_18872_11924# diff_8944_12928# GND efet w=300 l=116
+ ad=0 pd=0 as=159776 ps=5304 
M2683 diff_17252_11776# diff_17140_11656# GND GND efet w=220 l=112
+ ad=0 pd=0 as=0 ps=0 
M2684 Vdd Vdd diff_17792_11776# GND efet w=62 l=306
+ ad=0 pd=0 as=35920 ps=1360 
M2685 diff_6604_14548# diff_18784_11836# GND GND efet w=574 l=94
+ ad=0 pd=0 as=0 ps=0 
M2686 diff_13444_2608# diff_21968_13804# Vdd GND efet w=100 l=124
+ ad=0 pd=0 as=0 ps=0 
M2687 diff_21340_13480# diff_13444_2608# diff_21328_11812# GND efet w=220 l=106
+ ad=0 pd=0 as=17888 ps=752 
M2688 diff_21340_13480# diff_3808_28348# GND GND efet w=436 l=100
+ ad=0 pd=0 as=0 ps=0 
M2689 Vdd diff_18784_11836# diff_8944_12928# GND efet w=426 l=206
+ ad=0 pd=0 as=0 ps=0 
M2690 diff_6604_14548# diff_18872_11924# Vdd GND efet w=228 l=122
+ ad=0 pd=0 as=0 ps=0 
M2691 Vdd Vdd diff_18332_11776# GND efet w=56 l=324
+ ad=0 pd=0 as=39808 ps=1584 
M2692 diff_17792_11776# diff_17692_11632# GND GND efet w=214 l=112
+ ad=0 pd=0 as=0 ps=0 
M2693 GND diff_17452_11152# diff_17140_11656# GND efet w=460 l=100
+ ad=0 pd=0 as=35680 ps=1504 
M2694 GND diff_17992_11260# diff_17692_11632# GND efet w=454 l=94
+ ad=0 pd=0 as=32512 ps=1536 
M2695 GND diff_15592_16384# diff_16552_11020# GND efet w=118 l=94
+ ad=0 pd=0 as=29712 ps=1512 
M2696 diff_17140_11656# Vdd Vdd GND efet w=154 l=336
+ ad=0 pd=0 as=0 ps=0 
M2697 diff_16552_11020# diff_15292_15896# GND GND efet w=112 l=82
+ ad=0 pd=0 as=0 ps=0 
M2698 diff_9884_12392# Vdd diff_9884_12392# GND efet w=26 l=614
+ ad=0 pd=0 as=0 ps=0 
M2699 GND diff_16552_11020# diff_16636_10928# GND efet w=344 l=120
+ ad=0 pd=0 as=79504 ps=2328 
M2700 Vdd Vdd diff_16552_11020# GND efet w=52 l=568
+ ad=0 pd=0 as=0 ps=0 
M2701 diff_16636_10928# diff_5912_10948# GND GND efet w=334 l=82
+ ad=0 pd=0 as=0 ps=0 
M2702 diff_18332_11776# diff_18232_11632# GND GND efet w=208 l=118
+ ad=0 pd=0 as=0 ps=0 
M2703 Vdd Vdd diff_18872_11924# GND efet w=70 l=286
+ ad=0 pd=0 as=31264 ps=1240 
M2704 diff_18872_11924# diff_18784_11836# GND GND efet w=280 l=94
+ ad=0 pd=0 as=0 ps=0 
M2705 GND diff_18532_11416# diff_18232_11632# GND efet w=466 l=94
+ ad=0 pd=0 as=30736 ps=1504 
M2706 diff_17692_11632# Vdd Vdd GND efet w=84 l=240
+ ad=0 pd=0 as=0 ps=0 
M2707 GND diff_19240_11608# diff_18784_11836# GND efet w=526 l=94
+ ad=0 pd=0 as=31648 ps=1896 
M2708 Vdd Vdd diff_22504_12736# GND efet w=64 l=88
+ ad=0 pd=0 as=4352 ps=264 
M2709 diff_21824_12772# Vdd Vdd GND efet w=64 l=136
+ ad=3776 pd=360 as=0 ps=0 
M2710 diff_21544_11692# diff_21824_12772# diff_21544_11692# GND efet w=554 l=60
+ ad=265488 pd=7008 as=0 ps=0 
M2711 diff_21544_11692# diff_21824_12772# Vdd GND efet w=76 l=112
+ ad=0 pd=0 as=0 ps=0 
M2712 Vdd diff_22504_12736# diff_22216_9928# GND efet w=76 l=88
+ ad=0 pd=0 as=238944 ps=6024 
M2713 diff_22216_9928# diff_22504_12736# diff_22216_9928# GND efet w=444 l=278
+ ad=0 pd=0 as=0 ps=0 
M2714 Vdd diff_19136_10708# diff_3040_29500# GND efet w=382 l=142
+ ad=0 pd=0 as=0 ps=0 
M2715 diff_21544_11692# diff_13096_496# GND GND efet w=2092 l=88
+ ad=0 pd=0 as=0 ps=0 
M2716 GND diff_13096_496# diff_22216_9928# GND efet w=1882 l=82
+ ad=0 pd=0 as=0 ps=0 
M2717 diff_21544_11692# diff_21328_11812# GND GND efet w=808 l=88
+ ad=0 pd=0 as=0 ps=0 
M2718 GND diff_21544_11692# diff_22216_9928# GND efet w=610 l=44
+ ad=0 pd=0 as=0 ps=0 
M2719 diff_3040_29500# diff_18892_22660# diff_19240_11608# GND efet w=76 l=100
+ ad=0 pd=0 as=4688 ps=336 
M2720 Vdd diff_19136_10708# diff_3436_29560# GND efet w=382 l=130
+ ad=0 pd=0 as=0 ps=0 
M2721 diff_18232_11632# Vdd Vdd GND efet w=107 l=391
+ ad=0 pd=0 as=0 ps=0 
M2722 diff_18784_11836# Vdd Vdd GND efet w=101 l=386
+ ad=0 pd=0 as=0 ps=0 
M2723 diff_3436_29560# diff_18892_22660# diff_18532_11416# GND efet w=82 l=106
+ ad=0 pd=0 as=3968 ps=320 
M2724 GND diff_22216_9928# d3 GND efet w=10318 l=50
+ ad=0 pd=0 as=1.38446e+06 ps=31328 
M2725 diff_3244_29488# diff_18892_22660# diff_17992_11260# GND efet w=82 l=106
+ ad=0 pd=0 as=4112 ps=320 
M2726 d3 diff_21544_11692# Vdd GND efet w=5434 l=82
+ ad=0 pd=0 as=0 ps=0 
M2727 diff_16636_10928# diff_17356_10732# diff_16636_10928# GND efet w=308 l=384
+ ad=0 pd=0 as=0 ps=0 
M2728 diff_3808_28348# diff_18892_22660# diff_17452_11152# GND efet w=76 l=88
+ ad=0 pd=0 as=4880 ps=320 
M2729 Vdd diff_17356_10732# diff_16636_10928# GND efet w=64 l=160
+ ad=0 pd=0 as=0 ps=0 
M2730 diff_3244_29488# diff_19136_10708# Vdd GND efet w=376 l=100
+ ad=0 pd=0 as=0 ps=0 
M2731 diff_3808_28348# diff_19136_10708# Vdd GND efet w=322 l=94
+ ad=0 pd=0 as=0 ps=0 
M2732 Vdd Vdd diff_17356_10732# GND efet w=52 l=88
+ ad=0 pd=0 as=3536 ps=240 
M2733 diff_18400_10900# Vdd Vdd GND efet w=58 l=292
+ ad=72368 pd=1760 as=0 ps=0 
M2734 diff_19136_10708# Vdd Vdd GND efet w=88 l=170
+ ad=77200 pd=2016 as=0 ps=0 
M2735 diff_19136_10708# diff_18400_10900# GND GND efet w=436 l=76
+ ad=0 pd=0 as=0 ps=0 
M2736 Vdd Vdd diff_17428_9724# GND efet w=84 l=308
+ ad=0 pd=0 as=47872 ps=1352 
M2737 GND diff_10796_11596# diff_16576_8896# GND efet w=88 l=94
+ ad=0 pd=0 as=24736 ps=720 
M2738 diff_18268_10112# Vdd Vdd GND efet w=52 l=160
+ ad=93792 pd=3680 as=0 ps=0 
M2739 GND diff_17896_9496# diff_19360_10352# GND efet w=466 l=118
+ ad=0 pd=0 as=26864 ps=984 
M2740 GND diff_17896_9496# diff_18268_10112# GND efet w=346 l=82
+ ad=0 pd=0 as=0 ps=0 
M2741 GND diff_13112_11284# diff_13348_8620# GND efet w=112 l=88
+ ad=0 pd=0 as=77552 ps=2784 
M2742 Vdd Vdd diff_16576_8896# GND efet w=96 l=716
+ ad=0 pd=0 as=0 ps=0 
M2743 GND diff_9916_11896# diff_13180_9256# GND efet w=88 l=82
+ ad=0 pd=0 as=66960 ps=3328 
M2744 diff_16576_8896# diff_6772_10208# GND GND efet w=94 l=112
+ ad=0 pd=0 as=0 ps=0 
M2745 diff_5524_8116# diff_12064_8704# diff_11804_9160# GND efet w=112 l=88
+ ad=419376 pd=15360 as=120512 ps=4192 
M2746 diff_10628_9424# diff_7516_12484# diff_10252_9452# GND efet w=124 l=76
+ ad=96944 pd=3864 as=23696 ps=888 
M2747 diff_10252_9452# diff_5908_8188# Vdd GND efet w=106 l=100
+ ad=0 pd=0 as=0 ps=0 
M2748 diff_13348_8620# diff_14296_9472# diff_13348_8620# GND efet w=482 l=126
+ ad=0 pd=0 as=0 ps=0 
M2749 diff_10628_9424# diff_1840_19936# diff_10456_9200# GND efet w=58 l=94
+ ad=0 pd=0 as=181584 ps=6656 
M2750 diff_13268_9304# diff_13180_9256# diff_10456_9200# GND efet w=112 l=88
+ ad=46320 pd=1840 as=0 ps=0 
M2751 diff_10456_9200# Vdd Vdd GND efet w=76 l=280
+ ad=0 pd=0 as=0 ps=0 
M2752 diff_10456_9200# diff_10676_8788# GND GND efet w=334 l=88
+ ad=0 pd=0 as=0 ps=0 
M2753 diff_11804_9160# diff_11032_10744# diff_10628_9424# GND efet w=112 l=88
+ ad=0 pd=0 as=0 ps=0 
M2754 diff_3040_29500# diff_9748_9256# diff_5524_8116# GND efet w=466 l=76
+ ad=0 pd=0 as=0 ps=0 
M2755 GND diff_6772_10208# diff_13348_8620# GND efet w=106 l=106
+ ad=0 pd=0 as=0 ps=0 
M2756 diff_13180_9256# diff_14788_9016# diff_13180_9256# GND efet w=652 l=160
+ ad=0 pd=0 as=0 ps=0 
M2757 GND diff_6772_10208# diff_13180_9256# GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M2758 GND diff_10484_11956# diff_13168_4252# GND efet w=112 l=88
+ ad=0 pd=0 as=96256 ps=4176 
M2759 diff_11984_9020# diff_11896_8968# diff_10628_9424# GND efet w=76 l=100
+ ad=94208 pd=2624 as=0 ps=0 
M2760 GND diff_10628_9424# diff_10676_8788# GND efet w=484 l=88
+ ad=0 pd=0 as=220368 ps=6776 
M2761 diff_10676_8788# Vdd Vdd GND efet w=76 l=268
+ ad=0 pd=0 as=0 ps=0 
M2762 diff_9028_7480# diff_12064_8704# diff_10628_9424# GND efet w=52 l=88
+ ad=563264 pd=17328 as=0 ps=0 
M2763 diff_13348_8620# diff_14296_9472# Vdd GND efet w=46 l=394
+ ad=0 pd=0 as=0 ps=0 
M2764 GND diff_6772_10208# diff_13168_4252# GND efet w=114 l=112
+ ad=0 pd=0 as=0 ps=0 
M2765 GND diff_9964_12124# diff_11896_8968# GND efet w=102 l=82
+ ad=0 pd=0 as=35344 ps=912 
M2766 GND diff_9884_12392# diff_11860_4588# GND efet w=118 l=92
+ ad=0 pd=0 as=24832 ps=712 
M2767 GND diff_15940_9388# diff_11896_8968# GND efet w=100 l=100
+ ad=0 pd=0 as=0 ps=0 
M2768 Vdd Vdd diff_17200_9508# GND efet w=64 l=274
+ ad=0 pd=0 as=25264 ps=808 
M2769 diff_17428_9724# clk1 GND GND efet w=178 l=94
+ ad=0 pd=0 as=0 ps=0 
M2770 diff_17632_9892# clk1 diff_18268_10112# GND efet w=166 l=148
+ ad=8624 pd=480 as=0 ps=0 
M2771 diff_19360_10352# clk1 diff_18400_10900# GND efet w=376 l=88
+ ad=0 pd=0 as=0 ps=0 
M2772 GND diff_17428_9724# diff_17200_9508# GND efet w=236 l=124
+ ad=0 pd=0 as=0 ps=0 
M2773 GND diff_17632_10108# diff_17428_9724# GND efet w=196 l=112
+ ad=0 pd=0 as=0 ps=0 
M2774 diff_18268_10112# diff_13444_2608# diff_17632_10108# GND efet w=76 l=88
+ ad=0 pd=0 as=12416 ps=752 
M2775 diff_11200_2452# diff_17200_9508# Vdd GND efet w=334 l=116
+ ad=212016 pd=4432 as=0 ps=0 
M2776 diff_17428_9724# diff_17632_9892# GND GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M2777 GND diff_17428_9724# diff_11200_2452# GND efet w=370 l=94
+ ad=0 pd=0 as=0 ps=0 
M2778 GND diff_15940_9388# diff_11860_4588# GND efet w=112 l=100
+ ad=0 pd=0 as=0 ps=0 
M2779 diff_11860_4588# Vdd Vdd GND efet w=72 l=532
+ ad=0 pd=0 as=0 ps=0 
M2780 Vdd diff_14788_9016# diff_13180_9256# GND efet w=40 l=472
+ ad=0 pd=0 as=0 ps=0 
M2781 diff_11896_8968# Vdd Vdd GND efet w=64 l=652
+ ad=0 pd=0 as=0 ps=0 
M2782 diff_14788_9016# Vdd Vdd GND efet w=52 l=88
+ ad=7696 pd=528 as=0 ps=0 
M2783 diff_14296_9472# Vdd Vdd GND efet w=58 l=76
+ ad=3824 pd=312 as=0 ps=0 
M2784 diff_18400_10900# clk2 diff_19408_9944# GND efet w=364 l=124
+ ad=0 pd=0 as=32336 ps=1080 
M2785 diff_17896_9496# clk1 diff_18568_9736# GND efet w=82 l=100
+ ad=0 pd=0 as=5696 ps=336 
M2786 GND diff_17632_9892# diff_19408_9944# GND efet w=460 l=64
+ ad=0 pd=0 as=0 ps=0 
M2787 diff_17996_9392# diff_18568_9736# GND GND efet w=484 l=70
+ ad=149744 pd=4904 as=0 ps=0 
M2788 diff_17996_9392# diff_17896_9496# diff_17816_9236# GND efet w=1032 l=104
+ ad=0 pd=0 as=71648 ps=2256 
M2789 GND diff_4192_12940# diff_17996_9392# GND efet w=490 l=88
+ ad=0 pd=0 as=0 ps=0 
M2790 diff_17816_9236# diff_13444_2608# GND GND efet w=790 l=82
+ ad=0 pd=0 as=0 ps=0 
M2791 diff_17996_9392# Vdd Vdd GND efet w=114 l=224
+ ad=0 pd=0 as=0 ps=0 
M2792 GND diff_17996_9392# diff_18800_9028# GND efet w=308 l=120
+ ad=0 pd=0 as=27088 ps=1264 
M2793 GND diff_1840_19936# diff_13268_9304# GND efet w=76 l=76
+ ad=0 pd=0 as=0 ps=0 
M2794 diff_13268_9304# diff_16576_8896# Vdd GND efet w=66 l=118
+ ad=0 pd=0 as=0 ps=0 
M2795 GND diff_9676_8548# diff_5524_8116# GND efet w=436 l=76
+ ad=0 pd=0 as=0 ps=0 
M2796 diff_5524_8116# Vdd Vdd GND efet w=46 l=232
+ ad=0 pd=0 as=0 ps=0 
M2797 diff_10676_8788# diff_9916_2584# diff_9676_8548# GND efet w=64 l=76
+ ad=0 pd=0 as=28976 ps=1280 
M2798 diff_13268_9304# diff_13348_8620# diff_10676_8788# GND efet w=124 l=100
+ ad=0 pd=0 as=0 ps=0 
M2799 GND diff_5524_8116# diff_5644_7940# GND efet w=112 l=136
+ ad=0 pd=0 as=36048 ps=1576 
M2800 Vdd Vdd diff_6112_6628# GND efet w=52 l=412
+ ad=0 pd=0 as=55712 ps=2064 
M2801 GND diff_13112_11284# diff_17564_3592# GND efet w=100 l=88
+ ad=0 pd=0 as=99024 ps=3712 
M2802 diff_17564_3592# diff_1840_19936# GND GND efet w=134 l=70
+ ad=0 pd=0 as=0 ps=0 
M2803 diff_18800_9028# Vdd Vdd GND efet w=70 l=310
+ ad=0 pd=0 as=0 ps=0 
M2804 diff_13096_496# diff_18800_9028# Vdd GND efet w=538 l=94
+ ad=283760 pd=6160 as=0 ps=0 
M2805 GND diff_1840_19936# diff_13112_11284# GND efet w=106 l=88
+ ad=0 pd=0 as=0 ps=0 
M2806 diff_15248_8240# diff_13268_9304# diff_15092_8236# GND efet w=484 l=88
+ ad=40112 pd=1472 as=27104 ps=1032 
M2807 diff_15776_8224# diff_13268_9304# diff_16088_7840# GND efet w=502 l=82
+ ad=53888 pd=2448 as=102176 ps=3096 
M2808 GND diff_14444_7820# diff_9028_7480# GND efet w=496 l=88
+ ad=0 pd=0 as=0 ps=0 
M2809 GND diff_9604_8368# diff_6112_6160# GND efet w=478 l=94
+ ad=0 pd=0 as=93696 ps=2944 
M2810 diff_10676_8200# diff_9916_2584# diff_9604_8368# GND efet w=58 l=94
+ ad=202896 pd=6104 as=23744 ps=1056 
M2811 diff_6112_6160# Vdd Vdd GND efet w=46 l=262
+ ad=0 pd=0 as=0 ps=0 
M2812 diff_13148_8404# diff_12808_6016# diff_10676_8200# GND efet w=112 l=100
+ ad=113792 pd=4376 as=0 ps=0 
M2813 diff_9028_7480# diff_14332_8212# Vdd GND efet w=100 l=76
+ ad=0 pd=0 as=0 ps=0 
M2814 diff_15092_8236# diff_13148_8404# GND GND efet w=358 l=82
+ ad=0 pd=0 as=0 ps=0 
M2815 GND diff_4096_2464# diff_928_16456# GND efet w=634 l=82
+ ad=0 pd=0 as=0 ps=0 
M2816 Vdd diff_2860_7660# diff_2792_7532# GND efet w=40 l=220
+ ad=0 pd=0 as=0 ps=0 
M2817 diff_2416_8008# clk1 diff_3028_7132# GND efet w=124 l=76
+ ad=10400 pd=512 as=46192 ps=1776 
M2818 diff_3028_7132# diff_2804_7120# GND GND efet w=220 l=100
+ ad=0 pd=0 as=0 ps=0 
M2819 diff_2804_7120# clk2 diff_1132_21544# GND efet w=112 l=88
+ ad=10544 pd=464 as=944672 ps=30200 
M2820 Vdd Vdd diff_3028_7132# GND efet w=64 l=328
+ ad=0 pd=0 as=0 ps=0 
M2821 diff_2068_11368# diff_1132_21544# GND GND efet w=184 l=94
+ ad=0 pd=0 as=0 ps=0 
M2822 GND diff_6712_8284# diff_6244_8068# GND efet w=100 l=88
+ ad=0 pd=0 as=17248 ps=624 
M2823 diff_7028_7996# diff_5644_7940# GND GND efet w=226 l=88
+ ad=15776 pd=600 as=0 ps=0 
M2824 diff_7184_7996# diff_6712_8284# diff_7028_7996# GND efet w=232 l=88
+ ad=25008 pd=920 as=0 ps=0 
M2825 GND diff_7264_8080# diff_7184_7996# GND efet w=118 l=82
+ ad=0 pd=0 as=0 ps=0 
M2826 diff_6112_6628# diff_7504_8092# GND GND efet w=136 l=88
+ ad=0 pd=0 as=0 ps=0 
M2827 diff_5644_7940# diff_5524_7192# diff_5644_7384# GND efet w=226 l=76
+ ad=0 pd=0 as=79840 ps=3040 
M2828 Vdd diff_2792_6332# diff_1132_21544# GND efet w=310 l=94
+ ad=0 pd=0 as=0 ps=0 
M2829 diff_1132_21544# diff_2416_6808# GND GND efet w=316 l=100
+ ad=0 pd=0 as=0 ps=0 
M2830 diff_2792_6332# diff_2872_6400# diff_2792_6332# GND efet w=552 l=50
+ ad=81840 pd=2864 as=0 ps=0 
M2831 diff_2792_6332# diff_2416_6808# GND GND efet w=276 l=104
+ ad=0 pd=0 as=0 ps=0 
M2832 Vdd Vdd diff_2872_6400# GND efet w=40 l=100
+ ad=0 pd=0 as=4352 ps=312 
M2833 Vdd diff_2872_6400# diff_2792_6332# GND efet w=52 l=208
+ ad=0 pd=0 as=0 ps=0 
M2834 Vdd Vdd diff_4724_6472# GND efet w=64 l=352
+ ad=0 pd=0 as=47872 ps=1544 
M2835 Vdd Vdd diff_4672_2848# GND efet w=58 l=370
+ ad=0 pd=0 as=44080 ps=1456 
M2836 diff_4360_7024# Vdd Vdd GND efet w=52 l=364
+ ad=81888 pd=2584 as=0 ps=0 
M2837 GND diff_5692_7288# diff_5644_7384# GND efet w=280 l=82
+ ad=0 pd=0 as=0 ps=0 
M2838 diff_5644_7384# diff_5848_6916# GND GND efet w=304 l=88
+ ad=0 pd=0 as=0 ps=0 
M2839 diff_5644_7940# Vdd Vdd GND efet w=40 l=412
+ ad=0 pd=0 as=0 ps=0 
M2840 diff_5908_8188# Vdd Vdd GND efet w=44 l=278
+ ad=0 pd=0 as=0 ps=0 
M2841 diff_6244_8068# Vdd Vdd GND efet w=44 l=584
+ ad=0 pd=0 as=0 ps=0 
M2842 diff_10676_8200# Vdd Vdd GND efet w=76 l=304
+ ad=0 pd=0 as=0 ps=0 
M2843 diff_6412_6028# Vdd Vdd GND efet w=50 l=386
+ ad=70224 pd=2528 as=0 ps=0 
M2844 diff_6640_4576# Vdd Vdd GND efet w=68 l=416
+ ad=92032 pd=3224 as=0 ps=0 
M2845 diff_6856_6940# Vdd Vdd GND efet w=58 l=346
+ ad=90208 pd=3080 as=0 ps=0 
M2846 Vdd Vdd diff_5944_4600# GND efet w=58 l=418
+ ad=0 pd=0 as=139600 ps=4232 
M2847 diff_7184_7996# Vdd diff_7184_7996# GND efet w=26 l=422
+ ad=0 pd=0 as=0 ps=0 
M2848 diff_7396_4528# diff_7184_7996# diff_7204_5056# GND efet w=274 l=94
+ ad=50384 pd=1608 as=190848 ps=5088 
M2849 GND diff_6112_6160# diff_7660_12052# GND efet w=172 l=88
+ ad=0 pd=0 as=129488 ps=3744 
M2850 diff_5524_8116# diff_11032_10744# diff_10780_8056# GND efet w=52 l=94
+ ad=0 pd=0 as=83552 ps=3184 
M2851 diff_10676_8200# diff_10780_8056# GND GND efet w=502 l=88
+ ad=0 pd=0 as=0 ps=0 
M2852 diff_10456_7780# Vdd Vdd GND efet w=70 l=298
+ ad=179856 pd=6080 as=0 ps=0 
M2853 diff_6112_6160# diff_9004_4732# diff_3040_29500# GND efet w=352 l=82
+ ad=0 pd=0 as=0 ps=0 
M2854 diff_7660_12052# Vdd Vdd GND efet w=64 l=364
+ ad=0 pd=0 as=0 ps=0 
M2855 GND diff_9028_7480# diff_7216_13264# GND efet w=346 l=82
+ ad=0 pd=0 as=111344 ps=3672 
M2856 GND diff_1840_19936# diff_13148_8404# GND efet w=100 l=94
+ ad=0 pd=0 as=0 ps=0 
M2857 diff_10780_8056# diff_1840_19936# diff_10456_7780# GND efet w=52 l=88
+ ad=0 pd=0 as=0 ps=0 
M2858 diff_9028_7480# diff_11860_4588# diff_10780_8056# GND efet w=76 l=88
+ ad=0 pd=0 as=0 ps=0 
M2859 GND diff_14444_7820# diff_14332_8212# GND efet w=94 l=106
+ ad=0 pd=0 as=17056 ps=672 
M2860 diff_14444_7820# diff_15316_8272# diff_15248_8240# GND efet w=496 l=94
+ ad=60736 pd=2368 as=0 ps=0 
M2861 diff_15776_8224# diff_13148_8404# GND GND efet w=508 l=88
+ ad=0 pd=0 as=0 ps=0 
M2862 diff_16088_7840# diff_15316_8272# GND GND efet w=402 l=82
+ ad=0 pd=0 as=0 ps=0 
M2863 GND diff_10676_8200# diff_10456_7780# GND efet w=292 l=88
+ ad=0 pd=0 as=0 ps=0 
M2864 diff_9028_7144# diff_12064_8704# diff_10780_8056# GND efet w=76 l=88
+ ad=513296 pd=15736 as=0 ps=0 
M2865 diff_14332_8212# Vdd Vdd GND efet w=40 l=484
+ ad=0 pd=0 as=0 ps=0 
M2866 diff_16088_7840# diff_13148_8404# diff_15932_7840# GND efet w=558 l=140
+ ad=0 pd=0 as=50656 ps=1672 
M2867 diff_15932_7840# diff_15316_8272# diff_15776_8224# GND efet w=450 l=98
+ ad=0 pd=0 as=0 ps=0 
M2868 diff_17780_8368# diff_18284_8260# GND GND efet w=174 l=98
+ ad=54224 pd=1856 as=0 ps=0 
M2869 GND diff_17996_9392# diff_13096_496# GND efet w=784 l=64
+ ad=0 pd=0 as=0 ps=0 
M2870 diff_17780_8368# diff_17564_3592# diff_15316_8272# GND efet w=106 l=82
+ ad=0 pd=0 as=75248 ps=2592 
M2871 Vdd diff_18352_7784# diff_17780_8368# GND efet w=112 l=88
+ ad=0 pd=0 as=0 ps=0 
M2872 Vdd Vdd diff_15932_7840# GND efet w=40 l=544
+ ad=0 pd=0 as=0 ps=0 
M2873 diff_14444_7820# Vdd Vdd GND efet w=52 l=436
+ ad=0 pd=0 as=0 ps=0 
M2874 diff_14876_7768# diff_14776_7576# diff_14444_7820# GND efet w=292 l=100
+ ad=60784 pd=1896 as=0 ps=0 
M2875 GND diff_13148_8404# diff_14876_7768# GND efet w=286 l=106
+ ad=0 pd=0 as=0 ps=0 
M2876 diff_14876_7768# diff_13268_9304# GND GND efet w=352 l=100
+ ad=0 pd=0 as=0 ps=0 
M2877 GND diff_15316_8272# diff_14876_7768# GND efet w=286 l=94
+ ad=0 pd=0 as=0 ps=0 
M2878 diff_3040_29500# diff_8740_10168# diff_9028_7480# GND efet w=328 l=88
+ ad=0 pd=0 as=0 ps=0 
M2879 diff_13148_8404# diff_13168_4252# diff_10456_7780# GND efet w=112 l=100
+ ad=0 pd=0 as=0 ps=0 
M2880 diff_16520_7972# diff_15932_7840# GND GND efet w=88 l=88
+ ad=13264 pd=752 as=0 ps=0 
M2881 diff_18284_8260# Vdd Vdd GND efet w=32 l=384
+ ad=13456 pd=864 as=0 ps=0 
M2882 GND diff_18352_7784# diff_18284_8260# GND efet w=118 l=94
+ ad=0 pd=0 as=0 ps=0 
M2883 Vdd Vdd diff_16520_7972# GND efet w=52 l=514
+ ad=0 pd=0 as=0 ps=0 
M2884 diff_17744_7936# diff_13112_11284# diff_15316_8272# GND efet w=118 l=94
+ ad=60896 pd=2048 as=0 ps=0 
M2885 diff_17744_7936# diff_18284_8260# Vdd GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M2886 GND diff_18352_7784# diff_17744_7936# GND efet w=184 l=82
+ ad=0 pd=0 as=0 ps=0 
M2887 Vdd diff_1840_19936# diff_18832_7564# GND efet w=52 l=88
+ ad=0 pd=0 as=23248 ps=936 
M2888 diff_14776_7576# diff_16520_7972# GND GND efet w=160 l=76
+ ad=40096 pd=1104 as=0 ps=0 
M2889 diff_3040_29500# diff_19148_7324# diff_18832_7564# GND efet w=94 l=94
+ ad=0 pd=0 as=0 ps=0 
M2890 GND diff_18832_7564# diff_18352_7784# GND efet w=340 l=110
+ ad=0 pd=0 as=72384 ps=2656 
M2891 diff_18352_7784# diff_17972_7444# diff_18352_7784# GND efet w=414 l=158
+ ad=0 pd=0 as=0 ps=0 
M2892 diff_18352_7784# diff_17972_7444# Vdd GND efet w=40 l=388
+ ad=0 pd=0 as=0 ps=0 
M2893 Vdd diff_15932_7840# diff_14776_7576# GND efet w=112 l=88
+ ad=0 pd=0 as=0 ps=0 
M2894 GND diff_14396_6788# diff_9028_7144# GND efet w=514 l=106
+ ad=0 pd=0 as=0 ps=0 
M2895 Vdd diff_13312_7312# diff_12808_6016# GND efet w=40 l=370
+ ad=0 pd=0 as=0 ps=0 
M2896 diff_12808_6016# diff_13312_7312# diff_12808_6016# GND efet w=642 l=38
+ ad=0 pd=0 as=0 ps=0 
M2897 diff_7216_13264# Vdd Vdd GND efet w=64 l=376
+ ad=0 pd=0 as=0 ps=0 
M2898 Vdd Vdd diff_7396_4528# GND efet w=64 l=352
+ ad=0 pd=0 as=0 ps=0 
M2899 GND diff_4360_7024# diff_4672_2848# GND efet w=286 l=76
+ ad=0 pd=0 as=0 ps=0 
M2900 diff_4724_6472# diff_4432_7336# GND GND efet w=178 l=100
+ ad=0 pd=0 as=0 ps=0 
M2901 GND diff_4360_7024# diff_4252_4924# GND efet w=388 l=76
+ ad=0 pd=0 as=245264 ps=6832 
M2902 diff_4672_2848# diff_4724_6472# diff_4948_6352# GND efet w=94 l=94
+ ad=0 pd=0 as=28288 ps=1240 
M2903 diff_4360_7024# diff_4192_12940# GND GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M2904 GND diff_6112_6628# diff_7204_5056# GND efet w=304 l=100
+ ad=0 pd=0 as=0 ps=0 
M2905 GND diff_4948_6352# diff_4360_7024# GND efet w=412 l=76
+ ad=0 pd=0 as=0 ps=0 
M2906 diff_5944_4600# diff_6112_6628# GND GND efet w=136 l=100
+ ad=0 pd=0 as=0 ps=0 
M2907 diff_6412_6028# diff_6112_6628# GND GND efet w=112 l=88
+ ad=0 pd=0 as=0 ps=0 
M2908 GND diff_6112_6628# diff_6640_4576# GND efet w=136 l=100
+ ad=0 pd=0 as=0 ps=0 
M2909 diff_6856_6940# diff_6112_6628# GND GND efet w=142 l=106
+ ad=0 pd=0 as=0 ps=0 
M2910 Vdd Vdd diff_5924_6196# GND efet w=40 l=484
+ ad=0 pd=0 as=48336 ps=2064 
M2911 GND diff_9028_7144# diff_7216_13264# GND efet w=322 l=82
+ ad=0 pd=0 as=0 ps=0 
M2912 diff_9028_7144# diff_8740_10168# diff_3244_29488# GND efet w=322 l=88
+ ad=0 pd=0 as=0 ps=0 
M2913 Vdd Vdd diff_13312_7312# GND efet w=40 l=88
+ ad=0 pd=0 as=2720 ps=216 
M2914 diff_9028_7144# diff_14236_7000# Vdd GND efet w=120 l=104
+ ad=0 pd=0 as=0 ps=0 
M2915 Vdd Vdd diff_16876_7300# GND efet w=66 l=94
+ ad=0 pd=0 as=6080 ps=416 
M2916 diff_3244_29488# diff_9004_4732# diff_5848_6916# GND efet w=322 l=88
+ ad=0 pd=0 as=84768 ps=2736 
M2917 diff_13112_7048# diff_12808_6016# diff_10456_6980# GND efet w=112 l=100
+ ad=122480 pd=4040 as=158448 ps=5912 
M2918 diff_15236_7196# diff_14776_7576# diff_14972_7328# GND efet w=466 l=82
+ ad=43136 pd=1424 as=35168 ps=1320 
M2919 diff_14972_7328# diff_13112_7048# GND GND efet w=472 l=88
+ ad=0 pd=0 as=0 ps=0 
M2920 diff_14236_7000# diff_15316_7072# diff_15236_7196# GND efet w=490 l=88
+ ad=64384 pd=2152 as=0 ps=0 
M2921 GND diff_5848_6916# diff_7660_12052# GND efet w=184 l=76
+ ad=0 pd=0 as=0 ps=0 
M2922 diff_10456_6980# Vdd Vdd GND efet w=82 l=286
+ ad=0 pd=0 as=0 ps=0 
M2923 diff_10456_6980# diff_1840_19936# diff_10780_6688# GND efet w=64 l=88
+ ad=0 pd=0 as=75968 ps=3360 
M2924 diff_10456_6980# diff_10676_6568# GND GND efet w=298 l=88
+ ad=0 pd=0 as=0 ps=0 
M2925 diff_9028_7480# diff_11032_10744# diff_10780_6688# GND efet w=64 l=94
+ ad=0 pd=0 as=0 ps=0 
M2926 GND diff_14236_7000# diff_14396_6788# GND efet w=94 l=82
+ ad=0 pd=0 as=18784 ps=1184 
M2927 diff_15764_7268# diff_14776_7576# diff_16088_6640# GND efet w=496 l=76
+ ad=55424 pd=2496 as=98288 ps=3064 
M2928 diff_15764_7268# diff_13112_7048# GND GND efet w=538 l=94
+ ad=0 pd=0 as=0 ps=0 
M2929 diff_16088_6640# diff_15316_7072# GND GND efet w=394 l=82
+ ad=0 pd=0 as=0 ps=0 
M2930 diff_6856_6940# diff_5924_6196# GND GND efet w=136 l=88
+ ad=0 pd=0 as=0 ps=0 
M2931 diff_5924_6196# diff_6112_6160# GND GND efet w=112 l=76
+ ad=0 pd=0 as=0 ps=0 
M2932 Vdd Vdd diff_5716_5960# GND efet w=46 l=562
+ ad=0 pd=0 as=37728 ps=1816 
M2933 diff_3028_5932# diff_2804_5924# GND GND efet w=220 l=88
+ ad=44224 pd=1728 as=0 ps=0 
M2934 diff_2804_5924# clk2 diff_2140_5752# GND efet w=106 l=94
+ ad=9968 pd=440 as=0 ps=0 
M2935 diff_2416_6808# clk1 diff_3028_5932# GND efet w=112 l=88
+ ad=10304 pd=488 as=0 ps=0 
M2936 Vdd Vdd diff_3028_5932# GND efet w=58 l=304
+ ad=0 pd=0 as=0 ps=0 
M2937 diff_5924_6196# diff_4432_7336# diff_4948_6352# GND efet w=94 l=76
+ ad=0 pd=0 as=0 ps=0 
M2938 diff_15932_6640# diff_15316_7072# diff_15764_7268# GND efet w=462 l=110
+ ad=103632 pd=4008 as=0 ps=0 
M2939 diff_16088_6640# diff_13112_7048# diff_15932_6640# GND efet w=546 l=122
+ ad=0 pd=0 as=0 ps=0 
M2940 diff_15932_6640# diff_16876_7300# diff_15932_6640# GND efet w=402 l=184
+ ad=0 pd=0 as=0 ps=0 
M2941 diff_17972_7444# Vdd Vdd GND efet w=64 l=88
+ ad=12272 pd=536 as=0 ps=0 
M2942 GND diff_6772_10208# diff_19148_7324# GND efet w=190 l=106
+ ad=0 pd=0 as=37312 ps=1120 
M2943 diff_19148_7324# Vdd Vdd GND efet w=78 l=290
+ ad=0 pd=0 as=0 ps=0 
M2944 GND diff_13112_7048# diff_14864_6556# GND efet w=280 l=112
+ ad=0 pd=0 as=67984 ps=1944 
M2945 diff_14396_6788# Vdd Vdd GND efet w=56 l=402
+ ad=0 pd=0 as=0 ps=0 
M2946 GND diff_10780_6688# diff_10676_6568# GND efet w=484 l=88
+ ad=0 pd=0 as=206976 ps=6224 
M2947 diff_9028_7144# diff_11860_4588# diff_10780_6688# GND efet w=64 l=88
+ ad=0 pd=0 as=0 ps=0 
M2948 diff_10676_6568# Vdd Vdd GND efet w=76 l=268
+ ad=0 pd=0 as=0 ps=0 
M2949 diff_8704_5404# diff_12064_8704# diff_10780_6688# GND efet w=58 l=106
+ ad=563264 pd=17080 as=0 ps=0 
M2950 diff_5848_6916# Vdd Vdd GND efet w=52 l=268
+ ad=0 pd=0 as=0 ps=0 
M2951 diff_5848_6916# diff_9616_6388# GND GND efet w=472 l=88
+ ad=0 pd=0 as=0 ps=0 
M2952 diff_10676_6568# diff_9916_2584# diff_9616_6388# GND efet w=64 l=88
+ ad=0 pd=0 as=29792 ps=1112 
M2953 Vdd diff_1840_19936# diff_13112_7048# GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M2954 diff_14236_7000# Vdd Vdd GND efet w=38 l=558
+ ad=0 pd=0 as=0 ps=0 
M2955 diff_14864_6556# diff_14776_6328# diff_14236_7000# GND efet w=286 l=94
+ ad=0 pd=0 as=0 ps=0 
M2956 diff_14864_6556# diff_14776_7576# GND GND efet w=352 l=100
+ ad=0 pd=0 as=0 ps=0 
M2957 GND diff_15316_7072# diff_14864_6556# GND efet w=292 l=76
+ ad=0 pd=0 as=0 ps=0 
M2958 diff_13112_7048# diff_13168_4252# diff_10676_6568# GND efet w=124 l=94
+ ad=0 pd=0 as=0 ps=0 
M2959 diff_5944_4600# diff_6112_6160# GND GND efet w=142 l=94
+ ad=0 pd=0 as=0 ps=0 
M2960 GND diff_4364_5608# diff_4252_4924# GND efet w=400 l=88
+ ad=0 pd=0 as=0 ps=0 
M2961 GND diff_6112_6160# diff_6412_6028# GND efet w=112 l=76
+ ad=0 pd=0 as=0 ps=0 
M2962 GND diff_6112_6160# diff_6640_4576# GND efet w=154 l=82
+ ad=0 pd=0 as=0 ps=0 
M2963 diff_2068_11368# diff_2140_5752# GND GND efet w=184 l=100
+ ad=0 pd=0 as=0 ps=0 
M2964 GND diff_4924_5944# diff_4364_5608# GND efet w=316 l=88
+ ad=0 pd=0 as=69056 ps=2616 
M2965 GND diff_6112_6160# diff_7204_5056# GND efet w=292 l=88
+ ad=0 pd=0 as=0 ps=0 
M2966 GND diff_14432_5416# diff_8704_5404# GND efet w=496 l=76
+ ad=0 pd=0 as=0 ps=0 
M2967 GND diff_9616_6172# diff_5692_7288# GND efet w=460 l=88
+ ad=0 pd=0 as=85248 ps=2760 
M2968 diff_10676_5980# diff_9916_2584# diff_9616_6172# GND efet w=52 l=100
+ ad=183696 pd=5576 as=24176 ps=1056 
M2969 diff_5692_7288# Vdd Vdd GND efet w=64 l=232
+ ad=0 pd=0 as=0 ps=0 
M2970 Vdd diff_2800_5420# diff_2140_5752# GND efet w=334 l=82
+ ad=0 pd=0 as=0 ps=0 
M2971 diff_2140_5752# diff_2428_5596# GND GND efet w=304 l=88
+ ad=0 pd=0 as=0 ps=0 
M2972 diff_4364_5608# diff_4192_12940# GND GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M2973 diff_4364_5608# Vdd Vdd GND efet w=52 l=400
+ ad=0 pd=0 as=0 ps=0 
M2974 diff_5716_5960# diff_4432_7336# diff_4924_5944# GND efet w=94 l=118
+ ad=0 pd=0 as=16048 ps=1000 
M2975 diff_6640_4576# diff_5716_5960# GND GND efet w=136 l=76
+ ad=0 pd=0 as=0 ps=0 
M2976 GND diff_5848_6916# diff_5944_4600# GND efet w=196 l=94
+ ad=0 pd=0 as=0 ps=0 
M2977 GND diff_5848_6916# diff_6412_6028# GND efet w=106 l=94
+ ad=0 pd=0 as=0 ps=0 
M2978 diff_5716_5960# diff_5848_6916# GND GND efet w=112 l=76
+ ad=0 pd=0 as=0 ps=0 
M2979 diff_12896_6136# diff_12808_6016# diff_10676_5980# GND efet w=118 l=94
+ ad=137936 pd=5072 as=0 ps=0 
M2980 diff_8704_5404# diff_14332_5812# Vdd GND efet w=106 l=118
+ ad=0 pd=0 as=0 ps=0 
M2981 diff_10676_5980# Vdd Vdd GND efet w=76 l=334
+ ad=0 pd=0 as=0 ps=0 
M2982 GND diff_5848_6916# diff_6856_6940# GND efet w=148 l=76
+ ad=0 pd=0 as=0 ps=0 
M2983 GND diff_5848_6916# diff_7204_5056# GND efet w=292 l=76
+ ad=0 pd=0 as=0 ps=0 
M2984 GND diff_4364_5608# diff_4364_5440# GND efet w=184 l=88
+ ad=0 pd=0 as=55504 ps=1960 
M2985 diff_4364_5440# Vdd Vdd GND efet w=52 l=424
+ ad=0 pd=0 as=0 ps=0 
M2986 diff_2800_5420# diff_2872_5212# diff_2800_5420# GND efet w=564 l=44
+ ad=72528 pd=2792 as=0 ps=0 
M2987 diff_2800_5420# diff_2428_5596# GND GND efet w=258 l=122
+ ad=0 pd=0 as=0 ps=0 
M2988 Vdd Vdd diff_2872_5212# GND efet w=46 l=106
+ ad=0 pd=0 as=3680 ps=336 
M2989 Vdd diff_2872_5212# diff_2800_5420# GND efet w=40 l=196
+ ad=0 pd=0 as=0 ps=0 
M2990 diff_4364_5440# diff_4724_6472# diff_4924_5944# GND efet w=76 l=88
+ ad=0 pd=0 as=0 ps=0 
M2991 Vdd Vdd diff_5888_5404# GND efet w=46 l=598
+ ad=0 pd=0 as=25680 ps=1352 
M2992 diff_5888_5404# diff_4432_7336# diff_4924_4924# GND efet w=76 l=76
+ ad=0 pd=0 as=33152 ps=1288 
M2993 diff_6412_6028# diff_5888_5404# GND GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M2994 GND diff_5692_7288# diff_7660_12052# GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M2995 diff_9028_7144# diff_11032_10744# diff_10780_5824# GND efet w=52 l=112
+ ad=0 pd=0 as=80576 ps=3240 
M2996 diff_10676_5980# diff_10780_5824# GND GND efet w=526 l=88
+ ad=0 pd=0 as=0 ps=0 
M2997 diff_10456_5560# Vdd Vdd GND efet w=94 l=298
+ ad=178896 pd=6392 as=0 ps=0 
M2998 GND diff_8704_5404# diff_7216_13264# GND efet w=346 l=82
+ ad=0 pd=0 as=0 ps=0 
M2999 diff_5888_5404# diff_5692_7288# GND GND efet w=118 l=82
+ ad=0 pd=0 as=0 ps=0 
M3000 diff_5692_7288# diff_9004_4732# diff_3436_29560# GND efet w=316 l=106
+ ad=0 pd=0 as=0 ps=0 
M3001 diff_10780_5824# diff_1840_19936# diff_10456_5560# GND efet w=58 l=94
+ ad=0 pd=0 as=0 ps=0 
M3002 diff_8704_5404# diff_11860_4588# diff_10780_5824# GND efet w=58 l=88
+ ad=0 pd=0 as=0 ps=0 
M3003 Vdd diff_16876_7300# diff_15932_6640# GND efet w=40 l=418
+ ad=0 pd=0 as=0 ps=0 
M3004 diff_17780_7108# diff_17564_3592# diff_15316_7072# GND efet w=112 l=88
+ ad=50384 pd=1760 as=68576 ps=2448 
M3005 diff_17732_6584# diff_18212_7012# GND GND efet w=160 l=88
+ ad=61616 pd=1976 as=0 ps=0 
M3006 Vdd diff_18352_6464# diff_17732_6584# GND efet w=106 l=94
+ ad=0 pd=0 as=0 ps=0 
M3007 diff_19940_7264# diff_3436_29560# GND GND efet w=466 l=94
+ ad=76096 pd=1984 as=0 ps=0 
M3008 GND diff_4192_12940# d2 GND efet w=238 l=106
+ ad=0 pd=0 as=1.18643e+06 ps=27208 
M3009 Vdd Vdd diff_19940_7264# GND efet w=82 l=328
+ ad=0 pd=0 as=0 ps=0 
M3010 diff_21440_7492# Vdd Vdd GND efet w=52 l=124
+ ad=5888 pd=456 as=0 ps=0 
M3011 Vdd Vdd diff_22204_7420# GND efet w=52 l=118
+ ad=0 pd=0 as=4064 ps=288 
M3012 diff_21268_4636# diff_21440_7492# diff_21268_4636# GND efet w=572 l=78
+ ad=283296 pd=7248 as=0 ps=0 
M3013 Vdd diff_22204_7420# diff_21856_4648# GND efet w=76 l=94
+ ad=0 pd=0 as=235152 ps=5488 
M3014 diff_21268_4636# diff_21440_7492# Vdd GND efet w=94 l=142
+ ad=0 pd=0 as=0 ps=0 
M3015 diff_20152_7084# diff_13444_2608# diff_19940_7264# GND efet w=220 l=94
+ ad=13952 pd=624 as=0 ps=0 
M3016 diff_18212_7012# Vdd Vdd GND efet w=42 l=394
+ ad=15520 pd=1008 as=0 ps=0 
M3017 diff_16508_6772# diff_15932_6640# GND GND efet w=100 l=76
+ ad=13744 pd=776 as=0 ps=0 
M3018 Vdd Vdd diff_16508_6772# GND efet w=52 l=514
+ ad=0 pd=0 as=0 ps=0 
M3019 GND diff_18352_6464# diff_18212_7012# GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M3020 diff_21856_4648# diff_22204_7420# diff_21856_4648# GND efet w=334 l=388
+ ad=0 pd=0 as=0 ps=0 
M3021 Vdd diff_1840_19936# diff_18820_6424# GND efet w=58 l=76
+ ad=0 pd=0 as=20608 ps=792 
M3022 diff_17780_7108# diff_18212_7012# Vdd GND efet w=112 l=88
+ ad=0 pd=0 as=0 ps=0 
M3023 diff_17732_6584# diff_13112_11284# diff_15316_7072# GND efet w=142 l=94
+ ad=0 pd=0 as=0 ps=0 
M3024 GND diff_18352_6464# diff_17780_7108# GND efet w=160 l=88
+ ad=0 pd=0 as=0 ps=0 
M3025 diff_21268_4636# diff_13096_496# GND GND efet w=2164 l=100
+ ad=0 pd=0 as=0 ps=0 
M3026 diff_3244_29488# diff_19148_7324# diff_18820_6424# GND efet w=94 l=106
+ ad=0 pd=0 as=0 ps=0 
M3027 diff_14776_6328# diff_16508_6772# GND GND efet w=160 l=76
+ ad=40144 pd=1104 as=0 ps=0 
M3028 GND diff_18820_6424# diff_18352_6464# GND efet w=338 l=138
+ ad=0 pd=0 as=70656 ps=2536 
M3029 Vdd diff_15932_6640# diff_14776_6328# GND efet w=112 l=76
+ ad=0 pd=0 as=0 ps=0 
M3030 diff_18352_6464# diff_17972_6124# diff_18352_6464# GND efet w=402 l=164
+ ad=0 pd=0 as=0 ps=0 
M3031 diff_18352_6464# diff_17972_6124# Vdd GND efet w=40 l=352
+ ad=0 pd=0 as=0 ps=0 
M3032 diff_15236_5852# diff_14776_6328# diff_14960_6140# GND efet w=484 l=88
+ ad=46784 pd=1472 as=37616 ps=1344 
M3033 diff_14960_6140# diff_12896_6136# GND GND efet w=496 l=76
+ ad=0 pd=0 as=0 ps=0 
M3034 diff_14432_5416# diff_15316_5860# diff_15236_5852# GND efet w=532 l=82
+ ad=68080 pd=2368 as=0 ps=0 
M3035 diff_15764_5824# diff_12896_6136# GND GND efet w=526 l=82
+ ad=62960 pd=2424 as=0 ps=0 
M3036 GND diff_10676_5980# diff_10456_5560# GND efet w=292 l=88
+ ad=0 pd=0 as=0 ps=0 
M3037 GND diff_14432_5416# diff_14332_5812# GND efet w=76 l=94
+ ad=0 pd=0 as=14704 ps=648 
M3038 GND diff_1840_19936# diff_12896_6136# GND efet w=118 l=82
+ ad=0 pd=0 as=0 ps=0 
M3039 diff_8704_4912# diff_12064_8704# diff_10780_5824# GND efet w=70 l=94
+ ad=468544 pd=14016 as=0 ps=0 
M3040 GND diff_15316_5860# diff_16088_5440# GND efet w=430 l=82
+ ad=0 pd=0 as=107936 ps=3136 
M3041 diff_15932_5440# diff_15316_5860# diff_15764_5824# GND efet w=456 l=92
+ ad=64576 pd=2000 as=0 ps=0 
M3042 diff_16088_5440# diff_12896_6136# diff_15932_5440# GND efet w=552 l=116
+ ad=0 pd=0 as=0 ps=0 
M3043 diff_15764_5824# diff_14776_6328# diff_16088_5440# GND efet w=496 l=88
+ ad=0 pd=0 as=0 ps=0 
M3044 diff_21856_4648# diff_13096_496# GND GND efet w=1882 l=76
+ ad=0 pd=0 as=0 ps=0 
M3045 GND diff_20152_7084# diff_21268_4636# GND efet w=802 l=70
+ ad=0 pd=0 as=0 ps=0 
M3046 diff_3436_29560# diff_19148_7324# diff_18832_4924# GND efet w=154 l=140
+ ad=0 pd=0 as=42880 ps=1824 
M3047 GND diff_21268_4636# diff_21856_4648# GND efet w=604 l=88
+ ad=0 pd=0 as=0 ps=0 
M3048 diff_17972_6124# Vdd Vdd GND efet w=70 l=94
+ ad=12656 pd=528 as=0 ps=0 
M3049 Vdd Vdd diff_15932_5440# GND efet w=40 l=472
+ ad=0 pd=0 as=0 ps=0 
M3050 diff_14332_5812# Vdd Vdd GND efet w=62 l=548
+ ad=0 pd=0 as=0 ps=0 
M3051 diff_3436_29560# diff_8740_10168# diff_8704_5404# GND efet w=346 l=88
+ ad=0 pd=0 as=0 ps=0 
M3052 diff_12896_6136# diff_13168_4252# diff_10456_5560# GND efet w=112 l=88
+ ad=0 pd=0 as=0 ps=0 
M3053 diff_14432_5416# Vdd Vdd GND efet w=64 l=484
+ ad=0 pd=0 as=0 ps=0 
M3054 GND diff_4204_5056# diff_4252_4924# GND efet w=352 l=76
+ ad=0 pd=0 as=0 ps=0 
M3055 diff_3028_4720# diff_2804_4724# GND GND efet w=220 l=88
+ ad=42352 pd=1728 as=0 ps=0 
M3056 diff_2428_5596# clk1 diff_3028_4720# GND efet w=106 l=94
+ ad=8960 pd=464 as=0 ps=0 
M3057 diff_2804_4724# clk2 diff_2140_4552# GND efet w=124 l=88
+ ad=9056 pd=440 as=678432 ps=18720 
M3058 GND diff_4924_4924# diff_4204_5056# GND efet w=340 l=76
+ ad=0 pd=0 as=49056 ps=1720 
M3059 GND diff_5692_7288# diff_5944_4600# GND efet w=148 l=88
+ ad=0 pd=0 as=0 ps=0 
M3060 GND diff_5692_7288# diff_6640_4576# GND efet w=160 l=88
+ ad=0 pd=0 as=0 ps=0 
M3061 GND diff_5692_7288# diff_6856_6940# GND efet w=154 l=82
+ ad=0 pd=0 as=0 ps=0 
M3062 GND diff_5692_7288# diff_7204_5056# GND efet w=292 l=76
+ ad=0 pd=0 as=0 ps=0 
M3063 diff_14864_5368# diff_14776_5116# diff_14432_5416# GND efet w=280 l=94
+ ad=67504 pd=2040 as=0 ps=0 
M3064 GND diff_12896_6136# diff_14864_5368# GND efet w=292 l=76
+ ad=0 pd=0 as=0 ps=0 
M3065 diff_14864_5368# diff_14776_6328# GND GND efet w=352 l=88
+ ad=0 pd=0 as=0 ps=0 
M3066 GND diff_15316_5860# diff_14864_5368# GND efet w=328 l=100
+ ad=0 pd=0 as=0 ps=0 
M3067 diff_13168_4252# diff_13384_4948# diff_13168_4252# GND efet w=660 l=32
+ ad=0 pd=0 as=0 ps=0 
M3068 diff_17768_5812# diff_18212_5716# GND GND efet w=178 l=88
+ ad=55808 pd=1760 as=0 ps=0 
M3069 diff_17768_5812# diff_17564_3592# diff_15316_5860# GND efet w=124 l=82
+ ad=0 pd=0 as=76976 ps=2976 
M3070 Vdd diff_18392_5236# diff_17768_5812# GND efet w=112 l=100
+ ad=0 pd=0 as=0 ps=0 
M3071 GND diff_21856_4648# d2 GND efet w=9958 l=56
+ ad=0 pd=0 as=0 ps=0 
M3072 diff_18832_4924# diff_1840_19936# Vdd GND efet w=64 l=88
+ ad=0 pd=0 as=0 ps=0 
M3073 diff_19736_5548# diff_11200_2452# GND GND efet w=208 l=100
+ ad=55344 pd=1808 as=0 ps=0 
M3074 diff_16508_5572# diff_15932_5440# GND GND efet w=100 l=82
+ ad=13024 pd=752 as=0 ps=0 
M3075 Vdd Vdd diff_16508_5572# GND efet w=40 l=520
+ ad=0 pd=0 as=0 ps=0 
M3076 diff_14776_5116# diff_16508_5572# GND GND efet w=160 l=88
+ ad=39712 pd=1128 as=0 ps=0 
M3077 diff_18212_5716# Vdd Vdd GND efet w=34 l=378
+ ad=13888 pd=960 as=0 ps=0 
M3078 GND diff_18392_5236# diff_18212_5716# GND efet w=106 l=118
+ ad=0 pd=0 as=0 ps=0 
M3079 diff_17744_5272# diff_18212_5716# Vdd GND efet w=124 l=106
+ ad=51344 pd=1832 as=0 ps=0 
M3080 GND diff_18392_5236# diff_17744_5272# GND efet w=154 l=106
+ ad=0 pd=0 as=0 ps=0 
M3081 diff_6172_4720# Vdd diff_6172_4720# GND efet w=26 l=530
+ ad=21184 pd=952 as=0 ps=0 
M3082 Vdd diff_13384_4948# diff_13168_4252# GND efet w=46 l=370
+ ad=0 pd=0 as=0 ps=0 
M3083 Vdd Vdd diff_3028_4720# GND efet w=52 l=310
+ ad=0 pd=0 as=0 ps=0 
M3084 diff_2068_11368# diff_2140_4552# GND GND efet w=178 l=88
+ ad=0 pd=0 as=0 ps=0 
M3085 diff_4204_5056# Vdd Vdd GND efet w=64 l=352
+ ad=0 pd=0 as=0 ps=0 
M3086 diff_4592_4588# Vdd Vdd GND efet w=52 l=352
+ ad=59328 pd=2248 as=0 ps=0 
M3087 Vdd diff_2800_4264# diff_2140_4552# GND efet w=316 l=100
+ ad=0 pd=0 as=0 ps=0 
M3088 diff_2140_4552# diff_2428_4396# GND GND efet w=310 l=94
+ ad=0 pd=0 as=0 ps=0 
M3089 diff_4204_5056# diff_4192_12940# GND GND efet w=208 l=82
+ ad=0 pd=0 as=0 ps=0 
M3090 GND diff_4204_5056# diff_4592_4588# GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M3091 diff_2800_4264# diff_2872_4000# diff_2800_4264# GND efet w=552 l=44
+ ad=72256 pd=2840 as=0 ps=0 
M3092 diff_2800_4264# diff_2428_4396# GND GND efet w=220 l=88
+ ad=0 pd=0 as=0 ps=0 
M3093 Vdd Vdd diff_2872_4000# GND efet w=40 l=94
+ ad=0 pd=0 as=4496 ps=312 
M3094 diff_4924_4924# diff_4724_6472# diff_4592_4588# GND efet w=70 l=106
+ ad=0 pd=0 as=0 ps=0 
M3095 GND diff_6172_4720# diff_5944_4600# GND efet w=154 l=100
+ ad=0 pd=0 as=0 ps=0 
M3096 GND diff_5524_7192# diff_6412_6028# GND efet w=118 l=82
+ ad=0 pd=0 as=0 ps=0 
M3097 diff_6172_4720# diff_5524_7192# GND GND efet w=88 l=76
+ ad=0 pd=0 as=0 ps=0 
M3098 GND diff_8704_4912# diff_7216_13264# GND efet w=334 l=82
+ ad=0 pd=0 as=0 ps=0 
M3099 GND diff_5524_7192# diff_6640_4576# GND efet w=136 l=76
+ ad=0 pd=0 as=0 ps=0 
M3100 GND diff_5524_7192# diff_6856_6940# GND efet w=154 l=118
+ ad=0 pd=0 as=0 ps=0 
M3101 GND diff_5524_7192# diff_7204_5056# GND efet w=268 l=76
+ ad=0 pd=0 as=0 ps=0 
M3102 Vdd diff_2872_4000# diff_2800_4264# GND efet w=40 l=208
+ ad=0 pd=0 as=0 ps=0 
M3103 diff_8704_4912# diff_8740_10168# diff_3808_28348# GND efet w=328 l=88
+ ad=0 pd=0 as=0 ps=0 
M3104 Vdd Vdd diff_13384_4948# GND efet w=40 l=76
+ ad=0 pd=0 as=2240 ps=192 
M3105 diff_8704_4912# diff_14224_4612# Vdd GND efet w=150 l=98
+ ad=0 pd=0 as=0 ps=0 
M3106 diff_3808_28348# diff_9004_4732# diff_5524_7192# GND efet w=328 l=88
+ ad=0 pd=0 as=73008 ps=2136 
M3107 diff_13112_4720# diff_12808_6016# diff_10456_4760# GND efet w=124 l=106
+ ad=77072 pd=2720 as=163536 ps=6056 
M3108 GND diff_7396_4528# diff_6452_4072# GND efet w=526 l=106
+ ad=0 pd=0 as=237792 ps=5960 
M3109 GND diff_5944_4600# diff_6452_4072# GND efet w=592 l=88
+ ad=0 pd=0 as=0 ps=0 
M3110 diff_6452_4072# diff_6412_6028# GND GND efet w=544 l=88
+ ad=0 pd=0 as=0 ps=0 
M3111 GND diff_6640_4576# diff_6452_4072# GND efet w=610 l=94
+ ad=0 pd=0 as=0 ps=0 
M3112 diff_6452_4072# diff_6856_6940# GND GND efet w=490 l=82
+ ad=0 pd=0 as=0 ps=0 
M3113 diff_6452_4072# Vdd Vdd GND efet w=46 l=538
+ ad=0 pd=0 as=0 ps=0 
M3114 diff_1732_2884# diff_5392_3628# diff_1732_2884# GND efet w=624 l=56
+ ad=249840 pd=8064 as=0 ps=0 
M3115 diff_1732_2884# diff_4592_4588# GND GND efet w=370 l=94
+ ad=0 pd=0 as=0 ps=0 
M3116 diff_2428_4396# clk1 diff_3028_3520# GND efet w=106 l=76
+ ad=9536 pd=488 as=39712 ps=1728 
M3117 diff_3028_3520# diff_2816_3520# GND GND efet w=232 l=94
+ ad=0 pd=0 as=0 ps=0 
M3118 Vdd Vdd diff_3028_3520# GND efet w=58 l=316
+ ad=0 pd=0 as=0 ps=0 
M3119 diff_2816_3520# clk2 diff_2068_11368# GND efet w=100 l=88
+ ad=7952 pd=392 as=0 ps=0 
M3120 GND diff_4096_2464# diff_1732_2884# GND efet w=370 l=82
+ ad=0 pd=0 as=0 ps=0 
M3121 Vdd Vdd diff_5392_3628# GND efet w=58 l=94
+ ad=0 pd=0 as=4400 ps=336 
M3122 Vdd diff_5392_3628# diff_1732_2884# GND efet w=76 l=196
+ ad=0 pd=0 as=0 ps=0 
M3123 diff_6412_3304# Vdd Vdd GND efet w=40 l=544
+ ad=209440 pd=5376 as=0 ps=0 
M3124 Vdd Vdd diff_2068_11368# GND efet w=32 l=312
+ ad=0 pd=0 as=0 ps=0 
M3125 diff_3040_2836# diff_5392_2932# diff_3040_2836# GND efet w=624 l=80
+ ad=225104 pd=7440 as=0 ps=0 
M3126 diff_3040_2836# diff_4364_5440# GND GND efet w=364 l=88
+ ad=0 pd=0 as=0 ps=0 
M3127 diff_1732_1996# diff_1732_2884# GND GND efet w=388 l=148
+ ad=34624 pd=1672 as=0 ps=0 
M3128 Vdd diff_1732_2884# cm_ram3 GND efet w=1168 l=88
+ ad=0 pd=0 as=182624 ps=4888 
M3129 diff_1732_1996# Vdd Vdd GND efet w=38 l=186
+ ad=0 pd=0 as=0 ps=0 
M3130 Vdd Vdd diff_2788_2716# GND efet w=54 l=178
+ ad=0 pd=0 as=45088 ps=1792 
M3131 GND diff_4096_2464# diff_3040_2836# GND efet w=352 l=76
+ ad=0 pd=0 as=0 ps=0 
M3132 Vdd diff_3040_2836# cm_ram2 GND efet w=1162 l=94
+ ad=0 pd=0 as=169424 ps=4960 
M3133 GND diff_5908_8188# diff_6452_4072# GND efet w=496 l=76
+ ad=0 pd=0 as=0 ps=0 
M3134 GND diff_5524_7192# diff_7660_12052# GND efet w=184 l=88
+ ad=0 pd=0 as=0 ps=0 
M3135 diff_10456_4760# Vdd Vdd GND efet w=82 l=286
+ ad=0 pd=0 as=0 ps=0 
M3136 diff_5524_7192# diff_9592_4528# GND GND efet w=436 l=100
+ ad=0 pd=0 as=0 ps=0 
M3137 diff_5524_7192# Vdd Vdd GND efet w=64 l=280
+ ad=0 pd=0 as=0 ps=0 
M3138 diff_6412_3304# diff_6412_6028# GND GND efet w=502 l=82
+ ad=0 pd=0 as=0 ps=0 
M3139 GND diff_6640_4576# diff_6412_3304# GND efet w=484 l=88
+ ad=0 pd=0 as=0 ps=0 
M3140 diff_6412_3304# diff_6856_6940# GND GND efet w=496 l=82
+ ad=0 pd=0 as=0 ps=0 
M3141 GND diff_7396_4528# diff_6412_3304# GND efet w=484 l=88
+ ad=0 pd=0 as=0 ps=0 
M3142 diff_6412_3304# diff_7696_2656# GND GND efet w=490 l=82
+ ad=0 pd=0 as=0 ps=0 
M3143 Vdd Vdd diff_5392_2932# GND efet w=58 l=94
+ ad=0 pd=0 as=4544 ps=336 
M3144 GND diff_3040_2836# diff_2788_2716# GND efet w=328 l=100
+ ad=0 pd=0 as=0 ps=0 
M3145 Vdd diff_5392_2932# diff_3040_2836# GND efet w=76 l=196
+ ad=0 pd=0 as=0 ps=0 
M3146 diff_6476_3136# Vdd Vdd GND efet w=46 l=502
+ ad=189280 pd=4840 as=0 ps=0 
M3147 GND diff_5944_4600# diff_6476_3136# GND efet w=498 l=82
+ ad=0 pd=0 as=0 ps=0 
M3148 diff_6400_2620# Vdd Vdd GND efet w=46 l=556
+ ad=266880 pd=7848 as=0 ps=0 
M3149 diff_4252_4924# diff_5644_2212# diff_4252_4924# GND efet w=642 l=50
+ ad=0 pd=0 as=0 ps=0 
M3150 cm_ram2 diff_2788_2716# GND GND efet w=2176 l=112
+ ad=0 pd=0 as=0 ps=0 
M3151 cm_ram3 diff_1732_1996# GND GND efet w=2176 l=88
+ ad=0 pd=0 as=0 ps=0 
M3152 GND diff_4096_2464# diff_3568_1552# GND efet w=352 l=100
+ ad=0 pd=0 as=151776 ps=4064 
M3153 diff_4252_4924# diff_4096_2464# GND GND efet w=484 l=88
+ ad=0 pd=0 as=0 ps=0 
M3154 diff_3568_1552# diff_4136_2152# diff_3568_1552# GND efet w=612 l=44
+ ad=0 pd=0 as=0 ps=0 
M3155 diff_4136_2152# Vdd Vdd GND efet w=58 l=94
+ ad=3872 pd=264 as=0 ps=0 
M3156 diff_3568_1552# diff_4672_2848# GND GND efet w=382 l=82
+ ad=0 pd=0 as=0 ps=0 
M3157 diff_3436_29560# diff_7516_12484# diff_6412_3304# GND efet w=400 l=88
+ ad=0 pd=0 as=0 ps=0 
M3158 diff_3808_28348# diff_7516_12484# diff_6452_4072# GND efet w=400 l=112
+ ad=0 pd=0 as=0 ps=0 
M3159 diff_6476_3136# diff_6856_6940# GND GND efet w=538 l=94
+ ad=0 pd=0 as=0 ps=0 
M3160 GND diff_7396_4528# diff_6476_3136# GND efet w=490 l=94
+ ad=0 pd=0 as=0 ps=0 
M3161 diff_6476_3136# diff_7696_2656# GND GND efet w=484 l=88
+ ad=0 pd=0 as=0 ps=0 
M3162 diff_3244_29488# diff_7516_12484# diff_6476_3136# GND efet w=412 l=88
+ ad=0 pd=0 as=0 ps=0 
M3163 diff_3040_29500# diff_7516_12484# diff_6400_2620# GND efet w=454 l=88
+ ad=0 pd=0 as=0 ps=0 
M3164 diff_10456_4760# diff_1840_19936# diff_10780_4456# GND efet w=64 l=88
+ ad=0 pd=0 as=78656 ps=3288 
M3165 diff_10456_4760# diff_10676_4348# GND GND efet w=292 l=88
+ ad=0 pd=0 as=0 ps=0 
M3166 diff_8704_5404# diff_11032_10744# diff_10780_4456# GND efet w=64 l=88
+ ad=0 pd=0 as=0 ps=0 
M3167 GND diff_14384_4388# diff_8704_4912# GND efet w=538 l=82
+ ad=0 pd=0 as=0 ps=0 
M3168 Vdd diff_15932_5440# diff_14776_5116# GND efet w=118 l=82
+ ad=0 pd=0 as=0 ps=0 
M3169 Vdd Vdd diff_16900_4696# GND efet w=40 l=88
+ ad=0 pd=0 as=2864 ps=240 
M3170 diff_17744_5272# diff_13112_11284# diff_15316_5860# GND efet w=118 l=94
+ ad=0 pd=0 as=0 ps=0 
M3171 d2 diff_21268_4636# Vdd GND efet w=5290 l=106
+ ad=0 pd=0 as=0 ps=0 
M3172 Vdd Vdd diff_19736_5548# GND efet w=84 l=428
+ ad=0 pd=0 as=0 ps=0 
M3173 diff_19736_5548# diff_19552_4808# GND GND efet w=112 l=100
+ ad=0 pd=0 as=0 ps=0 
M3174 diff_18392_5236# diff_18020_4940# Vdd GND efet w=64 l=436
+ ad=60912 pd=2200 as=0 ps=0 
M3175 diff_14960_4928# diff_13112_4720# GND GND efet w=490 l=82
+ ad=37856 pd=1296 as=0 ps=0 
M3176 GND diff_14224_4612# diff_14384_4388# GND efet w=106 l=76
+ ad=0 pd=0 as=20080 ps=1080 
M3177 diff_15236_4640# diff_14776_5116# diff_14960_4928# GND efet w=460 l=88
+ ad=47408 pd=1496 as=0 ps=0 
M3178 diff_14224_4612# diff_15304_4708# diff_15236_4640# GND efet w=532 l=76
+ ad=67072 pd=2344 as=0 ps=0 
M3179 diff_15764_4612# diff_13112_4720# GND GND efet w=622 l=150
+ ad=48848 pd=2448 as=0 ps=0 
M3180 GND diff_15304_4708# diff_16076_4240# GND efet w=502 l=226
+ ad=0 pd=0 as=103472 ps=3040 
M3181 GND diff_10780_4456# diff_10676_4348# GND efet w=478 l=106
+ ad=0 pd=0 as=229104 ps=7160 
M3182 diff_8704_4912# diff_11860_4588# diff_10780_4456# GND efet w=70 l=82
+ ad=0 pd=0 as=0 ps=0 
M3183 diff_10676_4348# Vdd Vdd GND efet w=70 l=286
+ ad=0 pd=0 as=0 ps=0 
M3184 diff_8704_4912# diff_11032_10744# diff_11804_9160# GND efet w=118 l=94
+ ad=0 pd=0 as=0 ps=0 
M3185 diff_10676_4348# diff_9916_2584# diff_9592_4528# GND efet w=52 l=100
+ ad=0 pd=0 as=23792 ps=1056 
M3186 diff_11804_9160# diff_12064_8704# diff_10780_4456# GND efet w=100 l=106
+ ad=0 pd=0 as=0 ps=0 
M3187 diff_15920_4240# diff_15304_4708# diff_15764_4612# GND efet w=450 l=98
+ ad=84720 pd=4080 as=0 ps=0 
M3188 GND diff_13112_4720# diff_14852_4156# GND efet w=286 l=94
+ ad=0 pd=0 as=67552 ps=1944 
M3189 diff_16076_4240# diff_13112_4720# diff_15920_4240# GND efet w=534 l=134
+ ad=0 pd=0 as=0 ps=0 
M3190 diff_14384_4388# Vdd Vdd GND efet w=72 l=448
+ ad=0 pd=0 as=0 ps=0 
M3191 Vdd diff_1840_19936# diff_13112_4720# GND efet w=106 l=94
+ ad=0 pd=0 as=0 ps=0 
M3192 diff_14852_4156# diff_11984_9020# diff_14224_4612# GND efet w=304 l=76
+ ad=0 pd=0 as=0 ps=0 
M3193 diff_14224_4612# Vdd Vdd GND efet w=60 l=532
+ ad=0 pd=0 as=0 ps=0 
M3194 diff_13112_4720# diff_13168_4252# diff_10676_4348# GND efet w=124 l=82
+ ad=0 pd=0 as=0 ps=0 
M3195 diff_14852_4156# diff_14776_5116# GND GND efet w=352 l=76
+ ad=0 pd=0 as=0 ps=0 
M3196 GND diff_15304_4708# diff_14852_4156# GND efet w=304 l=88
+ ad=0 pd=0 as=0 ps=0 
M3197 diff_15764_4612# diff_14776_5116# diff_16076_4240# GND efet w=472 l=76
+ ad=0 pd=0 as=0 ps=0 
M3198 GND diff_18832_4924# diff_18392_5236# GND efet w=334 l=106
+ ad=0 pd=0 as=0 ps=0 
M3199 diff_18392_5236# diff_18020_4940# diff_18392_5236# GND efet w=372 l=170
+ ad=0 pd=0 as=0 ps=0 
M3200 diff_15920_4240# diff_16900_4696# diff_15920_4240# GND efet w=466 l=274
+ ad=0 pd=0 as=0 ps=0 
M3201 diff_18020_4940# Vdd Vdd GND efet w=90 l=104
+ ad=7568 pd=568 as=0 ps=0 
M3202 diff_3436_29560# diff_19552_4808# GND GND efet w=400 l=106
+ ad=0 pd=0 as=0 ps=0 
M3203 Vdd diff_19736_5548# diff_3436_29560# GND efet w=322 l=118
+ ad=0 pd=0 as=0 ps=0 
M3204 Vdd diff_16900_4696# diff_15920_4240# GND efet w=34 l=424
+ ad=0 pd=0 as=0 ps=0 
M3205 Vdd Vdd diff_19552_4808# GND efet w=72 l=320
+ ad=0 pd=0 as=95040 ps=2888 
M3206 diff_17768_4648# diff_18200_4528# GND GND efet w=166 l=100
+ ad=58928 pd=1832 as=0 ps=0 
M3207 diff_19552_4808# d2 GND GND efet w=580 l=94
+ ad=0 pd=0 as=0 ps=0 
M3208 diff_17768_4648# diff_13112_11284# diff_15304_4708# GND efet w=112 l=88
+ ad=0 pd=0 as=52640 ps=1944 
M3209 diff_19552_4808# diff_11200_2452# GND GND efet w=364 l=94
+ ad=0 pd=0 as=0 ps=0 
M3210 Vdd diff_18560_3808# diff_17768_4648# GND efet w=106 l=94
+ ad=0 pd=0 as=0 ps=0 
M3211 diff_16532_4372# diff_15920_4240# GND GND efet w=94 l=94
+ ad=10240 pd=680 as=0 ps=0 
M3212 Vdd Vdd diff_16532_4372# GND efet w=40 l=520
+ ad=0 pd=0 as=0 ps=0 
M3213 diff_11984_9020# diff_16532_4372# GND GND efet w=148 l=88
+ ad=0 pd=0 as=0 ps=0 
M3214 diff_18200_4528# Vdd Vdd GND efet w=50 l=366
+ ad=15520 pd=984 as=0 ps=0 
M3215 GND diff_18560_3808# diff_18200_4528# GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M3216 Vdd diff_1840_19936# diff_19072_3988# GND efet w=70 l=64
+ ad=0 pd=0 as=20272 ps=768 
M3217 diff_17744_4168# diff_17564_3592# diff_15304_4708# GND efet w=118 l=94
+ ad=45200 pd=1688 as=0 ps=0 
M3218 diff_17744_4168# diff_18200_4528# Vdd GND efet w=106 l=94
+ ad=0 pd=0 as=0 ps=0 
M3219 Vdd diff_15920_4240# diff_11984_9020# GND efet w=100 l=88
+ ad=0 pd=0 as=0 ps=0 
M3220 Vdd Vdd diff_18220_4012# GND efet w=46 l=70
+ ad=0 pd=0 as=2720 ps=216 
M3221 GND diff_18560_3808# diff_17744_4168# GND efet w=160 l=88
+ ad=0 pd=0 as=0 ps=0 
M3222 diff_3808_28348# diff_19148_7324# diff_19072_3988# GND efet w=108 l=116
+ ad=0 pd=0 as=0 ps=0 
M3223 d0 GND GND GND efet w=952 l=100
+ ad=1.27115e+06 pd=28200 as=0 ps=0 
M3224 diff_9916_2584# diff_9904_2116# diff_9916_2584# GND efet w=462 l=144
+ ad=0 pd=0 as=0 ps=0 
M3225 Vdd Vdd diff_5644_2212# GND efet w=58 l=94
+ ad=0 pd=0 as=3824 ps=264 
M3226 Vdd diff_5644_2212# diff_4252_4924# GND efet w=82 l=190
+ ad=0 pd=0 as=0 ps=0 
M3227 diff_3568_1552# diff_4136_2152# Vdd GND efet w=70 l=178
+ ad=0 pd=0 as=0 ps=0 
M3228 GND diff_5944_4600# diff_6400_2620# GND efet w=508 l=110
+ ad=0 pd=0 as=0 ps=0 
M3229 GND diff_6640_4576# diff_6400_2620# GND efet w=516 l=128
+ ad=0 pd=0 as=0 ps=0 
M3230 GND diff_7396_4528# diff_6400_2620# GND efet w=490 l=94
+ ad=0 pd=0 as=0 ps=0 
M3231 GND diff_5908_8188# diff_6400_2620# GND efet w=490 l=106
+ ad=0 pd=0 as=0 ps=0 
M3232 Vdd Vdd diff_17248_3544# GND efet w=52 l=70
+ ad=0 pd=0 as=3440 ps=288 
M3233 diff_18560_3808# diff_18220_4012# diff_18560_3808# GND efet w=552 l=44
+ ad=81504 pd=2840 as=0 ps=0 
M3234 GND diff_19072_3988# diff_18560_3808# GND efet w=310 l=106
+ ad=0 pd=0 as=0 ps=0 
M3235 diff_17564_3592# diff_17248_3544# diff_17564_3592# GND efet w=540 l=44
+ ad=0 pd=0 as=0 ps=0 
M3236 diff_18560_3808# diff_18220_4012# Vdd GND efet w=40 l=328
+ ad=0 pd=0 as=0 ps=0 
M3237 diff_11344_2752# d0 GND GND efet w=586 l=94
+ ad=118544 pd=3248 as=0 ps=0 
M3238 GND diff_11344_2752# diff_3040_29500# GND efet w=400 l=88
+ ad=0 pd=0 as=0 ps=0 
M3239 GND diff_11344_2752# diff_11728_2836# GND efet w=106 l=88
+ ad=0 pd=0 as=50976 ps=1912 
M3240 d1 GND GND GND efet w=940 l=112
+ ad=1.19502e+06 pd=28320 as=0 ps=0 
M3241 diff_9916_2584# diff_9904_2116# Vdd GND efet w=52 l=424
+ ad=0 pd=0 as=0 ps=0 
M3242 Vdd Vdd diff_9904_2116# GND efet w=64 l=100
+ ad=0 pd=0 as=8432 ps=456 
M3243 diff_11344_2752# diff_11200_2452# GND GND efet w=414 l=110
+ ad=0 pd=0 as=0 ps=0 
M3244 GND diff_11200_2452# diff_11728_2836# GND efet w=202 l=88
+ ad=0 pd=0 as=0 ps=0 
M3245 diff_3040_29500# diff_11728_2836# Vdd GND efet w=310 l=100
+ ad=0 pd=0 as=0 ps=0 
M3246 diff_11344_2752# Vdd Vdd GND efet w=76 l=298
+ ad=0 pd=0 as=0 ps=0 
M3247 diff_11728_2836# Vdd Vdd GND efet w=40 l=412
+ ad=0 pd=0 as=0 ps=0 
M3248 GND diff_3040_29500# diff_13532_2848# GND efet w=466 l=94
+ ad=0 pd=0 as=58480 ps=1816 
M3249 diff_16984_2740# d1 GND GND efet w=544 l=100
+ ad=103248 pd=3056 as=0 ps=0 
M3250 diff_17564_3592# diff_17248_3544# Vdd GND efet w=46 l=268
+ ad=0 pd=0 as=0 ps=0 
M3251 GND GND d2 GND efet w=814 l=118
+ ad=0 pd=0 as=0 ps=0 
M3252 diff_13532_2848# Vdd Vdd GND efet w=100 l=316
+ ad=0 pd=0 as=0 ps=0 
M3253 GND diff_16984_2740# diff_3244_29488# GND efet w=400 l=88
+ ad=0 pd=0 as=0 ps=0 
M3254 GND diff_16984_2740# diff_17356_2836# GND efet w=130 l=82
+ ad=0 pd=0 as=47712 ps=1608 
M3255 GND diff_11200_2452# diff_17356_2836# GND efet w=210 l=98
+ ad=0 pd=0 as=0 ps=0 
M3256 diff_13532_2848# diff_13444_2608# diff_12904_1408# GND efet w=220 l=88
+ ad=0 pd=0 as=21872 ps=752 
M3257 d0 diff_10924_1780# Vdd GND efet w=5506 l=82
+ ad=0 pd=0 as=0 ps=0 
M3258 diff_3556_676# diff_3568_1552# GND GND efet w=452 l=108
+ ad=35392 pd=1688 as=0 ps=0 
M3259 Vdd diff_3568_1552# cm_ram1 GND efet w=1168 l=88
+ ad=0 pd=0 as=178496 ps=4840 
M3260 Vdd Vdd diff_3556_676# GND efet w=52 l=184
+ ad=0 pd=0 as=0 ps=0 
M3261 Vdd Vdd diff_4624_1396# GND efet w=54 l=190
+ ad=0 pd=0 as=44848 ps=1744 
M3262 GND diff_12904_1408# diff_10924_1780# GND efet w=814 l=82
+ ad=0 pd=0 as=247488 ps=7176 
M3263 Vdd diff_4252_4924# cm_ram0 GND efet w=1168 l=88
+ ad=0 pd=0 as=173600 ps=4816 
M3264 GND diff_4252_4924# diff_4624_1396# GND efet w=352 l=88
+ ad=0 pd=0 as=0 ps=0 
M3265 cm_ram1 diff_3556_676# GND GND efet w=2158 l=94
+ ad=0 pd=0 as=0 ps=0 
M3266 cm_ram0 diff_4624_1396# GND GND efet w=2116 l=88
+ ad=0 pd=0 as=0 ps=0 
M3267 GND diff_11032_748# d0 GND efet w=10090 l=50
+ ad=0 pd=0 as=0 ps=0 
M3268 diff_10924_1780# diff_13096_496# GND GND efet w=2044 l=88
+ ad=0 pd=0 as=0 ps=0 
M3269 Vdd Vdd diff_13576_1552# GND efet w=70 l=94
+ ad=0 pd=0 as=5216 ps=360 
M3270 Vdd diff_13576_1552# diff_10924_1780# GND efet w=82 l=106
+ ad=0 pd=0 as=0 ps=0 
M3271 diff_10924_1780# diff_13576_1552# diff_10924_1780# GND efet w=632 l=44
+ ad=0 pd=0 as=0 ps=0 
M3272 GND diff_10924_1780# diff_11032_748# GND efet w=670 l=94
+ ad=0 pd=0 as=227904 ps=6024 
M3273 diff_11032_748# diff_13096_496# GND GND efet w=1888 l=88
+ ad=0 pd=0 as=0 ps=0 
M3274 Vdd diff_13612_688# diff_11032_748# GND efet w=76 l=88
+ ad=0 pd=0 as=0 ps=0 
M3275 diff_11032_748# diff_13612_688# diff_11032_748# GND efet w=468 l=284
+ ad=0 pd=0 as=0 ps=0 
M3276 Vdd Vdd diff_13612_688# GND efet w=76 l=100
+ ad=0 pd=0 as=3344 ps=288 
M3277 diff_16984_2740# diff_11200_2452# GND GND efet w=358 l=106
+ ad=0 pd=0 as=0 ps=0 
M3278 Vdd Vdd diff_17356_2836# GND efet w=46 l=454
+ ad=0 pd=0 as=0 ps=0 
M3279 diff_3244_29488# diff_17356_2836# Vdd GND efet w=316 l=88
+ ad=0 pd=0 as=0 ps=0 
M3280 diff_16984_2740# Vdd Vdd GND efet w=54 l=304
+ ad=0 pd=0 as=0 ps=0 
M3281 GND diff_3244_29488# diff_19124_2776# GND efet w=412 l=82
+ ad=0 pd=0 as=62128 ps=1888 
M3282 diff_19124_2776# diff_13444_2608# diff_18520_1384# GND efet w=220 l=94
+ ad=0 pd=0 as=6896 ps=648 
M3283 diff_19124_2776# Vdd Vdd GND efet w=82 l=298
+ ad=0 pd=0 as=0 ps=0 
M3284 diff_3808_28348# diff_20044_1600# GND GND efet w=400 l=94
+ ad=0 pd=0 as=0 ps=0 
M3285 Vdd diff_20236_1148# diff_3808_28348# GND efet w=322 l=94
+ ad=0 pd=0 as=0 ps=0 
M3286 GND diff_4192_12940# d3 GND efet w=232 l=112
+ ad=0 pd=0 as=0 ps=0 
M3287 Vdd diff_16516_1768# d1 GND efet w=5632 l=88
+ ad=0 pd=0 as=0 ps=0 
M3288 d0 diff_4192_12940# GND GND efet w=268 l=88
+ ad=0 pd=0 as=0 ps=0 
M3289 GND diff_18520_1384# diff_16516_1768# GND efet w=814 l=82
+ ad=0 pd=0 as=224112 ps=6760 
M3290 diff_16516_1768# diff_13096_496# GND GND efet w=2122 l=154
+ ad=0 pd=0 as=0 ps=0 
M3291 Vdd Vdd diff_19192_1444# GND efet w=52 l=88
+ ad=0 pd=0 as=4304 ps=288 
M3292 GND diff_16648_688# d1 GND efet w=10078 l=50
+ ad=0 pd=0 as=0 ps=0 
M3293 Vdd diff_19192_1444# diff_16516_1768# GND efet w=70 l=106
+ ad=0 pd=0 as=0 ps=0 
M3294 diff_16516_1768# diff_19192_1444# diff_16516_1768# GND efet w=612 l=56
+ ad=0 pd=0 as=0 ps=0 
M3295 Vdd Vdd diff_20236_1148# GND efet w=70 l=400
+ ad=0 pd=0 as=49056 ps=1808 
M3296 Vdd Vdd diff_20044_1600# GND efet w=64 l=292
+ ad=0 pd=0 as=96352 ps=3384 
M3297 GND diff_11200_2452# diff_20044_1600# GND efet w=456 l=116
+ ad=0 pd=0 as=0 ps=0 
M3298 GND diff_16516_1768# diff_16648_688# GND efet w=616 l=100
+ ad=0 pd=0 as=209280 ps=5760 
M3299 diff_16648_688# diff_13096_496# GND GND efet w=1894 l=82
+ ad=0 pd=0 as=0 ps=0 
M3300 Vdd diff_19216_760# diff_16648_688# GND efet w=76 l=112
+ ad=0 pd=0 as=0 ps=0 
M3301 diff_16648_688# diff_19216_760# diff_16648_688# GND efet w=456 l=308
+ ad=0 pd=0 as=0 ps=0 
M3302 Vdd Vdd diff_19216_760# GND efet w=52 l=106
+ ad=0 pd=0 as=3824 ps=264 
M3303 GND diff_20044_1600# diff_20236_1148# GND efet w=180 l=128
+ ad=0 pd=0 as=0 ps=0 
M3304 diff_20236_1148# diff_11200_2452# GND GND efet w=190 l=88
+ ad=0 pd=0 as=0 ps=0 
M3305 GND d3 diff_20044_1600# GND efet w=702 l=122
+ ad=0 pd=0 as=0 ps=0 
M3306 d3 GND GND GND efet w=1024 l=100
+ ad=0 pd=0 as=0 ps=0 
M3307 d1 diff_4192_12940# GND GND efet w=244 l=82
+ ad=0 pd=0 as=0 ps=0 
C0 metal_21064_28780# gnd! 321.5fF ;**FLOATING
C1 metal_20908_28744# gnd! 706.4fF ;**FLOATING
C2 metal_21004_29344# gnd! 290.8fF ;**FLOATING
C3 metal_20788_29368# gnd! 40.4fF ;**FLOATING
C4 metal_21736_29548# gnd! 67.6fF ;**FLOATING
C5 metal_22108_29524# gnd! 248.7fF ;**FLOATING
C6 metal_21004_29560# gnd! 618.0fF ;**FLOATING
C7 metal_22108_30016# gnd! 173.8fF ;**FLOATING
C8 metal_21736_29860# gnd! 123.3fF ;**FLOATING
C9 metal_880_29200# gnd! 13.2fF ;**FLOATING
C10 metal_880_29524# gnd! 308.1fF ;**FLOATING
C11 metal_880_29692# gnd! 13.2fF ;**FLOATING
C12 metal_880_29992# gnd! 295.0fF ;**FLOATING
C13 metal_20788_31228# gnd! 1967.4fF ;**FLOATING
C14 metal_16696_31396# gnd! 2368.1fF ;**FLOATING
C15 metal_10756_31708# gnd! 543.3fF ;**FLOATING
C16 metal_9856_31348# gnd! 548.1fF ;**FLOATING
C17 metal_9268_31708# gnd! 550.7fF ;**FLOATING
C18 metal_10348_31360# gnd! 544.2fF ;**FLOATING
C19 diff_19216_760# gnd! 1192.5fF
C20 diff_16648_688# gnd! 10893.2fF
C21 diff_19192_1444# gnd! 1225.4fF
C22 diff_16516_1768# gnd! 9491.0fF
C23 diff_18520_1384# gnd! 1403.1fF
C24 diff_19124_2776# gnd! 1069.6fF
C25 diff_13612_688# gnd! 1264.1fF
C26 diff_13576_1552# gnd! 1341.0fF
C27 diff_11032_748# gnd! 10897.6fF
C28 cm_ram0 gnd! 9877.1fF
C29 cm_ram1 gnd! 10061.5fF
C30 diff_4624_1396# gnd! 2646.6fF
C31 diff_3556_676# gnd! 2488.5fF
C32 diff_10924_1780# gnd! 9536.6fF
C33 diff_12904_1408# gnd! 1679.9fF
C34 diff_17356_2836# gnd! 1382.7fF
C35 diff_13532_2848# gnd! 1008.3fF
C36 diff_20236_1148# gnd! 2938.3fF
C37 diff_20044_1600# gnd! 4333.4fF
C38 diff_16984_2740# gnd! 2460.6fF
C39 diff_11728_2836# gnd! 1699.9fF
C40 diff_11344_2752# gnd! 2688.4fF
C41 diff_17248_3544# gnd! 1380.6fF
C42 diff_9904_2116# gnd! 1530.0fF
C43 d1 gnd! 30900.9fF
C44 d0 gnd! 32124.0fF
C45 diff_18220_4012# gnd! 1272.8fF
C46 diff_19072_3988# gnd! 796.7fF
C47 diff_17744_4168# gnd! 1109.4fF
C48 diff_16532_4372# gnd! 514.8fF
C49 diff_18560_3808# gnd! 2035.7fF
C50 diff_17768_4648# gnd! 1231.6fF
C51 diff_18200_4528# gnd! 829.4fF
C52 diff_15920_4240# gnd! 2929.3fF
C53 diff_14852_4156# gnd! 1361.9fF
C54 diff_16076_4240# gnd! 2034.1fF
C55 diff_15304_4708# gnd! 3837.5fF
C56 diff_15764_4612# gnd! 1236.2fF
C57 diff_15236_4640# gnd! 818.4fF
C58 diff_14960_4928# gnd! 657.5fF
C59 diff_19552_4808# gnd! 2457.9fF
C60 diff_18020_4940# gnd! 1374.7fF
C61 diff_16900_4696# gnd! 1327.9fF
C62 diff_10676_4348# gnd! 4580.9fF
C63 diff_4136_2152# gnd! 1057.8fF
C64 diff_3568_1552# gnd! 4878.8fF
C65 diff_5644_2212# gnd! 1298.7fF
C66 diff_6400_2620# gnd! 5825.8fF
C67 diff_6476_3136# gnd! 4116.1fF
C68 cm_ram2 gnd! 11792.2fF
C69 diff_9592_4528# gnd! 1132.3fF
C70 cm_ram3 gnd! 12788.5fF
C71 diff_2788_2716# gnd! 2628.6fF
C72 diff_1732_1996# gnd! 2490.1fF
C73 diff_5392_2932# gnd! 1335.4fF
C74 diff_6412_3304# gnd! 4513.6fF
C75 diff_3040_2836# gnd! 5735.1fF
C76 diff_3028_3520# gnd! 704.5fF
C77 diff_2816_3520# gnd! 457.3fF
C78 diff_5392_3628# gnd! 1332.6fF
C79 diff_1732_2884# gnd! 6371.7fF
C80 diff_6452_4072# gnd! 5039.9fF
C81 diff_10780_4456# gnd! 2042.3fF
C82 diff_13112_4720# gnd! 4700.6fF
C83 diff_14224_4612# gnd! 2289.3fF
C84 diff_10456_4760# gnd! 2858.8fF
C85 diff_2872_4000# gnd! 1259.8fF
C86 diff_2428_4396# gnd! 1210.8fF
C87 diff_2800_4264# gnd! 1935.5fF
C88 diff_4592_4588# gnd! 1685.0fF
C89 diff_6172_4720# gnd! 1657.5fF
C90 diff_17744_5272# gnd! 1200.6fF
C91 diff_16508_5572# gnd! 553.6fF
C92 diff_19736_5548# gnd! 1688.6fF
C93 diff_18392_5236# gnd! 1757.5fF
C94 diff_17768_5812# gnd! 1193.1fF
C95 diff_18212_5716# gnd! 836.9fF
C96 diff_15932_5440# gnd! 2451.0fF
C97 diff_14384_4388# gnd! 879.4fF
C98 diff_13384_4948# gnd! 1301.9fF
C99 diff_3028_4720# gnd! 746.8fF
C100 diff_4204_5056# gnd! 1894.4fF
C101 diff_2804_4724# gnd! 481.1fF
C102 diff_14776_5116# gnd! 3455.2fF
C103 diff_14864_5368# gnd! 1371.4fF
C104 diff_18832_4924# gnd! 1621.1fF
C105 diff_16088_5440# gnd! 2095.1fF
C106 diff_8704_4912# gnd! 9732.7fF
C107 diff_15316_5860# gnd! 4163.4fF
C108 diff_15764_5824# gnd! 1498.4fF
C109 diff_15236_5852# gnd! 807.4fF
C110 diff_14960_6140# gnd! 655.6fF
C111 diff_17972_6124# gnd! 1485.6fF
C112 diff_18820_6424# gnd! 868.3fF
C113 diff_20152_7084# gnd! 1785.1fF
C114 diff_21856_4648# gnd! 11293.4fF
C115 diff_16508_6772# gnd! 524.2fF
C116 diff_21268_4636# gnd! 10428.7fF
C117 diff_22204_7420# gnd! 1250.6fF
C118 diff_21440_7492# gnd! 1360.9fF
C119 diff_19940_7264# gnd! 1296.9fF
C120 diff_18352_6464# gnd! 1854.2fF
C121 diff_17732_6584# gnd! 1620.9fF
C122 diff_17780_7108# gnd! 1214.4fF
C123 diff_10456_5560# gnd! 3118.0fF
C124 diff_4924_4924# gnd! 2090.2fF
C125 diff_5888_5404# gnd! 1782.8fF
C126 diff_2872_5212# gnd! 1216.7fF
C127 diff_4364_5440# gnd! 2301.4fF
C128 diff_10780_5824# gnd! 2091.9fF
C129 diff_12896_6136# gnd! 5450.6fF
C130 diff_2428_5596# gnd! 1201.5fF
C131 diff_2800_5420# gnd! 1959.9fF
C132 diff_10676_5980# gnd! 3749.8fF
C133 diff_14332_5812# gnd! 626.2fF
C134 diff_9616_6172# gnd! 915.0fF
C135 diff_5716_5960# gnd! 1966.4fF
C136 diff_4924_5944# gnd! 1638.4fF
C137 diff_14432_5416# gnd! 2197.0fF
C138 diff_9616_6388# gnd! 998.6fF
C139 diff_8704_5404# gnd! 11539.9fF
C140 diff_14776_6328# gnd! 3448.1fF
C141 diff_14864_6556# gnd! 1351.7fF
C142 diff_18212_7012# gnd! 820.8fF
C143 d2 gnd! 31758.2fF
C144 diff_16876_7300# gnd! 1445.8fF
C145 diff_4364_5608# gnd! 2077.0fF
C146 diff_3028_5932# gnd! 776.7fF
C147 diff_16088_6640# gnd! 1940.4fF
C148 diff_10676_6568# gnd! 4168.2fF
C149 diff_10780_6688# gnd! 2037.5fF
C150 diff_15316_7072# gnd! 4053.1fF
C151 diff_15764_7268# gnd! 1367.3fF
C152 diff_15236_7196# gnd! 747.1fF
C153 diff_14972_7328# gnd! 615.5fF
C154 diff_15932_6640# gnd! 3097.9fF
C155 diff_13112_7048# gnd! 5277.8fF
C156 diff_10456_6980# gnd! 2771.7fF
C157 diff_14236_7000# gnd! 2293.9fF
C158 diff_5924_6196# gnd! 2125.2fF
C159 diff_2804_5924# gnd! 463.1fF
C160 diff_4252_4924# gnd! 7639.6fF
C161 diff_4948_6352# gnd! 1341.2fF
C162 diff_13312_7312# gnd! 1272.5fF
C163 diff_14396_6788# gnd! 893.0fF
C164 diff_17972_7444# gnd! 1459.1fF
C165 diff_19148_7324# gnd! 3247.5fF
C166 diff_18832_7564# gnd! 932.6fF
C167 diff_17744_7936# gnd! 1329.8fF
C168 diff_16520_7972# gnd! 516.2fF
C169 diff_15932_7840# gnd! 2347.8fF
C170 diff_14776_7576# gnd! 3511.3fF
C171 diff_14876_7768# gnd! 1233.2fF
C172 diff_18352_7784# gnd! 1876.3fF
C173 diff_17780_8368# gnd! 1174.6fF
C174 diff_18284_8260# gnd! 782.0fF
C175 diff_16088_7840# gnd! 2004.6fF
C176 diff_10456_7780# gnd! 3120.9fF
C177 diff_9028_7144# gnd! 10693.2fF
C178 diff_15316_8272# gnd! 4081.2fF
C179 diff_7204_5056# gnd! 4214.9fF
C180 diff_6856_6940# gnd! 3951.6fF
C181 diff_6640_4576# gnd! 4544.6fF
C182 diff_6412_6028# gnd! 3416.7fF
C183 diff_5944_4600# gnd! 5433.2fF
C184 diff_7396_4528# gnd! 3643.9fF
C185 diff_4672_2848# gnd! 3260.9fF
C186 diff_4724_6472# gnd! 2543.6fF
C187 diff_10780_8056# gnd! 2109.8fF
C188 diff_5848_6916# gnd! 6181.9fF
C189 diff_5692_7288# gnd! 6472.1fF
C190 diff_2872_6400# gnd! 1289.3fF
C191 diff_2416_6808# gnd! 1222.7fF
C192 diff_2792_6332# gnd! 2126.6fF
C193 diff_4360_7024# gnd! 2696.8fF
C194 diff_5644_7384# gnd! 1399.0fF
C195 diff_5524_7192# gnd! 5841.3fF
C196 diff_6112_6628# gnd! 2922.1fF
C197 diff_7184_7996# gnd! 1240.0fF
C198 diff_7028_7996# gnd! 276.4fF
C199 diff_3028_7132# gnd! 810.1fF
C200 diff_2804_7120# gnd! 494.7fF
C201 diff_6112_6160# gnd! 5837.5fF
C202 diff_9604_8368# gnd! 928.3fF
C203 diff_10676_8200# gnd! 4075.4fF
C204 diff_14444_7820# gnd! 2102.4fF
C205 diff_13148_8404# gnd! 5124.9fF
C206 diff_15776_8224# gnd! 1348.4fF
C207 diff_15248_8240# gnd! 700.7fF
C208 diff_14332_8212# gnd! 622.1fF
C209 diff_15092_8236# gnd! 474.9fF
C210 diff_9676_8548# gnd! 993.5fF
C211 diff_17564_3592# gnd! 4576.3fF
C212 diff_18800_9028# gnd! 1032.9fF
C213 diff_17816_9236# gnd! 1236.6fF
C214 diff_17996_9392# gnd! 3864.7fF
C215 diff_18568_9736# gnd! 558.2fF
C216 diff_19408_9944# gnd! 560.6fF
C217 diff_11200_2452# gnd! 18257.9fF
C218 diff_17632_9892# gnd! 1733.2fF
C219 diff_17632_10108# gnd! 582.4fF
C220 diff_17200_9508# gnd! 834.9fF
C221 diff_19360_10352# gnd! 469.2fF
C222 diff_9028_7480# gnd! 11343.3fF
C223 diff_11984_9020# gnd! 5089.1fF
C224 diff_14788_9016# gnd! 1734.0fF
C225 diff_10676_8788# gnd! 4439.3fF
C226 diff_13268_9304# gnd! 4720.3fF
C227 diff_10456_9200# gnd! 3171.6fF
C228 diff_11896_8968# gnd! 3542.9fF
C229 diff_14296_9472# gnd! 1437.6fF
C230 diff_10628_9424# gnd! 2726.7fF
C231 diff_10252_9452# gnd! 414.7fF
C232 diff_11804_9160# gnd! 4100.5fF
C233 diff_13168_4252# gnd! 6164.4fF
C234 diff_13348_8620# gnd! 2583.9fF
C235 diff_13180_9256# gnd! 2549.7fF
C236 diff_11860_4588# gnd! 5661.7fF
C237 diff_16576_8896# gnd! 1319.3fF
C238 diff_18268_10112# gnd! 1647.9fF
C239 diff_17428_9724# gnd! 1931.4fF
C240 diff_18400_10900# gnd! 2381.9fF
C241 diff_17356_10732# gnd! 1369.3fF
C242 d3 gnd! 35326.3fF
C243 diff_19136_10708# gnd! 3054.4fF
C244 diff_22216_9928# gnd! 11332.9fF
C245 diff_13096_496# gnd! 23420.4fF
C246 diff_22504_12736# gnd! 1236.5fF
C247 diff_21544_11692# gnd! 9824.8fF
C248 diff_21824_12772# gnd! 1162.7fF
C249 diff_19240_11608# gnd! 643.0fF
C250 diff_16552_11020# gnd! 1230.6fF
C251 diff_18532_11416# gnd! 1607.5fF
C252 diff_17992_11260# gnd! 1882.8fF
C253 diff_21328_11812# gnd! 2643.3fF
C254 diff_21340_13480# gnd! 1650.0fF
C255 diff_17452_11152# gnd! 2262.9fF
C256 diff_18784_11836# gnd! 2423.0fF
C257 diff_18872_11924# gnd! 2712.2fF
C258 diff_21968_13804# gnd! 1233.6fF
C259 diff_13444_2608# gnd! 13675.8fF
C260 diff_12808_6016# gnd! 5716.0fF
C261 diff_9916_2584# gnd! 5740.3fF
C262 diff_12628_10672# gnd! 510.5fF
C263 diff_12064_8704# gnd! 4901.2fF
C264 diff_11752_10888# gnd! 873.6fF
C265 diff_11032_10744# gnd! 6041.1fF
C266 diff_9220_9376# gnd! 1543.4fF
C267 diff_8680_9460# gnd! 1399.5fF
C268 diff_9748_9256# gnd! 2435.0fF
C269 diff_11176_10672# gnd! 741.4fF
C270 diff_13180_11488# gnd! 1434.9fF
C271 diff_13112_11284# gnd! 11607.2fF
C272 diff_8740_10168# gnd! 7276.5fF
C273 diff_9004_4732# gnd! 8980.7fF
C274 diff_9448_11188# gnd! 938.7fF
C275 diff_10796_11596# gnd! 3932.5fF
C276 diff_17692_11632# gnd! 2258.6fF
C277 diff_9184_10600# gnd! 2577.1fF
C278 diff_2860_7660# gnd! 1294.9fF
C279 diff_4100_7756# gnd! 1112.5fF
C280 diff_2416_8008# gnd! 1228.0fF
C281 diff_2792_7532# gnd! 2421.8fF
C282 diff_5644_7940# gnd! 1596.7fF
C283 diff_5908_8188# gnd! 7443.3fF
C284 diff_6244_8068# gnd! 1012.4fF
C285 diff_6652_8776# gnd! 400.5fF
C286 diff_6212_9136# gnd! 840.3fF
C287 diff_5944_8812# gnd! 420.3fF
C288 diff_7316_9668# gnd! 2366.4fF
C289 diff_5908_9436# gnd! 1772.4fF
C290 diff_4828_8656# gnd! 465.2fF
C291 diff_3028_8476# gnd! 763.1fF
C292 diff_2804_8464# gnd! 472.6fF
C293 diff_4772_9184# gnd! 680.6fF
C294 diff_4528_9016# gnd! 841.6fF
C295 diff_5872_10088# gnd! 1160.2fF
C296 diff_2860_8956# gnd! 1250.1fF
C297 diff_2416_9340# gnd! 1224.5fF
C298 diff_2788_9316# gnd! 2034.1fF
C299 diff_4672_9160# gnd! 2401.2fF
C300 diff_6772_10208# gnd! 10787.5fF
C301 diff_9448_11716# gnd! 2161.9fF
C302 diff_10484_11956# gnd! 5555.6fF
C303 diff_9916_11896# gnd! 4356.6fF
C304 diff_8752_10972# gnd! 1733.7fF
C305 diff_9964_12124# gnd! 6820.5fF
C306 diff_5996_10504# gnd! 316.5fF
C307 diff_5840_10504# gnd! 307.7fF
C308 diff_5516_10504# gnd! 276.4fF
C309 diff_5320_10684# gnd! 1237.5fF
C310 diff_5884_9412# gnd! 2898.3fF
C311 diff_6076_10456# gnd! 1434.5fF
C312 diff_4952_10516# gnd! 525.6fF
C313 diff_3028_9676# gnd! 783.2fF
C314 diff_2792_9668# gnd! 511.7fF
C315 diff_5108_10516# gnd! 603.6fF
C316 diff_5420_10876# gnd! 1844.2fF
C317 diff_9884_12392# gnd! 7292.6fF
C318 diff_4432_7336# gnd! 9362.8fF
C319 diff_8416_12352# gnd! 630.8fF
C320 diff_5912_10948# gnd! 9523.3fF
C321 diff_8672_12820# gnd! 634.6fF
C322 diff_6512_11944# gnd! 482.0fF
C323 diff_2860_10156# gnd! 1226.6fF
C324 diff_2416_10540# gnd! 1209.7fF
C325 diff_2780_10084# gnd! 2299.2fF
C326 diff_5476_11636# gnd! 1360.1fF
C327 diff_6344_12028# gnd! 296.0fF
C328 diff_3028_10888# gnd! 787.6fF
C329 diff_2792_10864# gnd! 491.4fF
C330 diff_2860_11344# gnd! 1191.4fF
C331 diff_2068_11368# gnd! 5954.8fF
C332 diff_2404_11752# gnd! 1168.8fF
C333 diff_2780_11284# gnd! 2127.4fF
C334 diff_6508_12124# gnd! 1624.3fF
C335 diff_5216_12100# gnd! 262.4fF
C336 diff_4576_11152# gnd! 5348.5fF
C337 diff_4360_8920# gnd! 4001.2fF
C338 diff_5600_12100# gnd! 617.6fF
C339 diff_6076_12268# gnd! 984.1fF
C340 diff_8500_13252# gnd! 10131.5fF
C341 diff_10204_13336# gnd! 6399.6fF
C342 diff_8396_13108# gnd! 541.4fF
C343 diff_7516_12484# gnd! 12569.9fF
C344 diff_6712_12448# gnd! 459.1fF
C345 diff_7004_12508# gnd! 521.2fF
C346 diff_4096_2464# gnd! 10557.2fF
C347 diff_7100_12928# gnd! 417.7fF
C348 diff_4120_12124# gnd! 2888.2fF
C349 diff_2860_12400# gnd! 1238.1fF
C350 diff_5792_12544# gnd! 751.6fF
C351 diff_6472_12712# gnd! 1235.2fF
C352 diff_7420_13000# gnd! 1618.8fF
C353 diff_5524_8116# gnd! 12338.3fF
C354 diff_17792_11776# gnd! 3238.4fF
C355 diff_18232_11632# gnd! 2847.8fF
C356 diff_8408_13540# gnd! 654.5fF
C357 diff_8944_13720# gnd! 7731.6fF
C358 diff_7660_12052# gnd! 7972.3fF
C359 diff_17140_11656# gnd! 2861.7fF
C360 diff_17252_11776# gnd! 3292.1fF
C361 diff_18332_11776# gnd! 3519.3fF
C362 diff_16900_14392# gnd! 413.5fF
C363 diff_8512_13708# gnd! 9917.7fF
C364 diff_7720_13960# gnd! 2223.0fF
C365 diff_7744_14056# gnd! 1350.4fF
C366 diff_8212_14116# gnd! 7768.3fF
C367 diff_7216_13264# gnd! 8349.3fF
C368 diff_7588_13816# gnd! 1202.3fF
C369 diff_7060_14084# gnd! 2469.1fF
C370 diff_5116_11728# gnd! 4543.4fF
C371 diff_4636_12124# gnd! 667.4fF
C372 diff_2780_12500# gnd! 2070.4fF
C373 diff_4300_13492# gnd! 3926.1fF
C374 diff_6604_14020# gnd! 1043.0fF
C375 diff_5240_13720# gnd! 460.3fF
C376 diff_5308_13696# gnd! 521.2fF
C377 diff_2428_12196# gnd! 1169.4fF
C378 diff_2752_13076# gnd! 1216.0fF
C379 diff_2608_13384# gnd! 781.5fF
C380 diff_3076_13504# gnd! 1175.5fF
C381 diff_2996_13528# gnd! 1962.7fF
C382 diff_5644_14008# gnd! 1027.3fF
C383 diff_6076_14080# gnd! 1661.1fF
C384 diff_18364_14864# gnd! 244.7fF
C385 diff_18032_14824# gnd! 606.3fF
C386 diff_17852_14980# gnd! 695.4fF
C387 diff_15940_9388# gnd! 4190.1fF
C388 diff_7012_10588# gnd! 9987.4fF
C389 diff_14872_12968# gnd! 2973.9fF
C390 diff_14572_12520# gnd! 3147.1fF
C391 diff_14164_12076# gnd! 2659.7fF
C392 diff_13960_12484# gnd! 2439.2fF
C393 diff_8212_13960# gnd! 10610.1fF
C394 diff_16636_10928# gnd! 6974.5fF
C395 diff_19000_15988# gnd! 815.7fF
C396 diff_17824_16204# gnd! 2926.5fF
C397 diff_13684_12616# gnd! 2918.2fF
C398 diff_13372_12532# gnd! 2680.6fF
C399 diff_13024_11248# gnd! 3291.7fF
C400 diff_12196_12148# gnd! 3644.3fF
C401 diff_11380_10888# gnd! 3817.9fF
C402 diff_11596_12508# gnd! 3687.1fF
C403 diff_10648_11020# gnd! 3088.6fF
C404 diff_12496_12980# gnd! 2974.7fF
C405 diff_12764_14728# gnd! 2855.5fF
C406 diff_6712_8284# gnd! 7880.8fF
C407 diff_7696_2656# gnd! 9691.8fF
C408 diff_7504_8092# gnd! 7108.0fF
C409 diff_7264_8080# gnd! 6043.6fF
C410 diff_8896_12352# gnd! 2385.6fF
C411 diff_6136_14144# gnd! 338.2fF
C412 diff_5584_14080# gnd! 519.7fF
C413 diff_6844_13916# gnd! 777.7fF
C414 diff_5512_12820# gnd! 8671.2fF
C415 diff_7744_12340# gnd! 6276.4fF
C416 diff_5536_14200# gnd! 300.6fF
C417 diff_6136_14300# gnd! 352.6fF
C418 diff_5020_13900# gnd! 1016.9fF
C419 diff_4120_13972# gnd! 2279.5fF
C420 diff_5704_12496# gnd! 2549.7fF
C421 diff_7472_14668# gnd! 336.3fF
C422 diff_8480_14848# gnd! 777.9fF
C423 diff_8044_14476# gnd! 538.6fF
C424 diff_4360_13720# gnd! 701.7fF
C425 diff_7576_16108# gnd! 6875.2fF
C426 diff_6604_14548# gnd! 14178.7fF
C427 diff_4976_15892# gnd! 206.3fF
C428 diff_4376_15940# gnd! 810.0fF
C429 diff_16852_15544# gnd! 4269.4fF
C430 diff_17824_15484# gnd! 3827.2fF
C431 diff_20848_16804# gnd! 963.9fF
C432 diff_16852_16108# gnd! 3095.1fF
C433 diff_20260_16504# gnd! 1596.3fF
C434 diff_19720_16504# gnd! 2002.9fF
C435 diff_19180_16528# gnd! 2271.3fF
C436 diff_20980_18032# gnd! 1548.8fF
C437 diff_18220_17272# gnd! 2705.9fF
C438 diff_18280_16804# gnd! 3132.7fF
C439 diff_6976_16348# gnd! 7510.8fF
C440 diff_5132_15892# gnd! 1773.3fF
C441 diff_7276_16504# gnd! 7602.2fF
C442 diff_17320_17404# gnd! 2482.8fF
C443 diff_17332_16324# gnd! 4874.8fF
C444 diff_6676_16672# gnd! 8954.0fF
C445 diff_6676_16900# gnd! 8897.1fF
C446 diff_15592_16384# gnd! 4840.0fF
C447 diff_5272_16192# gnd! 439.3fF
C448 diff_5204_16384# gnd! 688.0fF
C449 diff_5600_16228# gnd! 1586.6fF
C450 diff_5816_16240# gnd! 1737.5fF
C451 diff_9520_16492# gnd! 2953.4fF
C452 diff_20740_18548# gnd! 832.6fF
C453 diff_20348_18460# gnd! 220.4fF
C454 diff_20740_18704# gnd! 329.8fF
C455 diff_20740_18860# gnd! 377.6fF
C456 diff_17896_9496# gnd! 9616.8fF
C457 diff_19532_18580# gnd! 308.0fF
C458 diff_19688_18628# gnd! 1117.1fF
C459 diff_6904_14332# gnd! 3347.6fF
C460 diff_6976_17140# gnd! 8579.7fF
C461 diff_6556_14212# gnd! 3442.8fF
C462 diff_5812_16768# gnd! 2661.7fF
C463 diff_13252_16600# gnd! 3825.3fF
C464 diff_7384_14632# gnd! 2640.2fF
C465 diff_4720_16588# gnd! 1645.6fF
C466 diff_6676_17296# gnd! 8895.5fF
C467 diff_15292_15896# gnd! 5626.2fF
C468 diff_14992_15292# gnd! 4740.8fF
C469 diff_14644_15824# gnd! 5015.3fF
C470 diff_14164_15040# gnd! 4965.6fF
C471 diff_16144_12496# gnd! 7795.5fF
C472 diff_20656_19484# gnd! 290.4fF
C473 diff_18976_18112# gnd! 1444.5fF
C474 diff_20116_18580# gnd! 1163.2fF
C475 diff_20572_19660# gnd! 352.4fF
C476 diff_20572_19796# gnd! 893.7fF
C477 diff_19336_18748# gnd! 1225.4fF
C478 diff_16376_18520# gnd! 242.6fF
C479 diff_18040_19408# gnd! 473.0fF
C480 diff_18356_18196# gnd! 2726.3fF
C481 diff_17980_18148# gnd! 2904.0fF
C482 diff_18008_19060# gnd! 1984.8fF
C483 diff_17600_19420# gnd! 743.6fF
C484 diff_17084_19288# gnd! 242.6fF
C485 diff_16936_19336# gnd! 512.1fF
C486 diff_15992_18424# gnd! 339.0fF
C487 diff_9784_10948# gnd! 5880.6fF
C488 diff_11848_16852# gnd! 3238.8fF
C489 diff_13672_16400# gnd! 4201.4fF
C490 diff_16532_18520# gnd! 787.1fF
C491 diff_16376_19108# gnd! 242.6fF
C492 diff_15992_19108# gnd! 252.2fF
C493 diff_14176_18496# gnd! 2071.1fF
C494 diff_8920_12124# gnd! 6172.9fF
C495 diff_14516_18124# gnd! 769.9fF
C496 diff_14872_18520# gnd! 1188.1fF
C497 diff_14344_18676# gnd! 818.0fF
C498 diff_15316_19108# gnd! 837.4fF
C499 diff_15836_18652# gnd! 741.8fF
C500 diff_17452_19432# gnd! 600.6fF
C501 diff_14992_18404# gnd! 2288.7fF
C502 diff_15316_19232# gnd! 290.4fF
C503 diff_14344_18812# gnd! 701.8fF
C504 diff_7864_17452# gnd! 8255.3fF
C505 diff_8212_16444# gnd! 3401.4fF
C506 diff_7912_17540# gnd! 3233.1fF
C507 diff_11548_16012# gnd! 4209.1fF
C508 diff_13564_19468# gnd! 470.7fF
C509 diff_13004_19000# gnd! 477.7fF
C510 diff_8944_12928# gnd! 17746.9fF
C511 diff_13564_19592# gnd! 1480.8fF
C512 diff_12856_19024# gnd! 881.9fF
C513 diff_19900_20720# gnd! 699.2fF
C514 diff_19156_20272# gnd! 1530.8fF
C515 diff_18148_20656# gnd! 1513.9fF
C516 diff_18220_20996# gnd! 1280.6fF
C517 diff_18040_19532# gnd! 2422.6fF
C518 diff_19228_20764# gnd! 4196.7fF
C519 diff_15664_19120# gnd! 2071.9fF
C520 diff_12344_19228# gnd! 242.6fF
C521 diff_10664_18676# gnd! 1292.8fF
C522 diff_10564_18232# gnd! 3032.6fF
C523 diff_11828_19228# gnd! 202.5fF
C524 diff_12164_19364# gnd! 290.6fF
C525 diff_11884_18124# gnd! 7519.3fF
C526 diff_12100_17968# gnd! 7535.4fF
C527 diff_12028_18580# gnd! 4200.2fF
C528 diff_13744_19760# gnd! 1055.7fF
C529 diff_14128_19912# gnd! 1020.6fF
C530 diff_17080_20656# gnd! 1430.8fF
C531 diff_16300_20812# gnd! 2567.4fF
C532 diff_16732_20032# gnd! 1648.6fF
C533 diff_17452_19928# gnd! 1742.2fF
C534 diff_20092_21392# gnd! 314.9fF
C535 diff_19928_21736# gnd! 761.9fF
C536 diff_19648_21692# gnd! 441.7fF
C537 diff_18880_21544# gnd! 2305.0fF
C538 diff_18292_21404# gnd! 348.0fF
C539 diff_18220_21328# gnd! 624.6fF
C540 diff_18316_21548# gnd! 2431.6fF
C541 diff_18824_21640# gnd! 1122.8fF
C542 diff_17668_21404# gnd! 311.2fF
C543 diff_11984_19228# gnd! 1103.9fF
C544 diff_11524_19384# gnd! 836.7fF
C545 diff_11060_19228# gnd! 290.6fF
C546 diff_10904_19228# gnd! 290.4fF
C547 diff_10792_18352# gnd! 3502.3fF
C548 diff_8476_18188# gnd! 276.4fF
C549 diff_9064_18608# gnd! 206.3fF
C550 diff_10508_20008# gnd! 282.0fF
C551 diff_8476_18344# gnd! 1714.7fF
C552 diff_8308_18688# gnd! 958.4fF
C553 diff_8476_18004# gnd! 3350.9fF
C554 diff_7172_18664# gnd! 206.3fF
C555 diff_7160_18400# gnd! 920.1fF
C556 diff_10664_19996# gnd! 370.5fF
C557 diff_10972_20356# gnd! 2596.2fF
C558 diff_15856_21436# gnd! 311.7fF
C559 diff_15232_21416# gnd! 311.0fF
C560 diff_17516_21736# gnd! 741.2fF
C561 diff_17212_21704# gnd! 440.8fF
C562 diff_8908_18832# gnd! 9046.4fF
C563 diff_12416_19756# gnd! 1086.6fF
C564 diff_11600_20908# gnd! 280.7fF
C565 diff_11512_20872# gnd! 576.9fF
C566 diff_10264_20224# gnd! 1138.1fF
C567 diff_11216_20812# gnd! 280.1fF
C568 diff_11060_20488# gnd! 2678.3fF
C569 diff_15796_21328# gnd! 676.1fF
C570 diff_15116_21748# gnd! 701.7fF
C571 diff_16456_21556# gnd! 3743.6fF
C572 diff_15892_21560# gnd! 4630.3fF
C573 diff_14824_21716# gnd! 422.0fF
C574 diff_13468_21416# gnd! 304.3fF
C575 diff_13336_21568# gnd! 2835.6fF
C576 diff_13408_21340# gnd! 655.5fF
C577 diff_13492_21712# gnd! 4594.6fF
C578 diff_11068_21100# gnd! 489.9fF
C579 diff_11708_21568# gnd! 566.3fF
C580 diff_9080_19840# gnd! 1511.4fF
C581 diff_7228_18940# gnd! 3419.6fF
C582 diff_4408_17236# gnd! 1492.9fF
C583 diff_4936_17224# gnd! 1171.0fF
C584 diff_5624_18136# gnd! 318.5fF
C585 diff_5092_17944# gnd! 2086.2fF
C586 diff_5240_18248# gnd! 376.1fF
C587 diff_4712_18160# gnd! 329.2fF
C588 diff_4556_18160# gnd! 338.2fF
C589 diff_4456_14788# gnd! 6025.7fF
C590 diff_7324_19300# gnd! 826.2fF
C591 diff_7408_20204# gnd! 428.1fF
C592 diff_6496_19828# gnd! 1357.6fF
C593 diff_6688_20020# gnd! 577.0fF
C594 diff_4192_12940# gnd! 51221.5fF
C595 diff_7516_20284# gnd! 1721.8fF
C596 diff_7744_20500# gnd! 906.8fF
C597 diff_9592_20488# gnd! 1380.9fF
C598 diff_9280_20260# gnd! 812.4fF
C599 diff_8668_20836# gnd! 1116.0fF
C600 diff_5240_19432# gnd! 290.4fF
C601 diff_4928_19444# gnd! 276.4fF
C602 diff_4544_19444# gnd! 286.6fF
C603 diff_4376_19432# gnd! 329.8fF
C604 diff_5152_19192# gnd! 8571.6fF
C605 diff_5308_19396# gnd! 3404.0fF
C606 diff_4456_18616# gnd! 9235.1fF
C607 diff_3868_15448# gnd! 22453.8fF
C608 diff_5084_19444# gnd! 802.3fF
C609 diff_4928_19924# gnd! 290.4fF
C610 diff_4700_19924# gnd! 577.3fF
C611 diff_4996_19156# gnd! 9536.1fF
C612 diff_4576_17684# gnd! 2436.4fF
C613 diff_2212_11356# gnd! 18892.2fF
C614 diff_7084_20800# gnd! 525.4fF
C615 diff_7084_20632# gnd! 2752.1fF
C616 diff_8068_20716# gnd! 1265.4fF
C617 diff_6532_20236# gnd! 4044.9fF
C618 diff_6404_20440# gnd! 718.8fF
C619 diff_9932_21580# gnd! 2172.6fF
C620 diff_5656_20560# gnd! 1397.2fF
C621 diff_5704_20956# gnd! 3196.6fF
C622 diff_16400_21640# gnd! 1190.1fF
C623 diff_14068_21556# gnd! 3814.0fF
C624 diff_14012_21652# gnd! 1122.0fF
C625 diff_13816_22024# gnd! 6646.5fF
C626 diff_18892_22660# gnd! 9400.1fF
C627 diff_17068_22816# gnd! 1775.2fF
C628 diff_16420_22148# gnd! 3565.0fF
C629 diff_16576_22612# gnd! 1773.5fF
C630 diff_16108_22948# gnd! 1800.5fF
C631 diff_15616_22684# gnd! 1791.7fF
C632 diff_15172_22876# gnd! 1791.0fF
C633 diff_14680_22624# gnd! 1781.9fF
C634 diff_13360_22252# gnd! 4520.2fF
C635 diff_11600_22144# gnd! 280.7fF
C636 diff_8764_21368# gnd! 1731.0fF
C637 diff_11000_21736# gnd! 2367.6fF
C638 diff_11216_22036# gnd! 288.0fF
C639 diff_8272_21388# gnd! 1718.6fF
C640 diff_7816_21928# gnd! 1737.2fF
C641 diff_2104_10732# gnd! 28308.2fF
C642 diff_7324_21436# gnd! 1801.8fF
C643 diff_8344_22228# gnd! 2010.9fF
C644 diff_11512_22108# gnd! 606.0fF
C645 diff_11068_22336# gnd! 501.9fF
C646 diff_7492_22216# gnd! 1954.5fF
C647 diff_1696_20020# gnd! 893.2fF
C648 diff_2192_20392# gnd! 429.1fF
C649 diff_1912_20180# gnd! 700.1fF
C650 diff_2068_14080# gnd! 20587.0fF
C651 diff_1840_19936# gnd! 46798.6fF
C652 diff_3052_21280# gnd! 2248.5fF
C653 diff_3500_21460# gnd! 1646.3fF
C654 diff_11020_22492# gnd! 3217.0fF
C655 diff_11708_22792# gnd! 571.5fF
C656 diff_9932_21748# gnd! 2201.5fF
C657 diff_11224_22636# gnd! 1870.0fF
C658 diff_11000_22924# gnd! 1987.2fF
C659 diff_14236_22696# gnd! 1780.2fF
C660 diff_13744_22612# gnd! 1808.4fF
C661 diff_14320_23620# gnd! 3648.9fF
C662 diff_7840_22408# gnd! 2313.1fF
C663 diff_7492_22408# gnd! 2490.9fF
C664 diff_3872_22168# gnd! 1496.3fF
C665 diff_2392_18688# gnd! 24980.3fF
C666 diff_2072_21376# gnd! 1265.7fF
C667 diff_2344_20804# gnd! 1835.7fF
C668 diff_2284_21260# gnd! 1253.1fF
C669 diff_5824_22268# gnd! 490.8fF
C670 diff_6580_22360# gnd! 502.5fF
C671 diff_6208_22352# gnd! 486.8fF
C672 diff_12916_19724# gnd! 4302.4fF
C673 diff_11600_23524# gnd! 281.9fF
C674 diff_13352_23512# gnd! 3660.6fF
C675 diff_11512_23488# gnd! 595.9fF
C676 diff_10516_20840# gnd! 2718.6fF
C677 diff_11216_23416# gnd! 288.2fF
C678 diff_8740_22024# gnd! 2539.0fF
C679 diff_8320_21824# gnd! 2437.9fF
C680 diff_11068_23716# gnd! 488.7fF
C681 diff_13816_24004# gnd! 4290.4fF
C682 diff_14812_24004# gnd! 3567.7fF
C683 diff_13816_24208# gnd! 4015.8fF
C684 diff_18340_24112# gnd! 2647.9fF
C685 diff_8968_23872# gnd! 1650.4fF
C686 diff_6952_20728# gnd! 4666.4fF
C687 diff_3460_23104# gnd! 1224.3fF
C688 diff_6400_21080# gnd! 4155.3fF
C689 diff_7768_23620# gnd! 2530.5fF
C690 diff_7288_23632# gnd! 2638.1fF
C691 diff_8380_23308# gnd! 1081.8fF
C692 diff_7768_23848# gnd! 1175.8fF
C693 diff_7180_23308# gnd! 1425.7fF
C694 diff_4156_19880# gnd! 4413.1fF
C695 diff_13792_23696# gnd! 2083.6fF
C696 diff_11708_24184# gnd! 571.3fF
C697 diff_9412_21556# gnd! 2913.6fF
C698 diff_12848_24340# gnd! 1343.0fF
C699 diff_13816_24448# gnd! 1644.3fF
C700 diff_15472_24352# gnd! 3639.8fF
C701 diff_17068_23276# gnd! 3300.1fF
C702 diff_16636_23048# gnd! 3165.8fF
C703 diff_17668_25588# gnd! 1332.6fF
C704 diff_16120_23288# gnd! 3033.2fF
C705 diff_15676_23048# gnd! 3071.2fF
C706 diff_17092_24928# gnd! 1325.3fF
C707 diff_16504_25588# gnd! 1338.0fF
C708 diff_12848_24544# gnd! 1375.7fF
C709 diff_15124_23692# gnd! 2959.7fF
C710 diff_14740_23060# gnd! 2992.7fF
C711 diff_15928_24928# gnd! 1309.3fF
C712 diff_15328_25624# gnd! 1283.9fF
C713 diff_11600_24700# gnd! 291.8fF
C714 diff_11216_24704# gnd! 289.3fF
C715 diff_11000_24316# gnd! 2610.4fF
C716 diff_11512_24664# gnd! 687.5fF
C717 diff_11068_25000# gnd! 558.6fF
C718 diff_9392_24340# gnd! 224.6fF
C719 diff_8636_24304# gnd! 225.7fF
C720 diff_8264_24380# gnd! 242.0fF
C721 diff_9212_24604# gnd! 361.9fF
C722 diff_8704_24304# gnd! 357.2fF
C723 diff_9392_24904# gnd! 210.6fF
C724 diff_11020_25156# gnd! 3370.7fF
C725 diff_13972_25108# gnd! 11208.6fF
C726 diff_14164_25384# gnd! 2972.6fF
C727 diff_13708_25372# gnd! 2183.4fF
C728 diff_7508_24316# gnd! 217.7fF
C729 diff_8096_24604# gnd! 344.9fF
C730 diff_7588_24304# gnd! 345.7fF
C731 diff_9212_24748# gnd! 360.1fF
C732 diff_14752_24940# gnd! 1280.2fF
C733 diff_14164_25600# gnd! 1286.0fF
C734 diff_11708_25456# gnd! 583.0fF
C735 diff_9412_21772# gnd! 3306.4fF
C736 diff_13484_25336# gnd! 1357.4fF
C737 diff_13720_25264# gnd! 9350.7fF
C738 diff_17948_26108# gnd! 187.5fF
C739 diff_17204_26068# gnd! 214.0fF
C740 diff_17780_26356# gnd! 409.1fF
C741 diff_17272_26056# gnd! 373.9fF
C742 diff_16832_26180# gnd! 199.3fF
C743 diff_16076_26068# gnd! 231.9fF
C744 diff_15716_26116# gnd! 230.1fF
C745 diff_16664_26368# gnd! 367.6fF
C746 diff_16156_26056# gnd! 352.6fF
C747 diff_17948_26656# gnd! 213.6fF
C748 diff_17780_26512# gnd! 377.1fF
C749 diff_17948_26996# gnd! 178.7fF
C750 diff_17192_26816# gnd! 206.9fF
C751 diff_16832_26656# gnd! 213.1fF
C752 diff_14960_26068# gnd! 237.1fF
C753 diff_14600_26116# gnd! 229.4fF
C754 diff_11224_25648# gnd! 1894.5fF
C755 diff_10976_25588# gnd! 2062.2fF
C756 diff_15548_26368# gnd! 350.7fF
C757 diff_15040_26056# gnd! 339.5fF
C758 diff_17260_26836# gnd! 377.2fF
C759 diff_16664_26512# gnd! 357.9fF
C760 diff_16156_26512# gnd! 358.9fF
C761 diff_16076_26804# gnd! 207.1fF
C762 diff_15716_26668# gnd! 219.2fF
C763 diff_13844_26080# gnd! 209.8fF
C764 diff_14420_26368# gnd! 352.7fF
C765 diff_13912_26068# gnd! 355.8fF
C766 diff_15548_26512# gnd! 350.4fF
C767 diff_17192_26956# gnd! 212.5fF
C768 diff_16832_27004# gnd! 208.4fF
C769 diff_17780_27256# gnd! 376.4fF
C770 diff_17272_26944# gnd! 359.9fF
C771 diff_16076_26956# gnd! 235.1fF
C772 diff_15716_27004# gnd! 223.2fF
C773 diff_14960_26816# gnd! 219.2fF
C774 diff_14600_26668# gnd! 219.0fF
C775 diff_15028_26836# gnd! 377.6fF
C776 diff_16664_27256# gnd! 356.8fF
C777 diff_16144_26956# gnd! 350.3fF
C778 diff_17948_27544# gnd! 184.6fF
C779 diff_17780_27400# gnd! 382.7fF
C780 diff_17948_27880# gnd! 172.2fF
C781 diff_17192_27692# gnd! 231.7fF
C782 diff_16832_27556# gnd! 199.0fF
C783 diff_17272_27400# gnd! 337.6fF
C784 diff_14420_26524# gnd! 336.7fF
C785 diff_14960_26968# gnd! 228.6fF
C786 diff_14600_27004# gnd! 214.4fF
C787 diff_13844_26816# gnd! 209.8fF
C788 diff_12256_26224# gnd! 5236.7fF
C789 diff_13912_26836# gnd! 359.5fF
C790 diff_15548_27256# gnd! 353.6fF
C791 diff_15040_26944# gnd! 356.0fF
C792 diff_16664_27400# gnd! 357.5fF
C793 diff_16076_27692# gnd! 216.7fF
C794 diff_15716_27556# gnd! 209.8fF
C795 diff_16144_27724# gnd! 345.5fF
C796 diff_9392_25228# gnd! 219.0fF
C797 diff_8636_25028# gnd! 209.2fF
C798 diff_3856_18340# gnd! 6716.8fF
C799 diff_3952_23104# gnd! 575.3fF
C800 diff_3200_23188# gnd! 1293.2fF
C801 diff_4052_23284# gnd! 617.2fF
C802 diff_2140_4552# gnd! 31467.3fF
C803 diff_4436_22444# gnd! 3581.5fF
C804 diff_1232_22576# gnd! 4977.9fF
C805 cm_rom gnd! 14688.0fF
C806 diff_2140_5752# gnd! 32790.8fF
C807 diff_3952_23632# gnd! 507.3fF
C808 diff_3508_23020# gnd! 1071.8fF
C809 clk1 gnd! 66880.3fF
C810 clk2 gnd! 80492.1fF
C811 diff_1132_21544# gnd! 33238.8fF
C812 diff_4700_19432# gnd! 5768.2fF
C813 diff_6584_24388# gnd! 3673.1fF
C814 diff_8276_24904# gnd! 210.6fF
C815 diff_8704_25072# gnd! 363.4fF
C816 diff_8096_24748# gnd! 352.4fF
C817 diff_7508_25052# gnd! 217.7fF
C818 diff_4040_23804# gnd! 652.3fF
C819 diff_5792_24436# gnd! 3279.4fF
C820 diff_5428_24556# gnd! 3845.4fF
C821 diff_7588_25072# gnd! 346.6fF
C822 diff_6160_24964# gnd! 3642.9fF
C823 diff_8264_25240# gnd! 230.1fF
C824 diff_8636_25192# gnd! 225.0fF
C825 diff_9212_25492# gnd! 358.0fF
C826 diff_8704_25192# gnd! 344.1fF
C827 diff_7508_25192# gnd! 232.4fF
C828 diff_8096_25492# gnd! 340.4fF
C829 diff_9392_25792# gnd! 222.3fF
C830 diff_7588_25192# gnd! 352.6fF
C831 diff_9212_25636# gnd! 352.0fF
C832 diff_12236_26380# gnd! 4405.1fF
C833 diff_11800_26332# gnd! 4724.2fF
C834 diff_12680_26680# gnd! 4939.2fF
C835 diff_13844_26968# gnd! 212.1fF
C836 diff_14420_27256# gnd! 356.1fF
C837 diff_13912_26956# gnd! 357.4fF
C838 diff_15536_27428# gnd! 349.2fF
C839 diff_17192_27844# gnd! 229.2fF
C840 diff_16832_27892# gnd! 181.6fF
C841 diff_17780_28132# gnd! 414.9fF
C842 diff_17272_27832# gnd! 354.9fF
C843 diff_17948_28432# gnd! 180.6fF
C844 diff_16076_27844# gnd! 235.3fF
C845 diff_15716_27892# gnd! 201.7fF
C846 diff_14960_27692# gnd! 214.4fF
C847 diff_14600_27556# gnd! 214.4fF
C848 diff_15028_27712# gnd! 343.0fF
C849 diff_12680_27040# gnd! 5083.0fF
C850 diff_14420_27400# gnd! 361.9fF
C851 diff_16652_28144# gnd! 364.7fF
C852 diff_16144_27832# gnd! 339.4fF
C853 diff_17780_28288# gnd! 390.0fF
C854 diff_14960_27844# gnd! 226.9fF
C855 diff_13844_27692# gnd! 212.1fF
C856 diff_13912_27712# gnd! 340.5fF
C857 diff_14588_28028# gnd! 215.7fF
C858 diff_15536_28144# gnd! 362.3fF
C859 diff_15028_27832# gnd! 343.2fF
C860 diff_17192_28580# gnd! 223.0fF
C861 diff_17948_28768# gnd! 169.9fF
C862 diff_17272_28288# gnd! 339.4fF
C863 diff_16832_28432# gnd! 184.6fF
C864 diff_16652_28288# gnd! 371.8fF
C865 diff_17192_28732# gnd! 227.5fF
C866 diff_16832_28768# gnd! 174.5fF
C867 diff_16076_28580# gnd! 224.6fF
C868 diff_15704_28432# gnd! 222.8fF
C869 diff_13832_27860# gnd! 216.9fF
C870 diff_14420_28144# gnd! 350.4fF
C871 diff_13912_27832# gnd! 355.1fF
C872 diff_16144_28612# gnd! 335.3fF
C873 diff_15536_28288# gnd! 354.6fF
C874 diff_17780_29020# gnd! 411.2fF
C875 diff_17272_28708# gnd! 366.5fF
C876 diff_17632_26752# gnd! 3352.2fF
C877 diff_17440_26356# gnd! 3268.7fF
C878 diff_14948_28604# gnd! 219.4fF
C879 diff_14588_28444# gnd! 225.2fF
C880 diff_15028_28612# gnd! 349.7fF
C881 diff_14420_28288# gnd! 341.9fF
C882 diff_16076_28732# gnd! 216.7fF
C883 diff_15716_28780# gnd! 179.8fF
C884 diff_16652_29032# gnd! 388.0fF
C885 diff_16144_28720# gnd! 342.4fF
C886 diff_16516_26800# gnd! 3145.0fF
C887 diff_16312_25436# gnd! 3261.6fF
C888 diff_17948_29320# gnd! 169.3fF
C889 diff_17780_29176# gnd! 388.3fF
C890 diff_17932_25436# gnd! 3473.2fF
C891 diff_17152_20864# gnd! 7361.2fF
C892 diff_17192_29468# gnd! 186.9fF
C893 diff_14948_28736# gnd! 217.7fF
C894 diff_14588_28784# gnd! 219.6fF
C895 diff_13832_28604# gnd! 214.6fF
C896 diff_12236_27076# gnd! 4444.4fF
C897 diff_10996_26404# gnd! 1077.2fF
C898 diff_11180_26776# gnd! 2420.2fF
C899 diff_9392_26120# gnd! 218.2fF
C900 diff_8636_25916# gnd! 237.6fF
C901 diff_8264_25820# gnd! 246.5fF
C902 diff_8704_25960# gnd! 337.5fF
C903 diff_8096_25636# gnd! 340.5fF
C904 diff_8636_26080# gnd! 241.9fF
C905 diff_7508_25952# gnd! 210.8fF
C906 diff_7588_25948# gnd! 352.3fF
C907 diff_8264_26128# gnd! 258.8fF
C908 diff_9212_26380# gnd! 365.0fF
C909 diff_8704_26080# gnd! 348.4fF
C910 diff_7508_26080# gnd! 232.4fF
C911 diff_8096_26380# gnd! 321.5fF
C912 diff_7588_26080# gnd! 349.1fF
C913 diff_9392_26668# gnd! 230.7fF
C914 diff_9212_26524# gnd! 358.9fF
C915 diff_12256_27580# gnd! 5214.7fF
C916 diff_12256_27952# gnd! 5186.5fF
C917 diff_12680_28456# gnd! 4948.8fF
C918 diff_11180_26992# gnd! 2565.3fF
C919 diff_11800_27280# gnd! 4750.2fF
C920 diff_10996_27364# gnd! 1114.0fF
C921 diff_9392_27008# gnd! 234.6fF
C922 diff_8624_26828# gnd! 237.8fF
C923 diff_8264_26680# gnd! 247.6fF
C924 diff_8704_26848# gnd! 348.6fF
C925 diff_6152_25264# gnd! 3679.1fF
C926 diff_6152_25792# gnd! 3654.9fF
C927 diff_8096_26524# gnd! 322.2fF
C928 diff_8636_26968# gnd! 253.2fF
C929 diff_8276_27004# gnd! 235.3fF
C930 diff_7588_26848# gnd! 355.4fF
C931 diff_7508_26840# gnd! 208.4fF
C932 diff_6172_26164# gnd! 3704.8fF
C933 diff_6572_26696# gnd! 3588.8fF
C934 diff_9212_27268# gnd! 353.9fF
C935 diff_8704_26968# gnd! 331.8fF
C936 diff_7508_26968# gnd! 225.5fF
C937 diff_8096_27268# gnd! 348.8fF
C938 diff_7588_26968# gnd! 362.8fF
C939 diff_6584_27052# gnd! 3616.6fF
C940 diff_9392_27568# gnd! 226.9fF
C941 diff_9212_27412# gnd! 346.7fF
C942 diff_13900_28612# gnd! 352.1fF
C943 diff_15536_29032# gnd! 372.6fF
C944 diff_15028_28720# gnd! 349.8fF
C945 diff_13832_28732# gnd! 227.8fF
C946 diff_14420_29032# gnd! 364.5fF
C947 diff_13900_28732# gnd! 352.8fF
C948 diff_15388_25448# gnd! 3104.3fF
C949 diff_15148_25448# gnd! 3104.9fF
C950 diff_14224_25448# gnd! 3100.4fF
C951 diff_13972_25448# gnd! 3126.1fF
C952 diff_16832_29320# gnd! 177.2fF
C953 diff_17248_29488# gnd! 392.4fF
C954 diff_16652_29176# gnd! 402.1fF
C955 diff_17092_28684# gnd! 3342.2fF
C956 diff_16768_25436# gnd! 3320.7fF
C957 diff_16076_29492# gnd! 189.2fF
C958 diff_15716_29332# gnd! 175.8fF
C959 diff_16132_29488# gnd! 373.3fF
C960 diff_15536_29176# gnd! 394.4fF
C961 diff_15976_29452# gnd! 3210.1fF
C962 diff_15592_25448# gnd! 3308.0fF
C963 diff_14960_29468# gnd! 216.7fF
C964 diff_14600_29332# gnd! 180.4fF
C965 diff_15028_29188# gnd! 355.8fF
C966 diff_14860_29452# gnd! 3171.9fF
C967 diff_14420_29176# gnd! 387.8fF
C968 diff_14416_25448# gnd! 3208.7fF
C969 diff_13912_29200# gnd! 391.6fF
C970 diff_13844_29468# gnd! 189.8fF
C971 diff_12680_28816# gnd! 5014.9fF
C972 diff_12544_25804# gnd! 7678.2fF
C973 diff_12236_28156# gnd! 4419.9fF
C974 diff_9392_27908# gnd! 242.4fF
C975 diff_8636_27692# gnd! 235.3fF
C976 diff_8276_27568# gnd! 213.1fF
C977 diff_8704_27736# gnd! 340.6fF
C978 diff_8096_27412# gnd! 349.9fF
C979 diff_11800_28096# gnd! 4553.9fF
C980 diff_10996_28180# gnd! 1068.9fF
C981 diff_8636_27856# gnd! 250.9fF
C982 diff_8264_27920# gnd! 229.4fF
C983 diff_7588_27736# gnd! 369.6fF
C984 diff_7520_27716# gnd! 200.6fF
C985 diff_9224_28156# gnd! 349.8fF
C986 diff_8704_27856# gnd! 333.0fF
C987 diff_11180_28552# gnd! 2448.5fF
C988 diff_7508_27856# gnd! 225.7fF
C989 diff_8096_28156# gnd! 345.0fF
C990 diff_7588_27856# gnd! 370.2fF
C991 diff_9392_28444# gnd! 241.7fF
C992 diff_9224_28300# gnd! 340.0fF
C993 diff_12236_28852# gnd! 4438.4fF
C994 diff_12136_25792# gnd! 10485.9fF
C995 diff_9392_28796# gnd! 235.3fF
C996 diff_8636_28604# gnd! 242.4fF
C997 diff_8276_28444# gnd! 239.4fF
C998 diff_8716_28612# gnd! 334.1fF
C999 diff_11788_29092# gnd! 4776.6fF
C1000 diff_10996_29140# gnd! 1060.7fF
C1001 diff_11872_25876# gnd! 8356.1fF
C1002 diff_11180_28768# gnd! 2654.9fF
C1003 diff_12256_29344# gnd! 5048.5fF
C1004 diff_12328_25804# gnd! 7045.1fF
C1005 diff_13744_27736# gnd! 3224.4fF
C1006 diff_8096_28300# gnd! 343.7fF
C1007 diff_8636_28744# gnd! 254.0fF
C1008 diff_8276_28780# gnd! 241.9fF
C1009 diff_7520_28604# gnd! 198.5fF
C1010 diff_7588_28636# gnd! 373.9fF
C1011 diff_9224_29044# gnd! 358.4fF
C1012 diff_8704_28756# gnd! 342.2fF
C1013 diff_9028_23696# gnd! 4156.4fF
C1014 diff_8788_23696# gnd! 4265.1fF
C1015 diff_7508_28748# gnd! 225.5fF
C1016 diff_8096_29044# gnd! 350.4fF
C1017 diff_7588_28744# gnd! 376.8fF
C1018 diff_7816_23824# gnd! 4362.3fF
C1019 diff_7576_23716# gnd! 4312.6fF
C1020 diff_9392_29332# gnd! 234.9fF
C1021 diff_8680_20596# gnd! 8503.7fF
C1022 diff_9224_29188# gnd! 314.9fF
C1023 diff_9232_23696# gnd! 4449.1fF
C1024 diff_8636_29492# gnd! 186.9fF
C1025 diff_8276_29332# gnd! 226.9fF
C1026 diff_8704_29524# gnd! 385.2fF
C1027 diff_8096_29188# gnd! 322.6fF
C1028 diff_8548_23696# gnd! 4339.1fF
C1029 diff_8020_23696# gnd! 4378.6fF
C1030 diff_2836_23896# gnd! 1844.7fF
C1031 diff_928_16456# gnd! 16476.2fF
C1032 diff_928_20116# gnd! 8982.9fF
C1033 diff_2788_24040# gnd! 2714.3fF
C1034 diff_4204_24416# gnd! 4328.1fF
C1035 diff_3656_24604# gnd! 1303.4fF
C1036 diff_3608_24316# gnd! 1402.5fF
C1037 diff_4072_24796# gnd! 1206.7fF
C1038 diff_5396_25448# gnd! 3553.2fF
C1039 diff_2680_25420# gnd! 1966.8fF
C1040 diff_2476_25408# gnd! 1614.0fF
C1041 diff_2428_25492# gnd! 3012.4fF
C1042 diff_5408_25636# gnd! 3621.9fF
C1043 diff_5780_26516# gnd! 3384.3fF
C1044 diff_5428_26392# gnd! 3759.6fF
C1045 diff_5792_27100# gnd! 3307.4fF
C1046 diff_5428_27220# gnd! 3745.6fF
C1047 diff_6172_27580# gnd! 3723.2fF
C1048 diff_6164_27928# gnd! 3716.1fF
C1049 diff_6176_28456# gnd! 3673.2fF
C1050 diff_5144_23548# gnd! 5052.6fF
C1051 diff_6160_28852# gnd! 3701.9fF
C1052 diff_6020_23524# gnd! 4652.5fF
C1053 diff_2980_25568# gnd! 164.3fF
C1054 diff_2680_25568# gnd! 220.4fF
C1055 diff_2476_25568# gnd! 122.2fF
C1056 diff_2428_25648# gnd! 3157.0fF
C1057 diff_4072_26372# gnd! 1174.4fF
C1058 diff_4204_26720# gnd! 4265.2fF
C1059 diff_3136_26020# gnd! 2568.9fF
C1060 diff_3656_26524# gnd! 1352.2fF
C1061 diff_4204_27092# gnd! 4326.6fF
C1062 diff_3656_27268# gnd! 1338.2fF
C1063 diff_472_25516# gnd! 1015.6fF
C1064 diff_424_25492# gnd! 7981.9fF
C1065 diff_460_26224# gnd! 1025.9fF
C1066 diff_2984_25724# gnd! 2432.9fF
C1067 diff_5408_27856# gnd! 3484.4fF
C1068 diff_4084_27448# gnd! 1217.8fF
C1069 sync gnd! 26071.8fF
C1070 diff_424_25960# gnd! 10369.9fF
C1071 diff_2680_25724# gnd! 1548.4fF
C1072 diff_2476_25724# gnd! 1750.0fF
C1073 diff_2728_27904# gnd! 2788.2fF
C1074 diff_5408_28300# gnd! 3604.3fF
C1075 diff_5020_23836# gnd! 6213.5fF
C1076 diff_2740_24880# gnd! 5092.6fF
C1077 diff_2764_28012# gnd! 1221.7fF
C1078 diff_7520_29516# gnd! 210.0fF
C1079 diff_3088_28840# gnd! 2191.0fF
C1080 diff_4076_29024# gnd! 1282.2fF
C1081 diff_6496_23704# gnd! 5139.5fF
C1082 diff_5200_22772# gnd! 5874.6fF
C1083 diff_5212_23848# gnd! 5723.3fF
C1084 diff_5404_29068# gnd! 3723.9fF
C1085 Vdd gnd! 636263.0fF
C1086 diff_4204_29396# gnd! 4496.4fF
C1087 diff_7588_29524# gnd! 379.3fF
C1088 diff_7348_23696# gnd! 4432.5fF
C1089 diff_5792_29180# gnd! 3585.1fF
C1090 diff_6584_29296# gnd! 3685.2fF
C1091 diff_2860_29380# gnd! 2725.5fF
C1092 diff_3668_29188# gnd! 1320.0fF
C1093 diff_2656_22088# gnd! 11906.6fF
C1094 diff_3808_28348# gnd! 41154.0fF
C1095 diff_3436_29560# gnd! 42619.3fF
C1096 diff_3244_29488# gnd! 45673.5fF
C1097 diff_3040_29500# gnd! 46518.8fF
C1098 test gnd! 22334.6fF
C1099 reset gnd! 22637.5fF
