* SPICE3 file created from 4001.ext - technology: nmos

.option scale=0.001u

M1000 clk2 GND GND GND efet w=119880 l=8880
+ ad=1.91522e+09 pd=1.9092e+06 as=6.08391e+08 ps=4.84848e+07 
M1001 clk1 GND GND GND efet w=119880 l=8880
+ ad=-1.41856e+09 pd=1.45928e+06 as=0 ps=0 
M1002 d2 GND d2 GND efet w=218300 l=138380
+ ad=1.28561e+09 pd=3.69408e+06 as=0 ps=0 
M1003 d3 GND d3 GND efet w=220520 l=142080
+ ad=-8.99595e+08 pd=5.05568e+06 as=0 ps=0 
M1004 sync GND GND GND efet w=112480 l=8880
+ ad=-1.30823e+09 pd=3.22936e+06 as=0 ps=0 
M1005 GND diff_417360_2049800# d3 GND efet w=1151440 l=4440
+ ad=0 pd=0 as=0 ps=0 
M1006 GND diff_609760_2049800# d2 GND efet w=1149960 l=4440
+ ad=0 pd=0 as=0 ps=0 
M1007 Vdd diff_438080_1685720# d3 GND efet w=532060 l=12580
+ ad=-1.58224e+09 pd=1.88197e+07 as=0 ps=0 
M1008 GND diff_800680_2049800# d1 GND efet w=1149960 l=4440
+ ad=0 pd=0 as=1.15638e+09 ps=3.7444e+06 
M1009 GND diff_991600_2049800# d0 GND efet w=1149960 l=4440
+ ad=0 pd=0 as=9.43908e+08 ps=3.72072e+06 
M1010 GND diff_3001440_2148960# diff_3005880_2094200# GND efet w=439560 l=7400
+ ad=0 pd=0 as=1.24975e+09 ps=1.8204e+06 
M1011 GND clk1 diff_3223440_2120840# GND efet w=31080 l=8880
+ ad=0 pd=0 as=6.81214e+08 ps=112480 
M1012 GND sync diff_3001440_2148960# GND efet w=94720 l=8880
+ ad=0 pd=0 as=1.7783e+08 ps=748880 
M1013 diff_3455800_2137120# diff_3393640_2079400# GND GND efet w=34040 l=7400
+ ad=8.06067e+08 pd=224960 as=0 ps=0 
M1014 diff_3267840_1761200# diff_3455800_2137120# GND GND efet w=50320 l=7400
+ ad=1.16091e+09 pd=251600 as=0 ps=0 
M1015 GND diff_3001440_2148960# diff_3383280_2114920# GND efet w=50320 l=7400
+ ad=0 pd=0 as=5.95789e+08 ps=124320 
M1016 diff_3223440_2120840# Vdd Vdd GND efet w=8880 l=11840
+ ad=0 pd=0 as=0 ps=0 
M1017 diff_3001440_2148960# diff_3285600_2079400# GND GND efet w=57720 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1018 GND diff_1237280_2100120# diff_1243200_2079400# GND efet w=763680 l=8880
+ ad=0 pd=0 as=-5.38179e+08 ps=3.42768e+06 
M1019 Vdd diff_2043880_2100120# diff_1243200_2079400# GND efet w=793280 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1020 diff_1243200_2079400# diff_1238760_2072000# diff_1243200_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1021 diff_1243200_2079400# diff_1238760_2072000# diff_1268360_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1022 diff_1243200_2079400# diff_1238760_2072000# diff_1293520_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1023 diff_1243200_2079400# diff_1238760_2072000# diff_1318680_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1024 diff_1243200_2079400# diff_1238760_2072000# diff_1343840_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1025 diff_1243200_2079400# diff_1238760_2072000# diff_1369000_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1026 diff_1243200_2079400# diff_1238760_2072000# diff_1394160_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1027 diff_1243200_2079400# diff_1238760_2072000# diff_1419320_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1028 diff_1243200_2079400# diff_1238760_2072000# diff_1444480_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1029 diff_1243200_2079400# diff_1238760_2072000# diff_1469640_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1030 diff_1243200_2079400# diff_1238760_2072000# diff_1494800_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1031 diff_1243200_2079400# diff_1238760_2072000# diff_1519960_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1032 diff_1243200_2079400# diff_1238760_2072000# diff_1545120_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1033 diff_1243200_2079400# diff_1238760_2072000# diff_1570280_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1034 diff_1243200_2079400# diff_1238760_2072000# diff_1595440_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1035 diff_1243200_2079400# diff_1238760_2072000# diff_1620600_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1036 diff_1243200_2079400# diff_1238760_2072000# diff_1645760_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1037 diff_1243200_2079400# diff_1238760_2072000# diff_1670920_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1038 diff_1243200_2079400# diff_1238760_2072000# diff_1696080_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1039 diff_1243200_2079400# diff_1238760_2072000# diff_1721240_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1040 diff_1243200_2079400# diff_1238760_2072000# diff_1746400_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1041 diff_1243200_2079400# diff_1238760_2072000# diff_1771560_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1042 diff_1243200_2079400# diff_1238760_2072000# diff_1796720_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1043 diff_1243200_2079400# diff_1238760_2072000# diff_1821880_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1044 diff_1243200_2079400# diff_1238760_2072000# diff_1847040_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1045 diff_1243200_2079400# diff_1238760_2072000# diff_1872200_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1046 diff_1243200_2079400# diff_1238760_2072000# diff_1897360_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1047 diff_1243200_2079400# diff_1238760_2072000# diff_1922520_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1048 diff_1243200_2079400# diff_1238760_2072000# diff_1947680_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1049 diff_1243200_2079400# diff_1238760_2072000# diff_1972840_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1050 diff_1243200_2079400# diff_1238760_2072000# diff_1998000_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1051 diff_1243200_2079400# diff_1238760_2072000# diff_2023160_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1052 diff_1243200_2079400# diff_1238760_2072000# diff_2048320_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1053 diff_1243200_2079400# diff_1238760_2072000# diff_2073480_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1054 diff_1243200_2079400# diff_1238760_2072000# diff_2098640_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1055 diff_1243200_2079400# diff_1238760_2072000# diff_2123800_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1056 diff_1243200_2079400# diff_1238760_2072000# diff_2148960_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1057 diff_1243200_2079400# diff_1238760_2072000# diff_2174120_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1058 diff_1243200_2079400# diff_1238760_2072000# diff_2199280_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1059 diff_1243200_2079400# diff_1238760_2072000# diff_2224440_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1060 diff_1243200_2079400# diff_1238760_2072000# diff_2249600_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1061 diff_1243200_2079400# diff_1238760_2072000# diff_2274760_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1062 diff_1243200_2079400# diff_1238760_2072000# diff_2299920_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1063 diff_1243200_2079400# diff_1238760_2072000# diff_2325080_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1064 diff_1243200_2079400# diff_1238760_2072000# diff_2350240_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1065 diff_1243200_2079400# diff_1238760_2072000# diff_2375400_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1066 diff_1243200_2079400# diff_1238760_2072000# diff_2400560_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1067 diff_1243200_2079400# diff_1238760_2072000# diff_2425720_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1068 diff_1243200_2079400# diff_1238760_2072000# diff_2450880_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1069 diff_1243200_2079400# diff_1238760_2072000# diff_2476040_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1070 diff_1243200_2079400# diff_1238760_2072000# diff_2501200_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1071 diff_1243200_2079400# diff_1238760_2072000# diff_2526360_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1072 diff_1243200_2079400# diff_1238760_2072000# diff_2551520_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1073 diff_1243200_2079400# diff_1238760_2072000# diff_2576680_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1074 diff_1243200_2079400# diff_1238760_2072000# diff_2601840_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1075 diff_1243200_2079400# diff_1238760_2072000# diff_2627000_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1076 diff_1243200_2079400# diff_1238760_2072000# diff_2652160_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1077 diff_1243200_2079400# diff_1238760_2072000# diff_2677320_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1078 diff_1243200_2079400# diff_1238760_2072000# diff_2702480_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1079 diff_1243200_2079400# diff_1238760_2072000# diff_2727640_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1080 diff_1243200_2079400# diff_1238760_2072000# diff_2752800_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1081 diff_1243200_2079400# diff_1238760_2072000# diff_2777960_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1082 diff_1243200_2079400# diff_1238760_2072000# diff_2803120_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1083 diff_1243200_2079400# diff_1238760_2072000# diff_2828280_2051280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1084 diff_2920040_2064600# diff_2912640_526880# diff_1238760_2072000# GND efet w=110260 l=8880
+ ad=1.2117e+09 pd=849520 as=1.45443e+09 ps=284160 
M1085 Vdd Vdd diff_451400_1855920# GND efet w=11840 l=11840
+ ad=0 pd=0 as=3.78939e+08 ps=88800 
M1086 Vdd Vdd diff_528360_1858880# GND efet w=10360 l=13320
+ ad=0 pd=0 as=3.02275e+08 ps=82880 
M1087 diff_451400_1855920# diff_451400_1855920# diff_451400_1855920# GND efet w=2220 l=4440
+ ad=0 pd=0 as=0 ps=0 
M1088 Vdd diff_451400_1855920# diff_438080_1685720# GND efet w=10360 l=8880
+ ad=0 pd=0 as=3.07063e+08 ps=802160 
M1089 Vdd diff_528360_1858880# diff_417360_2049800# GND efet w=10360 l=8880
+ ad=0 pd=0 as=1.3256e+09 ps=947200 
M1090 diff_528360_1858880# diff_528360_1858880# diff_528360_1858880# GND efet w=2220 l=5920
+ ad=0 pd=0 as=0 ps=0 
M1091 Vdd diff_629000_1685720# d2 GND efet w=529840 l=13320
+ ad=0 pd=0 as=0 ps=0 
M1092 diff_451400_1855920# diff_451400_1855920# diff_451400_1855920# GND efet w=1480 l=4440
+ ad=0 pd=0 as=0 ps=0 
M1093 diff_438080_1685720# diff_451400_1855920# diff_438080_1685720# GND efet w=52540 l=17020
+ ad=0 pd=0 as=0 ps=0 
M1094 diff_528360_1858880# diff_528360_1858880# diff_528360_1858880# GND efet w=1480 l=7400
+ ad=0 pd=0 as=0 ps=0 
M1095 Vdd Vdd diff_642320_1854440# GND efet w=8880 l=11840
+ ad=0 pd=0 as=3.24179e+08 ps=91760 
M1096 Vdd Vdd diff_719280_1857400# GND efet w=11840 l=13320
+ ad=0 pd=0 as=3.35131e+08 ps=97680 
M1097 diff_642320_1854440# diff_642320_1854440# diff_642320_1854440# GND efet w=2960 l=3700
+ ad=0 pd=0 as=0 ps=0 
M1098 Vdd diff_642320_1854440# diff_629000_1685720# GND efet w=10360 l=8880
+ ad=0 pd=0 as=3.09254e+08 ps=802160 
M1099 Vdd diff_719280_1857400# diff_609760_2049800# GND efet w=10360 l=8880
+ ad=0 pd=0 as=1.41979e+09 ps=950160 
M1100 diff_719280_1857400# diff_719280_1857400# diff_719280_1857400# GND efet w=4440 l=5180
+ ad=0 pd=0 as=0 ps=0 
M1101 diff_642320_1854440# diff_642320_1854440# diff_642320_1854440# GND efet w=1480 l=5920
+ ad=0 pd=0 as=0 ps=0 
M1102 diff_417360_2049800# diff_528360_1858880# diff_417360_2049800# GND efet w=70300 l=8140
+ ad=0 pd=0 as=0 ps=0 
M1103 diff_629000_1685720# diff_642320_1854440# diff_629000_1685720# GND efet w=54020 l=17020
+ ad=0 pd=0 as=0 ps=0 
M1104 diff_719280_1857400# diff_719280_1857400# diff_719280_1857400# GND efet w=1480 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1105 Vdd diff_819920_1684240# d1 GND efet w=531320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1106 Vdd Vdd diff_830280_1857400# GND efet w=10360 l=13320
+ ad=0 pd=0 as=2.69419e+08 ps=79920 
M1107 Vdd Vdd diff_910200_1857400# GND efet w=10360 l=13320
+ ad=0 pd=0 as=2.91323e+08 ps=76960 
M1108 Vdd diff_1012320_1684240# d0 GND efet w=528360 l=12580
+ ad=0 pd=0 as=0 ps=0 
M1109 Vdd diff_830280_1857400# diff_819920_1684240# GND efet w=8880 l=8880
+ ad=0 pd=0 as=3.53062e+08 ps=858400 
M1110 diff_830280_1857400# diff_830280_1857400# diff_830280_1857400# GND efet w=2960 l=5920
+ ad=0 pd=0 as=0 ps=0 
M1111 diff_609760_2049800# diff_719280_1857400# diff_609760_2049800# GND efet w=70300 l=8140
+ ad=0 pd=0 as=0 ps=0 
M1112 Vdd diff_910200_1857400# diff_800680_2049800# GND efet w=9620 l=9620
+ ad=0 pd=0 as=1.26646e+09 ps=944240 
M1113 diff_910200_1857400# diff_910200_1857400# diff_910200_1857400# GND efet w=1480 l=2220
+ ad=0 pd=0 as=0 ps=0 
M1114 diff_830280_1857400# diff_830280_1857400# diff_830280_1857400# GND efet w=1480 l=5920
+ ad=0 pd=0 as=0 ps=0 
M1115 diff_910200_1857400# diff_910200_1857400# diff_910200_1857400# GND efet w=740 l=2220
+ ad=0 pd=0 as=0 ps=0 
M1116 Vdd Vdd diff_1025640_1855920# GND efet w=10360 l=11840
+ ad=0 pd=0 as=3.3075e+08 ps=82880 
M1117 Vdd Vdd diff_1093720_1907720# GND efet w=10360 l=11840
+ ad=0 pd=0 as=2.7161e+08 ps=74000 
M1118 diff_1025640_1855920# diff_1025640_1855920# diff_1025640_1855920# GND efet w=740 l=2220
+ ad=0 pd=0 as=0 ps=0 
M1119 Vdd diff_1025640_1855920# diff_1012320_1684240# GND efet w=8880 l=8880
+ ad=0 pd=0 as=3.37729e+08 ps=799200 
M1120 Vdd diff_1093720_1907720# diff_991600_2049800# GND efet w=8880 l=8880
+ ad=0 pd=0 as=1.36284e+09 ps=923520 
M1121 diff_1093720_1907720# diff_1093720_1907720# diff_1093720_1907720# GND efet w=1480 l=2220
+ ad=0 pd=0 as=0 ps=0 
M1122 diff_1243200_2051280# diff_1238760_2043880# diff_1243200_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1123 diff_1268360_2051280# diff_1238760_2043880# diff_1268360_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1124 diff_1293520_2051280# diff_1238760_2043880# diff_1293520_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1125 diff_1318680_2051280# diff_1238760_2043880# diff_1318680_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1126 diff_1343840_2051280# diff_1238760_2043880# diff_1343840_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1127 diff_1369000_2051280# diff_1238760_2043880# diff_1369000_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1128 diff_1394160_2051280# diff_1238760_2043880# diff_1394160_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1129 diff_1419320_2051280# diff_1238760_2043880# diff_1419320_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1130 diff_1444480_2051280# diff_1238760_2043880# diff_1444480_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1131 diff_1469640_2051280# diff_1238760_2043880# diff_1469640_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1132 diff_1494800_2051280# diff_1238760_2043880# diff_1494800_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1133 diff_1519960_2051280# diff_1238760_2043880# diff_1519960_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1134 diff_1545120_2051280# diff_1238760_2043880# diff_1545120_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1135 diff_1570280_2051280# diff_1238760_2043880# diff_1570280_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1136 diff_1595440_2051280# diff_1238760_2043880# diff_1595440_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1137 diff_1620600_2051280# diff_1238760_2043880# diff_1620600_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1138 diff_1645760_2051280# diff_1238760_2043880# diff_1645760_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1139 diff_1670920_2051280# diff_1238760_2043880# diff_1670920_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1140 diff_1696080_2051280# diff_1238760_2043880# diff_1696080_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1141 diff_1721240_2051280# diff_1238760_2043880# diff_1721240_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1142 diff_1746400_2051280# diff_1238760_2043880# diff_1746400_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1143 diff_1771560_2051280# diff_1238760_2043880# diff_1771560_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1144 diff_1796720_2051280# diff_1238760_2043880# diff_1796720_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1145 diff_1821880_2051280# diff_1238760_2043880# diff_1821880_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1146 diff_1847040_2051280# diff_1238760_2043880# diff_1847040_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1147 diff_1872200_2051280# diff_1238760_2043880# diff_1872200_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1148 diff_1897360_2051280# diff_1238760_2043880# diff_1897360_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1149 diff_1922520_2051280# diff_1238760_2043880# diff_1922520_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1150 diff_1947680_2051280# diff_1238760_2043880# diff_1947680_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1151 diff_1972840_2051280# diff_1238760_2043880# diff_1972840_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1152 diff_1998000_2051280# diff_1238760_2043880# diff_1998000_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1153 diff_2023160_2051280# diff_1238760_2043880# diff_2023160_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1154 diff_2048320_2051280# diff_1238760_2043880# diff_2048320_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1155 diff_2073480_2051280# diff_1238760_2043880# diff_2073480_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1156 diff_2098640_2051280# diff_1238760_2043880# diff_2098640_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1157 diff_2123800_2051280# diff_1238760_2043880# diff_2123800_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1158 diff_2148960_2051280# diff_1238760_2043880# diff_2148960_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1159 diff_2174120_2051280# diff_1238760_2043880# diff_2174120_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1160 diff_2199280_2051280# diff_1238760_2043880# diff_2199280_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1161 diff_2224440_2051280# diff_1238760_2043880# diff_2224440_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1162 diff_2249600_2051280# diff_1238760_2043880# diff_2249600_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1163 diff_2274760_2051280# diff_1238760_2043880# diff_2274760_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1164 diff_2299920_2051280# diff_1238760_2043880# diff_2299920_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1165 diff_2325080_2051280# diff_1238760_2043880# diff_2325080_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1166 diff_2350240_2051280# diff_1238760_2043880# diff_2350240_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1167 diff_2375400_2051280# diff_1238760_2043880# diff_2375400_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1168 diff_2400560_2051280# diff_1238760_2043880# diff_2400560_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1169 diff_2425720_2051280# diff_1238760_2043880# diff_2425720_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1170 diff_2450880_2051280# diff_1238760_2043880# diff_2450880_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1171 diff_2476040_2051280# diff_1238760_2043880# diff_2476040_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1172 diff_2501200_2051280# diff_1238760_2043880# diff_2501200_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1173 diff_2526360_2051280# diff_1238760_2043880# diff_2526360_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1174 diff_2551520_2051280# diff_1238760_2043880# diff_2551520_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1175 diff_2576680_2051280# diff_1238760_2043880# diff_2576680_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1176 diff_2601840_2051280# diff_1238760_2043880# diff_2601840_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1177 diff_2627000_2051280# diff_1238760_2043880# diff_2627000_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1178 diff_2652160_2051280# diff_1238760_2043880# diff_2652160_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1179 diff_2677320_2051280# diff_1238760_2043880# diff_2677320_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1180 diff_2702480_2051280# diff_1238760_2043880# diff_2702480_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1181 diff_2727640_2051280# diff_1238760_2043880# diff_2727640_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1182 diff_2752800_2051280# diff_1238760_2043880# diff_2752800_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1183 diff_2777960_2051280# diff_1238760_2043880# diff_2777960_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1184 diff_2803120_2051280# diff_1238760_2043880# diff_2803120_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1185 diff_2828280_2051280# diff_1238760_2043880# diff_2828280_2024640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1186 diff_1238760_2072000# Vdd Vdd GND efet w=7400 l=14800
+ ad=0 pd=0 as=0 ps=0 
M1187 diff_1243200_2024640# diff_1238760_2017240# diff_1243200_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1188 diff_1268360_2024640# diff_1238760_2017240# diff_1268360_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1189 diff_1293520_2024640# diff_1238760_2017240# diff_1293520_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1190 diff_1318680_2024640# diff_1238760_2017240# diff_1318680_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1191 diff_1343840_2024640# diff_1238760_2017240# diff_1343840_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1192 diff_1369000_2024640# diff_1238760_2017240# diff_1369000_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1193 diff_1394160_2024640# diff_1238760_2017240# diff_1394160_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1194 diff_1419320_2024640# diff_1238760_2017240# diff_1419320_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1195 diff_1444480_2024640# diff_1238760_2017240# diff_1444480_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1196 diff_1469640_2024640# diff_1238760_2017240# diff_1469640_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1197 diff_1494800_2024640# diff_1238760_2017240# diff_1494800_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1198 diff_1519960_2024640# diff_1238760_2017240# diff_1519960_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1199 diff_1545120_2024640# diff_1238760_2017240# diff_1545120_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1200 diff_1570280_2024640# diff_1238760_2017240# diff_1570280_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1201 diff_1595440_2024640# diff_1238760_2017240# diff_1595440_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1202 diff_1620600_2024640# diff_1238760_2017240# diff_1620600_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1203 diff_1645760_2024640# diff_1238760_2017240# diff_1645760_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1204 diff_1670920_2024640# diff_1238760_2017240# diff_1670920_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1205 diff_1696080_2024640# diff_1238760_2017240# diff_1696080_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1206 diff_1721240_2024640# diff_1238760_2017240# diff_1721240_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1207 diff_1746400_2024640# diff_1238760_2017240# diff_1746400_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1208 diff_1771560_2024640# diff_1238760_2017240# diff_1771560_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1209 diff_1796720_2024640# diff_1238760_2017240# diff_1796720_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1210 diff_1821880_2024640# diff_1238760_2017240# diff_1821880_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1211 diff_1847040_2024640# diff_1238760_2017240# diff_1847040_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1212 diff_1872200_2024640# diff_1238760_2017240# diff_1872200_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1213 diff_1897360_2024640# diff_1238760_2017240# diff_1897360_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1214 diff_1922520_2024640# diff_1238760_2017240# diff_1922520_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1215 diff_1947680_2024640# diff_1238760_2017240# diff_1947680_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1216 diff_1972840_2024640# diff_1238760_2017240# diff_1972840_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1217 diff_1998000_2024640# diff_1238760_2017240# diff_1998000_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1218 diff_2023160_2024640# diff_1238760_2017240# diff_2023160_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1219 diff_2048320_2024640# diff_1238760_2017240# diff_2048320_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1220 diff_2073480_2024640# diff_1238760_2017240# diff_2073480_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1221 diff_2098640_2024640# diff_1238760_2017240# diff_2098640_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1222 diff_2123800_2024640# diff_1238760_2017240# diff_2123800_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1223 diff_2148960_2024640# diff_1238760_2017240# diff_2148960_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1224 diff_2174120_2024640# diff_1238760_2017240# diff_2174120_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1225 diff_2199280_2024640# diff_1238760_2017240# diff_2199280_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1226 diff_2224440_2024640# diff_1238760_2017240# diff_2224440_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1227 diff_2249600_2024640# diff_1238760_2017240# diff_2249600_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1228 diff_2274760_2024640# diff_1238760_2017240# diff_2274760_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1229 diff_2299920_2024640# diff_1238760_2017240# diff_2299920_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1230 diff_2325080_2024640# diff_1238760_2017240# diff_2325080_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1231 diff_2350240_2024640# diff_1238760_2017240# diff_2350240_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1232 diff_2375400_2024640# diff_1238760_2017240# diff_2375400_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1233 diff_2400560_2024640# diff_1238760_2017240# diff_2400560_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1234 diff_2425720_2024640# diff_1238760_2017240# diff_2425720_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1235 diff_2450880_2024640# diff_1238760_2017240# diff_2450880_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1236 diff_2476040_2024640# diff_1238760_2017240# diff_2476040_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1237 diff_2501200_2024640# diff_1238760_2017240# diff_2501200_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1238 diff_2526360_2024640# diff_1238760_2017240# diff_2526360_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1239 diff_2551520_2024640# diff_1238760_2017240# diff_2551520_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1240 diff_2576680_2024640# diff_1238760_2017240# diff_2576680_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1241 diff_2601840_2024640# diff_1238760_2017240# diff_2601840_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1242 diff_2627000_2024640# diff_1238760_2017240# diff_2627000_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1243 diff_2652160_2024640# diff_1238760_2017240# diff_2652160_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1244 diff_2677320_2024640# diff_1238760_2017240# diff_2677320_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1245 diff_2702480_2024640# diff_1238760_2017240# diff_2702480_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1246 diff_2727640_2024640# diff_1238760_2017240# diff_2727640_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1247 diff_2752800_2024640# diff_1238760_2017240# diff_2752800_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1248 diff_2777960_2024640# diff_1238760_2017240# diff_2777960_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1249 diff_2803120_2024640# diff_1238760_2017240# diff_2803120_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1250 diff_2828280_2024640# diff_1238760_2017240# diff_2828280_1996520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1251 Vdd Vdd diff_1238760_1989120# GND efet w=7400 l=14800
+ ad=0 pd=0 as=1.29453e+09 ps=319680 
M1252 diff_1243200_1996520# diff_1238760_1989120# diff_1243200_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1253 diff_1268360_1996520# diff_1238760_1989120# diff_1268360_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1254 diff_1293520_1996520# diff_1238760_1989120# diff_1293520_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1255 diff_1318680_1996520# diff_1238760_1989120# diff_1318680_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1256 diff_1343840_1996520# diff_1238760_1989120# diff_1343840_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1257 diff_1369000_1996520# diff_1238760_1989120# diff_1369000_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1258 diff_1394160_1996520# diff_1238760_1989120# diff_1394160_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1259 diff_1419320_1996520# diff_1238760_1989120# diff_1419320_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1260 diff_1444480_1996520# diff_1238760_1989120# diff_1444480_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1261 diff_1469640_1996520# diff_1238760_1989120# diff_1469640_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1262 diff_1494800_1996520# diff_1238760_1989120# diff_1494800_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1263 diff_1519960_1996520# diff_1238760_1989120# diff_1519960_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1264 diff_1545120_1996520# diff_1238760_1989120# diff_1545120_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1265 diff_1570280_1996520# diff_1238760_1989120# diff_1570280_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1266 diff_1595440_1996520# diff_1238760_1989120# diff_1595440_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1267 diff_1620600_1996520# diff_1238760_1989120# diff_1620600_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1268 diff_1645760_1996520# diff_1238760_1989120# diff_1645760_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1269 diff_1670920_1996520# diff_1238760_1989120# diff_1670920_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1270 diff_1696080_1996520# diff_1238760_1989120# diff_1696080_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1271 diff_1721240_1996520# diff_1238760_1989120# diff_1721240_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1272 diff_1746400_1996520# diff_1238760_1989120# diff_1746400_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1273 diff_1771560_1996520# diff_1238760_1989120# diff_1771560_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1274 diff_1796720_1996520# diff_1238760_1989120# diff_1796720_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1275 diff_1821880_1996520# diff_1238760_1989120# diff_1821880_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1276 diff_1847040_1996520# diff_1238760_1989120# diff_1847040_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1277 diff_1872200_1996520# diff_1238760_1989120# diff_1872200_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1278 diff_1897360_1996520# diff_1238760_1989120# diff_1897360_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1279 diff_1922520_1996520# diff_1238760_1989120# diff_1922520_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1280 diff_1947680_1996520# diff_1238760_1989120# diff_1947680_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1281 diff_1972840_1996520# diff_1238760_1989120# diff_1972840_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1282 diff_1998000_1996520# diff_1238760_1989120# diff_1998000_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1283 diff_2023160_1996520# diff_1238760_1989120# diff_2023160_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1284 diff_2048320_1996520# diff_1238760_1989120# diff_2048320_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1285 diff_2073480_1996520# diff_1238760_1989120# diff_2073480_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1286 diff_2098640_1996520# diff_1238760_1989120# diff_2098640_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1287 diff_2123800_1996520# diff_1238760_1989120# diff_2123800_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1288 diff_2148960_1996520# diff_1238760_1989120# diff_2148960_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1289 diff_2174120_1996520# diff_1238760_1989120# diff_2174120_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1290 diff_2199280_1996520# diff_1238760_1989120# diff_2199280_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1291 diff_2224440_1996520# diff_1238760_1989120# diff_2224440_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1292 diff_2249600_1996520# diff_1238760_1989120# diff_2249600_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1293 diff_2274760_1996520# diff_1238760_1989120# diff_2274760_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1294 diff_2299920_1996520# diff_1238760_1989120# diff_2299920_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1295 diff_2325080_1996520# diff_1238760_1989120# diff_2325080_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1296 diff_2350240_1996520# diff_1238760_1989120# diff_2350240_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1297 diff_2375400_1996520# diff_1238760_1989120# diff_2375400_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1298 diff_2400560_1996520# diff_1238760_1989120# diff_2400560_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1299 diff_2425720_1996520# diff_1238760_1989120# diff_2425720_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1300 diff_2450880_1996520# diff_1238760_1989120# diff_2450880_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1301 diff_2476040_1996520# diff_1238760_1989120# diff_2476040_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1302 diff_2501200_1996520# diff_1238760_1989120# diff_2501200_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1303 diff_2526360_1996520# diff_1238760_1989120# diff_2526360_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1304 diff_2551520_1996520# diff_1238760_1989120# diff_2551520_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1305 diff_2576680_1996520# diff_1238760_1989120# diff_2576680_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1306 diff_2601840_1996520# diff_1238760_1989120# diff_2601840_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1307 diff_2627000_1996520# diff_1238760_1989120# diff_2627000_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1308 diff_2652160_1996520# diff_1238760_1989120# diff_2652160_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1309 diff_2677320_1996520# diff_1238760_1989120# diff_2677320_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1310 diff_2702480_1996520# diff_1238760_1989120# diff_2702480_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1311 diff_2727640_1996520# diff_1238760_1989120# diff_2727640_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1312 diff_2752800_1996520# diff_1238760_1989120# diff_2752800_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1313 diff_2777960_1996520# diff_1238760_1989120# diff_2777960_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1314 diff_2803120_1996520# diff_1238760_1989120# diff_2803120_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1315 diff_2828280_1996520# diff_1238760_1989120# diff_2828280_1969880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1316 diff_1238760_1989120# diff_2940760_526880# diff_2920040_2064600# GND efet w=91760 l=7400
+ ad=0 pd=0 as=0 ps=0 
M1317 diff_2920040_2064600# diff_2976280_1228400# diff_1238760_2043880# GND efet w=102120 l=8880
+ ad=0 pd=0 as=1.6428e+09 ps=275280 
M1318 diff_1238760_2043880# Vdd Vdd GND efet w=8880 l=14800
+ ad=0 pd=0 as=0 ps=0 
M1319 Vdd Vdd diff_1238760_2017240# GND efet w=8880 l=14800
+ ad=0 pd=0 as=1.43252e+09 ps=304880 
M1320 diff_1243200_1969880# diff_1238760_1962480# diff_1243200_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1321 diff_1268360_1969880# diff_1238760_1962480# diff_1268360_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1322 diff_1293520_1969880# diff_1238760_1962480# diff_1293520_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1323 diff_1318680_1969880# diff_1238760_1962480# diff_1318680_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1324 diff_1343840_1969880# diff_1238760_1962480# diff_1343840_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1325 diff_1369000_1969880# diff_1238760_1962480# diff_1369000_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1326 diff_1394160_1969880# diff_1238760_1962480# diff_1394160_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1327 diff_1419320_1969880# diff_1238760_1962480# diff_1419320_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1328 diff_1444480_1969880# diff_1238760_1962480# diff_1444480_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1329 diff_1469640_1969880# diff_1238760_1962480# diff_1469640_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1330 diff_1494800_1969880# diff_1238760_1962480# diff_1494800_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1331 diff_1519960_1969880# diff_1238760_1962480# diff_1519960_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1332 diff_1545120_1969880# diff_1238760_1962480# diff_1545120_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1333 diff_1570280_1969880# diff_1238760_1962480# diff_1570280_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1334 diff_1595440_1969880# diff_1238760_1962480# diff_1595440_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1335 diff_1620600_1969880# diff_1238760_1962480# diff_1620600_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1336 diff_1645760_1969880# diff_1238760_1962480# diff_1645760_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1337 diff_1670920_1969880# diff_1238760_1962480# diff_1670920_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1338 diff_1696080_1969880# diff_1238760_1962480# diff_1696080_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1339 diff_1721240_1969880# diff_1238760_1962480# diff_1721240_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1340 diff_1746400_1969880# diff_1238760_1962480# diff_1746400_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1341 diff_1771560_1969880# diff_1238760_1962480# diff_1771560_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1342 diff_1796720_1969880# diff_1238760_1962480# diff_1796720_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1343 diff_1821880_1969880# diff_1238760_1962480# diff_1821880_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1344 diff_1847040_1969880# diff_1238760_1962480# diff_1847040_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1345 diff_1872200_1969880# diff_1238760_1962480# diff_1872200_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1346 diff_1897360_1969880# diff_1238760_1962480# diff_1897360_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1347 diff_1922520_1969880# diff_1238760_1962480# diff_1922520_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1348 diff_1947680_1969880# diff_1238760_1962480# diff_1947680_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1349 diff_1972840_1969880# diff_1238760_1962480# diff_1972840_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1350 diff_1998000_1969880# diff_1238760_1962480# diff_1998000_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1351 diff_2023160_1969880# diff_1238760_1962480# diff_2023160_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1352 diff_2048320_1969880# diff_1238760_1962480# diff_2048320_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1353 diff_2073480_1969880# diff_1238760_1962480# diff_2073480_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1354 diff_2098640_1969880# diff_1238760_1962480# diff_2098640_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1355 diff_2123800_1969880# diff_1238760_1962480# diff_2123800_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1356 diff_2148960_1969880# diff_1238760_1962480# diff_2148960_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1357 diff_2174120_1969880# diff_1238760_1962480# diff_2174120_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1358 diff_2199280_1969880# diff_1238760_1962480# diff_2199280_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1359 diff_2224440_1969880# diff_1238760_1962480# diff_2224440_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1360 diff_2249600_1969880# diff_1238760_1962480# diff_2249600_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1361 diff_2274760_1969880# diff_1238760_1962480# diff_2274760_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1362 diff_2299920_1969880# diff_1238760_1962480# diff_2299920_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1363 diff_2325080_1969880# diff_1238760_1962480# diff_2325080_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1364 diff_2350240_1969880# diff_1238760_1962480# diff_2350240_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1365 diff_2375400_1969880# diff_1238760_1962480# diff_2375400_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1366 diff_2400560_1969880# diff_1238760_1962480# diff_2400560_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1367 diff_2425720_1969880# diff_1238760_1962480# diff_2425720_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1368 diff_2450880_1969880# diff_1238760_1962480# diff_2450880_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1369 diff_2476040_1969880# diff_1238760_1962480# diff_2476040_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1370 diff_2501200_1969880# diff_1238760_1962480# diff_2501200_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1371 diff_2526360_1969880# diff_1238760_1962480# diff_2526360_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1372 diff_2551520_1969880# diff_1238760_1962480# diff_2551520_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1373 diff_2576680_1969880# diff_1238760_1962480# diff_2576680_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1374 diff_2601840_1969880# diff_1238760_1962480# diff_2601840_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1375 diff_2627000_1969880# diff_1238760_1962480# diff_2627000_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1376 diff_2652160_1969880# diff_1238760_1962480# diff_2652160_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1377 diff_2677320_1969880# diff_1238760_1962480# diff_2677320_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1378 diff_2702480_1969880# diff_1238760_1962480# diff_2702480_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1379 diff_2727640_1969880# diff_1238760_1962480# diff_2727640_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1380 diff_2752800_1969880# diff_1238760_1962480# diff_2752800_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1381 diff_2777960_1969880# diff_1238760_1962480# diff_2777960_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1382 diff_2803120_1969880# diff_1238760_1962480# diff_2803120_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1383 diff_2828280_1969880# diff_1238760_1962480# diff_2828280_1941760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1384 diff_2920040_1955080# diff_2912640_526880# diff_1238760_1962480# GND efet w=108040 l=8140
+ ad=1.52054e+09 pd=902800 as=1.35367e+09 ps=278240 
M1385 diff_1238760_2017240# diff_2998480_1207680# diff_2920040_2064600# GND efet w=97680 l=7400
+ ad=0 pd=0 as=0 ps=0 
M1386 diff_1243200_1941760# diff_1238760_1934360# diff_1243200_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1387 diff_1268360_1941760# diff_1238760_1934360# diff_1268360_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1388 diff_1293520_1941760# diff_1238760_1934360# diff_1293520_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1389 diff_1318680_1941760# diff_1238760_1934360# diff_1318680_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1390 diff_1343840_1941760# diff_1238760_1934360# diff_1343840_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1391 diff_1369000_1941760# diff_1238760_1934360# diff_1369000_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1392 diff_1394160_1941760# diff_1238760_1934360# diff_1394160_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1393 diff_1419320_1941760# diff_1238760_1934360# diff_1419320_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1394 diff_1444480_1941760# diff_1238760_1934360# diff_1444480_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1395 diff_1469640_1941760# diff_1238760_1934360# diff_1469640_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1396 diff_1494800_1941760# diff_1238760_1934360# diff_1494800_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1397 diff_1519960_1941760# diff_1238760_1934360# diff_1519960_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1398 diff_1545120_1941760# diff_1238760_1934360# diff_1545120_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1399 diff_1570280_1941760# diff_1238760_1934360# diff_1570280_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1400 diff_1595440_1941760# diff_1238760_1934360# diff_1595440_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1401 diff_1620600_1941760# diff_1238760_1934360# diff_1620600_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1402 diff_1645760_1941760# diff_1238760_1934360# diff_1645760_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1403 diff_1670920_1941760# diff_1238760_1934360# diff_1670920_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1404 diff_1696080_1941760# diff_1238760_1934360# diff_1696080_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1405 diff_1721240_1941760# diff_1238760_1934360# diff_1721240_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1406 diff_1746400_1941760# diff_1238760_1934360# diff_1746400_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1407 diff_1771560_1941760# diff_1238760_1934360# diff_1771560_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1408 diff_1796720_1941760# diff_1238760_1934360# diff_1796720_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1409 diff_1821880_1941760# diff_1238760_1934360# diff_1821880_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1410 diff_1847040_1941760# diff_1238760_1934360# diff_1847040_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1411 diff_1872200_1941760# diff_1238760_1934360# diff_1872200_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1412 diff_1897360_1941760# diff_1238760_1934360# diff_1897360_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1413 diff_1922520_1941760# diff_1238760_1934360# diff_1922520_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1414 diff_1947680_1941760# diff_1238760_1934360# diff_1947680_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1415 diff_1972840_1941760# diff_1238760_1934360# diff_1972840_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1416 diff_1998000_1941760# diff_1238760_1934360# diff_1998000_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1417 diff_2023160_1941760# diff_1238760_1934360# diff_2023160_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1418 diff_2048320_1941760# diff_1238760_1934360# diff_2048320_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1419 diff_2073480_1941760# diff_1238760_1934360# diff_2073480_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1420 diff_2098640_1941760# diff_1238760_1934360# diff_2098640_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1421 diff_2123800_1941760# diff_1238760_1934360# diff_2123800_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1422 diff_2148960_1941760# diff_1238760_1934360# diff_2148960_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1423 diff_2174120_1941760# diff_1238760_1934360# diff_2174120_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1424 diff_2199280_1941760# diff_1238760_1934360# diff_2199280_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1425 diff_2224440_1941760# diff_1238760_1934360# diff_2224440_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1426 diff_2249600_1941760# diff_1238760_1934360# diff_2249600_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1427 diff_2274760_1941760# diff_1238760_1934360# diff_2274760_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1428 diff_2299920_1941760# diff_1238760_1934360# diff_2299920_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1429 diff_2325080_1941760# diff_1238760_1934360# diff_2325080_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1430 diff_2350240_1941760# diff_1238760_1934360# diff_2350240_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1431 diff_2375400_1941760# diff_1238760_1934360# diff_2375400_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1432 diff_2400560_1941760# diff_1238760_1934360# diff_2400560_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1433 diff_2425720_1941760# diff_1238760_1934360# diff_2425720_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1434 diff_2450880_1941760# diff_1238760_1934360# diff_2450880_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1435 diff_2476040_1941760# diff_1238760_1934360# diff_2476040_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1436 diff_2501200_1941760# diff_1238760_1934360# diff_2501200_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1437 diff_2526360_1941760# diff_1238760_1934360# diff_2526360_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1438 diff_2551520_1941760# diff_1238760_1934360# diff_2551520_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1439 diff_2576680_1941760# diff_1238760_1934360# diff_2576680_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1440 diff_2601840_1941760# diff_1238760_1934360# diff_2601840_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1441 diff_2627000_1941760# diff_1238760_1934360# diff_2627000_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1442 diff_2652160_1941760# diff_1238760_1934360# diff_2652160_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1443 diff_2677320_1941760# diff_1238760_1934360# diff_2677320_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1444 diff_2702480_1941760# diff_1238760_1934360# diff_2702480_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1445 diff_2727640_1941760# diff_1238760_1934360# diff_2727640_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1446 diff_2752800_1941760# diff_1238760_1934360# diff_2752800_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1447 diff_2777960_1941760# diff_1238760_1934360# diff_2777960_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1448 diff_2803120_1941760# diff_1238760_1934360# diff_2803120_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1449 diff_2828280_1941760# diff_1238760_1934360# diff_2828280_1915120# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1450 diff_1025640_1855920# diff_1025640_1855920# diff_1025640_1855920# GND efet w=740 l=2220
+ ad=0 pd=0 as=0 ps=0 
M1451 diff_438080_1685720# diff_417360_2049800# GND GND efet w=119880 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1452 diff_417360_2049800# diff_503200_1786360# GND GND efet w=230880 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1453 diff_819920_1684240# diff_830280_1857400# diff_819920_1684240# GND efet w=75480 l=4440
+ ad=0 pd=0 as=0 ps=0 
M1454 diff_800680_2049800# diff_910200_1857400# diff_800680_2049800# GND efet w=70300 l=9620
+ ad=0 pd=0 as=0 ps=0 
M1455 GND diff_233840_991600# diff_438080_1685720# GND efet w=233840 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1456 diff_629000_1685720# diff_609760_2049800# GND GND efet w=119880 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1457 diff_609760_2049800# diff_694120_1786360# GND GND efet w=232360 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1458 diff_1012320_1684240# diff_1025640_1855920# diff_1012320_1684240# GND efet w=52540 l=17020
+ ad=0 pd=0 as=0 ps=0 
M1459 diff_1093720_1907720# diff_1093720_1907720# diff_1093720_1907720# GND efet w=740 l=2220
+ ad=0 pd=0 as=0 ps=0 
M1460 diff_1238760_1962480# Vdd Vdd GND efet w=7400 l=16280
+ ad=0 pd=0 as=0 ps=0 
M1461 diff_1243200_1915120# diff_1238760_1907720# diff_1243200_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1462 diff_1268360_1915120# diff_1238760_1907720# diff_1268360_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1463 diff_1293520_1915120# diff_1238760_1907720# diff_1293520_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1464 diff_1318680_1915120# diff_1238760_1907720# diff_1318680_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1465 diff_1343840_1915120# diff_1238760_1907720# diff_1343840_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1466 diff_1369000_1915120# diff_1238760_1907720# diff_1369000_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1467 diff_1394160_1915120# diff_1238760_1907720# diff_1394160_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1468 diff_1419320_1915120# diff_1238760_1907720# diff_1419320_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1469 diff_1444480_1915120# diff_1238760_1907720# diff_1444480_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1470 diff_1469640_1915120# diff_1238760_1907720# diff_1469640_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1471 diff_1494800_1915120# diff_1238760_1907720# diff_1494800_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1472 diff_1519960_1915120# diff_1238760_1907720# diff_1519960_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1473 diff_1545120_1915120# diff_1238760_1907720# diff_1545120_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1474 diff_1570280_1915120# diff_1238760_1907720# diff_1570280_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1475 diff_1595440_1915120# diff_1238760_1907720# diff_1595440_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1476 diff_1620600_1915120# diff_1238760_1907720# diff_1620600_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1477 diff_1645760_1915120# diff_1238760_1907720# diff_1645760_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1478 diff_1670920_1915120# diff_1238760_1907720# diff_1670920_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1479 diff_1696080_1915120# diff_1238760_1907720# diff_1696080_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1480 diff_1721240_1915120# diff_1238760_1907720# diff_1721240_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1481 diff_1746400_1915120# diff_1238760_1907720# diff_1746400_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1482 diff_1771560_1915120# diff_1238760_1907720# diff_1771560_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1483 diff_1796720_1915120# diff_1238760_1907720# diff_1796720_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1484 diff_1821880_1915120# diff_1238760_1907720# diff_1821880_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1485 diff_1847040_1915120# diff_1238760_1907720# diff_1847040_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1486 diff_1872200_1915120# diff_1238760_1907720# diff_1872200_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1487 diff_1897360_1915120# diff_1238760_1907720# diff_1897360_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1488 diff_1922520_1915120# diff_1238760_1907720# diff_1922520_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1489 diff_1947680_1915120# diff_1238760_1907720# diff_1947680_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1490 diff_1972840_1915120# diff_1238760_1907720# diff_1972840_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1491 diff_1998000_1915120# diff_1238760_1907720# diff_1998000_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1492 diff_2023160_1915120# diff_1238760_1907720# diff_2023160_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1493 diff_2048320_1915120# diff_1238760_1907720# diff_2048320_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1494 diff_2073480_1915120# diff_1238760_1907720# diff_2073480_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1495 diff_2098640_1915120# diff_1238760_1907720# diff_2098640_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1496 diff_2123800_1915120# diff_1238760_1907720# diff_2123800_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1497 diff_2148960_1915120# diff_1238760_1907720# diff_2148960_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1498 diff_2174120_1915120# diff_1238760_1907720# diff_2174120_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1499 diff_2199280_1915120# diff_1238760_1907720# diff_2199280_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1500 diff_2224440_1915120# diff_1238760_1907720# diff_2224440_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1501 diff_2249600_1915120# diff_1238760_1907720# diff_2249600_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1502 diff_2274760_1915120# diff_1238760_1907720# diff_2274760_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1503 diff_2299920_1915120# diff_1238760_1907720# diff_2299920_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1504 diff_2325080_1915120# diff_1238760_1907720# diff_2325080_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1505 diff_2350240_1915120# diff_1238760_1907720# diff_2350240_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1506 diff_2375400_1915120# diff_1238760_1907720# diff_2375400_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1507 diff_2400560_1915120# diff_1238760_1907720# diff_2400560_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1508 diff_2425720_1915120# diff_1238760_1907720# diff_2425720_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1509 diff_2450880_1915120# diff_1238760_1907720# diff_2450880_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1510 diff_2476040_1915120# diff_1238760_1907720# diff_2476040_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1511 diff_2501200_1915120# diff_1238760_1907720# diff_2501200_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1512 diff_2526360_1915120# diff_1238760_1907720# diff_2526360_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1513 diff_2551520_1915120# diff_1238760_1907720# diff_2551520_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1514 diff_2576680_1915120# diff_1238760_1907720# diff_2576680_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1515 diff_2601840_1915120# diff_1238760_1907720# diff_2601840_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1516 diff_2627000_1915120# diff_1238760_1907720# diff_2627000_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1517 diff_2652160_1915120# diff_1238760_1907720# diff_2652160_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1518 diff_2677320_1915120# diff_1238760_1907720# diff_2677320_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1519 diff_2702480_1915120# diff_1238760_1907720# diff_2702480_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1520 diff_2727640_1915120# diff_1238760_1907720# diff_2727640_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1521 diff_2752800_1915120# diff_1238760_1907720# diff_2752800_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1522 diff_2777960_1915120# diff_1238760_1907720# diff_2777960_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1523 diff_2803120_1915120# diff_1238760_1907720# diff_2803120_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1524 diff_2828280_1915120# diff_1238760_1907720# diff_2828280_1887000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1525 diff_991600_2049800# diff_1093720_1907720# diff_991600_2049800# GND efet w=62160 l=12580
+ ad=0 pd=0 as=0 ps=0 
M1526 Vdd Vdd diff_1238760_1879600# GND efet w=7400 l=16280
+ ad=0 pd=0 as=1.29453e+09 ps=319680 
M1527 diff_1243200_1887000# diff_1238760_1879600# diff_1243200_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1528 diff_1268360_1887000# diff_1238760_1879600# diff_1268360_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1529 diff_1293520_1887000# diff_1238760_1879600# diff_1293520_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1530 diff_1318680_1887000# diff_1238760_1879600# diff_1318680_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1531 diff_1343840_1887000# diff_1238760_1879600# diff_1343840_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1532 diff_1369000_1887000# diff_1238760_1879600# diff_1369000_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1533 diff_1394160_1887000# diff_1238760_1879600# diff_1394160_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1534 diff_1419320_1887000# diff_1238760_1879600# diff_1419320_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1535 diff_1444480_1887000# diff_1238760_1879600# diff_1444480_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1536 diff_1469640_1887000# diff_1238760_1879600# diff_1469640_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1537 diff_1494800_1887000# diff_1238760_1879600# diff_1494800_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1538 diff_1519960_1887000# diff_1238760_1879600# diff_1519960_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1539 diff_1545120_1887000# diff_1238760_1879600# diff_1545120_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1540 diff_1570280_1887000# diff_1238760_1879600# diff_1570280_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1541 diff_1595440_1887000# diff_1238760_1879600# diff_1595440_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1542 diff_1620600_1887000# diff_1238760_1879600# diff_1620600_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1543 diff_1645760_1887000# diff_1238760_1879600# diff_1645760_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1544 diff_1670920_1887000# diff_1238760_1879600# diff_1670920_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1545 diff_1696080_1887000# diff_1238760_1879600# diff_1696080_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1546 diff_1721240_1887000# diff_1238760_1879600# diff_1721240_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1547 diff_1746400_1887000# diff_1238760_1879600# diff_1746400_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1548 diff_1771560_1887000# diff_1238760_1879600# diff_1771560_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1549 diff_1796720_1887000# diff_1238760_1879600# diff_1796720_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1550 diff_1821880_1887000# diff_1238760_1879600# diff_1821880_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1551 diff_1847040_1887000# diff_1238760_1879600# diff_1847040_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1552 diff_1872200_1887000# diff_1238760_1879600# diff_1872200_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1553 diff_1897360_1887000# diff_1238760_1879600# diff_1897360_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1554 diff_1922520_1887000# diff_1238760_1879600# diff_1922520_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1555 diff_1947680_1887000# diff_1238760_1879600# diff_1947680_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1556 diff_1972840_1887000# diff_1238760_1879600# diff_1972840_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1557 diff_1998000_1887000# diff_1238760_1879600# diff_1998000_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1558 diff_2023160_1887000# diff_1238760_1879600# diff_2023160_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1559 diff_2048320_1887000# diff_1238760_1879600# diff_2048320_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1560 diff_2073480_1887000# diff_1238760_1879600# diff_2073480_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1561 diff_2098640_1887000# diff_1238760_1879600# diff_2098640_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1562 diff_2123800_1887000# diff_1238760_1879600# diff_2123800_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1563 diff_2148960_1887000# diff_1238760_1879600# diff_2148960_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1564 diff_2174120_1887000# diff_1238760_1879600# diff_2174120_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1565 diff_2199280_1887000# diff_1238760_1879600# diff_2199280_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1566 diff_2224440_1887000# diff_1238760_1879600# diff_2224440_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1567 diff_2249600_1887000# diff_1238760_1879600# diff_2249600_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1568 diff_2274760_1887000# diff_1238760_1879600# diff_2274760_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1569 diff_2299920_1887000# diff_1238760_1879600# diff_2299920_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1570 diff_2325080_1887000# diff_1238760_1879600# diff_2325080_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1571 diff_2350240_1887000# diff_1238760_1879600# diff_2350240_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1572 diff_2375400_1887000# diff_1238760_1879600# diff_2375400_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1573 diff_2400560_1887000# diff_1238760_1879600# diff_2400560_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1574 diff_2425720_1887000# diff_1238760_1879600# diff_2425720_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1575 diff_2450880_1887000# diff_1238760_1879600# diff_2450880_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1576 diff_2476040_1887000# diff_1238760_1879600# diff_2476040_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1577 diff_2501200_1887000# diff_1238760_1879600# diff_2501200_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1578 diff_2526360_1887000# diff_1238760_1879600# diff_2526360_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1579 diff_2551520_1887000# diff_1238760_1879600# diff_2551520_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1580 diff_2576680_1887000# diff_1238760_1879600# diff_2576680_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1581 diff_2601840_1887000# diff_1238760_1879600# diff_2601840_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1582 diff_2627000_1887000# diff_1238760_1879600# diff_2627000_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1583 diff_2652160_1887000# diff_1238760_1879600# diff_2652160_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1584 diff_2677320_1887000# diff_1238760_1879600# diff_2677320_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1585 diff_2702480_1887000# diff_1238760_1879600# diff_2702480_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1586 diff_2727640_1887000# diff_1238760_1879600# diff_2727640_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1587 diff_2752800_1887000# diff_1238760_1879600# diff_2752800_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1588 diff_2777960_1887000# diff_1238760_1879600# diff_2777960_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1589 diff_2803120_1887000# diff_1238760_1879600# diff_2803120_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1590 diff_2828280_1887000# diff_1238760_1879600# diff_2828280_1860360# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1591 diff_1238760_1879600# diff_2940760_526880# diff_2920040_1955080# GND efet w=91760 l=7400
+ ad=0 pd=0 as=0 ps=0 
M1592 diff_2920040_1955080# diff_2976280_1228400# diff_1238760_1934360# GND efet w=104340 l=8140
+ ad=0 pd=0 as=1.70851e+09 ps=275280 
M1593 diff_1238760_1934360# Vdd Vdd GND efet w=8880 l=17760
+ ad=0 pd=0 as=0 ps=0 
M1594 Vdd Vdd diff_1238760_1907720# GND efet w=8880 l=16280
+ ad=0 pd=0 as=1.43252e+09 ps=304880 
M1595 diff_1243200_1860360# diff_1238760_1852960# diff_1243200_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1596 diff_1268360_1860360# diff_1238760_1852960# diff_1268360_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1597 diff_1293520_1860360# diff_1238760_1852960# diff_1293520_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1598 diff_1318680_1860360# diff_1238760_1852960# diff_1318680_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1599 diff_1343840_1860360# diff_1238760_1852960# diff_1343840_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1600 diff_1369000_1860360# diff_1238760_1852960# diff_1369000_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1601 diff_1394160_1860360# diff_1238760_1852960# diff_1394160_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1602 diff_1419320_1860360# diff_1238760_1852960# diff_1419320_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1603 diff_1444480_1860360# diff_1238760_1852960# diff_1444480_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1604 diff_1469640_1860360# diff_1238760_1852960# diff_1469640_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1605 diff_1494800_1860360# diff_1238760_1852960# diff_1494800_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1606 diff_1519960_1860360# diff_1238760_1852960# diff_1519960_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1607 diff_1545120_1860360# diff_1238760_1852960# diff_1545120_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1608 diff_1570280_1860360# diff_1238760_1852960# diff_1570280_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1609 diff_1595440_1860360# diff_1238760_1852960# diff_1595440_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1610 diff_1620600_1860360# diff_1238760_1852960# diff_1620600_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1611 diff_1645760_1860360# diff_1238760_1852960# diff_1645760_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1612 diff_1670920_1860360# diff_1238760_1852960# diff_1670920_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1613 diff_1696080_1860360# diff_1238760_1852960# diff_1696080_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1614 diff_1721240_1860360# diff_1238760_1852960# diff_1721240_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1615 diff_1746400_1860360# diff_1238760_1852960# diff_1746400_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1616 diff_1771560_1860360# diff_1238760_1852960# diff_1771560_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1617 diff_1796720_1860360# diff_1238760_1852960# diff_1796720_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1618 diff_1821880_1860360# diff_1238760_1852960# diff_1821880_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1619 diff_1847040_1860360# diff_1238760_1852960# diff_1847040_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1620 diff_1872200_1860360# diff_1238760_1852960# diff_1872200_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1621 diff_1897360_1860360# diff_1238760_1852960# diff_1897360_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1622 diff_1922520_1860360# diff_1238760_1852960# diff_1922520_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1623 diff_1947680_1860360# diff_1238760_1852960# diff_1947680_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1624 diff_1972840_1860360# diff_1238760_1852960# diff_1972840_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1625 diff_1998000_1860360# diff_1238760_1852960# diff_1998000_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1626 diff_2023160_1860360# diff_1238760_1852960# diff_2023160_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1627 diff_2048320_1860360# diff_1238760_1852960# diff_2048320_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1628 diff_2073480_1860360# diff_1238760_1852960# diff_2073480_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1629 diff_2098640_1860360# diff_1238760_1852960# diff_2098640_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1630 diff_2123800_1860360# diff_1238760_1852960# diff_2123800_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1631 diff_2148960_1860360# diff_1238760_1852960# diff_2148960_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1632 diff_2174120_1860360# diff_1238760_1852960# diff_2174120_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1633 diff_2199280_1860360# diff_1238760_1852960# diff_2199280_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1634 diff_2224440_1860360# diff_1238760_1852960# diff_2224440_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1635 diff_2249600_1860360# diff_1238760_1852960# diff_2249600_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1636 diff_2274760_1860360# diff_1238760_1852960# diff_2274760_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1637 diff_2299920_1860360# diff_1238760_1852960# diff_2299920_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1638 diff_2325080_1860360# diff_1238760_1852960# diff_2325080_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1639 diff_2350240_1860360# diff_1238760_1852960# diff_2350240_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1640 diff_2375400_1860360# diff_1238760_1852960# diff_2375400_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1641 diff_2400560_1860360# diff_1238760_1852960# diff_2400560_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1642 diff_2425720_1860360# diff_1238760_1852960# diff_2425720_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1643 diff_2450880_1860360# diff_1238760_1852960# diff_2450880_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1644 diff_2476040_1860360# diff_1238760_1852960# diff_2476040_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1645 diff_2501200_1860360# diff_1238760_1852960# diff_2501200_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1646 diff_2526360_1860360# diff_1238760_1852960# diff_2526360_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1647 diff_2551520_1860360# diff_1238760_1852960# diff_2551520_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1648 diff_2576680_1860360# diff_1238760_1852960# diff_2576680_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1649 diff_2601840_1860360# diff_1238760_1852960# diff_2601840_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1650 diff_2627000_1860360# diff_1238760_1852960# diff_2627000_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1651 diff_2652160_1860360# diff_1238760_1852960# diff_2652160_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1652 diff_2677320_1860360# diff_1238760_1852960# diff_2677320_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1653 diff_2702480_1860360# diff_1238760_1852960# diff_2702480_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1654 diff_2727640_1860360# diff_1238760_1852960# diff_2727640_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1655 diff_2752800_1860360# diff_1238760_1852960# diff_2752800_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1656 diff_2777960_1860360# diff_1238760_1852960# diff_2777960_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1657 diff_2803120_1860360# diff_1238760_1852960# diff_2803120_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1658 diff_2828280_1860360# diff_1238760_1852960# diff_2828280_1832240# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1659 diff_417360_2049800# diff_233840_991600# GND GND efet w=235320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1660 GND diff_233840_991600# diff_629000_1685720# GND efet w=233840 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1661 diff_819920_1684240# diff_800680_2049800# GND GND efet w=119880 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1662 diff_800680_2049800# diff_886520_1786360# GND GND efet w=232360 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1663 diff_609760_2049800# diff_233840_991600# GND GND efet w=235320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1664 GND diff_233840_991600# diff_819920_1684240# GND efet w=235320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1665 diff_1012320_1684240# diff_991600_2049800# GND GND efet w=119880 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1666 diff_991600_2049800# diff_1077440_1786360# GND GND efet w=232360 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1667 diff_2920040_1842600# diff_2912640_526880# diff_1238760_1852960# GND efet w=108780 l=8880
+ ad=1.57969e+09 pd=885040 as=1.43252e+09 ps=284160 
M1668 diff_1238760_1907720# diff_2998480_1207680# diff_2920040_1955080# GND efet w=97680 l=7400
+ ad=0 pd=0 as=0 ps=0 
M1669 diff_3005880_2094200# diff_3069520_1052280# diff_2920040_1955080# GND efet w=190920 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1670 diff_2920040_2064600# diff_3090240_1133680# diff_3005880_2094200# GND efet w=198320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1671 diff_3001440_2148960# Vdd Vdd GND efet w=8880 l=17760
+ ad=0 pd=0 as=0 ps=0 
M1672 diff_3393640_2079400# diff_3393640_2079400# diff_3393640_2079400# GND efet w=1480 l=2220
+ ad=1.30767e+09 pd=287120 as=0 ps=0 
M1673 diff_3383280_2114920# diff_3285600_1753800# diff_3383280_2100120# GND efet w=50320 l=7400
+ ad=0 pd=0 as=6.65882e+08 ps=148000 
M1674 diff_3393640_2079400# diff_3393640_2079400# diff_3393640_2079400# GND efet w=740 l=1480
+ ad=0 pd=0 as=0 ps=0 
M1675 GND diff_3307800_2085320# diff_3285600_2079400# GND efet w=28120 l=7400
+ ad=0 pd=0 as=1.13025e+09 ps=266400 
M1676 diff_3383280_2100120# diff_3267840_1873680# diff_3393640_2079400# GND efet w=51800 l=7400
+ ad=0 pd=0 as=0 ps=0 
M1677 diff_3285600_2079400# diff_3285600_2079400# diff_3285600_2079400# GND efet w=1480 l=1480
+ ad=0 pd=0 as=0 ps=0 
M1678 GND d3 diff_3488360_1339400# GND efet w=199800 l=7400
+ ad=0 pd=0 as=-1.51754e+09 ps=438080 
M1679 diff_3285600_2079400# Vdd Vdd GND efet w=8140 l=47360
+ ad=0 pd=0 as=0 ps=0 
M1680 diff_3307800_2085320# diff_3307800_2085320# diff_3307800_2085320# GND efet w=2220 l=5180
+ ad=2.1904e+08 pd=62160 as=0 ps=0 
M1681 Vdd Vdd Vdd GND efet w=740 l=1480
+ ad=0 pd=0 as=0 ps=0 
M1682 Vdd Vdd Vdd GND efet w=1480 l=2960
+ ad=0 pd=0 as=0 ps=0 
M1683 diff_3307800_2085320# diff_3307800_2085320# diff_3307800_2085320# GND efet w=1480 l=3700
+ ad=0 pd=0 as=0 ps=0 
M1684 Vdd Vdd diff_3393640_2079400# GND efet w=8880 l=39960
+ ad=0 pd=0 as=0 ps=0 
M1685 diff_3455800_2137120# Vdd Vdd GND efet w=7400 l=26640
+ ad=0 pd=0 as=0 ps=0 
M1686 diff_3267840_1761200# Vdd Vdd GND efet w=8880 l=14800
+ ad=0 pd=0 as=0 ps=0 
M1687 diff_3488360_1339400# Vdd Vdd GND efet w=11840 l=19240
+ ad=0 pd=0 as=0 ps=0 
M1688 diff_3307800_2085320# diff_3223440_2120840# diff_3343320_1672400# GND efet w=14800 l=8880
+ ad=0 pd=0 as=-1.88772e+09 ps=446960 
M1689 diff_3488360_1570280# Vdd Vdd GND efet w=11840 l=19240
+ ad=1.82679e+09 pd=242720 as=0 ps=0 
M1690 GND diff_3488360_1339400# diff_3488360_1570280# GND efet w=56240 l=7400
+ ad=0 pd=0 as=0 ps=0 
M1691 diff_3285600_2079400# diff_3267840_1873680# GND GND efet w=19240 l=7400
+ ad=0 pd=0 as=0 ps=0 
M1692 sync clk2 diff_3412880_1952120# GND efet w=14800 l=7400
+ ad=0 pd=0 as=2.32182e+08 ps=65120 
M1693 diff_3412880_1952120# diff_3412880_1952120# diff_3412880_1952120# GND efet w=1480 l=1480
+ ad=0 pd=0 as=0 ps=0 
M1694 diff_3412880_1952120# diff_3412880_1952120# diff_3412880_1952120# GND efet w=740 l=2220
+ ad=0 pd=0 as=0 ps=0 
M1695 GND diff_3267840_1873680# diff_2043880_2100120# GND efet w=362600 l=7400
+ ad=0 pd=0 as=-6.36592e+08 ps=1.31128e+06 
M1696 diff_2043880_2100120# diff_3196800_1889960# diff_2043880_2100120# GND efet w=68080 l=20720
+ ad=0 pd=0 as=0 ps=0 
M1697 diff_2043880_2100120# diff_3196800_1889960# Vdd GND efet w=19240 l=7400
+ ad=0 pd=0 as=0 ps=0 
M1698 diff_800680_2049800# diff_233840_991600# GND GND efet w=233840 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1699 GND diff_233840_991600# diff_1012320_1684240# GND efet w=233840 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1700 diff_1243200_1832240# diff_1238760_1824840# diff_1243200_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1701 diff_1268360_1832240# diff_1238760_1824840# diff_1268360_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1702 diff_1293520_1832240# diff_1238760_1824840# diff_1293520_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1703 diff_1318680_1832240# diff_1238760_1824840# diff_1318680_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1704 diff_1343840_1832240# diff_1238760_1824840# diff_1343840_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1705 diff_1369000_1832240# diff_1238760_1824840# diff_1369000_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1706 diff_1394160_1832240# diff_1238760_1824840# diff_1394160_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1707 diff_1419320_1832240# diff_1238760_1824840# diff_1419320_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1708 diff_1444480_1832240# diff_1238760_1824840# diff_1444480_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1709 diff_1469640_1832240# diff_1238760_1824840# diff_1469640_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1710 diff_1494800_1832240# diff_1238760_1824840# diff_1494800_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1711 diff_1519960_1832240# diff_1238760_1824840# diff_1519960_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1712 diff_1545120_1832240# diff_1238760_1824840# diff_1545120_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1713 diff_1570280_1832240# diff_1238760_1824840# diff_1570280_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1714 diff_1595440_1832240# diff_1238760_1824840# diff_1595440_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1715 diff_1620600_1832240# diff_1238760_1824840# diff_1620600_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1716 diff_1645760_1832240# diff_1238760_1824840# diff_1645760_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1717 diff_1670920_1832240# diff_1238760_1824840# diff_1670920_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1718 diff_1696080_1832240# diff_1238760_1824840# diff_1696080_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1719 diff_1721240_1832240# diff_1238760_1824840# diff_1721240_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1720 diff_1746400_1832240# diff_1238760_1824840# diff_1746400_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1721 diff_1771560_1832240# diff_1238760_1824840# diff_1771560_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1722 diff_1796720_1832240# diff_1238760_1824840# diff_1796720_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1723 diff_1821880_1832240# diff_1238760_1824840# diff_1821880_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1724 diff_1847040_1832240# diff_1238760_1824840# diff_1847040_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1725 diff_1872200_1832240# diff_1238760_1824840# diff_1872200_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1726 diff_1897360_1832240# diff_1238760_1824840# diff_1897360_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1727 diff_1922520_1832240# diff_1238760_1824840# diff_1922520_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1728 diff_1947680_1832240# diff_1238760_1824840# diff_1947680_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1729 diff_1972840_1832240# diff_1238760_1824840# diff_1972840_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1730 diff_1998000_1832240# diff_1238760_1824840# diff_1998000_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1731 diff_2023160_1832240# diff_1238760_1824840# diff_2023160_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1732 diff_2048320_1832240# diff_1238760_1824840# diff_2048320_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1733 diff_2073480_1832240# diff_1238760_1824840# diff_2073480_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1734 diff_2098640_1832240# diff_1238760_1824840# diff_2098640_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1735 diff_2123800_1832240# diff_1238760_1824840# diff_2123800_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1736 diff_2148960_1832240# diff_1238760_1824840# diff_2148960_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1737 diff_2174120_1832240# diff_1238760_1824840# diff_2174120_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1738 diff_2199280_1832240# diff_1238760_1824840# diff_2199280_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1739 diff_2224440_1832240# diff_1238760_1824840# diff_2224440_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1740 diff_2249600_1832240# diff_1238760_1824840# diff_2249600_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1741 diff_2274760_1832240# diff_1238760_1824840# diff_2274760_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1742 diff_2299920_1832240# diff_1238760_1824840# diff_2299920_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1743 diff_2325080_1832240# diff_1238760_1824840# diff_2325080_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1744 diff_2350240_1832240# diff_1238760_1824840# diff_2350240_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1745 diff_2375400_1832240# diff_1238760_1824840# diff_2375400_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1746 diff_2400560_1832240# diff_1238760_1824840# diff_2400560_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1747 diff_2425720_1832240# diff_1238760_1824840# diff_2425720_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1748 diff_2450880_1832240# diff_1238760_1824840# diff_2450880_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1749 diff_2476040_1832240# diff_1238760_1824840# diff_2476040_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1750 diff_2501200_1832240# diff_1238760_1824840# diff_2501200_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1751 diff_2526360_1832240# diff_1238760_1824840# diff_2526360_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1752 diff_2551520_1832240# diff_1238760_1824840# diff_2551520_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1753 diff_2576680_1832240# diff_1238760_1824840# diff_2576680_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1754 diff_2601840_1832240# diff_1238760_1824840# diff_2601840_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1755 diff_2627000_1832240# diff_1238760_1824840# diff_2627000_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1756 diff_2652160_1832240# diff_1238760_1824840# diff_2652160_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1757 diff_2677320_1832240# diff_1238760_1824840# diff_2677320_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1758 diff_2702480_1832240# diff_1238760_1824840# diff_2702480_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1759 diff_2727640_1832240# diff_1238760_1824840# diff_2727640_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1760 diff_2752800_1832240# diff_1238760_1824840# diff_2752800_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1761 diff_2777960_1832240# diff_1238760_1824840# diff_2777960_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1762 diff_2803120_1832240# diff_1238760_1824840# diff_2803120_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1763 diff_2828280_1832240# diff_1238760_1824840# diff_2828280_1805600# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1764 diff_1238760_1852960# Vdd Vdd GND efet w=7400 l=14800
+ ad=0 pd=0 as=0 ps=0 
M1765 diff_1243200_1805600# diff_1238760_1798200# diff_1243200_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1766 diff_1268360_1805600# diff_1238760_1798200# diff_1268360_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1767 diff_1293520_1805600# diff_1238760_1798200# diff_1293520_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1768 diff_1318680_1805600# diff_1238760_1798200# diff_1318680_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1769 diff_1343840_1805600# diff_1238760_1798200# diff_1343840_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1770 diff_1369000_1805600# diff_1238760_1798200# diff_1369000_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1771 diff_1394160_1805600# diff_1238760_1798200# diff_1394160_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1772 diff_1419320_1805600# diff_1238760_1798200# diff_1419320_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1773 diff_1444480_1805600# diff_1238760_1798200# diff_1444480_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1774 diff_1469640_1805600# diff_1238760_1798200# diff_1469640_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1775 diff_1494800_1805600# diff_1238760_1798200# diff_1494800_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1776 diff_1519960_1805600# diff_1238760_1798200# diff_1519960_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1777 diff_1545120_1805600# diff_1238760_1798200# diff_1545120_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1778 diff_1570280_1805600# diff_1238760_1798200# diff_1570280_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1779 diff_1595440_1805600# diff_1238760_1798200# diff_1595440_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1780 diff_1620600_1805600# diff_1238760_1798200# diff_1620600_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1781 diff_1645760_1805600# diff_1238760_1798200# diff_1645760_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1782 diff_1670920_1805600# diff_1238760_1798200# diff_1670920_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1783 diff_1696080_1805600# diff_1238760_1798200# diff_1696080_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1784 diff_1721240_1805600# diff_1238760_1798200# diff_1721240_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1785 diff_1746400_1805600# diff_1238760_1798200# diff_1746400_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1786 diff_1771560_1805600# diff_1238760_1798200# diff_1771560_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1787 diff_1796720_1805600# diff_1238760_1798200# diff_1796720_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1788 diff_1821880_1805600# diff_1238760_1798200# diff_1821880_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1789 diff_1847040_1805600# diff_1238760_1798200# diff_1847040_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1790 diff_1872200_1805600# diff_1238760_1798200# diff_1872200_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1791 diff_1897360_1805600# diff_1238760_1798200# diff_1897360_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1792 diff_1922520_1805600# diff_1238760_1798200# diff_1922520_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1793 diff_1947680_1805600# diff_1238760_1798200# diff_1947680_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1794 diff_1972840_1805600# diff_1238760_1798200# diff_1972840_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1795 diff_1998000_1805600# diff_1238760_1798200# diff_1998000_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1796 diff_2023160_1805600# diff_1238760_1798200# diff_2023160_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1797 diff_2048320_1805600# diff_1238760_1798200# diff_2048320_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1798 diff_2073480_1805600# diff_1238760_1798200# diff_2073480_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1799 diff_2098640_1805600# diff_1238760_1798200# diff_2098640_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1800 diff_2123800_1805600# diff_1238760_1798200# diff_2123800_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1801 diff_2148960_1805600# diff_1238760_1798200# diff_2148960_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1802 diff_2174120_1805600# diff_1238760_1798200# diff_2174120_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1803 diff_2199280_1805600# diff_1238760_1798200# diff_2199280_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1804 diff_2224440_1805600# diff_1238760_1798200# diff_2224440_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1805 diff_2249600_1805600# diff_1238760_1798200# diff_2249600_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1806 diff_2274760_1805600# diff_1238760_1798200# diff_2274760_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1807 diff_2299920_1805600# diff_1238760_1798200# diff_2299920_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1808 diff_2325080_1805600# diff_1238760_1798200# diff_2325080_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1809 diff_2350240_1805600# diff_1238760_1798200# diff_2350240_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1810 diff_2375400_1805600# diff_1238760_1798200# diff_2375400_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1811 diff_2400560_1805600# diff_1238760_1798200# diff_2400560_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1812 diff_2425720_1805600# diff_1238760_1798200# diff_2425720_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1813 diff_2450880_1805600# diff_1238760_1798200# diff_2450880_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1814 diff_2476040_1805600# diff_1238760_1798200# diff_2476040_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1815 diff_2501200_1805600# diff_1238760_1798200# diff_2501200_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1816 diff_2526360_1805600# diff_1238760_1798200# diff_2526360_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1817 diff_2551520_1805600# diff_1238760_1798200# diff_2551520_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1818 diff_2576680_1805600# diff_1238760_1798200# diff_2576680_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1819 diff_2601840_1805600# diff_1238760_1798200# diff_2601840_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1820 diff_2627000_1805600# diff_1238760_1798200# diff_2627000_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1821 diff_2652160_1805600# diff_1238760_1798200# diff_2652160_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1822 diff_2677320_1805600# diff_1238760_1798200# diff_2677320_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1823 diff_2702480_1805600# diff_1238760_1798200# diff_2702480_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1824 diff_2727640_1805600# diff_1238760_1798200# diff_2727640_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1825 diff_2752800_1805600# diff_1238760_1798200# diff_2752800_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1826 diff_2777960_1805600# diff_1238760_1798200# diff_2777960_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1827 diff_2803120_1805600# diff_1238760_1798200# diff_2803120_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1828 diff_2828280_1805600# diff_1238760_1798200# diff_2828280_1777480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1829 Vdd Vdd diff_1238760_1770080# GND efet w=7400 l=16280
+ ad=0 pd=0 as=1.29453e+09 ps=319680 
M1830 diff_1243200_1777480# diff_1238760_1770080# diff_1243200_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1831 diff_1268360_1777480# diff_1238760_1770080# diff_1268360_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1832 diff_1293520_1777480# diff_1238760_1770080# diff_1293520_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1833 diff_1318680_1777480# diff_1238760_1770080# diff_1318680_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1834 diff_1343840_1777480# diff_1238760_1770080# diff_1343840_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1835 diff_1369000_1777480# diff_1238760_1770080# diff_1369000_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1836 diff_1394160_1777480# diff_1238760_1770080# diff_1394160_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1837 diff_1419320_1777480# diff_1238760_1770080# diff_1419320_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1838 diff_1444480_1777480# diff_1238760_1770080# diff_1444480_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1839 diff_1469640_1777480# diff_1238760_1770080# diff_1469640_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1840 diff_1494800_1777480# diff_1238760_1770080# diff_1494800_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1841 diff_1519960_1777480# diff_1238760_1770080# diff_1519960_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1842 diff_1545120_1777480# diff_1238760_1770080# diff_1545120_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1843 diff_1570280_1777480# diff_1238760_1770080# diff_1570280_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1844 diff_1595440_1777480# diff_1238760_1770080# diff_1595440_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1845 diff_1620600_1777480# diff_1238760_1770080# diff_1620600_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1846 diff_1645760_1777480# diff_1238760_1770080# diff_1645760_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1847 diff_1670920_1777480# diff_1238760_1770080# diff_1670920_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1848 diff_1696080_1777480# diff_1238760_1770080# diff_1696080_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1849 diff_1721240_1777480# diff_1238760_1770080# diff_1721240_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1850 diff_1746400_1777480# diff_1238760_1770080# diff_1746400_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1851 diff_1771560_1777480# diff_1238760_1770080# diff_1771560_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1852 diff_1796720_1777480# diff_1238760_1770080# diff_1796720_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1853 diff_1821880_1777480# diff_1238760_1770080# diff_1821880_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1854 diff_1847040_1777480# diff_1238760_1770080# diff_1847040_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1855 diff_1872200_1777480# diff_1238760_1770080# diff_1872200_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1856 diff_1897360_1777480# diff_1238760_1770080# diff_1897360_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1857 diff_1922520_1777480# diff_1238760_1770080# diff_1922520_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1858 diff_1947680_1777480# diff_1238760_1770080# diff_1947680_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1859 diff_1972840_1777480# diff_1238760_1770080# diff_1972840_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1860 diff_1998000_1777480# diff_1238760_1770080# diff_1998000_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1861 diff_2023160_1777480# diff_1238760_1770080# diff_2023160_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1862 diff_2048320_1777480# diff_1238760_1770080# diff_2048320_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1863 diff_2073480_1777480# diff_1238760_1770080# diff_2073480_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1864 diff_2098640_1777480# diff_1238760_1770080# diff_2098640_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1865 diff_2123800_1777480# diff_1238760_1770080# diff_2123800_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1866 diff_2148960_1777480# diff_1238760_1770080# diff_2148960_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1867 diff_2174120_1777480# diff_1238760_1770080# diff_2174120_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1868 diff_2199280_1777480# diff_1238760_1770080# diff_2199280_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1869 diff_2224440_1777480# diff_1238760_1770080# diff_2224440_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1870 diff_2249600_1777480# diff_1238760_1770080# diff_2249600_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1871 diff_2274760_1777480# diff_1238760_1770080# diff_2274760_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1872 diff_2299920_1777480# diff_1238760_1770080# diff_2299920_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1873 diff_2325080_1777480# diff_1238760_1770080# diff_2325080_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1874 diff_2350240_1777480# diff_1238760_1770080# diff_2350240_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1875 diff_2375400_1777480# diff_1238760_1770080# diff_2375400_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1876 diff_2400560_1777480# diff_1238760_1770080# diff_2400560_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1877 diff_2425720_1777480# diff_1238760_1770080# diff_2425720_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1878 diff_2450880_1777480# diff_1238760_1770080# diff_2450880_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1879 diff_2476040_1777480# diff_1238760_1770080# diff_2476040_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1880 diff_2501200_1777480# diff_1238760_1770080# diff_2501200_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1881 diff_2526360_1777480# diff_1238760_1770080# diff_2526360_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1882 diff_2551520_1777480# diff_1238760_1770080# diff_2551520_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1883 diff_2576680_1777480# diff_1238760_1770080# diff_2576680_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1884 diff_2601840_1777480# diff_1238760_1770080# diff_2601840_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1885 diff_2627000_1777480# diff_1238760_1770080# diff_2627000_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1886 diff_2652160_1777480# diff_1238760_1770080# diff_2652160_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1887 diff_2677320_1777480# diff_1238760_1770080# diff_2677320_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1888 diff_2702480_1777480# diff_1238760_1770080# diff_2702480_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1889 diff_2727640_1777480# diff_1238760_1770080# diff_2727640_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1890 diff_2752800_1777480# diff_1238760_1770080# diff_2752800_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1891 diff_2777960_1777480# diff_1238760_1770080# diff_2777960_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1892 diff_2803120_1777480# diff_1238760_1770080# diff_2803120_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1893 diff_2828280_1777480# diff_1238760_1770080# diff_2828280_1750840# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1894 diff_991600_2049800# diff_233840_991600# GND GND efet w=235320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M1895 diff_1238760_1770080# diff_2940760_526880# diff_2920040_1842600# GND efet w=91760 l=7400
+ ad=0 pd=0 as=0 ps=0 
M1896 diff_2920040_1842600# diff_2976280_1228400# diff_1238760_1824840# GND efet w=103600 l=7400
+ ad=0 pd=0 as=1.7567e+09 ps=281200 
M1897 diff_1238760_1824840# Vdd Vdd GND efet w=8880 l=13320
+ ad=0 pd=0 as=0 ps=0 
M1898 Vdd Vdd diff_1238760_1798200# GND efet w=8880 l=14800
+ ad=0 pd=0 as=1.43252e+09 ps=304880 
M1899 diff_1243200_1750840# diff_1238760_1743440# diff_1243200_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1900 diff_1268360_1750840# diff_1238760_1743440# diff_1268360_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1901 diff_1293520_1750840# diff_1238760_1743440# diff_1293520_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1902 diff_1318680_1750840# diff_1238760_1743440# diff_1318680_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1903 diff_1343840_1750840# diff_1238760_1743440# diff_1343840_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1904 diff_1369000_1750840# diff_1238760_1743440# diff_1369000_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1905 diff_1394160_1750840# diff_1238760_1743440# diff_1394160_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1906 diff_1419320_1750840# diff_1238760_1743440# diff_1419320_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1907 diff_1444480_1750840# diff_1238760_1743440# diff_1444480_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1908 diff_1469640_1750840# diff_1238760_1743440# diff_1469640_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1909 diff_1494800_1750840# diff_1238760_1743440# diff_1494800_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1910 diff_1519960_1750840# diff_1238760_1743440# diff_1519960_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1911 diff_1545120_1750840# diff_1238760_1743440# diff_1545120_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1912 diff_1570280_1750840# diff_1238760_1743440# diff_1570280_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1913 diff_1595440_1750840# diff_1238760_1743440# diff_1595440_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1914 diff_1620600_1750840# diff_1238760_1743440# diff_1620600_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1915 diff_1645760_1750840# diff_1238760_1743440# diff_1645760_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1916 diff_1670920_1750840# diff_1238760_1743440# diff_1670920_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1917 diff_1696080_1750840# diff_1238760_1743440# diff_1696080_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1918 diff_1721240_1750840# diff_1238760_1743440# diff_1721240_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1919 diff_1746400_1750840# diff_1238760_1743440# diff_1746400_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1920 diff_1771560_1750840# diff_1238760_1743440# diff_1771560_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1921 diff_1796720_1750840# diff_1238760_1743440# diff_1796720_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1922 diff_1821880_1750840# diff_1238760_1743440# diff_1821880_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1923 diff_1847040_1750840# diff_1238760_1743440# diff_1847040_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1924 diff_1872200_1750840# diff_1238760_1743440# diff_1872200_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1925 diff_1897360_1750840# diff_1238760_1743440# diff_1897360_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1926 diff_1922520_1750840# diff_1238760_1743440# diff_1922520_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1927 diff_1947680_1750840# diff_1238760_1743440# diff_1947680_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1928 diff_1972840_1750840# diff_1238760_1743440# diff_1972840_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1929 diff_1998000_1750840# diff_1238760_1743440# diff_1998000_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1930 diff_2023160_1750840# diff_1238760_1743440# diff_2023160_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1931 diff_2048320_1750840# diff_1238760_1743440# diff_2048320_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1932 diff_2073480_1750840# diff_1238760_1743440# diff_2073480_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1933 diff_2098640_1750840# diff_1238760_1743440# diff_2098640_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1934 diff_2123800_1750840# diff_1238760_1743440# diff_2123800_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1935 diff_2148960_1750840# diff_1238760_1743440# diff_2148960_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1936 diff_2174120_1750840# diff_1238760_1743440# diff_2174120_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1937 diff_2199280_1750840# diff_1238760_1743440# diff_2199280_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1938 diff_2224440_1750840# diff_1238760_1743440# diff_2224440_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1939 diff_2249600_1750840# diff_1238760_1743440# diff_2249600_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1940 diff_2274760_1750840# diff_1238760_1743440# diff_2274760_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1941 diff_2299920_1750840# diff_1238760_1743440# diff_2299920_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1942 diff_2325080_1750840# diff_1238760_1743440# diff_2325080_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1943 diff_2350240_1750840# diff_1238760_1743440# diff_2350240_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1944 diff_2375400_1750840# diff_1238760_1743440# diff_2375400_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1945 diff_2400560_1750840# diff_1238760_1743440# diff_2400560_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1946 diff_2425720_1750840# diff_1238760_1743440# diff_2425720_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1947 diff_2450880_1750840# diff_1238760_1743440# diff_2450880_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1948 diff_2476040_1750840# diff_1238760_1743440# diff_2476040_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1949 diff_2501200_1750840# diff_1238760_1743440# diff_2501200_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1950 diff_2526360_1750840# diff_1238760_1743440# diff_2526360_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1951 diff_2551520_1750840# diff_1238760_1743440# diff_2551520_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1952 diff_2576680_1750840# diff_1238760_1743440# diff_2576680_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1953 diff_2601840_1750840# diff_1238760_1743440# diff_2601840_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1954 diff_2627000_1750840# diff_1238760_1743440# diff_2627000_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1955 diff_2652160_1750840# diff_1238760_1743440# diff_2652160_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1956 diff_2677320_1750840# diff_1238760_1743440# diff_2677320_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1957 diff_2702480_1750840# diff_1238760_1743440# diff_2702480_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1958 diff_2727640_1750840# diff_1238760_1743440# diff_2727640_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1959 diff_2752800_1750840# diff_1238760_1743440# diff_2752800_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1960 diff_2777960_1750840# diff_1238760_1743440# diff_2777960_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1961 diff_2803120_1750840# diff_1238760_1743440# diff_2803120_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1962 diff_2828280_1750840# diff_1238760_1743440# diff_2828280_1722720# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M1963 diff_2920040_1736040# diff_2912640_526880# diff_1238760_1743440# GND efet w=106560 l=7400
+ ad=1.52493e+09 pd=899840 as=1.47195e+09 ps=284160 
M1964 diff_1238760_1798200# diff_2998480_1207680# diff_2920040_1842600# GND efet w=97680 l=7400
+ ad=0 pd=0 as=0 ps=0 
M1965 diff_1243200_1722720# diff_1238760_1715320# diff_1243200_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1966 diff_1268360_1722720# diff_1238760_1715320# diff_1268360_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1967 diff_1293520_1722720# diff_1238760_1715320# diff_1293520_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1968 diff_1318680_1722720# diff_1238760_1715320# diff_1318680_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1969 diff_1343840_1722720# diff_1238760_1715320# diff_1343840_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1970 diff_1369000_1722720# diff_1238760_1715320# diff_1369000_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1971 diff_1394160_1722720# diff_1238760_1715320# diff_1394160_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1972 diff_1419320_1722720# diff_1238760_1715320# diff_1419320_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1973 diff_1444480_1722720# diff_1238760_1715320# diff_1444480_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1974 diff_1469640_1722720# diff_1238760_1715320# diff_1469640_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1975 diff_1494800_1722720# diff_1238760_1715320# diff_1494800_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1976 diff_1519960_1722720# diff_1238760_1715320# diff_1519960_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1977 diff_1545120_1722720# diff_1238760_1715320# diff_1545120_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1978 diff_1570280_1722720# diff_1238760_1715320# diff_1570280_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1979 diff_1595440_1722720# diff_1238760_1715320# diff_1595440_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1980 diff_1620600_1722720# diff_1238760_1715320# diff_1620600_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1981 diff_1645760_1722720# diff_1238760_1715320# diff_1645760_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1982 diff_1670920_1722720# diff_1238760_1715320# diff_1670920_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1983 diff_1696080_1722720# diff_1238760_1715320# diff_1696080_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1984 diff_1721240_1722720# diff_1238760_1715320# diff_1721240_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1985 diff_1746400_1722720# diff_1238760_1715320# diff_1746400_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1986 diff_1771560_1722720# diff_1238760_1715320# diff_1771560_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1987 diff_1796720_1722720# diff_1238760_1715320# diff_1796720_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1988 diff_1821880_1722720# diff_1238760_1715320# diff_1821880_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1989 diff_1847040_1722720# diff_1238760_1715320# diff_1847040_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1990 diff_1872200_1722720# diff_1238760_1715320# diff_1872200_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1991 diff_1897360_1722720# diff_1238760_1715320# diff_1897360_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1992 diff_1922520_1722720# diff_1238760_1715320# diff_1922520_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1993 diff_1947680_1722720# diff_1238760_1715320# diff_1947680_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1994 diff_1972840_1722720# diff_1238760_1715320# diff_1972840_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1995 diff_1998000_1722720# diff_1238760_1715320# diff_1998000_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1996 diff_2023160_1722720# diff_1238760_1715320# diff_2023160_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1997 diff_2048320_1722720# diff_1238760_1715320# diff_2048320_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1998 diff_2073480_1722720# diff_1238760_1715320# diff_2073480_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M1999 diff_2098640_1722720# diff_1238760_1715320# diff_2098640_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2000 diff_2123800_1722720# diff_1238760_1715320# diff_2123800_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2001 diff_2148960_1722720# diff_1238760_1715320# diff_2148960_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2002 diff_2174120_1722720# diff_1238760_1715320# diff_2174120_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2003 diff_2199280_1722720# diff_1238760_1715320# diff_2199280_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2004 diff_2224440_1722720# diff_1238760_1715320# diff_2224440_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2005 diff_2249600_1722720# diff_1238760_1715320# diff_2249600_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2006 diff_2274760_1722720# diff_1238760_1715320# diff_2274760_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2007 diff_2299920_1722720# diff_1238760_1715320# diff_2299920_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2008 diff_2325080_1722720# diff_1238760_1715320# diff_2325080_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2009 diff_2350240_1722720# diff_1238760_1715320# diff_2350240_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2010 diff_2375400_1722720# diff_1238760_1715320# diff_2375400_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2011 diff_2400560_1722720# diff_1238760_1715320# diff_2400560_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2012 diff_2425720_1722720# diff_1238760_1715320# diff_2425720_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2013 diff_2450880_1722720# diff_1238760_1715320# diff_2450880_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2014 diff_2476040_1722720# diff_1238760_1715320# diff_2476040_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2015 diff_2501200_1722720# diff_1238760_1715320# diff_2501200_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2016 diff_2526360_1722720# diff_1238760_1715320# diff_2526360_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2017 diff_2551520_1722720# diff_1238760_1715320# diff_2551520_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2018 diff_2576680_1722720# diff_1238760_1715320# diff_2576680_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2019 diff_2601840_1722720# diff_1238760_1715320# diff_2601840_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2020 diff_2627000_1722720# diff_1238760_1715320# diff_2627000_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2021 diff_2652160_1722720# diff_1238760_1715320# diff_2652160_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2022 diff_2677320_1722720# diff_1238760_1715320# diff_2677320_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2023 diff_2702480_1722720# diff_1238760_1715320# diff_2702480_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2024 diff_2727640_1722720# diff_1238760_1715320# diff_2727640_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2025 diff_2752800_1722720# diff_1238760_1715320# diff_2752800_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2026 diff_2777960_1722720# diff_1238760_1715320# diff_2777960_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2027 diff_2803120_1722720# diff_1238760_1715320# diff_2803120_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2028 diff_2828280_1722720# diff_1238760_1715320# diff_2828280_1696080# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2029 diff_1238760_1743440# Vdd Vdd GND efet w=7400 l=14800
+ ad=0 pd=0 as=0 ps=0 
M2030 diff_1243200_1696080# diff_1238760_1688680# diff_1243200_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2031 diff_1268360_1696080# diff_1238760_1688680# diff_1268360_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2032 diff_1293520_1696080# diff_1238760_1688680# diff_1293520_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2033 diff_1318680_1696080# diff_1238760_1688680# diff_1318680_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2034 diff_1343840_1696080# diff_1238760_1688680# diff_1343840_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2035 diff_1369000_1696080# diff_1238760_1688680# diff_1369000_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2036 diff_1394160_1696080# diff_1238760_1688680# diff_1394160_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2037 diff_1419320_1696080# diff_1238760_1688680# diff_1419320_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2038 diff_1444480_1696080# diff_1238760_1688680# diff_1444480_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2039 diff_1469640_1696080# diff_1238760_1688680# diff_1469640_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2040 diff_1494800_1696080# diff_1238760_1688680# diff_1494800_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2041 diff_1519960_1696080# diff_1238760_1688680# diff_1519960_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2042 diff_1545120_1696080# diff_1238760_1688680# diff_1545120_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2043 diff_1570280_1696080# diff_1238760_1688680# diff_1570280_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2044 diff_1595440_1696080# diff_1238760_1688680# diff_1595440_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2045 diff_1620600_1696080# diff_1238760_1688680# diff_1620600_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2046 diff_1645760_1696080# diff_1238760_1688680# diff_1645760_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2047 diff_1670920_1696080# diff_1238760_1688680# diff_1670920_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2048 diff_1696080_1696080# diff_1238760_1688680# diff_1696080_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2049 diff_1721240_1696080# diff_1238760_1688680# diff_1721240_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2050 diff_1746400_1696080# diff_1238760_1688680# diff_1746400_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2051 diff_1771560_1696080# diff_1238760_1688680# diff_1771560_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2052 diff_1796720_1696080# diff_1238760_1688680# diff_1796720_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2053 diff_1821880_1696080# diff_1238760_1688680# diff_1821880_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2054 diff_1847040_1696080# diff_1238760_1688680# diff_1847040_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2055 diff_1872200_1696080# diff_1238760_1688680# diff_1872200_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2056 diff_1897360_1696080# diff_1238760_1688680# diff_1897360_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2057 diff_1922520_1696080# diff_1238760_1688680# diff_1922520_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2058 diff_1947680_1696080# diff_1238760_1688680# diff_1947680_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2059 diff_1972840_1696080# diff_1238760_1688680# diff_1972840_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2060 diff_1998000_1696080# diff_1238760_1688680# diff_1998000_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2061 diff_2023160_1696080# diff_1238760_1688680# diff_2023160_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2062 diff_2048320_1696080# diff_1238760_1688680# diff_2048320_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2063 diff_2073480_1696080# diff_1238760_1688680# diff_2073480_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2064 diff_2098640_1696080# diff_1238760_1688680# diff_2098640_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2065 diff_2123800_1696080# diff_1238760_1688680# diff_2123800_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2066 diff_2148960_1696080# diff_1238760_1688680# diff_2148960_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2067 diff_2174120_1696080# diff_1238760_1688680# diff_2174120_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2068 diff_2199280_1696080# diff_1238760_1688680# diff_2199280_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2069 diff_2224440_1696080# diff_1238760_1688680# diff_2224440_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2070 diff_2249600_1696080# diff_1238760_1688680# diff_2249600_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2071 diff_2274760_1696080# diff_1238760_1688680# diff_2274760_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2072 diff_2299920_1696080# diff_1238760_1688680# diff_2299920_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2073 diff_2325080_1696080# diff_1238760_1688680# diff_2325080_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2074 diff_2350240_1696080# diff_1238760_1688680# diff_2350240_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2075 diff_2375400_1696080# diff_1238760_1688680# diff_2375400_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2076 diff_2400560_1696080# diff_1238760_1688680# diff_2400560_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2077 diff_2425720_1696080# diff_1238760_1688680# diff_2425720_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2078 diff_2450880_1696080# diff_1238760_1688680# diff_2450880_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2079 diff_2476040_1696080# diff_1238760_1688680# diff_2476040_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2080 diff_2501200_1696080# diff_1238760_1688680# diff_2501200_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2081 diff_2526360_1696080# diff_1238760_1688680# diff_2526360_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2082 diff_2551520_1696080# diff_1238760_1688680# diff_2551520_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2083 diff_2576680_1696080# diff_1238760_1688680# diff_2576680_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2084 diff_2601840_1696080# diff_1238760_1688680# diff_2601840_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2085 diff_2627000_1696080# diff_1238760_1688680# diff_2627000_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2086 diff_2652160_1696080# diff_1238760_1688680# diff_2652160_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2087 diff_2677320_1696080# diff_1238760_1688680# diff_2677320_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2088 diff_2702480_1696080# diff_1238760_1688680# diff_2702480_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2089 diff_2727640_1696080# diff_1238760_1688680# diff_2727640_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2090 diff_2752800_1696080# diff_1238760_1688680# diff_2752800_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2091 diff_2777960_1696080# diff_1238760_1688680# diff_2777960_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2092 diff_2803120_1696080# diff_1238760_1688680# diff_2803120_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2093 diff_2828280_1696080# diff_1238760_1688680# diff_2828280_1667960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2094 d3 clk2 diff_411440_1660560# GND efet w=14800 l=8880
+ ad=0 pd=0 as=1.53328e+08 ps=50320 
M2095 d2 clk2 diff_602360_1660560# GND efet w=14800 l=8880
+ ad=0 pd=0 as=1.53328e+08 ps=50320 
M2096 d1 clk2 diff_794760_1660560# GND efet w=14800 l=8880
+ ad=0 pd=0 as=1.53328e+08 ps=50320 
M2097 d0 clk2 diff_985680_1660560# GND efet w=14800 l=8880
+ ad=0 pd=0 as=1.53328e+08 ps=50320 
M2098 Vdd Vdd diff_1238760_1660560# GND efet w=7400 l=16280
+ ad=0 pd=0 as=1.29453e+09 ps=319680 
M2099 diff_411440_1660560# diff_190920_1013800# diff_411440_1576200# GND efet w=14800 l=8880
+ ad=0 pd=0 as=-1.78915e+09 ps=438080 
M2100 diff_602360_1660560# diff_190920_1013800# diff_602360_1574720# GND efet w=14800 l=8880
+ ad=0 pd=0 as=-1.84391e+09 ps=435120 
M2101 diff_794760_1660560# diff_190920_1013800# diff_794760_1574720# GND efet w=14800 l=8880
+ ad=0 pd=0 as=-1.75629e+09 ps=435120 
M2102 diff_985680_1660560# diff_190920_1013800# diff_985680_1574720# GND efet w=14800 l=8880
+ ad=0 pd=0 as=-1.77163e+09 ps=441040 
M2103 diff_1243200_1667960# diff_1238760_1660560# diff_1243200_1628000# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2104 diff_1268360_1667960# diff_1238760_1660560# diff_1263920_1558440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2105 diff_1293520_1667960# diff_1238760_1660560# diff_1293520_1630960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2106 diff_1318680_1667960# diff_1238760_1660560# diff_1318680_1580640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2107 diff_1343840_1667960# diff_1238760_1660560# diff_1343840_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2108 diff_1369000_1667960# diff_1238760_1660560# diff_1369000_1556960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2109 diff_1394160_1667960# diff_1238760_1660560# diff_1394160_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2110 diff_1419320_1667960# diff_1238760_1660560# diff_1419320_1580640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2111 diff_1444480_1667960# diff_1238760_1660560# diff_1444480_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2112 diff_1469640_1667960# diff_1238760_1660560# diff_1469640_1556960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2113 diff_1494800_1667960# diff_1238760_1660560# diff_1494800_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2114 diff_1519960_1667960# diff_1238760_1660560# diff_1519960_1580640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2115 diff_1545120_1667960# diff_1238760_1660560# diff_1545120_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2116 diff_1570280_1667960# diff_1238760_1660560# diff_1570280_1556960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2117 diff_1595440_1667960# diff_1238760_1660560# diff_1595440_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2118 diff_1620600_1667960# diff_1238760_1660560# diff_1620600_1580640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2119 diff_1645760_1667960# diff_1238760_1660560# diff_1645760_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2120 diff_1670920_1667960# diff_1238760_1660560# diff_1670920_1556960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2121 diff_1696080_1667960# diff_1238760_1660560# diff_1696080_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2122 diff_1721240_1667960# diff_1238760_1660560# diff_1721240_1580640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2123 diff_1746400_1667960# diff_1238760_1660560# diff_1746400_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2124 diff_1771560_1667960# diff_1238760_1660560# diff_1771560_1556960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2125 diff_1796720_1667960# diff_1238760_1660560# diff_1796720_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2126 diff_1821880_1667960# diff_1238760_1660560# diff_1821880_1580640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2127 diff_1847040_1667960# diff_1238760_1660560# diff_1847040_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2128 diff_1872200_1667960# diff_1238760_1660560# diff_1872200_1556960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2129 diff_1897360_1667960# diff_1238760_1660560# diff_1897360_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2130 diff_1922520_1667960# diff_1238760_1660560# diff_1922520_1580640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2131 diff_1947680_1667960# diff_1238760_1660560# diff_1947680_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2132 diff_1972840_1667960# diff_1238760_1660560# diff_1972840_1556960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2133 diff_1998000_1667960# diff_1238760_1660560# diff_1998000_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2134 diff_2023160_1667960# diff_1238760_1660560# diff_2023160_1580640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2135 diff_2048320_1667960# diff_1238760_1660560# diff_2048320_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2136 diff_2073480_1667960# diff_1238760_1660560# diff_2073480_1556960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2137 diff_2098640_1667960# diff_1238760_1660560# diff_2098640_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2138 diff_2123800_1667960# diff_1238760_1660560# diff_2123800_1580640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2139 diff_2148960_1667960# diff_1238760_1660560# diff_2148960_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2140 diff_2174120_1667960# diff_1238760_1660560# diff_2174120_1556960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2141 diff_2199280_1667960# diff_1238760_1660560# diff_2199280_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2142 diff_2224440_1667960# diff_1238760_1660560# diff_2224440_1580640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2143 diff_2249600_1667960# diff_1238760_1660560# diff_2249600_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2144 diff_2274760_1667960# diff_1238760_1660560# diff_2274760_1556960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2145 diff_2299920_1667960# diff_1238760_1660560# diff_2299920_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2146 diff_2325080_1667960# diff_1238760_1660560# diff_2325080_1580640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2147 diff_2350240_1667960# diff_1238760_1660560# diff_2350240_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2148 diff_2375400_1667960# diff_1238760_1660560# diff_2375400_1556960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2149 diff_2400560_1667960# diff_1238760_1660560# diff_2400560_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2150 diff_2425720_1667960# diff_1238760_1660560# diff_2425720_1580640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2151 diff_2450880_1667960# diff_1238760_1660560# diff_2450880_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2152 diff_2476040_1667960# diff_1238760_1660560# diff_2476040_1556960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2153 diff_2501200_1667960# diff_1238760_1660560# diff_2501200_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2154 diff_2526360_1667960# diff_1238760_1660560# diff_2526360_1580640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2155 diff_2551520_1667960# diff_1238760_1660560# diff_2551520_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2156 diff_2576680_1667960# diff_1238760_1660560# diff_2576680_1556960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2157 diff_2601840_1667960# diff_1238760_1660560# diff_2601840_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2158 diff_2627000_1667960# diff_1238760_1660560# diff_2627000_1580640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2159 diff_2652160_1667960# diff_1238760_1660560# diff_2652160_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2160 diff_2677320_1667960# diff_1238760_1660560# diff_2677320_1556960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2161 diff_2702480_1667960# diff_1238760_1660560# diff_2702480_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2162 diff_2727640_1667960# diff_1238760_1660560# diff_2727640_1580640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2163 diff_2752800_1667960# diff_1238760_1660560# diff_2752800_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2164 diff_2777960_1667960# diff_1238760_1660560# diff_2777960_1556960# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2165 diff_2803120_1667960# diff_1238760_1660560# diff_2803120_1629480# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2166 diff_2828280_1667960# diff_1238760_1660560# diff_2828280_1580640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=1.92755e+08 ps=56240 
M2167 diff_346320_1623560# diff_190920_1013800# GND GND efet w=22200 l=8880
+ ad=3.92082e+08 pd=88800 as=0 ps=0 
M2168 diff_411440_1576200# diff_411440_1576200# diff_411440_1576200# GND efet w=4440 l=4440
+ ad=0 pd=0 as=0 ps=0 
M2169 Vdd Vdd diff_346320_1623560# GND efet w=5180 l=51060
+ ad=0 pd=0 as=0 ps=0 
M2170 GND GND sync GND efet w=142820 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2171 diff_414400_1443000# diff_411440_1576200# GND GND efet w=94720 l=8880
+ ad=1.14339e+09 pd=272320 as=0 ps=0 
M2172 diff_602360_1574720# diff_602360_1574720# diff_602360_1574720# GND efet w=4440 l=4440
+ ad=0 pd=0 as=0 ps=0 
M2173 diff_411440_1576200# diff_411440_1576200# diff_411440_1576200# GND efet w=2960 l=2960
+ ad=0 pd=0 as=0 ps=0 
M2174 GND diff_414400_1443000# diff_438080_1602840# GND efet w=62160 l=7400
+ ad=0 pd=0 as=2.09183e+09 ps=426240 
M2175 diff_438080_1602840# diff_346320_1623560# diff_411440_1576200# GND efet w=14800 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2176 diff_606800_1443000# diff_602360_1574720# GND GND efet w=94720 l=8880
+ ad=1.13244e+09 pd=272320 as=0 ps=0 
M2177 diff_794760_1574720# diff_794760_1574720# diff_794760_1574720# GND efet w=2960 l=2960
+ ad=0 pd=0 as=0 ps=0 
M2178 diff_602360_1574720# diff_602360_1574720# diff_602360_1574720# GND efet w=2960 l=2960
+ ad=0 pd=0 as=0 ps=0 
M2179 GND diff_606800_1443000# diff_627520_1602840# GND efet w=62160 l=7400
+ ad=0 pd=0 as=2.09402e+09 ps=423280 
M2180 diff_627520_1602840# diff_346320_1623560# diff_602360_1574720# GND efet w=14800 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2181 diff_797720_1443000# diff_794760_1574720# GND GND efet w=93240 l=8880
+ ad=1.2091e+09 pd=269360 as=0 ps=0 
M2182 diff_1238760_1660560# diff_2940760_526880# diff_2920040_1736040# GND efet w=91760 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2183 diff_2920040_1736040# diff_2976280_1228400# diff_1238760_1715320# GND efet w=105080 l=7400
+ ad=0 pd=0 as=1.74575e+09 ps=281200 
M2184 diff_1238760_1715320# Vdd Vdd GND efet w=8880 l=13320
+ ad=0 pd=0 as=0 ps=0 
M2185 Vdd Vdd diff_1238760_1688680# GND efet w=8880 l=16280
+ ad=0 pd=0 as=1.43252e+09 ps=304880 
M2186 diff_985680_1574720# diff_985680_1574720# diff_985680_1574720# GND efet w=4440 l=4440
+ ad=0 pd=0 as=0 ps=0 
M2187 diff_794760_1574720# diff_794760_1574720# diff_794760_1574720# GND efet w=1480 l=1480
+ ad=0 pd=0 as=0 ps=0 
M2188 GND diff_797720_1443000# diff_821400_1602840# GND efet w=62160 l=8880
+ ad=0 pd=0 as=2.04145e+09 ps=420320 
M2189 diff_821400_1602840# diff_346320_1623560# diff_794760_1574720# GND efet w=14800 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2190 diff_988640_1443000# diff_985680_1574720# GND GND efet w=94720 l=8880
+ ad=1.13244e+09 pd=269360 as=0 ps=0 
M2191 diff_985680_1574720# diff_985680_1574720# diff_985680_1574720# GND efet w=2960 l=2960
+ ad=0 pd=0 as=0 ps=0 
M2192 GND diff_988640_1443000# diff_1012320_1602840# GND efet w=62160 l=7400
+ ad=0 pd=0 as=2.08088e+09 ps=423280 
M2193 diff_1012320_1602840# diff_346320_1623560# diff_985680_1574720# GND efet w=14800 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2194 diff_411440_1576200# cl GND GND efet w=44400 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2195 GND cl diff_411440_1576200# GND efet w=44400 l=10360
+ ad=0 pd=0 as=0 ps=0 
M2196 diff_411440_1576200# diff_321160_969400# GND GND efet w=58460 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2197 diff_414400_1443000# Vdd Vdd GND efet w=7400 l=19240
+ ad=0 pd=0 as=0 ps=0 
M2198 diff_438080_1602840# Vdd Vdd GND efet w=7400 l=17760
+ ad=0 pd=0 as=0 ps=0 
M2199 Vdd Vdd Vdd GND efet w=2960 l=2960
+ ad=0 pd=0 as=0 ps=0 
M2200 Vdd Vdd Vdd GND efet w=2220 l=2960
+ ad=0 pd=0 as=0 ps=0 
M2201 diff_602360_1574720# cl GND GND efet w=44400 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2202 GND cl diff_602360_1574720# GND efet w=44400 l=10360
+ ad=0 pd=0 as=0 ps=0 
M2203 GND diff_1243200_1628000# diff_1229880_1524400# GND efet w=35520 l=7400
+ ad=0 pd=0 as=1.20472e+09 ps=239760 
M2204 diff_1274280_1562880# diff_1263920_1558440# GND GND efet w=56980 l=8880
+ ad=5.60742e+08 pd=130240 as=0 ps=0 
M2205 GND diff_1293520_1630960# diff_1278720_1482960# GND efet w=48840 l=7400
+ ad=0 pd=0 as=1.14777e+09 ps=236800 
M2206 diff_1326080_1583600# diff_1318680_1580640# GND GND efet w=48840 l=7400
+ ad=9.74728e+08 pd=230880 as=0 ps=0 
M2207 GND diff_1343840_1629480# diff_1324600_1456320# GND efet w=43660 l=8880
+ ad=0 pd=0 as=1.01635e+09 ps=216080 
M2208 GND diff_1394160_1629480# diff_1376400_1481480# GND efet w=48840 l=7400
+ ad=0 pd=0 as=1.15434e+09 ps=242720 
M2209 diff_1426720_1583600# diff_1419320_1580640# GND GND efet w=48840 l=7400
+ ad=1.00539e+09 pd=230880 as=0 ps=0 
M2210 diff_1376400_1561400# diff_1369000_1556960# GND GND efet w=43660 l=8140
+ ad=5.01602e+08 pd=115440 as=0 ps=0 
M2211 GND diff_1444480_1629480# diff_1425240_1456320# GND efet w=43660 l=8880
+ ad=0 pd=0 as=1.02511e+09 ps=216080 
M2212 GND diff_1494800_1629480# diff_1477040_1482960# GND efet w=48840 l=7400
+ ad=0 pd=0 as=1.18063e+09 ps=242720 
M2213 diff_1527360_1583600# diff_1519960_1580640# GND GND efet w=48840 l=7400
+ ad=9.96632e+08 pd=230880 as=0 ps=0 
M2214 diff_1477040_1561400# diff_1469640_1556960# GND GND efet w=43660 l=8140
+ ad=5.01602e+08 pd=115440 as=0 ps=0 
M2215 GND diff_1545120_1629480# diff_1524400_1456320# GND efet w=43660 l=8880
+ ad=0 pd=0 as=1.0733e+09 ps=219040 
M2216 GND diff_1595440_1629480# diff_1576200_1482960# GND efet w=48840 l=7400
+ ad=0 pd=0 as=1.2091e+09 ps=242720 
M2217 diff_1628000_1583600# diff_1620600_1580640# GND GND efet w=48840 l=7400
+ ad=1.04482e+09 pd=233840 as=0 ps=0 
M2218 diff_1577680_1561400# diff_1570280_1556960# GND GND efet w=43660 l=8140
+ ad=5.01602e+08 pd=115440 as=0 ps=0 
M2219 GND diff_1645760_1629480# diff_1625040_1456320# GND efet w=43660 l=8880
+ ad=0 pd=0 as=1.08206e+09 ps=219040 
M2220 GND diff_1696080_1629480# diff_1676840_1481480# GND efet w=48840 l=7400
+ ad=0 pd=0 as=1.23977e+09 ps=248640 
M2221 diff_1728640_1583600# diff_1721240_1580640# GND GND efet w=48840 l=7400
+ ad=9.06826e+08 pd=227920 as=0 ps=0 
M2222 diff_1678320_1561400# diff_1670920_1556960# GND GND efet w=43660 l=8140
+ ad=5.01602e+08 pd=115440 as=0 ps=0 
M2223 GND diff_1746400_1629480# diff_1727160_1456320# GND efet w=43660 l=8880
+ ad=0 pd=0 as=9.59395e+08 ps=213120 
M2224 GND diff_1796720_1629480# diff_1778960_1482960# GND efet w=48840 l=7400
+ ad=0 pd=0 as=1.0952e+09 ps=236800 
M2225 diff_1829280_1583600# diff_1821880_1580640# GND GND efet w=48840 l=7400
+ ad=9.44062e+08 pd=227920 as=0 ps=0 
M2226 diff_1778960_1561400# diff_1771560_1556960# GND GND efet w=43660 l=8140
+ ad=5.01602e+08 pd=115440 as=0 ps=0 
M2227 GND diff_1847040_1629480# diff_1827800_1456320# GND efet w=43660 l=8880
+ ad=0 pd=0 as=9.68157e+08 ps=213120 
M2228 GND diff_1897360_1629480# diff_1879600_1482960# GND efet w=48840 l=7400
+ ad=0 pd=0 as=1.12368e+09 ps=239760 
M2229 diff_1929920_1583600# diff_1922520_1580640# GND GND efet w=48840 l=7400
+ ad=9.06826e+08 pd=227920 as=0 ps=0 
M2230 diff_1879600_1561400# diff_1872200_1556960# GND GND efet w=43660 l=8140
+ ad=5.01602e+08 pd=115440 as=0 ps=0 
M2231 GND diff_1947680_1629480# diff_1928440_1456320# GND efet w=43660 l=8880
+ ad=0 pd=0 as=9.59395e+08 ps=213120 
M2232 GND diff_1998000_1629480# diff_1980240_1482960# GND efet w=48840 l=7400
+ ad=0 pd=0 as=1.0952e+09 ps=236800 
M2233 diff_2030560_1583600# diff_2023160_1580640# GND GND efet w=48840 l=7400
+ ad=9.50634e+08 pd=227920 as=0 ps=0 
M2234 diff_1980240_1561400# diff_1972840_1556960# GND GND efet w=43660 l=8140
+ ad=5.01602e+08 pd=115440 as=0 ps=0 
M2235 GND diff_2048320_1629480# diff_2029080_1456320# GND efet w=43660 l=8880
+ ad=0 pd=0 as=9.68157e+08 ps=213120 
M2236 GND diff_2098640_1629480# diff_2080880_1482960# GND efet w=48840 l=7400
+ ad=0 pd=0 as=1.12368e+09 ps=239760 
M2237 diff_2131200_1583600# diff_2123800_1580640# GND GND efet w=48840 l=7400
+ ad=9.68157e+08 pd=230880 as=0 ps=0 
M2238 diff_2080880_1561400# diff_2073480_1556960# GND GND efet w=43660 l=8140
+ ad=5.01602e+08 pd=115440 as=0 ps=0 
M2239 GND diff_2148960_1629480# diff_2131200_1456320# GND efet w=43660 l=8880
+ ad=0 pd=0 as=1.01635e+09 ps=216080 
M2240 GND diff_2199280_1629480# diff_2183000_1482960# GND efet w=48840 l=7400
+ ad=0 pd=0 as=1.15215e+09 ps=239760 
M2241 diff_2231840_1583600# diff_2224440_1580640# GND GND efet w=48840 l=7400
+ ad=1.00977e+09 pd=230880 as=0 ps=0 
M2242 diff_2181520_1561400# diff_2174120_1556960# GND GND efet w=43660 l=8140
+ ad=5.01602e+08 pd=115440 as=0 ps=0 
M2243 GND diff_2249600_1629480# diff_2231840_1456320# GND efet w=43660 l=8880
+ ad=0 pd=0 as=1.02511e+09 ps=216080 
M2244 GND diff_2299920_1629480# diff_2283640_1482960# GND efet w=48840 l=7400
+ ad=0 pd=0 as=1.18063e+09 ps=242720 
M2245 diff_2332480_1583600# diff_2325080_1580640# GND GND efet w=48840 l=7400
+ ad=9.65966e+08 pd=230880 as=0 ps=0 
M2246 diff_2282160_1561400# diff_2274760_1556960# GND GND efet w=43660 l=8140
+ ad=5.01602e+08 pd=115440 as=0 ps=0 
M2247 GND diff_2350240_1629480# diff_2331000_1456320# GND efet w=43660 l=8880
+ ad=0 pd=0 as=1.01635e+09 ps=216080 
M2248 GND diff_2400560_1629480# diff_2382800_1482960# GND efet w=48840 l=7400
+ ad=0 pd=0 as=1.15215e+09 ps=239760 
M2249 diff_2433120_1583600# diff_2425720_1580640# GND GND efet w=48840 l=7400
+ ad=1.00539e+09 pd=230880 as=0 ps=0 
M2250 diff_2382800_1561400# diff_2375400_1556960# GND GND efet w=43660 l=8140
+ ad=5.01602e+08 pd=115440 as=0 ps=0 
M2251 GND diff_2450880_1629480# diff_2431640_1456320# GND efet w=43660 l=8880
+ ad=0 pd=0 as=1.02511e+09 ps=216080 
M2252 GND diff_2501200_1629480# diff_2483440_1482960# GND efet w=48840 l=7400
+ ad=0 pd=0 as=1.18063e+09 ps=242720 
M2253 diff_2533760_1583600# diff_2526360_1580640# GND GND efet w=48840 l=7400
+ ad=9.65966e+08 pd=230880 as=0 ps=0 
M2254 diff_2483440_1561400# diff_2476040_1556960# GND GND efet w=43660 l=8140
+ ad=5.01602e+08 pd=115440 as=0 ps=0 
M2255 GND diff_2551520_1629480# diff_2532280_1456320# GND efet w=43660 l=8880
+ ad=0 pd=0 as=1.01635e+09 ps=216080 
M2256 GND diff_2601840_1629480# diff_2584080_1482960# GND efet w=48840 l=7400
+ ad=0 pd=0 as=1.15215e+09 ps=239760 
M2257 diff_2634400_1583600# diff_2627000_1580640# GND GND efet w=48840 l=7400
+ ad=1.00539e+09 pd=230880 as=0 ps=0 
M2258 diff_2584080_1561400# diff_2576680_1556960# GND GND efet w=43660 l=8140
+ ad=5.01602e+08 pd=115440 as=0 ps=0 
M2259 GND diff_2652160_1629480# diff_2632920_1456320# GND efet w=43660 l=8880
+ ad=0 pd=0 as=1.02511e+09 ps=216080 
M2260 GND diff_2702480_1629480# diff_2684720_1482960# GND efet w=48840 l=7400
+ ad=0 pd=0 as=1.18063e+09 ps=242720 
M2261 diff_2735040_1583600# diff_2727640_1580640# GND GND efet w=48840 l=7400
+ ad=9.39682e+08 pd=224960 as=0 ps=0 
M2262 diff_2684720_1561400# diff_2677320_1556960# GND GND efet w=43660 l=8140
+ ad=5.01602e+08 pd=115440 as=0 ps=0 
M2263 GND diff_2752800_1629480# diff_2735040_1456320# GND efet w=43660 l=8880
+ ad=0 pd=0 as=1.0032e+09 ps=213120 
M2264 GND diff_2803120_1629480# diff_2786840_1482960# GND efet w=48840 l=7400
+ ad=0 pd=0 as=1.11929e+09 ps=236800 
M2265 diff_2835680_1583600# diff_2828280_1580640# GND GND efet w=48840 l=7400
+ ad=1.22224e+09 pd=307840 as=0 ps=0 
M2266 diff_2785360_1561400# diff_2777960_1556960# GND GND efet w=43660 l=8140
+ ad=5.01602e+08 pd=115440 as=0 ps=0 
M2267 diff_602360_1574720# diff_321160_969400# GND GND efet w=56980 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2268 diff_606800_1443000# Vdd Vdd GND efet w=7400 l=19240
+ ad=0 pd=0 as=0 ps=0 
M2269 diff_627520_1602840# Vdd Vdd GND efet w=7400 l=17760
+ ad=0 pd=0 as=0 ps=0 
M2270 Vdd Vdd Vdd GND efet w=2960 l=2960
+ ad=0 pd=0 as=0 ps=0 
M2271 Vdd Vdd Vdd GND efet w=1480 l=2960
+ ad=0 pd=0 as=0 ps=0 
M2272 diff_794760_1574720# cl GND GND efet w=44400 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2273 GND cl diff_794760_1574720# GND efet w=44400 l=10360
+ ad=0 pd=0 as=0 ps=0 
M2274 diff_794760_1574720# diff_321160_969400# GND GND efet w=59940 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2275 diff_797720_1443000# Vdd Vdd GND efet w=7400 l=19240
+ ad=0 pd=0 as=0 ps=0 
M2276 diff_821400_1602840# Vdd Vdd GND efet w=7400 l=17760
+ ad=0 pd=0 as=0 ps=0 
M2277 Vdd Vdd Vdd GND efet w=1480 l=1480
+ ad=0 pd=0 as=0 ps=0 
M2278 Vdd Vdd Vdd GND efet w=1480 l=1480
+ ad=0 pd=0 as=0 ps=0 
M2279 diff_985680_1574720# cl GND GND efet w=44400 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2280 GND cl diff_985680_1574720# GND efet w=44400 l=10360
+ ad=0 pd=0 as=0 ps=0 
M2281 diff_985680_1574720# diff_321160_969400# GND GND efet w=59940 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2282 diff_1232840_1500720# diff_1293520_1043400# diff_1274280_1562880# GND efet w=38480 l=8880
+ ad=-1.20431e+09 pd=592000 as=0 ps=0 
M2283 diff_1329040_1488880# diff_1293520_1043400# diff_1376400_1561400# GND efet w=37000 l=7400
+ ad=-1.72344e+09 pd=503200 as=0 ps=0 
M2284 diff_1429680_1488880# diff_1293520_1043400# diff_1477040_1561400# GND efet w=37000 l=7400
+ ad=-1.62268e+09 pd=565360 as=0 ps=0 
M2285 diff_1528840_1490360# diff_1293520_1043400# diff_1577680_1561400# GND efet w=37000 l=7400
+ ad=-1.83077e+09 pd=497280 as=0 ps=0 
M2286 diff_1629480_1490360# diff_1293520_1043400# diff_1678320_1561400# GND efet w=37000 l=7400
+ ad=-1.56135e+09 pd=577200 as=0 ps=0 
M2287 diff_1731600_1487400# diff_1293520_1043400# diff_1778960_1561400# GND efet w=37000 l=7400
+ ad=-1.64239e+09 pd=509120 as=0 ps=0 
M2288 diff_1832240_1487400# diff_1293520_1043400# diff_1879600_1561400# GND efet w=37000 l=7400
+ ad=-1.46935e+09 pd=580160 as=0 ps=0 
M2289 diff_1932880_1487400# diff_1293520_1043400# diff_1980240_1561400# GND efet w=37000 l=7400
+ ad=-1.64239e+09 pd=509120 as=0 ps=0 
M2290 diff_2033520_1487400# diff_1293520_1043400# diff_2080880_1561400# GND efet w=37000 l=7400
+ ad=-1.5263e+09 pd=571280 as=0 ps=0 
M2291 diff_2135640_1488880# diff_1293520_1043400# diff_2181520_1561400# GND efet w=37000 l=7400
+ ad=-1.71906e+09 pd=503200 as=0 ps=0 
M2292 diff_2236280_1488880# diff_1293520_1043400# diff_2282160_1561400# GND efet w=37000 l=7400
+ ad=-1.55697e+09 pd=568320 as=0 ps=0 
M2293 diff_2335440_1488880# diff_1293520_1043400# diff_2382800_1561400# GND efet w=37000 l=7400
+ ad=-1.72782e+09 pd=503200 as=0 ps=0 
M2294 diff_2436080_1488880# diff_1293520_1043400# diff_2483440_1561400# GND efet w=37000 l=7400
+ ad=-1.55697e+09 pd=571280 as=0 ps=0 
M2295 diff_2536720_1488880# diff_1293520_1043400# diff_2584080_1561400# GND efet w=37000 l=7400
+ ad=-1.72782e+09 pd=503200 as=0 ps=0 
M2296 diff_2637360_1488880# diff_1293520_1043400# diff_2684720_1561400# GND efet w=37000 l=7400
+ ad=-1.52192e+09 pd=574240 as=0 ps=0 
M2297 diff_2739480_1487400# diff_1293520_1043400# diff_2785360_1561400# GND efet w=37000 l=7400
+ ad=-1.58763e+09 pd=523920 as=0 ps=0 
M2298 diff_1238760_1688680# diff_2998480_1207680# diff_2920040_1736040# GND efet w=97680 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2299 diff_3005880_2094200# diff_3023640_1207680# diff_2920040_1736040# GND efet w=190920 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2300 diff_2920040_1842600# diff_3045840_1124800# diff_3005880_2094200# GND efet w=190920 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2301 diff_1232840_1500720# diff_1226920_1511080# diff_1229880_1524400# GND efet w=50320 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2302 diff_988640_1443000# Vdd Vdd GND efet w=7400 l=19240
+ ad=0 pd=0 as=0 ps=0 
M2303 diff_1012320_1602840# Vdd Vdd GND efet w=7400 l=17760
+ ad=0 pd=0 as=0 ps=0 
M2304 diff_1628000_1583600# diff_1226920_1511080# diff_1629480_1490360# GND efet w=42180 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2305 diff_1527360_1583600# diff_1226920_1511080# diff_1528840_1490360# GND efet w=38480 l=8140
+ ad=0 pd=0 as=0 ps=0 
M2306 diff_1728640_1583600# diff_1226920_1511080# diff_1731600_1487400# GND efet w=38480 l=8140
+ ad=0 pd=0 as=0 ps=0 
M2307 diff_1829280_1583600# diff_1226920_1511080# diff_1832240_1487400# GND efet w=39960 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2308 diff_1929920_1583600# diff_1226920_1511080# diff_1932880_1487400# GND efet w=38480 l=8140
+ ad=0 pd=0 as=0 ps=0 
M2309 diff_1326080_1583600# diff_1226920_1511080# diff_1329040_1488880# GND efet w=37740 l=8140
+ ad=0 pd=0 as=0 ps=0 
M2310 diff_1426720_1583600# diff_1226920_1511080# diff_1429680_1488880# GND efet w=38480 l=8140
+ ad=0 pd=0 as=0 ps=0 
M2311 diff_2030560_1583600# diff_1226920_1511080# diff_2033520_1487400# GND efet w=38480 l=8140
+ ad=0 pd=0 as=0 ps=0 
M2312 diff_2332480_1583600# diff_1226920_1511080# diff_2335440_1488880# GND efet w=37740 l=8140
+ ad=0 pd=0 as=0 ps=0 
M2313 diff_2433120_1583600# diff_1226920_1511080# diff_2436080_1488880# GND efet w=38480 l=8140
+ ad=0 pd=0 as=0 ps=0 
M2314 diff_2533760_1583600# diff_1226920_1511080# diff_2536720_1488880# GND efet w=37740 l=8140
+ ad=0 pd=0 as=0 ps=0 
M2315 diff_2634400_1583600# diff_1226920_1511080# diff_2637360_1488880# GND efet w=38480 l=8140
+ ad=0 pd=0 as=0 ps=0 
M2316 Vdd Vdd Vdd GND efet w=1480 l=1480
+ ad=0 pd=0 as=0 ps=0 
M2317 Vdd Vdd Vdd GND efet w=1480 l=1480
+ ad=0 pd=0 as=0 ps=0 
M2318 diff_1278720_1482960# diff_1274280_1133680# diff_1232840_1500720# GND efet w=35520 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2319 diff_1376400_1481480# diff_1274280_1133680# diff_1329040_1488880# GND efet w=42180 l=8140
+ ad=0 pd=0 as=0 ps=0 
M2320 diff_1477040_1482960# diff_1274280_1133680# diff_1429680_1488880# GND efet w=41440 l=10360
+ ad=0 pd=0 as=0 ps=0 
M2321 diff_1576200_1482960# diff_1274280_1133680# diff_1528840_1490360# GND efet w=41440 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2322 diff_1676840_1481480# diff_1274280_1133680# diff_1629480_1490360# GND efet w=42920 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2323 diff_1778960_1482960# diff_1274280_1133680# diff_1731600_1487400# GND efet w=41440 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2324 diff_1879600_1482960# diff_1274280_1133680# diff_1832240_1487400# GND efet w=42180 l=10360
+ ad=0 pd=0 as=0 ps=0 
M2325 diff_2131200_1583600# diff_1226920_1511080# diff_2135640_1488880# GND efet w=37000 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2326 diff_2231840_1583600# diff_1226920_1511080# diff_2236280_1488880# GND efet w=37740 l=8140
+ ad=0 pd=0 as=0 ps=0 
M2327 diff_1980240_1482960# diff_1274280_1133680# diff_1932880_1487400# GND efet w=41440 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2328 diff_2080880_1482960# diff_1274280_1133680# diff_2033520_1487400# GND efet w=41440 l=10360
+ ad=0 pd=0 as=0 ps=0 
M2329 diff_2183000_1482960# diff_1274280_1133680# diff_2135640_1488880# GND efet w=40700 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2330 diff_2283640_1482960# diff_1274280_1133680# diff_2236280_1488880# GND efet w=40700 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2331 diff_2382800_1482960# diff_1274280_1133680# diff_2335440_1488880# GND efet w=41440 l=10360
+ ad=0 pd=0 as=0 ps=0 
M2332 diff_2483440_1482960# diff_1274280_1133680# diff_2436080_1488880# GND efet w=41440 l=10360
+ ad=0 pd=0 as=0 ps=0 
M2333 diff_2735040_1583600# diff_1226920_1511080# diff_2739480_1487400# GND efet w=35520 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2334 diff_2584080_1482960# diff_1274280_1133680# diff_2536720_1488880# GND efet w=41440 l=10360
+ ad=0 pd=0 as=0 ps=0 
M2335 diff_2684720_1482960# diff_1274280_1133680# diff_2637360_1488880# GND efet w=41440 l=10360
+ ad=0 pd=0 as=0 ps=0 
M2336 diff_2786840_1482960# diff_1274280_1133680# diff_2739480_1487400# GND efet w=39220 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2337 GND diff_414400_1443000# diff_415880_1340880# GND efet w=69560 l=7400
+ ad=0 pd=0 as=1.69537e+09 ps=319680 
M2338 GND diff_606800_1443000# diff_608280_1340880# GND efet w=69560 l=7400
+ ad=0 pd=0 as=1.69975e+09 ps=313760 
M2339 Vdd Vdd diff_415880_1340880# GND efet w=8880 l=16280
+ ad=0 pd=0 as=0 ps=0 
M2340 GND diff_797720_1443000# diff_799200_1340880# GND efet w=69560 l=7400
+ ad=0 pd=0 as=1.7808e+09 ps=319680 
M2341 diff_415880_1340880# diff_415880_1340880# diff_415880_1340880# GND efet w=2220 l=2220
+ ad=0 pd=0 as=0 ps=0 
M2342 diff_415880_1340880# diff_415880_1340880# diff_415880_1340880# GND efet w=4440 l=4440
+ ad=0 pd=0 as=0 ps=0 
M2343 Vdd Vdd diff_608280_1340880# GND efet w=8880 l=13320
+ ad=0 pd=0 as=0 ps=0 
M2344 GND diff_988640_1443000# diff_990120_1340880# GND efet w=69560 l=7400
+ ad=0 pd=0 as=1.78299e+09 ps=328560 
M2345 diff_608280_1340880# diff_608280_1340880# diff_608280_1340880# GND efet w=4440 l=5180
+ ad=0 pd=0 as=0 ps=0 
M2346 Vdd Vdd diff_799200_1340880# GND efet w=8880 l=13320
+ ad=0 pd=0 as=0 ps=0 
M2347 diff_1324600_1456320# diff_1311280_1160320# diff_1232840_1500720# GND efet w=38480 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2348 diff_1425240_1456320# diff_1311280_1160320# diff_1329040_1488880# GND efet w=38480 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2349 diff_1524400_1456320# diff_1311280_1160320# diff_1429680_1488880# GND efet w=38480 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2350 diff_1625040_1456320# diff_1311280_1160320# diff_1528840_1490360# GND efet w=38480 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2351 diff_1727160_1456320# diff_1311280_1160320# diff_1629480_1490360# GND efet w=38480 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2352 diff_1827800_1456320# diff_1311280_1160320# diff_1731600_1487400# GND efet w=38480 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2353 diff_1928440_1456320# diff_1311280_1160320# diff_1832240_1487400# GND efet w=38480 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2354 diff_2029080_1456320# diff_1311280_1160320# diff_1932880_1487400# GND efet w=38480 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2355 diff_2131200_1456320# diff_1311280_1160320# diff_2033520_1487400# GND efet w=38480 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2356 diff_2231840_1456320# diff_1311280_1160320# diff_2135640_1488880# GND efet w=38480 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2357 diff_2331000_1456320# diff_1311280_1160320# diff_2236280_1488880# GND efet w=38480 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2358 diff_2431640_1456320# diff_1311280_1160320# diff_2335440_1488880# GND efet w=38480 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2359 diff_2532280_1456320# diff_1311280_1160320# diff_2436080_1488880# GND efet w=38480 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2360 diff_2632920_1456320# diff_1311280_1160320# diff_2536720_1488880# GND efet w=38480 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2361 diff_2735040_1456320# diff_1311280_1160320# diff_2637360_1488880# GND efet w=37000 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2362 diff_2835680_1583600# diff_1311280_1160320# diff_2739480_1487400# GND efet w=56980 l=8140
+ ad=0 pd=0 as=0 ps=0 
M2363 diff_799200_1340880# diff_799200_1340880# diff_799200_1340880# GND efet w=5920 l=5920
+ ad=0 pd=0 as=0 ps=0 
M2364 diff_990120_1340880# diff_990120_1340880# diff_990120_1340880# GND efet w=2960 l=2960
+ ad=0 pd=0 as=0 ps=0 
M2365 Vdd Vdd diff_990120_1340880# GND efet w=8880 l=13320
+ ad=0 pd=0 as=0 ps=0 
M2366 diff_990120_1340880# diff_990120_1340880# diff_990120_1340880# GND efet w=5180 l=5180
+ ad=0 pd=0 as=0 ps=0 
M2367 diff_1232840_1500720# diff_1247640_1422280# diff_1253560_1194360# GND efet w=50320 l=8880
+ ad=0 pd=0 as=1.09342e+09 ps=852480 
M2368 diff_1329040_1488880# diff_1386760_1422280# diff_1253560_1194360# GND efet w=50320 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2369 diff_1528840_1490360# diff_1386760_1422280# diff_1456320_1215080# GND efet w=50320 l=7400
+ ad=0 pd=0 as=7.62666e+08 ps=808080 
M2370 diff_1731600_1487400# diff_1386760_1422280# diff_1656120_1383800# GND efet w=50320 l=7400
+ ad=0 pd=0 as=1.37379e+09 ps=864320 
M2371 diff_1932880_1487400# diff_1386760_1422280# diff_1858880_1213600# GND efet w=50320 l=7400
+ ad=0 pd=0 as=1.43512e+09 ps=855440 
M2372 diff_2135640_1488880# diff_1386760_1422280# diff_2060160_1213600# GND efet w=50320 l=7400
+ ad=0 pd=0 as=9.66374e+08 ps=814000 
M2373 diff_2335440_1488880# diff_1386760_1422280# diff_2262920_1213600# GND efet w=50320 l=7400
+ ad=0 pd=0 as=8.54663e+08 ps=784400 
M2374 diff_2536720_1488880# diff_1386760_1422280# diff_2462720_1213600# GND efet w=50320 l=7400
+ ad=0 pd=0 as=1.41322e+09 ps=882080 
M2375 diff_2739480_1487400# diff_1386760_1422280# diff_2664000_1215080# GND efet w=42920 l=7400
+ ad=0 pd=0 as=2.10686e+08 ps=710400 
M2376 Vdd diff_415880_1340880# io3 GND efet w=217560 l=8880
+ ad=0 pd=0 as=-1.92592e+09 ps=2.39168e+06 
M2377 d3 GND d3 GND efet w=218300 l=138380
+ ad=0 pd=0 as=0 ps=0 
M2378 GND diff_414400_1443000# io3 GND efet w=222740 l=10360
+ ad=0 pd=0 as=0 ps=0 
M2379 Vdd diff_608280_1340880# io2 GND efet w=219040 l=8880
+ ad=0 pd=0 as=1.61555e+09 ps=2.37688e+06 
M2380 io2 GND io2 GND efet w=216820 l=132460
+ ad=0 pd=0 as=0 ps=0 
M2381 GND diff_606800_1443000# io2 GND efet w=222740 l=10360
+ ad=0 pd=0 as=0 ps=0 
M2382 Vdd diff_799200_1340880# io1 GND efet w=219040 l=8880
+ ad=0 pd=0 as=1.09642e+09 ps=2.28512e+06 
M2383 GND diff_797720_1443000# io1 GND efet w=222740 l=10360
+ ad=0 pd=0 as=0 ps=0 
M2384 Vdd diff_990120_1340880# io0 GND efet w=217560 l=8880
+ ad=0 pd=0 as=1.58926e+09 ps=2.38872e+06 
M2385 diff_612720_1192880# diff_501720_853960# diff_503200_1786360# GND efet w=28120 l=8880
+ ad=1.36024e+09 pd=284160 as=1.90346e+09 ps=402560 
M2386 diff_670440_1255040# diff_550560_1112960# diff_612720_1192880# GND efet w=28120 l=8880
+ ad=1.65813e+09 pd=301920 as=0 ps=0 
M2387 diff_799200_1192880# diff_501720_853960# diff_694120_1786360# GND efet w=28120 l=8880
+ ad=1.461e+09 pd=296000 as=1.53109e+09 ps=322640 
M2388 diff_842120_1275760# diff_550560_1112960# diff_799200_1192880# GND efet w=28120 l=8880
+ ad=1.55956e+09 pd=266400 as=0 ps=0 
M2389 io1 GND io1 GND efet w=206460 l=154660
+ ad=0 pd=0 as=0 ps=0 
M2390 io3 GND io3 GND efet w=184260 l=86580
+ ad=0 pd=0 as=0 ps=0 
M2391 diff_612720_1192880# diff_507640_1070040# io3 GND efet w=26640 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2392 GND diff_988640_1443000# io0 GND efet w=222740 l=10360
+ ad=0 pd=0 as=0 ps=0 
M2393 diff_1429680_1488880# diff_1247640_1422280# diff_1456320_1215080# GND efet w=48840 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2394 diff_1629480_1490360# diff_1247640_1422280# diff_1656120_1383800# GND efet w=50320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2395 diff_1832240_1487400# diff_1247640_1422280# diff_1858880_1213600# GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2396 diff_2033520_1487400# diff_1247640_1422280# diff_2060160_1213600# GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2397 diff_2236280_1488880# diff_1247640_1422280# diff_2262920_1213600# GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2398 diff_2436080_1488880# diff_1247640_1422280# diff_2462720_1213600# GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2399 diff_2637360_1488880# diff_1247640_1422280# diff_2664000_1215080# GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2400 diff_1111480_1194360# diff_501720_853960# diff_1077440_1786360# GND efet w=26640 l=8880
+ ad=-1.96e+09 pd=497280 as=4.29318e+08 ps=85840 
M2401 diff_1192880_1336440# diff_550560_1112960# diff_1111480_1194360# GND efet w=26640 l=8880
+ ad=1.10177e+09 pd=198320 as=0 ps=0 
M2402 diff_990120_1192880# diff_501720_853960# diff_886520_1786360# GND efet w=28120 l=8880
+ ad=1.57709e+09 pd=325600 as=1.34929e+09 ps=287120 
M2403 diff_1022680_1281680# diff_550560_1112960# diff_990120_1192880# GND efet w=28120 l=8880
+ ad=-1.80886e+09 pd=423280 as=0 ps=0 
M2404 io0 GND io0 GND efet w=219040 l=159840
+ ad=0 pd=0 as=0 ps=0 
M2405 io3 GND io3 GND efet w=34780 l=42180
+ ad=0 pd=0 as=0 ps=0 
M2406 GND diff_507640_1070040# diff_550560_1112960# GND efet w=20720 l=8880
+ ad=0 pd=0 as=1.9845e+09 ps=526880 
M2407 diff_609760_1096680# io3 GND GND efet w=42920 l=8880
+ ad=1.27043e+09 pd=224960 as=0 ps=0 
M2408 GND io3 diff_609760_1096680# GND efet w=42920 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2409 diff_799200_1192880# diff_507640_1070040# io2 GND efet w=28120 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2410 diff_1456320_1215080# diff_695600_586080# diff_1232840_1340880# GND efet w=28120 l=7400
+ ad=0 pd=0 as=-1.8921e+09 ps=408480 
M2411 diff_1192880_1336440# diff_1232840_1340880# GND GND efet w=62160 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2412 diff_1232840_1340880# diff_1232840_1340880# diff_1232840_1340880# GND efet w=1480 l=1480
+ ad=0 pd=0 as=0 ps=0 
M2413 diff_1192880_1336440# Vdd Vdd GND efet w=11840 l=31080
+ ad=0 pd=0 as=0 ps=0 
M2414 diff_1232840_1340880# diff_1232840_1340880# diff_1232840_1340880# GND efet w=1480 l=2960
+ ad=0 pd=0 as=0 ps=0 
M2415 diff_1858880_1213600# diff_695600_586080# diff_1657600_1243200# GND efet w=29600 l=7400
+ ad=0 pd=0 as=-2.01695e+09 ps=390720 
M2416 diff_2262920_1213600# diff_695600_586080# diff_2060160_1243200# GND efet w=26640 l=7400
+ ad=0 pd=0 as=-1.53725e+09 ps=411440 
M2417 Vdd Vdd Vdd GND efet w=2960 l=3700
+ ad=0 pd=0 as=0 ps=0 
M2418 Vdd Vdd Vdd GND efet w=2960 l=3700
+ ad=0 pd=0 as=0 ps=0 
M2419 diff_550560_1112960# diff_550560_1112960# diff_550560_1112960# GND efet w=2960 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2420 Vdd Vdd Vdd GND efet w=1480 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2421 Vdd Vdd diff_1456320_1215080# GND efet w=8140 l=79920
+ ad=0 pd=0 as=0 ps=0 
M2422 Vdd Vdd diff_1253560_1194360# GND efet w=7400 l=81400
+ ad=0 pd=0 as=0 ps=0 
M2423 Vdd Vdd Vdd GND efet w=1480 l=6660
+ ad=0 pd=0 as=0 ps=0 
M2424 diff_1657600_1243200# diff_1657600_1243200# diff_1657600_1243200# GND efet w=3700 l=3700
+ ad=0 pd=0 as=0 ps=0 
M2425 diff_1657600_1243200# diff_1657600_1243200# diff_1657600_1243200# GND efet w=1480 l=2960
+ ad=0 pd=0 as=0 ps=0 
M2426 diff_1858880_1213600# Vdd Vdd GND efet w=7400 l=79920
+ ad=0 pd=0 as=0 ps=0 
M2427 Vdd Vdd diff_1022680_1281680# GND efet w=10360 l=29600
+ ad=0 pd=0 as=0 ps=0 
M2428 Vdd Vdd Vdd GND efet w=1480 l=5920
+ ad=0 pd=0 as=0 ps=0 
M2429 Vdd Vdd diff_1656120_1383800# GND efet w=7400 l=79920
+ ad=0 pd=0 as=0 ps=0 
M2430 Vdd Vdd Vdd GND efet w=2960 l=5920
+ ad=0 pd=0 as=0 ps=0 
M2431 diff_1022680_1281680# diff_1657600_1243200# GND GND efet w=51800 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2432 diff_2060160_1213600# Vdd Vdd GND efet w=8140 l=83620
+ ad=0 pd=0 as=0 ps=0 
M2433 Vdd Vdd diff_842120_1275760# GND efet w=10360 l=48840
+ ad=0 pd=0 as=0 ps=0 
M2434 diff_2664000_1215080# diff_695600_586080# diff_2462720_1243200# GND efet w=29600 l=8880
+ ad=0 pd=0 as=-1.64677e+09 ps=396640 
M2435 diff_2262920_1213600# Vdd Vdd GND efet w=6660 l=82140
+ ad=0 pd=0 as=0 ps=0 
M2436 diff_842120_1275760# diff_2060160_1243200# GND GND efet w=62160 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2437 Vdd Vdd Vdd GND efet w=1480 l=3700
+ ad=0 pd=0 as=0 ps=0 
M2438 diff_1657600_1243200# diff_769600_586080# diff_1656120_1383800# GND efet w=28120 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2439 diff_2462720_1213600# Vdd Vdd GND efet w=9620 l=83620
+ ad=0 pd=0 as=0 ps=0 
M2440 diff_2060160_1243200# diff_769600_586080# diff_2060160_1213600# GND efet w=29600 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2441 diff_2462720_1243200# diff_769600_586080# diff_2462720_1213600# GND efet w=29600 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2442 Vdd Vdd diff_670440_1255040# GND efet w=10360 l=31080
+ ad=0 pd=0 as=0 ps=0 
M2443 diff_2664000_1215080# Vdd Vdd GND efet w=8880 l=87320
+ ad=0 pd=0 as=0 ps=0 
M2444 diff_670440_1255040# diff_2462720_1243200# GND GND efet w=50320 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2445 Vdd Vdd diff_550560_1112960# GND efet w=8880 l=54760
+ ad=0 pd=0 as=0 ps=0 
M2446 diff_550560_1112960# diff_550560_1112960# diff_550560_1112960# GND efet w=2220 l=8140
+ ad=0 pd=0 as=0 ps=0 
M2447 diff_1232840_1340880# diff_769600_586080# diff_1253560_1194360# GND efet w=28120 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2448 io3 Vdd Vdd GND efet w=10360 l=14800
+ ad=0 pd=0 as=0 ps=0 
M2449 diff_700040_1055240# diff_700040_1055240# diff_700040_1055240# GND efet w=2220 l=4440
+ ad=3.04466e+08 pd=94720 as=0 ps=0 
M2450 diff_507640_1070040# diff_507640_1070040# diff_507640_1070040# GND efet w=740 l=2220
+ ad=-1.46278e+09 pd=674880 as=0 ps=0 
M2451 diff_507640_1070040# diff_507640_1070040# diff_507640_1070040# GND efet w=740 l=1480
+ ad=0 pd=0 as=0 ps=0 
M2452 diff_700040_1055240# diff_700040_1055240# diff_700040_1055240# GND efet w=2220 l=6660
+ ad=0 pd=0 as=0 ps=0 
M2453 diff_507640_1070040# diff_507640_1070040# diff_507640_1070040# GND efet w=1480 l=4440
+ ad=0 pd=0 as=0 ps=0 
M2454 diff_797720_1095200# io2 GND GND efet w=42920 l=8880
+ ad=1.28357e+09 pd=227920 as=0 ps=0 
M2455 GND io2 diff_797720_1095200# GND efet w=42920 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2456 diff_990120_1192880# diff_507640_1070040# io1 GND efet w=28120 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2457 diff_1111480_1194360# diff_507640_1070040# io0 GND efet w=28120 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2458 io2 Vdd Vdd GND efet w=10360 l=14800
+ ad=0 pd=0 as=0 ps=0 
M2459 diff_700040_1055240# Vdd Vdd GND efet w=8880 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2460 diff_507640_1070040# clk1 diff_507640_1052280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=4.4027e+08 ps=136160 
M2461 diff_507640_1052280# diff_507640_1052280# diff_507640_1052280# GND efet w=2220 l=5180
+ ad=0 pd=0 as=0 ps=0 
M2462 GND diff_507640_1052280# diff_550560_1112960# GND efet w=45140 l=8140
+ ad=0 pd=0 as=0 ps=0 
M2463 Vdd Vdd diff_609760_1096680# GND efet w=8880 l=26640
+ ad=0 pd=0 as=0 ps=0 
M2464 diff_507640_1052280# diff_507640_1052280# diff_507640_1052280# GND efet w=2220 l=2960
+ ad=0 pd=0 as=0 ps=0 
M2465 Vdd Vdd Vdd GND efet w=1480 l=4440
+ ad=0 pd=0 as=0 ps=0 
M2466 Vdd diff_700040_1055240# diff_507640_1070040# GND efet w=11100 l=26640
+ ad=0 pd=0 as=0 ps=0 
M2467 Vdd Vdd diff_593480_988640# GND efet w=8880 l=17760
+ ad=0 pd=0 as=1.25072e+09 ps=272320 
M2468 diff_507640_1070040# diff_700040_1055240# diff_507640_1070040# GND efet w=57720 l=3700
+ ad=0 pd=0 as=0 ps=0 
M2469 diff_988640_1095200# io1 GND GND efet w=42920 l=8880
+ ad=1.27043e+09 pd=224960 as=0 ps=0 
M2470 GND io1 diff_988640_1095200# GND efet w=42920 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2471 diff_1456320_1215080# diff_1250600_1186960# diff_1429680_1120360# GND efet w=48840 l=8880
+ ad=0 pd=0 as=-1.71906e+09 ps=559440 
M2472 diff_1656120_1383800# diff_1250600_1186960# diff_1629480_1115920# GND efet w=48100 l=8140
+ ad=0 pd=0 as=-1.6862e+09 ps=568320 
M2473 diff_2664000_1215080# diff_1250600_1186960# diff_2637360_1120360# GND efet w=50320 l=8880
+ ad=0 pd=0 as=-1.68839e+09 ps=565360 
M2474 diff_1858880_1213600# diff_1250600_1186960# diff_1832240_1118880# GND efet w=48840 l=7400
+ ad=0 pd=0 as=-1.57449e+09 ps=571280 
M2475 diff_2060160_1213600# diff_1250600_1186960# diff_2033520_1120360# GND efet w=48840 l=7400
+ ad=0 pd=0 as=-1.62268e+09 ps=565360 
M2476 diff_1253560_1194360# diff_1250600_1186960# diff_1232840_1105560# GND efet w=50320 l=8880
+ ad=0 pd=0 as=-1.31164e+09 ps=583120 
M2477 diff_1253560_1194360# diff_1386760_1188440# diff_1329040_1118880# GND efet w=50320 l=7400
+ ad=0 pd=0 as=-1.81762e+09 ps=497280 
M2478 diff_1456320_1215080# diff_1386760_1188440# diff_1528840_1118880# GND efet w=50320 l=7400
+ ad=0 pd=0 as=-1.92495e+09 ps=491360 
M2479 diff_1656120_1383800# diff_1386760_1188440# diff_1731600_1118880# GND efet w=50320 l=7400
+ ad=0 pd=0 as=-1.73658e+09 ps=503200 
M2480 diff_1858880_1213600# diff_1386760_1188440# diff_1932880_1118880# GND efet w=50320 l=7400
+ ad=0 pd=0 as=-1.73658e+09 ps=503200 
M2481 diff_2262920_1213600# diff_1250600_1186960# diff_2236280_1120360# GND efet w=48840 l=7400
+ ad=0 pd=0 as=-1.65334e+09 ps=562400 
M2482 diff_2060160_1213600# diff_1386760_1188440# diff_2135640_1118880# GND efet w=50320 l=7400
+ ad=0 pd=0 as=-1.81324e+09 ps=497280 
M2483 diff_2462720_1213600# diff_1250600_1186960# diff_2436080_1120360# GND efet w=48840 l=7400
+ ad=0 pd=0 as=-1.66211e+09 ps=562400 
M2484 diff_2262920_1213600# diff_1386760_1188440# diff_2335440_1118880# GND efet w=50320 l=7400
+ ad=0 pd=0 as=-1.82201e+09 ps=497280 
M2485 diff_2462720_1213600# diff_1386760_1188440# diff_2536720_1118880# GND efet w=50320 l=7400
+ ad=0 pd=0 as=-1.82201e+09 ps=497280 
M2486 diff_2664000_1215080# diff_1386760_1188440# diff_2739480_1118880# GND efet w=42920 l=5920
+ ad=0 pd=0 as=-1.70153e+09 ps=515040 
M2487 diff_2835680_1022680# diff_1311280_1160320# diff_2739480_1118880# GND efet w=54020 l=8140
+ ad=1.30767e+09 pd=307840 as=0 ps=0 
M2488 diff_1232840_1105560# diff_1311280_1160320# diff_1324600_1144040# GND efet w=38480 l=7400
+ ad=0 pd=0 as=1.07549e+09 ps=219040 
M2489 diff_1329040_1118880# diff_1311280_1160320# diff_1425240_1144040# GND efet w=38480 l=7400
+ ad=0 pd=0 as=1.08425e+09 ps=219040 
M2490 diff_1429680_1120360# diff_1311280_1160320# diff_1524400_1142560# GND efet w=38480 l=7400
+ ad=0 pd=0 as=1.13244e+09 ps=222000 
M2491 diff_1528840_1118880# diff_1311280_1160320# diff_1625040_1142560# GND efet w=38480 l=7400
+ ad=0 pd=0 as=1.1412e+09 ps=222000 
M2492 diff_1629480_1115920# diff_1311280_1160320# diff_1727160_1145520# GND efet w=38480 l=7400
+ ad=0 pd=0 as=1.01854e+09 ps=216080 
M2493 diff_1731600_1118880# diff_1311280_1160320# diff_1827800_1145520# GND efet w=38480 l=7400
+ ad=0 pd=0 as=1.0273e+09 ps=216080 
M2494 diff_1832240_1118880# diff_1311280_1160320# diff_1928440_1145520# GND efet w=38480 l=7400
+ ad=0 pd=0 as=1.01854e+09 ps=216080 
M2495 diff_1932880_1118880# diff_1311280_1160320# diff_2029080_1145520# GND efet w=38480 l=7400
+ ad=0 pd=0 as=1.0273e+09 ps=216080 
M2496 diff_2033520_1120360# diff_1311280_1160320# diff_2131200_1144040# GND efet w=38480 l=7400
+ ad=0 pd=0 as=1.07549e+09 ps=219040 
M2497 diff_2135640_1118880# diff_1311280_1160320# diff_2231840_1144040# GND efet w=38480 l=7400
+ ad=0 pd=0 as=1.08425e+09 ps=219040 
M2498 diff_2236280_1120360# diff_1311280_1160320# diff_2331000_1144040# GND efet w=38480 l=7400
+ ad=0 pd=0 as=1.07549e+09 ps=219040 
M2499 diff_2335440_1118880# diff_1311280_1160320# diff_2431640_1144040# GND efet w=38480 l=7400
+ ad=0 pd=0 as=1.08425e+09 ps=219040 
M2500 diff_2436080_1120360# diff_1311280_1160320# diff_2532280_1144040# GND efet w=38480 l=7400
+ ad=0 pd=0 as=1.07549e+09 ps=219040 
M2501 diff_2536720_1118880# diff_1311280_1160320# diff_2632920_1144040# GND efet w=38480 l=7400
+ ad=0 pd=0 as=1.08425e+09 ps=219040 
M2502 diff_2637360_1120360# diff_1311280_1160320# diff_2735040_1144040# GND efet w=37000 l=7400
+ ad=0 pd=0 as=1.06015e+09 ps=216080 
M2503 io1 Vdd Vdd GND efet w=10360 l=14800
+ ad=0 pd=0 as=0 ps=0 
M2504 diff_1108520_1095200# io0 GND GND efet w=42920 l=8880
+ ad=1.28357e+09 pd=227920 as=0 ps=0 
M2505 GND io0 diff_1108520_1095200# GND efet w=42920 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2506 io0 Vdd Vdd GND efet w=10360 l=14800
+ ad=0 pd=0 as=0 ps=0 
M2507 Vdd Vdd diff_797720_1095200# GND efet w=8880 l=28120
+ ad=0 pd=0 as=0 ps=0 
M2508 Vdd Vdd diff_988640_1095200# GND efet w=8880 l=26640
+ ad=0 pd=0 as=0 ps=0 
M2509 Vdd Vdd diff_1108520_1095200# GND efet w=8880 l=25160
+ ad=0 pd=0 as=0 ps=0 
M2510 GND diff_612720_984200# diff_593480_988640# GND efet w=75480 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2511 diff_593480_988640# diff_501720_853960# diff_552040_951640# GND efet w=14800 l=8880
+ ad=0 pd=0 as=2.54086e+08 ps=65120 
M2512 diff_1329040_1118880# diff_1274280_1133680# diff_1376400_1118880# GND efet w=42180 l=8140
+ ad=0 pd=0 as=1.20253e+09 ps=245680 
M2513 diff_1429680_1120360# diff_1274280_1133680# diff_1477040_1118880# GND efet w=41440 l=10360
+ ad=0 pd=0 as=1.22881e+09 ps=245680 
M2514 diff_1629480_1115920# diff_1274280_1133680# diff_1676840_1117400# GND efet w=42920 l=7400
+ ad=0 pd=0 as=1.28796e+09 ps=251600 
M2515 diff_1528840_1118880# diff_1274280_1133680# diff_1576200_1117400# GND efet w=41440 l=9620
+ ad=0 pd=0 as=1.25729e+09 ps=245680 
M2516 diff_1731600_1118880# diff_1274280_1133680# diff_1778960_1120360# GND efet w=41440 l=9620
+ ad=0 pd=0 as=1.14339e+09 ps=239760 
M2517 diff_1832240_1118880# diff_1274280_1133680# diff_1879600_1120360# GND efet w=42180 l=10360
+ ad=0 pd=0 as=1.17186e+09 ps=242720 
M2518 diff_1932880_1118880# diff_1274280_1133680# diff_1980240_1120360# GND efet w=41440 l=9620
+ ad=0 pd=0 as=1.14339e+09 ps=239760 
M2519 diff_2033520_1120360# diff_1274280_1133680# diff_2080880_1120360# GND efet w=41440 l=10360
+ ad=0 pd=0 as=1.17186e+09 ps=242720 
M2520 diff_2135640_1118880# diff_1274280_1133680# diff_2183000_1118880# GND efet w=40700 l=9620
+ ad=0 pd=0 as=1.20034e+09 ps=242720 
M2521 diff_2335440_1118880# diff_1274280_1133680# diff_2382800_1118880# GND efet w=41440 l=10360
+ ad=0 pd=0 as=1.20034e+09 ps=242720 
M2522 diff_2236280_1120360# diff_1274280_1133680# diff_2283640_1118880# GND efet w=40700 l=9620
+ ad=0 pd=0 as=1.22881e+09 ps=245680 
M2523 diff_2436080_1120360# diff_1274280_1133680# diff_2483440_1118880# GND efet w=41440 l=10360
+ ad=0 pd=0 as=1.22881e+09 ps=245680 
M2524 diff_2536720_1118880# diff_1274280_1133680# diff_2584080_1118880# GND efet w=41440 l=10360
+ ad=0 pd=0 as=1.20034e+09 ps=242720 
M2525 diff_2637360_1120360# diff_1274280_1133680# diff_2684720_1118880# GND efet w=41440 l=10360
+ ad=0 pd=0 as=1.22881e+09 ps=245680 
M2526 diff_2739480_1118880# diff_1274280_1133680# diff_2786840_1118880# GND efet w=39960 l=10360
+ ad=0 pd=0 as=1.1631e+09 ps=239760 
M2527 diff_507640_1070040# diff_507640_1070040# diff_507640_1070040# GND efet w=1480 l=1480
+ ad=0 pd=0 as=0 ps=0 
M2528 diff_1232840_1105560# diff_1274280_1133680# diff_1278720_1114440# GND efet w=35520 l=7400
+ ad=0 pd=0 as=1.19158e+09 ps=239760 
M2529 diff_1329040_1118880# diff_1226920_1511080# diff_1326080_1019720# GND efet w=37740 l=8140
+ ad=0 pd=0 as=1.02073e+09 ps=233840 
M2530 diff_1429680_1120360# diff_1226920_1511080# diff_1426720_1022680# GND efet w=38480 l=8140
+ ad=0 pd=0 as=1.05139e+09 ps=233840 
M2531 diff_1629480_1115920# diff_1226920_1511080# diff_1628000_1022680# GND efet w=42180 l=7400
+ ad=0 pd=0 as=1.09082e+09 ps=236800 
M2532 diff_1528840_1118880# diff_1226920_1511080# diff_1527360_1022680# GND efet w=38480 l=8140
+ ad=0 pd=0 as=1.04263e+09 ps=233840 
M2533 diff_1731600_1118880# diff_1226920_1511080# diff_1728640_1022680# GND efet w=38480 l=8140
+ ad=0 pd=0 as=9.52824e+08 ps=230880 
M2534 diff_1832240_1118880# diff_1226920_1511080# diff_1829280_1022680# GND efet w=39960 l=7400
+ ad=0 pd=0 as=9.90061e+08 ps=230880 
M2535 diff_1932880_1118880# diff_1226920_1511080# diff_1929920_1022680# GND efet w=38480 l=8140
+ ad=0 pd=0 as=9.52824e+08 ps=230880 
M2536 diff_2033520_1120360# diff_1226920_1511080# diff_2030560_1022680# GND efet w=38480 l=8140
+ ad=0 pd=0 as=9.96632e+08 ps=230880 
M2537 diff_2135640_1118880# diff_1226920_1511080# diff_2131200_1022680# GND efet w=37000 l=7400
+ ad=0 pd=0 as=1.01416e+09 ps=233840 
M2538 diff_2236280_1120360# diff_1226920_1511080# diff_2231840_1022680# GND efet w=37740 l=8140
+ ad=0 pd=0 as=1.05577e+09 ps=233840 
M2539 diff_2335440_1118880# diff_1226920_1511080# diff_2332480_1022680# GND efet w=37740 l=8140
+ ad=0 pd=0 as=1.01196e+09 ps=233840 
M2540 diff_2436080_1120360# diff_1226920_1511080# diff_2433120_1022680# GND efet w=38480 l=8140
+ ad=0 pd=0 as=1.05139e+09 ps=233840 
M2541 diff_2536720_1118880# diff_1226920_1511080# diff_2533760_1022680# GND efet w=37740 l=8140
+ ad=0 pd=0 as=1.01196e+09 ps=233840 
M2542 diff_2637360_1120360# diff_1226920_1511080# diff_2634400_1022680# GND efet w=38480 l=8140
+ ad=0 pd=0 as=1.05139e+09 ps=233840 
M2543 diff_2739480_1118880# diff_1226920_1511080# diff_2735040_1022680# GND efet w=35520 l=7400
+ ad=0 pd=0 as=9.8349e+08 ps=227920 
M2544 diff_1232840_1105560# diff_1226920_1511080# diff_1229880_1031560# GND efet w=47360 l=5920
+ ad=0 pd=0 as=1.277e+09 ps=239760 
M2545 diff_1274280_1049320# diff_1263920_1047840# GND GND efet w=57720 l=8880
+ ad=5.54171e+08 pd=130240 as=0 ps=0 
M2546 diff_507640_1070040# diff_507640_1070040# diff_507640_1070040# GND efet w=740 l=2220
+ ad=0 pd=0 as=0 ps=0 
M2547 GND diff_552040_951640# diff_233840_991600# GND efet w=112480 l=8880
+ ad=0 pd=0 as=-4.50408e+08 ps=1.45632e+06 
M2548 diff_233840_991600# diff_519480_898360# Vdd GND efet w=102860 l=8140
+ ad=0 pd=0 as=0 ps=0 
M2549 diff_688200_944240# diff_504680_587560# diff_661560_957560# GND efet w=44400 l=8880
+ ad=1.31424e+09 pd=281200 as=1.28576e+09 ps=272320 
M2550 diff_661560_957560# diff_418840_657120# diff_612720_984200# GND efet w=48840 l=8880
+ ad=0 pd=0 as=9.15587e+08 ps=186480 
M2551 GND diff_1243200_956080# diff_1229880_1031560# GND efet w=35520 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2552 diff_1232840_1105560# diff_1293520_1043400# diff_1274280_1049320# GND efet w=38480 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2553 GND diff_1343840_956080# diff_1324600_1144040# GND efet w=43660 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2554 diff_1376400_1047840# diff_1369000_956080# GND GND efet w=44400 l=8880
+ ad=5.05982e+08 pd=115440 as=0 ps=0 
M2555 diff_1329040_1118880# diff_1293520_1043400# diff_1376400_1047840# GND efet w=37000 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2556 GND diff_1444480_956080# diff_1425240_1144040# GND efet w=43660 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2557 diff_1477040_1047840# diff_1469640_956080# GND GND efet w=44400 l=8880
+ ad=5.05982e+08 pd=115440 as=0 ps=0 
M2558 diff_1429680_1120360# diff_1293520_1043400# diff_1477040_1047840# GND efet w=37000 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2559 GND diff_1545120_956080# diff_1524400_1142560# GND efet w=43660 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2560 diff_1577680_1047840# diff_1570280_956080# GND GND efet w=44400 l=8880
+ ad=5.05982e+08 pd=115440 as=0 ps=0 
M2561 diff_1528840_1118880# diff_1293520_1043400# diff_1577680_1047840# GND efet w=37000 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2562 GND diff_1645760_956080# diff_1625040_1142560# GND efet w=43660 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2563 diff_1678320_1047840# diff_1670920_956080# GND GND efet w=44400 l=8880
+ ad=5.05982e+08 pd=115440 as=0 ps=0 
M2564 diff_1629480_1115920# diff_1293520_1043400# diff_1678320_1047840# GND efet w=37000 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2565 GND diff_1746400_956080# diff_1727160_1145520# GND efet w=43660 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2566 diff_1778960_1047840# diff_1771560_956080# GND GND efet w=44400 l=8880
+ ad=5.05982e+08 pd=115440 as=0 ps=0 
M2567 diff_1731600_1118880# diff_1293520_1043400# diff_1778960_1047840# GND efet w=37000 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2568 GND diff_1847040_956080# diff_1827800_1145520# GND efet w=43660 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2569 diff_1879600_1047840# diff_1872200_956080# GND GND efet w=44400 l=8880
+ ad=5.05982e+08 pd=115440 as=0 ps=0 
M2570 diff_1832240_1118880# diff_1293520_1043400# diff_1879600_1047840# GND efet w=37000 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2571 GND diff_1947680_956080# diff_1928440_1145520# GND efet w=43660 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2572 diff_1980240_1047840# diff_1972840_956080# GND GND efet w=44400 l=8880
+ ad=5.05982e+08 pd=115440 as=0 ps=0 
M2573 diff_1932880_1118880# diff_1293520_1043400# diff_1980240_1047840# GND efet w=37000 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2574 GND diff_2048320_956080# diff_2029080_1145520# GND efet w=43660 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2575 diff_2080880_1047840# diff_2073480_956080# GND GND efet w=44400 l=8880
+ ad=5.05982e+08 pd=115440 as=0 ps=0 
M2576 diff_2033520_1120360# diff_1293520_1043400# diff_2080880_1047840# GND efet w=37000 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2577 GND diff_2148960_956080# diff_2131200_1144040# GND efet w=43660 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2578 diff_2181520_1047840# diff_2174120_956080# GND GND efet w=44400 l=8880
+ ad=5.05982e+08 pd=115440 as=0 ps=0 
M2579 diff_2135640_1118880# diff_1293520_1043400# diff_2181520_1047840# GND efet w=37000 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2580 GND diff_2249600_956080# diff_2231840_1144040# GND efet w=43660 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2581 diff_2282160_1047840# diff_2274760_956080# GND GND efet w=44400 l=8880
+ ad=5.05982e+08 pd=115440 as=0 ps=0 
M2582 diff_2236280_1120360# diff_1293520_1043400# diff_2282160_1047840# GND efet w=37000 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2583 GND diff_2350240_956080# diff_2331000_1144040# GND efet w=43660 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2584 diff_2382800_1047840# diff_2375400_956080# GND GND efet w=44400 l=8880
+ ad=5.05982e+08 pd=115440 as=0 ps=0 
M2585 diff_2335440_1118880# diff_1293520_1043400# diff_2382800_1047840# GND efet w=37000 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2586 GND diff_2450880_956080# diff_2431640_1144040# GND efet w=43660 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2587 diff_2483440_1047840# diff_2476040_956080# GND GND efet w=44400 l=8880
+ ad=5.05982e+08 pd=115440 as=0 ps=0 
M2588 diff_2436080_1120360# diff_1293520_1043400# diff_2483440_1047840# GND efet w=37000 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2589 GND diff_2551520_956080# diff_2532280_1144040# GND efet w=43660 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2590 diff_2584080_1047840# diff_2576680_956080# GND GND efet w=44400 l=8880
+ ad=5.05982e+08 pd=115440 as=0 ps=0 
M2591 diff_2536720_1118880# diff_1293520_1043400# diff_2584080_1047840# GND efet w=37000 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2592 GND diff_2652160_956080# diff_2632920_1144040# GND efet w=43660 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2593 diff_2684720_1047840# diff_2677320_956080# GND GND efet w=44400 l=8880
+ ad=5.05982e+08 pd=115440 as=0 ps=0 
M2594 diff_2637360_1120360# diff_1293520_1043400# diff_2684720_1047840# GND efet w=37000 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2595 GND diff_2752800_956080# diff_2735040_1144040# GND efet w=43660 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2596 diff_2785360_1047840# diff_2777960_956080# GND GND efet w=44400 l=8880
+ ad=5.05982e+08 pd=115440 as=0 ps=0 
M2597 diff_2739480_1118880# diff_1293520_1043400# diff_2785360_1047840# GND efet w=37000 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2598 diff_3196800_1889960# Vdd Vdd GND efet w=16280 l=8880
+ ad=2.38754e+08 pd=71040 as=0 ps=0 
M2599 diff_3196800_1889960# diff_3196800_1889960# diff_3196800_1889960# GND efet w=2220 l=6660
+ ad=0 pd=0 as=0 ps=0 
M2600 diff_3196800_1889960# diff_3196800_1889960# diff_3196800_1889960# GND efet w=2220 l=2220
+ ad=0 pd=0 as=0 ps=0 
M2601 Vdd Vdd Vdd GND efet w=740 l=2220
+ ad=0 pd=0 as=0 ps=0 
M2602 GND diff_3412880_1952120# diff_3267840_1873680# GND efet w=99160 l=7400
+ ad=0 pd=0 as=1.99107e+09 ps=310800 
M2603 Vdd Vdd diff_3267840_1873680# GND efet w=10360 l=20720
+ ad=0 pd=0 as=0 ps=0 
M2604 Vdd Vdd Vdd GND efet w=740 l=1480
+ ad=0 pd=0 as=0 ps=0 
M2605 GND d2 diff_3469120_1237280# GND efet w=241240 l=7400
+ ad=0 pd=0 as=-1.18679e+09 ps=488400 
M2606 diff_3469120_1237280# Vdd Vdd GND efet w=10360 l=20720
+ ad=0 pd=0 as=0 ps=0 
M2607 diff_3267840_1873680# clk1 diff_3414360_1900320# GND efet w=16280 l=7400
+ ad=0 pd=0 as=2.56277e+08 ps=68080 
M2608 Vdd Vdd diff_3469120_1398600# GND efet w=10360 l=20720
+ ad=0 pd=0 as=1.66251e+09 ps=281200 
M2609 diff_3414360_1900320# diff_3414360_1900320# diff_3414360_1900320# GND efet w=2220 l=2220
+ ad=0 pd=0 as=0 ps=0 
M2610 GND diff_3414360_1900320# diff_3343320_1672400# GND efet w=54760 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2611 Vdd Vdd diff_3343320_1672400# GND efet w=11840 l=23680
+ ad=0 pd=0 as=0 ps=0 
M2612 Vdd Vdd Vdd GND efet w=2960 l=5920
+ ad=0 pd=0 as=0 ps=0 
M2613 Vdd Vdd Vdd GND efet w=2960 l=3700
+ ad=0 pd=0 as=0 ps=0 
M2614 diff_3343320_1672400# clk2 diff_3414360_1847040# GND efet w=14800 l=7400
+ ad=0 pd=0 as=2.10278e+08 ps=59200 
M2615 diff_1237280_2100120# diff_3193840_1805600# Vdd GND efet w=19240 l=7400
+ ad=1.59283e+09 pd=911680 as=0 ps=0 
M2616 GND diff_3267840_1761200# diff_1237280_2100120# GND efet w=365560 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2617 diff_1237280_2100120# diff_3193840_1805600# diff_1237280_2100120# GND efet w=50320 l=5920
+ ad=0 pd=0 as=0 ps=0 
M2618 diff_3193840_1805600# Vdd Vdd GND efet w=14800 l=7400
+ ad=2.65038e+08 pd=74000 as=0 ps=0 
M2619 diff_3193840_1805600# diff_3193840_1805600# diff_3193840_1805600# GND efet w=1480 l=5920
+ ad=0 pd=0 as=0 ps=0 
M2620 diff_3193840_1805600# diff_3193840_1805600# diff_3193840_1805600# GND efet w=2220 l=2220
+ ad=0 pd=0 as=0 ps=0 
M2621 diff_3414360_1847040# diff_3414360_1847040# diff_3414360_1847040# GND efet w=1480 l=2960
+ ad=0 pd=0 as=0 ps=0 
M2622 GND diff_3414360_1847040# diff_3285600_1753800# GND efet w=54760 l=8880
+ ad=0 pd=0 as=-1.90962e+09 ps=414400 
M2623 Vdd Vdd diff_3285600_1753800# GND efet w=10360 l=22200
+ ad=0 pd=0 as=0 ps=0 
M2624 Vdd Vdd Vdd GND efet w=740 l=2220
+ ad=0 pd=0 as=0 ps=0 
M2625 GND diff_3469120_1237280# diff_3469120_1398600# GND efet w=54760 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2626 diff_3285600_1753800# clk1 diff_3412880_1796720# GND efet w=17760 l=7400
+ ad=0 pd=0 as=2.54086e+08 ps=65120 
M2627 GND diff_3412880_1796720# diff_3358120_1041920# GND efet w=54760 l=7400
+ ad=0 pd=0 as=1.72823e+09 ps=278240 
M2628 Vdd Vdd diff_3358120_1041920# GND efet w=10360 l=20720
+ ad=0 pd=0 as=0 ps=0 
M2629 Vdd Vdd Vdd GND efet w=1480 l=1480
+ ad=0 pd=0 as=0 ps=0 
M2630 Vdd Vdd Vdd GND efet w=1480 l=2220
+ ad=0 pd=0 as=0 ps=0 
M2631 GND diff_3285600_1753800# diff_3239720_1740480# GND efet w=16280 l=7400
+ ad=0 pd=0 as=7.33784e+08 ps=171680 
M2632 diff_3239720_1740480# Vdd Vdd GND efet w=8880 l=44400
+ ad=0 pd=0 as=0 ps=0 
M2633 diff_3213080_1693120# Vdd Vdd GND efet w=8880 l=22200
+ ad=1.08863e+09 pd=216080 as=0 ps=0 
M2634 diff_3340360_1716800# diff_3285600_1753800# diff_3208640_1687200# GND efet w=19240 l=7400
+ ad=4.31509e+08 pd=109520 as=7.84163e+08 ps=168720 
M2635 diff_3213080_1693120# diff_3208640_1687200# GND GND efet w=75480 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2636 diff_3208640_1687200# diff_3208640_1687200# diff_3208640_1687200# GND efet w=3700 l=3700
+ ad=0 pd=0 as=0 ps=0 
M2637 diff_3208640_1687200# diff_3208640_1687200# diff_3208640_1687200# GND efet w=2220 l=2220
+ ad=0 pd=0 as=0 ps=0 
M2638 diff_3340360_1716800# diff_3223440_2120840# diff_3343320_1672400# GND efet w=16280 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2639 diff_3208640_1687200# diff_3239720_1740480# GND GND efet w=14800 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2640 diff_3377360_1571760# diff_3343320_1672400# diff_3115400_1533280# GND efet w=25160 l=7400
+ ad=8.65208e+08 pd=168720 as=4.42461e+08 ps=85840 
M2641 diff_3421760_1613200# clk2 diff_3377360_1571760# GND efet w=25160 l=7400
+ ad=1.50919e+09 pd=201280 as=0 ps=0 
M2642 GND diff_3167200_1580640# diff_1386760_1422280# GND efet w=173160 l=7400
+ ad=0 pd=0 as=-1.32259e+09 ps=488400 
M2643 diff_3377360_1571760# diff_3358120_1041920# diff_3167200_1580640# GND efet w=23680 l=7400
+ ad=0 pd=0 as=3.8113e+08 ps=79920 
M2644 GND diff_507640_1070040# diff_661560_957560# GND efet w=33300 l=9620
+ ad=0 pd=0 as=0 ps=0 
M2645 diff_688200_944240# diff_695600_586080# GND GND efet w=45880 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2646 GND diff_769600_586080# diff_688200_944240# GND efet w=44400 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2647 diff_1018240_964960# d3 GND GND efet w=45140 l=8140
+ ad=1.34929e+09 pd=260480 as=0 ps=0 
M2648 GND diff_864320_837680# diff_858400_964960# GND efet w=26640 l=8880
+ ad=0 pd=0 as=5.21315e+08 ps=100640 
M2649 GND diff_858400_964960# diff_190920_1013800# GND efet w=20720 l=8880
+ ad=0 pd=0 as=-7.509e+08 ps=908720 
M2650 diff_1006400_970880# clk2 diff_864320_837680# GND efet w=13320 l=8880
+ ad=1.57709e+08 pd=50320 as=5.21315e+08 ps=136160 
M2651 Vdd diff_1018240_964960# diff_1006400_970880# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2652 diff_1018240_964960# Vdd Vdd GND efet w=8880 l=41440
+ ad=0 pd=0 as=0 ps=0 
M2653 GND diff_856920_686720# diff_1018240_964960# GND efet w=22200 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2654 GND diff_1133680_519480# diff_1018240_964960# GND efet w=22200 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2655 GND diff_1293520_956080# diff_1278720_1114440# GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2656 diff_1326080_1019720# diff_1318680_956080# GND GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2657 GND diff_1394160_956080# diff_1376400_1118880# GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2658 diff_1426720_1022680# diff_1419320_956080# GND GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2659 GND diff_1494800_956080# diff_1477040_1118880# GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2660 diff_1527360_1022680# diff_1519960_956080# GND GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2661 GND diff_1595440_956080# diff_1576200_1117400# GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2662 diff_1628000_1022680# diff_1620600_956080# GND GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2663 GND diff_1696080_956080# diff_1676840_1117400# GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2664 diff_1728640_1022680# diff_1721240_956080# GND GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2665 GND diff_1796720_956080# diff_1778960_1120360# GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2666 diff_1829280_1022680# diff_1821880_956080# GND GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2667 GND diff_1897360_956080# diff_1879600_1120360# GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2668 diff_1929920_1022680# diff_1922520_956080# GND GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2669 GND diff_1998000_956080# diff_1980240_1120360# GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2670 diff_2030560_1022680# diff_2023160_956080# GND GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2671 GND diff_2098640_956080# diff_2080880_1120360# GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2672 diff_2131200_1022680# diff_2123800_956080# GND GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2673 GND diff_2199280_956080# diff_2183000_1118880# GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2674 diff_2231840_1022680# diff_2224440_956080# GND GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2675 GND diff_2299920_956080# diff_2283640_1118880# GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2676 diff_2332480_1022680# diff_2325080_956080# GND GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2677 GND diff_2400560_956080# diff_2382800_1118880# GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2678 diff_2433120_1022680# diff_2425720_956080# GND GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2679 GND diff_2501200_956080# diff_2483440_1118880# GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2680 diff_2533760_1022680# diff_2526360_956080# GND GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2681 GND diff_2601840_956080# diff_2584080_1118880# GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2682 diff_2634400_1022680# diff_2627000_956080# GND GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2683 GND diff_2702480_956080# diff_2684720_1118880# GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2684 diff_2735040_1022680# diff_2727640_956080# GND GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2685 GND diff_2803120_956080# diff_2786840_1118880# GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2686 diff_2835680_1022680# diff_2828280_956080# GND GND efet w=48840 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2687 GND diff_593480_988640# diff_614200_882080# GND efet w=59940 l=8140
+ ad=0 pd=0 as=5.93598e+08 ps=153920 
M2688 diff_614200_882080# diff_501720_853960# diff_519480_898360# GND efet w=13320 l=7400
+ ad=0 pd=0 as=4.75317e+08 ps=124320 
M2689 diff_614200_882080# Vdd Vdd GND efet w=8880 l=19240
+ ad=0 pd=0 as=0 ps=0 
M2690 Vdd Vdd Vdd GND efet w=1480 l=5920
+ ad=0 pd=0 as=0 ps=0 
M2691 Vdd Vdd Vdd GND efet w=2220 l=5920
+ ad=0 pd=0 as=0 ps=0 
M2692 Vdd Vdd diff_612720_984200# GND efet w=8880 l=82880
+ ad=0 pd=0 as=0 ps=0 
M2693 Vdd Vdd Vdd GND efet w=2220 l=4440
+ ad=0 pd=0 as=0 ps=0 
M2694 Vdd Vdd Vdd GND efet w=2220 l=6660
+ ad=0 pd=0 as=0 ps=0 
M2695 diff_321160_969400# Vdd Vdd GND efet w=11840 l=22200
+ ad=1.44785e+09 pd=263440 as=0 ps=0 
M2696 diff_501720_853960# diff_592000_757760# Vdd GND efet w=10360 l=10360
+ ad=1.49604e+09 pd=296000 as=0 ps=0 
M2697 diff_501720_853960# diff_592000_757760# diff_501720_853960# GND efet w=56980 l=28860
+ ad=0 pd=0 as=0 ps=0 
M2698 diff_592000_757760# Vdd Vdd GND efet w=10360 l=8880
+ ad=2.738e+08 pd=71040 as=0 ps=0 
M2699 Vdd Vdd diff_418840_657120# GND efet w=10360 l=22200
+ ad=0 pd=0 as=2.11593e+09 ps=361120 
M2700 diff_321160_969400# diff_418840_657120# GND GND efet w=106560 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2701 GND clk2 diff_501720_853960# GND efet w=56240 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2702 Vdd Vdd Vdd GND efet w=3700 l=4440
+ ad=0 pd=0 as=0 ps=0 
M2703 reset GND reset GND efet w=224960 l=139120
+ ad=1.14818e+09 pd=1.07744e+06 as=0 ps=0 
M2704 diff_418840_657120# reset GND GND efet w=178340 l=8140
+ ad=0 pd=0 as=0 ps=0 
M2705 Vdd Vdd Vdd GND efet w=2220 l=2960
+ ad=0 pd=0 as=0 ps=0 
M2706 sync clk2 diff_350760_574240# GND efet w=14800 l=8880
+ ad=0 pd=0 as=2.7599e+08 ps=74000 
M2707 diff_350760_574240# diff_350760_574240# diff_350760_574240# GND efet w=2960 l=5180
+ ad=0 pd=0 as=0 ps=0 
M2708 diff_350760_574240# diff_350760_574240# diff_350760_574240# GND efet w=1480 l=5920
+ ad=0 pd=0 as=0 ps=0 
M2709 GND diff_350760_574240# diff_356680_563880# GND efet w=49580 l=8140
+ ad=0 pd=0 as=1.69537e+09 ps=364080 
M2710 Vdd Vdd Vdd GND efet w=740 l=2220
+ ad=0 pd=0 as=0 ps=0 
M2711 Vdd Vdd diff_504680_587560# GND efet w=11100 l=43660
+ ad=0 pd=0 as=5.71694e+08 ps=124320 
M2712 Vdd Vdd diff_605320_617160# GND efet w=10360 l=79920
+ ad=0 pd=0 as=6.37406e+08 ps=121360 
M2713 diff_190920_1013800# diff_856920_939800# GND GND efet w=20720 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2714 diff_190920_1013800# Vdd Vdd GND efet w=8880 l=41440
+ ad=0 pd=0 as=0 ps=0 
M2715 Vdd Vdd Vdd GND efet w=1480 l=4440
+ ad=0 pd=0 as=0 ps=0 
M2716 Vdd Vdd Vdd GND efet w=1480 l=2960
+ ad=0 pd=0 as=0 ps=0 
M2717 diff_858400_964960# Vdd Vdd GND efet w=8880 l=62160
+ ad=0 pd=0 as=0 ps=0 
M2718 diff_864320_837680# diff_417360_463240# GND GND efet w=14800 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2719 diff_864320_837680# diff_864320_837680# diff_864320_837680# GND efet w=2220 l=2220
+ ad=0 pd=0 as=0 ps=0 
M2720 diff_864320_837680# diff_864320_837680# diff_864320_837680# GND efet w=740 l=2220
+ ad=0 pd=0 as=0 ps=0 
M2721 diff_1115920_948680# Vdd Vdd GND efet w=8880 l=63640
+ ad=8.89302e+08 pd=216080 as=0 ps=0 
M2722 GND d3 diff_1115920_948680# GND efet w=35520 l=8140
+ ad=0 pd=0 as=0 ps=0 
M2723 diff_1243200_956080# diff_1238760_948680# diff_1243200_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2724 diff_1263920_1047840# diff_1238760_948680# diff_1268360_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2725 diff_1293520_956080# diff_1238760_948680# diff_1293520_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2726 diff_1318680_956080# diff_1238760_948680# diff_1318680_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2727 diff_1343840_956080# diff_1238760_948680# diff_1343840_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2728 diff_1369000_956080# diff_1238760_948680# diff_1369000_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2729 diff_1394160_956080# diff_1238760_948680# diff_1394160_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2730 diff_1419320_956080# diff_1238760_948680# diff_1419320_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2731 diff_1444480_956080# diff_1238760_948680# diff_1444480_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2732 diff_1469640_956080# diff_1238760_948680# diff_1469640_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2733 diff_1494800_956080# diff_1238760_948680# diff_1494800_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2734 diff_1519960_956080# diff_1238760_948680# diff_1519960_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2735 diff_1545120_956080# diff_1238760_948680# diff_1545120_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2736 diff_1570280_956080# diff_1238760_948680# diff_1570280_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2737 diff_1595440_956080# diff_1238760_948680# diff_1595440_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2738 diff_1620600_956080# diff_1238760_948680# diff_1620600_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2739 diff_1645760_956080# diff_1238760_948680# diff_1645760_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2740 diff_1670920_956080# diff_1238760_948680# diff_1670920_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2741 diff_1696080_956080# diff_1238760_948680# diff_1696080_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2742 diff_1721240_956080# diff_1238760_948680# diff_1721240_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2743 diff_1746400_956080# diff_1238760_948680# diff_1746400_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2744 diff_1771560_956080# diff_1238760_948680# diff_1771560_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2745 diff_1796720_956080# diff_1238760_948680# diff_1796720_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2746 diff_1821880_956080# diff_1238760_948680# diff_1821880_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2747 diff_1847040_956080# diff_1238760_948680# diff_1847040_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2748 diff_1872200_956080# diff_1238760_948680# diff_1872200_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2749 diff_1897360_956080# diff_1238760_948680# diff_1897360_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2750 diff_1922520_956080# diff_1238760_948680# diff_1922520_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2751 diff_1947680_956080# diff_1238760_948680# diff_1947680_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2752 diff_1972840_956080# diff_1238760_948680# diff_1972840_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2753 diff_1998000_956080# diff_1238760_948680# diff_1998000_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2754 diff_2023160_956080# diff_1238760_948680# diff_2023160_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2755 diff_2048320_956080# diff_1238760_948680# diff_2048320_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2756 diff_2073480_956080# diff_1238760_948680# diff_2073480_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2757 diff_2098640_956080# diff_1238760_948680# diff_2098640_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2758 diff_2123800_956080# diff_1238760_948680# diff_2123800_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2759 diff_2148960_956080# diff_1238760_948680# diff_2148960_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2760 diff_2174120_956080# diff_1238760_948680# diff_2174120_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2761 diff_2199280_956080# diff_1238760_948680# diff_2199280_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2762 diff_2224440_956080# diff_1238760_948680# diff_2224440_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2763 diff_2249600_956080# diff_1238760_948680# diff_2249600_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2764 diff_2274760_956080# diff_1238760_948680# diff_2274760_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2765 diff_2299920_956080# diff_1238760_948680# diff_2299920_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2766 diff_2325080_956080# diff_1238760_948680# diff_2325080_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2767 diff_2350240_956080# diff_1238760_948680# diff_2350240_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2768 diff_2375400_956080# diff_1238760_948680# diff_2375400_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2769 diff_2400560_956080# diff_1238760_948680# diff_2400560_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2770 diff_2425720_956080# diff_1238760_948680# diff_2425720_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2771 diff_2450880_956080# diff_1238760_948680# diff_2450880_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2772 diff_2476040_956080# diff_1238760_948680# diff_2476040_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2773 diff_2501200_956080# diff_1238760_948680# diff_2501200_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2774 diff_2526360_956080# diff_1238760_948680# diff_2526360_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2775 diff_2551520_956080# diff_1238760_948680# diff_2551520_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2776 diff_2576680_956080# diff_1238760_948680# diff_2576680_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2777 diff_2601840_956080# diff_1238760_948680# diff_2601840_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2778 diff_2627000_956080# diff_1238760_948680# diff_2627000_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2779 diff_2652160_956080# diff_1238760_948680# diff_2652160_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2780 diff_2677320_956080# diff_1238760_948680# diff_2677320_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2781 diff_2702480_956080# diff_1238760_948680# diff_2702480_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2782 diff_2727640_956080# diff_1238760_948680# diff_2727640_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2783 diff_2752800_956080# diff_1238760_948680# diff_2752800_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2784 diff_2777960_956080# diff_1238760_948680# diff_2777960_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2785 diff_2803120_956080# diff_1238760_948680# diff_2803120_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2786 diff_2828280_956080# diff_1238760_948680# diff_2828280_927960# GND efet w=13320 l=8880
+ ad=1.73042e+08 pd=53280 as=2.56277e+08 ps=65120 
M2787 GND diff_3115400_1533280# diff_2998480_1207680# GND efet w=150960 l=7400
+ ad=0 pd=0 as=-1.71249e+09 ps=408480 
M2788 Vdd Vdd diff_1386760_1422280# GND efet w=8880 l=17760
+ ad=0 pd=0 as=0 ps=0 
M2789 Vdd Vdd diff_2998480_1207680# GND efet w=8880 l=17760
+ ad=0 pd=0 as=0 ps=0 
M2790 diff_3377360_1515520# diff_3358120_1041920# diff_3121320_1481480# GND efet w=23680 l=7400
+ ad=8.93683e+08 pd=171680 as=4.16176e+08 ps=82880 
M2791 Vdd Vdd diff_1386760_1188440# GND efet w=8880 l=17760
+ ad=0 pd=0 as=-1.5942e+09 ps=396640 
M2792 diff_1386760_1188440# diff_3121320_1481480# GND GND efet w=150960 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2793 GND diff_3121320_1453360# diff_2912640_526880# GND efet w=150960 l=7400
+ ad=0 pd=0 as=-1.25031e+09 ps=408480 
M2794 Vdd Vdd diff_2912640_526880# GND efet w=8880 l=17760
+ ad=0 pd=0 as=0 ps=0 
M2795 Vdd Vdd diff_2940760_526880# GND efet w=8880 l=17760
+ ad=0 pd=0 as=-1.26783e+09 ps=402560 
M2796 diff_3421760_1613200# Vdd Vdd GND efet w=10360 l=41440
+ ad=0 pd=0 as=0 ps=0 
M2797 diff_3476520_1593960# diff_3469120_1398600# diff_3421760_1613200# GND efet w=44400 l=7400
+ ad=5.25696e+08 pd=112480 as=0 ps=0 
M2798 GND diff_3488360_1570280# diff_3476520_1593960# GND efet w=44400 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2799 Vdd Vdd Vdd GND efet w=1480 l=2960
+ ad=0 pd=0 as=0 ps=0 
M2800 Vdd Vdd Vdd GND efet w=1480 l=2960
+ ad=0 pd=0 as=0 ps=0 
M2801 Vdd Vdd diff_3421760_1466680# GND efet w=10360 l=41440
+ ad=0 pd=0 as=1.79613e+09 ps=260480 
M2802 diff_3377360_1515520# diff_3343320_1672400# diff_3121320_1453360# GND efet w=26640 l=7400
+ ad=0 pd=0 as=5.08173e+08 ps=91760 
M2803 diff_3421760_1466680# clk2 diff_3377360_1515520# GND efet w=26640 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2804 diff_3504640_1514040# diff_3488360_1570280# diff_3421760_1466680# GND efet w=42920 l=7400
+ ad=5.08173e+08 pd=109520 as=0 ps=0 
M2805 GND diff_3469120_1237280# diff_3504640_1514040# GND efet w=42920 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2806 GND diff_3488360_1339400# diff_3476520_1401560# GND efet w=44400 l=7400
+ ad=0 pd=0 as=1.50261e+09 ps=245680 
M2807 diff_3377360_1374920# diff_3343320_1672400# diff_3121320_1397120# GND efet w=23680 l=7400
+ ad=8.60827e+08 pd=168720 as=4.16176e+08 ps=82880 
M2808 diff_3421760_1422280# clk2 diff_3377360_1374920# GND efet w=23680 l=7400
+ ad=1.36243e+09 pd=189440 as=0 ps=0 
M2809 diff_2940760_526880# diff_3121320_1397120# GND GND efet w=150960 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2810 GND diff_3122800_1370480# diff_1247640_1422280# GND efet w=150960 l=7400
+ ad=0 pd=0 as=-1.4343e+09 ps=399600 
M2811 diff_3377360_1374920# diff_3358120_1041920# diff_3122800_1370480# GND efet w=25160 l=7400
+ ad=0 pd=0 as=4.42461e+08 ps=85840 
M2812 Vdd Vdd diff_1247640_1422280# GND efet w=8880 l=17760
+ ad=0 pd=0 as=0 ps=0 
M2813 diff_3377360_1329040# diff_3358120_1041920# diff_3121320_1305360# GND efet w=23680 l=7400
+ ad=8.36733e+08 pd=165760 as=4.16176e+08 ps=82880 
M2814 Vdd Vdd diff_1250600_1186960# GND efet w=8880 l=17760
+ ad=0 pd=0 as=-1.3905e+09 ps=399600 
M2815 diff_1250600_1186960# diff_3121320_1305360# GND GND efet w=150960 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2816 GND diff_3121320_1277240# diff_2976280_1228400# GND efet w=150960 l=7400
+ ad=0 pd=0 as=-1.34012e+09 ps=399600 
M2817 Vdd Vdd diff_2976280_1228400# GND efet w=8880 l=17760
+ ad=0 pd=0 as=0 ps=0 
M2818 Vdd Vdd diff_3045840_1124800# GND efet w=8880 l=17760
+ ad=0 pd=0 as=-1.32698e+09 ps=402560 
M2819 diff_3045840_1124800# diff_3121320_1222480# GND GND efet w=150960 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2820 GND diff_3121320_1194360# diff_1274280_1133680# GND efet w=150960 l=7400
+ ad=0 pd=0 as=-1.47811e+09 ps=402560 
M2821 diff_3421760_1422280# Vdd Vdd GND efet w=8880 l=41440
+ ad=0 pd=0 as=0 ps=0 
M2822 diff_3476520_1401560# diff_3469120_1398600# diff_3421760_1422280# GND efet w=44400 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2823 diff_3534240_1386760# diff_3469120_1237280# diff_3421760_1283160# GND efet w=45880 l=7400
+ ad=6.11122e+08 pd=118400 as=1.80489e+09 ps=266400 
M2824 GND diff_3488360_1339400# diff_3534240_1386760# GND efet w=45880 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2825 Vdd Vdd Vdd GND efet w=2220 l=5180
+ ad=0 pd=0 as=0 ps=0 
M2826 Vdd Vdd Vdd GND efet w=2220 l=5180
+ ad=0 pd=0 as=0 ps=0 
M2827 Vdd Vdd diff_3421760_1283160# GND efet w=8880 l=41440
+ ad=0 pd=0 as=0 ps=0 
M2828 diff_3377360_1329040# diff_3343320_1672400# diff_3121320_1277240# GND efet w=23680 l=7400
+ ad=0 pd=0 as=4.16176e+08 ps=82880 
M2829 diff_3421760_1283160# clk2 diff_3377360_1329040# GND efet w=23680 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2830 diff_3377360_1189920# diff_3343320_1672400# diff_3121320_1222480# GND efet w=25160 l=7400
+ ad=8.89302e+08 pd=171680 as=4.42461e+08 ps=85840 
M2831 diff_3421760_1235800# clk2 diff_3377360_1189920# GND efet w=25160 l=7400
+ ad=1.80708e+09 pd=266400 as=0 ps=0 
M2832 d1 GND d1 GND efet w=219040 l=137640
+ ad=0 pd=0 as=0 ps=0 
M2833 GND diff_3488360_1339400# diff_3492800_1326080# GND efet w=78440 l=7400
+ ad=0 pd=0 as=9.2873e+08 ps=180560 
M2834 diff_3492800_1326080# diff_3469120_1237280# diff_3492800_1302400# GND efet w=78440 l=7400
+ ad=0 pd=0 as=-1.3664e+09 ps=432160 
M2835 diff_1133680_519480# diff_3469120_1237280# diff_3513520_1223960# GND efet w=57720 l=7400
+ ad=5.07863e+07 pd=740000 as=6.83405e+08 ps=139120 
M2836 diff_3377360_1189920# diff_3358120_1041920# diff_3121320_1194360# GND efet w=25160 l=7400
+ ad=0 pd=0 as=4.42461e+08 ps=85840 
M2837 Vdd Vdd diff_1274280_1133680# GND efet w=7400 l=17760
+ ad=0 pd=0 as=0 ps=0 
M2838 Vdd Vdd diff_1311280_1160320# GND efet w=7400 l=17760
+ ad=0 pd=0 as=-1.61173e+09 ps=399600 
M2839 diff_3377360_1142560# diff_3358120_1041920# diff_3119840_1129240# GND efet w=26640 l=7400
+ ad=9.13397e+08 pd=174640 as=4.68746e+08 ps=88800 
M2840 diff_1311280_1160320# diff_3119840_1129240# GND GND efet w=149480 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2841 GND diff_3119840_1102600# diff_3023640_1207680# GND efet w=149480 l=7400
+ ad=0 pd=0 as=-1.30945e+09 ps=399600 
M2842 Vdd Vdd diff_3023640_1207680# GND efet w=10360 l=17760
+ ad=0 pd=0 as=0 ps=0 
M2843 Vdd Vdd Vdd GND efet w=7400 l=5920
+ ad=0 pd=0 as=0 ps=0 
M2844 diff_1243200_927960# diff_1238760_920560# diff_1243200_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2845 diff_1268360_927960# diff_1238760_920560# diff_1268360_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2846 diff_1293520_927960# diff_1238760_920560# diff_1293520_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2847 diff_1318680_927960# diff_1238760_920560# diff_1318680_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2848 diff_1343840_927960# diff_1238760_920560# diff_1343840_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2849 diff_1369000_927960# diff_1238760_920560# diff_1369000_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2850 diff_1394160_927960# diff_1238760_920560# diff_1394160_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2851 diff_1419320_927960# diff_1238760_920560# diff_1419320_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2852 diff_1444480_927960# diff_1238760_920560# diff_1444480_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2853 diff_1469640_927960# diff_1238760_920560# diff_1469640_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2854 diff_1494800_927960# diff_1238760_920560# diff_1494800_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2855 diff_1519960_927960# diff_1238760_920560# diff_1519960_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2856 diff_1545120_927960# diff_1238760_920560# diff_1545120_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2857 diff_1570280_927960# diff_1238760_920560# diff_1570280_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2858 diff_1595440_927960# diff_1238760_920560# diff_1595440_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2859 diff_1620600_927960# diff_1238760_920560# diff_1620600_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2860 diff_1645760_927960# diff_1238760_920560# diff_1645760_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2861 diff_1670920_927960# diff_1238760_920560# diff_1670920_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2862 diff_1696080_927960# diff_1238760_920560# diff_1696080_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2863 diff_1721240_927960# diff_1238760_920560# diff_1721240_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2864 diff_1746400_927960# diff_1238760_920560# diff_1746400_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2865 diff_1771560_927960# diff_1238760_920560# diff_1771560_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2866 diff_1796720_927960# diff_1238760_920560# diff_1796720_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2867 diff_1821880_927960# diff_1238760_920560# diff_1821880_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2868 diff_1847040_927960# diff_1238760_920560# diff_1847040_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2869 diff_1872200_927960# diff_1238760_920560# diff_1872200_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2870 diff_1897360_927960# diff_1238760_920560# diff_1897360_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2871 diff_1922520_927960# diff_1238760_920560# diff_1922520_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2872 diff_1947680_927960# diff_1238760_920560# diff_1947680_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2873 diff_1972840_927960# diff_1238760_920560# diff_1972840_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2874 diff_1998000_927960# diff_1238760_920560# diff_1998000_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2875 diff_2023160_927960# diff_1238760_920560# diff_2023160_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2876 diff_2048320_927960# diff_1238760_920560# diff_2048320_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2877 diff_2073480_927960# diff_1238760_920560# diff_2073480_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2878 diff_2098640_927960# diff_1238760_920560# diff_2098640_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2879 diff_2123800_927960# diff_1238760_920560# diff_2123800_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2880 diff_2148960_927960# diff_1238760_920560# diff_2148960_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2881 diff_2174120_927960# diff_1238760_920560# diff_2174120_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2882 diff_2199280_927960# diff_1238760_920560# diff_2199280_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2883 diff_2224440_927960# diff_1238760_920560# diff_2224440_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2884 diff_2249600_927960# diff_1238760_920560# diff_2249600_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2885 diff_2274760_927960# diff_1238760_920560# diff_2274760_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2886 diff_2299920_927960# diff_1238760_920560# diff_2299920_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2887 diff_2325080_927960# diff_1238760_920560# diff_2325080_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2888 diff_2350240_927960# diff_1238760_920560# diff_2350240_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2889 diff_2375400_927960# diff_1238760_920560# diff_2375400_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2890 diff_2400560_927960# diff_1238760_920560# diff_2400560_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2891 diff_2425720_927960# diff_1238760_920560# diff_2425720_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2892 diff_2450880_927960# diff_1238760_920560# diff_2450880_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2893 diff_2476040_927960# diff_1238760_920560# diff_2476040_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2894 diff_2501200_927960# diff_1238760_920560# diff_2501200_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2895 diff_2526360_927960# diff_1238760_920560# diff_2526360_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2896 diff_2551520_927960# diff_1238760_920560# diff_2551520_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2897 diff_2576680_927960# diff_1238760_920560# diff_2576680_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2898 diff_2601840_927960# diff_1238760_920560# diff_2601840_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2899 diff_2627000_927960# diff_1238760_920560# diff_2627000_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2900 diff_2652160_927960# diff_1238760_920560# diff_2652160_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2901 diff_2677320_927960# diff_1238760_920560# diff_2677320_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2902 diff_2702480_927960# diff_1238760_920560# diff_2702480_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2903 diff_2727640_927960# diff_1238760_920560# diff_2727640_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2904 diff_2752800_927960# diff_1238760_920560# diff_2752800_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2905 diff_2777960_927960# diff_1238760_920560# diff_2777960_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2906 diff_2803120_927960# diff_1238760_920560# diff_2803120_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2907 diff_2828280_927960# diff_1238760_920560# diff_2828280_901320# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2908 diff_1238760_948680# Vdd Vdd GND efet w=7400 l=16280
+ ad=1.43033e+09 pd=322640 as=0 ps=0 
M2909 Vdd Vdd Vdd GND efet w=2960 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2910 Vdd Vdd Vdd GND efet w=1480 l=5920
+ ad=0 pd=0 as=0 ps=0 
M2911 diff_1068560_852480# Vdd Vdd GND efet w=8880 l=62160
+ ad=9.44062e+08 pd=183520 as=0 ps=0 
M2912 diff_507640_1070040# diff_1036000_463240# GND GND efet w=26640 l=7400
+ ad=0 pd=0 as=0 ps=0 
M2913 GND diff_1068560_852480# diff_507640_1070040# GND efet w=28120 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2914 diff_1243200_901320# diff_1238760_893920# diff_1243200_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2915 diff_1268360_901320# diff_1238760_893920# diff_1268360_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2916 diff_1293520_901320# diff_1238760_893920# diff_1293520_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2917 diff_1318680_901320# diff_1238760_893920# diff_1318680_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2918 diff_1343840_901320# diff_1238760_893920# diff_1343840_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2919 diff_1369000_901320# diff_1238760_893920# diff_1369000_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2920 diff_1394160_901320# diff_1238760_893920# diff_1394160_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2921 diff_1419320_901320# diff_1238760_893920# diff_1419320_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2922 diff_1444480_901320# diff_1238760_893920# diff_1444480_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2923 diff_1469640_901320# diff_1238760_893920# diff_1469640_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2924 diff_1494800_901320# diff_1238760_893920# diff_1494800_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2925 diff_1519960_901320# diff_1238760_893920# diff_1519960_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2926 diff_1545120_901320# diff_1238760_893920# diff_1545120_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2927 diff_1570280_901320# diff_1238760_893920# diff_1570280_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2928 diff_1595440_901320# diff_1238760_893920# diff_1595440_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2929 diff_1620600_901320# diff_1238760_893920# diff_1620600_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2930 diff_1645760_901320# diff_1238760_893920# diff_1645760_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2931 diff_1670920_901320# diff_1238760_893920# diff_1670920_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2932 diff_1696080_901320# diff_1238760_893920# diff_1696080_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2933 diff_1721240_901320# diff_1238760_893920# diff_1721240_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2934 diff_1746400_901320# diff_1238760_893920# diff_1746400_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2935 diff_1771560_901320# diff_1238760_893920# diff_1771560_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2936 diff_1796720_901320# diff_1238760_893920# diff_1796720_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2937 diff_1821880_901320# diff_1238760_893920# diff_1821880_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2938 diff_1847040_901320# diff_1238760_893920# diff_1847040_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2939 diff_1872200_901320# diff_1238760_893920# diff_1872200_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2940 diff_1897360_901320# diff_1238760_893920# diff_1897360_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2941 diff_1922520_901320# diff_1238760_893920# diff_1922520_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2942 diff_1947680_901320# diff_1238760_893920# diff_1947680_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2943 diff_1972840_901320# diff_1238760_893920# diff_1972840_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2944 diff_1998000_901320# diff_1238760_893920# diff_1998000_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2945 diff_2023160_901320# diff_1238760_893920# diff_2023160_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2946 diff_2048320_901320# diff_1238760_893920# diff_2048320_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2947 diff_2073480_901320# diff_1238760_893920# diff_2073480_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2948 diff_2098640_901320# diff_1238760_893920# diff_2098640_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2949 diff_2123800_901320# diff_1238760_893920# diff_2123800_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2950 diff_2148960_901320# diff_1238760_893920# diff_2148960_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2951 diff_2174120_901320# diff_1238760_893920# diff_2174120_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2952 diff_2199280_901320# diff_1238760_893920# diff_2199280_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2953 diff_2224440_901320# diff_1238760_893920# diff_2224440_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2954 diff_2249600_901320# diff_1238760_893920# diff_2249600_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2955 diff_2274760_901320# diff_1238760_893920# diff_2274760_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2956 diff_2299920_901320# diff_1238760_893920# diff_2299920_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2957 diff_2325080_901320# diff_1238760_893920# diff_2325080_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2958 diff_2350240_901320# diff_1238760_893920# diff_2350240_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2959 diff_2375400_901320# diff_1238760_893920# diff_2375400_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2960 diff_2400560_901320# diff_1238760_893920# diff_2400560_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2961 diff_2425720_901320# diff_1238760_893920# diff_2425720_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2962 diff_2450880_901320# diff_1238760_893920# diff_2450880_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2963 diff_2476040_901320# diff_1238760_893920# diff_2476040_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2964 diff_2501200_901320# diff_1238760_893920# diff_2501200_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2965 diff_2526360_901320# diff_1238760_893920# diff_2526360_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2966 diff_2551520_901320# diff_1238760_893920# diff_2551520_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2967 diff_2576680_901320# diff_1238760_893920# diff_2576680_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2968 diff_2601840_901320# diff_1238760_893920# diff_2601840_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2969 diff_2627000_901320# diff_1238760_893920# diff_2627000_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2970 diff_2652160_901320# diff_1238760_893920# diff_2652160_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2971 diff_2677320_901320# diff_1238760_893920# diff_2677320_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2972 diff_2702480_901320# diff_1238760_893920# diff_2702480_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2973 diff_2727640_901320# diff_1238760_893920# diff_2727640_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2974 diff_2752800_901320# diff_1238760_893920# diff_2752800_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2975 diff_2777960_901320# diff_1238760_893920# diff_2777960_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2976 diff_2803120_901320# diff_1238760_893920# diff_2803120_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2977 diff_2828280_901320# diff_1238760_893920# diff_2828280_873200# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M2978 Vdd Vdd diff_1238760_865800# GND efet w=7400 l=14800
+ ad=0 pd=0 as=1.32738e+09 ps=281200 
M2979 diff_2920040_858400# diff_2912640_526880# diff_1238760_865800# GND efet w=106560 l=7400
+ ad=1.25113e+09 pd=896880 as=0 ps=0 
M2980 diff_1068560_852480# diff_1068560_852480# diff_1068560_852480# GND efet w=2220 l=2960
+ ad=0 pd=0 as=0 ps=0 
M2981 diff_1068560_852480# diff_1068560_852480# diff_1068560_852480# GND efet w=2960 l=2960
+ ad=0 pd=0 as=0 ps=0 
M2982 GND diff_1115920_809560# diff_1068560_852480# GND efet w=25160 l=8880
+ ad=0 pd=0 as=0 ps=0 
M2983 diff_1243200_873200# diff_1238760_865800# diff_1243200_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2984 diff_1268360_873200# diff_1238760_865800# diff_1268360_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2985 diff_1293520_873200# diff_1238760_865800# diff_1293520_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2986 diff_1318680_873200# diff_1238760_865800# diff_1318680_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2987 diff_1343840_873200# diff_1238760_865800# diff_1343840_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2988 diff_1369000_873200# diff_1238760_865800# diff_1369000_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2989 diff_1394160_873200# diff_1238760_865800# diff_1394160_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2990 diff_1419320_873200# diff_1238760_865800# diff_1419320_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2991 diff_1444480_873200# diff_1238760_865800# diff_1444480_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2992 diff_1469640_873200# diff_1238760_865800# diff_1469640_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2993 diff_1494800_873200# diff_1238760_865800# diff_1494800_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2994 diff_1519960_873200# diff_1238760_865800# diff_1519960_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2995 diff_1545120_873200# diff_1238760_865800# diff_1545120_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2996 diff_1570280_873200# diff_1238760_865800# diff_1570280_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2997 diff_1595440_873200# diff_1238760_865800# diff_1595440_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2998 diff_1620600_873200# diff_1238760_865800# diff_1620600_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M2999 diff_1645760_873200# diff_1238760_865800# diff_1645760_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3000 diff_1670920_873200# diff_1238760_865800# diff_1670920_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3001 diff_1696080_873200# diff_1238760_865800# diff_1696080_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3002 diff_1721240_873200# diff_1238760_865800# diff_1721240_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3003 diff_1746400_873200# diff_1238760_865800# diff_1746400_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3004 diff_1771560_873200# diff_1238760_865800# diff_1771560_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3005 diff_1796720_873200# diff_1238760_865800# diff_1796720_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3006 diff_1821880_873200# diff_1238760_865800# diff_1821880_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3007 diff_1847040_873200# diff_1238760_865800# diff_1847040_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3008 diff_1872200_873200# diff_1238760_865800# diff_1872200_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3009 diff_1897360_873200# diff_1238760_865800# diff_1897360_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3010 diff_1922520_873200# diff_1238760_865800# diff_1922520_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3011 diff_1947680_873200# diff_1238760_865800# diff_1947680_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3012 diff_1972840_873200# diff_1238760_865800# diff_1972840_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3013 diff_1998000_873200# diff_1238760_865800# diff_1998000_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3014 diff_2023160_873200# diff_1238760_865800# diff_2023160_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3015 diff_2048320_873200# diff_1238760_865800# diff_2048320_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3016 diff_2073480_873200# diff_1238760_865800# diff_2073480_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3017 diff_2098640_873200# diff_1238760_865800# diff_2098640_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3018 diff_2123800_873200# diff_1238760_865800# diff_2123800_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3019 diff_2148960_873200# diff_1238760_865800# diff_2148960_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3020 diff_2174120_873200# diff_1238760_865800# diff_2174120_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3021 diff_2199280_873200# diff_1238760_865800# diff_2199280_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3022 diff_2224440_873200# diff_1238760_865800# diff_2224440_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3023 diff_2249600_873200# diff_1238760_865800# diff_2249600_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3024 diff_2274760_873200# diff_1238760_865800# diff_2274760_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3025 diff_2299920_873200# diff_1238760_865800# diff_2299920_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3026 diff_2325080_873200# diff_1238760_865800# diff_2325080_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3027 diff_2350240_873200# diff_1238760_865800# diff_2350240_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3028 diff_2375400_873200# diff_1238760_865800# diff_2375400_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3029 diff_2400560_873200# diff_1238760_865800# diff_2400560_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3030 diff_2425720_873200# diff_1238760_865800# diff_2425720_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3031 diff_2450880_873200# diff_1238760_865800# diff_2450880_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3032 diff_2476040_873200# diff_1238760_865800# diff_2476040_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3033 diff_2501200_873200# diff_1238760_865800# diff_2501200_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3034 diff_2526360_873200# diff_1238760_865800# diff_2526360_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3035 diff_2551520_873200# diff_1238760_865800# diff_2551520_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3036 diff_2576680_873200# diff_1238760_865800# diff_2576680_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3037 diff_2601840_873200# diff_1238760_865800# diff_2601840_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3038 diff_2627000_873200# diff_1238760_865800# diff_2627000_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3039 diff_2652160_873200# diff_1238760_865800# diff_2652160_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3040 diff_2677320_873200# diff_1238760_865800# diff_2677320_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3041 diff_2702480_873200# diff_1238760_865800# diff_2702480_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3042 diff_2727640_873200# diff_1238760_865800# diff_2727640_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3043 diff_2752800_873200# diff_1238760_865800# diff_2752800_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3044 diff_2777960_873200# diff_1238760_865800# diff_2777960_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3045 diff_2803120_873200# diff_1238760_865800# diff_2803120_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3046 diff_2828280_873200# diff_1238760_865800# diff_2828280_846560# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3047 diff_1238760_948680# diff_2940760_526880# diff_2920040_858400# GND efet w=91760 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3048 diff_1238760_920560# Vdd Vdd GND efet w=8880 l=16280
+ ad=1.57709e+09 pd=307840 as=0 ps=0 
M3049 Vdd Vdd diff_1238760_893920# GND efet w=8880 l=13320
+ ad=0 pd=0 as=1.60118e+09 ps=278240 
M3050 diff_2920040_858400# diff_2976280_1228400# diff_1238760_893920# GND efet w=105080 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3051 diff_1243200_846560# diff_1238760_839160# diff_1243200_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3052 diff_1268360_846560# diff_1238760_839160# diff_1268360_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3053 diff_1293520_846560# diff_1238760_839160# diff_1293520_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3054 diff_1318680_846560# diff_1238760_839160# diff_1318680_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3055 diff_1343840_846560# diff_1238760_839160# diff_1343840_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3056 diff_1369000_846560# diff_1238760_839160# diff_1369000_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3057 diff_1394160_846560# diff_1238760_839160# diff_1394160_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3058 diff_1419320_846560# diff_1238760_839160# diff_1419320_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3059 diff_1444480_846560# diff_1238760_839160# diff_1444480_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3060 diff_1469640_846560# diff_1238760_839160# diff_1469640_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3061 diff_1494800_846560# diff_1238760_839160# diff_1494800_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3062 diff_1519960_846560# diff_1238760_839160# diff_1519960_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3063 diff_1545120_846560# diff_1238760_839160# diff_1545120_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3064 diff_1570280_846560# diff_1238760_839160# diff_1570280_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3065 diff_1595440_846560# diff_1238760_839160# diff_1595440_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3066 diff_1620600_846560# diff_1238760_839160# diff_1620600_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3067 diff_1645760_846560# diff_1238760_839160# diff_1645760_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3068 diff_1670920_846560# diff_1238760_839160# diff_1670920_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3069 diff_1696080_846560# diff_1238760_839160# diff_1696080_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3070 diff_1721240_846560# diff_1238760_839160# diff_1721240_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3071 diff_1746400_846560# diff_1238760_839160# diff_1746400_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3072 diff_1771560_846560# diff_1238760_839160# diff_1771560_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3073 diff_1796720_846560# diff_1238760_839160# diff_1796720_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3074 diff_1821880_846560# diff_1238760_839160# diff_1821880_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3075 diff_1847040_846560# diff_1238760_839160# diff_1847040_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3076 diff_1872200_846560# diff_1238760_839160# diff_1872200_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3077 diff_1897360_846560# diff_1238760_839160# diff_1897360_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3078 diff_1922520_846560# diff_1238760_839160# diff_1922520_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3079 diff_1947680_846560# diff_1238760_839160# diff_1947680_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3080 diff_1972840_846560# diff_1238760_839160# diff_1972840_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3081 diff_1998000_846560# diff_1238760_839160# diff_1998000_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3082 diff_2023160_846560# diff_1238760_839160# diff_2023160_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3083 diff_2048320_846560# diff_1238760_839160# diff_2048320_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3084 diff_2073480_846560# diff_1238760_839160# diff_2073480_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3085 diff_2098640_846560# diff_1238760_839160# diff_2098640_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3086 diff_2123800_846560# diff_1238760_839160# diff_2123800_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3087 diff_2148960_846560# diff_1238760_839160# diff_2148960_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3088 diff_2174120_846560# diff_1238760_839160# diff_2174120_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3089 diff_2199280_846560# diff_1238760_839160# diff_2199280_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3090 diff_2224440_846560# diff_1238760_839160# diff_2224440_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3091 diff_2249600_846560# diff_1238760_839160# diff_2249600_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3092 diff_2274760_846560# diff_1238760_839160# diff_2274760_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3093 diff_2299920_846560# diff_1238760_839160# diff_2299920_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3094 diff_2325080_846560# diff_1238760_839160# diff_2325080_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3095 diff_2350240_846560# diff_1238760_839160# diff_2350240_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3096 diff_2375400_846560# diff_1238760_839160# diff_2375400_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3097 diff_2400560_846560# diff_1238760_839160# diff_2400560_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3098 diff_2425720_846560# diff_1238760_839160# diff_2425720_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3099 diff_2450880_846560# diff_1238760_839160# diff_2450880_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3100 diff_2476040_846560# diff_1238760_839160# diff_2476040_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3101 diff_2501200_846560# diff_1238760_839160# diff_2501200_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3102 diff_2526360_846560# diff_1238760_839160# diff_2526360_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3103 diff_2551520_846560# diff_1238760_839160# diff_2551520_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3104 diff_2576680_846560# diff_1238760_839160# diff_2576680_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3105 diff_2601840_846560# diff_1238760_839160# diff_2601840_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3106 diff_2627000_846560# diff_1238760_839160# diff_2627000_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3107 diff_2652160_846560# diff_1238760_839160# diff_2652160_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3108 diff_2677320_846560# diff_1238760_839160# diff_2677320_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3109 diff_2702480_846560# diff_1238760_839160# diff_2702480_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3110 diff_2727640_846560# diff_1238760_839160# diff_2727640_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3111 diff_2752800_846560# diff_1238760_839160# diff_2752800_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3112 diff_2777960_846560# diff_1238760_839160# diff_2777960_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3113 diff_2803120_846560# diff_1238760_839160# diff_2803120_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3114 diff_2828280_846560# diff_1238760_839160# diff_2828280_818440# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3115 diff_1238760_920560# diff_2998480_1207680# diff_2920040_858400# GND efet w=97680 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3116 diff_2920040_748880# diff_2912640_526880# diff_1238760_756280# GND efet w=108780 l=8880
+ ad=1.87101e+09 pd=888000 as=1.28796e+09 ps=281200 
M3117 diff_1099640_809560# clk2 Vdd GND efet w=14800 l=8880
+ ad=1.0952e+08 pd=44400 as=0 ps=0 
M3118 diff_1115920_809560# diff_1107040_787360# diff_1099640_809560# GND efet w=14800 l=8880
+ ad=7.00928e+08 pd=124320 as=0 ps=0 
M3119 GND diff_417360_463240# diff_1115920_809560# GND efet w=14800 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3120 diff_1243200_818440# diff_1238760_811040# diff_1243200_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3121 diff_1268360_818440# diff_1238760_811040# diff_1268360_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3122 diff_1293520_818440# diff_1238760_811040# diff_1293520_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3123 diff_1318680_818440# diff_1238760_811040# diff_1318680_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3124 diff_1343840_818440# diff_1238760_811040# diff_1343840_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3125 diff_1369000_818440# diff_1238760_811040# diff_1369000_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3126 diff_1394160_818440# diff_1238760_811040# diff_1394160_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3127 diff_1419320_818440# diff_1238760_811040# diff_1419320_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3128 diff_1444480_818440# diff_1238760_811040# diff_1444480_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3129 diff_1469640_818440# diff_1238760_811040# diff_1469640_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3130 diff_1494800_818440# diff_1238760_811040# diff_1494800_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3131 diff_1519960_818440# diff_1238760_811040# diff_1519960_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3132 diff_1545120_818440# diff_1238760_811040# diff_1545120_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3133 diff_1570280_818440# diff_1238760_811040# diff_1570280_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3134 diff_1595440_818440# diff_1238760_811040# diff_1595440_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3135 diff_1620600_818440# diff_1238760_811040# diff_1620600_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3136 diff_1645760_818440# diff_1238760_811040# diff_1645760_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3137 diff_1670920_818440# diff_1238760_811040# diff_1670920_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3138 diff_1696080_818440# diff_1238760_811040# diff_1696080_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3139 diff_1721240_818440# diff_1238760_811040# diff_1721240_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3140 diff_1746400_818440# diff_1238760_811040# diff_1746400_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3141 diff_1771560_818440# diff_1238760_811040# diff_1771560_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3142 diff_1796720_818440# diff_1238760_811040# diff_1796720_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3143 diff_1821880_818440# diff_1238760_811040# diff_1821880_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3144 diff_1847040_818440# diff_1238760_811040# diff_1847040_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3145 diff_1872200_818440# diff_1238760_811040# diff_1872200_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3146 diff_1897360_818440# diff_1238760_811040# diff_1897360_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3147 diff_1922520_818440# diff_1238760_811040# diff_1922520_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3148 diff_1947680_818440# diff_1238760_811040# diff_1947680_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3149 diff_1972840_818440# diff_1238760_811040# diff_1972840_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3150 diff_1998000_818440# diff_1238760_811040# diff_1998000_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3151 diff_2023160_818440# diff_1238760_811040# diff_2023160_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3152 diff_2048320_818440# diff_1238760_811040# diff_2048320_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3153 diff_2073480_818440# diff_1238760_811040# diff_2073480_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3154 diff_2098640_818440# diff_1238760_811040# diff_2098640_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3155 diff_2123800_818440# diff_1238760_811040# diff_2123800_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3156 diff_2148960_818440# diff_1238760_811040# diff_2148960_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3157 diff_2174120_818440# diff_1238760_811040# diff_2174120_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3158 diff_2199280_818440# diff_1238760_811040# diff_2199280_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3159 diff_2224440_818440# diff_1238760_811040# diff_2224440_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3160 diff_2249600_818440# diff_1238760_811040# diff_2249600_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3161 diff_2274760_818440# diff_1238760_811040# diff_2274760_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3162 diff_2299920_818440# diff_1238760_811040# diff_2299920_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3163 diff_2325080_818440# diff_1238760_811040# diff_2325080_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3164 diff_2350240_818440# diff_1238760_811040# diff_2350240_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3165 diff_2375400_818440# diff_1238760_811040# diff_2375400_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3166 diff_2400560_818440# diff_1238760_811040# diff_2400560_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3167 diff_2425720_818440# diff_1238760_811040# diff_2425720_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3168 diff_2450880_818440# diff_1238760_811040# diff_2450880_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3169 diff_2476040_818440# diff_1238760_811040# diff_2476040_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3170 diff_2501200_818440# diff_1238760_811040# diff_2501200_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3171 diff_2526360_818440# diff_1238760_811040# diff_2526360_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3172 diff_2551520_818440# diff_1238760_811040# diff_2551520_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3173 diff_2576680_818440# diff_1238760_811040# diff_2576680_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3174 diff_2601840_818440# diff_1238760_811040# diff_2601840_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3175 diff_2627000_818440# diff_1238760_811040# diff_2627000_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3176 diff_2652160_818440# diff_1238760_811040# diff_2652160_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3177 diff_2677320_818440# diff_1238760_811040# diff_2677320_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3178 diff_2702480_818440# diff_1238760_811040# diff_2702480_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3179 diff_2727640_818440# diff_1238760_811040# diff_2727640_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3180 diff_2752800_818440# diff_1238760_811040# diff_2752800_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3181 diff_2777960_818440# diff_1238760_811040# diff_2777960_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3182 diff_2803120_818440# diff_1238760_811040# diff_2803120_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3183 diff_2828280_818440# diff_1238760_811040# diff_2828280_791800# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3184 diff_1238760_839160# Vdd Vdd GND efet w=7400 l=16280
+ ad=1.43033e+09 pd=322640 as=0 ps=0 
M3185 diff_856920_939800# diff_920560_771080# GND GND efet w=14800 l=8880
+ ad=3.76749e+08 pd=85840 as=0 ps=0 
M3186 Vdd Vdd diff_856920_939800# GND efet w=9620 l=62900
+ ad=0 pd=0 as=0 ps=0 
M3187 diff_695600_586080# diff_695600_586080# diff_695600_586080# GND efet w=3700 l=4440
+ ad=1.70413e+09 pd=316720 as=0 ps=0 
M3188 diff_695600_586080# diff_695600_586080# diff_695600_586080# GND efet w=3700 l=5180
+ ad=0 pd=0 as=0 ps=0 
M3189 Vdd Vdd diff_695600_586080# GND efet w=11840 l=20720
+ ad=0 pd=0 as=0 ps=0 
M3190 diff_1243200_791800# diff_1238760_784400# diff_1243200_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3191 diff_1268360_791800# diff_1238760_784400# diff_1268360_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3192 diff_1293520_791800# diff_1238760_784400# diff_1293520_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3193 diff_1318680_791800# diff_1238760_784400# diff_1318680_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3194 diff_1343840_791800# diff_1238760_784400# diff_1343840_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3195 diff_1369000_791800# diff_1238760_784400# diff_1369000_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3196 diff_1394160_791800# diff_1238760_784400# diff_1394160_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3197 diff_1419320_791800# diff_1238760_784400# diff_1419320_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3198 diff_1444480_791800# diff_1238760_784400# diff_1444480_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3199 diff_1469640_791800# diff_1238760_784400# diff_1469640_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3200 diff_1494800_791800# diff_1238760_784400# diff_1494800_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3201 diff_1519960_791800# diff_1238760_784400# diff_1519960_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3202 diff_1545120_791800# diff_1238760_784400# diff_1545120_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3203 diff_1570280_791800# diff_1238760_784400# diff_1570280_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3204 diff_1595440_791800# diff_1238760_784400# diff_1595440_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3205 diff_1620600_791800# diff_1238760_784400# diff_1620600_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3206 diff_1645760_791800# diff_1238760_784400# diff_1645760_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3207 diff_1670920_791800# diff_1238760_784400# diff_1670920_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3208 diff_1696080_791800# diff_1238760_784400# diff_1696080_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3209 diff_1721240_791800# diff_1238760_784400# diff_1721240_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3210 diff_1746400_791800# diff_1238760_784400# diff_1746400_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3211 diff_1771560_791800# diff_1238760_784400# diff_1771560_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3212 diff_1796720_791800# diff_1238760_784400# diff_1796720_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3213 diff_1821880_791800# diff_1238760_784400# diff_1821880_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3214 diff_1847040_791800# diff_1238760_784400# diff_1847040_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3215 diff_1872200_791800# diff_1238760_784400# diff_1872200_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3216 diff_1897360_791800# diff_1238760_784400# diff_1897360_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3217 diff_1922520_791800# diff_1238760_784400# diff_1922520_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3218 diff_1947680_791800# diff_1238760_784400# diff_1947680_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3219 diff_1972840_791800# diff_1238760_784400# diff_1972840_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3220 diff_1998000_791800# diff_1238760_784400# diff_1998000_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3221 diff_2023160_791800# diff_1238760_784400# diff_2023160_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3222 diff_2048320_791800# diff_1238760_784400# diff_2048320_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3223 diff_2073480_791800# diff_1238760_784400# diff_2073480_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3224 diff_2098640_791800# diff_1238760_784400# diff_2098640_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3225 diff_2123800_791800# diff_1238760_784400# diff_2123800_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3226 diff_2148960_791800# diff_1238760_784400# diff_2148960_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3227 diff_2174120_791800# diff_1238760_784400# diff_2174120_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3228 diff_2199280_791800# diff_1238760_784400# diff_2199280_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3229 diff_2224440_791800# diff_1238760_784400# diff_2224440_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3230 diff_2249600_791800# diff_1238760_784400# diff_2249600_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3231 diff_2274760_791800# diff_1238760_784400# diff_2274760_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3232 diff_2299920_791800# diff_1238760_784400# diff_2299920_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3233 diff_2325080_791800# diff_1238760_784400# diff_2325080_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3234 diff_2350240_791800# diff_1238760_784400# diff_2350240_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3235 diff_2375400_791800# diff_1238760_784400# diff_2375400_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3236 diff_2400560_791800# diff_1238760_784400# diff_2400560_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3237 diff_2425720_791800# diff_1238760_784400# diff_2425720_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3238 diff_2450880_791800# diff_1238760_784400# diff_2450880_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3239 diff_2476040_791800# diff_1238760_784400# diff_2476040_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3240 diff_2501200_791800# diff_1238760_784400# diff_2501200_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3241 diff_2526360_791800# diff_1238760_784400# diff_2526360_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3242 diff_2551520_791800# diff_1238760_784400# diff_2551520_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3243 diff_2576680_791800# diff_1238760_784400# diff_2576680_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3244 diff_2601840_791800# diff_1238760_784400# diff_2601840_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3245 diff_2627000_791800# diff_1238760_784400# diff_2627000_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3246 diff_2652160_791800# diff_1238760_784400# diff_2652160_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3247 diff_2677320_791800# diff_1238760_784400# diff_2677320_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3248 diff_2702480_791800# diff_1238760_784400# diff_2702480_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3249 diff_2727640_791800# diff_1238760_784400# diff_2727640_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3250 diff_2752800_791800# diff_1238760_784400# diff_2752800_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3251 diff_2777960_791800# diff_1238760_784400# diff_2777960_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3252 diff_2803120_791800# diff_1238760_784400# diff_2803120_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3253 diff_2828280_791800# diff_1238760_784400# diff_2828280_763680# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3254 Vdd Vdd diff_1238760_756280# GND efet w=7400 l=14800
+ ad=0 pd=0 as=0 ps=0 
M3255 Vdd Vdd diff_769600_586080# GND efet w=11840 l=20720
+ ad=0 pd=0 as=1.29453e+09 ps=233840 
M3256 Vdd Vdd Vdd GND efet w=5180 l=5180
+ ad=0 pd=0 as=0 ps=0 
M3257 Vdd Vdd diff_856920_686720# GND efet w=8880 l=78440
+ ad=0 pd=0 as=1.31205e+09 ps=257520 
M3258 diff_856920_686720# cm diff_856920_608280# GND efet w=96200 l=8880
+ ad=0 pd=0 as=1.08644e+09 ps=213120 
M3259 diff_498760_580160# diff_417360_463240# Vdd GND efet w=16280 l=7400
+ ad=3.8551e+08 pd=79920 as=0 ps=0 
M3260 diff_586080_617160# clk2 diff_498760_580160# GND efet w=16280 l=8880
+ ad=1.68661e+08 pd=53280 as=0 ps=0 
M3261 diff_605320_617160# diff_590520_580160# diff_586080_617160# GND efet w=16280 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3262 Vdd Vdd diff_852480_600880# GND efet w=10360 l=62160
+ ad=0 pd=0 as=1.55299e+09 ps=272320 
M3263 Vdd Vdd diff_932400_560920# GND efet w=8880 l=62160
+ ad=0 pd=0 as=7.27213e+08 ps=159840 
M3264 Vdd Vdd Vdd GND efet w=4440 l=4440
+ ad=0 pd=0 as=0 ps=0 
M3265 diff_1107040_787360# Vdd Vdd GND efet w=8880 l=42920
+ ad=9.70347e+08 pd=201280 as=0 ps=0 
M3266 GND diff_856920_686720# diff_1107040_787360# GND efet w=22200 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3267 diff_1107040_787360# diff_1115920_948680# GND GND efet w=26640 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3268 GND diff_1133680_519480# diff_1107040_787360# GND efet w=22200 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3269 diff_1243200_763680# diff_1238760_756280# diff_1243200_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3270 diff_1268360_763680# diff_1238760_756280# diff_1268360_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3271 diff_1293520_763680# diff_1238760_756280# diff_1293520_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3272 diff_1318680_763680# diff_1238760_756280# diff_1318680_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3273 diff_1343840_763680# diff_1238760_756280# diff_1343840_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3274 diff_1369000_763680# diff_1238760_756280# diff_1369000_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3275 diff_1394160_763680# diff_1238760_756280# diff_1394160_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3276 diff_1419320_763680# diff_1238760_756280# diff_1419320_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3277 diff_1444480_763680# diff_1238760_756280# diff_1444480_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3278 diff_1469640_763680# diff_1238760_756280# diff_1469640_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3279 diff_1494800_763680# diff_1238760_756280# diff_1494800_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3280 diff_1519960_763680# diff_1238760_756280# diff_1519960_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3281 diff_1545120_763680# diff_1238760_756280# diff_1545120_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3282 diff_1570280_763680# diff_1238760_756280# diff_1570280_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3283 diff_1595440_763680# diff_1238760_756280# diff_1595440_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3284 diff_1620600_763680# diff_1238760_756280# diff_1620600_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3285 diff_1645760_763680# diff_1238760_756280# diff_1645760_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3286 diff_1670920_763680# diff_1238760_756280# diff_1670920_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3287 diff_1696080_763680# diff_1238760_756280# diff_1696080_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3288 diff_1721240_763680# diff_1238760_756280# diff_1721240_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3289 diff_1746400_763680# diff_1238760_756280# diff_1746400_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3290 diff_1771560_763680# diff_1238760_756280# diff_1771560_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3291 diff_1796720_763680# diff_1238760_756280# diff_1796720_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3292 diff_1821880_763680# diff_1238760_756280# diff_1821880_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3293 diff_1847040_763680# diff_1238760_756280# diff_1847040_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3294 diff_1872200_763680# diff_1238760_756280# diff_1872200_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3295 diff_1897360_763680# diff_1238760_756280# diff_1897360_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3296 diff_1922520_763680# diff_1238760_756280# diff_1922520_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3297 diff_1947680_763680# diff_1238760_756280# diff_1947680_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3298 diff_1972840_763680# diff_1238760_756280# diff_1972840_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3299 diff_1998000_763680# diff_1238760_756280# diff_1998000_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3300 diff_2023160_763680# diff_1238760_756280# diff_2023160_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3301 diff_2048320_763680# diff_1238760_756280# diff_2048320_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3302 diff_2073480_763680# diff_1238760_756280# diff_2073480_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3303 diff_2098640_763680# diff_1238760_756280# diff_2098640_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3304 diff_2123800_763680# diff_1238760_756280# diff_2123800_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3305 diff_2148960_763680# diff_1238760_756280# diff_2148960_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3306 diff_2174120_763680# diff_1238760_756280# diff_2174120_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3307 diff_2199280_763680# diff_1238760_756280# diff_2199280_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3308 diff_2224440_763680# diff_1238760_756280# diff_2224440_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3309 diff_2249600_763680# diff_1238760_756280# diff_2249600_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3310 diff_2274760_763680# diff_1238760_756280# diff_2274760_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3311 diff_2299920_763680# diff_1238760_756280# diff_2299920_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3312 diff_2325080_763680# diff_1238760_756280# diff_2325080_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3313 diff_2350240_763680# diff_1238760_756280# diff_2350240_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3314 diff_2375400_763680# diff_1238760_756280# diff_2375400_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3315 diff_2400560_763680# diff_1238760_756280# diff_2400560_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3316 diff_2425720_763680# diff_1238760_756280# diff_2425720_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3317 diff_2450880_763680# diff_1238760_756280# diff_2450880_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3318 diff_2476040_763680# diff_1238760_756280# diff_2476040_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3319 diff_2501200_763680# diff_1238760_756280# diff_2501200_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3320 diff_2526360_763680# diff_1238760_756280# diff_2526360_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3321 diff_2551520_763680# diff_1238760_756280# diff_2551520_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3322 diff_2576680_763680# diff_1238760_756280# diff_2576680_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3323 diff_2601840_763680# diff_1238760_756280# diff_2601840_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3324 diff_2627000_763680# diff_1238760_756280# diff_2627000_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3325 diff_2652160_763680# diff_1238760_756280# diff_2652160_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3326 diff_2677320_763680# diff_1238760_756280# diff_2677320_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3327 diff_2702480_763680# diff_1238760_756280# diff_2702480_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3328 diff_2727640_763680# diff_1238760_756280# diff_2727640_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3329 diff_2752800_763680# diff_1238760_756280# diff_2752800_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3330 diff_2777960_763680# diff_1238760_756280# diff_2777960_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3331 diff_2803120_763680# diff_1238760_756280# diff_2803120_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3332 diff_2828280_763680# diff_1238760_756280# diff_2828280_737040# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3333 Vdd Vdd diff_999000_629000# GND efet w=8880 l=63640
+ ad=0 pd=0 as=9.79109e+08 ps=213120 
M3334 diff_1238760_839160# diff_2940760_526880# diff_2920040_748880# GND efet w=91760 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3335 diff_1238760_811040# Vdd Vdd GND efet w=8880 l=14800
+ ad=1.57709e+09 pd=307840 as=0 ps=0 
M3336 Vdd Vdd diff_1238760_784400# GND efet w=8880 l=13320
+ ad=0 pd=0 as=1.61213e+09 ps=278240 
M3337 diff_2920040_748880# diff_2976280_1228400# diff_1238760_784400# GND efet w=103600 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3338 diff_1243200_737040# diff_1238760_729640# diff_1243200_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3339 diff_1268360_737040# diff_1238760_729640# diff_1268360_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3340 diff_1293520_737040# diff_1238760_729640# diff_1293520_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3341 diff_1318680_737040# diff_1238760_729640# diff_1318680_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3342 diff_1343840_737040# diff_1238760_729640# diff_1343840_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3343 diff_1369000_737040# diff_1238760_729640# diff_1369000_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3344 diff_1394160_737040# diff_1238760_729640# diff_1394160_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3345 diff_1419320_737040# diff_1238760_729640# diff_1419320_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3346 diff_1444480_737040# diff_1238760_729640# diff_1444480_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3347 diff_1469640_737040# diff_1238760_729640# diff_1469640_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3348 diff_1494800_737040# diff_1238760_729640# diff_1494800_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3349 diff_1519960_737040# diff_1238760_729640# diff_1519960_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3350 diff_1545120_737040# diff_1238760_729640# diff_1545120_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3351 diff_1570280_737040# diff_1238760_729640# diff_1570280_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3352 diff_1595440_737040# diff_1238760_729640# diff_1595440_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3353 diff_1620600_737040# diff_1238760_729640# diff_1620600_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3354 diff_1645760_737040# diff_1238760_729640# diff_1645760_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3355 diff_1670920_737040# diff_1238760_729640# diff_1670920_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3356 diff_1696080_737040# diff_1238760_729640# diff_1696080_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3357 diff_1721240_737040# diff_1238760_729640# diff_1721240_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3358 diff_1746400_737040# diff_1238760_729640# diff_1746400_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3359 diff_1771560_737040# diff_1238760_729640# diff_1771560_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3360 diff_1796720_737040# diff_1238760_729640# diff_1796720_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3361 diff_1821880_737040# diff_1238760_729640# diff_1821880_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3362 diff_1847040_737040# diff_1238760_729640# diff_1847040_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3363 diff_1872200_737040# diff_1238760_729640# diff_1872200_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3364 diff_1897360_737040# diff_1238760_729640# diff_1897360_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3365 diff_1922520_737040# diff_1238760_729640# diff_1922520_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3366 diff_1947680_737040# diff_1238760_729640# diff_1947680_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3367 diff_1972840_737040# diff_1238760_729640# diff_1972840_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3368 diff_1998000_737040# diff_1238760_729640# diff_1998000_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3369 diff_2023160_737040# diff_1238760_729640# diff_2023160_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3370 diff_2048320_737040# diff_1238760_729640# diff_2048320_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3371 diff_2073480_737040# diff_1238760_729640# diff_2073480_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3372 diff_2098640_737040# diff_1238760_729640# diff_2098640_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3373 diff_2123800_737040# diff_1238760_729640# diff_2123800_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3374 diff_2148960_737040# diff_1238760_729640# diff_2148960_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3375 diff_2174120_737040# diff_1238760_729640# diff_2174120_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3376 diff_2199280_737040# diff_1238760_729640# diff_2199280_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3377 diff_2224440_737040# diff_1238760_729640# diff_2224440_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3378 diff_2249600_737040# diff_1238760_729640# diff_2249600_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3379 diff_2274760_737040# diff_1238760_729640# diff_2274760_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3380 diff_2299920_737040# diff_1238760_729640# diff_2299920_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3381 diff_2325080_737040# diff_1238760_729640# diff_2325080_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3382 diff_2350240_737040# diff_1238760_729640# diff_2350240_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3383 diff_2375400_737040# diff_1238760_729640# diff_2375400_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3384 diff_2400560_737040# diff_1238760_729640# diff_2400560_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3385 diff_2425720_737040# diff_1238760_729640# diff_2425720_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3386 diff_2450880_737040# diff_1238760_729640# diff_2450880_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3387 diff_2476040_737040# diff_1238760_729640# diff_2476040_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3388 diff_2501200_737040# diff_1238760_729640# diff_2501200_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3389 diff_2526360_737040# diff_1238760_729640# diff_2526360_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3390 diff_2551520_737040# diff_1238760_729640# diff_2551520_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3391 diff_2576680_737040# diff_1238760_729640# diff_2576680_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3392 diff_2601840_737040# diff_1238760_729640# diff_2601840_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3393 diff_2627000_737040# diff_1238760_729640# diff_2627000_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3394 diff_2652160_737040# diff_1238760_729640# diff_2652160_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3395 diff_2677320_737040# diff_1238760_729640# diff_2677320_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3396 diff_2702480_737040# diff_1238760_729640# diff_2702480_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3397 diff_2727640_737040# diff_1238760_729640# diff_2727640_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3398 diff_2752800_737040# diff_1238760_729640# diff_2752800_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3399 diff_2777960_737040# diff_1238760_729640# diff_2777960_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3400 diff_2803120_737040# diff_1238760_729640# diff_2803120_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3401 diff_2828280_737040# diff_1238760_729640# diff_2828280_708920# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3402 diff_1238760_811040# diff_2998480_1207680# diff_2920040_748880# GND efet w=97680 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3403 diff_3093200_531320# diff_3023640_1207680# diff_2920040_858400# GND efet w=190920 l=8880
+ ad=-1.95919e+09 pd=1.38824e+06 as=0 ps=0 
M3404 diff_2920040_748880# diff_3045840_1124800# diff_3093200_531320# GND efet w=190920 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3405 diff_2920040_640840# diff_2912640_526880# diff_1238760_646760# GND efet w=108040 l=8140
+ ad=1.24674e+09 pd=899840 as=1.2091e+09 ps=275280 
M3406 diff_1243200_708920# diff_1238760_701520# diff_1243200_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3407 diff_1268360_708920# diff_1238760_701520# diff_1268360_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3408 diff_1293520_708920# diff_1238760_701520# diff_1293520_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3409 diff_1318680_708920# diff_1238760_701520# diff_1318680_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3410 diff_1343840_708920# diff_1238760_701520# diff_1343840_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3411 diff_1369000_708920# diff_1238760_701520# diff_1369000_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3412 diff_1394160_708920# diff_1238760_701520# diff_1394160_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3413 diff_1419320_708920# diff_1238760_701520# diff_1419320_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3414 diff_1444480_708920# diff_1238760_701520# diff_1444480_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3415 diff_1469640_708920# diff_1238760_701520# diff_1469640_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3416 diff_1494800_708920# diff_1238760_701520# diff_1494800_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3417 diff_1519960_708920# diff_1238760_701520# diff_1519960_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3418 diff_1545120_708920# diff_1238760_701520# diff_1545120_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3419 diff_1570280_708920# diff_1238760_701520# diff_1570280_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3420 diff_1595440_708920# diff_1238760_701520# diff_1595440_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3421 diff_1620600_708920# diff_1238760_701520# diff_1620600_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3422 diff_1645760_708920# diff_1238760_701520# diff_1645760_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3423 diff_1670920_708920# diff_1238760_701520# diff_1670920_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3424 diff_1696080_708920# diff_1238760_701520# diff_1696080_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3425 diff_1721240_708920# diff_1238760_701520# diff_1721240_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3426 diff_1746400_708920# diff_1238760_701520# diff_1746400_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3427 diff_1771560_708920# diff_1238760_701520# diff_1771560_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3428 diff_1796720_708920# diff_1238760_701520# diff_1796720_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3429 diff_1821880_708920# diff_1238760_701520# diff_1821880_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3430 diff_1847040_708920# diff_1238760_701520# diff_1847040_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3431 diff_1872200_708920# diff_1238760_701520# diff_1872200_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3432 diff_1897360_708920# diff_1238760_701520# diff_1897360_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3433 diff_1922520_708920# diff_1238760_701520# diff_1922520_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3434 diff_1947680_708920# diff_1238760_701520# diff_1947680_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3435 diff_1972840_708920# diff_1238760_701520# diff_1972840_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3436 diff_1998000_708920# diff_1238760_701520# diff_1998000_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3437 diff_2023160_708920# diff_1238760_701520# diff_2023160_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3438 diff_2048320_708920# diff_1238760_701520# diff_2048320_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3439 diff_2073480_708920# diff_1238760_701520# diff_2073480_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3440 diff_2098640_708920# diff_1238760_701520# diff_2098640_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3441 diff_2123800_708920# diff_1238760_701520# diff_2123800_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3442 diff_2148960_708920# diff_1238760_701520# diff_2148960_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3443 diff_2174120_708920# diff_1238760_701520# diff_2174120_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3444 diff_2199280_708920# diff_1238760_701520# diff_2199280_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3445 diff_2224440_708920# diff_1238760_701520# diff_2224440_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3446 diff_2249600_708920# diff_1238760_701520# diff_2249600_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3447 diff_2274760_708920# diff_1238760_701520# diff_2274760_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3448 diff_2299920_708920# diff_1238760_701520# diff_2299920_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3449 diff_2325080_708920# diff_1238760_701520# diff_2325080_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3450 diff_2350240_708920# diff_1238760_701520# diff_2350240_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3451 diff_2375400_708920# diff_1238760_701520# diff_2375400_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3452 diff_2400560_708920# diff_1238760_701520# diff_2400560_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3453 diff_2425720_708920# diff_1238760_701520# diff_2425720_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3454 diff_2450880_708920# diff_1238760_701520# diff_2450880_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3455 diff_2476040_708920# diff_1238760_701520# diff_2476040_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3456 diff_2501200_708920# diff_1238760_701520# diff_2501200_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3457 diff_2526360_708920# diff_1238760_701520# diff_2526360_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3458 diff_2551520_708920# diff_1238760_701520# diff_2551520_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3459 diff_2576680_708920# diff_1238760_701520# diff_2576680_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3460 diff_2601840_708920# diff_1238760_701520# diff_2601840_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3461 diff_2627000_708920# diff_1238760_701520# diff_2627000_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3462 diff_2652160_708920# diff_1238760_701520# diff_2652160_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3463 diff_2677320_708920# diff_1238760_701520# diff_2677320_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3464 diff_2702480_708920# diff_1238760_701520# diff_2702480_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3465 diff_2727640_708920# diff_1238760_701520# diff_2727640_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3466 diff_2752800_708920# diff_1238760_701520# diff_2752800_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3467 diff_2777960_708920# diff_1238760_701520# diff_2777960_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3468 diff_2803120_708920# diff_1238760_701520# diff_2803120_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3469 diff_2828280_708920# diff_1238760_701520# diff_2828280_682280# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3470 diff_1238760_729640# Vdd Vdd GND efet w=7400 l=16280
+ ad=1.43033e+09 pd=322640 as=0 ps=0 
M3471 diff_957560_602360# Vdd Vdd GND efet w=9620 l=107300
+ ad=5.51981e+08 pd=133200 as=0 ps=0 
M3472 diff_1243200_682280# diff_1238760_674880# diff_1243200_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3473 diff_1268360_682280# diff_1238760_674880# diff_1268360_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3474 diff_1293520_682280# diff_1238760_674880# diff_1293520_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3475 diff_1318680_682280# diff_1238760_674880# diff_1318680_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3476 diff_1343840_682280# diff_1238760_674880# diff_1343840_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3477 diff_1369000_682280# diff_1238760_674880# diff_1369000_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3478 diff_1394160_682280# diff_1238760_674880# diff_1394160_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3479 diff_1419320_682280# diff_1238760_674880# diff_1419320_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3480 diff_1444480_682280# diff_1238760_674880# diff_1444480_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3481 diff_1469640_682280# diff_1238760_674880# diff_1469640_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3482 diff_1494800_682280# diff_1238760_674880# diff_1494800_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3483 diff_1519960_682280# diff_1238760_674880# diff_1519960_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3484 diff_1545120_682280# diff_1238760_674880# diff_1545120_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3485 diff_1570280_682280# diff_1238760_674880# diff_1570280_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3486 diff_1595440_682280# diff_1238760_674880# diff_1595440_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3487 diff_1620600_682280# diff_1238760_674880# diff_1620600_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3488 diff_1645760_682280# diff_1238760_674880# diff_1645760_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3489 diff_1670920_682280# diff_1238760_674880# diff_1670920_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3490 diff_1696080_682280# diff_1238760_674880# diff_1696080_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3491 diff_1721240_682280# diff_1238760_674880# diff_1721240_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3492 diff_1746400_682280# diff_1238760_674880# diff_1746400_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3493 diff_1771560_682280# diff_1238760_674880# diff_1771560_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3494 diff_1796720_682280# diff_1238760_674880# diff_1796720_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3495 diff_1821880_682280# diff_1238760_674880# diff_1821880_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3496 diff_1847040_682280# diff_1238760_674880# diff_1847040_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3497 diff_1872200_682280# diff_1238760_674880# diff_1872200_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3498 diff_1897360_682280# diff_1238760_674880# diff_1897360_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3499 diff_1922520_682280# diff_1238760_674880# diff_1922520_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3500 diff_1947680_682280# diff_1238760_674880# diff_1947680_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3501 diff_1972840_682280# diff_1238760_674880# diff_1972840_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3502 diff_1998000_682280# diff_1238760_674880# diff_1998000_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3503 diff_2023160_682280# diff_1238760_674880# diff_2023160_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3504 diff_2048320_682280# diff_1238760_674880# diff_2048320_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3505 diff_2073480_682280# diff_1238760_674880# diff_2073480_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3506 diff_2098640_682280# diff_1238760_674880# diff_2098640_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3507 diff_2123800_682280# diff_1238760_674880# diff_2123800_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3508 diff_2148960_682280# diff_1238760_674880# diff_2148960_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3509 diff_2174120_682280# diff_1238760_674880# diff_2174120_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3510 diff_2199280_682280# diff_1238760_674880# diff_2199280_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3511 diff_2224440_682280# diff_1238760_674880# diff_2224440_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3512 diff_2249600_682280# diff_1238760_674880# diff_2249600_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3513 diff_2274760_682280# diff_1238760_674880# diff_2274760_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3514 diff_2299920_682280# diff_1238760_674880# diff_2299920_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3515 diff_2325080_682280# diff_1238760_674880# diff_2325080_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3516 diff_2350240_682280# diff_1238760_674880# diff_2350240_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3517 diff_2375400_682280# diff_1238760_674880# diff_2375400_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3518 diff_2400560_682280# diff_1238760_674880# diff_2400560_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3519 diff_2425720_682280# diff_1238760_674880# diff_2425720_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3520 diff_2450880_682280# diff_1238760_674880# diff_2450880_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3521 diff_2476040_682280# diff_1238760_674880# diff_2476040_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3522 diff_2501200_682280# diff_1238760_674880# diff_2501200_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3523 diff_2526360_682280# diff_1238760_674880# diff_2526360_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3524 diff_2551520_682280# diff_1238760_674880# diff_2551520_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3525 diff_2576680_682280# diff_1238760_674880# diff_2576680_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3526 diff_2601840_682280# diff_1238760_674880# diff_2601840_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3527 diff_2627000_682280# diff_1238760_674880# diff_2627000_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3528 diff_2652160_682280# diff_1238760_674880# diff_2652160_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3529 diff_2677320_682280# diff_1238760_674880# diff_2677320_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3530 diff_2702480_682280# diff_1238760_674880# diff_2702480_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3531 diff_2727640_682280# diff_1238760_674880# diff_2727640_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3532 diff_2752800_682280# diff_1238760_674880# diff_2752800_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3533 diff_2777960_682280# diff_1238760_674880# diff_2777960_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3534 diff_2803120_682280# diff_1238760_674880# diff_2803120_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3535 diff_2828280_682280# diff_1238760_674880# diff_2828280_654160# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3536 diff_504680_587560# diff_498760_580160# GND GND efet w=39960 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3537 diff_605320_617160# diff_612720_606800# diff_617160_592000# GND efet w=23680 l=8880
+ ad=0 pd=0 as=4.70936e+08 ps=109520 
M3538 diff_962000_550560# diff_957560_602360# diff_852480_600880# GND efet w=16280 l=8880
+ ad=1.33176e+09 pd=242720 as=0 ps=0 
M3539 diff_612720_606800# diff_999000_629000# diff_962000_550560# GND efet w=16280 l=8880
+ ad=1.59242e+09 pd=296000 as=0 ps=0 
M3540 diff_617160_592000# cm GND GND efet w=41440 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3541 diff_856920_608280# diff_852480_600880# diff_856920_590520# GND efet w=37000 l=8880
+ ad=0 pd=0 as=3.52654e+08 ps=103600 
M3542 diff_852480_600880# diff_852480_600880# diff_852480_600880# GND efet w=1480 l=1480
+ ad=0 pd=0 as=0 ps=0 
M3543 diff_852480_600880# diff_852480_600880# diff_852480_600880# GND efet w=2220 l=3700
+ ad=0 pd=0 as=0 ps=0 
M3544 diff_856920_590520# diff_852480_583120# GND GND efet w=42920 l=8140
+ ad=0 pd=0 as=0 ps=0 
M3545 diff_695600_586080# diff_679320_560920# GND GND efet w=56240 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3546 diff_769600_586080# diff_766640_578680# GND GND efet w=56240 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3547 diff_417360_463240# diff_396640_491360# GND GND efet w=25160 l=8880
+ ad=1.3471e+09 pd=251600 as=0 ps=0 
M3548 diff_472120_463240# diff_452880_491360# GND GND efet w=23680 l=8880
+ ad=1.13901e+09 pd=236800 as=0 ps=0 
M3549 diff_529840_463240# diff_510600_491360# GND GND efet w=25160 l=8880
+ ad=1.04263e+09 pd=230880 as=0 ps=0 
M3550 diff_396640_491360# clk1 diff_356680_563880# GND efet w=13320 l=8880
+ ad=2.10278e+08 pd=68080 as=0 ps=0 
M3551 diff_396640_491360# diff_396640_491360# diff_396640_491360# GND efet w=1480 l=6660
+ ad=0 pd=0 as=0 ps=0 
M3552 diff_396640_491360# diff_396640_491360# diff_396640_491360# GND efet w=2220 l=2960
+ ad=0 pd=0 as=0 ps=0 
M3553 diff_452880_491360# clk2 diff_417360_463240# GND efet w=14800 l=8880
+ ad=2.25611e+08 pd=65120 as=0 ps=0 
M3554 diff_452880_491360# diff_452880_491360# diff_452880_491360# GND efet w=2220 l=3700
+ ad=0 pd=0 as=0 ps=0 
M3555 diff_452880_491360# diff_452880_491360# diff_452880_491360# GND efet w=740 l=1480
+ ad=0 pd=0 as=0 ps=0 
M3556 diff_510600_491360# clk1 diff_472120_463240# GND efet w=14800 l=8880
+ ad=2.1685e+08 pd=68080 as=0 ps=0 
M3557 diff_510600_491360# diff_510600_491360# diff_510600_491360# GND efet w=2960 l=5180
+ ad=0 pd=0 as=0 ps=0 
M3558 GND diff_932400_560920# diff_852480_600880# GND efet w=16280 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3559 diff_584600_463240# diff_566840_491360# GND GND efet w=23680 l=8880
+ ad=1.12587e+09 pd=236800 as=0 ps=0 
M3560 diff_590520_580160# diff_624560_491360# GND GND efet w=25160 l=8880
+ ad=1.30548e+09 pd=260480 as=0 ps=0 
M3561 diff_679320_560920# diff_679320_491360# GND GND efet w=23680 l=8880
+ ad=1.32957e+09 pd=260480 as=0 ps=0 
M3562 diff_756280_463240# diff_737040_491360# GND GND efet w=25160 l=8880
+ ad=1.04263e+09 pd=230880 as=0 ps=0 
M3563 diff_766640_578680# diff_793280_491360# GND GND efet w=23680 l=8880
+ ad=1.29891e+09 pd=260480 as=0 ps=0 
M3564 diff_932400_560920# diff_962000_550560# GND GND efet w=26640 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3565 diff_957560_602360# diff_957560_602360# diff_957560_602360# GND efet w=740 l=2220
+ ad=0 pd=0 as=0 ps=0 
M3566 diff_999000_629000# diff_957560_602360# GND GND efet w=14800 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3567 diff_957560_602360# diff_957560_602360# diff_957560_602360# GND efet w=1480 l=1480
+ ad=0 pd=0 as=0 ps=0 
M3568 diff_962000_550560# diff_962000_550560# diff_962000_550560# GND efet w=2220 l=6660
+ ad=0 pd=0 as=0 ps=0 
M3569 diff_962000_550560# diff_962000_550560# diff_962000_550560# GND efet w=2220 l=5180
+ ad=0 pd=0 as=0 ps=0 
M3570 diff_1115920_572760# clk2 diff_957560_602360# GND efet w=28120 l=8880
+ ad=4.4027e+08 pd=97680 as=0 ps=0 
M3571 diff_1138120_565360# diff_920560_771080# diff_1115920_572760# GND efet w=35520 l=8880
+ ad=1.415e+09 pd=245680 as=0 ps=0 
M3572 Vdd Vdd diff_1238760_646760# GND efet w=7400 l=16280
+ ad=0 pd=0 as=0 ps=0 
M3573 diff_1243200_654160# diff_1238760_646760# diff_1243200_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3574 diff_1268360_654160# diff_1238760_646760# diff_1268360_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3575 diff_1293520_654160# diff_1238760_646760# diff_1293520_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3576 diff_1318680_654160# diff_1238760_646760# diff_1318680_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3577 diff_1343840_654160# diff_1238760_646760# diff_1343840_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3578 diff_1369000_654160# diff_1238760_646760# diff_1369000_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3579 diff_1394160_654160# diff_1238760_646760# diff_1394160_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3580 diff_1419320_654160# diff_1238760_646760# diff_1419320_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3581 diff_1444480_654160# diff_1238760_646760# diff_1444480_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3582 diff_1469640_654160# diff_1238760_646760# diff_1469640_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3583 diff_1494800_654160# diff_1238760_646760# diff_1494800_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3584 diff_1519960_654160# diff_1238760_646760# diff_1519960_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3585 diff_1545120_654160# diff_1238760_646760# diff_1545120_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3586 diff_1570280_654160# diff_1238760_646760# diff_1570280_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3587 diff_1595440_654160# diff_1238760_646760# diff_1595440_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3588 diff_1620600_654160# diff_1238760_646760# diff_1620600_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3589 diff_1645760_654160# diff_1238760_646760# diff_1645760_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3590 diff_1670920_654160# diff_1238760_646760# diff_1670920_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3591 diff_1696080_654160# diff_1238760_646760# diff_1696080_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3592 diff_1721240_654160# diff_1238760_646760# diff_1721240_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3593 diff_1746400_654160# diff_1238760_646760# diff_1746400_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3594 diff_1771560_654160# diff_1238760_646760# diff_1771560_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3595 diff_1796720_654160# diff_1238760_646760# diff_1796720_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3596 diff_1821880_654160# diff_1238760_646760# diff_1821880_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3597 diff_1847040_654160# diff_1238760_646760# diff_1847040_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3598 diff_1872200_654160# diff_1238760_646760# diff_1872200_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3599 diff_1897360_654160# diff_1238760_646760# diff_1897360_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3600 diff_1922520_654160# diff_1238760_646760# diff_1922520_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3601 diff_1947680_654160# diff_1238760_646760# diff_1947680_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3602 diff_1972840_654160# diff_1238760_646760# diff_1972840_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3603 diff_1998000_654160# diff_1238760_646760# diff_1998000_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3604 diff_2023160_654160# diff_1238760_646760# diff_2023160_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3605 diff_2048320_654160# diff_1238760_646760# diff_2048320_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3606 diff_2073480_654160# diff_1238760_646760# diff_2073480_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3607 diff_2098640_654160# diff_1238760_646760# diff_2098640_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3608 diff_2123800_654160# diff_1238760_646760# diff_2123800_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3609 diff_2148960_654160# diff_1238760_646760# diff_2148960_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3610 diff_2174120_654160# diff_1238760_646760# diff_2174120_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3611 diff_2199280_654160# diff_1238760_646760# diff_2199280_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3612 diff_2224440_654160# diff_1238760_646760# diff_2224440_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3613 diff_2249600_654160# diff_1238760_646760# diff_2249600_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3614 diff_2274760_654160# diff_1238760_646760# diff_2274760_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3615 diff_2299920_654160# diff_1238760_646760# diff_2299920_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3616 diff_2325080_654160# diff_1238760_646760# diff_2325080_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3617 diff_2350240_654160# diff_1238760_646760# diff_2350240_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3618 diff_2375400_654160# diff_1238760_646760# diff_2375400_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3619 diff_2400560_654160# diff_1238760_646760# diff_2400560_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3620 diff_2425720_654160# diff_1238760_646760# diff_2425720_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3621 diff_2450880_654160# diff_1238760_646760# diff_2450880_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3622 diff_2476040_654160# diff_1238760_646760# diff_2476040_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3623 diff_2501200_654160# diff_1238760_646760# diff_2501200_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3624 diff_2526360_654160# diff_1238760_646760# diff_2526360_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3625 diff_2551520_654160# diff_1238760_646760# diff_2551520_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3626 diff_2576680_654160# diff_1238760_646760# diff_2576680_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3627 diff_2601840_654160# diff_1238760_646760# diff_2601840_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3628 diff_2627000_654160# diff_1238760_646760# diff_2627000_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3629 diff_2652160_654160# diff_1238760_646760# diff_2652160_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3630 diff_2677320_654160# diff_1238760_646760# diff_2677320_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3631 diff_2702480_654160# diff_1238760_646760# diff_2702480_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3632 diff_2727640_654160# diff_1238760_646760# diff_2727640_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3633 diff_2752800_654160# diff_1238760_646760# diff_2752800_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3634 diff_2777960_654160# diff_1238760_646760# diff_2777960_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3635 diff_2803120_654160# diff_1238760_646760# diff_2803120_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3636 diff_2828280_654160# diff_1238760_646760# diff_2828280_627520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3637 diff_1238760_729640# diff_2940760_526880# diff_2920040_640840# GND efet w=91760 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3638 diff_1238760_701520# Vdd Vdd GND efet w=8880 l=16280
+ ad=1.57709e+09 pd=307840 as=0 ps=0 
M3639 Vdd Vdd diff_1238760_674880# GND efet w=8880 l=17760
+ ad=0 pd=0 as=1.56395e+09 ps=272320 
M3640 diff_2920040_640840# diff_2976280_1228400# diff_1238760_674880# GND efet w=104340 l=8140
+ ad=0 pd=0 as=0 ps=0 
M3641 diff_1243200_627520# diff_1238760_620120# diff_1243200_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3642 diff_1268360_627520# diff_1238760_620120# diff_1268360_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3643 diff_1293520_627520# diff_1238760_620120# diff_1293520_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3644 diff_1318680_627520# diff_1238760_620120# diff_1318680_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3645 diff_1343840_627520# diff_1238760_620120# diff_1343840_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3646 diff_1369000_627520# diff_1238760_620120# diff_1369000_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3647 diff_1394160_627520# diff_1238760_620120# diff_1394160_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3648 diff_1419320_627520# diff_1238760_620120# diff_1419320_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3649 diff_1444480_627520# diff_1238760_620120# diff_1444480_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3650 diff_1469640_627520# diff_1238760_620120# diff_1469640_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3651 diff_1494800_627520# diff_1238760_620120# diff_1494800_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3652 diff_1519960_627520# diff_1238760_620120# diff_1519960_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3653 diff_1545120_627520# diff_1238760_620120# diff_1545120_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3654 diff_1570280_627520# diff_1238760_620120# diff_1570280_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3655 diff_1595440_627520# diff_1238760_620120# diff_1595440_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3656 diff_1620600_627520# diff_1238760_620120# diff_1620600_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3657 diff_1645760_627520# diff_1238760_620120# diff_1645760_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3658 diff_1670920_627520# diff_1238760_620120# diff_1670920_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3659 diff_1696080_627520# diff_1238760_620120# diff_1696080_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3660 diff_1721240_627520# diff_1238760_620120# diff_1721240_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3661 diff_1746400_627520# diff_1238760_620120# diff_1746400_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3662 diff_1771560_627520# diff_1238760_620120# diff_1771560_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3663 diff_1796720_627520# diff_1238760_620120# diff_1796720_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3664 diff_1821880_627520# diff_1238760_620120# diff_1821880_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3665 diff_1847040_627520# diff_1238760_620120# diff_1847040_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3666 diff_1872200_627520# diff_1238760_620120# diff_1872200_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3667 diff_1897360_627520# diff_1238760_620120# diff_1897360_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3668 diff_1922520_627520# diff_1238760_620120# diff_1922520_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3669 diff_1947680_627520# diff_1238760_620120# diff_1947680_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3670 diff_1972840_627520# diff_1238760_620120# diff_1972840_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3671 diff_1998000_627520# diff_1238760_620120# diff_1998000_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3672 diff_2023160_627520# diff_1238760_620120# diff_2023160_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3673 diff_2048320_627520# diff_1238760_620120# diff_2048320_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3674 diff_2073480_627520# diff_1238760_620120# diff_2073480_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3675 diff_2098640_627520# diff_1238760_620120# diff_2098640_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3676 diff_2123800_627520# diff_1238760_620120# diff_2123800_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3677 diff_2148960_627520# diff_1238760_620120# diff_2148960_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3678 diff_2174120_627520# diff_1238760_620120# diff_2174120_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3679 diff_2199280_627520# diff_1238760_620120# diff_2199280_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3680 diff_2224440_627520# diff_1238760_620120# diff_2224440_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3681 diff_2249600_627520# diff_1238760_620120# diff_2249600_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3682 diff_2274760_627520# diff_1238760_620120# diff_2274760_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3683 diff_2299920_627520# diff_1238760_620120# diff_2299920_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3684 diff_2325080_627520# diff_1238760_620120# diff_2325080_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3685 diff_2350240_627520# diff_1238760_620120# diff_2350240_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3686 diff_2375400_627520# diff_1238760_620120# diff_2375400_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3687 diff_2400560_627520# diff_1238760_620120# diff_2400560_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3688 diff_2425720_627520# diff_1238760_620120# diff_2425720_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3689 diff_2450880_627520# diff_1238760_620120# diff_2450880_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3690 diff_2476040_627520# diff_1238760_620120# diff_2476040_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3691 diff_2501200_627520# diff_1238760_620120# diff_2501200_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3692 diff_2526360_627520# diff_1238760_620120# diff_2526360_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3693 diff_2551520_627520# diff_1238760_620120# diff_2551520_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3694 diff_2576680_627520# diff_1238760_620120# diff_2576680_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3695 diff_2601840_627520# diff_1238760_620120# diff_2601840_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3696 diff_2627000_627520# diff_1238760_620120# diff_2627000_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3697 diff_2652160_627520# diff_1238760_620120# diff_2652160_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3698 diff_2677320_627520# diff_1238760_620120# diff_2677320_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3699 diff_2702480_627520# diff_1238760_620120# diff_2702480_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3700 diff_2727640_627520# diff_1238760_620120# diff_2727640_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3701 diff_2752800_627520# diff_1238760_620120# diff_2752800_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3702 diff_2777960_627520# diff_1238760_620120# diff_2777960_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3703 diff_2803120_627520# diff_1238760_620120# diff_2803120_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3704 diff_2828280_627520# diff_1238760_620120# diff_2828280_599400# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3705 diff_1238760_701520# diff_2998480_1207680# diff_2920040_640840# GND efet w=97680 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3706 Vdd Vdd Vdd GND efet w=6660 l=9620
+ ad=0 pd=0 as=0 ps=0 
M3707 Vdd Vdd diff_3069520_1052280# GND efet w=8880 l=17760
+ ad=0 pd=0 as=-5.99762e+08 ps=520960 
M3708 diff_3421760_1235800# Vdd Vdd GND efet w=8880 l=39960
+ ad=0 pd=0 as=0 ps=0 
M3709 diff_3513520_1223960# diff_3427680_599400# diff_3513520_1204720# GND efet w=57720 l=7400
+ ad=0 pd=0 as=6.83405e+08 ps=139120 
M3710 Vdd Vdd Vdd GND efet w=2960 l=5920
+ ad=0 pd=0 as=0 ps=0 
M3711 Vdd Vdd Vdd GND efet w=2220 l=5180
+ ad=0 pd=0 as=0 ps=0 
M3712 Vdd Vdd diff_3421760_1096680# GND efet w=8880 l=39960
+ ad=0 pd=0 as=1.48728e+09 ps=198320 
M3713 diff_3513520_1204720# diff_3369960_677840# GND GND efet w=57720 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3714 diff_3377360_1142560# diff_3343320_1672400# diff_3119840_1102600# GND efet w=25160 l=7400
+ ad=0 pd=0 as=4.79698e+08 ps=88800 
M3715 diff_3421760_1096680# clk2 diff_3377360_1142560# GND efet w=25160 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3716 diff_3476520_1096680# diff_3377360_680800# diff_3421760_1096680# GND efet w=45880 l=7400
+ ad=1.461e+09 pd=245680 as=0 ps=0 
M3717 diff_3377360_1003440# diff_3343320_1672400# diff_3204200_809560# GND efet w=25160 l=7400
+ ad=8.89302e+08 pd=171680 as=4.42461e+08 ps=85840 
M3718 diff_3421760_1050800# clk2 diff_3377360_1003440# GND efet w=25160 l=7400
+ ad=1.75889e+09 pd=260480 as=0 ps=0 
M3719 Vdd Vdd diff_1293520_1043400# GND efet w=8880 l=16280
+ ad=0 pd=0 as=-1.53944e+09 ps=399600 
M3720 Vdd Vdd diff_1226920_1511080# GND efet w=8880 l=16280
+ ad=0 pd=0 as=-1.08822e+09 ps=405520 
M3721 Vdd Vdd diff_3090240_1133680# GND efet w=10360 l=16280
+ ad=0 pd=0 as=-1.26783e+09 ps=402560 
M3722 diff_3377360_1003440# diff_3358120_1041920# diff_3227880_973840# GND efet w=25160 l=7400
+ ad=0 pd=0 as=4.42461e+08 ps=85840 
M3723 GND diff_3204200_809560# diff_3069520_1052280# GND efet w=152440 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3724 diff_1293520_1043400# diff_3227880_973840# GND GND efet w=152440 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3725 GND diff_3287080_973840# diff_1226920_1511080# GND efet w=152440 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3726 diff_3090240_1133680# diff_3313720_973840# GND GND efet w=152440 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3727 diff_3377360_957560# diff_3358120_1041920# diff_3287080_973840# GND efet w=25160 l=7400
+ ad=9.17778e+08 pd=174640 as=4.42461e+08 ps=85840 
M3728 diff_3421760_1050800# Vdd Vdd GND efet w=8880 l=41440
+ ad=0 pd=0 as=0 ps=0 
M3729 Vdd Vdd Vdd GND efet w=3700 l=8140
+ ad=0 pd=0 as=0 ps=0 
M3730 Vdd Vdd Vdd GND efet w=1480 l=5920
+ ad=0 pd=0 as=0 ps=0 
M3731 Vdd Vdd diff_3421760_910200# GND efet w=8880 l=39960
+ ad=0 pd=0 as=1.54423e+09 ps=198320 
M3732 diff_3534240_1110000# diff_3369960_677840# diff_3421760_1235800# GND efet w=47360 l=7400
+ ad=5.60742e+08 pd=118400 as=0 ps=0 
M3733 GND diff_3393640_557960# diff_3534240_1110000# GND efet w=47360 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3734 d0 GND d0 GND efet w=221260 l=138380
+ ad=0 pd=0 as=0 ps=0 
M3735 GND diff_3393640_557960# diff_3476520_1096680# GND efet w=44400 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3736 diff_3504640_985680# diff_3427680_599400# diff_3421760_1050800# GND efet w=44400 l=7400
+ ad=5.25696e+08 pd=112480 as=0 ps=0 
M3737 GND diff_3369960_677840# diff_3504640_985680# GND efet w=44400 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3738 diff_3377360_957560# diff_3343320_1672400# diff_3313720_973840# GND efet w=26640 l=7400
+ ad=0 pd=0 as=5.03792e+08 ps=91760 
M3739 diff_3421760_910200# clk2 diff_3377360_957560# GND efet w=26640 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3740 diff_3476520_910200# diff_3377360_680800# diff_3421760_910200# GND efet w=47360 l=7400
+ ad=5.60742e+08 pd=118400 as=0 ps=0 
M3741 GND diff_3427680_599400# diff_3476520_910200# GND efet w=47360 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3742 Vdd Vdd Vdd GND efet w=2960 l=5180
+ ad=0 pd=0 as=0 ps=0 
M3743 Vdd Vdd Vdd GND efet w=2960 l=5920
+ ad=0 pd=0 as=0 ps=0 
M3744 diff_3369960_677840# Vdd Vdd GND efet w=13320 l=20720
+ ad=-1.65115e+09 pd=417360 as=0 ps=0 
M3745 GND diff_3001440_2148960# diff_3093200_531320# GND efet w=371480 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3746 diff_2920040_531320# diff_2912640_526880# diff_1238760_537240# GND efet w=110260 l=8880
+ ad=1.47893e+09 pd=852480 as=1.30986e+09 ps=281200 
M3747 diff_1243200_599400# diff_1238760_592000# diff_1243200_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3748 diff_1268360_599400# diff_1238760_592000# diff_1268360_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3749 diff_1293520_599400# diff_1238760_592000# diff_1293520_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3750 diff_1318680_599400# diff_1238760_592000# diff_1318680_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3751 diff_1343840_599400# diff_1238760_592000# diff_1343840_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3752 diff_1369000_599400# diff_1238760_592000# diff_1369000_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3753 diff_1394160_599400# diff_1238760_592000# diff_1394160_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3754 diff_1419320_599400# diff_1238760_592000# diff_1419320_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3755 diff_1444480_599400# diff_1238760_592000# diff_1444480_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3756 diff_1469640_599400# diff_1238760_592000# diff_1469640_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3757 diff_1494800_599400# diff_1238760_592000# diff_1494800_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3758 diff_1519960_599400# diff_1238760_592000# diff_1519960_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3759 diff_1545120_599400# diff_1238760_592000# diff_1545120_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3760 diff_1570280_599400# diff_1238760_592000# diff_1570280_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3761 diff_1595440_599400# diff_1238760_592000# diff_1595440_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3762 diff_1620600_599400# diff_1238760_592000# diff_1620600_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3763 diff_1645760_599400# diff_1238760_592000# diff_1645760_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3764 diff_1670920_599400# diff_1238760_592000# diff_1670920_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3765 diff_1696080_599400# diff_1238760_592000# diff_1696080_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3766 diff_1721240_599400# diff_1238760_592000# diff_1721240_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3767 diff_1746400_599400# diff_1238760_592000# diff_1746400_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3768 diff_1771560_599400# diff_1238760_592000# diff_1771560_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3769 diff_1796720_599400# diff_1238760_592000# diff_1796720_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3770 diff_1821880_599400# diff_1238760_592000# diff_1821880_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3771 diff_1847040_599400# diff_1238760_592000# diff_1847040_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3772 diff_1872200_599400# diff_1238760_592000# diff_1872200_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3773 diff_1897360_599400# diff_1238760_592000# diff_1897360_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3774 diff_1922520_599400# diff_1238760_592000# diff_1922520_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3775 diff_1947680_599400# diff_1238760_592000# diff_1947680_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3776 diff_1972840_599400# diff_1238760_592000# diff_1972840_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3777 diff_1998000_599400# diff_1238760_592000# diff_1998000_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3778 diff_2023160_599400# diff_1238760_592000# diff_2023160_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3779 diff_2048320_599400# diff_1238760_592000# diff_2048320_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3780 diff_2073480_599400# diff_1238760_592000# diff_2073480_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3781 diff_2098640_599400# diff_1238760_592000# diff_2098640_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3782 diff_2123800_599400# diff_1238760_592000# diff_2123800_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3783 diff_2148960_599400# diff_1238760_592000# diff_2148960_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3784 diff_2174120_599400# diff_1238760_592000# diff_2174120_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3785 diff_2199280_599400# diff_1238760_592000# diff_2199280_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3786 diff_2224440_599400# diff_1238760_592000# diff_2224440_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3787 diff_2249600_599400# diff_1238760_592000# diff_2249600_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3788 diff_2274760_599400# diff_1238760_592000# diff_2274760_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3789 diff_2299920_599400# diff_1238760_592000# diff_2299920_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3790 diff_2325080_599400# diff_1238760_592000# diff_2325080_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3791 diff_2350240_599400# diff_1238760_592000# diff_2350240_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3792 diff_2375400_599400# diff_1238760_592000# diff_2375400_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3793 diff_2400560_599400# diff_1238760_592000# diff_2400560_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3794 diff_2425720_599400# diff_1238760_592000# diff_2425720_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3795 diff_2450880_599400# diff_1238760_592000# diff_2450880_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3796 diff_2476040_599400# diff_1238760_592000# diff_2476040_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3797 diff_2501200_599400# diff_1238760_592000# diff_2501200_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3798 diff_2526360_599400# diff_1238760_592000# diff_2526360_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3799 diff_2551520_599400# diff_1238760_592000# diff_2551520_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3800 diff_2576680_599400# diff_1238760_592000# diff_2576680_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3801 diff_2601840_599400# diff_1238760_592000# diff_2601840_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3802 diff_2627000_599400# diff_1238760_592000# diff_2627000_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3803 diff_2652160_599400# diff_1238760_592000# diff_2652160_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3804 diff_2677320_599400# diff_1238760_592000# diff_2677320_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3805 diff_2702480_599400# diff_1238760_592000# diff_2702480_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3806 diff_2727640_599400# diff_1238760_592000# diff_2727640_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3807 diff_2752800_599400# diff_1238760_592000# diff_2752800_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3808 diff_2777960_599400# diff_1238760_592000# diff_2777960_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3809 diff_2803120_599400# diff_1238760_592000# diff_2803120_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3810 diff_2828280_599400# diff_1238760_592000# diff_2828280_572760# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.36563e+08 ps=62160 
M3811 diff_1238760_620120# Vdd Vdd GND efet w=7400 l=14800
+ ad=1.43033e+09 pd=322640 as=0 ps=0 
M3812 GND cm diff_1138120_565360# GND efet w=82880 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3813 diff_852480_583120# clk1 GND GND efet w=25160 l=8880
+ ad=1.26386e+09 pd=254560 as=0 ps=0 
M3814 diff_923520_463240# diff_904280_491360# GND GND efet w=23680 l=8880
+ ad=1.13901e+09 pd=236800 as=0 ps=0 
M3815 diff_981240_463240# diff_962000_491360# GND GND efet w=25160 l=8880
+ ad=1.04263e+09 pd=230880 as=0 ps=0 
M3816 diff_510600_491360# diff_510600_491360# diff_510600_491360# GND efet w=1480 l=2220
+ ad=0 pd=0 as=0 ps=0 
M3817 diff_566840_491360# clk2 diff_529840_463240# GND efet w=14800 l=8880
+ ad=2.10278e+08 pd=59200 as=0 ps=0 
M3818 diff_566840_491360# diff_566840_491360# diff_566840_491360# GND efet w=1480 l=2220
+ ad=0 pd=0 as=0 ps=0 
M3819 diff_624560_491360# clk1 diff_584600_463240# GND efet w=14800 l=8880
+ ad=1.94946e+08 pd=65120 as=0 ps=0 
M3820 diff_624560_491360# diff_624560_491360# diff_624560_491360# GND efet w=2960 l=5180
+ ad=0 pd=0 as=0 ps=0 
M3821 diff_624560_491360# diff_624560_491360# diff_624560_491360# GND efet w=1480 l=2220
+ ad=0 pd=0 as=0 ps=0 
M3822 diff_679320_491360# clk2 diff_590520_580160# GND efet w=14800 l=8880
+ ad=2.25611e+08 pd=65120 as=0 ps=0 
M3823 diff_679320_491360# diff_679320_491360# diff_679320_491360# GND efet w=2220 l=3700
+ ad=0 pd=0 as=0 ps=0 
M3824 diff_679320_491360# diff_679320_491360# diff_679320_491360# GND efet w=740 l=1480
+ ad=0 pd=0 as=0 ps=0 
M3825 diff_737040_491360# clk1 diff_679320_560920# GND efet w=14800 l=8880
+ ad=2.1685e+08 pd=68080 as=0 ps=0 
M3826 diff_737040_491360# diff_737040_491360# diff_737040_491360# GND efet w=2960 l=5180
+ ad=0 pd=0 as=0 ps=0 
M3827 diff_737040_491360# diff_737040_491360# diff_737040_491360# GND efet w=1480 l=2220
+ ad=0 pd=0 as=0 ps=0 
M3828 diff_793280_491360# clk2 diff_756280_463240# GND efet w=14800 l=8880
+ ad=2.10278e+08 pd=59200 as=0 ps=0 
M3829 diff_793280_491360# diff_793280_491360# diff_793280_491360# GND efet w=1480 l=2220
+ ad=0 pd=0 as=0 ps=0 
M3830 clk1 clk1 diff_766640_578680# GND efet w=12580 l=11100
+ ad=0 pd=0 as=0 ps=0 
M3831 clk1 clk1 clk1 GND efet w=2960 l=5920
+ ad=0 pd=0 as=0 ps=0 
M3832 clk1 clk1 clk1 GND efet w=2220 l=2960
+ ad=0 pd=0 as=0 ps=0 
M3833 diff_904280_491360# clk2 diff_852480_583120# GND efet w=14800 l=8880
+ ad=2.25611e+08 pd=65120 as=0 ps=0 
M3834 diff_904280_491360# diff_904280_491360# diff_904280_491360# GND efet w=2220 l=3700
+ ad=0 pd=0 as=0 ps=0 
M3835 diff_904280_491360# diff_904280_491360# diff_904280_491360# GND efet w=740 l=1480
+ ad=0 pd=0 as=0 ps=0 
M3836 diff_962000_491360# clk1 diff_923520_463240# GND efet w=14800 l=8880
+ ad=2.1685e+08 pd=68080 as=0 ps=0 
M3837 diff_962000_491360# diff_962000_491360# diff_962000_491360# GND efet w=2960 l=5180
+ ad=0 pd=0 as=0 ps=0 
M3838 diff_1036000_463240# diff_1018240_491360# GND GND efet w=23680 l=8880
+ ad=1.26167e+09 pd=257520 as=0 ps=0 
M3839 diff_920560_771080# diff_1075960_491360# GND GND efet w=25160 l=7400
+ ad=1.14777e+09 pd=245680 as=0 ps=0 
M3840 diff_1243200_572760# diff_1238760_565360# diff_1243200_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3841 diff_1268360_572760# diff_1238760_565360# diff_1268360_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3842 diff_1293520_572760# diff_1238760_565360# diff_1293520_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3843 diff_1318680_572760# diff_1238760_565360# diff_1318680_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3844 diff_1343840_572760# diff_1238760_565360# diff_1343840_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3845 diff_1369000_572760# diff_1238760_565360# diff_1369000_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3846 diff_1394160_572760# diff_1238760_565360# diff_1394160_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3847 diff_1419320_572760# diff_1238760_565360# diff_1419320_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3848 diff_1444480_572760# diff_1238760_565360# diff_1444480_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3849 diff_1469640_572760# diff_1238760_565360# diff_1469640_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3850 diff_1494800_572760# diff_1238760_565360# diff_1494800_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3851 diff_1519960_572760# diff_1238760_565360# diff_1519960_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3852 diff_1545120_572760# diff_1238760_565360# diff_1545120_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3853 diff_1570280_572760# diff_1238760_565360# diff_1570280_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3854 diff_1595440_572760# diff_1238760_565360# diff_1595440_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3855 diff_1620600_572760# diff_1238760_565360# diff_1620600_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3856 diff_1645760_572760# diff_1238760_565360# diff_1645760_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3857 diff_1670920_572760# diff_1238760_565360# diff_1670920_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3858 diff_1696080_572760# diff_1238760_565360# diff_1696080_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3859 diff_1721240_572760# diff_1238760_565360# diff_1721240_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3860 diff_1746400_572760# diff_1238760_565360# diff_1746400_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3861 diff_1771560_572760# diff_1238760_565360# diff_1771560_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3862 diff_1796720_572760# diff_1238760_565360# diff_1796720_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3863 diff_1821880_572760# diff_1238760_565360# diff_1821880_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3864 diff_1847040_572760# diff_1238760_565360# diff_1847040_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3865 diff_1872200_572760# diff_1238760_565360# diff_1872200_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3866 diff_1897360_572760# diff_1238760_565360# diff_1897360_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3867 diff_1922520_572760# diff_1238760_565360# diff_1922520_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3868 diff_1947680_572760# diff_1238760_565360# diff_1947680_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3869 diff_1972840_572760# diff_1238760_565360# diff_1972840_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3870 diff_1998000_572760# diff_1238760_565360# diff_1998000_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3871 diff_2023160_572760# diff_1238760_565360# diff_2023160_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3872 diff_2048320_572760# diff_1238760_565360# diff_2048320_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3873 diff_2073480_572760# diff_1238760_565360# diff_2073480_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3874 diff_2098640_572760# diff_1238760_565360# diff_2098640_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3875 diff_2123800_572760# diff_1238760_565360# diff_2123800_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3876 diff_2148960_572760# diff_1238760_565360# diff_2148960_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3877 diff_2174120_572760# diff_1238760_565360# diff_2174120_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3878 diff_2199280_572760# diff_1238760_565360# diff_2199280_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3879 diff_2224440_572760# diff_1238760_565360# diff_2224440_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3880 diff_2249600_572760# diff_1238760_565360# diff_2249600_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3881 diff_2274760_572760# diff_1238760_565360# diff_2274760_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3882 diff_2299920_572760# diff_1238760_565360# diff_2299920_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3883 diff_2325080_572760# diff_1238760_565360# diff_2325080_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3884 diff_2350240_572760# diff_1238760_565360# diff_2350240_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3885 diff_2375400_572760# diff_1238760_565360# diff_2375400_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3886 diff_2400560_572760# diff_1238760_565360# diff_2400560_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3887 diff_2425720_572760# diff_1238760_565360# diff_2425720_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3888 diff_2450880_572760# diff_1238760_565360# diff_2450880_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3889 diff_2476040_572760# diff_1238760_565360# diff_2476040_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3890 diff_2501200_572760# diff_1238760_565360# diff_2501200_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3891 diff_2526360_572760# diff_1238760_565360# diff_2526360_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3892 diff_2551520_572760# diff_1238760_565360# diff_2551520_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3893 diff_2576680_572760# diff_1238760_565360# diff_2576680_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3894 diff_2601840_572760# diff_1238760_565360# diff_2601840_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3895 diff_2627000_572760# diff_1238760_565360# diff_2627000_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3896 diff_2652160_572760# diff_1238760_565360# diff_2652160_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3897 diff_2677320_572760# diff_1238760_565360# diff_2677320_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3898 diff_2702480_572760# diff_1238760_565360# diff_2702480_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3899 diff_2727640_572760# diff_1238760_565360# diff_2727640_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3900 diff_2752800_572760# diff_1238760_565360# diff_2752800_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3901 diff_2777960_572760# diff_1238760_565360# diff_2777960_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3902 diff_2803120_572760# diff_1238760_565360# diff_2803120_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3903 diff_2828280_572760# diff_1238760_565360# diff_2828280_544640# GND efet w=13320 l=8880
+ ad=0 pd=0 as=2.56277e+08 ps=65120 
M3904 diff_962000_491360# diff_962000_491360# diff_962000_491360# GND efet w=1480 l=2220
+ ad=0 pd=0 as=0 ps=0 
M3905 diff_1018240_491360# clk2 diff_981240_463240# GND efet w=14800 l=8880
+ ad=2.10278e+08 pd=59200 as=0 ps=0 
M3906 diff_1018240_491360# diff_1018240_491360# diff_1018240_491360# GND efet w=1480 l=2220
+ ad=0 pd=0 as=0 ps=0 
M3907 diff_1075960_491360# clk1 diff_1036000_463240# GND efet w=14800 l=8880
+ ad=1.99326e+08 pd=68080 as=0 ps=0 
M3908 diff_1075960_491360# diff_1075960_491360# diff_1075960_491360# GND efet w=2960 l=3700
+ ad=0 pd=0 as=0 ps=0 
M3909 diff_1075960_491360# diff_1075960_491360# diff_1075960_491360# GND efet w=1480 l=2220
+ ad=0 pd=0 as=0 ps=0 
M3910 Vdd Vdd diff_356680_563880# GND efet w=9620 l=43660
+ ad=0 pd=0 as=0 ps=0 
M3911 diff_417360_463240# Vdd Vdd GND efet w=8880 l=42920
+ ad=0 pd=0 as=0 ps=0 
M3912 Vdd Vdd diff_472120_463240# GND efet w=9620 l=45140
+ ad=0 pd=0 as=0 ps=0 
M3913 diff_529840_463240# Vdd Vdd GND efet w=8880 l=41440
+ ad=0 pd=0 as=0 ps=0 
M3914 Vdd Vdd diff_584600_463240# GND efet w=9620 l=46620
+ ad=0 pd=0 as=0 ps=0 
M3915 diff_590520_580160# Vdd Vdd GND efet w=8880 l=41440
+ ad=0 pd=0 as=0 ps=0 
M3916 Vdd Vdd diff_679320_560920# GND efet w=9620 l=45140
+ ad=0 pd=0 as=0 ps=0 
M3917 diff_756280_463240# Vdd Vdd GND efet w=8880 l=41440
+ ad=0 pd=0 as=0 ps=0 
M3918 Vdd Vdd diff_766640_578680# GND efet w=9620 l=46620
+ ad=0 pd=0 as=0 ps=0 
M3919 diff_852480_583120# Vdd Vdd GND efet w=8880 l=42920
+ ad=0 pd=0 as=0 ps=0 
M3920 Vdd Vdd diff_923520_463240# GND efet w=9620 l=45140
+ ad=0 pd=0 as=0 ps=0 
M3921 diff_981240_463240# Vdd Vdd GND efet w=8880 l=41440
+ ad=0 pd=0 as=0 ps=0 
M3922 Vdd Vdd diff_1036000_463240# GND efet w=9620 l=46620
+ ad=0 pd=0 as=0 ps=0 
M3923 diff_920560_771080# Vdd Vdd GND efet w=8880 l=41440
+ ad=0 pd=0 as=0 ps=0 
M3924 cl GND GND GND efet w=121360 l=8880
+ ad=1.93672e+09 pd=1.19288e+06 as=0 ps=0 
M3925 Vdd Vdd diff_1238760_537240# GND efet w=7400 l=14800
+ ad=0 pd=0 as=0 ps=0 
M3926 diff_1243200_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=-4.76848e+08 ps=3.42472e+06 
M3927 diff_1268360_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3928 diff_1293520_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3929 diff_1318680_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3930 diff_1343840_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3931 diff_1369000_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3932 diff_1394160_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3933 diff_1419320_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3934 diff_1444480_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3935 diff_1469640_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3936 diff_1494800_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3937 diff_1519960_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3938 diff_1545120_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3939 diff_1570280_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3940 diff_1595440_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3941 diff_1620600_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3942 diff_1645760_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3943 diff_1670920_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3944 diff_1696080_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3945 diff_1721240_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3946 diff_1746400_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3947 diff_1771560_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3948 diff_1796720_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3949 diff_1821880_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3950 diff_1847040_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3951 diff_1872200_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3952 diff_1897360_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3953 diff_1922520_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3954 diff_1947680_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3955 diff_1972840_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3956 diff_1998000_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3957 diff_2023160_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3958 diff_2048320_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3959 diff_2073480_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3960 diff_2098640_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3961 diff_2123800_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3962 diff_2148960_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3963 diff_2174120_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3964 diff_2199280_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3965 diff_2224440_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3966 diff_2249600_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3967 diff_2274760_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3968 diff_2299920_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3969 diff_2325080_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3970 diff_2350240_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3971 diff_2375400_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3972 diff_2400560_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3973 diff_2425720_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3974 diff_2450880_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3975 diff_2476040_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3976 diff_2501200_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3977 diff_2526360_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3978 diff_2551520_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3979 diff_2576680_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3980 diff_2601840_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3981 diff_2627000_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3982 diff_2652160_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3983 diff_2677320_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3984 diff_2702480_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3985 diff_2727640_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3986 diff_2752800_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3987 diff_2777960_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3988 diff_2803120_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3989 diff_2828280_544640# diff_1238760_537240# diff_1243200_516520# GND efet w=13320 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3990 diff_1238760_620120# diff_2940760_526880# diff_2920040_531320# GND efet w=91760 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3991 diff_1238760_592000# Vdd Vdd GND efet w=8880 l=14800
+ ad=1.57709e+09 pd=307840 as=0 ps=0 
M3992 Vdd Vdd diff_1238760_565360# GND efet w=8880 l=14800
+ ad=0 pd=0 as=1.49823e+09 ps=272320 
M3993 diff_2920040_531320# diff_2976280_1228400# diff_1238760_565360# GND efet w=102120 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3994 diff_1238760_592000# diff_2998480_1207680# diff_2920040_531320# GND efet w=97680 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3995 diff_3093200_531320# diff_3069520_1052280# diff_2920040_640840# GND efet w=190920 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3996 diff_2920040_531320# diff_3090240_1133680# diff_3093200_531320# GND efet w=199800 l=8880
+ ad=0 pd=0 as=0 ps=0 
M3997 diff_3369960_677840# d0 GND GND efet w=211640 l=7400
+ ad=0 pd=0 as=0 ps=0 
M3998 diff_3526840_754800# diff_3369960_677840# diff_1173640_538720# GND efet w=102120 l=7400
+ ad=1.26386e+09 pd=230880 as=7.34191e+08 ps=867280 
M3999 diff_3492800_1302400# diff_3393640_557960# diff_3526840_754800# GND efet w=103600 l=7400
+ ad=0 pd=0 as=0 ps=0 
M4000 diff_3377360_680800# diff_3369960_677840# GND GND efet w=54760 l=7400
+ ad=1.10177e+09 pd=189440 as=0 ps=0 
M4001 diff_3377360_680800# Vdd Vdd GND efet w=8880 l=20720
+ ad=0 pd=0 as=0 ps=0 
M4002 diff_3427680_599400# Vdd Vdd GND efet w=11840 l=20720
+ ad=8.82731e+08 pd=153920 as=0 ps=0 
M4003 Vdd Vdd diff_3393640_557960# GND efet w=8880 l=22200
+ ad=0 pd=0 as=-1.01375e+09 ps=639360 
M4004 GND diff_3393640_557960# diff_3427680_599400# GND efet w=54760 l=7400
+ ad=0 pd=0 as=0 ps=0 
M4005 diff_3393640_557960# d1 GND GND efet w=211640 l=7400
+ ad=0 pd=0 as=0 ps=0 
M4006 GND diff_1173640_538720# diff_612720_606800# GND efet w=23680 l=8880
+ ad=0 pd=0 as=0 ps=0 
M4007 diff_1243200_516520# diff_1237280_2100120# GND GND efet w=763680 l=8880
+ ad=0 pd=0 as=0 ps=0 
M4008 diff_1243200_516520# diff_2043880_2100120# Vdd GND efet w=793280 l=8880
+ ad=0 pd=0 as=0 ps=0 
M4009 Vdd Vdd Vdd GND efet w=3700 l=5920
+ ad=0 pd=0 as=0 ps=0 
M4010 Vdd Vdd Vdd GND efet w=2960 l=8140
+ ad=0 pd=0 as=0 ps=0 
M4011 Vdd Vdd diff_612720_606800# GND efet w=10360 l=41440
+ ad=0 pd=0 as=0 ps=0 
M4012 Vdd Vdd Vdd GND efet w=740 l=2220
+ ad=0 pd=0 as=0 ps=0 
M4013 Vdd Vdd Vdd GND efet w=2960 l=3700
+ ad=0 pd=0 as=0 ps=0 
M4014 diff_1133680_519480# Vdd Vdd GND efet w=9620 l=51060
+ ad=0 pd=0 as=0 ps=0 
M4015 Vdd Vdd diff_1173640_538720# GND efet w=11100 l=42180
+ ad=0 pd=0 as=0 ps=0 
M4016 cm GND GND GND efet w=122840 l=8880
+ ad=1.0518e+09 pd=950160 as=0 ps=0 
C0 metal_2255520_227920# gnd! 8.9fF ;**FLOATING
C1 metal_2233320_232360# gnd! 11.4fF ;**FLOATING
C2 metal_2107520_192400# gnd! 10.8fF ;**FLOATING
C3 metal_2100120_192400# gnd! 4.5fF ;**FLOATING
C4 metal_2132680_220520# gnd! 32.1fF ;**FLOATING
C5 metal_2043880_205720# gnd! 12.6fF ;**FLOATING
C6 metal_2212600_193880# gnd! 16.2fF ;**FLOATING
C7 metal_2199280_227920# gnd! 8.9fF ;**FLOATING
C8 metal_2033520_201280# gnd! 27.9fF ;**FLOATING
C9 metal_507640_201280# gnd! 28.7fF ;**FLOATING
C10 metal_445480_210160# gnd! 60.5fF ;**FLOATING
C11 metal_384800_213120# gnd! 63.3fF ;**FLOATING
C12 metal_327080_223480# gnd! 57.6fF ;**FLOATING
C13 diff_3233800_85840# gnd! 2311.4fF ;**FLOATING
C14 diff_3526840_754800# gnd! 149.5fF
C15 diff_1243200_516520# gnd! 2148.9fF
C16 diff_1173640_538720# gnd! 844.7fF
C17 diff_2828280_544640# gnd! 38.4fF
C18 diff_2803120_544640# gnd! 38.4fF
C19 diff_2777960_544640# gnd! 38.4fF
C20 diff_2752800_544640# gnd! 38.4fF
C21 diff_2727640_544640# gnd! 38.4fF
C22 diff_2702480_544640# gnd! 38.4fF
C23 diff_2677320_544640# gnd! 38.4fF
C24 diff_2652160_544640# gnd! 38.4fF
C25 diff_2627000_544640# gnd! 38.4fF
C26 diff_2601840_544640# gnd! 38.4fF
C27 diff_2576680_544640# gnd! 38.4fF
C28 diff_2551520_544640# gnd! 38.4fF
C29 diff_2526360_544640# gnd! 38.4fF
C30 diff_2501200_544640# gnd! 38.4fF
C31 diff_2476040_544640# gnd! 38.4fF
C32 diff_2450880_544640# gnd! 38.4fF
C33 diff_2425720_544640# gnd! 38.4fF
C34 diff_2400560_544640# gnd! 38.4fF
C35 diff_2375400_544640# gnd! 38.4fF
C36 diff_2350240_544640# gnd! 38.4fF
C37 diff_2325080_544640# gnd! 38.4fF
C38 diff_2299920_544640# gnd! 38.4fF
C39 diff_2274760_544640# gnd! 38.4fF
C40 diff_2249600_544640# gnd! 38.4fF
C41 diff_2224440_544640# gnd! 38.4fF
C42 diff_2199280_544640# gnd! 38.4fF
C43 diff_2174120_544640# gnd! 38.4fF
C44 diff_2148960_544640# gnd! 38.4fF
C45 diff_2123800_544640# gnd! 38.4fF
C46 diff_2098640_544640# gnd! 38.4fF
C47 diff_2073480_544640# gnd! 38.4fF
C48 diff_2048320_544640# gnd! 38.4fF
C49 diff_2023160_544640# gnd! 38.4fF
C50 diff_1998000_544640# gnd! 38.4fF
C51 diff_1972840_544640# gnd! 38.4fF
C52 diff_1947680_544640# gnd! 38.4fF
C53 diff_1922520_544640# gnd! 38.4fF
C54 diff_1897360_544640# gnd! 38.4fF
C55 diff_1872200_544640# gnd! 38.4fF
C56 diff_1847040_544640# gnd! 38.4fF
C57 diff_1821880_544640# gnd! 38.4fF
C58 diff_1796720_544640# gnd! 38.4fF
C59 diff_1771560_544640# gnd! 38.4fF
C60 diff_1746400_544640# gnd! 38.4fF
C61 diff_1721240_544640# gnd! 38.4fF
C62 diff_1696080_544640# gnd! 38.4fF
C63 diff_1670920_544640# gnd! 38.4fF
C64 diff_1645760_544640# gnd! 38.4fF
C65 diff_1620600_544640# gnd! 38.4fF
C66 diff_1595440_544640# gnd! 38.4fF
C67 diff_1570280_544640# gnd! 38.4fF
C68 diff_1545120_544640# gnd! 38.4fF
C69 diff_1519960_544640# gnd! 38.4fF
C70 diff_1494800_544640# gnd! 38.4fF
C71 diff_1469640_544640# gnd! 38.4fF
C72 diff_1444480_544640# gnd! 38.4fF
C73 diff_1419320_544640# gnd! 38.4fF
C74 diff_1394160_544640# gnd! 38.4fF
C75 diff_1369000_544640# gnd! 38.4fF
C76 diff_1343840_544640# gnd! 38.4fF
C77 diff_1318680_544640# gnd! 38.4fF
C78 diff_1293520_544640# gnd! 38.4fF
C79 diff_1268360_544640# gnd! 38.4fF
C80 diff_1243200_544640# gnd! 38.4fF
C81 diff_1238760_565360# gnd! 954.5fF
C82 diff_2828280_572760# gnd! 36.1fF
C83 diff_2803120_572760# gnd! 36.1fF
C84 diff_2777960_572760# gnd! 36.1fF
C85 diff_2752800_572760# gnd! 36.1fF
C86 diff_2727640_572760# gnd! 36.1fF
C87 diff_2702480_572760# gnd! 36.1fF
C88 diff_2677320_572760# gnd! 36.1fF
C89 diff_2652160_572760# gnd! 36.1fF
C90 diff_2627000_572760# gnd! 36.1fF
C91 diff_2601840_572760# gnd! 36.1fF
C92 diff_2576680_572760# gnd! 36.1fF
C93 diff_2551520_572760# gnd! 36.1fF
C94 diff_2526360_572760# gnd! 36.1fF
C95 diff_2501200_572760# gnd! 36.1fF
C96 diff_2476040_572760# gnd! 36.1fF
C97 diff_2450880_572760# gnd! 36.1fF
C98 diff_2425720_572760# gnd! 36.1fF
C99 diff_2400560_572760# gnd! 36.1fF
C100 diff_2375400_572760# gnd! 36.1fF
C101 diff_2350240_572760# gnd! 36.1fF
C102 diff_2325080_572760# gnd! 36.1fF
C103 diff_2299920_572760# gnd! 36.1fF
C104 diff_2274760_572760# gnd! 36.1fF
C105 diff_2249600_572760# gnd! 36.1fF
C106 diff_2224440_572760# gnd! 36.1fF
C107 diff_2199280_572760# gnd! 36.1fF
C108 diff_2174120_572760# gnd! 36.1fF
C109 diff_2148960_572760# gnd! 36.1fF
C110 diff_2123800_572760# gnd! 36.1fF
C111 diff_2098640_572760# gnd! 36.1fF
C112 diff_2073480_572760# gnd! 36.1fF
C113 diff_2048320_572760# gnd! 36.1fF
C114 diff_2023160_572760# gnd! 36.1fF
C115 diff_1998000_572760# gnd! 36.1fF
C116 diff_1972840_572760# gnd! 36.1fF
C117 diff_1947680_572760# gnd! 36.1fF
C118 diff_1922520_572760# gnd! 36.1fF
C119 diff_1897360_572760# gnd! 36.1fF
C120 diff_1872200_572760# gnd! 36.1fF
C121 diff_1847040_572760# gnd! 36.1fF
C122 diff_1821880_572760# gnd! 36.1fF
C123 diff_1796720_572760# gnd! 36.1fF
C124 diff_1771560_572760# gnd! 36.1fF
C125 diff_1746400_572760# gnd! 36.1fF
C126 diff_1721240_572760# gnd! 36.1fF
C127 diff_1696080_572760# gnd! 36.1fF
C128 diff_1670920_572760# gnd! 36.1fF
C129 diff_1645760_572760# gnd! 36.1fF
C130 diff_1620600_572760# gnd! 36.1fF
C131 diff_1595440_572760# gnd! 36.1fF
C132 diff_1570280_572760# gnd! 36.1fF
C133 diff_1545120_572760# gnd! 36.1fF
C134 diff_1519960_572760# gnd! 36.1fF
C135 diff_1494800_572760# gnd! 36.1fF
C136 diff_1469640_572760# gnd! 36.1fF
C137 diff_1444480_572760# gnd! 36.1fF
C138 diff_1419320_572760# gnd! 36.1fF
C139 diff_1394160_572760# gnd! 36.1fF
C140 diff_1369000_572760# gnd! 36.1fF
C141 diff_1343840_572760# gnd! 36.1fF
C142 diff_1318680_572760# gnd! 36.1fF
C143 diff_1293520_572760# gnd! 36.1fF
C144 diff_1268360_572760# gnd! 36.1fF
C145 diff_981240_463240# gnd! 127.4fF
C146 diff_923520_463240# gnd! 137.6fF
C147 diff_1075960_491360# gnd! 56.1fF
C148 diff_1018240_491360# gnd! 61.4fF
C149 diff_962000_491360# gnd! 62.6fF
C150 diff_904280_491360# gnd! 62.9fF
C151 diff_1243200_572760# gnd! 36.1fF
C152 diff_1238760_592000# gnd! 986.1fF
C153 diff_2828280_599400# gnd! 38.4fF
C154 diff_2803120_599400# gnd! 38.4fF
C155 diff_2777960_599400# gnd! 38.4fF
C156 diff_2752800_599400# gnd! 38.4fF
C157 diff_2727640_599400# gnd! 38.4fF
C158 diff_2702480_599400# gnd! 38.4fF
C159 diff_2677320_599400# gnd! 38.4fF
C160 diff_2652160_599400# gnd! 38.4fF
C161 diff_2627000_599400# gnd! 38.4fF
C162 diff_2601840_599400# gnd! 38.4fF
C163 diff_2576680_599400# gnd! 38.4fF
C164 diff_2551520_599400# gnd! 38.4fF
C165 diff_2526360_599400# gnd! 38.4fF
C166 diff_2501200_599400# gnd! 38.4fF
C167 diff_2476040_599400# gnd! 38.4fF
C168 diff_2450880_599400# gnd! 38.4fF
C169 diff_2425720_599400# gnd! 38.4fF
C170 diff_2400560_599400# gnd! 38.4fF
C171 diff_2375400_599400# gnd! 38.4fF
C172 diff_2350240_599400# gnd! 38.4fF
C173 diff_2325080_599400# gnd! 38.4fF
C174 diff_2299920_599400# gnd! 38.4fF
C175 diff_2274760_599400# gnd! 38.4fF
C176 diff_2249600_599400# gnd! 38.4fF
C177 diff_2224440_599400# gnd! 38.4fF
C178 diff_2199280_599400# gnd! 38.4fF
C179 diff_2174120_599400# gnd! 38.4fF
C180 diff_2148960_599400# gnd! 38.4fF
C181 diff_2123800_599400# gnd! 38.4fF
C182 diff_2098640_599400# gnd! 38.4fF
C183 diff_2073480_599400# gnd! 38.4fF
C184 diff_2048320_599400# gnd! 38.4fF
C185 diff_2023160_599400# gnd! 38.4fF
C186 diff_1998000_599400# gnd! 38.4fF
C187 diff_1972840_599400# gnd! 38.4fF
C188 diff_1947680_599400# gnd! 38.4fF
C189 diff_1922520_599400# gnd! 38.4fF
C190 diff_1897360_599400# gnd! 38.4fF
C191 diff_1872200_599400# gnd! 38.4fF
C192 diff_1847040_599400# gnd! 38.4fF
C193 diff_1821880_599400# gnd! 38.4fF
C194 diff_1796720_599400# gnd! 38.4fF
C195 diff_1771560_599400# gnd! 38.4fF
C196 diff_1746400_599400# gnd! 38.4fF
C197 diff_1721240_599400# gnd! 38.4fF
C198 diff_1696080_599400# gnd! 38.4fF
C199 diff_1670920_599400# gnd! 38.4fF
C200 diff_1645760_599400# gnd! 38.4fF
C201 diff_1620600_599400# gnd! 38.4fF
C202 diff_1595440_599400# gnd! 38.4fF
C203 diff_1570280_599400# gnd! 38.4fF
C204 diff_1545120_599400# gnd! 38.4fF
C205 diff_1519960_599400# gnd! 38.4fF
C206 diff_1494800_599400# gnd! 38.4fF
C207 diff_1469640_599400# gnd! 38.4fF
C208 diff_1444480_599400# gnd! 38.4fF
C209 diff_1419320_599400# gnd! 38.4fF
C210 diff_1394160_599400# gnd! 38.4fF
C211 diff_1369000_599400# gnd! 38.4fF
C212 diff_1343840_599400# gnd! 38.4fF
C213 diff_1318680_599400# gnd! 38.4fF
C214 diff_1293520_599400# gnd! 38.4fF
C215 diff_1268360_599400# gnd! 38.4fF
C216 diff_1243200_599400# gnd! 38.4fF
C217 diff_2920040_531320# gnd! 769.9fF
C218 diff_1238760_537240# gnd! 903.1fF
C219 diff_3476520_910200# gnd! 67.9fF
C220 diff_3421760_910200# gnd! 174.3fF
C221 diff_3504640_985680# gnd! 63.8fF
C222 diff_3534240_1110000# gnd! 67.9fF
C223 diff_3377360_957560# gnd! 136.5fF
C224 diff_3313720_973840# gnd! 171.0fF
C225 diff_3287080_973840# gnd! 166.3fF
C226 diff_3227880_973840# gnd! 184.3fF
C227 diff_3421760_1050800# gnd! 244.1fF
C228 diff_3377360_1003440# gnd! 132.9fF
C229 diff_3204200_809560# gnd! 208.3fF
C230 diff_3476520_1096680# gnd! 216.3fF
C231 diff_3421760_1096680# gnd! 168.6fF
C232 diff_3377360_680800# gnd! 326.3fF
C233 diff_3393640_557960# gnd! 810.5fF
C234 diff_3369960_677840# gnd! 686.5fF
C235 diff_3513520_1204720# gnd! 82.3fF
C236 diff_3427680_599400# gnd! 493.7fF
C237 diff_3513520_1223960# gnd! 82.3fF
C238 diff_1238760_620120# gnd! 939.9fF
C239 diff_2828280_627520# gnd! 36.1fF
C240 diff_2803120_627520# gnd! 36.1fF
C241 diff_2777960_627520# gnd! 36.1fF
C242 diff_2752800_627520# gnd! 36.1fF
C243 diff_2727640_627520# gnd! 36.1fF
C244 diff_2702480_627520# gnd! 36.1fF
C245 diff_2677320_627520# gnd! 36.1fF
C246 diff_2652160_627520# gnd! 36.1fF
C247 diff_2627000_627520# gnd! 36.1fF
C248 diff_2601840_627520# gnd! 36.1fF
C249 diff_2576680_627520# gnd! 36.1fF
C250 diff_2551520_627520# gnd! 36.1fF
C251 diff_2526360_627520# gnd! 36.1fF
C252 diff_2501200_627520# gnd! 36.1fF
C253 diff_2476040_627520# gnd! 36.1fF
C254 diff_2450880_627520# gnd! 36.1fF
C255 diff_2425720_627520# gnd! 36.1fF
C256 diff_2400560_627520# gnd! 36.1fF
C257 diff_2375400_627520# gnd! 36.1fF
C258 diff_2350240_627520# gnd! 36.1fF
C259 diff_2325080_627520# gnd! 36.1fF
C260 diff_2299920_627520# gnd! 36.1fF
C261 diff_2274760_627520# gnd! 36.1fF
C262 diff_2249600_627520# gnd! 36.1fF
C263 diff_2224440_627520# gnd! 36.1fF
C264 diff_2199280_627520# gnd! 36.1fF
C265 diff_2174120_627520# gnd! 36.1fF
C266 diff_2148960_627520# gnd! 36.1fF
C267 diff_2123800_627520# gnd! 36.1fF
C268 diff_2098640_627520# gnd! 36.1fF
C269 diff_2073480_627520# gnd! 36.1fF
C270 diff_2048320_627520# gnd! 36.1fF
C271 diff_2023160_627520# gnd! 36.1fF
C272 diff_1998000_627520# gnd! 36.1fF
C273 diff_1972840_627520# gnd! 36.1fF
C274 diff_1947680_627520# gnd! 36.1fF
C275 diff_1922520_627520# gnd! 36.1fF
C276 diff_1897360_627520# gnd! 36.1fF
C277 diff_1872200_627520# gnd! 36.1fF
C278 diff_1847040_627520# gnd! 36.1fF
C279 diff_1821880_627520# gnd! 36.1fF
C280 diff_1796720_627520# gnd! 36.1fF
C281 diff_1771560_627520# gnd! 36.1fF
C282 diff_1746400_627520# gnd! 36.1fF
C283 diff_1721240_627520# gnd! 36.1fF
C284 diff_1696080_627520# gnd! 36.1fF
C285 diff_1670920_627520# gnd! 36.1fF
C286 diff_1645760_627520# gnd! 36.1fF
C287 diff_1620600_627520# gnd! 36.1fF
C288 diff_1595440_627520# gnd! 36.1fF
C289 diff_1570280_627520# gnd! 36.1fF
C290 diff_1545120_627520# gnd! 36.1fF
C291 diff_1519960_627520# gnd! 36.1fF
C292 diff_1494800_627520# gnd! 36.1fF
C293 diff_1469640_627520# gnd! 36.1fF
C294 diff_1444480_627520# gnd! 36.1fF
C295 diff_1419320_627520# gnd! 36.1fF
C296 diff_1394160_627520# gnd! 36.1fF
C297 diff_1369000_627520# gnd! 36.1fF
C298 diff_1343840_627520# gnd! 36.1fF
C299 diff_1318680_627520# gnd! 36.1fF
C300 diff_1293520_627520# gnd! 36.1fF
C301 diff_1268360_627520# gnd! 36.1fF
C302 diff_1243200_627520# gnd! 36.1fF
C303 diff_2828280_654160# gnd! 38.4fF
C304 diff_2803120_654160# gnd! 38.4fF
C305 diff_2777960_654160# gnd! 38.4fF
C306 diff_2752800_654160# gnd! 38.4fF
C307 diff_2727640_654160# gnd! 38.4fF
C308 diff_2702480_654160# gnd! 38.4fF
C309 diff_2677320_654160# gnd! 38.4fF
C310 diff_2652160_654160# gnd! 38.4fF
C311 diff_2627000_654160# gnd! 38.4fF
C312 diff_2601840_654160# gnd! 38.4fF
C313 diff_2576680_654160# gnd! 38.4fF
C314 diff_2551520_654160# gnd! 38.4fF
C315 diff_2526360_654160# gnd! 38.4fF
C316 diff_2501200_654160# gnd! 38.4fF
C317 diff_2476040_654160# gnd! 38.4fF
C318 diff_2450880_654160# gnd! 38.4fF
C319 diff_2425720_654160# gnd! 38.4fF
C320 diff_2400560_654160# gnd! 38.4fF
C321 diff_2375400_654160# gnd! 38.4fF
C322 diff_2350240_654160# gnd! 38.4fF
C323 diff_2325080_654160# gnd! 38.4fF
C324 diff_2299920_654160# gnd! 38.4fF
C325 diff_2274760_654160# gnd! 38.4fF
C326 diff_2249600_654160# gnd! 38.4fF
C327 diff_2224440_654160# gnd! 38.4fF
C328 diff_2199280_654160# gnd! 38.4fF
C329 diff_2174120_654160# gnd! 38.4fF
C330 diff_2148960_654160# gnd! 38.4fF
C331 diff_2123800_654160# gnd! 38.4fF
C332 diff_2098640_654160# gnd! 38.4fF
C333 diff_2073480_654160# gnd! 38.4fF
C334 diff_2048320_654160# gnd! 38.4fF
C335 diff_2023160_654160# gnd! 38.4fF
C336 diff_1998000_654160# gnd! 38.4fF
C337 diff_1972840_654160# gnd! 38.4fF
C338 diff_1947680_654160# gnd! 38.4fF
C339 diff_1922520_654160# gnd! 38.4fF
C340 diff_1897360_654160# gnd! 38.4fF
C341 diff_1872200_654160# gnd! 38.4fF
C342 diff_1847040_654160# gnd! 38.4fF
C343 diff_1821880_654160# gnd! 38.4fF
C344 diff_1796720_654160# gnd! 38.4fF
C345 diff_1771560_654160# gnd! 38.4fF
C346 diff_1746400_654160# gnd! 38.4fF
C347 diff_1721240_654160# gnd! 38.4fF
C348 diff_1696080_654160# gnd! 38.4fF
C349 diff_1670920_654160# gnd! 38.4fF
C350 diff_1645760_654160# gnd! 38.4fF
C351 diff_1620600_654160# gnd! 38.4fF
C352 diff_1595440_654160# gnd! 38.4fF
C353 diff_1570280_654160# gnd! 38.4fF
C354 diff_1545120_654160# gnd! 38.4fF
C355 diff_1519960_654160# gnd! 38.4fF
C356 diff_1494800_654160# gnd! 38.4fF
C357 diff_1469640_654160# gnd! 38.4fF
C358 diff_1444480_654160# gnd! 38.4fF
C359 diff_1419320_654160# gnd! 38.4fF
C360 diff_1394160_654160# gnd! 38.4fF
C361 diff_1369000_654160# gnd! 38.4fF
C362 diff_1343840_654160# gnd! 38.4fF
C363 diff_1318680_654160# gnd! 38.4fF
C364 diff_1293520_654160# gnd! 38.4fF
C365 diff_1268360_654160# gnd! 38.4fF
C366 diff_1138120_565360# gnd! 166.1fF
C367 diff_1115920_572760# gnd! 53.8fF
C368 diff_756280_463240# gnd! 127.4fF
C369 diff_584600_463240# gnd! 136.3fF
C370 diff_793280_491360# gnd! 62.0fF
C371 diff_737040_491360# gnd! 62.0fF
C372 diff_679320_491360# gnd! 63.5fF
C373 diff_624560_491360# gnd! 59.5fF
C374 diff_566840_491360# gnd! 62.0fF
C375 diff_529840_463240# gnd! 127.4fF
C376 diff_472120_463240# gnd! 137.6fF
C377 diff_510600_491360# gnd! 62.0fF
C378 diff_452880_491360# gnd! 63.5fF
C379 diff_396640_491360# gnd! 60.8fF
C380 diff_766640_578680# gnd! 215.0fF
C381 diff_679320_560920# gnd! 227.5fF
C382 diff_852480_583120# gnd! 205.2fF
C383 diff_856920_590520# gnd! 45.6fF
C384 diff_617160_592000# gnd! 58.0fF
C385 diff_962000_550560# gnd! 207.8fF
C386 diff_356680_563880# gnd! 205.9fF
C387 diff_999000_629000# gnd! 160.3fF
C388 diff_1243200_654160# gnd! 38.4fF
C389 diff_1238760_674880# gnd! 962.2fF
C390 diff_2828280_682280# gnd! 36.1fF
C391 diff_2803120_682280# gnd! 36.1fF
C392 diff_2777960_682280# gnd! 36.1fF
C393 diff_2752800_682280# gnd! 36.1fF
C394 diff_2727640_682280# gnd! 36.1fF
C395 diff_2702480_682280# gnd! 36.1fF
C396 diff_2677320_682280# gnd! 36.1fF
C397 diff_2652160_682280# gnd! 36.1fF
C398 diff_2627000_682280# gnd! 36.1fF
C399 diff_2601840_682280# gnd! 36.1fF
C400 diff_2576680_682280# gnd! 36.1fF
C401 diff_2551520_682280# gnd! 36.1fF
C402 diff_2526360_682280# gnd! 36.1fF
C403 diff_2501200_682280# gnd! 36.1fF
C404 diff_2476040_682280# gnd! 36.1fF
C405 diff_2450880_682280# gnd! 36.1fF
C406 diff_2425720_682280# gnd! 36.1fF
C407 diff_2400560_682280# gnd! 36.1fF
C408 diff_2375400_682280# gnd! 36.1fF
C409 diff_2350240_682280# gnd! 36.1fF
C410 diff_2325080_682280# gnd! 36.1fF
C411 diff_2299920_682280# gnd! 36.1fF
C412 diff_2274760_682280# gnd! 36.1fF
C413 diff_2249600_682280# gnd! 36.1fF
C414 diff_2224440_682280# gnd! 36.1fF
C415 diff_2199280_682280# gnd! 36.1fF
C416 diff_2174120_682280# gnd! 36.1fF
C417 diff_2148960_682280# gnd! 36.1fF
C418 diff_2123800_682280# gnd! 36.1fF
C419 diff_2098640_682280# gnd! 36.1fF
C420 diff_2073480_682280# gnd! 36.1fF
C421 diff_2048320_682280# gnd! 36.1fF
C422 diff_2023160_682280# gnd! 36.1fF
C423 diff_1998000_682280# gnd! 36.1fF
C424 diff_1972840_682280# gnd! 36.1fF
C425 diff_1947680_682280# gnd! 36.1fF
C426 diff_1922520_682280# gnd! 36.1fF
C427 diff_1897360_682280# gnd! 36.1fF
C428 diff_1872200_682280# gnd! 36.1fF
C429 diff_1847040_682280# gnd! 36.1fF
C430 diff_1821880_682280# gnd! 36.1fF
C431 diff_1796720_682280# gnd! 36.1fF
C432 diff_1771560_682280# gnd! 36.1fF
C433 diff_1746400_682280# gnd! 36.1fF
C434 diff_1721240_682280# gnd! 36.1fF
C435 diff_1696080_682280# gnd! 36.1fF
C436 diff_1670920_682280# gnd! 36.1fF
C437 diff_1645760_682280# gnd! 36.1fF
C438 diff_1620600_682280# gnd! 36.1fF
C439 diff_1595440_682280# gnd! 36.1fF
C440 diff_1570280_682280# gnd! 36.1fF
C441 diff_1545120_682280# gnd! 36.1fF
C442 diff_1519960_682280# gnd! 36.1fF
C443 diff_1494800_682280# gnd! 36.1fF
C444 diff_1469640_682280# gnd! 36.1fF
C445 diff_1444480_682280# gnd! 36.1fF
C446 diff_1419320_682280# gnd! 36.1fF
C447 diff_1394160_682280# gnd! 36.1fF
C448 diff_1369000_682280# gnd! 36.1fF
C449 diff_1343840_682280# gnd! 36.1fF
C450 diff_1318680_682280# gnd! 36.1fF
C451 diff_1293520_682280# gnd! 36.1fF
C452 diff_1268360_682280# gnd! 36.1fF
C453 diff_1243200_682280# gnd! 36.1fF
C454 diff_1238760_701520# gnd! 984.6fF
C455 diff_2828280_708920# gnd! 38.4fF
C456 diff_2803120_708920# gnd! 38.4fF
C457 diff_2777960_708920# gnd! 38.4fF
C458 diff_2752800_708920# gnd! 38.4fF
C459 diff_2727640_708920# gnd! 38.4fF
C460 diff_2702480_708920# gnd! 38.4fF
C461 diff_2677320_708920# gnd! 38.4fF
C462 diff_2652160_708920# gnd! 38.4fF
C463 diff_2627000_708920# gnd! 38.4fF
C464 diff_2601840_708920# gnd! 38.4fF
C465 diff_2576680_708920# gnd! 38.4fF
C466 diff_2551520_708920# gnd! 38.4fF
C467 diff_2526360_708920# gnd! 38.4fF
C468 diff_2501200_708920# gnd! 38.4fF
C469 diff_2476040_708920# gnd! 38.4fF
C470 diff_2450880_708920# gnd! 38.4fF
C471 diff_2425720_708920# gnd! 38.4fF
C472 diff_2400560_708920# gnd! 38.4fF
C473 diff_2375400_708920# gnd! 38.4fF
C474 diff_2350240_708920# gnd! 38.4fF
C475 diff_2325080_708920# gnd! 38.4fF
C476 diff_2299920_708920# gnd! 38.4fF
C477 diff_2274760_708920# gnd! 38.4fF
C478 diff_2249600_708920# gnd! 38.4fF
C479 diff_2224440_708920# gnd! 38.4fF
C480 diff_2199280_708920# gnd! 38.4fF
C481 diff_2174120_708920# gnd! 38.4fF
C482 diff_2148960_708920# gnd! 38.4fF
C483 diff_2123800_708920# gnd! 38.4fF
C484 diff_2098640_708920# gnd! 38.4fF
C485 diff_2073480_708920# gnd! 38.4fF
C486 diff_2048320_708920# gnd! 38.4fF
C487 diff_2023160_708920# gnd! 38.4fF
C488 diff_1998000_708920# gnd! 38.4fF
C489 diff_1972840_708920# gnd! 38.4fF
C490 diff_1947680_708920# gnd! 38.4fF
C491 diff_1922520_708920# gnd! 38.4fF
C492 diff_1897360_708920# gnd! 38.4fF
C493 diff_1872200_708920# gnd! 38.4fF
C494 diff_1847040_708920# gnd! 38.4fF
C495 diff_1821880_708920# gnd! 38.4fF
C496 diff_1796720_708920# gnd! 38.4fF
C497 diff_1771560_708920# gnd! 38.4fF
C498 diff_1746400_708920# gnd! 38.4fF
C499 diff_1721240_708920# gnd! 38.4fF
C500 diff_1696080_708920# gnd! 38.4fF
C501 diff_1670920_708920# gnd! 38.4fF
C502 diff_1645760_708920# gnd! 38.4fF
C503 diff_1620600_708920# gnd! 38.4fF
C504 diff_1595440_708920# gnd! 38.4fF
C505 diff_1570280_708920# gnd! 38.4fF
C506 diff_1545120_708920# gnd! 38.4fF
C507 diff_1519960_708920# gnd! 38.4fF
C508 diff_1494800_708920# gnd! 38.4fF
C509 diff_1469640_708920# gnd! 38.4fF
C510 diff_1444480_708920# gnd! 38.4fF
C511 diff_1419320_708920# gnd! 38.4fF
C512 diff_1394160_708920# gnd! 38.4fF
C513 diff_1369000_708920# gnd! 38.4fF
C514 diff_1343840_708920# gnd! 38.4fF
C515 diff_1318680_708920# gnd! 38.4fF
C516 diff_1293520_708920# gnd! 38.4fF
C517 diff_1268360_708920# gnd! 38.4fF
C518 diff_1243200_708920# gnd! 38.4fF
C519 diff_2920040_640840# gnd! 713.2fF
C520 diff_1238760_646760# gnd! 894.7fF
C521 diff_3093200_531320# gnd! 1018.3fF
C522 diff_1238760_729640# gnd! 938.4fF
C523 diff_2828280_737040# gnd! 36.1fF
C524 diff_2803120_737040# gnd! 36.1fF
C525 diff_2777960_737040# gnd! 36.1fF
C526 diff_2752800_737040# gnd! 36.1fF
C527 diff_2727640_737040# gnd! 36.1fF
C528 diff_2702480_737040# gnd! 36.1fF
C529 diff_2677320_737040# gnd! 36.1fF
C530 diff_2652160_737040# gnd! 36.1fF
C531 diff_2627000_737040# gnd! 36.1fF
C532 diff_2601840_737040# gnd! 36.1fF
C533 diff_2576680_737040# gnd! 36.1fF
C534 diff_2551520_737040# gnd! 36.1fF
C535 diff_2526360_737040# gnd! 36.1fF
C536 diff_2501200_737040# gnd! 36.1fF
C537 diff_2476040_737040# gnd! 36.1fF
C538 diff_2450880_737040# gnd! 36.1fF
C539 diff_2425720_737040# gnd! 36.1fF
C540 diff_2400560_737040# gnd! 36.1fF
C541 diff_2375400_737040# gnd! 36.1fF
C542 diff_2350240_737040# gnd! 36.1fF
C543 diff_2325080_737040# gnd! 36.1fF
C544 diff_2299920_737040# gnd! 36.1fF
C545 diff_2274760_737040# gnd! 36.1fF
C546 diff_2249600_737040# gnd! 36.1fF
C547 diff_2224440_737040# gnd! 36.1fF
C548 diff_2199280_737040# gnd! 36.1fF
C549 diff_2174120_737040# gnd! 36.1fF
C550 diff_2148960_737040# gnd! 36.1fF
C551 diff_2123800_737040# gnd! 36.1fF
C552 diff_2098640_737040# gnd! 36.1fF
C553 diff_2073480_737040# gnd! 36.1fF
C554 diff_2048320_737040# gnd! 36.1fF
C555 diff_2023160_737040# gnd! 36.1fF
C556 diff_1998000_737040# gnd! 36.1fF
C557 diff_1972840_737040# gnd! 36.1fF
C558 diff_1947680_737040# gnd! 36.1fF
C559 diff_1922520_737040# gnd! 36.1fF
C560 diff_1897360_737040# gnd! 36.1fF
C561 diff_1872200_737040# gnd! 36.1fF
C562 diff_1847040_737040# gnd! 36.1fF
C563 diff_1821880_737040# gnd! 36.1fF
C564 diff_1796720_737040# gnd! 36.1fF
C565 diff_1771560_737040# gnd! 36.1fF
C566 diff_1746400_737040# gnd! 36.1fF
C567 diff_1721240_737040# gnd! 36.1fF
C568 diff_1696080_737040# gnd! 36.1fF
C569 diff_1670920_737040# gnd! 36.1fF
C570 diff_1645760_737040# gnd! 36.1fF
C571 diff_1620600_737040# gnd! 36.1fF
C572 diff_1595440_737040# gnd! 36.1fF
C573 diff_1570280_737040# gnd! 36.1fF
C574 diff_1545120_737040# gnd! 36.1fF
C575 diff_1519960_737040# gnd! 36.1fF
C576 diff_1494800_737040# gnd! 36.1fF
C577 diff_1469640_737040# gnd! 36.1fF
C578 diff_1444480_737040# gnd! 36.1fF
C579 diff_1419320_737040# gnd! 36.1fF
C580 diff_1394160_737040# gnd! 36.1fF
C581 diff_1369000_737040# gnd! 36.1fF
C582 diff_1343840_737040# gnd! 36.1fF
C583 diff_1318680_737040# gnd! 36.1fF
C584 diff_1293520_737040# gnd! 36.1fF
C585 diff_1268360_737040# gnd! 36.1fF
C586 diff_957560_602360# gnd! 158.1fF
C587 diff_852480_600880# gnd! 216.9fF
C588 diff_932400_560920# gnd! 154.5fF
C589 diff_1243200_737040# gnd! 36.1fF
C590 diff_856920_608280# gnd! 130.0fF
C591 diff_586080_617160# gnd! 22.2fF
C592 diff_498760_580160# gnd! 101.1fF
C593 diff_605320_617160# gnd! 75.9fF
C594 diff_590520_580160# gnd! 223.3fF
C595 diff_612720_606800# gnd! 536.3fF
C596 cm gnd! 1498.0fF
C597 diff_2920040_748880# gnd! 808.0fF
C598 diff_2828280_763680# gnd! 38.4fF
C599 diff_2803120_763680# gnd! 38.4fF
C600 diff_2777960_763680# gnd! 38.4fF
C601 diff_2752800_763680# gnd! 38.4fF
C602 diff_2727640_763680# gnd! 38.4fF
C603 diff_2702480_763680# gnd! 38.4fF
C604 diff_2677320_763680# gnd! 38.4fF
C605 diff_2652160_763680# gnd! 38.4fF
C606 diff_2627000_763680# gnd! 38.4fF
C607 diff_2601840_763680# gnd! 38.4fF
C608 diff_2576680_763680# gnd! 38.4fF
C609 diff_2551520_763680# gnd! 38.4fF
C610 diff_2526360_763680# gnd! 38.4fF
C611 diff_2501200_763680# gnd! 38.4fF
C612 diff_2476040_763680# gnd! 38.4fF
C613 diff_2450880_763680# gnd! 38.4fF
C614 diff_2425720_763680# gnd! 38.4fF
C615 diff_2400560_763680# gnd! 38.4fF
C616 diff_2375400_763680# gnd! 38.4fF
C617 diff_2350240_763680# gnd! 38.4fF
C618 diff_2325080_763680# gnd! 38.4fF
C619 diff_2299920_763680# gnd! 38.4fF
C620 diff_2274760_763680# gnd! 38.4fF
C621 diff_2249600_763680# gnd! 38.4fF
C622 diff_2224440_763680# gnd! 38.4fF
C623 diff_2199280_763680# gnd! 38.4fF
C624 diff_2174120_763680# gnd! 38.4fF
C625 diff_2148960_763680# gnd! 38.4fF
C626 diff_2123800_763680# gnd! 38.4fF
C627 diff_2098640_763680# gnd! 38.4fF
C628 diff_2073480_763680# gnd! 38.4fF
C629 diff_2048320_763680# gnd! 38.4fF
C630 diff_2023160_763680# gnd! 38.4fF
C631 diff_1998000_763680# gnd! 38.4fF
C632 diff_1972840_763680# gnd! 38.4fF
C633 diff_1947680_763680# gnd! 38.4fF
C634 diff_1922520_763680# gnd! 38.4fF
C635 diff_1897360_763680# gnd! 38.4fF
C636 diff_1872200_763680# gnd! 38.4fF
C637 diff_1847040_763680# gnd! 38.4fF
C638 diff_1821880_763680# gnd! 38.4fF
C639 diff_1796720_763680# gnd! 38.4fF
C640 diff_1771560_763680# gnd! 38.4fF
C641 diff_1746400_763680# gnd! 38.4fF
C642 diff_1721240_763680# gnd! 38.4fF
C643 diff_1696080_763680# gnd! 38.4fF
C644 diff_1670920_763680# gnd! 38.4fF
C645 diff_1645760_763680# gnd! 38.4fF
C646 diff_1620600_763680# gnd! 38.4fF
C647 diff_1595440_763680# gnd! 38.4fF
C648 diff_1570280_763680# gnd! 38.4fF
C649 diff_1545120_763680# gnd! 38.4fF
C650 diff_1519960_763680# gnd! 38.4fF
C651 diff_1494800_763680# gnd! 38.4fF
C652 diff_1469640_763680# gnd! 38.4fF
C653 diff_1444480_763680# gnd! 38.4fF
C654 diff_1419320_763680# gnd! 38.4fF
C655 diff_1394160_763680# gnd! 38.4fF
C656 diff_1369000_763680# gnd! 38.4fF
C657 diff_1343840_763680# gnd! 38.4fF
C658 diff_1318680_763680# gnd! 38.4fF
C659 diff_1293520_763680# gnd! 38.4fF
C660 diff_1268360_763680# gnd! 38.4fF
C661 diff_1243200_763680# gnd! 38.4fF
C662 diff_1238760_784400# gnd! 968.7fF
C663 diff_2828280_791800# gnd! 36.1fF
C664 diff_2803120_791800# gnd! 36.1fF
C665 diff_2777960_791800# gnd! 36.1fF
C666 diff_2752800_791800# gnd! 36.1fF
C667 diff_2727640_791800# gnd! 36.1fF
C668 diff_2702480_791800# gnd! 36.1fF
C669 diff_2677320_791800# gnd! 36.1fF
C670 diff_2652160_791800# gnd! 36.1fF
C671 diff_2627000_791800# gnd! 36.1fF
C672 diff_2601840_791800# gnd! 36.1fF
C673 diff_2576680_791800# gnd! 36.1fF
C674 diff_2551520_791800# gnd! 36.1fF
C675 diff_2526360_791800# gnd! 36.1fF
C676 diff_2501200_791800# gnd! 36.1fF
C677 diff_2476040_791800# gnd! 36.1fF
C678 diff_2450880_791800# gnd! 36.1fF
C679 diff_2425720_791800# gnd! 36.1fF
C680 diff_2400560_791800# gnd! 36.1fF
C681 diff_2375400_791800# gnd! 36.1fF
C682 diff_2350240_791800# gnd! 36.1fF
C683 diff_2325080_791800# gnd! 36.1fF
C684 diff_2299920_791800# gnd! 36.1fF
C685 diff_2274760_791800# gnd! 36.1fF
C686 diff_2249600_791800# gnd! 36.1fF
C687 diff_2224440_791800# gnd! 36.1fF
C688 diff_2199280_791800# gnd! 36.1fF
C689 diff_2174120_791800# gnd! 36.1fF
C690 diff_2148960_791800# gnd! 36.1fF
C691 diff_2123800_791800# gnd! 36.1fF
C692 diff_2098640_791800# gnd! 36.1fF
C693 diff_2073480_791800# gnd! 36.1fF
C694 diff_2048320_791800# gnd! 36.1fF
C695 diff_2023160_791800# gnd! 36.1fF
C696 diff_1998000_791800# gnd! 36.1fF
C697 diff_1972840_791800# gnd! 36.1fF
C698 diff_1947680_791800# gnd! 36.1fF
C699 diff_1922520_791800# gnd! 36.1fF
C700 diff_1897360_791800# gnd! 36.1fF
C701 diff_1872200_791800# gnd! 36.1fF
C702 diff_1847040_791800# gnd! 36.1fF
C703 diff_1821880_791800# gnd! 36.1fF
C704 diff_1796720_791800# gnd! 36.1fF
C705 diff_1771560_791800# gnd! 36.1fF
C706 diff_1746400_791800# gnd! 36.1fF
C707 diff_1721240_791800# gnd! 36.1fF
C708 diff_1696080_791800# gnd! 36.1fF
C709 diff_1670920_791800# gnd! 36.1fF
C710 diff_1645760_791800# gnd! 36.1fF
C711 diff_1620600_791800# gnd! 36.1fF
C712 diff_1595440_791800# gnd! 36.1fF
C713 diff_1570280_791800# gnd! 36.1fF
C714 diff_1545120_791800# gnd! 36.1fF
C715 diff_1519960_791800# gnd! 36.1fF
C716 diff_1494800_791800# gnd! 36.1fF
C717 diff_1469640_791800# gnd! 36.1fF
C718 diff_1444480_791800# gnd! 36.1fF
C719 diff_1419320_791800# gnd! 36.1fF
C720 diff_1394160_791800# gnd! 36.1fF
C721 diff_1369000_791800# gnd! 36.1fF
C722 diff_1343840_791800# gnd! 36.1fF
C723 diff_1318680_791800# gnd! 36.1fF
C724 diff_1293520_791800# gnd! 36.1fF
C725 diff_1268360_791800# gnd! 36.1fF
C726 diff_1243200_791800# gnd! 36.1fF
C727 diff_920560_771080# gnd! 355.1fF
C728 diff_1238760_811040# gnd! 985.6fF
C729 diff_2828280_818440# gnd! 38.4fF
C730 diff_2803120_818440# gnd! 38.4fF
C731 diff_2777960_818440# gnd! 38.4fF
C732 diff_2752800_818440# gnd! 38.4fF
C733 diff_2727640_818440# gnd! 38.4fF
C734 diff_2702480_818440# gnd! 38.4fF
C735 diff_2677320_818440# gnd! 38.4fF
C736 diff_2652160_818440# gnd! 38.4fF
C737 diff_2627000_818440# gnd! 38.4fF
C738 diff_2601840_818440# gnd! 38.4fF
C739 diff_2576680_818440# gnd! 38.4fF
C740 diff_2551520_818440# gnd! 38.4fF
C741 diff_2526360_818440# gnd! 38.4fF
C742 diff_2501200_818440# gnd! 38.4fF
C743 diff_2476040_818440# gnd! 38.4fF
C744 diff_2450880_818440# gnd! 38.4fF
C745 diff_2425720_818440# gnd! 38.4fF
C746 diff_2400560_818440# gnd! 38.4fF
C747 diff_2375400_818440# gnd! 38.4fF
C748 diff_2350240_818440# gnd! 38.4fF
C749 diff_2325080_818440# gnd! 38.4fF
C750 diff_2299920_818440# gnd! 38.4fF
C751 diff_2274760_818440# gnd! 38.4fF
C752 diff_2249600_818440# gnd! 38.4fF
C753 diff_2224440_818440# gnd! 38.4fF
C754 diff_2199280_818440# gnd! 38.4fF
C755 diff_2174120_818440# gnd! 38.4fF
C756 diff_2148960_818440# gnd! 38.4fF
C757 diff_2123800_818440# gnd! 38.4fF
C758 diff_2098640_818440# gnd! 38.4fF
C759 diff_2073480_818440# gnd! 38.4fF
C760 diff_2048320_818440# gnd! 38.4fF
C761 diff_2023160_818440# gnd! 38.4fF
C762 diff_1998000_818440# gnd! 38.4fF
C763 diff_1972840_818440# gnd! 38.4fF
C764 diff_1947680_818440# gnd! 38.4fF
C765 diff_1922520_818440# gnd! 38.4fF
C766 diff_1897360_818440# gnd! 38.4fF
C767 diff_1872200_818440# gnd! 38.4fF
C768 diff_1847040_818440# gnd! 38.4fF
C769 diff_1821880_818440# gnd! 38.4fF
C770 diff_1796720_818440# gnd! 38.4fF
C771 diff_1771560_818440# gnd! 38.4fF
C772 diff_1746400_818440# gnd! 38.4fF
C773 diff_1721240_818440# gnd! 38.4fF
C774 diff_1696080_818440# gnd! 38.4fF
C775 diff_1670920_818440# gnd! 38.4fF
C776 diff_1645760_818440# gnd! 38.4fF
C777 diff_1620600_818440# gnd! 38.4fF
C778 diff_1595440_818440# gnd! 38.4fF
C779 diff_1570280_818440# gnd! 38.4fF
C780 diff_1545120_818440# gnd! 38.4fF
C781 diff_1519960_818440# gnd! 38.4fF
C782 diff_1494800_818440# gnd! 38.4fF
C783 diff_1469640_818440# gnd! 38.4fF
C784 diff_1444480_818440# gnd! 38.4fF
C785 diff_1419320_818440# gnd! 38.4fF
C786 diff_1394160_818440# gnd! 38.4fF
C787 diff_1369000_818440# gnd! 38.4fF
C788 diff_1343840_818440# gnd! 38.4fF
C789 diff_1318680_818440# gnd! 38.4fF
C790 diff_1293520_818440# gnd! 38.4fF
C791 diff_1268360_818440# gnd! 38.4fF
C792 diff_1099640_809560# gnd! 15.4fF
C793 diff_1107040_787360# gnd! 184.8fF
C794 diff_1243200_818440# gnd! 38.4fF
C795 diff_1238760_756280# gnd! 902.5fF
C796 diff_1238760_839160# gnd! 939.9fF
C797 diff_2828280_846560# gnd! 36.1fF
C798 diff_2803120_846560# gnd! 36.1fF
C799 diff_2777960_846560# gnd! 36.1fF
C800 diff_2752800_846560# gnd! 36.1fF
C801 diff_2727640_846560# gnd! 36.1fF
C802 diff_2702480_846560# gnd! 36.1fF
C803 diff_2677320_846560# gnd! 36.1fF
C804 diff_2652160_846560# gnd! 36.1fF
C805 diff_2627000_846560# gnd! 36.1fF
C806 diff_2601840_846560# gnd! 36.1fF
C807 diff_2576680_846560# gnd! 36.1fF
C808 diff_2551520_846560# gnd! 36.1fF
C809 diff_2526360_846560# gnd! 36.1fF
C810 diff_2501200_846560# gnd! 36.1fF
C811 diff_2476040_846560# gnd! 36.1fF
C812 diff_2450880_846560# gnd! 36.1fF
C813 diff_2425720_846560# gnd! 36.1fF
C814 diff_2400560_846560# gnd! 36.1fF
C815 diff_2375400_846560# gnd! 36.1fF
C816 diff_2350240_846560# gnd! 36.1fF
C817 diff_2325080_846560# gnd! 36.1fF
C818 diff_2299920_846560# gnd! 36.1fF
C819 diff_2274760_846560# gnd! 36.1fF
C820 diff_2249600_846560# gnd! 36.1fF
C821 diff_2224440_846560# gnd! 36.1fF
C822 diff_2199280_846560# gnd! 36.1fF
C823 diff_2174120_846560# gnd! 36.1fF
C824 diff_2148960_846560# gnd! 36.1fF
C825 diff_2123800_846560# gnd! 36.1fF
C826 diff_2098640_846560# gnd! 36.1fF
C827 diff_2073480_846560# gnd! 36.1fF
C828 diff_2048320_846560# gnd! 36.1fF
C829 diff_2023160_846560# gnd! 36.1fF
C830 diff_1998000_846560# gnd! 36.1fF
C831 diff_1972840_846560# gnd! 36.1fF
C832 diff_1947680_846560# gnd! 36.1fF
C833 diff_1922520_846560# gnd! 36.1fF
C834 diff_1897360_846560# gnd! 36.1fF
C835 diff_1872200_846560# gnd! 36.1fF
C836 diff_1847040_846560# gnd! 36.1fF
C837 diff_1821880_846560# gnd! 36.1fF
C838 diff_1796720_846560# gnd! 36.1fF
C839 diff_1771560_846560# gnd! 36.1fF
C840 diff_1746400_846560# gnd! 36.1fF
C841 diff_1721240_846560# gnd! 36.1fF
C842 diff_1696080_846560# gnd! 36.1fF
C843 diff_1670920_846560# gnd! 36.1fF
C844 diff_1645760_846560# gnd! 36.1fF
C845 diff_1620600_846560# gnd! 36.1fF
C846 diff_1595440_846560# gnd! 36.1fF
C847 diff_1570280_846560# gnd! 36.1fF
C848 diff_1545120_846560# gnd! 36.1fF
C849 diff_1519960_846560# gnd! 36.1fF
C850 diff_1494800_846560# gnd! 36.1fF
C851 diff_1469640_846560# gnd! 36.1fF
C852 diff_1444480_846560# gnd! 36.1fF
C853 diff_1419320_846560# gnd! 36.1fF
C854 diff_1394160_846560# gnd! 36.1fF
C855 diff_1369000_846560# gnd! 36.1fF
C856 diff_1343840_846560# gnd! 36.1fF
C857 diff_1318680_846560# gnd! 36.1fF
C858 diff_1293520_846560# gnd! 36.1fF
C859 diff_1268360_846560# gnd! 36.1fF
C860 diff_1243200_846560# gnd! 36.1fF
C861 diff_2920040_858400# gnd! 710.9fF
C862 diff_2828280_873200# gnd! 38.4fF
C863 diff_2803120_873200# gnd! 38.4fF
C864 diff_2777960_873200# gnd! 38.4fF
C865 diff_2752800_873200# gnd! 38.4fF
C866 diff_2727640_873200# gnd! 38.4fF
C867 diff_2702480_873200# gnd! 38.4fF
C868 diff_2677320_873200# gnd! 38.4fF
C869 diff_2652160_873200# gnd! 38.4fF
C870 diff_2627000_873200# gnd! 38.4fF
C871 diff_2601840_873200# gnd! 38.4fF
C872 diff_2576680_873200# gnd! 38.4fF
C873 diff_2551520_873200# gnd! 38.4fF
C874 diff_2526360_873200# gnd! 38.4fF
C875 diff_2501200_873200# gnd! 38.4fF
C876 diff_2476040_873200# gnd! 38.4fF
C877 diff_2450880_873200# gnd! 38.4fF
C878 diff_2425720_873200# gnd! 38.4fF
C879 diff_2400560_873200# gnd! 38.4fF
C880 diff_2375400_873200# gnd! 38.4fF
C881 diff_2350240_873200# gnd! 38.4fF
C882 diff_2325080_873200# gnd! 38.4fF
C883 diff_2299920_873200# gnd! 38.4fF
C884 diff_2274760_873200# gnd! 38.4fF
C885 diff_2249600_873200# gnd! 38.4fF
C886 diff_2224440_873200# gnd! 38.4fF
C887 diff_2199280_873200# gnd! 38.4fF
C888 diff_2174120_873200# gnd! 38.4fF
C889 diff_2148960_873200# gnd! 38.4fF
C890 diff_2123800_873200# gnd! 38.4fF
C891 diff_2098640_873200# gnd! 38.4fF
C892 diff_2073480_873200# gnd! 38.4fF
C893 diff_2048320_873200# gnd! 38.4fF
C894 diff_2023160_873200# gnd! 38.4fF
C895 diff_1998000_873200# gnd! 38.4fF
C896 diff_1972840_873200# gnd! 38.4fF
C897 diff_1947680_873200# gnd! 38.4fF
C898 diff_1922520_873200# gnd! 38.4fF
C899 diff_1897360_873200# gnd! 38.4fF
C900 diff_1872200_873200# gnd! 38.4fF
C901 diff_1847040_873200# gnd! 38.4fF
C902 diff_1821880_873200# gnd! 38.4fF
C903 diff_1796720_873200# gnd! 38.4fF
C904 diff_1771560_873200# gnd! 38.4fF
C905 diff_1746400_873200# gnd! 38.4fF
C906 diff_1721240_873200# gnd! 38.4fF
C907 diff_1696080_873200# gnd! 38.4fF
C908 diff_1670920_873200# gnd! 38.4fF
C909 diff_1645760_873200# gnd! 38.4fF
C910 diff_1620600_873200# gnd! 38.4fF
C911 diff_1595440_873200# gnd! 38.4fF
C912 diff_1570280_873200# gnd! 38.4fF
C913 diff_1545120_873200# gnd! 38.4fF
C914 diff_1519960_873200# gnd! 38.4fF
C915 diff_1494800_873200# gnd! 38.4fF
C916 diff_1469640_873200# gnd! 38.4fF
C917 diff_1444480_873200# gnd! 38.4fF
C918 diff_1419320_873200# gnd! 38.4fF
C919 diff_1394160_873200# gnd! 38.4fF
C920 diff_1369000_873200# gnd! 38.4fF
C921 diff_1343840_873200# gnd! 38.4fF
C922 diff_1318680_873200# gnd! 38.4fF
C923 diff_1293520_873200# gnd! 38.4fF
C924 diff_1268360_873200# gnd! 38.4fF
C925 diff_1115920_809560# gnd! 116.2fF
C926 diff_1243200_873200# gnd! 38.4fF
C927 diff_1238760_893920# gnd! 966.5fF
C928 diff_2828280_901320# gnd! 36.1fF
C929 diff_2803120_901320# gnd! 36.1fF
C930 diff_2777960_901320# gnd! 36.1fF
C931 diff_2752800_901320# gnd! 36.1fF
C932 diff_2727640_901320# gnd! 36.1fF
C933 diff_2702480_901320# gnd! 36.1fF
C934 diff_2677320_901320# gnd! 36.1fF
C935 diff_2652160_901320# gnd! 36.1fF
C936 diff_2627000_901320# gnd! 36.1fF
C937 diff_2601840_901320# gnd! 36.1fF
C938 diff_2576680_901320# gnd! 36.1fF
C939 diff_2551520_901320# gnd! 36.1fF
C940 diff_2526360_901320# gnd! 36.1fF
C941 diff_2501200_901320# gnd! 36.1fF
C942 diff_2476040_901320# gnd! 36.1fF
C943 diff_2450880_901320# gnd! 36.1fF
C944 diff_2425720_901320# gnd! 36.1fF
C945 diff_2400560_901320# gnd! 36.1fF
C946 diff_2375400_901320# gnd! 36.1fF
C947 diff_2350240_901320# gnd! 36.1fF
C948 diff_2325080_901320# gnd! 36.1fF
C949 diff_2299920_901320# gnd! 36.1fF
C950 diff_2274760_901320# gnd! 36.1fF
C951 diff_2249600_901320# gnd! 36.1fF
C952 diff_2224440_901320# gnd! 36.1fF
C953 diff_2199280_901320# gnd! 36.1fF
C954 diff_2174120_901320# gnd! 36.1fF
C955 diff_2148960_901320# gnd! 36.1fF
C956 diff_2123800_901320# gnd! 36.1fF
C957 diff_2098640_901320# gnd! 36.1fF
C958 diff_2073480_901320# gnd! 36.1fF
C959 diff_2048320_901320# gnd! 36.1fF
C960 diff_2023160_901320# gnd! 36.1fF
C961 diff_1998000_901320# gnd! 36.1fF
C962 diff_1972840_901320# gnd! 36.1fF
C963 diff_1947680_901320# gnd! 36.1fF
C964 diff_1922520_901320# gnd! 36.1fF
C965 diff_1897360_901320# gnd! 36.1fF
C966 diff_1872200_901320# gnd! 36.1fF
C967 diff_1847040_901320# gnd! 36.1fF
C968 diff_1821880_901320# gnd! 36.1fF
C969 diff_1796720_901320# gnd! 36.1fF
C970 diff_1771560_901320# gnd! 36.1fF
C971 diff_1746400_901320# gnd! 36.1fF
C972 diff_1721240_901320# gnd! 36.1fF
C973 diff_1696080_901320# gnd! 36.1fF
C974 diff_1670920_901320# gnd! 36.1fF
C975 diff_1645760_901320# gnd! 36.1fF
C976 diff_1620600_901320# gnd! 36.1fF
C977 diff_1595440_901320# gnd! 36.1fF
C978 diff_1570280_901320# gnd! 36.1fF
C979 diff_1545120_901320# gnd! 36.1fF
C980 diff_1519960_901320# gnd! 36.1fF
C981 diff_1494800_901320# gnd! 36.1fF
C982 diff_1469640_901320# gnd! 36.1fF
C983 diff_1444480_901320# gnd! 36.1fF
C984 diff_1419320_901320# gnd! 36.1fF
C985 diff_1394160_901320# gnd! 36.1fF
C986 diff_1369000_901320# gnd! 36.1fF
C987 diff_1343840_901320# gnd! 36.1fF
C988 diff_1318680_901320# gnd! 36.1fF
C989 diff_1293520_901320# gnd! 36.1fF
C990 diff_1268360_901320# gnd! 36.1fF
C991 diff_1243200_901320# gnd! 36.1fF
C992 diff_1238760_920560# gnd! 985.6fF
C993 diff_2828280_927960# gnd! 38.4fF
C994 diff_2803120_927960# gnd! 38.4fF
C995 diff_2777960_927960# gnd! 38.4fF
C996 diff_2752800_927960# gnd! 38.4fF
C997 diff_2727640_927960# gnd! 38.4fF
C998 diff_2702480_927960# gnd! 38.4fF
C999 diff_2677320_927960# gnd! 38.4fF
C1000 diff_2652160_927960# gnd! 38.4fF
C1001 diff_2627000_927960# gnd! 38.4fF
C1002 diff_2601840_927960# gnd! 38.4fF
C1003 diff_2576680_927960# gnd! 38.4fF
C1004 diff_2551520_927960# gnd! 38.4fF
C1005 diff_2526360_927960# gnd! 38.4fF
C1006 diff_2501200_927960# gnd! 38.4fF
C1007 diff_2476040_927960# gnd! 38.4fF
C1008 diff_2450880_927960# gnd! 38.4fF
C1009 diff_2425720_927960# gnd! 38.4fF
C1010 diff_2400560_927960# gnd! 38.4fF
C1011 diff_2375400_927960# gnd! 38.4fF
C1012 diff_2350240_927960# gnd! 38.4fF
C1013 diff_2325080_927960# gnd! 38.4fF
C1014 diff_2299920_927960# gnd! 38.4fF
C1015 diff_2274760_927960# gnd! 38.4fF
C1016 diff_2249600_927960# gnd! 38.4fF
C1017 diff_2224440_927960# gnd! 38.4fF
C1018 diff_2199280_927960# gnd! 38.4fF
C1019 diff_2174120_927960# gnd! 38.4fF
C1020 diff_2148960_927960# gnd! 38.4fF
C1021 diff_2123800_927960# gnd! 38.4fF
C1022 diff_2098640_927960# gnd! 38.4fF
C1023 diff_2073480_927960# gnd! 38.4fF
C1024 diff_2048320_927960# gnd! 38.4fF
C1025 diff_2023160_927960# gnd! 38.4fF
C1026 diff_1998000_927960# gnd! 38.4fF
C1027 diff_1972840_927960# gnd! 38.4fF
C1028 diff_1947680_927960# gnd! 38.4fF
C1029 diff_1922520_927960# gnd! 38.4fF
C1030 diff_1897360_927960# gnd! 38.4fF
C1031 diff_1872200_927960# gnd! 38.4fF
C1032 diff_1847040_927960# gnd! 38.4fF
C1033 diff_1821880_927960# gnd! 38.4fF
C1034 diff_1796720_927960# gnd! 38.4fF
C1035 diff_1771560_927960# gnd! 38.4fF
C1036 diff_1746400_927960# gnd! 38.4fF
C1037 diff_1721240_927960# gnd! 38.4fF
C1038 diff_1696080_927960# gnd! 38.4fF
C1039 diff_1670920_927960# gnd! 38.4fF
C1040 diff_1645760_927960# gnd! 38.4fF
C1041 diff_1620600_927960# gnd! 38.4fF
C1042 diff_1595440_927960# gnd! 38.4fF
C1043 diff_1570280_927960# gnd! 38.4fF
C1044 diff_1545120_927960# gnd! 38.4fF
C1045 diff_1519960_927960# gnd! 38.4fF
C1046 diff_1494800_927960# gnd! 38.4fF
C1047 diff_1469640_927960# gnd! 38.4fF
C1048 diff_1444480_927960# gnd! 38.4fF
C1049 diff_1419320_927960# gnd! 38.4fF
C1050 diff_1394160_927960# gnd! 38.4fF
C1051 diff_1369000_927960# gnd! 38.4fF
C1052 diff_1343840_927960# gnd! 38.4fF
C1053 diff_1318680_927960# gnd! 38.4fF
C1054 diff_1293520_927960# gnd! 38.4fF
C1055 diff_1268360_927960# gnd! 38.4fF
C1056 diff_1243200_927960# gnd! 38.4fF
C1057 diff_1068560_852480# gnd! 144.7fF
C1058 diff_1036000_463240# gnd! 317.1fF
C1059 diff_1238760_865800# gnd! 906.6fF
C1060 diff_3119840_1102600# gnd! 162.0fF
C1061 diff_3377360_1142560# gnd! 135.5fF
C1062 diff_3119840_1129240# gnd! 160.4fF
C1063 diff_3492800_1302400# gnd! 429.4fF
C1064 diff_3492800_1326080# gnd! 110.9fF
C1065 diff_3421760_1235800# gnd! 276.2fF
C1066 diff_3377360_1189920# gnd! 136.8fF
C1067 diff_3534240_1386760# gnd! 73.0fF
C1068 diff_3421760_1283160# gnd! 271.7fF
C1069 diff_3121320_1194360# gnd! 152.7fF
C1070 diff_3121320_1222480# gnd! 165.1fF
C1071 diff_3121320_1277240# gnd! 157.4fF
C1072 diff_3377360_1329040# gnd! 127.9fF
C1073 diff_3121320_1305360# gnd! 156.3fF
C1074 diff_3122800_1370480# gnd! 153.0fF
C1075 diff_3421760_1422280# gnd! 155.2fF
C1076 diff_3377360_1374920# gnd! 126.7fF
C1077 diff_3121320_1397120# gnd! 163.8fF
C1078 diff_3476520_1401560# gnd! 220.2fF
C1079 diff_3504640_1514040# gnd! 61.8fF
C1080 diff_3421760_1466680# gnd! 245.6fF
C1081 diff_3476520_1593960# gnd! 63.8fF
C1082 diff_3121320_1453360# gnd! 171.3fF
C1083 diff_3377360_1515520# gnd! 134.4fF
C1084 diff_3121320_1481480# gnd! 161.0fF
C1085 diff_1238760_948680# gnd! 939.9fF
C1086 diff_1115920_948680# gnd! 190.8fF
C1087 diff_350760_574240# gnd! 88.1fF
C1088 diff_417360_463240# gnd! 648.9fF
C1089 reset gnd! 1123.0fF
C1090 diff_592000_757760# gnd! 137.9fF
C1091 diff_614200_882080# gnd! 74.8fF
C1092 diff_856920_939800# gnd! 203.5fF
C1093 diff_2828280_956080# gnd! 61.6fF
C1094 diff_2803120_956080# gnd! 62.5fF
C1095 diff_2727640_956080# gnd! 61.6fF
C1096 diff_2702480_956080# gnd! 62.5fF
C1097 diff_2627000_956080# gnd! 61.6fF
C1098 diff_2601840_956080# gnd! 62.5fF
C1099 diff_2526360_956080# gnd! 61.6fF
C1100 diff_2501200_956080# gnd! 62.5fF
C1101 diff_2425720_956080# gnd! 61.6fF
C1102 diff_2400560_956080# gnd! 62.5fF
C1103 diff_2325080_956080# gnd! 61.6fF
C1104 diff_2299920_956080# gnd! 62.5fF
C1105 diff_2224440_956080# gnd! 61.6fF
C1106 diff_2199280_956080# gnd! 62.5fF
C1107 diff_2123800_956080# gnd! 61.6fF
C1108 diff_2098640_956080# gnd! 62.5fF
C1109 diff_2023160_956080# gnd! 61.6fF
C1110 diff_1998000_956080# gnd! 62.5fF
C1111 diff_1922520_956080# gnd! 61.6fF
C1112 diff_1897360_956080# gnd! 62.5fF
C1113 diff_1821880_956080# gnd! 61.6fF
C1114 diff_1796720_956080# gnd! 62.5fF
C1115 diff_1721240_956080# gnd! 61.6fF
C1116 diff_1696080_956080# gnd! 62.5fF
C1117 diff_1620600_956080# gnd! 61.6fF
C1118 diff_1595440_956080# gnd! 62.5fF
C1119 diff_1519960_956080# gnd! 61.6fF
C1120 diff_1494800_956080# gnd! 62.5fF
C1121 diff_1419320_956080# gnd! 61.6fF
C1122 diff_1394160_956080# gnd! 62.5fF
C1123 diff_1318680_956080# gnd! 60.0fF
C1124 diff_1293520_956080# gnd! 61.2fF
C1125 diff_1006400_970880# gnd! 20.8fF
C1126 diff_858400_964960# gnd! 103.4fF
C1127 diff_864320_837680# gnd! 220.8fF
C1128 diff_856920_686720# gnd! 398.0fF
C1129 diff_1133680_519480# gnd! 796.6fF
C1130 diff_1018240_964960# gnd! 248.3fF
C1131 diff_3421760_1613200# gnd! 171.0fF
C1132 diff_3377360_1571760# gnd! 132.0fF
C1133 diff_3115400_1533280# gnd! 213.5fF
C1134 diff_3167200_1580640# gnd! 132.3fF
C1135 diff_3340360_1716800# gnd! 54.1fF
C1136 diff_3213080_1693120# gnd! 135.8fF
C1137 diff_3208640_1687200# gnd! 145.1fF
C1138 diff_3239720_1740480# gnd! 134.4fF
C1139 diff_3358120_1041920# gnd! 550.1fF
C1140 diff_3412880_1796720# gnd! 73.9fF
C1141 diff_3193840_1805600# gnd! 118.4fF
C1142 diff_3469120_1398600# gnd! 454.4fF
C1143 diff_3414360_1847040# gnd! 74.1fF
C1144 diff_3414360_1900320# gnd! 72.1fF
C1145 diff_2777960_956080# gnd! 79.5fF
C1146 diff_2752800_956080# gnd! 79.4fF
C1147 diff_2785360_1047840# gnd! 62.0fF
C1148 diff_2677320_956080# gnd! 79.5fF
C1149 diff_2652160_956080# gnd! 79.4fF
C1150 diff_2684720_1047840# gnd! 62.0fF
C1151 diff_2576680_956080# gnd! 79.5fF
C1152 diff_2551520_956080# gnd! 79.4fF
C1153 diff_2584080_1047840# gnd! 62.0fF
C1154 diff_2476040_956080# gnd! 79.5fF
C1155 diff_2450880_956080# gnd! 79.4fF
C1156 diff_2483440_1047840# gnd! 62.0fF
C1157 diff_2375400_956080# gnd! 79.5fF
C1158 diff_2350240_956080# gnd! 79.4fF
C1159 diff_2382800_1047840# gnd! 62.0fF
C1160 diff_2274760_956080# gnd! 79.5fF
C1161 diff_2249600_956080# gnd! 79.4fF
C1162 diff_2282160_1047840# gnd! 62.0fF
C1163 diff_2174120_956080# gnd! 79.5fF
C1164 diff_2148960_956080# gnd! 79.4fF
C1165 diff_2181520_1047840# gnd! 62.0fF
C1166 diff_2073480_956080# gnd! 79.5fF
C1167 diff_2048320_956080# gnd! 79.4fF
C1168 diff_2080880_1047840# gnd! 62.0fF
C1169 diff_1972840_956080# gnd! 79.5fF
C1170 diff_1947680_956080# gnd! 79.4fF
C1171 diff_1980240_1047840# gnd! 62.0fF
C1172 diff_1872200_956080# gnd! 79.5fF
C1173 diff_1847040_956080# gnd! 79.4fF
C1174 diff_1879600_1047840# gnd! 62.0fF
C1175 diff_1771560_956080# gnd! 79.5fF
C1176 diff_1746400_956080# gnd! 79.4fF
C1177 diff_1778960_1047840# gnd! 62.0fF
C1178 diff_1670920_956080# gnd! 79.5fF
C1179 diff_1645760_956080# gnd! 79.4fF
C1180 diff_1678320_1047840# gnd! 62.0fF
C1181 diff_1570280_956080# gnd! 79.5fF
C1182 diff_1545120_956080# gnd! 79.4fF
C1183 diff_1577680_1047840# gnd! 62.0fF
C1184 diff_1469640_956080# gnd! 79.5fF
C1185 diff_1444480_956080# gnd! 79.4fF
C1186 diff_1477040_1047840# gnd! 62.0fF
C1187 diff_1369000_956080# gnd! 79.5fF
C1188 diff_1343840_956080# gnd! 79.4fF
C1189 diff_1376400_1047840# gnd! 62.0fF
C1190 diff_688200_944240# gnd! 201.3fF
C1191 diff_519480_898360# gnd! 147.1fF
C1192 diff_661560_957560# gnd! 188.2fF
C1193 diff_418840_657120# gnd! 588.5fF
C1194 diff_504680_587560# gnd! 315.7fF
C1195 diff_1243200_956080# gnd! 71.6fF
C1196 diff_1274280_1049320# gnd! 68.1fF
C1197 diff_1263920_1047840# gnd! 83.0fF
C1198 diff_1229880_1031560# gnd! 151.7fF
C1199 diff_2735040_1022680# gnd! 161.7fF
C1200 diff_2533760_1022680# gnd! 165.1fF
C1201 diff_2332480_1022680# gnd! 165.1fF
C1202 diff_2131200_1022680# gnd! 165.3fF
C1203 diff_1929920_1022680# gnd! 158.9fF
C1204 diff_1728640_1022680# gnd! 158.9fF
C1205 diff_1527360_1022680# gnd! 168.2fF
C1206 diff_1326080_1019720# gnd! 166.0fF
C1207 diff_2634400_1022680# gnd! 169.1fF
C1208 diff_2786840_1118880# gnd! 180.8fF
C1209 diff_2433120_1022680# gnd! 169.1fF
C1210 diff_2684720_1118880# gnd! 188.0fF
C1211 diff_2584080_1118880# gnd! 184.8fF
C1212 diff_2483440_1118880# gnd! 188.0fF
C1213 diff_2231840_1022680# gnd! 169.5fF
C1214 diff_2382800_1118880# gnd! 184.8fF
C1215 diff_2283640_1118880# gnd! 188.0fF
C1216 diff_2030560_1022680# gnd! 163.3fF
C1217 diff_2183000_1118880# gnd! 184.8fF
C1218 diff_2080880_1120360# gnd! 182.0fF
C1219 diff_1829280_1022680# gnd! 162.6fF
C1220 diff_1980240_1120360# gnd! 178.8fF
C1221 diff_1879600_1120360# gnd! 182.0fF
C1222 diff_1628000_1022680# gnd! 173.3fF
C1223 diff_1778960_1120360# gnd! 178.8fF
C1224 diff_1426720_1022680# gnd! 169.1fF
C1225 diff_1576200_1117400# gnd! 190.8fF
C1226 diff_1477040_1118880# gnd! 188.0fF
C1227 diff_1278720_1114440# gnd! 183.8fF
C1228 diff_1676840_1117400# gnd! 192.0fF
C1229 diff_1376400_1118880# gnd! 185.3fF
C1230 diff_2735040_1144040# gnd! 165.2fF
C1231 diff_2632920_1144040# gnd! 167.9fF
C1232 diff_2532280_1144040# gnd! 167.0fF
C1233 diff_2431640_1144040# gnd! 167.9fF
C1234 diff_2331000_1144040# gnd! 167.0fF
C1235 diff_2231840_1144040# gnd! 167.9fF
C1236 diff_2131200_1144040# gnd! 167.0fF
C1237 diff_2029080_1145520# gnd! 161.9fF
C1238 diff_1928440_1145520# gnd! 161.0fF
C1239 diff_1827800_1145520# gnd! 161.9fF
C1240 diff_1727160_1145520# gnd! 161.0fF
C1241 diff_1625040_1142560# gnd! 172.6fF
C1242 diff_1524400_1142560# gnd! 173.0fF
C1243 diff_552040_951640# gnd! 117.3fF
C1244 diff_612720_984200# gnd! 203.5fF
C1245 diff_1108520_1095200# gnd! 164.2fF
C1246 diff_1425240_1144040# gnd! 167.9fF
C1247 diff_1324600_1144040# gnd! 167.0fF
C1248 diff_2835680_1022680# gnd! 201.3fF
C1249 diff_2536720_1118880# gnd! 382.6fF
C1250 diff_2335440_1118880# gnd! 383.3fF
C1251 diff_2135640_1118880# gnd! 384.2fF
C1252 diff_1932880_1118880# gnd! 391.1fF
C1253 diff_1731600_1118880# gnd! 389.2fF
C1254 diff_1528840_1118880# gnd! 369.7fF
C1255 diff_1329040_1118880# gnd! 380.4fF
C1256 diff_1232840_1105560# gnd! 464.9fF
C1257 diff_2739480_1118880# gnd! 391.3fF
C1258 diff_2637360_1120360# gnd! 426.3fF
C1259 diff_2436080_1120360# gnd! 423.8fF
C1260 diff_2236280_1120360# gnd! 427.5fF
C1261 diff_2033520_1120360# gnd! 426.5fF
C1262 diff_1832240_1118880# gnd! 432.7fF
C1263 diff_1629480_1115920# gnd! 420.7fF
C1264 diff_1429680_1120360# gnd! 416.9fF
C1265 diff_1386760_1188440# gnd! 1142.5fF
C1266 diff_988640_1095200# gnd! 162.6fF
C1267 diff_593480_988640# gnd! 224.6fF
C1268 diff_797720_1095200# gnd! 164.2fF
C1269 diff_507640_1052280# gnd! 90.3fF
C1270 diff_700040_1055240# gnd! 151.5fF
C1271 diff_1250600_1186960# gnd! 1243.9fF
C1272 diff_2462720_1243200# gnd! 442.1fF
C1273 diff_2060160_1243200# gnd! 494.7fF
C1274 diff_769600_586080# gnd! 1071.7fF
C1275 diff_1657600_1243200# gnd! 433.2fF
C1276 diff_1232840_1340880# gnd! 397.9fF
C1277 diff_609760_1096680# gnd! 162.6fF
C1278 diff_1022680_1281680# gnd! 586.1fF
C1279 diff_990120_1192880# gnd! 190.3fF
C1280 diff_1192880_1336440# gnd! 159.3fF
C1281 diff_1111480_1194360# gnd! 283.2fF
C1282 diff_2664000_1215080# gnd! 698.5fF
C1283 diff_2462720_1213600# gnd! 830.0fF
C1284 diff_695600_586080# gnd! 1279.2fF
C1285 diff_2262920_1213600# gnd! 787.5fF
C1286 diff_2060160_1213600# gnd! 790.8fF
C1287 diff_1858880_1213600# gnd! 854.7fF
C1288 diff_1656120_1383800# gnd! 814.6fF
C1289 diff_1456320_1215080# gnd! 752.8fF
C1290 diff_507640_1070040# gnd! 1019.9fF
C1291 diff_842120_1275760# gnd! 613.5fF
C1292 diff_799200_1192880# gnd! 175.7fF
C1293 diff_670440_1255040# gnd! 713.5fF
C1294 diff_612720_1192880# gnd! 164.4fF
C1295 io0 gnd! 2145.5fF
C1296 diff_550560_1112960# gnd! 676.8fF
C1297 diff_501720_853960# gnd! 760.7fF
C1298 io1 gnd! 2391.3fF
C1299 io2 gnd! 2923.7fF
C1300 io3 gnd! 2757.9fF
C1301 diff_1253560_1194360# gnd! 793.5fF
C1302 diff_1247640_1422280# gnd! 1208.1fF
C1303 diff_990120_1340880# gnd! 331.1fF
C1304 diff_799200_1340880# gnd! 330.2fF
C1305 diff_608280_1340880# gnd! 322.0fF
C1306 diff_415880_1340880# gnd! 322.4fF
C1307 diff_1311280_1160320# gnd! 1751.2fF
C1308 diff_1274280_1133680# gnd! 1903.8fF
C1309 diff_1226920_1511080# gnd! 1863.5fF
C1310 diff_2739480_1487400# gnd! 397.7fF
C1311 diff_2785360_1561400# gnd! 61.6fF
C1312 diff_2637360_1488880# gnd! 435.0fF
C1313 diff_2735040_1456320# gnd! 154.9fF
C1314 diff_2684720_1561400# gnd! 61.6fF
C1315 diff_2536720_1488880# gnd! 380.5fF
C1316 diff_2632920_1456320# gnd! 157.1fF
C1317 diff_2584080_1561400# gnd! 61.6fF
C1318 diff_2436080_1488880# gnd! 430.7fF
C1319 diff_2532280_1456320# gnd! 156.5fF
C1320 diff_2483440_1561400# gnd! 61.6fF
C1321 diff_2335440_1488880# gnd! 380.5fF
C1322 diff_2431640_1456320# gnd! 157.1fF
C1323 diff_2382800_1561400# gnd! 61.6fF
C1324 diff_2236280_1488880# gnd! 428.3fF
C1325 diff_2331000_1456320# gnd! 156.5fF
C1326 diff_2282160_1561400# gnd! 61.6fF
C1327 diff_2135640_1488880# gnd! 381.2fF
C1328 diff_2231840_1456320# gnd! 157.1fF
C1329 diff_2181520_1561400# gnd! 61.6fF
C1330 diff_2033520_1487400# gnd! 431.6fF
C1331 diff_2131200_1456320# gnd! 156.5fF
C1332 diff_2080880_1561400# gnd! 61.6fF
C1333 diff_1932880_1487400# gnd! 389.6fF
C1334 diff_2029080_1456320# gnd! 151.1fF
C1335 diff_1980240_1561400# gnd! 61.6fF
C1336 diff_1832240_1487400# gnd! 437.5fF
C1337 diff_1928440_1456320# gnd! 150.5fF
C1338 diff_1879600_1561400# gnd! 61.6fF
C1339 diff_1731600_1487400# gnd! 389.6fF
C1340 diff_1827800_1456320# gnd! 151.1fF
C1341 diff_1778960_1561400# gnd! 61.6fF
C1342 diff_1629480_1490360# gnd! 428.3fF
C1343 diff_1727160_1456320# gnd! 150.5fF
C1344 diff_1678320_1561400# gnd! 61.6fF
C1345 diff_1528840_1490360# gnd! 369.1fF
C1346 diff_1625040_1456320# gnd! 158.6fF
C1347 diff_1577680_1561400# gnd! 61.6fF
C1348 diff_1429680_1488880# gnd! 421.4fF
C1349 diff_1524400_1456320# gnd! 162.5fF
C1350 diff_1477040_1561400# gnd! 61.6fF
C1351 diff_1329040_1488880# gnd! 380.9fF
C1352 diff_1425240_1456320# gnd! 157.1fF
C1353 diff_1376400_1561400# gnd! 61.6fF
C1354 diff_1324600_1456320# gnd! 156.5fF
C1355 diff_1232840_1500720# gnd! 462.0fF
C1356 diff_1274280_1562880# gnd! 69.0fF
C1357 diff_1293520_1043400# gnd! 716.3fF
C1358 diff_2835680_1583600# gnd! 193.2fF
C1359 diff_2786840_1482960# gnd! 173.4fF
C1360 diff_2735040_1583600# gnd! 151.5fF
C1361 diff_2684720_1482960# gnd! 180.6fF
C1362 diff_2634400_1583600# gnd! 159.9fF
C1363 diff_2584080_1482960# gnd! 177.2fF
C1364 diff_2533760_1583600# gnd! 154.7fF
C1365 diff_2483440_1482960# gnd! 180.6fF
C1366 diff_2433120_1583600# gnd! 159.9fF
C1367 diff_2382800_1482960# gnd! 177.2fF
C1368 diff_2332480_1583600# gnd! 154.7fF
C1369 diff_2283640_1482960# gnd! 180.6fF
C1370 diff_2231840_1583600# gnd! 160.4fF
C1371 diff_2183000_1482960# gnd! 177.2fF
C1372 diff_2131200_1583600# gnd! 154.9fF
C1373 diff_2080880_1482960# gnd! 174.6fF
C1374 diff_2030560_1583600# gnd! 154.2fF
C1375 diff_1980240_1482960# gnd! 171.2fF
C1376 diff_1929920_1583600# gnd! 148.5fF
C1377 diff_1879600_1482960# gnd! 174.6fF
C1378 diff_1829280_1583600# gnd! 153.0fF
C1379 diff_1778960_1482960# gnd! 171.2fF
C1380 diff_1728640_1583600# gnd! 148.5fF
C1381 diff_1676840_1481480# gnd! 187.1fF
C1382 diff_1628000_1583600# gnd! 164.3fF
C1383 diff_1576200_1482960# gnd! 183.2fF
C1384 diff_1527360_1583600# gnd! 157.8fF
C1385 diff_1477040_1482960# gnd! 180.6fF
C1386 diff_1426720_1583600# gnd! 160.5fF
C1387 diff_1376400_1481480# gnd! 177.7fF
C1388 diff_1326080_1583600# gnd! 155.6fF
C1389 diff_1278720_1482960# gnd! 176.4fF
C1390 diff_1386760_1422280# gnd! 1187.0fF
C1391 diff_321160_969400# gnd! 877.4fF
C1392 cl gnd! 1854.2fF
C1393 diff_1229880_1524400# gnd! 144.4fF
C1394 diff_1012320_1602840# gnd! 304.1fF
C1395 diff_1154400_1582120# gnd! 37.0fF ;**FLOATING
C1396 diff_821400_1602840# gnd! 299.4fF
C1397 diff_988640_1443000# gnd! 463.9fF
C1398 diff_2828280_1580640# gnd! 63.9fF
C1399 diff_2803120_1629480# gnd! 64.8fF
C1400 diff_2777960_1556960# gnd! 81.8fF
C1401 diff_2752800_1629480# gnd! 81.7fF
C1402 diff_2727640_1580640# gnd! 63.9fF
C1403 diff_2702480_1629480# gnd! 64.8fF
C1404 diff_2677320_1556960# gnd! 81.8fF
C1405 diff_2652160_1629480# gnd! 81.7fF
C1406 diff_2627000_1580640# gnd! 63.9fF
C1407 diff_2601840_1629480# gnd! 64.8fF
C1408 diff_2576680_1556960# gnd! 81.8fF
C1409 diff_2551520_1629480# gnd! 81.7fF
C1410 diff_2526360_1580640# gnd! 63.9fF
C1411 diff_2501200_1629480# gnd! 64.8fF
C1412 diff_2476040_1556960# gnd! 81.8fF
C1413 diff_2450880_1629480# gnd! 81.7fF
C1414 diff_2425720_1580640# gnd! 63.9fF
C1415 diff_2400560_1629480# gnd! 64.8fF
C1416 diff_2375400_1556960# gnd! 81.8fF
C1417 diff_2350240_1629480# gnd! 81.7fF
C1418 diff_2325080_1580640# gnd! 63.9fF
C1419 diff_2299920_1629480# gnd! 64.8fF
C1420 diff_2274760_1556960# gnd! 81.8fF
C1421 diff_2249600_1629480# gnd! 81.7fF
C1422 diff_2224440_1580640# gnd! 63.9fF
C1423 diff_2199280_1629480# gnd! 64.8fF
C1424 diff_2174120_1556960# gnd! 81.8fF
C1425 diff_2148960_1629480# gnd! 81.7fF
C1426 diff_2123800_1580640# gnd! 63.9fF
C1427 diff_2098640_1629480# gnd! 64.8fF
C1428 diff_2073480_1556960# gnd! 81.8fF
C1429 diff_2048320_1629480# gnd! 81.7fF
C1430 diff_2023160_1580640# gnd! 63.9fF
C1431 diff_1998000_1629480# gnd! 64.8fF
C1432 diff_1972840_1556960# gnd! 81.8fF
C1433 diff_1947680_1629480# gnd! 81.7fF
C1434 diff_1922520_1580640# gnd! 63.9fF
C1435 diff_1897360_1629480# gnd! 64.8fF
C1436 diff_1872200_1556960# gnd! 81.8fF
C1437 diff_1847040_1629480# gnd! 81.7fF
C1438 diff_1821880_1580640# gnd! 63.9fF
C1439 diff_1796720_1629480# gnd! 64.8fF
C1440 diff_1771560_1556960# gnd! 81.8fF
C1441 diff_1746400_1629480# gnd! 81.7fF
C1442 diff_1721240_1580640# gnd! 63.9fF
C1443 diff_1696080_1629480# gnd! 64.8fF
C1444 diff_1670920_1556960# gnd! 81.8fF
C1445 diff_1645760_1629480# gnd! 81.7fF
C1446 diff_1620600_1580640# gnd! 63.9fF
C1447 diff_1595440_1629480# gnd! 64.8fF
C1448 diff_1570280_1556960# gnd! 81.8fF
C1449 diff_1545120_1629480# gnd! 81.7fF
C1450 diff_1519960_1580640# gnd! 63.9fF
C1451 diff_1494800_1629480# gnd! 64.8fF
C1452 diff_1469640_1556960# gnd! 81.8fF
C1453 diff_1444480_1629480# gnd! 81.7fF
C1454 diff_1419320_1580640# gnd! 63.9fF
C1455 diff_1394160_1629480# gnd! 64.8fF
C1456 diff_1369000_1556960# gnd! 81.8fF
C1457 diff_1343840_1629480# gnd! 81.7fF
C1458 diff_1318680_1580640# gnd! 62.3fF
C1459 diff_1293520_1630960# gnd! 63.5fF
C1460 diff_1263920_1558440# gnd! 85.3fF
C1461 diff_985680_1574720# gnd! 454.3fF
C1462 diff_627520_1602840# gnd! 304.5fF
C1463 diff_797720_1443000# gnd! 478.6fF
C1464 diff_794760_1574720# gnd! 452.9fF
C1465 diff_438080_1602840# gnd! 305.5fF
C1466 diff_606800_1443000# gnd! 462.9fF
C1467 diff_602360_1574720# gnd! 442.7fF
C1468 diff_414400_1443000# gnd! 465.0fF
C1469 diff_411440_1576200# gnd! 450.9fF
C1470 diff_346320_1623560# gnd! 206.4fF
C1471 diff_1243200_1628000# gnd! 75.3fF
C1472 diff_1238760_1660560# gnd! 926.2fF
C1473 diff_2828280_1667960# gnd! 38.4fF
C1474 diff_2803120_1667960# gnd! 38.4fF
C1475 diff_2777960_1667960# gnd! 38.4fF
C1476 diff_2752800_1667960# gnd! 38.4fF
C1477 diff_2727640_1667960# gnd! 38.4fF
C1478 diff_2702480_1667960# gnd! 38.4fF
C1479 diff_2677320_1667960# gnd! 38.4fF
C1480 diff_2652160_1667960# gnd! 38.4fF
C1481 diff_2627000_1667960# gnd! 38.4fF
C1482 diff_2601840_1667960# gnd! 38.4fF
C1483 diff_2576680_1667960# gnd! 38.4fF
C1484 diff_2551520_1667960# gnd! 38.4fF
C1485 diff_2526360_1667960# gnd! 38.4fF
C1486 diff_2501200_1667960# gnd! 38.4fF
C1487 diff_2476040_1667960# gnd! 38.4fF
C1488 diff_2450880_1667960# gnd! 38.4fF
C1489 diff_2425720_1667960# gnd! 38.4fF
C1490 diff_2400560_1667960# gnd! 38.4fF
C1491 diff_2375400_1667960# gnd! 38.4fF
C1492 diff_2350240_1667960# gnd! 38.4fF
C1493 diff_2325080_1667960# gnd! 38.4fF
C1494 diff_2299920_1667960# gnd! 38.4fF
C1495 diff_2274760_1667960# gnd! 38.4fF
C1496 diff_2249600_1667960# gnd! 38.4fF
C1497 diff_2224440_1667960# gnd! 38.4fF
C1498 diff_2199280_1667960# gnd! 38.4fF
C1499 diff_2174120_1667960# gnd! 38.4fF
C1500 diff_2148960_1667960# gnd! 38.4fF
C1501 diff_2123800_1667960# gnd! 38.4fF
C1502 diff_2098640_1667960# gnd! 38.4fF
C1503 diff_2073480_1667960# gnd! 38.4fF
C1504 diff_2048320_1667960# gnd! 38.4fF
C1505 diff_2023160_1667960# gnd! 38.4fF
C1506 diff_1998000_1667960# gnd! 38.4fF
C1507 diff_1972840_1667960# gnd! 38.4fF
C1508 diff_1947680_1667960# gnd! 38.4fF
C1509 diff_1922520_1667960# gnd! 38.4fF
C1510 diff_1897360_1667960# gnd! 38.4fF
C1511 diff_1872200_1667960# gnd! 38.4fF
C1512 diff_1847040_1667960# gnd! 38.4fF
C1513 diff_1821880_1667960# gnd! 38.4fF
C1514 diff_1796720_1667960# gnd! 38.4fF
C1515 diff_1771560_1667960# gnd! 38.4fF
C1516 diff_1746400_1667960# gnd! 38.4fF
C1517 diff_1721240_1667960# gnd! 38.4fF
C1518 diff_1696080_1667960# gnd! 38.4fF
C1519 diff_1670920_1667960# gnd! 38.4fF
C1520 diff_1645760_1667960# gnd! 38.4fF
C1521 diff_1620600_1667960# gnd! 38.4fF
C1522 diff_1595440_1667960# gnd! 38.4fF
C1523 diff_1570280_1667960# gnd! 38.4fF
C1524 diff_1545120_1667960# gnd! 38.4fF
C1525 diff_1519960_1667960# gnd! 38.4fF
C1526 diff_1494800_1667960# gnd! 38.4fF
C1527 diff_1469640_1667960# gnd! 38.4fF
C1528 diff_1444480_1667960# gnd! 38.4fF
C1529 diff_1419320_1667960# gnd! 38.4fF
C1530 diff_1394160_1667960# gnd! 38.4fF
C1531 diff_1369000_1667960# gnd! 38.4fF
C1532 diff_1343840_1667960# gnd! 38.4fF
C1533 diff_1318680_1667960# gnd! 38.4fF
C1534 diff_1293520_1667960# gnd! 38.4fF
C1535 diff_1268360_1667960# gnd! 38.4fF
C1536 diff_985680_1660560# gnd! 20.4fF
C1537 diff_794760_1660560# gnd! 20.4fF
C1538 diff_602360_1660560# gnd! 20.4fF
C1539 diff_411440_1660560# gnd! 20.4fF
C1540 diff_190920_1013800# gnd! 927.2fF
C1541 diff_1243200_1667960# gnd! 38.4fF
C1542 diff_1238760_1688680# gnd! 973.7fF
C1543 diff_2828280_1696080# gnd! 36.1fF
C1544 diff_2803120_1696080# gnd! 36.1fF
C1545 diff_2777960_1696080# gnd! 36.1fF
C1546 diff_2752800_1696080# gnd! 36.1fF
C1547 diff_2727640_1696080# gnd! 36.1fF
C1548 diff_2702480_1696080# gnd! 36.1fF
C1549 diff_2677320_1696080# gnd! 36.1fF
C1550 diff_2652160_1696080# gnd! 36.1fF
C1551 diff_2627000_1696080# gnd! 36.1fF
C1552 diff_2601840_1696080# gnd! 36.1fF
C1553 diff_2576680_1696080# gnd! 36.1fF
C1554 diff_2551520_1696080# gnd! 36.1fF
C1555 diff_2526360_1696080# gnd! 36.1fF
C1556 diff_2501200_1696080# gnd! 36.1fF
C1557 diff_2476040_1696080# gnd! 36.1fF
C1558 diff_2450880_1696080# gnd! 36.1fF
C1559 diff_2425720_1696080# gnd! 36.1fF
C1560 diff_2400560_1696080# gnd! 36.1fF
C1561 diff_2375400_1696080# gnd! 36.1fF
C1562 diff_2350240_1696080# gnd! 36.1fF
C1563 diff_2325080_1696080# gnd! 36.1fF
C1564 diff_2299920_1696080# gnd! 36.1fF
C1565 diff_2274760_1696080# gnd! 36.1fF
C1566 diff_2249600_1696080# gnd! 36.1fF
C1567 diff_2224440_1696080# gnd! 36.1fF
C1568 diff_2199280_1696080# gnd! 36.1fF
C1569 diff_2174120_1696080# gnd! 36.1fF
C1570 diff_2148960_1696080# gnd! 36.1fF
C1571 diff_2123800_1696080# gnd! 36.1fF
C1572 diff_2098640_1696080# gnd! 36.1fF
C1573 diff_2073480_1696080# gnd! 36.1fF
C1574 diff_2048320_1696080# gnd! 36.1fF
C1575 diff_2023160_1696080# gnd! 36.1fF
C1576 diff_1998000_1696080# gnd! 36.1fF
C1577 diff_1972840_1696080# gnd! 36.1fF
C1578 diff_1947680_1696080# gnd! 36.1fF
C1579 diff_1922520_1696080# gnd! 36.1fF
C1580 diff_1897360_1696080# gnd! 36.1fF
C1581 diff_1872200_1696080# gnd! 36.1fF
C1582 diff_1847040_1696080# gnd! 36.1fF
C1583 diff_1821880_1696080# gnd! 36.1fF
C1584 diff_1796720_1696080# gnd! 36.1fF
C1585 diff_1771560_1696080# gnd! 36.1fF
C1586 diff_1746400_1696080# gnd! 36.1fF
C1587 diff_1721240_1696080# gnd! 36.1fF
C1588 diff_1696080_1696080# gnd! 36.1fF
C1589 diff_1670920_1696080# gnd! 36.1fF
C1590 diff_1645760_1696080# gnd! 36.1fF
C1591 diff_1620600_1696080# gnd! 36.1fF
C1592 diff_1595440_1696080# gnd! 36.1fF
C1593 diff_1570280_1696080# gnd! 36.1fF
C1594 diff_1545120_1696080# gnd! 36.1fF
C1595 diff_1519960_1696080# gnd! 36.1fF
C1596 diff_1494800_1696080# gnd! 36.1fF
C1597 diff_1469640_1696080# gnd! 36.1fF
C1598 diff_1444480_1696080# gnd! 36.1fF
C1599 diff_1419320_1696080# gnd! 36.1fF
C1600 diff_1394160_1696080# gnd! 36.1fF
C1601 diff_1369000_1696080# gnd! 36.1fF
C1602 diff_1343840_1696080# gnd! 36.1fF
C1603 diff_1318680_1696080# gnd! 36.1fF
C1604 diff_1293520_1696080# gnd! 36.1fF
C1605 diff_1268360_1696080# gnd! 36.1fF
C1606 diff_1243200_1696080# gnd! 36.1fF
C1607 diff_1238760_1715320# gnd! 981.4fF
C1608 diff_2920040_1736040# gnd! 740.2fF
C1609 diff_2828280_1722720# gnd! 38.4fF
C1610 diff_2803120_1722720# gnd! 38.4fF
C1611 diff_2777960_1722720# gnd! 38.4fF
C1612 diff_2752800_1722720# gnd! 38.4fF
C1613 diff_2727640_1722720# gnd! 38.4fF
C1614 diff_2702480_1722720# gnd! 38.4fF
C1615 diff_2677320_1722720# gnd! 38.4fF
C1616 diff_2652160_1722720# gnd! 38.4fF
C1617 diff_2627000_1722720# gnd! 38.4fF
C1618 diff_2601840_1722720# gnd! 38.4fF
C1619 diff_2576680_1722720# gnd! 38.4fF
C1620 diff_2551520_1722720# gnd! 38.4fF
C1621 diff_2526360_1722720# gnd! 38.4fF
C1622 diff_2501200_1722720# gnd! 38.4fF
C1623 diff_2476040_1722720# gnd! 38.4fF
C1624 diff_2450880_1722720# gnd! 38.4fF
C1625 diff_2425720_1722720# gnd! 38.4fF
C1626 diff_2400560_1722720# gnd! 38.4fF
C1627 diff_2375400_1722720# gnd! 38.4fF
C1628 diff_2350240_1722720# gnd! 38.4fF
C1629 diff_2325080_1722720# gnd! 38.4fF
C1630 diff_2299920_1722720# gnd! 38.4fF
C1631 diff_2274760_1722720# gnd! 38.4fF
C1632 diff_2249600_1722720# gnd! 38.4fF
C1633 diff_2224440_1722720# gnd! 38.4fF
C1634 diff_2199280_1722720# gnd! 38.4fF
C1635 diff_2174120_1722720# gnd! 38.4fF
C1636 diff_2148960_1722720# gnd! 38.4fF
C1637 diff_2123800_1722720# gnd! 38.4fF
C1638 diff_2098640_1722720# gnd! 38.4fF
C1639 diff_2073480_1722720# gnd! 38.4fF
C1640 diff_2048320_1722720# gnd! 38.4fF
C1641 diff_2023160_1722720# gnd! 38.4fF
C1642 diff_1998000_1722720# gnd! 38.4fF
C1643 diff_1972840_1722720# gnd! 38.4fF
C1644 diff_1947680_1722720# gnd! 38.4fF
C1645 diff_1922520_1722720# gnd! 38.4fF
C1646 diff_1897360_1722720# gnd! 38.4fF
C1647 diff_1872200_1722720# gnd! 38.4fF
C1648 diff_1847040_1722720# gnd! 38.4fF
C1649 diff_1821880_1722720# gnd! 38.4fF
C1650 diff_1796720_1722720# gnd! 38.4fF
C1651 diff_1771560_1722720# gnd! 38.4fF
C1652 diff_1746400_1722720# gnd! 38.4fF
C1653 diff_1721240_1722720# gnd! 38.4fF
C1654 diff_1696080_1722720# gnd! 38.4fF
C1655 diff_1670920_1722720# gnd! 38.4fF
C1656 diff_1645760_1722720# gnd! 38.4fF
C1657 diff_1620600_1722720# gnd! 38.4fF
C1658 diff_1595440_1722720# gnd! 38.4fF
C1659 diff_1570280_1722720# gnd! 38.4fF
C1660 diff_1545120_1722720# gnd! 38.4fF
C1661 diff_1519960_1722720# gnd! 38.4fF
C1662 diff_1494800_1722720# gnd! 38.4fF
C1663 diff_1469640_1722720# gnd! 38.4fF
C1664 diff_1444480_1722720# gnd! 38.4fF
C1665 diff_1419320_1722720# gnd! 38.4fF
C1666 diff_1394160_1722720# gnd! 38.4fF
C1667 diff_1369000_1722720# gnd! 38.4fF
C1668 diff_1343840_1722720# gnd! 38.4fF
C1669 diff_1318680_1722720# gnd! 38.4fF
C1670 diff_1293520_1722720# gnd! 38.4fF
C1671 diff_1268360_1722720# gnd! 38.4fF
C1672 diff_1243200_1722720# gnd! 38.4fF
C1673 diff_1238760_1743440# gnd! 920.4fF
C1674 diff_2828280_1750840# gnd! 36.1fF
C1675 diff_2803120_1750840# gnd! 36.1fF
C1676 diff_2777960_1750840# gnd! 36.1fF
C1677 diff_2752800_1750840# gnd! 36.1fF
C1678 diff_2727640_1750840# gnd! 36.1fF
C1679 diff_2702480_1750840# gnd! 36.1fF
C1680 diff_2677320_1750840# gnd! 36.1fF
C1681 diff_2652160_1750840# gnd! 36.1fF
C1682 diff_2627000_1750840# gnd! 36.1fF
C1683 diff_2601840_1750840# gnd! 36.1fF
C1684 diff_2576680_1750840# gnd! 36.1fF
C1685 diff_2551520_1750840# gnd! 36.1fF
C1686 diff_2526360_1750840# gnd! 36.1fF
C1687 diff_2501200_1750840# gnd! 36.1fF
C1688 diff_2476040_1750840# gnd! 36.1fF
C1689 diff_2450880_1750840# gnd! 36.1fF
C1690 diff_2425720_1750840# gnd! 36.1fF
C1691 diff_2400560_1750840# gnd! 36.1fF
C1692 diff_2375400_1750840# gnd! 36.1fF
C1693 diff_2350240_1750840# gnd! 36.1fF
C1694 diff_2325080_1750840# gnd! 36.1fF
C1695 diff_2299920_1750840# gnd! 36.1fF
C1696 diff_2274760_1750840# gnd! 36.1fF
C1697 diff_2249600_1750840# gnd! 36.1fF
C1698 diff_2224440_1750840# gnd! 36.1fF
C1699 diff_2199280_1750840# gnd! 36.1fF
C1700 diff_2174120_1750840# gnd! 36.1fF
C1701 diff_2148960_1750840# gnd! 36.1fF
C1702 diff_2123800_1750840# gnd! 36.1fF
C1703 diff_2098640_1750840# gnd! 36.1fF
C1704 diff_2073480_1750840# gnd! 36.1fF
C1705 diff_2048320_1750840# gnd! 36.1fF
C1706 diff_2023160_1750840# gnd! 36.1fF
C1707 diff_1998000_1750840# gnd! 36.1fF
C1708 diff_1972840_1750840# gnd! 36.1fF
C1709 diff_1947680_1750840# gnd! 36.1fF
C1710 diff_1922520_1750840# gnd! 36.1fF
C1711 diff_1897360_1750840# gnd! 36.1fF
C1712 diff_1872200_1750840# gnd! 36.1fF
C1713 diff_1847040_1750840# gnd! 36.1fF
C1714 diff_1821880_1750840# gnd! 36.1fF
C1715 diff_1796720_1750840# gnd! 36.1fF
C1716 diff_1771560_1750840# gnd! 36.1fF
C1717 diff_1746400_1750840# gnd! 36.1fF
C1718 diff_1721240_1750840# gnd! 36.1fF
C1719 diff_1696080_1750840# gnd! 36.1fF
C1720 diff_1670920_1750840# gnd! 36.1fF
C1721 diff_1645760_1750840# gnd! 36.1fF
C1722 diff_1620600_1750840# gnd! 36.1fF
C1723 diff_1595440_1750840# gnd! 36.1fF
C1724 diff_1570280_1750840# gnd! 36.1fF
C1725 diff_1545120_1750840# gnd! 36.1fF
C1726 diff_1519960_1750840# gnd! 36.1fF
C1727 diff_1494800_1750840# gnd! 36.1fF
C1728 diff_1469640_1750840# gnd! 36.1fF
C1729 diff_1444480_1750840# gnd! 36.1fF
C1730 diff_1419320_1750840# gnd! 36.1fF
C1731 diff_1394160_1750840# gnd! 36.1fF
C1732 diff_1369000_1750840# gnd! 36.1fF
C1733 diff_1343840_1750840# gnd! 36.1fF
C1734 diff_1318680_1750840# gnd! 36.1fF
C1735 diff_1293520_1750840# gnd! 36.1fF
C1736 diff_1268360_1750840# gnd! 36.1fF
C1737 diff_1243200_1750840# gnd! 36.1fF
C1738 diff_1238760_1770080# gnd! 927.2fF
C1739 diff_2828280_1777480# gnd! 38.4fF
C1740 diff_2803120_1777480# gnd! 38.4fF
C1741 diff_2777960_1777480# gnd! 38.4fF
C1742 diff_2752800_1777480# gnd! 38.4fF
C1743 diff_2727640_1777480# gnd! 38.4fF
C1744 diff_2702480_1777480# gnd! 38.4fF
C1745 diff_2677320_1777480# gnd! 38.4fF
C1746 diff_2652160_1777480# gnd! 38.4fF
C1747 diff_2627000_1777480# gnd! 38.4fF
C1748 diff_2601840_1777480# gnd! 38.4fF
C1749 diff_2576680_1777480# gnd! 38.4fF
C1750 diff_2551520_1777480# gnd! 38.4fF
C1751 diff_2526360_1777480# gnd! 38.4fF
C1752 diff_2501200_1777480# gnd! 38.4fF
C1753 diff_2476040_1777480# gnd! 38.4fF
C1754 diff_2450880_1777480# gnd! 38.4fF
C1755 diff_2425720_1777480# gnd! 38.4fF
C1756 diff_2400560_1777480# gnd! 38.4fF
C1757 diff_2375400_1777480# gnd! 38.4fF
C1758 diff_2350240_1777480# gnd! 38.4fF
C1759 diff_2325080_1777480# gnd! 38.4fF
C1760 diff_2299920_1777480# gnd! 38.4fF
C1761 diff_2274760_1777480# gnd! 38.4fF
C1762 diff_2249600_1777480# gnd! 38.4fF
C1763 diff_2224440_1777480# gnd! 38.4fF
C1764 diff_2199280_1777480# gnd! 38.4fF
C1765 diff_2174120_1777480# gnd! 38.4fF
C1766 diff_2148960_1777480# gnd! 38.4fF
C1767 diff_2123800_1777480# gnd! 38.4fF
C1768 diff_2098640_1777480# gnd! 38.4fF
C1769 diff_2073480_1777480# gnd! 38.4fF
C1770 diff_2048320_1777480# gnd! 38.4fF
C1771 diff_2023160_1777480# gnd! 38.4fF
C1772 diff_1998000_1777480# gnd! 38.4fF
C1773 diff_1972840_1777480# gnd! 38.4fF
C1774 diff_1947680_1777480# gnd! 38.4fF
C1775 diff_1922520_1777480# gnd! 38.4fF
C1776 diff_1897360_1777480# gnd! 38.4fF
C1777 diff_1872200_1777480# gnd! 38.4fF
C1778 diff_1847040_1777480# gnd! 38.4fF
C1779 diff_1821880_1777480# gnd! 38.4fF
C1780 diff_1796720_1777480# gnd! 38.4fF
C1781 diff_1771560_1777480# gnd! 38.4fF
C1782 diff_1746400_1777480# gnd! 38.4fF
C1783 diff_1721240_1777480# gnd! 38.4fF
C1784 diff_1696080_1777480# gnd! 38.4fF
C1785 diff_1670920_1777480# gnd! 38.4fF
C1786 diff_1645760_1777480# gnd! 38.4fF
C1787 diff_1620600_1777480# gnd! 38.4fF
C1788 diff_1595440_1777480# gnd! 38.4fF
C1789 diff_1570280_1777480# gnd! 38.4fF
C1790 diff_1545120_1777480# gnd! 38.4fF
C1791 diff_1519960_1777480# gnd! 38.4fF
C1792 diff_1494800_1777480# gnd! 38.4fF
C1793 diff_1469640_1777480# gnd! 38.4fF
C1794 diff_1444480_1777480# gnd! 38.4fF
C1795 diff_1419320_1777480# gnd! 38.4fF
C1796 diff_1394160_1777480# gnd! 38.4fF
C1797 diff_1369000_1777480# gnd! 38.4fF
C1798 diff_1343840_1777480# gnd! 38.4fF
C1799 diff_1318680_1777480# gnd! 38.4fF
C1800 diff_1293520_1777480# gnd! 38.4fF
C1801 diff_1268360_1777480# gnd! 38.4fF
C1802 diff_1243200_1777480# gnd! 38.4fF
C1803 diff_1238760_1798200# gnd! 975.6fF
C1804 diff_2828280_1805600# gnd! 36.1fF
C1805 diff_2803120_1805600# gnd! 36.1fF
C1806 diff_2777960_1805600# gnd! 36.1fF
C1807 diff_2752800_1805600# gnd! 36.1fF
C1808 diff_2727640_1805600# gnd! 36.1fF
C1809 diff_2702480_1805600# gnd! 36.1fF
C1810 diff_2677320_1805600# gnd! 36.1fF
C1811 diff_2652160_1805600# gnd! 36.1fF
C1812 diff_2627000_1805600# gnd! 36.1fF
C1813 diff_2601840_1805600# gnd! 36.1fF
C1814 diff_2576680_1805600# gnd! 36.1fF
C1815 diff_2551520_1805600# gnd! 36.1fF
C1816 diff_2526360_1805600# gnd! 36.1fF
C1817 diff_2501200_1805600# gnd! 36.1fF
C1818 diff_2476040_1805600# gnd! 36.1fF
C1819 diff_2450880_1805600# gnd! 36.1fF
C1820 diff_2425720_1805600# gnd! 36.1fF
C1821 diff_2400560_1805600# gnd! 36.1fF
C1822 diff_2375400_1805600# gnd! 36.1fF
C1823 diff_2350240_1805600# gnd! 36.1fF
C1824 diff_2325080_1805600# gnd! 36.1fF
C1825 diff_2299920_1805600# gnd! 36.1fF
C1826 diff_2274760_1805600# gnd! 36.1fF
C1827 diff_2249600_1805600# gnd! 36.1fF
C1828 diff_2224440_1805600# gnd! 36.1fF
C1829 diff_2199280_1805600# gnd! 36.1fF
C1830 diff_2174120_1805600# gnd! 36.1fF
C1831 diff_2148960_1805600# gnd! 36.1fF
C1832 diff_2123800_1805600# gnd! 36.1fF
C1833 diff_2098640_1805600# gnd! 36.1fF
C1834 diff_2073480_1805600# gnd! 36.1fF
C1835 diff_2048320_1805600# gnd! 36.1fF
C1836 diff_2023160_1805600# gnd! 36.1fF
C1837 diff_1998000_1805600# gnd! 36.1fF
C1838 diff_1972840_1805600# gnd! 36.1fF
C1839 diff_1947680_1805600# gnd! 36.1fF
C1840 diff_1922520_1805600# gnd! 36.1fF
C1841 diff_1897360_1805600# gnd! 36.1fF
C1842 diff_1872200_1805600# gnd! 36.1fF
C1843 diff_1847040_1805600# gnd! 36.1fF
C1844 diff_1821880_1805600# gnd! 36.1fF
C1845 diff_1796720_1805600# gnd! 36.1fF
C1846 diff_1771560_1805600# gnd! 36.1fF
C1847 diff_1746400_1805600# gnd! 36.1fF
C1848 diff_1721240_1805600# gnd! 36.1fF
C1849 diff_1696080_1805600# gnd! 36.1fF
C1850 diff_1670920_1805600# gnd! 36.1fF
C1851 diff_1645760_1805600# gnd! 36.1fF
C1852 diff_1620600_1805600# gnd! 36.1fF
C1853 diff_1595440_1805600# gnd! 36.1fF
C1854 diff_1570280_1805600# gnd! 36.1fF
C1855 diff_1545120_1805600# gnd! 36.1fF
C1856 diff_1519960_1805600# gnd! 36.1fF
C1857 diff_1494800_1805600# gnd! 36.1fF
C1858 diff_1469640_1805600# gnd! 36.1fF
C1859 diff_1444480_1805600# gnd! 36.1fF
C1860 diff_1419320_1805600# gnd! 36.1fF
C1861 diff_1394160_1805600# gnd! 36.1fF
C1862 diff_1369000_1805600# gnd! 36.1fF
C1863 diff_1343840_1805600# gnd! 36.1fF
C1864 diff_1318680_1805600# gnd! 36.1fF
C1865 diff_1293520_1805600# gnd! 36.1fF
C1866 diff_1268360_1805600# gnd! 36.1fF
C1867 diff_1243200_1805600# gnd! 36.1fF
C1868 diff_1238760_1824840# gnd! 982.6fF
C1869 diff_3023640_1207680# gnd! 941.1fF
C1870 diff_3045840_1124800# gnd! 748.1fF
C1871 diff_3196800_1889960# gnd! 118.3fF
C1872 diff_3469120_1237280# gnd! 870.5fF
C1873 diff_3412880_1952120# gnd! 80.9fF
C1874 diff_3343320_1672400# gnd! 804.1fF
C1875 diff_3488360_1570280# gnd! 464.5fF
C1876 diff_3488360_1339400# gnd! 862.6fF
C1877 diff_3307800_2085320# gnd! 80.1fF
C1878 diff_3267840_1873680# gnd! 572.8fF
C1879 diff_3383280_2100120# gnd! 81.4fF
C1880 diff_3285600_1753800# gnd! 367.3fF
C1881 diff_3383280_2114920# gnd! 72.0fF
C1882 diff_2920040_1842600# gnd! 784.4fF
C1883 diff_2828280_1832240# gnd! 38.4fF
C1884 diff_2803120_1832240# gnd! 38.4fF
C1885 diff_2777960_1832240# gnd! 38.4fF
C1886 diff_2752800_1832240# gnd! 38.4fF
C1887 diff_2727640_1832240# gnd! 38.4fF
C1888 diff_2702480_1832240# gnd! 38.4fF
C1889 diff_2677320_1832240# gnd! 38.4fF
C1890 diff_2652160_1832240# gnd! 38.4fF
C1891 diff_2627000_1832240# gnd! 38.4fF
C1892 diff_2601840_1832240# gnd! 38.4fF
C1893 diff_2576680_1832240# gnd! 38.4fF
C1894 diff_2551520_1832240# gnd! 38.4fF
C1895 diff_2526360_1832240# gnd! 38.4fF
C1896 diff_2501200_1832240# gnd! 38.4fF
C1897 diff_2476040_1832240# gnd! 38.4fF
C1898 diff_2450880_1832240# gnd! 38.4fF
C1899 diff_2425720_1832240# gnd! 38.4fF
C1900 diff_2400560_1832240# gnd! 38.4fF
C1901 diff_2375400_1832240# gnd! 38.4fF
C1902 diff_2350240_1832240# gnd! 38.4fF
C1903 diff_2325080_1832240# gnd! 38.4fF
C1904 diff_2299920_1832240# gnd! 38.4fF
C1905 diff_2274760_1832240# gnd! 38.4fF
C1906 diff_2249600_1832240# gnd! 38.4fF
C1907 diff_2224440_1832240# gnd! 38.4fF
C1908 diff_2199280_1832240# gnd! 38.4fF
C1909 diff_2174120_1832240# gnd! 38.4fF
C1910 diff_2148960_1832240# gnd! 38.4fF
C1911 diff_2123800_1832240# gnd! 38.4fF
C1912 diff_2098640_1832240# gnd! 38.4fF
C1913 diff_2073480_1832240# gnd! 38.4fF
C1914 diff_2048320_1832240# gnd! 38.4fF
C1915 diff_2023160_1832240# gnd! 38.4fF
C1916 diff_1998000_1832240# gnd! 38.4fF
C1917 diff_1972840_1832240# gnd! 38.4fF
C1918 diff_1947680_1832240# gnd! 38.4fF
C1919 diff_1922520_1832240# gnd! 38.4fF
C1920 diff_1897360_1832240# gnd! 38.4fF
C1921 diff_1872200_1832240# gnd! 38.4fF
C1922 diff_1847040_1832240# gnd! 38.4fF
C1923 diff_1821880_1832240# gnd! 38.4fF
C1924 diff_1796720_1832240# gnd! 38.4fF
C1925 diff_1771560_1832240# gnd! 38.4fF
C1926 diff_1746400_1832240# gnd! 38.4fF
C1927 diff_1721240_1832240# gnd! 38.4fF
C1928 diff_1696080_1832240# gnd! 38.4fF
C1929 diff_1670920_1832240# gnd! 38.4fF
C1930 diff_1645760_1832240# gnd! 38.4fF
C1931 diff_1620600_1832240# gnd! 38.4fF
C1932 diff_1595440_1832240# gnd! 38.4fF
C1933 diff_1570280_1832240# gnd! 38.4fF
C1934 diff_1545120_1832240# gnd! 38.4fF
C1935 diff_1519960_1832240# gnd! 38.4fF
C1936 diff_1494800_1832240# gnd! 38.4fF
C1937 diff_1469640_1832240# gnd! 38.4fF
C1938 diff_1444480_1832240# gnd! 38.4fF
C1939 diff_1419320_1832240# gnd! 38.4fF
C1940 diff_1394160_1832240# gnd! 38.4fF
C1941 diff_1369000_1832240# gnd! 38.4fF
C1942 diff_1343840_1832240# gnd! 38.4fF
C1943 diff_1318680_1832240# gnd! 38.4fF
C1944 diff_1293520_1832240# gnd! 38.4fF
C1945 diff_1268360_1832240# gnd! 38.4fF
C1946 diff_1077440_1786360# gnd! 227.2fF
C1947 diff_1243200_1832240# gnd! 38.4fF
C1948 diff_886520_1786360# gnd! 464.3fF
C1949 diff_1238760_1852960# gnd! 916.2fF
C1950 diff_2828280_1860360# gnd! 36.1fF
C1951 diff_2803120_1860360# gnd! 36.1fF
C1952 diff_2777960_1860360# gnd! 36.1fF
C1953 diff_2752800_1860360# gnd! 36.1fF
C1954 diff_2727640_1860360# gnd! 36.1fF
C1955 diff_2702480_1860360# gnd! 36.1fF
C1956 diff_2677320_1860360# gnd! 36.1fF
C1957 diff_2652160_1860360# gnd! 36.1fF
C1958 diff_2627000_1860360# gnd! 36.1fF
C1959 diff_2601840_1860360# gnd! 36.1fF
C1960 diff_2576680_1860360# gnd! 36.1fF
C1961 diff_2551520_1860360# gnd! 36.1fF
C1962 diff_2526360_1860360# gnd! 36.1fF
C1963 diff_2501200_1860360# gnd! 36.1fF
C1964 diff_2476040_1860360# gnd! 36.1fF
C1965 diff_2450880_1860360# gnd! 36.1fF
C1966 diff_2425720_1860360# gnd! 36.1fF
C1967 diff_2400560_1860360# gnd! 36.1fF
C1968 diff_2375400_1860360# gnd! 36.1fF
C1969 diff_2350240_1860360# gnd! 36.1fF
C1970 diff_2325080_1860360# gnd! 36.1fF
C1971 diff_2299920_1860360# gnd! 36.1fF
C1972 diff_2274760_1860360# gnd! 36.1fF
C1973 diff_2249600_1860360# gnd! 36.1fF
C1974 diff_2224440_1860360# gnd! 36.1fF
C1975 diff_2199280_1860360# gnd! 36.1fF
C1976 diff_2174120_1860360# gnd! 36.1fF
C1977 diff_2148960_1860360# gnd! 36.1fF
C1978 diff_2123800_1860360# gnd! 36.1fF
C1979 diff_2098640_1860360# gnd! 36.1fF
C1980 diff_2073480_1860360# gnd! 36.1fF
C1981 diff_2048320_1860360# gnd! 36.1fF
C1982 diff_2023160_1860360# gnd! 36.1fF
C1983 diff_1998000_1860360# gnd! 36.1fF
C1984 diff_1972840_1860360# gnd! 36.1fF
C1985 diff_1947680_1860360# gnd! 36.1fF
C1986 diff_1922520_1860360# gnd! 36.1fF
C1987 diff_1897360_1860360# gnd! 36.1fF
C1988 diff_1872200_1860360# gnd! 36.1fF
C1989 diff_1847040_1860360# gnd! 36.1fF
C1990 diff_1821880_1860360# gnd! 36.1fF
C1991 diff_1796720_1860360# gnd! 36.1fF
C1992 diff_1771560_1860360# gnd! 36.1fF
C1993 diff_1746400_1860360# gnd! 36.1fF
C1994 diff_1721240_1860360# gnd! 36.1fF
C1995 diff_1696080_1860360# gnd! 36.1fF
C1996 diff_1670920_1860360# gnd! 36.1fF
C1997 diff_1645760_1860360# gnd! 36.1fF
C1998 diff_1620600_1860360# gnd! 36.1fF
C1999 diff_1595440_1860360# gnd! 36.1fF
C2000 diff_1570280_1860360# gnd! 36.1fF
C2001 diff_1545120_1860360# gnd! 36.1fF
C2002 diff_1519960_1860360# gnd! 36.1fF
C2003 diff_1494800_1860360# gnd! 36.1fF
C2004 diff_1469640_1860360# gnd! 36.1fF
C2005 diff_1444480_1860360# gnd! 36.1fF
C2006 diff_1419320_1860360# gnd! 36.1fF
C2007 diff_1394160_1860360# gnd! 36.1fF
C2008 diff_1369000_1860360# gnd! 36.1fF
C2009 diff_1343840_1860360# gnd! 36.1fF
C2010 diff_1318680_1860360# gnd! 36.1fF
C2011 diff_1293520_1860360# gnd! 36.1fF
C2012 diff_1268360_1860360# gnd! 36.1fF
C2013 diff_1243200_1860360# gnd! 36.1fF
C2014 diff_1238760_1879600# gnd! 927.6fF
C2015 diff_2828280_1887000# gnd! 38.4fF
C2016 diff_2803120_1887000# gnd! 38.4fF
C2017 diff_2777960_1887000# gnd! 38.4fF
C2018 diff_2752800_1887000# gnd! 38.4fF
C2019 diff_2727640_1887000# gnd! 38.4fF
C2020 diff_2702480_1887000# gnd! 38.4fF
C2021 diff_2677320_1887000# gnd! 38.4fF
C2022 diff_2652160_1887000# gnd! 38.4fF
C2023 diff_2627000_1887000# gnd! 38.4fF
C2024 diff_2601840_1887000# gnd! 38.4fF
C2025 diff_2576680_1887000# gnd! 38.4fF
C2026 diff_2551520_1887000# gnd! 38.4fF
C2027 diff_2526360_1887000# gnd! 38.4fF
C2028 diff_2501200_1887000# gnd! 38.4fF
C2029 diff_2476040_1887000# gnd! 38.4fF
C2030 diff_2450880_1887000# gnd! 38.4fF
C2031 diff_2425720_1887000# gnd! 38.4fF
C2032 diff_2400560_1887000# gnd! 38.4fF
C2033 diff_2375400_1887000# gnd! 38.4fF
C2034 diff_2350240_1887000# gnd! 38.4fF
C2035 diff_2325080_1887000# gnd! 38.4fF
C2036 diff_2299920_1887000# gnd! 38.4fF
C2037 diff_2274760_1887000# gnd! 38.4fF
C2038 diff_2249600_1887000# gnd! 38.4fF
C2039 diff_2224440_1887000# gnd! 38.4fF
C2040 diff_2199280_1887000# gnd! 38.4fF
C2041 diff_2174120_1887000# gnd! 38.4fF
C2042 diff_2148960_1887000# gnd! 38.4fF
C2043 diff_2123800_1887000# gnd! 38.4fF
C2044 diff_2098640_1887000# gnd! 38.4fF
C2045 diff_2073480_1887000# gnd! 38.4fF
C2046 diff_2048320_1887000# gnd! 38.4fF
C2047 diff_2023160_1887000# gnd! 38.4fF
C2048 diff_1998000_1887000# gnd! 38.4fF
C2049 diff_1972840_1887000# gnd! 38.4fF
C2050 diff_1947680_1887000# gnd! 38.4fF
C2051 diff_1922520_1887000# gnd! 38.4fF
C2052 diff_1897360_1887000# gnd! 38.4fF
C2053 diff_1872200_1887000# gnd! 38.4fF
C2054 diff_1847040_1887000# gnd! 38.4fF
C2055 diff_1821880_1887000# gnd! 38.4fF
C2056 diff_1796720_1887000# gnd! 38.4fF
C2057 diff_1771560_1887000# gnd! 38.4fF
C2058 diff_1746400_1887000# gnd! 38.4fF
C2059 diff_1721240_1887000# gnd! 38.4fF
C2060 diff_1696080_1887000# gnd! 38.4fF
C2061 diff_1670920_1887000# gnd! 38.4fF
C2062 diff_1645760_1887000# gnd! 38.4fF
C2063 diff_1620600_1887000# gnd! 38.4fF
C2064 diff_1595440_1887000# gnd! 38.4fF
C2065 diff_1570280_1887000# gnd! 38.4fF
C2066 diff_1545120_1887000# gnd! 38.4fF
C2067 diff_1519960_1887000# gnd! 38.4fF
C2068 diff_1494800_1887000# gnd! 38.4fF
C2069 diff_1469640_1887000# gnd! 38.4fF
C2070 diff_1444480_1887000# gnd! 38.4fF
C2071 diff_1419320_1887000# gnd! 38.4fF
C2072 diff_1394160_1887000# gnd! 38.4fF
C2073 diff_1369000_1887000# gnd! 38.4fF
C2074 diff_1343840_1887000# gnd! 38.4fF
C2075 diff_1318680_1887000# gnd! 38.4fF
C2076 diff_1293520_1887000# gnd! 38.4fF
C2077 diff_1268360_1887000# gnd! 38.4fF
C2078 diff_1243200_1887000# gnd! 38.4fF
C2079 diff_1238760_1907720# gnd! 974.7fF
C2080 diff_2828280_1915120# gnd! 36.1fF
C2081 diff_2803120_1915120# gnd! 36.1fF
C2082 diff_2777960_1915120# gnd! 36.1fF
C2083 diff_2752800_1915120# gnd! 36.1fF
C2084 diff_2727640_1915120# gnd! 36.1fF
C2085 diff_2702480_1915120# gnd! 36.1fF
C2086 diff_2677320_1915120# gnd! 36.1fF
C2087 diff_2652160_1915120# gnd! 36.1fF
C2088 diff_2627000_1915120# gnd! 36.1fF
C2089 diff_2601840_1915120# gnd! 36.1fF
C2090 diff_2576680_1915120# gnd! 36.1fF
C2091 diff_2551520_1915120# gnd! 36.1fF
C2092 diff_2526360_1915120# gnd! 36.1fF
C2093 diff_2501200_1915120# gnd! 36.1fF
C2094 diff_2476040_1915120# gnd! 36.1fF
C2095 diff_2450880_1915120# gnd! 36.1fF
C2096 diff_2425720_1915120# gnd! 36.1fF
C2097 diff_2400560_1915120# gnd! 36.1fF
C2098 diff_2375400_1915120# gnd! 36.1fF
C2099 diff_2350240_1915120# gnd! 36.1fF
C2100 diff_2325080_1915120# gnd! 36.1fF
C2101 diff_2299920_1915120# gnd! 36.1fF
C2102 diff_2274760_1915120# gnd! 36.1fF
C2103 diff_2249600_1915120# gnd! 36.1fF
C2104 diff_2224440_1915120# gnd! 36.1fF
C2105 diff_2199280_1915120# gnd! 36.1fF
C2106 diff_2174120_1915120# gnd! 36.1fF
C2107 diff_2148960_1915120# gnd! 36.1fF
C2108 diff_2123800_1915120# gnd! 36.1fF
C2109 diff_2098640_1915120# gnd! 36.1fF
C2110 diff_2073480_1915120# gnd! 36.1fF
C2111 diff_2048320_1915120# gnd! 36.1fF
C2112 diff_2023160_1915120# gnd! 36.1fF
C2113 diff_1998000_1915120# gnd! 36.1fF
C2114 diff_1972840_1915120# gnd! 36.1fF
C2115 diff_1947680_1915120# gnd! 36.1fF
C2116 diff_1922520_1915120# gnd! 36.1fF
C2117 diff_1897360_1915120# gnd! 36.1fF
C2118 diff_1872200_1915120# gnd! 36.1fF
C2119 diff_1847040_1915120# gnd! 36.1fF
C2120 diff_1821880_1915120# gnd! 36.1fF
C2121 diff_1796720_1915120# gnd! 36.1fF
C2122 diff_1771560_1915120# gnd! 36.1fF
C2123 diff_1746400_1915120# gnd! 36.1fF
C2124 diff_1721240_1915120# gnd! 36.1fF
C2125 diff_1696080_1915120# gnd! 36.1fF
C2126 diff_1670920_1915120# gnd! 36.1fF
C2127 diff_1645760_1915120# gnd! 36.1fF
C2128 diff_1620600_1915120# gnd! 36.1fF
C2129 diff_1595440_1915120# gnd! 36.1fF
C2130 diff_1570280_1915120# gnd! 36.1fF
C2131 diff_1545120_1915120# gnd! 36.1fF
C2132 diff_1519960_1915120# gnd! 36.1fF
C2133 diff_1494800_1915120# gnd! 36.1fF
C2134 diff_1469640_1915120# gnd! 36.1fF
C2135 diff_1444480_1915120# gnd! 36.1fF
C2136 diff_1419320_1915120# gnd! 36.1fF
C2137 diff_1394160_1915120# gnd! 36.1fF
C2138 diff_1369000_1915120# gnd! 36.1fF
C2139 diff_1343840_1915120# gnd! 36.1fF
C2140 diff_1318680_1915120# gnd! 36.1fF
C2141 diff_1293520_1915120# gnd! 36.1fF
C2142 diff_1268360_1915120# gnd! 36.1fF
C2143 diff_1243200_1915120# gnd! 36.1fF
C2144 diff_694120_1786360# gnd! 486.6fF
C2145 diff_503200_1786360# gnd! 532.9fF
C2146 diff_1238760_1934360# gnd! 977.0fF
C2147 diff_2920040_1955080# gnd! 747.3fF
C2148 diff_2828280_1941760# gnd! 38.4fF
C2149 diff_2803120_1941760# gnd! 38.4fF
C2150 diff_2777960_1941760# gnd! 38.4fF
C2151 diff_2752800_1941760# gnd! 38.4fF
C2152 diff_2727640_1941760# gnd! 38.4fF
C2153 diff_2702480_1941760# gnd! 38.4fF
C2154 diff_2677320_1941760# gnd! 38.4fF
C2155 diff_2652160_1941760# gnd! 38.4fF
C2156 diff_2627000_1941760# gnd! 38.4fF
C2157 diff_2601840_1941760# gnd! 38.4fF
C2158 diff_2576680_1941760# gnd! 38.4fF
C2159 diff_2551520_1941760# gnd! 38.4fF
C2160 diff_2526360_1941760# gnd! 38.4fF
C2161 diff_2501200_1941760# gnd! 38.4fF
C2162 diff_2476040_1941760# gnd! 38.4fF
C2163 diff_2450880_1941760# gnd! 38.4fF
C2164 diff_2425720_1941760# gnd! 38.4fF
C2165 diff_2400560_1941760# gnd! 38.4fF
C2166 diff_2375400_1941760# gnd! 38.4fF
C2167 diff_2350240_1941760# gnd! 38.4fF
C2168 diff_2325080_1941760# gnd! 38.4fF
C2169 diff_2299920_1941760# gnd! 38.4fF
C2170 diff_2274760_1941760# gnd! 38.4fF
C2171 diff_2249600_1941760# gnd! 38.4fF
C2172 diff_2224440_1941760# gnd! 38.4fF
C2173 diff_2199280_1941760# gnd! 38.4fF
C2174 diff_2174120_1941760# gnd! 38.4fF
C2175 diff_2148960_1941760# gnd! 38.4fF
C2176 diff_2123800_1941760# gnd! 38.4fF
C2177 diff_2098640_1941760# gnd! 38.4fF
C2178 diff_2073480_1941760# gnd! 38.4fF
C2179 diff_2048320_1941760# gnd! 38.4fF
C2180 diff_2023160_1941760# gnd! 38.4fF
C2181 diff_1998000_1941760# gnd! 38.4fF
C2182 diff_1972840_1941760# gnd! 38.4fF
C2183 diff_1947680_1941760# gnd! 38.4fF
C2184 diff_1922520_1941760# gnd! 38.4fF
C2185 diff_1897360_1941760# gnd! 38.4fF
C2186 diff_1872200_1941760# gnd! 38.4fF
C2187 diff_1847040_1941760# gnd! 38.4fF
C2188 diff_1821880_1941760# gnd! 38.4fF
C2189 diff_1796720_1941760# gnd! 38.4fF
C2190 diff_1771560_1941760# gnd! 38.4fF
C2191 diff_1746400_1941760# gnd! 38.4fF
C2192 diff_1721240_1941760# gnd! 38.4fF
C2193 diff_1696080_1941760# gnd! 38.4fF
C2194 diff_1670920_1941760# gnd! 38.4fF
C2195 diff_1645760_1941760# gnd! 38.4fF
C2196 diff_1620600_1941760# gnd! 38.4fF
C2197 diff_1595440_1941760# gnd! 38.4fF
C2198 diff_1570280_1941760# gnd! 38.4fF
C2199 diff_1545120_1941760# gnd! 38.4fF
C2200 diff_1519960_1941760# gnd! 38.4fF
C2201 diff_1494800_1941760# gnd! 38.4fF
C2202 diff_1469640_1941760# gnd! 38.4fF
C2203 diff_1444480_1941760# gnd! 38.4fF
C2204 diff_1419320_1941760# gnd! 38.4fF
C2205 diff_1394160_1941760# gnd! 38.4fF
C2206 diff_1369000_1941760# gnd! 38.4fF
C2207 diff_1343840_1941760# gnd! 38.4fF
C2208 diff_1318680_1941760# gnd! 38.4fF
C2209 diff_1293520_1941760# gnd! 38.4fF
C2210 diff_1268360_1941760# gnd! 38.4fF
C2211 diff_1243200_1941760# gnd! 38.4fF
C2212 diff_1238760_1962480# gnd! 907.6fF
C2213 diff_2828280_1969880# gnd! 36.1fF
C2214 diff_2803120_1969880# gnd! 36.1fF
C2215 diff_2777960_1969880# gnd! 36.1fF
C2216 diff_2752800_1969880# gnd! 36.1fF
C2217 diff_2727640_1969880# gnd! 36.1fF
C2218 diff_2702480_1969880# gnd! 36.1fF
C2219 diff_2677320_1969880# gnd! 36.1fF
C2220 diff_2652160_1969880# gnd! 36.1fF
C2221 diff_2627000_1969880# gnd! 36.1fF
C2222 diff_2601840_1969880# gnd! 36.1fF
C2223 diff_2576680_1969880# gnd! 36.1fF
C2224 diff_2551520_1969880# gnd! 36.1fF
C2225 diff_2526360_1969880# gnd! 36.1fF
C2226 diff_2501200_1969880# gnd! 36.1fF
C2227 diff_2476040_1969880# gnd! 36.1fF
C2228 diff_2450880_1969880# gnd! 36.1fF
C2229 diff_2425720_1969880# gnd! 36.1fF
C2230 diff_2400560_1969880# gnd! 36.1fF
C2231 diff_2375400_1969880# gnd! 36.1fF
C2232 diff_2350240_1969880# gnd! 36.1fF
C2233 diff_2325080_1969880# gnd! 36.1fF
C2234 diff_2299920_1969880# gnd! 36.1fF
C2235 diff_2274760_1969880# gnd! 36.1fF
C2236 diff_2249600_1969880# gnd! 36.1fF
C2237 diff_2224440_1969880# gnd! 36.1fF
C2238 diff_2199280_1969880# gnd! 36.1fF
C2239 diff_2174120_1969880# gnd! 36.1fF
C2240 diff_2148960_1969880# gnd! 36.1fF
C2241 diff_2123800_1969880# gnd! 36.1fF
C2242 diff_2098640_1969880# gnd! 36.1fF
C2243 diff_2073480_1969880# gnd! 36.1fF
C2244 diff_2048320_1969880# gnd! 36.1fF
C2245 diff_2023160_1969880# gnd! 36.1fF
C2246 diff_1998000_1969880# gnd! 36.1fF
C2247 diff_1972840_1969880# gnd! 36.1fF
C2248 diff_1947680_1969880# gnd! 36.1fF
C2249 diff_1922520_1969880# gnd! 36.1fF
C2250 diff_1897360_1969880# gnd! 36.1fF
C2251 diff_1872200_1969880# gnd! 36.1fF
C2252 diff_1847040_1969880# gnd! 36.1fF
C2253 diff_1821880_1969880# gnd! 36.1fF
C2254 diff_1796720_1969880# gnd! 36.1fF
C2255 diff_1771560_1969880# gnd! 36.1fF
C2256 diff_1746400_1969880# gnd! 36.1fF
C2257 diff_1721240_1969880# gnd! 36.1fF
C2258 diff_1696080_1969880# gnd! 36.1fF
C2259 diff_1670920_1969880# gnd! 36.1fF
C2260 diff_1645760_1969880# gnd! 36.1fF
C2261 diff_1620600_1969880# gnd! 36.1fF
C2262 diff_1595440_1969880# gnd! 36.1fF
C2263 diff_1570280_1969880# gnd! 36.1fF
C2264 diff_1545120_1969880# gnd! 36.1fF
C2265 diff_1519960_1969880# gnd! 36.1fF
C2266 diff_1494800_1969880# gnd! 36.1fF
C2267 diff_1469640_1969880# gnd! 36.1fF
C2268 diff_1444480_1969880# gnd! 36.1fF
C2269 diff_1419320_1969880# gnd! 36.1fF
C2270 diff_1394160_1969880# gnd! 36.1fF
C2271 diff_1369000_1969880# gnd! 36.1fF
C2272 diff_1343840_1969880# gnd! 36.1fF
C2273 diff_1318680_1969880# gnd! 36.1fF
C2274 diff_1293520_1969880# gnd! 36.1fF
C2275 diff_1268360_1969880# gnd! 36.1fF
C2276 diff_1243200_1969880# gnd! 36.1fF
C2277 diff_1238760_1989120# gnd! 925.4fF
C2278 diff_2828280_1996520# gnd! 38.4fF
C2279 diff_2803120_1996520# gnd! 38.4fF
C2280 diff_2777960_1996520# gnd! 38.4fF
C2281 diff_2752800_1996520# gnd! 38.4fF
C2282 diff_2727640_1996520# gnd! 38.4fF
C2283 diff_2702480_1996520# gnd! 38.4fF
C2284 diff_2677320_1996520# gnd! 38.4fF
C2285 diff_2652160_1996520# gnd! 38.4fF
C2286 diff_2627000_1996520# gnd! 38.4fF
C2287 diff_2601840_1996520# gnd! 38.4fF
C2288 diff_2576680_1996520# gnd! 38.4fF
C2289 diff_2551520_1996520# gnd! 38.4fF
C2290 diff_2526360_1996520# gnd! 38.4fF
C2291 diff_2501200_1996520# gnd! 38.4fF
C2292 diff_2476040_1996520# gnd! 38.4fF
C2293 diff_2450880_1996520# gnd! 38.4fF
C2294 diff_2425720_1996520# gnd! 38.4fF
C2295 diff_2400560_1996520# gnd! 38.4fF
C2296 diff_2375400_1996520# gnd! 38.4fF
C2297 diff_2350240_1996520# gnd! 38.4fF
C2298 diff_2325080_1996520# gnd! 38.4fF
C2299 diff_2299920_1996520# gnd! 38.4fF
C2300 diff_2274760_1996520# gnd! 38.4fF
C2301 diff_2249600_1996520# gnd! 38.4fF
C2302 diff_2224440_1996520# gnd! 38.4fF
C2303 diff_2199280_1996520# gnd! 38.4fF
C2304 diff_2174120_1996520# gnd! 38.4fF
C2305 diff_2148960_1996520# gnd! 38.4fF
C2306 diff_2123800_1996520# gnd! 38.4fF
C2307 diff_2098640_1996520# gnd! 38.4fF
C2308 diff_2073480_1996520# gnd! 38.4fF
C2309 diff_2048320_1996520# gnd! 38.4fF
C2310 diff_2023160_1996520# gnd! 38.4fF
C2311 diff_1998000_1996520# gnd! 38.4fF
C2312 diff_1972840_1996520# gnd! 38.4fF
C2313 diff_1947680_1996520# gnd! 38.4fF
C2314 diff_1922520_1996520# gnd! 38.4fF
C2315 diff_1897360_1996520# gnd! 38.4fF
C2316 diff_1872200_1996520# gnd! 38.4fF
C2317 diff_1847040_1996520# gnd! 38.4fF
C2318 diff_1821880_1996520# gnd! 38.4fF
C2319 diff_1796720_1996520# gnd! 38.4fF
C2320 diff_1771560_1996520# gnd! 38.4fF
C2321 diff_1746400_1996520# gnd! 38.4fF
C2322 diff_1721240_1996520# gnd! 38.4fF
C2323 diff_1696080_1996520# gnd! 38.4fF
C2324 diff_1670920_1996520# gnd! 38.4fF
C2325 diff_1645760_1996520# gnd! 38.4fF
C2326 diff_1620600_1996520# gnd! 38.4fF
C2327 diff_1595440_1996520# gnd! 38.4fF
C2328 diff_1570280_1996520# gnd! 38.4fF
C2329 diff_1545120_1996520# gnd! 38.4fF
C2330 diff_1519960_1996520# gnd! 38.4fF
C2331 diff_1494800_1996520# gnd! 38.4fF
C2332 diff_1469640_1996520# gnd! 38.4fF
C2333 diff_1444480_1996520# gnd! 38.4fF
C2334 diff_1419320_1996520# gnd! 38.4fF
C2335 diff_1394160_1996520# gnd! 38.4fF
C2336 diff_1369000_1996520# gnd! 38.4fF
C2337 diff_1343840_1996520# gnd! 38.4fF
C2338 diff_1318680_1996520# gnd! 38.4fF
C2339 diff_1293520_1996520# gnd! 38.4fF
C2340 diff_1268360_1996520# gnd! 38.4fF
C2341 diff_1243200_1996520# gnd! 38.4fF
C2342 diff_1238760_2017240# gnd! 973.6fF
C2343 diff_2828280_2024640# gnd! 36.1fF
C2344 diff_2803120_2024640# gnd! 36.1fF
C2345 diff_2777960_2024640# gnd! 36.1fF
C2346 diff_2752800_2024640# gnd! 36.1fF
C2347 diff_2727640_2024640# gnd! 36.1fF
C2348 diff_2702480_2024640# gnd! 36.1fF
C2349 diff_2677320_2024640# gnd! 36.1fF
C2350 diff_2652160_2024640# gnd! 36.1fF
C2351 diff_2627000_2024640# gnd! 36.1fF
C2352 diff_2601840_2024640# gnd! 36.1fF
C2353 diff_2576680_2024640# gnd! 36.1fF
C2354 diff_2551520_2024640# gnd! 36.1fF
C2355 diff_2526360_2024640# gnd! 36.1fF
C2356 diff_2501200_2024640# gnd! 36.1fF
C2357 diff_2476040_2024640# gnd! 36.1fF
C2358 diff_2450880_2024640# gnd! 36.1fF
C2359 diff_2425720_2024640# gnd! 36.1fF
C2360 diff_2400560_2024640# gnd! 36.1fF
C2361 diff_2375400_2024640# gnd! 36.1fF
C2362 diff_2350240_2024640# gnd! 36.1fF
C2363 diff_2325080_2024640# gnd! 36.1fF
C2364 diff_2299920_2024640# gnd! 36.1fF
C2365 diff_2274760_2024640# gnd! 36.1fF
C2366 diff_2249600_2024640# gnd! 36.1fF
C2367 diff_2224440_2024640# gnd! 36.1fF
C2368 diff_2199280_2024640# gnd! 36.1fF
C2369 diff_2174120_2024640# gnd! 36.1fF
C2370 diff_2148960_2024640# gnd! 36.1fF
C2371 diff_2123800_2024640# gnd! 36.1fF
C2372 diff_2098640_2024640# gnd! 36.1fF
C2373 diff_2073480_2024640# gnd! 36.1fF
C2374 diff_2048320_2024640# gnd! 36.1fF
C2375 diff_2023160_2024640# gnd! 36.1fF
C2376 diff_1998000_2024640# gnd! 36.1fF
C2377 diff_1972840_2024640# gnd! 36.1fF
C2378 diff_1947680_2024640# gnd! 36.1fF
C2379 diff_1922520_2024640# gnd! 36.1fF
C2380 diff_1897360_2024640# gnd! 36.1fF
C2381 diff_1872200_2024640# gnd! 36.1fF
C2382 diff_1847040_2024640# gnd! 36.1fF
C2383 diff_1821880_2024640# gnd! 36.1fF
C2384 diff_1796720_2024640# gnd! 36.1fF
C2385 diff_1771560_2024640# gnd! 36.1fF
C2386 diff_1746400_2024640# gnd! 36.1fF
C2387 diff_1721240_2024640# gnd! 36.1fF
C2388 diff_1696080_2024640# gnd! 36.1fF
C2389 diff_1670920_2024640# gnd! 36.1fF
C2390 diff_1645760_2024640# gnd! 36.1fF
C2391 diff_1620600_2024640# gnd! 36.1fF
C2392 diff_1595440_2024640# gnd! 36.1fF
C2393 diff_1570280_2024640# gnd! 36.1fF
C2394 diff_1545120_2024640# gnd! 36.1fF
C2395 diff_1519960_2024640# gnd! 36.1fF
C2396 diff_1494800_2024640# gnd! 36.1fF
C2397 diff_1469640_2024640# gnd! 36.1fF
C2398 diff_1444480_2024640# gnd! 36.1fF
C2399 diff_1419320_2024640# gnd! 36.1fF
C2400 diff_1394160_2024640# gnd! 36.1fF
C2401 diff_1369000_2024640# gnd! 36.1fF
C2402 diff_1343840_2024640# gnd! 36.1fF
C2403 diff_1318680_2024640# gnd! 36.1fF
C2404 diff_1293520_2024640# gnd! 36.1fF
C2405 diff_1268360_2024640# gnd! 36.1fF
C2406 diff_1243200_2024640# gnd! 36.1fF
C2407 diff_1093720_1907720# gnd! 132.3fF
C2408 diff_1025640_1855920# gnd! 135.7fF
C2409 diff_1012320_1684240# gnd! 912.9fF
C2410 diff_910200_1857400# gnd! 132.8fF
C2411 diff_830280_1857400# gnd! 146.3fF
C2412 diff_819920_1684240# gnd! 898.7fF
C2413 diff_233840_991600# gnd! 2583.8fF
C2414 diff_719280_1857400# gnd! 142.0fF
C2415 diff_642320_1854440# gnd! 134.8fF
C2416 diff_629000_1685720# gnd! 916.9fF
C2417 diff_528360_1858880# gnd! 136.3fF
C2418 diff_451400_1855920# gnd! 141.4fF
C2419 diff_1238760_2043880# gnd! 970.6fF
C2420 diff_3090240_1133680# gnd! 630.9fF
C2421 diff_3069520_1052280# gnd! 858.8fF
C2422 diff_2920040_2064600# gnd! 740.5fF
C2423 diff_2828280_2051280# gnd! 38.4fF
C2424 diff_2803120_2051280# gnd! 38.4fF
C2425 diff_2777960_2051280# gnd! 38.4fF
C2426 diff_2752800_2051280# gnd! 38.4fF
C2427 diff_2727640_2051280# gnd! 38.4fF
C2428 diff_2702480_2051280# gnd! 38.4fF
C2429 diff_2677320_2051280# gnd! 38.4fF
C2430 diff_2652160_2051280# gnd! 38.4fF
C2431 diff_2627000_2051280# gnd! 38.4fF
C2432 diff_2601840_2051280# gnd! 38.4fF
C2433 diff_2576680_2051280# gnd! 38.4fF
C2434 diff_2551520_2051280# gnd! 38.4fF
C2435 diff_2526360_2051280# gnd! 38.4fF
C2436 diff_2501200_2051280# gnd! 38.4fF
C2437 diff_2476040_2051280# gnd! 38.4fF
C2438 diff_2450880_2051280# gnd! 38.4fF
C2439 diff_2425720_2051280# gnd! 38.4fF
C2440 diff_2400560_2051280# gnd! 38.4fF
C2441 diff_2375400_2051280# gnd! 38.4fF
C2442 diff_2350240_2051280# gnd! 38.4fF
C2443 diff_2325080_2051280# gnd! 38.4fF
C2444 diff_2299920_2051280# gnd! 38.4fF
C2445 diff_2274760_2051280# gnd! 38.4fF
C2446 diff_2249600_2051280# gnd! 38.4fF
C2447 diff_2224440_2051280# gnd! 38.4fF
C2448 diff_2199280_2051280# gnd! 38.4fF
C2449 diff_2174120_2051280# gnd! 38.4fF
C2450 diff_2148960_2051280# gnd! 38.4fF
C2451 diff_2123800_2051280# gnd! 38.4fF
C2452 diff_2098640_2051280# gnd! 38.4fF
C2453 diff_2073480_2051280# gnd! 38.4fF
C2454 diff_2048320_2051280# gnd! 38.4fF
C2455 diff_2023160_2051280# gnd! 38.4fF
C2456 diff_1998000_2051280# gnd! 38.4fF
C2457 diff_1972840_2051280# gnd! 38.4fF
C2458 diff_1947680_2051280# gnd! 38.4fF
C2459 diff_1922520_2051280# gnd! 38.4fF
C2460 diff_1897360_2051280# gnd! 38.4fF
C2461 diff_1872200_2051280# gnd! 38.4fF
C2462 diff_1847040_2051280# gnd! 38.4fF
C2463 diff_1821880_2051280# gnd! 38.4fF
C2464 diff_1796720_2051280# gnd! 38.4fF
C2465 diff_1771560_2051280# gnd! 38.4fF
C2466 diff_1746400_2051280# gnd! 38.4fF
C2467 diff_1721240_2051280# gnd! 38.4fF
C2468 diff_1696080_2051280# gnd! 38.4fF
C2469 diff_1670920_2051280# gnd! 38.4fF
C2470 diff_1645760_2051280# gnd! 38.4fF
C2471 diff_1620600_2051280# gnd! 38.4fF
C2472 diff_1595440_2051280# gnd! 38.4fF
C2473 diff_1570280_2051280# gnd! 38.4fF
C2474 diff_1545120_2051280# gnd! 38.4fF
C2475 diff_1519960_2051280# gnd! 38.4fF
C2476 diff_1494800_2051280# gnd! 38.4fF
C2477 diff_1469640_2051280# gnd! 38.4fF
C2478 diff_1444480_2051280# gnd! 38.4fF
C2479 diff_1419320_2051280# gnd! 38.4fF
C2480 diff_1394160_2051280# gnd! 38.4fF
C2481 diff_1369000_2051280# gnd! 38.4fF
C2482 diff_1343840_2051280# gnd! 38.4fF
C2483 diff_1318680_2051280# gnd! 38.4fF
C2484 diff_1293520_2051280# gnd! 38.4fF
C2485 diff_1268360_2051280# gnd! 38.4fF
C2486 diff_1243200_2051280# gnd! 38.4fF
C2487 diff_1238760_2072000# gnd! 917.2fF
C2488 diff_2998480_1207680# gnd! 1057.6fF
C2489 diff_2976280_1228400# gnd! 1117.1fF
C2490 diff_2940760_526880# gnd! 873.4fF
C2491 diff_2912640_526880# gnd! 913.9fF
C2492 diff_1243200_2079400# gnd! 1412.9fF
C2493 diff_2043880_2100120# gnd! 1441.3fF
C2494 diff_3285600_2079400# gnd! 227.5fF
C2495 diff_3267840_1761200# gnd! 445.2fF
C2496 diff_3223440_2120840# gnd! 356.7fF
C2497 diff_3005880_2094200# gnd! 1310.0fF
C2498 diff_1237280_2100120# gnd! 1110.8fF
C2499 diff_3001440_2148960# gnd! 1224.7fF
C2500 diff_3393640_2079400# gnd! 189.6fF
C2501 diff_3455800_2137120# gnd! 149.1fF
C2502 diff_991600_2049800# gnd! 1447.1fF
C2503 diff_800680_2049800# gnd! 1450.3fF
C2504 Vdd gnd! 23696.8fF
C2505 diff_438080_1685720# gnd! 916.9fF
C2506 diff_609760_2049800# gnd! 1465.9fF
C2507 diff_417360_2049800# gnd! 1464.8fF
C2508 d0 gnd! 3114.4fF
C2509 d1 gnd! 3416.0fF
C2510 d3 gnd! 4969.7fF
C2511 sync gnd! 2859.3fF
C2512 d2 gnd! 3698.9fF
C2513 clk1 gnd! 3035.7fF
C2514 clk2 gnd! 4412.4fF
