* SPICE3 file created from 4002.ext - technology: nmos

.option scale=0.001u

M1000 diff_289200_2884800# diff_358800_2898000# GND GND efet w=77400 l=7200
+ ad=-1.31993e+09 pd=585600 as=8.96681e+08 ps=7.19088e+07 
M1001 d1 GND GND GND efet w=105600 l=8400
+ ad=7.42371e+08 pd=3.0336e+06 as=0 ps=0 
M1002 GND diff_87600_2288400# diff_289200_2884800# GND efet w=215400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1003 GND d1 diff_97200_2845200# GND efet w=55800 l=6600
+ ad=0 pd=0 as=1.31616e+09 ps=290400 
M1004 GND diff_87600_2288400# diff_358800_2898000# GND efet w=223200 l=6600
+ ad=0 pd=0 as=-4.22807e+08 ps=760800 
M1005 diff_358800_2898000# diff_457200_2878800# GND GND efet w=211800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1006 diff_289200_2884800# diff_289200_2857200# diff_289200_2884800# GND efet w=40200 l=13200
+ ad=0 pd=0 as=0 ps=0 
M1007 GND diff_97200_2845200# diff_165600_2822400# GND efet w=22200 l=7800
+ ad=0 pd=0 as=1.43856e+09 ps=273600 
M1008 diff_97200_2845200# diff_97200_2845200# diff_97200_2845200# GND efet w=2400 l=4800
+ ad=0 pd=0 as=0 ps=0 
M1009 diff_97200_2845200# diff_97200_2845200# diff_97200_2845200# GND efet w=1800 l=1800
+ ad=0 pd=0 as=0 ps=0 
M1010 diff_165600_2822400# diff_165600_2822400# diff_165600_2822400# GND efet w=3600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M1011 diff_165600_2822400# diff_165600_2822400# diff_165600_2822400# GND efet w=1200 l=4800
+ ad=0 pd=0 as=0 ps=0 
M1012 diff_97200_2845200# Vdd Vdd GND efet w=9600 l=35400
+ ad=0 pd=0 as=5.66981e+08 ps=3.49416e+07 
M1013 GND diff_132000_2799600# diff_97200_2845200# GND efet w=34800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1014 diff_165600_2822400# diff_132000_2799600# GND GND efet w=36600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1015 GND diff_289200_2884800# d1 GND efet w=1123800 l=4200
+ ad=0 pd=0 as=0 ps=0 
M1016 diff_358800_2898000# diff_386400_2857200# diff_358800_2898000# GND efet w=42600 l=13200
+ ad=0 pd=0 as=0 ps=0 
M1017 diff_289200_2884800# diff_289200_2857200# Vdd GND efet w=11400 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1018 diff_289200_2857200# diff_289200_2857200# diff_289200_2857200# GND efet w=3000 l=4200
+ ad=2.2032e+08 pd=76800 as=0 ps=0 
M1019 diff_289200_2857200# diff_289200_2857200# diff_289200_2857200# GND efet w=1800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1020 diff_358800_2898000# diff_386400_2857200# Vdd GND efet w=11400 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1021 diff_386400_2857200# diff_386400_2857200# diff_386400_2857200# GND efet w=3000 l=4200
+ ad=2.1168e+08 pd=72000 as=0 ps=0 
M1022 diff_386400_2857200# diff_386400_2857200# diff_386400_2857200# GND efet w=1800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1023 diff_289200_2857200# Vdd Vdd GND efet w=9600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1024 Vdd Vdd Vdd GND efet w=2400 l=4800
+ ad=0 pd=0 as=0 ps=0 
M1025 Vdd Vdd Vdd GND efet w=1200 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1026 Vdd Vdd diff_165600_2822400# GND efet w=8400 l=37800
+ ad=0 pd=0 as=0 ps=0 
M1027 diff_252000_2766000# diff_165600_2822400# Vdd GND efet w=38400 l=9600
+ ad=1.38458e+08 pd=2.8128e+06 as=0 ps=0 
M1028 GND diff_97200_2845200# diff_252000_2766000# GND efet w=38400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1029 d0 GND GND GND efet w=108000 l=8400
+ ad=2.57091e+08 pd=3.0504e+06 as=0 ps=0 
M1030 GND diff_87600_2288400# diff_1262400_2888400# GND efet w=211200 l=7200
+ ad=0 pd=0 as=-1.32857e+09 ps=578400 
M1031 GND d0 diff_943200_2844000# GND efet w=55200 l=7200
+ ad=0 pd=0 as=1.27728e+09 ps=285600 
M1032 diff_1262400_2888400# diff_1330800_2899200# GND GND efet w=75600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1033 GND diff_87600_2288400# diff_1330800_2899200# GND efet w=217800 l=7800
+ ad=0 pd=0 as=-4.64567e+08 ps=717600 
M1034 diff_1330800_2899200# diff_1429200_2878800# GND GND efet w=212400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1035 GND diff_943200_2844000# diff_1009200_2812800# GND efet w=21600 l=7200
+ ad=0 pd=0 as=1.46016e+09 ps=288000 
M1036 diff_943200_2844000# diff_943200_2844000# diff_943200_2844000# GND efet w=2400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M1037 diff_1009200_2812800# diff_1009200_2812800# diff_1009200_2812800# GND efet w=6000 l=4800
+ ad=0 pd=0 as=0 ps=0 
M1038 d1 diff_358800_2898000# Vdd GND efet w=606000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1039 diff_457200_2878800# diff_457200_2878800# diff_457200_2878800# GND efet w=2400 l=9600
+ ad=9.9648e+08 pd=223200 as=0 ps=0 
M1040 diff_386400_2857200# Vdd Vdd GND efet w=8400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1041 diff_457200_2878800# diff_457200_2878800# diff_457200_2878800# GND efet w=3000 l=4800
+ ad=0 pd=0 as=0 ps=0 
M1042 diff_1009200_2812800# diff_1009200_2812800# diff_1009200_2812800# GND efet w=1800 l=5400
+ ad=0 pd=0 as=0 ps=0 
M1043 diff_943200_2844000# Vdd Vdd GND efet w=9000 l=35400
+ ad=0 pd=0 as=0 ps=0 
M1044 GND diff_132000_2799600# diff_943200_2844000# GND efet w=34800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1045 diff_1009200_2812800# diff_132000_2799600# GND GND efet w=34800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1046 diff_1262400_2888400# diff_1261200_2857200# diff_1262400_2888400# GND efet w=36600 l=31800
+ ad=0 pd=0 as=0 ps=0 
M1047 GND diff_1262400_2888400# d0 GND efet w=1115400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M1048 diff_1330800_2899200# diff_1358400_2856000# diff_1330800_2899200# GND efet w=34200 l=33600
+ ad=0 pd=0 as=0 ps=0 
M1049 o0 diff_1916400_2860800# GND GND efet w=198000 l=7200
+ ad=-4.61687e+08 pd=691200 as=0 ps=0 
M1050 diff_1916400_2860800# diff_2017200_2959200# GND GND efet w=110400 l=7200
+ ad=1.37088e+09 pd=283200 as=0 ps=0 
M1051 diff_1923600_2864400# diff_1916400_2860800# GND GND efet w=48000 l=7200
+ ad=9.3744e+08 pd=172800 as=0 ps=0 
M1052 diff_2016000_2904000# diff_1916400_2860800# GND GND efet w=24000 l=7200
+ ad=5.6736e+08 pd=136800 as=0 ps=0 
M1053 diff_2017200_2959200# diff_2050800_2889600# diff_2016000_2904000# GND efet w=13200 l=7200
+ ad=1.47024e+09 pd=319200 as=0 ps=0 
M1054 GND diff_2077200_2900400# diff_2017200_2959200# GND efet w=25200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1055 diff_1923600_2864400# diff_1923600_2864400# diff_1923600_2864400# GND efet w=3600 l=4800
+ ad=0 pd=0 as=0 ps=0 
M1056 diff_1923600_2864400# diff_1923600_2864400# diff_1923600_2864400# GND efet w=1200 l=2400
+ ad=0 pd=0 as=0 ps=0 
M1057 o0 diff_1923600_2864400# Vdd GND efet w=211800 l=6600
+ ad=0 pd=0 as=0 ps=0 
M1058 d0 diff_1330800_2899200# Vdd GND efet w=609000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1059 diff_1262400_2888400# diff_1261200_2857200# Vdd GND efet w=10200 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1060 diff_1261200_2857200# diff_1261200_2857200# diff_1261200_2857200# GND efet w=2400 l=4200
+ ad=2.1024e+08 pd=69600 as=0 ps=0 
M1061 diff_1261200_2857200# diff_1261200_2857200# diff_1261200_2857200# GND efet w=1200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M1062 diff_1358400_2856000# diff_1358400_2856000# diff_1358400_2856000# GND efet w=2400 l=4200
+ ad=1.9728e+08 pd=67200 as=0 ps=0 
M1063 diff_1358400_2856000# diff_1358400_2856000# diff_1358400_2856000# GND efet w=1800 l=5400
+ ad=0 pd=0 as=0 ps=0 
M1064 Vdd Vdd Vdd GND efet w=2400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M1065 diff_457200_2878800# diff_222000_1082400# diff_252000_2766000# GND efet w=29400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1066 Vdd Vdd diff_1009200_2812800# GND efet w=8400 l=37200
+ ad=0 pd=0 as=0 ps=0 
M1067 diff_349200_1096800# diff_1009200_2812800# Vdd GND efet w=37200 l=7200
+ ad=-1.0409e+09 pd=2.4816e+06 as=0 ps=0 
M1068 GND diff_943200_2844000# diff_349200_1096800# GND efet w=39000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1069 diff_1261200_2857200# Vdd Vdd GND efet w=10200 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1070 diff_1330800_2899200# diff_1358400_2856000# Vdd GND efet w=9600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1071 Vdd Vdd diff_1358400_2856000# GND efet w=7800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1072 Vdd Vdd Vdd GND efet w=1200 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1073 diff_1923600_2864400# Vdd Vdd GND efet w=9600 l=19200
+ ad=0 pd=0 as=0 ps=0 
M1074 diff_2016000_2904000# Vdd Vdd GND efet w=7200 l=30000
+ ad=0 pd=0 as=0 ps=0 
M1075 GND diff_2074800_2772000# diff_2050800_2889600# GND efet w=13200 l=7200
+ ad=0 pd=0 as=2.9664e+08 ps=74400 
M1076 diff_2050800_2889600# Vdd Vdd GND efet w=7800 l=57000
+ ad=0 pd=0 as=0 ps=0 
M1077 Vdd Vdd Vdd GND efet w=4800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1078 Vdd Vdd Vdd GND efet w=5400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M1079 diff_1916400_2860800# Vdd Vdd GND efet w=11400 l=18600
+ ad=0 pd=0 as=0 ps=0 
M1080 GND diff_2415600_2852400# diff_2373600_2752800# GND efet w=49200 l=7200
+ ad=0 pd=0 as=1.15056e+09 ps=187200 
M1081 GND diff_2415600_2852400# o1 GND efet w=202800 l=6000
+ ad=0 pd=0 as=-1.70807e+08 ps=708000 
M1082 diff_2017200_2959200# diff_2074800_2772000# diff_2104800_2774400# GND efet w=19200 l=6600
+ ad=0 pd=0 as=2.88e+08 ps=79200 
M1083 Vdd diff_68400_2361600# d2 GND efet w=623400 l=6600
+ ad=0 pd=0 as=1.76045e+09 ps=3.0696e+06 
M1084 GND diff_69600_2534400# d2 GND efet w=1144200 l=4200
+ ad=0 pd=0 as=0 ps=0 
M1085 diff_1429200_2878800# diff_222000_1082400# diff_349200_1096800# GND efet w=26400 l=7200
+ ad=8.208e+08 pd=170400 as=0 ps=0 
M1086 diff_2104800_2774400# clk2 diff_349200_1096800# GND efet w=18000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1087 diff_2373600_2752800# Vdd Vdd GND efet w=10800 l=19200
+ ad=0 pd=0 as=0 ps=0 
M1088 diff_2373600_2752800# diff_2373600_2752800# diff_2373600_2752800# GND efet w=4200 l=4200
+ ad=0 pd=0 as=0 ps=0 
M1089 o1 diff_2373600_2752800# Vdd GND efet w=209400 l=6600
+ ad=0 pd=0 as=0 ps=0 
M1090 GND diff_2415600_2852400# diff_2454000_2737200# GND efet w=26400 l=8400
+ ad=0 pd=0 as=6.5952e+08 ps=146400 
M1091 diff_2454000_2737200# Vdd Vdd GND efet w=10800 l=28800
+ ad=0 pd=0 as=0 ps=0 
M1092 Vdd Vdd Vdd GND efet w=3600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1093 Vdd Vdd Vdd GND efet w=3600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1094 GND diff_2346000_2652000# diff_2415600_2852400# GND efet w=111600 l=5400
+ ad=0 pd=0 as=1.4112e+09 ps=276000 
M1095 diff_2454000_2737200# diff_2424000_2713200# diff_2346000_2652000# GND efet w=14400 l=8400
+ ad=0 pd=0 as=1.6344e+09 ps=326400 
M1096 diff_2424000_2713200# Vdd Vdd GND efet w=8400 l=57600
+ ad=3.456e+08 pd=79200 as=0 ps=0 
M1097 diff_2424000_2713200# diff_2074800_2772000# GND GND efet w=15000 l=6600
+ ad=0 pd=0 as=0 ps=0 
M1098 diff_2346000_2652000# diff_2077200_2900400# GND GND efet w=25200 l=6600
+ ad=0 pd=0 as=0 ps=0 
M1099 Vdd Vdd Vdd GND efet w=3000 l=4200
+ ad=0 pd=0 as=0 ps=0 
M1100 Vdd Vdd Vdd GND efet w=2400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1101 diff_487200_2602800# diff_326400_2457600# diff_349200_1096800# GND efet w=38400 l=7200
+ ad=9.8928e+08 pd=228000 as=0 ps=0 
M1102 diff_487200_2602800# diff_523200_1467600# diff_506400_2604000# GND efet w=38400 l=7200
+ ad=0 pd=0 as=1.73808e+09 ps=340800 
M1103 diff_548400_2601600# diff_426000_1591200# diff_487200_2602800# GND efet w=46200 l=7800
+ ad=-1.12121e+09 pd=864000 as=0 ps=0 
M1104 diff_2325600_2644800# clk2 diff_252000_2766000# GND efet w=20400 l=7200
+ ad=3.2112e+08 pd=81600 as=0 ps=0 
M1105 diff_2346000_2652000# diff_2074800_2772000# diff_2325600_2644800# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1106 diff_567600_2590800# Vdd Vdd GND efet w=8400 l=30000
+ ad=9.1872e+08 pd=225600 as=0 ps=0 
M1107 Vdd diff_663600_2611200# diff_506400_2604000# GND efet w=15600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1108 diff_567600_2590800# diff_423600_2420400# diff_548400_2601600# GND efet w=32400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1109 diff_487200_2554800# diff_326400_2457600# diff_252000_2766000# GND efet w=38400 l=7200
+ ad=9.8928e+08 pd=228000 as=0 ps=0 
M1110 diff_567600_2553600# diff_423600_2420400# diff_548400_2534400# GND efet w=31800 l=7800
+ ad=9.216e+08 pd=218400 as=-1.08521e+09 ps=885600 
M1111 diff_506400_2604000# diff_567600_2590800# GND GND efet w=55200 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1112 diff_567600_2590800# diff_663600_2611200# GND GND efet w=27000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1113 GND diff_567600_2553600# diff_506400_2533200# GND efet w=54000 l=8400
+ ad=0 pd=0 as=1.7352e+09 ps=333600 
M1114 diff_813600_2584800# diff_804000_2611200# GND GND efet w=22800 l=7200
+ ad=2.4048e+08 pd=72000 as=0 ps=0 
M1115 diff_548400_2601600# diff_843600_1497600# diff_804000_2611200# GND efet w=9600 l=7200
+ ad=0 pd=0 as=2.6928e+08 ps=74400 
M1116 diff_880800_2613600# diff_872400_1458000# diff_548400_2601600# GND efet w=9600 l=7200
+ ad=2.6208e+08 pd=74400 as=0 ps=0 
M1117 diff_663600_2611200# diff_807600_1443600# diff_813600_2584800# GND efet w=21600 l=8400
+ ad=-2.11857e+09 pd=1.5408e+06 as=0 ps=0 
M1118 diff_664800_2534400# diff_807600_1443600# diff_813600_2542800# GND efet w=22200 l=9600
+ ad=1.88839e+09 pd=1.548e+06 as=2.4192e+08 ps=74400 
M1119 diff_68400_2361600# diff_87600_2492400# GND GND efet w=215400 l=6600
+ ad=-3.53687e+08 pd=787200 as=0 ps=0 
M1120 diff_87600_2492400# diff_87600_2492400# diff_87600_2492400# GND efet w=1800 l=6600
+ ad=1.1592e+09 pd=218400 as=0 ps=0 
M1121 diff_87600_2492400# diff_87600_2492400# diff_87600_2492400# GND efet w=3000 l=4200
+ ad=0 pd=0 as=0 ps=0 
M1122 diff_230400_2126400# diff_222000_1082400# diff_87600_2492400# GND efet w=27600 l=7200
+ ad=-1.05242e+09 pd=2.484e+06 as=0 ps=0 
M1123 diff_487200_2491200# diff_326400_2457600# diff_230400_2126400# GND efet w=38400 l=7200
+ ad=9.6048e+08 pd=228000 as=0 ps=0 
M1124 diff_487200_2554800# diff_523200_1467600# diff_506400_2533200# GND efet w=38400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1125 diff_548400_2534400# diff_426000_1591200# diff_487200_2554800# GND efet w=45000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1126 GND diff_664800_2534400# diff_567600_2553600# GND efet w=26400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1127 GND diff_326400_2457600# diff_440400_2446800# GND efet w=52200 l=7800
+ ad=0 pd=0 as=5.7456e+08 ps=127200 
M1128 diff_487200_2491200# diff_523200_1467600# diff_506400_2467200# GND efet w=37200 l=7200
+ ad=0 pd=0 as=1.7136e+09 ps=324000 
M1129 diff_548400_2460000# diff_426000_1591200# diff_487200_2491200# GND efet w=45000 l=7800
+ ad=-1.17881e+09 pd=859200 as=0 ps=0 
M1130 Vdd diff_664800_2534400# diff_506400_2533200# GND efet w=15000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1131 diff_813600_2542800# diff_804000_2528400# GND GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1132 diff_567600_2553600# Vdd Vdd GND efet w=7200 l=27600
+ ad=0 pd=0 as=0 ps=0 
M1133 Vdd Vdd Vdd GND efet w=6000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M1134 Vdd Vdd Vdd GND efet w=4200 l=11400
+ ad=0 pd=0 as=0 ps=0 
M1135 diff_567600_2450400# Vdd Vdd GND efet w=7200 l=27600
+ ad=9.6912e+08 pd=232800 as=0 ps=0 
M1136 diff_567600_2450400# diff_423600_2420400# diff_548400_2460000# GND efet w=32400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1137 diff_440400_2446800# diff_426000_1591200# diff_423600_2420400# GND efet w=48600 l=7800
+ ad=0 pd=0 as=9.864e+08 ps=204000 
M1138 diff_68400_2361600# diff_87600_2288400# GND GND efet w=215400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1139 Vdd diff_162000_2388000# diff_68400_2361600# GND efet w=10800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1140 Vdd Vdd diff_423600_2420400# GND efet w=12000 l=39000
+ ad=0 pd=0 as=0 ps=0 
M1141 diff_68400_2361600# diff_162000_2388000# diff_68400_2361600# GND efet w=48600 l=18000
+ ad=0 pd=0 as=0 ps=0 
M1142 diff_162000_2388000# diff_162000_2388000# diff_162000_2388000# GND efet w=3000 l=7800
+ ad=2.376e+08 pd=76800 as=0 ps=0 
M1143 Vdd Vdd diff_162000_2388000# GND efet w=9600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1144 diff_162000_2388000# diff_162000_2388000# diff_162000_2388000# GND efet w=1800 l=3600
+ ad=0 pd=0 as=0 ps=0 
M1145 Vdd Vdd Vdd GND efet w=2400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1146 Vdd Vdd Vdd GND efet w=1800 l=3600
+ ad=0 pd=0 as=0 ps=0 
M1147 Vdd diff_663600_2470800# diff_506400_2467200# GND efet w=13200 l=6600
+ ad=0 pd=0 as=0 ps=0 
M1148 diff_506400_2467200# diff_567600_2450400# GND GND efet w=52200 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1149 diff_951600_2584800# diff_940800_2611200# GND GND efet w=22800 l=9600
+ ad=2.376e+08 pd=74400 as=0 ps=0 
M1150 diff_904800_2581200# diff_894000_1458000# diff_663600_2611200# GND efet w=21600 l=7200
+ ad=2.6496e+08 pd=76800 as=0 ps=0 
M1151 GND diff_880800_2613600# diff_904800_2581200# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1152 diff_548400_2601600# diff_981600_1458000# diff_940800_2611200# GND efet w=10200 l=7200
+ ad=0 pd=0 as=2.6784e+08 ps=74400 
M1153 diff_1017600_2613600# diff_1009200_1458000# diff_548400_2601600# GND efet w=9600 l=7200
+ ad=2.592e+08 pd=76800 as=0 ps=0 
M1154 diff_663600_2611200# diff_945600_1442400# diff_951600_2584800# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1155 diff_904800_2547600# diff_894000_1458000# diff_664800_2534400# GND efet w=21600 l=7200
+ ad=2.6784e+08 pd=76800 as=0 ps=0 
M1156 diff_664800_2534400# diff_945600_1442400# diff_950400_2565600# GND efet w=21600 l=9000
+ ad=0 pd=0 as=2.4336e+08 ps=79200 
M1157 GND diff_880800_2528400# diff_904800_2547600# GND efet w=23400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1158 diff_548400_2534400# diff_843600_1497600# diff_804000_2528400# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6928e+08 ps=76800 
M1159 diff_880800_2528400# diff_872400_1458000# diff_548400_2534400# GND efet w=8400 l=7200
+ ad=2.448e+08 pd=74400 as=0 ps=0 
M1160 diff_567600_2450400# diff_663600_2470800# GND GND efet w=26400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1161 diff_567600_2410800# diff_423600_2420400# diff_548400_2392800# GND efet w=32400 l=7800
+ ad=9.6768e+08 pd=232800 as=-1.14281e+09 ps=866400 
M1162 diff_813600_2443200# diff_804000_2469600# GND GND efet w=22800 l=7200
+ ad=2.3184e+08 pd=72000 as=0 ps=0 
M1163 diff_548400_2460000# diff_843600_1497600# diff_804000_2469600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.5344e+08 ps=74400 
M1164 diff_880800_2472000# diff_872400_1458000# diff_548400_2460000# GND efet w=8400 l=7200
+ ad=2.5056e+08 pd=74400 as=0 ps=0 
M1165 diff_663600_2470800# diff_807600_1443600# diff_813600_2443200# GND efet w=21600 l=8400
+ ad=-2.09841e+09 pd=1.5432e+06 as=0 ps=0 
M1166 diff_664800_2392800# diff_807600_1443600# diff_813600_2401200# GND efet w=22200 l=7800
+ ad=2.01799e+09 pd=1.5528e+06 as=2.4336e+08 ps=76800 
M1167 GND diff_567600_2410800# diff_506400_2392800# GND efet w=50400 l=7200
+ ad=0 pd=0 as=1.68624e+09 ps=326400 
M1168 GND diff_664800_2392800# diff_567600_2410800# GND efet w=26400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1169 diff_69600_2534400# diff_68400_2361600# GND GND efet w=79200 l=6000
+ ad=-1.13129e+09 pd=609600 as=0 ps=0 
M1170 diff_487200_2368800# diff_326400_2457600# diff_231600_1357200# GND efet w=38400 l=7200
+ ad=9.6768e+08 pd=228000 as=-8.76219e+07 ps=2.7168e+06 
M1171 diff_487200_2368800# diff_523200_1467600# diff_506400_2392800# GND efet w=37800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1172 diff_548400_2392800# diff_426000_1591200# diff_487200_2368800# GND efet w=45600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1173 diff_506400_2392800# diff_664800_2392800# Vdd GND efet w=13800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1174 diff_813600_2401200# diff_804000_2386800# GND GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1175 diff_69600_2534400# diff_87600_2288400# GND GND efet w=216000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1176 Vdd diff_162000_2286000# diff_69600_2534400# GND efet w=11400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1177 diff_69600_2534400# diff_162000_2286000# diff_69600_2534400# GND efet w=40200 l=16800
+ ad=0 pd=0 as=0 ps=0 
M1178 diff_162000_2286000# diff_162000_2286000# diff_162000_2286000# GND efet w=2400 l=7200
+ ad=2.2464e+08 pd=76800 as=0 ps=0 
M1179 Vdd Vdd diff_162000_2286000# GND efet w=8400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1180 diff_487200_2312400# diff_327600_1404000# diff_349200_1096800# GND efet w=38400 l=7200
+ ad=1.10448e+09 pd=252000 as=0 ps=0 
M1181 diff_487200_2312400# diff_523200_1467600# diff_506400_2320800# GND efet w=39600 l=7200
+ ad=0 pd=0 as=1.6704e+09 ps=336000 
M1182 diff_567600_2410800# Vdd Vdd GND efet w=7200 l=27600
+ ad=0 pd=0 as=0 ps=0 
M1183 Vdd Vdd Vdd GND efet w=3600 l=10800
+ ad=0 pd=0 as=0 ps=0 
M1184 Vdd Vdd Vdd GND efet w=6000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M1185 diff_548400_2319600# diff_426000_1591200# diff_487200_2312400# GND efet w=45000 l=7800
+ ad=-1.18169e+09 pd=866400 as=0 ps=0 
M1186 diff_567600_2308800# Vdd Vdd GND efet w=7200 l=28800
+ ad=8.928e+08 pd=218400 as=0 ps=0 
M1187 Vdd diff_664800_2328000# diff_506400_2320800# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1188 diff_567600_2308800# diff_423600_2138400# diff_548400_2319600# GND efet w=32400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1189 diff_162000_2286000# diff_162000_2286000# diff_162000_2286000# GND efet w=3000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M1190 diff_487200_2258400# diff_327600_1404000# diff_252000_2766000# GND efet w=37200 l=7200
+ ad=9.5616e+08 pd=230400 as=0 ps=0 
M1191 diff_567600_2274000# diff_423600_2138400# diff_548400_2252400# GND efet w=31800 l=7800
+ ad=8.9136e+08 pd=216000 as=-1.18889e+09 ps=859200 
M1192 diff_506400_2320800# diff_567600_2308800# GND GND efet w=54600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1193 diff_950400_2565600# diff_940800_2528400# GND GND efet w=23400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1194 diff_904800_2439600# diff_894000_1458000# diff_663600_2470800# GND efet w=21600 l=7200
+ ad=2.6352e+08 pd=74400 as=0 ps=0 
M1195 GND diff_880800_2472000# diff_904800_2439600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1196 diff_950400_2443200# diff_940800_2470800# GND GND efet w=23400 l=7800
+ ad=2.592e+08 pd=74400 as=0 ps=0 
M1197 diff_1042800_2581200# diff_1032000_1458000# diff_663600_2611200# GND efet w=21600 l=7200
+ ad=2.3904e+08 pd=74400 as=0 ps=0 
M1198 GND diff_1017600_2613600# diff_1042800_2581200# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1199 diff_1088400_2584800# diff_1078800_2611200# GND GND efet w=22800 l=7200
+ ad=2.376e+08 pd=72000 as=0 ps=0 
M1200 diff_548400_2601600# diff_1118400_1497600# diff_1078800_2611200# GND efet w=9600 l=7200
+ ad=0 pd=0 as=2.6928e+08 ps=74400 
M1201 diff_1155600_2613600# diff_1147200_1458000# diff_548400_2601600# GND efet w=11400 l=6600
+ ad=2.5776e+08 pd=72000 as=0 ps=0 
M1202 diff_663600_2611200# diff_1082400_1443600# diff_1088400_2584800# GND efet w=21600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1203 diff_1042800_2546400# diff_1032000_1458000# diff_664800_2534400# GND efet w=21600 l=8400
+ ad=2.3904e+08 pd=74400 as=0 ps=0 
M1204 diff_664800_2534400# diff_1082400_1443600# diff_1088400_2542800# GND efet w=21600 l=9000
+ ad=0 pd=0 as=2.376e+08 ps=72000 
M1205 diff_548400_2534400# diff_981600_1458000# diff_940800_2528400# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.7216e+08 ps=76800 
M1206 diff_1017600_2528400# diff_1009200_1458000# diff_548400_2534400# GND efet w=8400 l=7200
+ ad=2.592e+08 pd=76800 as=0 ps=0 
M1207 diff_548400_2460000# diff_981600_1458000# diff_940800_2470800# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.5056e+08 ps=76800 
M1208 diff_1017600_2472000# diff_1009200_1458000# diff_548400_2460000# GND efet w=8400 l=7200
+ ad=2.5776e+08 pd=79200 as=0 ps=0 
M1209 diff_663600_2470800# diff_945600_1442400# diff_950400_2443200# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1210 diff_904800_2406000# diff_894000_1458000# diff_664800_2392800# GND efet w=21600 l=7200
+ ad=2.7072e+08 pd=76800 as=0 ps=0 
M1211 GND diff_880800_2386800# diff_904800_2406000# GND efet w=23400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1212 diff_548400_2392800# diff_843600_1497600# diff_804000_2386800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.7072e+08 ps=76800 
M1213 diff_880800_2386800# diff_872400_1458000# diff_548400_2392800# GND efet w=8400 l=7200
+ ad=2.5632e+08 pd=72000 as=0 ps=0 
M1214 diff_548400_2319600# diff_843600_1497600# diff_804000_2328000# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.7072e+08 ps=74400 
M1215 diff_880800_2330400# diff_872400_1458000# diff_548400_2319600# GND efet w=8400 l=7200
+ ad=2.592e+08 pd=72000 as=0 ps=0 
M1216 diff_567600_2308800# diff_664800_2328000# GND GND efet w=27000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1217 diff_813600_2301600# diff_804000_2328000# GND GND efet w=22800 l=7200
+ ad=2.3328e+08 pd=72000 as=0 ps=0 
M1218 GND diff_567600_2274000# diff_506400_2251200# GND efet w=50400 l=8400
+ ad=0 pd=0 as=1.6488e+09 ps=321600 
M1219 diff_664800_2328000# diff_807600_1443600# diff_813600_2301600# GND efet w=21600 l=8400
+ ad=-2.10993e+09 pd=1.5432e+06 as=0 ps=0 
M1220 diff_487200_2209200# diff_327600_1404000# diff_230400_2126400# GND efet w=37200 l=7200
+ ad=9.72e+08 pd=228000 as=0 ps=0 
M1221 diff_487200_2258400# diff_523200_1467600# diff_506400_2251200# GND efet w=37200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1222 diff_548400_2252400# diff_426000_1591200# diff_487200_2258400# GND efet w=46800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1223 GND diff_327600_1404000# diff_440400_2163600# GND efet w=56400 l=7200
+ ad=0 pd=0 as=5.2992e+08 ps=122400 
M1224 diff_487200_2209200# diff_523200_1467600# diff_506400_2186400# GND efet w=38400 l=7200
+ ad=0 pd=0 as=1.6776e+09 ps=328800 
M1225 diff_548400_2178000# diff_426000_1591200# diff_487200_2209200# GND efet w=45600 l=7200
+ ad=-1.15289e+09 pd=866400 as=0 ps=0 
M1226 GND diff_664800_2251200# diff_567600_2274000# GND efet w=26400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1227 diff_506400_2251200# diff_664800_2251200# Vdd GND efet w=13800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1228 diff_813600_2259600# diff_804000_2245200# GND GND efet w=24000 l=7200
+ ad=2.4192e+08 pd=74400 as=0 ps=0 
M1229 diff_664800_2251200# diff_807600_1443600# diff_813600_2259600# GND efet w=21600 l=8400
+ ad=1.84231e+09 pd=1.5288e+06 as=0 ps=0 
M1230 diff_567600_2274000# Vdd Vdd GND efet w=6000 l=26400
+ ad=0 pd=0 as=0 ps=0 
M1231 Vdd Vdd Vdd GND efet w=6000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M1232 Vdd Vdd Vdd GND efet w=3600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1233 diff_568800_2167200# Vdd Vdd GND efet w=6000 l=26400
+ ad=9.6912e+08 pd=232800 as=0 ps=0 
M1234 diff_568800_2167200# diff_423600_2138400# diff_548400_2178000# GND efet w=33600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1235 diff_440400_2163600# diff_426000_1591200# diff_423600_2138400# GND efet w=46800 l=8400
+ ad=0 pd=0 as=9.6192e+08 ps=204000 
M1236 GND diff_163200_2012400# diff_230400_2126400# GND efet w=38400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1237 d2 GND GND GND efet w=105600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1238 diff_230400_2126400# diff_170400_2043600# Vdd GND efet w=38400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1239 Vdd Vdd diff_423600_2138400# GND efet w=12000 l=38400
+ ad=0 pd=0 as=0 ps=0 
M1240 Vdd Vdd Vdd GND efet w=2400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1241 Vdd Vdd Vdd GND efet w=1800 l=3600
+ ad=0 pd=0 as=0 ps=0 
M1242 Vdd diff_664800_2186400# diff_506400_2186400# GND efet w=13800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1243 diff_506400_2186400# diff_568800_2167200# GND GND efet w=52800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1244 diff_950400_2408400# diff_940800_2386800# GND GND efet w=25800 l=9000
+ ad=2.5776e+08 pd=79200 as=0 ps=0 
M1245 diff_664800_2392800# diff_945600_1442400# diff_950400_2408400# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1246 diff_904800_2298000# diff_894000_1458000# diff_664800_2328000# GND efet w=21600 l=7200
+ ad=2.6496e+08 pd=76800 as=0 ps=0 
M1247 GND diff_880800_2330400# diff_904800_2298000# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1248 diff_951600_2301600# diff_940800_2329200# GND GND efet w=22800 l=8400
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1249 GND diff_1017600_2528400# diff_1042800_2546400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1250 diff_1088400_2542800# diff_1077600_2532000# GND GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1251 diff_1042800_2439600# diff_1032000_1458000# diff_663600_2470800# GND efet w=21600 l=7200
+ ad=2.376e+08 pd=72000 as=0 ps=0 
M1252 GND diff_1017600_2472000# diff_1042800_2439600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1253 diff_1088400_2443200# diff_1078800_2469600# GND GND efet w=22800 l=7200
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1254 diff_1179600_2581200# diff_1168800_1458000# diff_663600_2611200# GND efet w=21600 l=7200
+ ad=2.6496e+08 pd=74400 as=0 ps=0 
M1255 GND diff_1155600_2613600# diff_1179600_2581200# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1256 diff_1226400_2584800# diff_1215600_2611200# GND GND efet w=22800 l=8400
+ ad=2.376e+08 pd=74400 as=0 ps=0 
M1257 diff_548400_2601600# diff_1256400_1458000# diff_1215600_2611200# GND efet w=9600 l=7800
+ ad=0 pd=0 as=2.5776e+08 ps=76800 
M1258 diff_1292400_2613600# diff_1284000_1458000# diff_548400_2601600# GND efet w=9600 l=7200
+ ad=2.5344e+08 pd=74400 as=0 ps=0 
M1259 diff_663600_2611200# diff_1220400_1442400# diff_1226400_2584800# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1260 diff_1179600_2547600# diff_1168800_1458000# diff_664800_2534400# GND efet w=21600 l=7200
+ ad=2.6496e+08 pd=74400 as=0 ps=0 
M1261 diff_548400_2534400# diff_1118400_1497600# diff_1077600_2532000# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.664e+08 ps=74400 
M1262 diff_1155600_2528400# diff_1147200_1458000# diff_548400_2534400# GND efet w=9600 l=7200
+ ad=2.5344e+08 pd=72000 as=0 ps=0 
M1263 diff_548400_2460000# diff_1118400_1497600# diff_1078800_2469600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6784e+08 ps=74400 
M1264 diff_1155600_2472000# diff_1147200_1458000# diff_548400_2460000# GND efet w=9000 l=7200
+ ad=2.5056e+08 pd=74400 as=0 ps=0 
M1265 diff_663600_2470800# diff_1082400_1443600# diff_1088400_2443200# GND efet w=21600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1266 diff_1042800_2404800# diff_1032000_1458000# diff_664800_2392800# GND efet w=21600 l=7200
+ ad=2.4624e+08 pd=74400 as=0 ps=0 
M1267 diff_1017600_2386800# diff_1009200_1458000# diff_548400_2392800# GND efet w=8400 l=7800
+ ad=2.592e+08 pd=76800 as=0 ps=0 
M1268 diff_548400_2392800# diff_981600_1458000# diff_940800_2386800# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.664e+08 ps=76800 
M1269 diff_548400_2319600# diff_981600_1458000# diff_940800_2329200# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.6208e+08 ps=76800 
M1270 diff_1017600_2330400# diff_1009200_1458000# diff_548400_2319600# GND efet w=8400 l=7200
+ ad=2.6208e+08 pd=76800 as=0 ps=0 
M1271 diff_664800_2328000# diff_945600_1442400# diff_951600_2301600# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1272 diff_904800_2264400# diff_894000_1458000# diff_664800_2251200# GND efet w=20400 l=7200
+ ad=2.6496e+08 pd=74400 as=0 ps=0 
M1273 diff_664800_2251200# diff_945600_1442400# diff_951600_2259600# GND efet w=21000 l=9000
+ ad=0 pd=0 as=2.4048e+08 ps=74400 
M1274 GND diff_880800_2245200# diff_904800_2264400# GND efet w=23400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1275 diff_548400_2252400# diff_843600_1497600# diff_804000_2245200# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6352e+08 ps=74400 
M1276 diff_880800_2245200# diff_872400_1458000# diff_548400_2252400# GND efet w=8400 l=7200
+ ad=2.5776e+08 pd=74400 as=0 ps=0 
M1277 diff_548400_2178000# diff_843600_1497600# diff_804000_2187600# GND efet w=9600 l=7200
+ ad=0 pd=0 as=2.6064e+08 ps=74400 
M1278 diff_880800_2188800# diff_872400_1458000# diff_548400_2178000# GND efet w=9600 l=7200
+ ad=2.5632e+08 pd=72000 as=0 ps=0 
M1279 diff_951600_2259600# diff_940800_2246400# GND GND efet w=24000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1280 diff_568800_2167200# diff_664800_2186400# GND GND efet w=27000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1281 diff_568800_2127600# diff_423600_2138400# diff_548400_2109600# GND efet w=33600 l=8400
+ ad=9.36e+08 pd=232800 as=-1.15433e+09 ps=876000 
M1282 GND diff_568800_2127600# diff_506400_2109600# GND efet w=52200 l=7200
+ ad=0 pd=0 as=1.68624e+09 ps=324000 
M1283 diff_813600_2160000# diff_804000_2187600# GND GND efet w=24000 l=8400
+ ad=2.6064e+08 pd=74400 as=0 ps=0 
M1284 diff_664800_2186400# diff_807600_1443600# diff_813600_2160000# GND efet w=21000 l=7800
+ ad=2.07991e+09 pd=1.5408e+06 as=0 ps=0 
M1285 diff_487200_2085600# diff_327600_1404000# diff_231600_1357200# GND efet w=39000 l=7800
+ ad=9.9504e+08 pd=228000 as=0 ps=0 
M1286 diff_170400_2043600# diff_163200_2012400# GND GND efet w=21600 l=7200
+ ad=1.50624e+09 pd=276000 as=0 ps=0 
M1287 diff_170400_2043600# diff_170400_2043600# diff_170400_2043600# GND efet w=2400 l=3600
+ ad=0 pd=0 as=0 ps=0 
M1288 diff_170400_2043600# diff_170400_2043600# diff_170400_2043600# GND efet w=2400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1289 Vdd Vdd diff_170400_2043600# GND efet w=8400 l=37200
+ ad=0 pd=0 as=0 ps=0 
M1290 diff_487200_2085600# diff_523200_1467600# diff_506400_2109600# GND efet w=38400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1291 diff_548400_2109600# diff_426000_1591200# diff_487200_2085600# GND efet w=45000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1292 GND diff_664800_2109600# diff_568800_2127600# GND efet w=27600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1293 diff_813600_2119200# diff_804000_2103600# GND GND efet w=22800 l=7200
+ ad=2.6064e+08 pd=74400 as=0 ps=0 
M1294 diff_664800_2109600# diff_807600_1443600# diff_813600_2119200# GND efet w=21600 l=7200
+ ad=-2.14305e+09 pd=1.5504e+06 as=0 ps=0 
M1295 diff_506400_2109600# diff_664800_2109600# Vdd GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1296 diff_568800_2127600# Vdd Vdd GND efet w=6000 l=26400
+ ad=0 pd=0 as=0 ps=0 
M1297 diff_163200_2012400# diff_163200_2012400# diff_163200_2012400# GND efet w=2400 l=7200
+ ad=1.19808e+09 pd=280800 as=0 ps=0 
M1298 diff_163200_2012400# diff_163200_2012400# diff_163200_2012400# GND efet w=1800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1299 diff_163200_2012400# d2 GND GND efet w=56400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1300 diff_170400_2043600# diff_132000_2799600# GND GND efet w=34800 l=6600
+ ad=0 pd=0 as=0 ps=0 
M1301 diff_487200_2029200# diff_331200_1510800# diff_349200_1096800# GND efet w=38400 l=7200
+ ad=1.09728e+09 pd=247200 as=0 ps=0 
M1302 diff_487200_2029200# diff_523200_1467600# diff_506400_2037600# GND efet w=38400 l=7200
+ ad=0 pd=0 as=1.68192e+09 ps=326400 
M1303 Vdd Vdd Vdd GND efet w=6000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M1304 diff_548400_2036400# diff_426000_1591200# diff_487200_2029200# GND efet w=45000 l=7800
+ ad=-1.10969e+09 pd=864000 as=0 ps=0 
M1305 Vdd Vdd Vdd GND efet w=3600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1306 diff_568800_2025600# Vdd Vdd GND efet w=6600 l=27000
+ ad=8.7552e+08 pd=218400 as=0 ps=0 
M1307 Vdd diff_664800_2044800# diff_506400_2037600# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1308 diff_568800_2025600# diff_423600_1854000# diff_548400_2036400# GND efet w=31800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1309 GND diff_132000_2799600# diff_163200_2012400# GND efet w=34800 l=6600
+ ad=0 pd=0 as=0 ps=0 
M1310 GND GND GND GND efet w=600 l=1800
+ ad=0 pd=0 as=0 ps=0 
M1311 Vdd Vdd Vdd GND efet w=2400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1312 Vdd Vdd Vdd GND efet w=1800 l=4800
+ ad=0 pd=0 as=0 ps=0 
M1313 Vdd Vdd diff_163200_2012400# GND efet w=8400 l=36000
+ ad=0 pd=0 as=0 ps=0 
M1314 diff_487200_1975200# diff_331200_1510800# diff_252000_2766000# GND efet w=37200 l=7200
+ ad=9.7344e+08 pd=223200 as=0 ps=0 
M1315 diff_506400_2037600# diff_568800_2025600# GND GND efet w=52800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1316 diff_568800_2025600# diff_664800_2044800# GND GND efet w=28200 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1317 diff_813600_2018400# diff_804000_2044800# GND GND efet w=24600 l=7800
+ ad=2.6496e+08 pd=76800 as=0 ps=0 
M1318 diff_904800_2156400# diff_894000_1458000# diff_664800_2186400# GND efet w=22800 l=7800
+ ad=2.4336e+08 pd=76800 as=0 ps=0 
M1319 GND diff_880800_2188800# diff_904800_2156400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1320 diff_951600_2160000# diff_940800_2187600# GND GND efet w=22800 l=8400
+ ad=2.3472e+08 pd=74400 as=0 ps=0 
M1321 GND diff_1017600_2386800# diff_1042800_2404800# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1322 diff_1088400_2401200# diff_1078800_2386800# GND GND efet w=23400 l=7800
+ ad=2.4336e+08 pd=74400 as=0 ps=0 
M1323 diff_664800_2392800# diff_1082400_1443600# diff_1088400_2401200# GND efet w=23400 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1324 GND diff_1155600_2528400# diff_1179600_2547600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1325 diff_1226400_2542800# diff_1215600_2528400# GND GND efet w=22800 l=8400
+ ad=2.376e+08 pd=74400 as=0 ps=0 
M1326 diff_664800_2534400# diff_1220400_1442400# diff_1226400_2542800# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1327 diff_1179600_2439600# diff_1168800_1458000# diff_663600_2470800# GND efet w=21600 l=7200
+ ad=2.6208e+08 pd=74400 as=0 ps=0 
M1328 GND diff_1155600_2472000# diff_1179600_2439600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1329 diff_1226400_2443200# diff_1215600_2470800# GND GND efet w=22800 l=8400
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1330 diff_1317600_2581200# diff_1306800_1458000# diff_663600_2611200# GND efet w=21600 l=7200
+ ad=2.3904e+08 pd=74400 as=0 ps=0 
M1331 GND diff_1292400_2613600# diff_1317600_2581200# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1332 diff_1363200_2584800# diff_1353600_2611200# GND GND efet w=22800 l=7200
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1333 diff_548400_2601600# diff_1393200_1496400# diff_1353600_2611200# GND efet w=9600 l=7200
+ ad=0 pd=0 as=2.6928e+08 ps=74400 
M1334 diff_1430400_2613600# diff_1422000_1458000# diff_548400_2601600# GND efet w=9600 l=7800
+ ad=2.5776e+08 pd=72000 as=0 ps=0 
M1335 diff_663600_2611200# diff_1357200_1444800# diff_1363200_2584800# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1336 diff_1317600_2547600# diff_1306800_1458000# diff_664800_2534400# GND efet w=21000 l=7800
+ ad=2.376e+08 pd=74400 as=0 ps=0 
M1337 diff_548400_2534400# diff_1256400_1458000# diff_1215600_2528400# GND efet w=8400 l=9600
+ ad=0 pd=0 as=2.5056e+08 ps=74400 
M1338 diff_1292400_2528400# diff_1284000_1458000# diff_548400_2534400# GND efet w=8400 l=8400
+ ad=2.5488e+08 pd=76800 as=0 ps=0 
M1339 diff_548400_2460000# diff_1256400_1458000# diff_1215600_2470800# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.52e+08 ps=74400 
M1340 diff_1292400_2472000# diff_1284000_1458000# diff_548400_2460000# GND efet w=8400 l=7200
+ ad=2.5776e+08 pd=76800 as=0 ps=0 
M1341 diff_663600_2470800# diff_1220400_1442400# diff_1226400_2443200# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1342 diff_1179600_2406000# diff_1168800_1458000# diff_664800_2392800# GND efet w=21000 l=7200
+ ad=2.664e+08 pd=74400 as=0 ps=0 
M1343 diff_664800_2392800# diff_1220400_1442400# diff_1226400_2401200# GND efet w=21600 l=9600
+ ad=0 pd=0 as=2.3904e+08 ps=74400 
M1344 diff_548400_2392800# diff_1118400_1497600# diff_1078800_2386800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.664e+08 ps=74400 
M1345 diff_1155600_2386800# diff_1147200_1458000# diff_548400_2392800# GND efet w=9600 l=8400
+ ad=2.5632e+08 pd=72000 as=0 ps=0 
M1346 diff_1042800_2298000# diff_1032000_1458000# diff_664800_2328000# GND efet w=21600 l=7200
+ ad=2.3904e+08 pd=74400 as=0 ps=0 
M1347 GND diff_1017600_2330400# diff_1042800_2298000# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1348 diff_1088400_2300400# diff_1078800_2328000# GND GND efet w=22800 l=7200
+ ad=2.3904e+08 pd=74400 as=0 ps=0 
M1349 diff_548400_2319600# diff_1118400_1497600# diff_1078800_2328000# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6928e+08 ps=74400 
M1350 diff_1155600_2330400# diff_1147200_1458000# diff_548400_2319600# GND efet w=8400 l=8400
+ ad=2.592e+08 pd=72000 as=0 ps=0 
M1351 diff_664800_2328000# diff_1082400_1443600# diff_1088400_2300400# GND efet w=21600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1352 diff_1042800_2263200# diff_1032000_1458000# diff_664800_2251200# GND efet w=21600 l=9600
+ ad=2.4192e+08 pd=74400 as=0 ps=0 
M1353 diff_664800_2251200# diff_1082400_1443600# diff_1088400_2259600# GND efet w=21000 l=10200
+ ad=0 pd=0 as=2.4336e+08 ps=74400 
M1354 diff_548400_2252400# diff_981600_1458000# diff_940800_2246400# GND efet w=9600 l=8400
+ ad=0 pd=0 as=2.6928e+08 ps=81600 
M1355 diff_1017600_2245200# diff_1009200_1458000# diff_548400_2252400# GND efet w=8400 l=7200
+ ad=2.736e+08 pd=79200 as=0 ps=0 
M1356 diff_548400_2178000# diff_981600_1458000# diff_940800_2187600# GND efet w=10800 l=7800
+ ad=0 pd=0 as=2.664e+08 ps=81600 
M1357 diff_1017600_2188800# diff_1009200_1458000# diff_548400_2178000# GND efet w=9600 l=7200
+ ad=2.592e+08 pd=76800 as=0 ps=0 
M1358 diff_664800_2186400# diff_945600_1442400# diff_951600_2160000# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1359 diff_904800_2138400# diff_894000_1458000# diff_664800_2109600# GND efet w=24000 l=8400
+ ad=2.448e+08 pd=76800 as=0 ps=0 
M1360 GND diff_880800_2104800# diff_904800_2138400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1361 diff_951600_2119200# diff_940800_2103600# GND GND efet w=22800 l=8400
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1362 diff_664800_2109600# diff_945600_1442400# diff_951600_2119200# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1363 diff_548400_2109600# diff_843600_1497600# diff_804000_2103600# GND efet w=9600 l=7800
+ ad=0 pd=0 as=2.7072e+08 ps=74400 
M1364 diff_880800_2104800# diff_872400_1458000# diff_548400_2109600# GND efet w=8400 l=7200
+ ad=2.5488e+08 pd=72000 as=0 ps=0 
M1365 diff_548400_2036400# diff_843600_1497600# diff_804000_2044800# GND efet w=9000 l=9000
+ ad=0 pd=0 as=2.7072e+08 ps=76800 
M1366 diff_880800_2047200# diff_872400_1458000# diff_548400_2036400# GND efet w=9000 l=7800
+ ad=2.5776e+08 pd=72000 as=0 ps=0 
M1367 diff_568800_1984800# diff_423600_1854000# diff_548400_1968000# GND efet w=32400 l=9600
+ ad=8.8992e+08 pd=216000 as=-1.10393e+09 ps=907200 
M1368 GND diff_568800_1984800# diff_506400_1968000# GND efet w=51600 l=7200
+ ad=0 pd=0 as=1.63584e+09 ps=326400 
M1369 diff_664800_2044800# diff_807600_1443600# diff_813600_2018400# GND efet w=21600 l=7200
+ ad=2.13751e+09 pd=1.5408e+06 as=0 ps=0 
M1370 Vdd diff_68400_1594800# d3 GND efet w=612600 l=6600
+ ad=0 pd=0 as=1.51277e+09 ps=3.0288e+06 
M1371 GND diff_69600_1911600# d3 GND efet w=1146600 l=4200
+ ad=0 pd=0 as=0 ps=0 
M1372 diff_487200_1924800# diff_331200_1510800# diff_230400_2126400# GND efet w=38400 l=7200
+ ad=1.00368e+09 pd=232800 as=0 ps=0 
M1373 diff_487200_1975200# diff_523200_1467600# diff_506400_1968000# GND efet w=37200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1374 diff_548400_1968000# diff_426000_1591200# diff_487200_1975200# GND efet w=45000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1375 diff_487200_1924800# diff_523200_1467600# diff_506400_1902000# GND efet w=40800 l=7200
+ ad=0 pd=0 as=1.6704e+09 ps=328800 
M1376 GND diff_664800_1966800# diff_568800_1984800# GND efet w=26400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1377 diff_506400_1968000# diff_664800_1966800# Vdd GND efet w=14400 l=6600
+ ad=0 pd=0 as=0 ps=0 
M1378 diff_813600_1976400# diff_804000_1962000# GND GND efet w=24000 l=7200
+ ad=2.7072e+08 pd=76800 as=0 ps=0 
M1379 diff_664800_1966800# diff_807600_1443600# diff_813600_1976400# GND efet w=21600 l=7200
+ ad=1.87975e+09 pd=1.536e+06 as=0 ps=0 
M1380 Vdd Vdd Vdd GND efet w=6000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M1381 GND diff_331200_1510800# diff_440400_1879200# GND efet w=52800 l=6600
+ ad=0 pd=0 as=5.4576e+08 ps=124800 
M1382 diff_548400_1893600# diff_426000_1591200# diff_487200_1924800# GND efet w=46200 l=7800
+ ad=-1.12841e+09 pd=876000 as=0 ps=0 
M1383 diff_568800_1984800# Vdd Vdd GND efet w=7200 l=26400
+ ad=0 pd=0 as=0 ps=0 
M1384 Vdd Vdd Vdd GND efet w=3600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1385 diff_568800_1882800# Vdd Vdd GND efet w=7800 l=27000
+ ad=9.8352e+08 pd=232800 as=0 ps=0 
M1386 diff_568800_1882800# diff_423600_1854000# diff_548400_1893600# GND efet w=33000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1387 Vdd diff_664800_1902000# diff_506400_1902000# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1388 diff_440400_1879200# diff_426000_1591200# diff_423600_1854000# GND efet w=51000 l=7800
+ ad=0 pd=0 as=9.8496e+08 ps=211200 
M1389 Vdd Vdd diff_423600_1854000# GND efet w=11400 l=39000
+ ad=0 pd=0 as=0 ps=0 
M1390 Vdd Vdd Vdd GND efet w=2400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1391 Vdd Vdd Vdd GND efet w=2400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M1392 diff_506400_1902000# diff_568800_1882800# GND GND efet w=51600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1393 diff_568800_1882800# diff_664800_1902000# GND GND efet w=27000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1394 diff_813600_1876800# diff_804000_1903200# GND GND efet w=22800 l=7200
+ ad=2.6352e+08 pd=74400 as=0 ps=0 
M1395 diff_906000_2014800# diff_894000_1458000# diff_664800_2044800# GND efet w=21600 l=8400
+ ad=2.3904e+08 pd=74400 as=0 ps=0 
M1396 GND diff_880800_2047200# diff_906000_2014800# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1397 diff_951600_2018400# diff_940800_2044800# GND GND efet w=24600 l=7800
+ ad=2.376e+08 pd=74400 as=0 ps=0 
M1398 GND diff_1017600_2245200# diff_1042800_2263200# GND efet w=24600 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1399 diff_1088400_2259600# diff_1078800_2245200# GND GND efet w=24000 l=9600
+ ad=0 pd=0 as=0 ps=0 
M1400 diff_1042800_2156400# diff_1032000_1458000# diff_664800_2186400# GND efet w=21600 l=7200
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1401 GND diff_1017600_2188800# diff_1042800_2156400# GND efet w=23400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1402 diff_1088400_2160000# diff_1078800_2187600# GND GND efet w=22800 l=7200
+ ad=2.3328e+08 pd=72000 as=0 ps=0 
M1403 GND diff_1155600_2386800# diff_1179600_2406000# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1404 diff_1226400_2401200# diff_1215600_2386800# GND GND efet w=22800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1405 diff_1179600_2298000# diff_1168800_1458000# diff_664800_2328000# GND efet w=26400 l=7200
+ ad=2.592e+08 pd=84000 as=0 ps=0 
M1406 GND diff_1155600_2330400# diff_1179600_2298000# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1407 diff_1226400_2301600# diff_1215600_2329200# GND GND efet w=22800 l=8400
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1408 GND diff_1292400_2528400# diff_1317600_2547600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1409 diff_1363200_2542800# diff_1353600_2528400# GND GND efet w=22800 l=7200
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1410 diff_664800_2534400# diff_1357200_1444800# diff_1363200_2542800# GND efet w=21000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1411 diff_1317600_2439600# diff_1306800_1458000# diff_663600_2470800# GND efet w=21600 l=7200
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1412 GND diff_1292400_2472000# diff_1317600_2439600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1413 diff_1363200_2443200# diff_1353600_2469600# GND GND efet w=22800 l=7200
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1414 diff_1454400_2581200# diff_1443600_1458000# diff_663600_2611200# GND efet w=21600 l=7200
+ ad=2.6352e+08 pd=74400 as=0 ps=0 
M1415 GND diff_1430400_2613600# diff_1454400_2581200# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1416 diff_1501200_2584800# diff_1490400_2612400# GND GND efet w=22800 l=8400
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1417 diff_548400_2601600# diff_1531200_1458000# diff_1490400_2612400# GND efet w=10200 l=8400
+ ad=0 pd=0 as=2.5776e+08 ps=76800 
M1418 diff_1567200_2613600# diff_1558800_1458000# diff_548400_2601600# GND efet w=9000 l=7800
+ ad=2.6784e+08 pd=74400 as=0 ps=0 
M1419 diff_663600_2611200# diff_1495200_1443600# diff_1501200_2584800# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1420 diff_1454400_2547600# diff_1443600_1458000# diff_664800_2534400# GND efet w=21000 l=7800
+ ad=2.6208e+08 pd=74400 as=0 ps=0 
M1421 diff_548400_2534400# diff_1393200_1496400# diff_1353600_2528400# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6208e+08 ps=74400 
M1422 diff_1430400_2528400# diff_1422000_1458000# diff_548400_2534400# GND efet w=8400 l=8400
+ ad=2.5488e+08 pd=74400 as=0 ps=0 
M1423 diff_548400_2460000# diff_1393200_1496400# diff_1353600_2469600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6352e+08 ps=74400 
M1424 diff_1430400_2472000# diff_1422000_1458000# diff_548400_2460000# GND efet w=8400 l=8400
+ ad=2.5488e+08 pd=72000 as=0 ps=0 
M1425 diff_663600_2470800# diff_1357200_1444800# diff_1363200_2443200# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1426 diff_1317600_2406000# diff_1306800_1458000# diff_664800_2392800# GND efet w=21600 l=7200
+ ad=2.4336e+08 pd=74400 as=0 ps=0 
M1427 diff_548400_2392800# diff_1256400_1458000# diff_1215600_2386800# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.5632e+08 ps=76800 
M1428 diff_1292400_2386800# diff_1284000_1458000# diff_548400_2392800# GND efet w=8400 l=7200
+ ad=2.592e+08 pd=76800 as=0 ps=0 
M1429 diff_548400_2319600# diff_1256400_1458000# diff_1215600_2329200# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.6064e+08 ps=76800 
M1430 diff_1292400_2330400# diff_1284000_1458000# diff_548400_2319600# GND efet w=8400 l=7200
+ ad=2.5776e+08 pd=76800 as=0 ps=0 
M1431 diff_664800_2328000# diff_1220400_1442400# diff_1226400_2301600# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1432 diff_1179600_2268000# diff_1168800_1458000# diff_664800_2251200# GND efet w=22800 l=8400
+ ad=2.592e+08 pd=76800 as=0 ps=0 
M1433 GND diff_1155600_2245200# diff_1179600_2268000# GND efet w=23400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1434 diff_1226400_2259600# diff_1215600_2246400# GND GND efet w=24000 l=8400
+ ad=2.3472e+08 pd=74400 as=0 ps=0 
M1435 diff_664800_2251200# diff_1220400_1442400# diff_1226400_2259600# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1436 diff_548400_2252400# diff_1118400_1497600# diff_1078800_2245200# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.7072e+08 ps=76800 
M1437 diff_1155600_2245200# diff_1147200_1458000# diff_548400_2252400# GND efet w=9600 l=7800
+ ad=2.5488e+08 pd=72000 as=0 ps=0 
M1438 diff_548400_2178000# diff_1118400_1497600# diff_1078800_2187600# GND efet w=9600 l=7200
+ ad=0 pd=0 as=2.7504e+08 ps=76800 
M1439 diff_1155600_2188800# diff_1147200_1458000# diff_548400_2178000# GND efet w=9600 l=7200
+ ad=2.4336e+08 pd=69600 as=0 ps=0 
M1440 diff_664800_2186400# diff_1082400_1443600# diff_1088400_2160000# GND efet w=21600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1441 diff_1042800_2122800# diff_1032000_1458000# diff_664800_2109600# GND efet w=21600 l=7200
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1442 diff_548400_2109600# diff_981600_1458000# diff_940800_2103600# GND efet w=10200 l=7200
+ ad=0 pd=0 as=2.6928e+08 ps=81600 
M1443 diff_1017600_2103600# diff_1009200_1458000# diff_548400_2109600# GND efet w=8400 l=7200
+ ad=2.5632e+08 pd=76800 as=0 ps=0 
M1444 diff_548400_2036400# diff_981600_1458000# diff_940800_2044800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6784e+08 ps=74400 
M1445 diff_1017600_2048400# diff_1009200_1458000# diff_548400_2036400# GND efet w=8400 l=7200
+ ad=2.52e+08 pd=74400 as=0 ps=0 
M1446 diff_664800_2044800# diff_945600_1442400# diff_951600_2018400# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1447 diff_906000_1977600# diff_894000_1458000# diff_664800_1966800# GND efet w=22200 l=9000
+ ad=2.448e+08 pd=74400 as=0 ps=0 
M1448 diff_548400_1968000# diff_843600_1497600# diff_804000_1962000# GND efet w=12600 l=15600
+ ad=0 pd=0 as=2.6352e+08 ps=74400 
M1449 diff_880800_1962000# diff_872400_1458000# diff_548400_1968000# GND efet w=8400 l=7200
+ ad=2.6496e+08 pd=74400 as=0 ps=0 
M1450 diff_548400_1893600# diff_843600_1497600# diff_804000_1903200# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.6496e+08 ps=74400 
M1451 diff_880800_1904400# diff_872400_1458000# diff_548400_1893600# GND efet w=8400 l=7200
+ ad=2.5632e+08 pd=72000 as=0 ps=0 
M1452 diff_664800_1902000# diff_807600_1443600# diff_813600_1876800# GND efet w=20400 l=7200
+ ad=2.04823e+09 pd=1.5288e+06 as=0 ps=0 
M1453 diff_568800_1843200# diff_423600_1854000# diff_548400_1826400# GND efet w=31800 l=7200
+ ad=9.6912e+08 pd=232800 as=-1.17305e+09 ps=868800 
M1454 GND diff_568800_1843200# diff_506400_1825200# GND efet w=51600 l=8400
+ ad=0 pd=0 as=1.6848e+09 ps=324000 
M1455 GND diff_664800_1825200# diff_568800_1843200# GND efet w=27600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1456 diff_487200_1801200# diff_331200_1510800# diff_231600_1357200# GND efet w=39000 l=7800
+ ad=1.01088e+09 pd=230400 as=0 ps=0 
M1457 diff_487200_1801200# diff_523200_1467600# diff_506400_1825200# GND efet w=38400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1458 diff_548400_1826400# diff_426000_1591200# diff_487200_1801200# GND efet w=45000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1459 diff_506400_1825200# diff_664800_1825200# Vdd GND efet w=13800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1460 diff_813600_1834800# diff_804000_1819200# GND GND efet w=22800 l=7200
+ ad=2.6064e+08 pd=74400 as=0 ps=0 
M1461 diff_664800_1825200# diff_807600_1443600# diff_813600_1834800# GND efet w=21600 l=7200
+ ad=2.14615e+09 pd=1.5384e+06 as=0 ps=0 
M1462 diff_568800_1843200# Vdd Vdd GND efet w=6600 l=27600
+ ad=0 pd=0 as=0 ps=0 
M1463 diff_68400_1594800# diff_88800_1684800# GND GND efet w=218400 l=7200
+ ad=-2.75927e+08 pd=796800 as=0 ps=0 
M1464 diff_487200_1740000# diff_436800_1612800# diff_349200_1096800# GND efet w=37200 l=7200
+ ad=1.15344e+09 pd=259200 as=0 ps=0 
M1465 diff_487200_1740000# diff_523200_1467600# diff_506400_1747200# GND efet w=39600 l=7200
+ ad=0 pd=0 as=1.7064e+09 ps=336000 
M1466 Vdd Vdd Vdd GND efet w=6600 l=4200
+ ad=0 pd=0 as=0 ps=0 
M1467 diff_548400_1752000# diff_426000_1591200# diff_487200_1740000# GND efet w=45000 l=7800
+ ad=-1.13561e+09 pd=859200 as=0 ps=0 
M1468 Vdd Vdd Vdd GND efet w=3600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1469 diff_568800_1741200# Vdd Vdd GND efet w=6000 l=26400
+ ad=8.8272e+08 pd=216000 as=0 ps=0 
M1470 Vdd diff_664800_1760400# diff_506400_1747200# GND efet w=13800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1471 diff_88800_1684800# diff_88800_1684800# diff_88800_1684800# GND efet w=2400 l=4800
+ ad=1.1808e+09 pd=216000 as=0 ps=0 
M1472 diff_88800_1684800# diff_88800_1684800# diff_88800_1684800# GND efet w=3600 l=4800
+ ad=0 pd=0 as=0 ps=0 
M1473 diff_231600_1357200# diff_222000_1082400# diff_88800_1684800# GND efet w=27600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1474 diff_487200_1690800# diff_436800_1612800# diff_252000_2766000# GND efet w=37200 l=7200
+ ad=9.7056e+08 pd=228000 as=0 ps=0 
M1475 diff_568800_1741200# diff_423600_1570800# diff_548400_1752000# GND efet w=31200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1476 diff_568800_1701600# diff_423600_1570800# diff_548400_1684800# GND efet w=31800 l=7800
+ ad=8.7408e+08 pd=216000 as=-1.13417e+09 ps=866400 
M1477 diff_506400_1747200# diff_568800_1741200# GND GND efet w=50400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1478 diff_568800_1741200# diff_664800_1760400# GND GND efet w=26400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1479 GND diff_568800_1701600# diff_506400_1683600# GND efet w=51600 l=7200
+ ad=0 pd=0 as=1.6416e+09 ps=324000 
M1480 diff_813600_1734000# diff_804000_1760400# GND GND efet w=25800 l=7800
+ ad=2.6784e+08 pd=79200 as=0 ps=0 
M1481 GND diff_880800_1962000# diff_906000_1977600# GND efet w=23400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1482 diff_951600_1976400# diff_940800_1962000# GND GND efet w=26400 l=7200
+ ad=2.4336e+08 pd=74400 as=0 ps=0 
M1483 diff_664800_1966800# diff_945600_1442400# diff_951600_1976400# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1484 diff_906000_1872000# diff_894000_1458000# diff_664800_1902000# GND efet w=22200 l=9000
+ ad=2.4768e+08 pd=74400 as=0 ps=0 
M1485 GND diff_880800_1904400# diff_906000_1872000# GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1486 diff_951600_1875600# diff_940800_1903200# GND GND efet w=25800 l=7800
+ ad=2.4048e+08 pd=74400 as=0 ps=0 
M1487 GND diff_1017600_2103600# diff_1042800_2122800# GND efet w=22800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1488 diff_1088400_2119200# diff_1078800_2103600# GND GND efet w=22800 l=7200
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1489 diff_664800_2109600# diff_1082400_1443600# diff_1088400_2119200# GND efet w=21600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1490 diff_1180800_2156400# diff_1168800_1458000# diff_664800_2186400# GND efet w=21600 l=8400
+ ad=2.376e+08 pd=72000 as=0 ps=0 
M1491 GND diff_1155600_2188800# diff_1180800_2156400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1492 diff_1226400_2160000# diff_1215600_2187600# GND GND efet w=22800 l=8400
+ ad=2.3472e+08 pd=74400 as=0 ps=0 
M1493 diff_664800_2392800# diff_1357200_1444800# diff_1363200_2401200# GND efet w=21600 l=9600
+ ad=0 pd=0 as=2.3904e+08 ps=74400 
M1494 GND diff_1292400_2386800# diff_1317600_2406000# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1495 diff_1363200_2401200# diff_1353600_2386800# GND GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1496 diff_1317600_2298000# diff_1306800_1458000# diff_664800_2328000# GND efet w=21600 l=7200
+ ad=2.376e+08 pd=74400 as=0 ps=0 
M1497 GND diff_1292400_2330400# diff_1317600_2298000# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1498 diff_1363200_2301600# diff_1353600_2328000# GND GND efet w=22800 l=7200
+ ad=2.3328e+08 pd=72000 as=0 ps=0 
M1499 GND diff_1430400_2528400# diff_1454400_2547600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1500 diff_1501200_2542800# diff_1490400_2528400# GND GND efet w=22800 l=8400
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1501 diff_664800_2534400# diff_1495200_1443600# diff_1501200_2542800# GND efet w=21000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1502 diff_1454400_2439600# diff_1443600_1458000# diff_663600_2470800# GND efet w=21600 l=7200
+ ad=2.6064e+08 pd=74400 as=0 ps=0 
M1503 GND diff_1430400_2472000# diff_1454400_2439600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1504 diff_1501200_2443200# diff_1490400_2470800# GND GND efet w=22800 l=8400
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1505 diff_1592400_2581200# diff_1581600_1458000# diff_663600_2611200# GND efet w=21600 l=7200
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1506 GND diff_1567200_2613600# diff_1592400_2581200# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1507 diff_1638000_2584800# diff_1628400_2611200# GND GND efet w=22800 l=7200
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1508 diff_548400_2601600# diff_1668000_1497600# diff_1628400_2611200# GND efet w=9000 l=7800
+ ad=0 pd=0 as=2.5632e+08 ps=76800 
M1509 diff_1705200_2613600# diff_1696800_1458000# diff_548400_2601600# GND efet w=9000 l=7800
+ ad=2.5488e+08 pd=74400 as=0 ps=0 
M1510 diff_663600_2611200# diff_1633200_1442400# diff_1638000_2584800# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1511 diff_1592400_2547600# diff_1581600_1458000# diff_664800_2534400# GND efet w=21000 l=7800
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1512 diff_548400_2534400# diff_1531200_1458000# diff_1490400_2528400# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.52e+08 ps=72000 
M1513 diff_1567200_2528400# diff_1558800_1458000# diff_548400_2534400# GND efet w=8400 l=7200
+ ad=2.6496e+08 pd=74400 as=0 ps=0 
M1514 diff_548400_2460000# diff_1531200_1458000# diff_1490400_2470800# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.4768e+08 ps=76800 
M1515 diff_1567200_2472000# diff_1558800_1458000# diff_548400_2460000# GND efet w=8400 l=7200
+ ad=2.5344e+08 pd=74400 as=0 ps=0 
M1516 diff_663600_2470800# diff_1495200_1443600# diff_1501200_2443200# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1517 diff_1454400_2406000# diff_1443600_1458000# diff_664800_2392800# GND efet w=20400 l=7200
+ ad=2.6064e+08 pd=74400 as=0 ps=0 
M1518 diff_548400_2392800# diff_1393200_1496400# diff_1353600_2386800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6352e+08 ps=74400 
M1519 diff_1430400_2386800# diff_1422000_1458000# diff_548400_2392800# GND efet w=8400 l=8400
+ ad=2.5344e+08 pd=72000 as=0 ps=0 
M1520 diff_548400_2319600# diff_1393200_1496400# diff_1353600_2328000# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.664e+08 ps=74400 
M1521 diff_1430400_2330400# diff_1422000_1458000# diff_548400_2319600# GND efet w=8400 l=8400
+ ad=2.5488e+08 pd=74400 as=0 ps=0 
M1522 diff_664800_2328000# diff_1357200_1444800# diff_1363200_2301600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1523 diff_1317600_2264400# diff_1306800_1458000# diff_664800_2251200# GND efet w=20400 l=7200
+ ad=2.376e+08 pd=74400 as=0 ps=0 
M1524 diff_548400_2252400# diff_1256400_1458000# diff_1215600_2246400# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.5488e+08 ps=76800 
M1525 diff_1292400_2245200# diff_1284000_1458000# diff_548400_2252400# GND efet w=8400 l=7200
+ ad=2.5488e+08 pd=76800 as=0 ps=0 
M1526 diff_548400_2178000# diff_1256400_1458000# diff_1215600_2187600# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.5776e+08 ps=76800 
M1527 diff_1292400_2188800# diff_1284000_1458000# diff_548400_2178000# GND efet w=8400 l=7200
+ ad=2.6064e+08 pd=76800 as=0 ps=0 
M1528 diff_664800_2186400# diff_1220400_1442400# diff_1226400_2160000# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1529 diff_1180800_2120400# diff_1168800_1458000# diff_664800_2109600# GND efet w=21600 l=8400
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1530 diff_548400_2109600# diff_1118400_1497600# diff_1078800_2103600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6496e+08 ps=74400 
M1531 diff_1155600_2103600# diff_1147200_1458000# diff_548400_2109600# GND efet w=8400 l=7200
+ ad=2.5632e+08 pd=72000 as=0 ps=0 
M1532 diff_1042800_2014800# diff_1032000_1458000# diff_664800_2044800# GND efet w=21600 l=7200
+ ad=2.3904e+08 pd=74400 as=0 ps=0 
M1533 GND diff_1017600_2048400# diff_1042800_2014800# GND efet w=22800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1534 diff_1088400_2018400# diff_1078800_2044800# GND GND efet w=22800 l=7200
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1535 diff_548400_2036400# diff_1118400_1497600# diff_1078800_2044800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6784e+08 ps=74400 
M1536 diff_1155600_2048400# diff_1147200_1458000# diff_548400_2036400# GND efet w=8400 l=7200
+ ad=2.5632e+08 pd=72000 as=0 ps=0 
M1537 diff_664800_2044800# diff_1082400_1443600# diff_1088400_2018400# GND efet w=21600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1538 diff_1042800_1981200# diff_1032000_1458000# diff_664800_1966800# GND efet w=22200 l=7800
+ ad=2.4336e+08 pd=74400 as=0 ps=0 
M1539 diff_664800_1966800# diff_1082400_1443600# diff_1088400_1976400# GND efet w=22200 l=9000
+ ad=0 pd=0 as=2.448e+08 ps=76800 
M1540 GND diff_1017600_1962000# diff_1042800_1981200# GND efet w=23400 l=10200
+ ad=0 pd=0 as=0 ps=0 
M1541 diff_548400_1968000# diff_981600_1458000# diff_940800_1962000# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.808e+08 ps=79200 
M1542 diff_1017600_1962000# diff_1009200_1458000# diff_548400_1968000# GND efet w=8400 l=7200
+ ad=2.6208e+08 pd=79200 as=0 ps=0 
M1543 diff_548400_1893600# diff_981600_1458000# diff_940800_1903200# GND efet w=9000 l=7800
+ ad=0 pd=0 as=2.7072e+08 ps=81600 
M1544 diff_1017600_1905600# diff_1009200_1458000# diff_548400_1893600# GND efet w=8400 l=7200
+ ad=2.5488e+08 pd=76800 as=0 ps=0 
M1545 diff_664800_1902000# diff_945600_1442400# diff_951600_1875600# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1546 diff_906000_1836000# diff_894000_1458000# diff_664800_1825200# GND efet w=21600 l=8400
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1547 diff_548400_1826400# diff_843600_1497600# diff_804000_1819200# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.6928e+08 ps=76800 
M1548 diff_880800_1820400# diff_872400_1458000# diff_548400_1826400# GND efet w=8400 l=7200
+ ad=2.6064e+08 pd=74400 as=0 ps=0 
M1549 GND diff_880800_1820400# diff_906000_1836000# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1550 diff_951600_1834800# diff_940800_1819200# GND GND efet w=22800 l=7200
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1551 diff_664800_1825200# diff_945600_1442400# diff_951600_1834800# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1552 diff_548400_1752000# diff_843600_1497600# diff_804000_1760400# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.664e+08 ps=74400 
M1553 diff_880800_1762800# diff_872400_1458000# diff_548400_1752000# GND efet w=8400 l=7200
+ ad=2.5776e+08 pd=72000 as=0 ps=0 
M1554 diff_664800_1760400# diff_807600_1443600# diff_813600_1734000# GND efet w=21600 l=7200
+ ad=2.11015e+09 pd=1.5384e+06 as=0 ps=0 
M1555 diff_487200_1690800# diff_523200_1467600# diff_506400_1683600# GND efet w=39000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1556 diff_68400_1594800# diff_87600_2288400# GND GND efet w=218400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1557 Vdd diff_162000_1621200# diff_68400_1594800# GND efet w=10800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1558 diff_68400_1594800# diff_162000_1621200# diff_68400_1594800# GND efet w=49800 l=16800
+ ad=0 pd=0 as=0 ps=0 
M1559 diff_162000_1621200# diff_162000_1621200# diff_162000_1621200# GND efet w=2400 l=8400
+ ad=2.2896e+08 pd=81600 as=0 ps=0 
M1560 Vdd Vdd diff_162000_1621200# GND efet w=8400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1561 diff_162000_1621200# diff_162000_1621200# diff_162000_1621200# GND efet w=3600 l=4200
+ ad=0 pd=0 as=0 ps=0 
M1562 diff_69600_1911600# diff_68400_1594800# GND GND efet w=79200 l=6000
+ ad=-1.16873e+09 pd=607200 as=0 ps=0 
M1563 diff_69600_1911600# diff_87600_2288400# GND GND efet w=214800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1564 diff_69600_1911600# diff_162000_1520400# diff_69600_1911600# GND efet w=39000 l=18600
+ ad=0 pd=0 as=0 ps=0 
M1565 Vdd diff_162000_1520400# diff_69600_1911600# GND efet w=10800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1566 diff_162000_1520400# diff_162000_1520400# diff_162000_1520400# GND efet w=2400 l=9600
+ ad=2.1168e+08 pd=69600 as=0 ps=0 
M1567 Vdd Vdd diff_162000_1520400# GND efet w=8400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1568 diff_162000_1520400# diff_162000_1520400# diff_162000_1520400# GND efet w=600 l=3000
+ ad=0 pd=0 as=0 ps=0 
M1569 diff_487200_1641600# diff_436800_1612800# diff_230400_2126400# GND efet w=37200 l=7200
+ ad=9.4176e+08 pd=225600 as=0 ps=0 
M1570 diff_548400_1684800# diff_426000_1591200# diff_487200_1690800# GND efet w=45600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1571 GND diff_436800_1612800# diff_440400_1596000# GND efet w=52800 l=6600
+ ad=0 pd=0 as=5.5584e+08 ps=124800 
M1572 diff_487200_1641600# diff_523200_1467600# diff_506400_1618800# GND efet w=38400 l=8400
+ ad=0 pd=0 as=1.67328e+09 ps=326400 
M1573 diff_548400_1610400# diff_426000_1591200# diff_487200_1641600# GND efet w=45000 l=7800
+ ad=-1.21769e+09 pd=861600 as=0 ps=0 
M1574 GND diff_664800_1683600# diff_568800_1701600# GND efet w=28200 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1575 diff_506400_1683600# diff_664800_1683600# Vdd GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1576 diff_813600_1692000# diff_804000_1677600# GND GND efet w=25200 l=7200
+ ad=2.664e+08 pd=79200 as=0 ps=0 
M1577 diff_664800_1683600# diff_807600_1443600# diff_813600_1692000# GND efet w=21600 l=7200
+ ad=1.87255e+09 pd=1.5552e+06 as=0 ps=0 
M1578 diff_568800_1701600# Vdd Vdd GND efet w=6000 l=26400
+ ad=0 pd=0 as=0 ps=0 
M1579 Vdd Vdd Vdd GND efet w=6000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M1580 Vdd Vdd Vdd GND efet w=3600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1581 diff_568800_1599600# Vdd Vdd GND efet w=7200 l=27600
+ ad=9.2736e+08 pd=228000 as=0 ps=0 
M1582 diff_568800_1599600# diff_423600_1570800# diff_548400_1610400# GND efet w=34200 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1583 diff_440400_1596000# diff_426000_1591200# diff_423600_1570800# GND efet w=46800 l=7200
+ ad=0 pd=0 as=1.0008e+09 ps=204000 
M1584 Vdd Vdd diff_423600_1570800# GND efet w=12000 l=39600
+ ad=0 pd=0 as=0 ps=0 
M1585 Vdd Vdd Vdd GND efet w=1800 l=5400
+ ad=0 pd=0 as=0 ps=0 
M1586 Vdd Vdd Vdd GND efet w=1200 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1587 Vdd Vdd Vdd GND efet w=3000 l=4200
+ ad=0 pd=0 as=0 ps=0 
M1588 Vdd diff_664800_1620000# diff_506400_1618800# GND efet w=13800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1589 diff_506400_1618800# diff_568800_1599600# GND GND efet w=51600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1590 diff_568800_1599600# diff_664800_1620000# GND GND efet w=26400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1591 diff_568800_1560000# diff_423600_1570800# diff_548400_1543200# GND efet w=32400 l=7200
+ ad=9.648e+08 pd=230400 as=-1.15001e+09 ps=861600 
M1592 diff_813600_1597200# diff_804000_1620000# GND GND efet w=25200 l=7800
+ ad=2.3616e+08 pd=76800 as=0 ps=0 
M1593 GND diff_880800_1762800# diff_906000_1730400# GND efet w=23400 l=7800
+ ad=0 pd=0 as=2.376e+08 ps=74400 
M1594 diff_951600_1734000# diff_940800_1761600# GND GND efet w=25800 l=7800
+ ad=2.4336e+08 pd=74400 as=0 ps=0 
M1595 diff_906000_1730400# diff_894000_1458000# diff_664800_1760400# GND efet w=23400 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1596 diff_1088400_1976400# diff_1078800_1960800# GND GND efet w=22800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1597 GND diff_1155600_2103600# diff_1180800_2120400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1598 diff_1226400_2119200# diff_1215600_2103600# GND GND efet w=22800 l=7800
+ ad=2.3328e+08 pd=72000 as=0 ps=0 
M1599 diff_664800_2109600# diff_1220400_1442400# diff_1226400_2119200# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1600 diff_1180800_2014800# diff_1168800_1458000# diff_664800_2044800# GND efet w=21600 l=8400
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1601 GND diff_1155600_2048400# diff_1180800_2014800# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1602 diff_1226400_2018400# diff_1215600_2044800# GND GND efet w=25800 l=7800
+ ad=2.3616e+08 pd=74400 as=0 ps=0 
M1603 GND diff_1292400_2245200# diff_1317600_2264400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1604 diff_1363200_2259600# diff_1353600_2245200# GND GND efet w=22800 l=7200
+ ad=2.376e+08 pd=72000 as=0 ps=0 
M1605 diff_664800_2251200# diff_1357200_1444800# diff_1363200_2259600# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1606 GND diff_1430400_2386800# diff_1454400_2406000# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1607 diff_1500000_2420400# diff_1490400_2386800# GND GND efet w=24000 l=7800
+ ad=2.3328e+08 pd=76800 as=0 ps=0 
M1608 diff_664800_2392800# diff_1495200_1443600# diff_1500000_2420400# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1609 diff_1454400_2298000# diff_1443600_1458000# diff_664800_2328000# GND efet w=21600 l=7200
+ ad=2.592e+08 pd=74400 as=0 ps=0 
M1610 GND diff_1430400_2330400# diff_1454400_2298000# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1611 diff_1501200_2301600# diff_1490400_2329200# GND GND efet w=22800 l=8400
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1612 GND diff_1567200_2528400# diff_1592400_2547600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1613 diff_1638000_2542800# diff_1628400_2528400# GND GND efet w=22800 l=7200
+ ad=2.376e+08 pd=74400 as=0 ps=0 
M1614 diff_664800_2534400# diff_1633200_1442400# diff_1638000_2542800# GND efet w=21000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1615 diff_1592400_2439600# diff_1581600_1458000# diff_663600_2470800# GND efet w=21600 l=7200
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1616 GND diff_1567200_2472000# diff_1592400_2439600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1617 diff_1638000_2443200# diff_1628400_2470800# GND GND efet w=22800 l=7200
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1618 diff_1729200_2588400# diff_1719600_1458000# diff_663600_2611200# GND efet w=25800 l=7800
+ ad=2.4768e+08 pd=84000 as=0 ps=0 
M1619 GND diff_1705200_2613600# diff_1729200_2588400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1620 diff_1776000_2584800# diff_1765200_2612400# GND GND efet w=22800 l=7200
+ ad=2.376e+08 pd=74400 as=0 ps=0 
M1621 diff_548400_2601600# diff_1806000_1496400# diff_1765200_2612400# GND efet w=9600 l=7200
+ ad=0 pd=0 as=2.664e+08 ps=76800 
M1622 diff_1842000_2622000# diff_1834800_1458000# diff_548400_2601600# GND efet w=10200 l=7800
+ ad=2.592e+08 pd=79200 as=0 ps=0 
M1623 diff_663600_2611200# diff_1770000_1443600# diff_1776000_2584800# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1624 diff_1729200_2547600# diff_1719600_1458000# diff_664800_2534400# GND efet w=25200 l=7800
+ ad=2.5776e+08 pd=84000 as=0 ps=0 
M1625 diff_548400_2534400# diff_1668000_1497600# diff_1628400_2528400# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.5056e+08 ps=74400 
M1626 diff_1705200_2528400# diff_1696800_1458000# diff_548400_2534400# GND efet w=8400 l=7200
+ ad=2.5488e+08 pd=76800 as=0 ps=0 
M1627 diff_548400_2460000# diff_1668000_1497600# diff_1628400_2470800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.52e+08 ps=76800 
M1628 diff_1705200_2472000# diff_1696800_1458000# diff_548400_2460000# GND efet w=8400 l=7200
+ ad=2.5056e+08 pd=74400 as=0 ps=0 
M1629 diff_663600_2470800# diff_1633200_1442400# diff_1638000_2443200# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1630 diff_1592400_2406000# diff_1581600_1458000# diff_664800_2392800# GND efet w=20400 l=7800
+ ad=2.4048e+08 pd=74400 as=0 ps=0 
M1631 diff_548400_2392800# diff_1531200_1458000# diff_1490400_2386800# GND efet w=8400 l=7800
+ ad=0 pd=0 as=2.5488e+08 ps=72000 
M1632 diff_1567200_2386800# diff_1558800_1458000# diff_548400_2392800# GND efet w=8400 l=7200
+ ad=2.6496e+08 pd=74400 as=0 ps=0 
M1633 diff_548400_2319600# diff_1531200_1458000# diff_1490400_2329200# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.592e+08 ps=74400 
M1634 diff_1567200_2330400# diff_1558800_1458000# diff_548400_2319600# GND efet w=8400 l=7200
+ ad=2.6064e+08 pd=76800 as=0 ps=0 
M1635 diff_664800_2328000# diff_1495200_1443600# diff_1501200_2301600# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1636 diff_1454400_2264400# diff_1443600_1458000# diff_664800_2251200# GND efet w=20400 l=7200
+ ad=2.6208e+08 pd=74400 as=0 ps=0 
M1637 diff_548400_2252400# diff_1393200_1496400# diff_1353600_2245200# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6496e+08 ps=76800 
M1638 diff_1430400_2245200# diff_1422000_1458000# diff_548400_2252400# GND efet w=8400 l=8400
+ ad=2.52e+08 pd=72000 as=0 ps=0 
M1639 diff_1317600_2156400# diff_1306800_1458000# diff_664800_2186400# GND efet w=21600 l=7200
+ ad=2.3616e+08 pd=74400 as=0 ps=0 
M1640 GND diff_1292400_2188800# diff_1317600_2156400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1641 diff_1363200_2160000# diff_1353600_2187600# GND GND efet w=22800 l=7200
+ ad=2.3328e+08 pd=72000 as=0 ps=0 
M1642 diff_548400_2178000# diff_1393200_1496400# diff_1353600_2187600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.592e+08 ps=79200 
M1643 diff_1430400_2188800# diff_1422000_1458000# diff_548400_2178000# GND efet w=8400 l=8400
+ ad=2.5632e+08 pd=72000 as=0 ps=0 
M1644 diff_664800_2186400# diff_1357200_1444800# diff_1363200_2160000# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1645 diff_1317600_2122800# diff_1306800_1458000# diff_664800_2109600# GND efet w=21600 l=7200
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1646 diff_1292400_2104800# diff_1284000_1458000# diff_548400_2109600# GND efet w=10800 l=12600
+ ad=2.592e+08 pd=84000 as=0 ps=0 
M1647 diff_548400_2109600# diff_1256400_1458000# diff_1215600_2103600# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.592e+08 ps=76800 
M1648 diff_548400_2036400# diff_1256400_1458000# diff_1215600_2044800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.7072e+08 ps=79200 
M1649 diff_1292400_2047200# diff_1284000_1458000# diff_548400_2036400# GND efet w=8400 l=7200
+ ad=2.5776e+08 pd=74400 as=0 ps=0 
M1650 diff_664800_2044800# diff_1220400_1442400# diff_1226400_2018400# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1651 diff_1180800_1980000# diff_1168800_1458000# diff_664800_1966800# GND efet w=21600 l=9600
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1652 diff_664800_1966800# diff_1220400_1442400# diff_1226400_1976400# GND efet w=21000 l=9000
+ ad=0 pd=0 as=2.3616e+08 ps=74400 
M1653 diff_548400_1968000# diff_1118400_1497600# diff_1078800_1960800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.7648e+08 ps=76800 
M1654 diff_1155600_1962000# diff_1147200_1458000# diff_548400_1968000# GND efet w=8400 l=7200
+ ad=2.6496e+08 pd=74400 as=0 ps=0 
M1655 diff_1042800_1872000# diff_1032000_1458000# diff_664800_1902000# GND efet w=21600 l=7200
+ ad=2.4624e+08 pd=74400 as=0 ps=0 
M1656 GND diff_1017600_1905600# diff_1042800_1872000# GND efet w=24000 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1657 diff_1088400_1875600# diff_1078800_1903200# GND GND efet w=24000 l=7200
+ ad=2.4624e+08 pd=76800 as=0 ps=0 
M1658 diff_548400_1893600# diff_1118400_1497600# diff_1078800_1903200# GND efet w=9000 l=7200
+ ad=0 pd=0 as=2.6928e+08 ps=76800 
M1659 diff_1155600_1904400# diff_1147200_1458000# diff_548400_1893600# GND efet w=8400 l=7200
+ ad=2.5632e+08 pd=72000 as=0 ps=0 
M1660 diff_664800_1902000# diff_1082400_1443600# diff_1088400_1875600# GND efet w=22800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1661 diff_1042800_1838400# diff_1032000_1458000# diff_664800_1825200# GND efet w=21600 l=7200
+ ad=2.376e+08 pd=72000 as=0 ps=0 
M1662 diff_548400_1826400# diff_981600_1458000# diff_940800_1819200# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6928e+08 ps=81600 
M1663 diff_1017600_1820400# diff_1009200_1458000# diff_548400_1826400# GND efet w=8400 l=7200
+ ad=2.5632e+08 pd=79200 as=0 ps=0 
M1664 diff_548400_1752000# diff_981600_1458000# diff_940800_1761600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.7072e+08 ps=79200 
M1665 diff_1017600_1764000# diff_1009200_1458000# diff_548400_1752000# GND efet w=8400 l=7200
+ ad=2.6496e+08 pd=74400 as=0 ps=0 
M1666 diff_664800_1760400# diff_945600_1442400# diff_951600_1734000# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1667 diff_906000_1693200# diff_894000_1458000# diff_664800_1683600# GND efet w=22800 l=10200
+ ad=2.4192e+08 pd=72000 as=0 ps=0 
M1668 diff_548400_1684800# diff_843600_1497600# diff_804000_1677600# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.6496e+08 ps=74400 
M1669 diff_880800_1677600# diff_872400_1458000# diff_548400_1684800# GND efet w=8400 l=7200
+ ad=2.5488e+08 pd=72000 as=0 ps=0 
M1670 GND diff_880800_1677600# diff_906000_1693200# GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1671 diff_951600_1692000# diff_940800_1677600# GND GND efet w=25800 l=7800
+ ad=2.4336e+08 pd=74400 as=0 ps=0 
M1672 diff_664800_1683600# diff_945600_1442400# diff_951600_1692000# GND efet w=22200 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1673 diff_548400_1610400# diff_843600_1497600# diff_804000_1620000# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.6496e+08 ps=74400 
M1674 diff_880800_1621200# diff_872400_1458000# diff_548400_1610400# GND efet w=8400 l=7200
+ ad=2.5776e+08 pd=72000 as=0 ps=0 
M1675 diff_664800_1620000# diff_807600_1443600# diff_813600_1597200# GND efet w=21600 l=7200
+ ad=1.92151e+09 pd=1.5288e+06 as=0 ps=0 
M1676 GND diff_568800_1560000# diff_506400_1542000# GND efet w=51600 l=7200
+ ad=0 pd=0 as=1.71792e+09 ps=326400 
M1677 diff_487200_1521600# diff_436800_1612800# diff_231600_1357200# GND efet w=40200 l=9000
+ ad=9.288e+08 pd=228000 as=0 ps=0 
M1678 diff_487200_1521600# diff_523200_1467600# diff_506400_1542000# GND efet w=37200 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1679 diff_548400_1543200# diff_426000_1591200# diff_487200_1521600# GND efet w=45000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1680 GND diff_664800_1543200# diff_568800_1560000# GND efet w=26400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1681 diff_506400_1542000# diff_664800_1543200# Vdd GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1682 diff_814800_1551600# diff_804000_1537200# GND GND efet w=22800 l=8400
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1683 diff_664800_1543200# diff_807600_1443600# diff_814800_1551600# GND efet w=21600 l=7200
+ ad=1.99207e+09 pd=1.5432e+06 as=0 ps=0 
M1684 diff_568800_1560000# Vdd Vdd GND efet w=6600 l=27000
+ ad=0 pd=0 as=0 ps=0 
M1685 Vdd Vdd Vdd GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M1686 Vdd Vdd Vdd GND efet w=1800 l=6600
+ ad=0 pd=0 as=0 ps=0 
M1687 diff_906000_1588800# diff_894000_1458000# diff_664800_1620000# GND efet w=21600 l=8400
+ ad=2.376e+08 pd=72000 as=0 ps=0 
M1688 GND diff_880800_1621200# diff_906000_1588800# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1689 diff_951600_1592400# diff_940800_1620000# GND GND efet w=25800 l=7800
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1690 GND diff_1017600_1820400# diff_1042800_1838400# GND efet w=22800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1691 diff_1088400_1834800# diff_1078800_1819200# GND GND efet w=22800 l=7200
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1692 diff_664800_1825200# diff_1082400_1443600# diff_1088400_1834800# GND efet w=21600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1693 GND diff_1155600_1962000# diff_1180800_1980000# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1694 diff_1226400_1976400# diff_1215600_1962000# GND GND efet w=25200 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1695 GND diff_1292400_2104800# diff_1317600_2122800# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1696 diff_1363200_2119200# diff_1353600_2103600# GND GND efet w=22800 l=7200
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1697 diff_664800_2109600# diff_1357200_1444800# diff_1363200_2119200# GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1698 GND diff_1430400_2245200# diff_1454400_2264400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1699 diff_1501200_2259600# diff_1490400_2246400# GND GND efet w=22800 l=8400
+ ad=2.3328e+08 pd=74400 as=0 ps=0 
M1700 diff_664800_2251200# diff_1495200_1443600# diff_1501200_2259600# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1701 diff_1454400_2156400# diff_1443600_1458000# diff_664800_2186400# GND efet w=21600 l=7200
+ ad=2.6064e+08 pd=74400 as=0 ps=0 
M1702 GND diff_1430400_2188800# diff_1454400_2156400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1703 diff_1501200_2160000# diff_1490400_2187600# GND GND efet w=22800 l=8400
+ ad=2.3472e+08 pd=74400 as=0 ps=0 
M1704 GND diff_1567200_2386800# diff_1592400_2406000# GND efet w=22800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1705 diff_1638000_2401200# diff_1628400_2386800# GND GND efet w=22800 l=7200
+ ad=2.3616e+08 pd=74400 as=0 ps=0 
M1706 diff_664800_2392800# diff_1633200_1442400# diff_1638000_2401200# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1707 diff_1592400_2298000# diff_1581600_1458000# diff_664800_2328000# GND efet w=21600 l=7200
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1708 GND diff_1567200_2330400# diff_1592400_2298000# GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1709 diff_1638000_2301600# diff_1628400_2328000# GND GND efet w=22800 l=7200
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1710 GND diff_1705200_2528400# diff_1729200_2547600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1711 diff_1776000_2542800# diff_1765200_2529600# GND GND efet w=22800 l=7200
+ ad=2.376e+08 pd=74400 as=0 ps=0 
M1712 diff_664800_2534400# diff_1770000_1443600# diff_1776000_2542800# GND efet w=21000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1713 diff_1729200_2439600# diff_1719600_1458000# diff_663600_2470800# GND efet w=21600 l=7200
+ ad=2.6208e+08 pd=74400 as=0 ps=0 
M1714 GND diff_1705200_2472000# diff_1729200_2439600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1715 diff_1776000_2443200# diff_1765200_2470800# GND GND efet w=22800 l=7200
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1716 diff_1867200_2581200# diff_1856400_1458000# diff_663600_2611200# GND efet w=21600 l=7200
+ ad=2.6208e+08 pd=76800 as=0 ps=0 
M1717 GND diff_1842000_2622000# diff_1867200_2581200# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1718 diff_1914000_2584800# diff_1903200_2612400# GND GND efet w=22800 l=7200
+ ad=2.376e+08 pd=74400 as=0 ps=0 
M1719 diff_548400_2601600# diff_1944000_1496400# diff_1903200_2612400# GND efet w=7800 l=7800
+ ad=0 pd=0 as=2.6496e+08 ps=74400 
M1720 diff_1980000_2614800# diff_1972800_1458000# diff_548400_2601600# GND efet w=8400 l=7200
+ ad=2.6208e+08 pd=79200 as=0 ps=0 
M1721 diff_663600_2611200# diff_1908000_1442400# diff_1914000_2584800# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1722 diff_1867200_2547600# diff_1856400_1458000# diff_664800_2534400# GND efet w=20400 l=7200
+ ad=2.664e+08 pd=76800 as=0 ps=0 
M1723 diff_548400_2534400# diff_1806000_1496400# diff_1765200_2529600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6496e+08 ps=74400 
M1724 diff_1843200_2528400# diff_1834800_1458000# diff_548400_2534400# GND efet w=8400 l=8400
+ ad=2.5488e+08 pd=76800 as=0 ps=0 
M1725 diff_548400_2460000# diff_1806000_1496400# diff_1765200_2470800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6496e+08 ps=74400 
M1726 diff_1842000_2472000# diff_1834800_1458000# diff_548400_2460000# GND efet w=9000 l=7800
+ ad=2.5344e+08 pd=84000 as=0 ps=0 
M1727 diff_663600_2470800# diff_1770000_1443600# diff_1776000_2443200# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1728 diff_1729200_2407200# diff_1719600_1458000# diff_664800_2392800# GND efet w=20400 l=7200
+ ad=2.6064e+08 pd=76800 as=0 ps=0 
M1729 diff_664800_2392800# diff_1770000_1443600# diff_1776000_2401200# GND efet w=21600 l=8400
+ ad=0 pd=0 as=2.3904e+08 ps=74400 
M1730 diff_548400_2392800# diff_1668000_1497600# diff_1628400_2386800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.5344e+08 ps=76800 
M1731 diff_1705200_2386800# diff_1696800_1458000# diff_548400_2392800# GND efet w=8400 l=7200
+ ad=2.592e+08 pd=76800 as=0 ps=0 
M1732 diff_548400_2319600# diff_1668000_1497600# diff_1628400_2328000# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.4048e+08 ps=74400 
M1733 diff_1705200_2330400# diff_1696800_1458000# diff_548400_2319600# GND efet w=8400 l=7200
+ ad=2.3904e+08 pd=72000 as=0 ps=0 
M1734 diff_664800_2328000# diff_1633200_1442400# diff_1638000_2301600# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1735 diff_1592400_2264400# diff_1581600_1458000# diff_664800_2251200# GND efet w=20400 l=7200
+ ad=2.3616e+08 pd=74400 as=0 ps=0 
M1736 diff_548400_2252400# diff_1531200_1458000# diff_1490400_2246400# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.5056e+08 ps=74400 
M1737 diff_1567200_2245200# diff_1558800_1458000# diff_548400_2252400# GND efet w=8400 l=7200
+ ad=2.6064e+08 pd=74400 as=0 ps=0 
M1738 diff_548400_2178000# diff_1531200_1458000# diff_1490400_2187600# GND efet w=9600 l=7200
+ ad=0 pd=0 as=2.4912e+08 ps=74400 
M1739 diff_1567200_2188800# diff_1558800_1458000# diff_548400_2178000# GND efet w=8400 l=7200
+ ad=2.6496e+08 pd=74400 as=0 ps=0 
M1740 diff_664800_2186400# diff_1495200_1443600# diff_1501200_2160000# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1741 diff_1454400_2124000# diff_1443600_1458000# diff_664800_2109600# GND efet w=21600 l=7200
+ ad=2.592e+08 pd=74400 as=0 ps=0 
M1742 diff_548400_2109600# diff_1393200_1496400# diff_1353600_2103600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6352e+08 ps=74400 
M1743 diff_1430400_2104800# diff_1422000_1458000# diff_548400_2109600# GND efet w=9600 l=7200
+ ad=2.6208e+08 pd=74400 as=0 ps=0 
M1744 diff_1317600_2014800# diff_1306800_1458000# diff_664800_2044800# GND efet w=21600 l=7200
+ ad=2.3904e+08 pd=74400 as=0 ps=0 
M1745 GND diff_1292400_2047200# diff_1317600_2014800# GND efet w=27000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1746 diff_1363200_2018400# diff_1353600_2044800# GND GND efet w=22800 l=7200
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1747 diff_548400_2036400# diff_1393200_1496400# diff_1353600_2044800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.664e+08 ps=74400 
M1748 diff_1430400_2048400# diff_1422000_1458000# diff_548400_2036400# GND efet w=8400 l=7200
+ ad=2.592e+08 pd=74400 as=0 ps=0 
M1749 diff_664800_2044800# diff_1357200_1444800# diff_1363200_2018400# GND efet w=21600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1750 diff_1317600_1981200# diff_1306800_1458000# diff_664800_1966800# GND efet w=21600 l=7800
+ ad=2.3904e+08 pd=74400 as=0 ps=0 
M1751 GND diff_1292400_1962000# diff_1317600_1981200# GND efet w=27000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1752 diff_548400_1968000# diff_1256400_1458000# diff_1215600_1962000# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6352e+08 ps=76800 
M1753 diff_1292400_1962000# diff_1284000_1458000# diff_548400_1968000# GND efet w=8400 l=7200
+ ad=2.6928e+08 pd=76800 as=0 ps=0 
M1754 diff_1180800_1872000# diff_1168800_1458000# diff_664800_1902000# GND efet w=21600 l=8400
+ ad=2.448e+08 pd=74400 as=0 ps=0 
M1755 GND diff_1155600_1904400# diff_1180800_1872000# GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1756 diff_1226400_1875600# diff_1215600_1903200# GND GND efet w=24600 l=7800
+ ad=2.4048e+08 pd=74400 as=0 ps=0 
M1757 diff_548400_1893600# diff_1256400_1458000# diff_1215600_1903200# GND efet w=9600 l=7200
+ ad=0 pd=0 as=2.736e+08 ps=79200 
M1758 diff_1292400_1904400# diff_1284000_1458000# diff_548400_1893600# GND efet w=9600 l=7200
+ ad=2.7504e+08 pd=79200 as=0 ps=0 
M1759 diff_664800_1902000# diff_1220400_1442400# diff_1226400_1875600# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1760 diff_1180800_1837200# diff_1168800_1458000# diff_664800_1825200# GND efet w=22200 l=9000
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1761 diff_548400_1826400# diff_1118400_1497600# diff_1078800_1819200# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.664e+08 ps=74400 
M1762 diff_1155600_1819200# diff_1147200_1458000# diff_548400_1826400# GND efet w=8400 l=7200
+ ad=2.6064e+08 pd=74400 as=0 ps=0 
M1763 diff_1042800_1730400# diff_1032000_1458000# diff_664800_1760400# GND efet w=21600 l=7200
+ ad=2.3904e+08 pd=74400 as=0 ps=0 
M1764 GND diff_1017600_1764000# diff_1042800_1730400# GND efet w=22800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1765 diff_1088400_1734000# diff_1078800_1761600# GND GND efet w=22800 l=7200
+ ad=2.4048e+08 pd=74400 as=0 ps=0 
M1766 diff_548400_1752000# diff_1118400_1497600# diff_1078800_1761600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6784e+08 ps=74400 
M1767 diff_1155600_1762800# diff_1147200_1458000# diff_548400_1752000# GND efet w=8400 l=7200
+ ad=2.5488e+08 pd=74400 as=0 ps=0 
M1768 diff_664800_1760400# diff_1082400_1443600# diff_1088400_1734000# GND efet w=22800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1769 diff_1042800_1696800# diff_1032000_1458000# diff_664800_1683600# GND efet w=21600 l=7800
+ ad=2.448e+08 pd=74400 as=0 ps=0 
M1770 diff_548400_1684800# diff_981600_1458000# diff_940800_1677600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6208e+08 ps=76800 
M1771 diff_1017600_1677600# diff_1009200_1458000# diff_548400_1684800# GND efet w=9000 l=7200
+ ad=2.6352e+08 pd=74400 as=0 ps=0 
M1772 diff_548400_1610400# diff_981600_1458000# diff_940800_1620000# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6928e+08 ps=79200 
M1773 diff_1018800_1621200# diff_1009200_1458000# diff_548400_1610400# GND efet w=8400 l=8400
+ ad=2.5776e+08 pd=76800 as=0 ps=0 
M1774 diff_664800_1620000# diff_945600_1442400# diff_951600_1592400# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1775 diff_906000_1551600# diff_894000_1458000# diff_664800_1543200# GND efet w=24000 l=8400
+ ad=2.448e+08 pd=74400 as=0 ps=0 
M1776 diff_548400_1543200# diff_843600_1497600# diff_804000_1537200# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.6496e+08 ps=74400 
M1777 diff_880800_1536000# diff_872400_1458000# diff_548400_1543200# GND efet w=9000 l=7800
+ ad=2.5632e+08 pd=72000 as=0 ps=0 
M1778 GND diff_880800_1536000# diff_906000_1551600# GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1779 diff_951600_1550400# diff_940800_1537200# GND GND efet w=24600 l=7800
+ ad=2.4192e+08 pd=74400 as=0 ps=0 
M1780 diff_664800_1543200# diff_945600_1442400# diff_951600_1550400# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1781 GND diff_1017600_1677600# diff_1042800_1696800# GND efet w=24000 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1782 diff_1088400_1692000# diff_1078800_1677600# GND GND efet w=24000 l=7200
+ ad=2.448e+08 pd=74400 as=0 ps=0 
M1783 diff_664800_1683600# diff_1082400_1443600# diff_1088400_1692000# GND efet w=22200 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1784 GND diff_1155600_1819200# diff_1180800_1837200# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1785 diff_1226400_1834800# diff_1215600_1819200# GND GND efet w=24600 l=7800
+ ad=2.3328e+08 pd=72000 as=0 ps=0 
M1786 diff_664800_1825200# diff_1220400_1442400# diff_1226400_1834800# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1787 diff_1180800_1730400# diff_1168800_1458000# diff_664800_1760400# GND efet w=21600 l=8400
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1788 GND diff_1155600_1762800# diff_1180800_1730400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1789 diff_1226400_1734000# diff_1215600_1761600# GND GND efet w=27000 l=7800
+ ad=2.376e+08 pd=74400 as=0 ps=0 
M1790 diff_1363200_1976400# diff_1353600_1962000# GND GND efet w=22800 l=7200
+ ad=2.4048e+08 pd=72000 as=0 ps=0 
M1791 diff_664800_1966800# diff_1357200_1444800# diff_1363200_1976400# GND efet w=21600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1792 GND diff_1430400_2104800# diff_1454400_2124000# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1793 diff_1501200_2119200# diff_1490400_2103600# GND GND efet w=22800 l=7800
+ ad=2.3328e+08 pd=72000 as=0 ps=0 
M1794 diff_664800_2109600# diff_1495200_1443600# diff_1501200_2119200# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1795 diff_1454400_2014800# diff_1443600_1458000# diff_664800_2044800# GND efet w=21600 l=7200
+ ad=2.6064e+08 pd=74400 as=0 ps=0 
M1796 GND diff_1430400_2048400# diff_1454400_2014800# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1797 diff_1501200_2018400# diff_1490400_2044800# GND GND efet w=24000 l=7800
+ ad=2.3328e+08 pd=72000 as=0 ps=0 
M1798 GND diff_1567200_2245200# diff_1592400_2264400# GND efet w=25800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1799 diff_1638000_2259600# diff_1628400_2245200# GND GND efet w=22800 l=7200
+ ad=2.376e+08 pd=74400 as=0 ps=0 
M1800 diff_664800_2251200# diff_1633200_1442400# diff_1638000_2259600# GND efet w=21000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1801 GND diff_1705200_2386800# diff_1729200_2407200# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1802 diff_1776000_2401200# diff_1765200_2388000# GND GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1803 diff_1729200_2298000# diff_1719600_1458000# diff_664800_2328000# GND efet w=22800 l=7200
+ ad=2.5776e+08 pd=76800 as=0 ps=0 
M1804 GND diff_1705200_2330400# diff_1729200_2298000# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1805 diff_1776000_2301600# diff_1765200_2329200# GND GND efet w=22800 l=7200
+ ad=2.376e+08 pd=72000 as=0 ps=0 
M1806 GND diff_1843200_2528400# diff_1867200_2547600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1807 diff_1914000_2542800# diff_1903200_2529600# GND GND efet w=22800 l=7200
+ ad=2.4048e+08 pd=74400 as=0 ps=0 
M1808 diff_664800_2534400# diff_1908000_1442400# diff_1914000_2542800# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1809 diff_1867200_2439600# diff_1856400_1458000# diff_663600_2470800# GND efet w=21600 l=7200
+ ad=2.6352e+08 pd=76800 as=0 ps=0 
M1810 GND diff_1842000_2472000# diff_1867200_2439600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1811 diff_1914000_2443200# diff_1903200_2470800# GND GND efet w=23400 l=7800
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1812 diff_2005200_2581200# diff_1994400_1460400# diff_663600_2611200# GND efet w=21600 l=7200
+ ad=2.6064e+08 pd=76800 as=0 ps=0 
M1813 GND diff_1980000_2614800# diff_2005200_2581200# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1814 diff_2052000_2584800# diff_2041200_2612400# GND GND efet w=25200 l=7200
+ ad=2.3184e+08 pd=72000 as=0 ps=0 
M1815 diff_548400_2601600# diff_2082000_1496400# diff_2041200_2612400# GND efet w=7200 l=7200
+ ad=0 pd=0 as=2.5776e+08 ps=74400 
M1816 diff_2118000_2614800# diff_2110800_1458000# diff_548400_2601600# GND efet w=7200 l=7200
+ ad=2.5488e+08 pd=76800 as=0 ps=0 
M1817 diff_663600_2611200# diff_2046000_1444800# diff_2052000_2584800# GND efet w=21000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1818 diff_2005200_2548800# diff_1994400_1460400# diff_664800_2534400# GND efet w=20400 l=7200
+ ad=2.6064e+08 pd=76800 as=0 ps=0 
M1819 diff_548400_2534400# diff_1944000_1496400# diff_1903200_2529600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6064e+08 ps=74400 
M1820 diff_1980000_2528400# diff_1972800_1458000# diff_548400_2534400# GND efet w=8400 l=7200
+ ad=2.5776e+08 pd=76800 as=0 ps=0 
M1821 diff_548400_2460000# diff_1944000_1496400# diff_1903200_2470800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.5776e+08 ps=79200 
M1822 diff_1980000_2472000# diff_1972800_1458000# diff_548400_2460000# GND efet w=8400 l=7200
+ ad=2.592e+08 pd=76800 as=0 ps=0 
M1823 diff_663600_2470800# diff_1908000_1442400# diff_1914000_2443200# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1824 diff_664800_2392800# diff_1908000_1442400# diff_1914000_2401200# GND efet w=21600 l=8400
+ ad=0 pd=0 as=2.3472e+08 ps=74400 
M1825 diff_1867200_2407200# diff_1856400_1458000# diff_664800_2392800# GND efet w=20400 l=7200
+ ad=2.5776e+08 pd=76800 as=0 ps=0 
M1826 GND diff_1842000_2389200# diff_1867200_2407200# GND efet w=23400 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1827 diff_548400_2392800# diff_1806000_1496400# diff_1765200_2388000# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.7504e+08 ps=76800 
M1828 diff_1842000_2389200# diff_1834800_1458000# diff_548400_2392800# GND efet w=10800 l=7800
+ ad=2.5776e+08 pd=81600 as=0 ps=0 
M1829 diff_548400_2319600# diff_1806000_1496400# diff_1765200_2329200# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.5488e+08 ps=76800 
M1830 diff_1842000_2334000# diff_1834800_1458000# diff_548400_2319600# GND efet w=9600 l=7200
+ ad=2.5344e+08 pd=76800 as=0 ps=0 
M1831 diff_664800_2328000# diff_1770000_1443600# diff_1776000_2301600# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1832 diff_1729200_2264400# diff_1719600_1458000# diff_664800_2251200# GND efet w=21600 l=7200
+ ad=2.52e+08 pd=79200 as=0 ps=0 
M1833 diff_548400_2252400# diff_1668000_1497600# diff_1628400_2245200# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.5344e+08 ps=76800 
M1834 diff_1705200_2245200# diff_1696800_1458000# diff_548400_2252400# GND efet w=8400 l=7200
+ ad=2.6496e+08 pd=76800 as=0 ps=0 
M1835 diff_548400_2178000# diff_1668000_1497600# diff_1628400_2187600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.5056e+08 ps=74400 
M1836 diff_1705200_2188800# diff_1696800_1458000# diff_548400_2178000# GND efet w=8400 l=7200
+ ad=2.5344e+08 pd=74400 as=0 ps=0 
M1837 diff_1592400_2156400# diff_1581600_1458000# diff_664800_2186400# GND efet w=21600 l=7200
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1838 GND diff_1567200_2188800# diff_1592400_2156400# GND efet w=24600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1839 diff_1638000_2160000# diff_1628400_2187600# GND GND efet w=22800 l=7200
+ ad=2.3616e+08 pd=74400 as=0 ps=0 
M1840 diff_664800_2186400# diff_1633200_1442400# diff_1638000_2160000# GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1841 diff_1592400_2122800# diff_1581600_1458000# diff_664800_2109600# GND efet w=21600 l=7200
+ ad=2.376e+08 pd=72000 as=0 ps=0 
M1842 diff_664800_2109600# diff_1633200_1442400# diff_1638000_2119200# GND efet w=24000 l=7200
+ ad=0 pd=0 as=2.4768e+08 ps=76800 
M1843 diff_548400_2109600# diff_1531200_1458000# diff_1490400_2103600# GND efet w=7200 l=7200
+ ad=0 pd=0 as=2.6928e+08 ps=76800 
M1844 diff_1567200_2103600# diff_1558800_1458000# diff_548400_2109600# GND efet w=7200 l=7200
+ ad=2.664e+08 pd=74400 as=0 ps=0 
M1845 diff_548400_2036400# diff_1531200_1458000# diff_1490400_2044800# GND efet w=9600 l=7200
+ ad=0 pd=0 as=2.6784e+08 ps=74400 
M1846 diff_1567200_2047200# diff_1558800_1458000# diff_548400_2036400# GND efet w=8400 l=7200
+ ad=2.664e+08 pd=74400 as=0 ps=0 
M1847 diff_664800_2044800# diff_1495200_1443600# diff_1501200_2018400# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1848 diff_1454400_1981200# diff_1443600_1458000# diff_664800_1966800# GND efet w=21000 l=7800
+ ad=2.6208e+08 pd=74400 as=0 ps=0 
M1849 diff_548400_1968000# diff_1393200_1496400# diff_1353600_1962000# GND efet w=9600 l=7200
+ ad=0 pd=0 as=2.736e+08 ps=79200 
M1850 diff_1430400_1960800# diff_1422000_1458000# diff_548400_1968000# GND efet w=8400 l=7200
+ ad=2.736e+08 pd=76800 as=0 ps=0 
M1851 diff_1317600_1872000# diff_1306800_1458000# diff_664800_1902000# GND efet w=21600 l=7200
+ ad=2.232e+08 pd=74400 as=0 ps=0 
M1852 GND diff_1292400_1904400# diff_1317600_1872000# GND efet w=24600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1853 diff_1363200_1875600# diff_1353600_1903200# GND GND efet w=24000 l=7200
+ ad=2.4624e+08 pd=74400 as=0 ps=0 
M1854 diff_548400_1893600# diff_1393200_1496400# diff_1353600_1903200# GND efet w=9600 l=7200
+ ad=0 pd=0 as=2.6784e+08 ps=74400 
M1855 diff_1430400_1904400# diff_1422000_1458000# diff_548400_1893600# GND efet w=9600 l=7200
+ ad=2.6064e+08 pd=76800 as=0 ps=0 
M1856 diff_664800_1902000# diff_1357200_1444800# diff_1363200_1875600# GND efet w=21600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1857 diff_1317600_1838400# diff_1306800_1458000# diff_664800_1825200# GND efet w=21600 l=7200
+ ad=2.376e+08 pd=72000 as=0 ps=0 
M1858 diff_548400_1826400# diff_1256400_1458000# diff_1215600_1819200# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.664e+08 ps=79200 
M1859 diff_1292400_1820400# diff_1284000_1458000# diff_548400_1826400# GND efet w=8400 l=7200
+ ad=2.5632e+08 pd=74400 as=0 ps=0 
M1860 diff_548400_1752000# diff_1256400_1458000# diff_1215600_1761600# GND efet w=9000 l=7200
+ ad=0 pd=0 as=2.6064e+08 ps=79200 
M1861 diff_1292400_1764000# diff_1284000_1458000# diff_548400_1752000# GND efet w=8400 l=7200
+ ad=2.4048e+08 pd=74400 as=0 ps=0 
M1862 diff_664800_1760400# diff_1220400_1442400# diff_1226400_1734000# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1863 diff_1180800_1694400# diff_1168800_1458000# diff_664800_1683600# GND efet w=21600 l=9600
+ ad=2.3904e+08 pd=72000 as=0 ps=0 
M1864 GND diff_1155600_1677600# diff_1180800_1694400# GND efet w=23400 l=9000
+ ad=0 pd=0 as=0 ps=0 
M1865 diff_548400_1684800# diff_1118400_1497600# diff_1078800_1677600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6496e+08 ps=74400 
M1866 diff_1155600_1677600# diff_1147200_1458000# diff_548400_1684800# GND efet w=8400 l=7200
+ ad=2.6064e+08 pd=74400 as=0 ps=0 
M1867 diff_1042800_1588800# diff_1032000_1458000# diff_664800_1620000# GND efet w=21600 l=7200
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1868 GND diff_1018800_1621200# diff_1042800_1588800# GND efet w=22800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1869 diff_1088400_1592400# diff_1078800_1620000# GND GND efet w=22800 l=7200
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1870 diff_548400_1610400# diff_1118400_1497600# diff_1078800_1620000# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.664e+08 ps=74400 
M1871 diff_1155600_1621200# diff_1147200_1458000# diff_548400_1610400# GND efet w=8400 l=7200
+ ad=2.5488e+08 pd=72000 as=0 ps=0 
M1872 diff_664800_1620000# diff_1082400_1443600# diff_1088400_1592400# GND efet w=21600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1873 diff_1042800_1555200# diff_1032000_1458000# diff_664800_1543200# GND efet w=21600 l=7200
+ ad=2.4336e+08 pd=74400 as=0 ps=0 
M1874 diff_548400_1543200# diff_981600_1458000# diff_940800_1537200# GND efet w=9600 l=8400
+ ad=0 pd=0 as=2.7072e+08 ps=79200 
M1875 diff_1018800_1528800# diff_1009200_1458000# diff_548400_1543200# GND efet w=9000 l=9000
+ ad=2.5776e+08 pd=74400 as=0 ps=0 
M1876 GND diff_1018800_1528800# diff_1042800_1555200# GND efet w=24000 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1877 diff_1088400_1550400# diff_1078800_1537200# GND GND efet w=24000 l=7200
+ ad=2.4912e+08 pd=79200 as=0 ps=0 
M1878 diff_664800_1543200# diff_1082400_1443600# diff_1088400_1550400# GND efet w=24000 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1879 diff_1226400_1692000# diff_1215600_1677600# GND GND efet w=24000 l=9600
+ ad=2.4048e+08 pd=74400 as=0 ps=0 
M1880 diff_664800_1683600# diff_1220400_1442400# diff_1226400_1692000# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1881 diff_1180800_1588800# diff_1168800_1458000# diff_664800_1620000# GND efet w=21600 l=8400
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1882 GND diff_1155600_1621200# diff_1180800_1588800# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1883 diff_1226400_1592400# diff_1215600_1620000# GND GND efet w=22800 l=7800
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1884 GND diff_1292400_1820400# diff_1317600_1838400# GND efet w=23400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1885 diff_1363200_1834800# diff_1353600_1819200# GND GND efet w=22800 l=7200
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1886 diff_664800_1825200# diff_1357200_1444800# diff_1363200_1834800# GND efet w=21600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1887 GND diff_1430400_1960800# diff_1454400_1981200# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1888 diff_1501200_1976400# diff_1490400_1962000# GND GND efet w=22800 l=7800
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1889 diff_664800_1966800# diff_1495200_1443600# diff_1501200_1976400# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1890 diff_1454400_1872000# diff_1443600_1458000# diff_664800_1902000# GND efet w=21600 l=7200
+ ad=2.7216e+08 pd=76800 as=0 ps=0 
M1891 GND diff_1430400_1904400# diff_1454400_1872000# GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1892 diff_1501200_1875600# diff_1490400_1903200# GND GND efet w=24600 l=7800
+ ad=2.4192e+08 pd=74400 as=0 ps=0 
M1893 GND diff_1567200_2103600# diff_1592400_2122800# GND efet w=22800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1894 diff_1638000_2119200# diff_1628400_2103600# GND GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1895 GND diff_1567200_2047200# diff_1592400_2014800# GND efet w=24000 l=7800
+ ad=0 pd=0 as=2.376e+08 ps=74400 
M1896 diff_1592400_2014800# diff_1581600_1458000# diff_664800_2044800# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1897 diff_1638000_2018400# diff_1628400_2044800# GND GND efet w=22800 l=7200
+ ad=2.6352e+08 pd=76800 as=0 ps=0 
M1898 GND diff_1705200_2245200# diff_1729200_2264400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1899 diff_1776000_2259600# diff_1765200_2246400# GND GND efet w=22800 l=7200
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1900 diff_664800_2251200# diff_1770000_1443600# diff_1776000_2259600# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1901 diff_1729200_2158800# diff_1719600_1458000# diff_664800_2186400# GND efet w=22800 l=7800
+ ad=2.4048e+08 pd=76800 as=0 ps=0 
M1902 GND diff_1705200_2188800# diff_1729200_2158800# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1903 diff_1776000_2160000# diff_1765200_2188800# GND GND efet w=22800 l=7200
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1904 diff_1914000_2401200# diff_1903200_2386800# GND GND efet w=24000 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1905 diff_1867200_2298000# diff_1856400_1458000# diff_664800_2328000# GND efet w=21600 l=7200
+ ad=2.6352e+08 pd=76800 as=0 ps=0 
M1906 GND diff_1842000_2334000# diff_1867200_2298000# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1907 diff_1914000_2301600# diff_1903200_2329200# GND GND efet w=24000 l=7200
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1908 GND diff_1980000_2528400# diff_2005200_2548800# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1909 diff_2052000_2542800# diff_2041200_2528400# GND GND efet w=24600 l=7800
+ ad=2.3904e+08 pd=74400 as=0 ps=0 
M1910 diff_664800_2534400# diff_2046000_1444800# diff_2052000_2542800# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1911 diff_2005200_2439600# diff_1994400_1460400# diff_663600_2470800# GND efet w=21600 l=7200
+ ad=2.6064e+08 pd=76800 as=0 ps=0 
M1912 GND diff_1980000_2472000# diff_2005200_2439600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1913 diff_2050800_2456400# diff_2041200_2470800# GND GND efet w=25200 l=7800
+ ad=2.3472e+08 pd=76800 as=0 ps=0 
M1914 Vdd diff_1892400_663600# diff_548400_2601600# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1915 diff_2143200_2581200# diff_2133600_1458000# diff_663600_2611200# GND efet w=21600 l=7200
+ ad=2.6928e+08 pd=76800 as=0 ps=0 
M1916 GND diff_2118000_2614800# diff_2143200_2581200# GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1917 Vdd diff_2224800_1584000# diff_663600_2611200# GND efet w=14400 l=6600
+ ad=0 pd=0 as=0 ps=0 
M1918 diff_2415600_2852400# Vdd Vdd GND efet w=10800 l=19200
+ ad=0 pd=0 as=0 ps=0 
M1919 Vdd Vdd Vdd GND efet w=5400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M1920 Vdd Vdd Vdd GND efet w=4200 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1921 diff_2414400_2601600# Vdd Vdd GND efet w=13200 l=18600
+ ad=1.25424e+09 pd=261600 as=0 ps=0 
M1922 diff_2325600_2576400# clk2 diff_230400_2126400# GND efet w=19200 l=7200
+ ad=2.736e+08 pd=76800 as=0 ps=0 
M1923 diff_2344800_2570400# diff_2074800_2772000# diff_2325600_2576400# GND efet w=19200 l=7200
+ ad=1.67184e+09 pd=326400 as=0 ps=0 
M1924 diff_2143200_2548800# diff_2133600_1458000# diff_664800_2534400# GND efet w=20400 l=7200
+ ad=2.1024e+08 pd=64800 as=0 ps=0 
M1925 GND diff_2118000_2528400# diff_2143200_2548800# GND efet w=16800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1926 diff_548400_2534400# diff_2082000_1496400# diff_2041200_2528400# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.5776e+08 ps=74400 
M1927 diff_2118000_2528400# diff_2110800_1458000# diff_548400_2534400# GND efet w=8400 l=7200
+ ad=2.5776e+08 pd=76800 as=0 ps=0 
M1928 diff_548400_2460000# diff_2082000_1496400# diff_2041200_2470800# GND efet w=7800 l=9000
+ ad=0 pd=0 as=2.4192e+08 ps=86400 
M1929 diff_2118000_2472000# diff_2110800_1458000# diff_548400_2460000# GND efet w=8400 l=8400
+ ad=2.5344e+08 pd=74400 as=0 ps=0 
M1930 diff_663600_2470800# diff_2046000_1444800# diff_2050800_2456400# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1931 diff_2005200_2407200# diff_1994400_1460400# diff_664800_2392800# GND efet w=21000 l=7800
+ ad=2.52e+08 pd=76800 as=0 ps=0 
M1932 diff_548400_2392800# diff_1944000_1496400# diff_1903200_2386800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6352e+08 ps=74400 
M1933 diff_1980000_2386800# diff_1972800_1458000# diff_548400_2392800# GND efet w=8400 l=7200
+ ad=2.6208e+08 pd=76800 as=0 ps=0 
M1934 diff_548400_2319600# diff_1944000_1496400# diff_1903200_2329200# GND efet w=9000 l=7800
+ ad=0 pd=0 as=2.6784e+08 ps=74400 
M1935 diff_1980000_2330400# diff_1972800_1458000# diff_548400_2319600# GND efet w=8400 l=7200
+ ad=2.6208e+08 pd=76800 as=0 ps=0 
M1936 diff_664800_2328000# diff_1908000_1442400# diff_1914000_2301600# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1937 diff_1867200_2265600# diff_1856400_1458000# diff_664800_2251200# GND efet w=20400 l=7200
+ ad=2.592e+08 pd=74400 as=0 ps=0 
M1938 diff_548400_2252400# diff_1806000_1496400# diff_1765200_2246400# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6208e+08 ps=76800 
M1939 diff_1842000_2251200# diff_1834800_1458000# diff_548400_2252400# GND efet w=10200 l=7200
+ ad=2.5776e+08 pd=79200 as=0 ps=0 
M1940 diff_548400_2178000# diff_1806000_1496400# diff_1765200_2188800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6496e+08 ps=74400 
M1941 diff_1843200_2188800# diff_1834800_1458000# diff_548400_2178000# GND efet w=8400 l=8400
+ ad=2.5632e+08 pd=76800 as=0 ps=0 
M1942 diff_664800_2186400# diff_1770000_1443600# diff_1776000_2160000# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1943 diff_1730400_2122800# diff_1719600_1458000# diff_664800_2109600# GND efet w=21600 l=8400
+ ad=2.4336e+08 pd=74400 as=0 ps=0 
M1944 diff_548400_2109600# diff_1668000_1497600# diff_1628400_2103600# GND efet w=7800 l=7800
+ ad=0 pd=0 as=2.5344e+08 ps=74400 
M1945 diff_1705200_2103600# diff_1696800_1458000# diff_548400_2109600# GND efet w=8400 l=8400
+ ad=2.5488e+08 pd=74400 as=0 ps=0 
M1946 GND diff_1705200_2103600# diff_1730400_2122800# GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1947 diff_1776000_2118000# diff_1765200_2109600# GND GND efet w=24000 l=7200
+ ad=2.4048e+08 pd=74400 as=0 ps=0 
M1948 diff_664800_2109600# diff_1770000_1443600# diff_1776000_2118000# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1949 diff_1705200_2047200# diff_1696800_1458000# diff_548400_2036400# GND efet w=9600 l=8400
+ ad=2.52e+08 pd=74400 as=0 ps=0 
M1950 diff_548400_2036400# diff_1668000_1497600# diff_1628400_2044800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.5344e+08 ps=74400 
M1951 diff_664800_2044800# diff_1633200_1442400# diff_1638000_2018400# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1952 diff_1592400_1981200# diff_1581600_1458000# diff_664800_1966800# GND efet w=20400 l=7200
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1953 diff_548400_1968000# diff_1531200_1458000# diff_1490400_1962000# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.592e+08 ps=74400 
M1954 diff_1567200_1962000# diff_1558800_1458000# diff_548400_1968000# GND efet w=8400 l=7200
+ ad=2.6064e+08 pd=79200 as=0 ps=0 
M1955 diff_548400_1893600# diff_1531200_1458000# diff_1490400_1903200# GND efet w=9000 l=7800
+ ad=0 pd=0 as=2.6784e+08 ps=74400 
M1956 diff_1567200_1904400# diff_1558800_1458000# diff_548400_1893600# GND efet w=9600 l=7200
+ ad=2.7072e+08 pd=79200 as=0 ps=0 
M1957 diff_664800_1902000# diff_1495200_1443600# diff_1501200_1875600# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1958 diff_1454400_1839600# diff_1443600_1458000# diff_664800_1825200# GND efet w=21600 l=7200
+ ad=2.6208e+08 pd=74400 as=0 ps=0 
M1959 diff_548400_1826400# diff_1393200_1496400# diff_1353600_1819200# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6496e+08 ps=74400 
M1960 diff_1430400_1819200# diff_1422000_1458000# diff_548400_1826400# GND efet w=8400 l=7200
+ ad=2.6208e+08 pd=74400 as=0 ps=0 
M1961 GND diff_1292400_1764000# diff_1317600_1730400# GND efet w=25800 l=7800
+ ad=0 pd=0 as=2.3904e+08 ps=74400 
M1962 diff_1317600_1730400# diff_1306800_1458000# diff_664800_1760400# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1963 diff_1363200_1734000# diff_1353600_1760400# GND GND efet w=22800 l=7200
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M1964 diff_548400_1752000# diff_1393200_1496400# diff_1353600_1760400# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6352e+08 ps=74400 
M1965 diff_1430400_1764000# diff_1422000_1458000# diff_548400_1752000# GND efet w=8400 l=7200
+ ad=2.5056e+08 pd=74400 as=0 ps=0 
M1966 diff_664800_1760400# diff_1357200_1444800# diff_1363200_1734000# GND efet w=21600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1967 diff_1317600_1696800# diff_1306800_1458000# diff_664800_1683600# GND efet w=20400 l=7200
+ ad=2.3904e+08 pd=74400 as=0 ps=0 
M1968 diff_548400_1684800# diff_1256400_1458000# diff_1215600_1677600# GND efet w=9600 l=8400
+ ad=0 pd=0 as=2.592e+08 ps=79200 
M1969 diff_1292400_1677600# diff_1284000_1458000# diff_548400_1684800# GND efet w=8400 l=7200
+ ad=2.6064e+08 pd=76800 as=0 ps=0 
M1970 diff_548400_1610400# diff_1256400_1458000# diff_1215600_1620000# GND efet w=10200 l=7800
+ ad=0 pd=0 as=2.592e+08 ps=84000 
M1971 diff_1292400_1621200# diff_1284000_1458000# diff_548400_1610400# GND efet w=8400 l=7200
+ ad=2.52e+08 pd=79200 as=0 ps=0 
M1972 diff_664800_1620000# diff_1220400_1442400# diff_1226400_1592400# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1973 diff_1180800_1554000# diff_1168800_1458000# diff_664800_1543200# GND efet w=21600 l=8400
+ ad=2.4192e+08 pd=74400 as=0 ps=0 
M1974 diff_548400_1543200# diff_1118400_1497600# diff_1078800_1537200# GND efet w=9000 l=7800
+ ad=0 pd=0 as=2.6928e+08 ps=74400 
M1975 diff_1155600_1536000# diff_1147200_1458000# diff_548400_1543200# GND efet w=9600 l=7200
+ ad=2.5632e+08 pd=72000 as=0 ps=0 
M1976 GND diff_1155600_1536000# diff_1180800_1554000# GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1977 diff_1226400_1550400# diff_1215600_1537200# GND GND efet w=25800 l=7800
+ ad=2.376e+08 pd=76800 as=0 ps=0 
M1978 diff_664800_1543200# diff_1220400_1442400# diff_1226400_1550400# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1979 GND diff_1292400_1677600# diff_1317600_1696800# GND efet w=23400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1980 diff_1363200_1692000# diff_1353600_1677600# GND GND efet w=22800 l=7200
+ ad=2.376e+08 pd=72000 as=0 ps=0 
M1981 diff_664800_1683600# diff_1357200_1444800# diff_1363200_1692000# GND efet w=20400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1982 diff_1317600_1588800# diff_1306800_1458000# diff_664800_1620000# GND efet w=21600 l=7200
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M1983 GND diff_1292400_1621200# diff_1317600_1588800# GND efet w=24000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1984 diff_1363200_1592400# diff_1353600_1620000# GND GND efet w=22800 l=7200
+ ad=2.3328e+08 pd=72000 as=0 ps=0 
M1985 GND diff_1430400_1819200# diff_1454400_1839600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1986 diff_1501200_1834800# diff_1490400_1819200# GND GND efet w=25200 l=7800
+ ad=2.3328e+08 pd=74400 as=0 ps=0 
M1987 diff_664800_1825200# diff_1495200_1443600# diff_1501200_1834800# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1988 diff_1454400_1730400# diff_1443600_1458000# diff_664800_1760400# GND efet w=22800 l=7200
+ ad=2.592e+08 pd=76800 as=0 ps=0 
M1989 GND diff_1430400_1764000# diff_1454400_1730400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1990 diff_1501200_1734000# diff_1490400_1761600# GND GND efet w=22800 l=8400
+ ad=2.3328e+08 pd=72000 as=0 ps=0 
M1991 GND diff_1567200_1962000# diff_1592400_1981200# GND efet w=22800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1992 diff_1638000_1976400# diff_1628400_1962000# GND GND efet w=22800 l=7200
+ ad=2.5632e+08 pd=76800 as=0 ps=0 
M1993 diff_664800_1966800# diff_1633200_1442400# diff_1638000_1976400# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1994 diff_1592400_1872000# diff_1581600_1458000# diff_664800_1902000# GND efet w=21600 l=7200
+ ad=2.4624e+08 pd=74400 as=0 ps=0 
M1995 GND diff_1567200_1904400# diff_1592400_1872000# GND efet w=24000 l=8400
+ ad=0 pd=0 as=0 ps=0 
M1996 diff_1638000_1875600# diff_1628400_1903200# GND GND efet w=24000 l=7200
+ ad=2.6928e+08 pd=79200 as=0 ps=0 
M1997 diff_1730400_2014800# diff_1719600_1458000# diff_664800_2044800# GND efet w=21600 l=8400
+ ad=2.1888e+08 pd=72000 as=0 ps=0 
M1998 GND diff_1705200_2047200# diff_1730400_2014800# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1999 diff_1776000_2018400# diff_1766400_2044800# GND GND efet w=22800 l=7200
+ ad=2.376e+08 pd=74400 as=0 ps=0 
M2000 GND diff_1842000_2251200# diff_1867200_2265600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2001 diff_1914000_2259600# diff_1903200_2246400# GND GND efet w=27000 l=7800
+ ad=2.3904e+08 pd=72000 as=0 ps=0 
M2002 diff_664800_2251200# diff_1908000_1442400# diff_1914000_2259600# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2003 diff_1867200_2156400# diff_1856400_1458000# diff_664800_2186400# GND efet w=21600 l=7200
+ ad=2.5776e+08 pd=76800 as=0 ps=0 
M2004 GND diff_1843200_2188800# diff_1867200_2156400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2005 diff_1914000_2160000# diff_1903200_2187600# GND GND efet w=25200 l=7200
+ ad=2.3184e+08 pd=72000 as=0 ps=0 
M2006 GND diff_1980000_2386800# diff_2005200_2407200# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2007 diff_2052000_2402400# diff_2041200_2386800# GND GND efet w=22200 l=7800
+ ad=2.232e+08 pd=69600 as=0 ps=0 
M2008 diff_664800_2392800# diff_2046000_1444800# diff_2052000_2402400# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2009 diff_2005200_2298000# diff_1994400_1460400# diff_664800_2328000# GND efet w=21600 l=7200
+ ad=2.6208e+08 pd=76800 as=0 ps=0 
M2010 GND diff_1980000_2330400# diff_2005200_2298000# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2011 diff_2052000_2301600# diff_2041200_2329200# GND GND efet w=27000 l=7800
+ ad=2.3184e+08 pd=72000 as=0 ps=0 
M2012 Vdd diff_2224800_1584000# diff_664800_2534400# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2013 Vdd diff_1892400_663600# diff_548400_2534400# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2014 GND diff_2074800_2772000# diff_2424000_2518800# GND efet w=15600 l=6000
+ ad=0 pd=0 as=3.8736e+08 ps=84000 
M2015 GND diff_2077200_2900400# diff_2344800_2570400# GND efet w=28200 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2016 diff_2424000_2518800# Vdd Vdd GND efet w=8400 l=57600
+ ad=0 pd=0 as=0 ps=0 
M2017 Vdd Vdd Vdd GND efet w=6000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2018 diff_2344800_2570400# diff_2424000_2518800# diff_2455200_2494800# GND efet w=14400 l=7200
+ ad=0 pd=0 as=6.3792e+08 ps=139200 
M2019 diff_2414400_2601600# diff_2344800_2570400# GND GND efet w=112200 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2020 Vdd Vdd Vdd GND efet w=4200 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2021 diff_2455200_2494800# Vdd Vdd GND efet w=10800 l=28200
+ ad=0 pd=0 as=0 ps=0 
M2022 Vdd diff_1892400_663600# diff_548400_2460000# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2023 diff_2143200_2439600# diff_2133600_1458000# diff_663600_2470800# GND efet w=21600 l=7200
+ ad=2.6064e+08 pd=74400 as=0 ps=0 
M2024 GND diff_2118000_2472000# diff_2143200_2439600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2025 Vdd diff_2224800_1584000# diff_663600_2470800# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2026 o2 diff_2374800_2434800# Vdd GND efet w=207000 l=6600
+ ad=-3.79607e+08 pd=698400 as=0 ps=0 
M2027 diff_2143200_2407200# diff_2133600_1458000# diff_664800_2392800# GND efet w=21600 l=7200
+ ad=2.592e+08 pd=76800 as=0 ps=0 
M2028 diff_548400_2392800# diff_2082000_1496400# diff_2041200_2386800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6208e+08 ps=74400 
M2029 diff_2118000_2386800# diff_2110800_1458000# diff_548400_2392800# GND efet w=8400 l=7200
+ ad=2.592e+08 pd=76800 as=0 ps=0 
M2030 diff_548400_2319600# diff_2082000_1496400# diff_2041200_2329200# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6352e+08 ps=74400 
M2031 diff_2118000_2330400# diff_2110800_1458000# diff_548400_2319600# GND efet w=8400 l=7200
+ ad=2.592e+08 pd=76800 as=0 ps=0 
M2032 diff_664800_2328000# diff_2046000_1444800# diff_2052000_2301600# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2033 diff_2005200_2265600# diff_1994400_1460400# diff_664800_2251200# GND efet w=20400 l=7200
+ ad=2.6064e+08 pd=76800 as=0 ps=0 
M2034 diff_548400_2252400# diff_1944000_1496400# diff_1903200_2246400# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.664e+08 ps=76800 
M2035 diff_1980000_2245200# diff_1972800_1458000# diff_548400_2252400# GND efet w=8400 l=7200
+ ad=2.5776e+08 pd=76800 as=0 ps=0 
M2036 diff_548400_2178000# diff_1944000_1496400# diff_1903200_2187600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6352e+08 ps=74400 
M2037 diff_1980000_2190000# diff_1972800_1458000# diff_548400_2178000# GND efet w=7200 l=7200
+ ad=2.6064e+08 pd=76800 as=0 ps=0 
M2038 diff_664800_2186400# diff_1908000_1442400# diff_1914000_2160000# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2039 diff_1867200_2124000# diff_1856400_1458000# diff_664800_2109600# GND efet w=21600 l=7200
+ ad=2.6064e+08 pd=74400 as=0 ps=0 
M2040 diff_548400_2109600# diff_1806000_1496400# diff_1765200_2109600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6496e+08 ps=79200 
M2041 diff_1843200_2103600# diff_1834800_1458000# diff_548400_2109600# GND efet w=9000 l=8400
+ ad=2.6064e+08 pd=76800 as=0 ps=0 
M2042 diff_548400_2036400# diff_1806000_1496400# diff_1766400_2044800# GND efet w=9600 l=7200
+ ad=0 pd=0 as=2.7072e+08 ps=76800 
M2043 diff_1843200_2047200# diff_1834800_1458000# diff_548400_2036400# GND efet w=9600 l=7200
+ ad=2.6208e+08 pd=76800 as=0 ps=0 
M2044 diff_664800_2044800# diff_1770000_1443600# diff_1776000_2018400# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2045 diff_1730400_1981200# diff_1719600_1458000# diff_664800_1966800# GND efet w=21000 l=9000
+ ad=2.376e+08 pd=74400 as=0 ps=0 
M2046 diff_548400_1968000# diff_1668000_1497600# diff_1628400_1962000# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.4048e+08 ps=74400 
M2047 diff_1705200_1962000# diff_1696800_1458000# diff_548400_1968000# GND efet w=8400 l=7200
+ ad=2.3904e+08 pd=74400 as=0 ps=0 
M2048 diff_548400_1893600# diff_1668000_1497600# diff_1628400_1903200# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.52e+08 ps=74400 
M2049 diff_1705200_1904400# diff_1696800_1458000# diff_548400_1893600# GND efet w=8400 l=7200
+ ad=2.664e+08 pd=79200 as=0 ps=0 
M2050 diff_664800_1902000# diff_1633200_1442400# diff_1638000_1875600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2051 diff_1592400_1838400# diff_1581600_1458000# diff_664800_1825200# GND efet w=21600 l=7200
+ ad=2.4048e+08 pd=74400 as=0 ps=0 
M2052 diff_664800_1825200# diff_1633200_1442400# diff_1638000_1833600# GND efet w=27000 l=7200
+ ad=0 pd=0 as=2.5632e+08 ps=86400 
M2053 diff_548400_1826400# diff_1531200_1458000# diff_1490400_1819200# GND efet w=9000 l=7800
+ ad=0 pd=0 as=2.664e+08 ps=74400 
M2054 diff_1567200_1819200# diff_1558800_1458000# diff_548400_1826400# GND efet w=9600 l=8400
+ ad=2.664e+08 pd=74400 as=0 ps=0 
M2055 diff_548400_1752000# diff_1531200_1458000# diff_1490400_1761600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6208e+08 ps=74400 
M2056 diff_1567200_1764000# diff_1558800_1458000# diff_548400_1752000# GND efet w=8400 l=7200
+ ad=2.6496e+08 pd=74400 as=0 ps=0 
M2057 diff_664800_1760400# diff_1495200_1443600# diff_1501200_1734000# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2058 diff_1454400_1696800# diff_1443600_1458000# diff_664800_1683600# GND efet w=20400 l=7200
+ ad=2.6208e+08 pd=74400 as=0 ps=0 
M2059 diff_548400_1684800# diff_1393200_1496400# diff_1353600_1677600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6928e+08 ps=76800 
M2060 diff_1430400_1677600# diff_1422000_1458000# diff_548400_1684800# GND efet w=9000 l=7800
+ ad=2.5344e+08 pd=72000 as=0 ps=0 
M2061 diff_548400_1610400# diff_1393200_1496400# diff_1353600_1620000# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6496e+08 ps=74400 
M2062 diff_1430400_1621200# diff_1422000_1458000# diff_548400_1610400# GND efet w=8400 l=7200
+ ad=2.5344e+08 pd=72000 as=0 ps=0 
M2063 diff_664800_1620000# diff_1357200_1444800# diff_1363200_1592400# GND efet w=21600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2064 diff_1317600_1555200# diff_1306800_1458000# diff_664800_1543200# GND efet w=21600 l=7200
+ ad=2.3616e+08 pd=74400 as=0 ps=0 
M2065 diff_548400_1543200# diff_1256400_1458000# diff_1215600_1537200# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6928e+08 ps=79200 
M2066 diff_1292400_1536000# diff_1284000_1458000# diff_548400_1543200# GND efet w=8400 l=7200
+ ad=2.5776e+08 pd=76800 as=0 ps=0 
M2067 GND diff_1292400_1536000# diff_1317600_1555200# GND efet w=22800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2068 diff_1363200_1551600# diff_1353600_1537200# GND GND efet w=22800 l=7200
+ ad=2.3184e+08 pd=72000 as=0 ps=0 
M2069 diff_664800_1543200# diff_1357200_1444800# diff_1363200_1551600# GND efet w=21600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2070 GND diff_1430400_1677600# diff_1454400_1696800# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2071 diff_1501200_1692000# diff_1490400_1677600# GND GND efet w=22800 l=8400
+ ad=2.3328e+08 pd=74400 as=0 ps=0 
M2072 diff_664800_1683600# diff_1495200_1443600# diff_1501200_1692000# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2073 diff_1454400_1588800# diff_1443600_1458000# diff_664800_1620000# GND efet w=21600 l=7200
+ ad=2.6208e+08 pd=74400 as=0 ps=0 
M2074 GND diff_1430400_1621200# diff_1454400_1588800# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2075 diff_1501200_1592400# diff_1490400_1620000# GND GND efet w=22800 l=8400
+ ad=2.3328e+08 pd=72000 as=0 ps=0 
M2076 GND diff_1567200_1819200# diff_1592400_1838400# GND efet w=23400 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2077 diff_1638000_1833600# diff_1628400_1819200# GND GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2078 GND diff_1705200_1962000# diff_1730400_1981200# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2079 diff_1776000_1976400# diff_1766400_1960800# GND GND efet w=22800 l=7200
+ ad=2.3616e+08 pd=74400 as=0 ps=0 
M2080 diff_664800_1966800# diff_1770000_1443600# diff_1776000_1976400# GND efet w=21000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2081 diff_1730400_1872000# diff_1719600_1458000# diff_664800_1902000# GND efet w=21600 l=8400
+ ad=2.448e+08 pd=74400 as=0 ps=0 
M2082 GND diff_1705200_1904400# diff_1730400_1872000# GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2083 diff_1776000_1875600# diff_1765200_1904400# GND GND efet w=24000 l=7200
+ ad=2.4624e+08 pd=74400 as=0 ps=0 
M2084 GND diff_1843200_2103600# diff_1867200_2124000# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2085 diff_1914000_2119200# diff_1903200_2103600# GND GND efet w=22800 l=7200
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M2086 diff_664800_2109600# diff_1908000_1442400# diff_1914000_2119200# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2087 diff_1867200_2014800# diff_1856400_1458000# diff_664800_2044800# GND efet w=21600 l=7200
+ ad=2.6208e+08 pd=76800 as=0 ps=0 
M2088 GND diff_1843200_2047200# diff_1867200_2014800# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2089 diff_1914000_2018400# diff_1903200_2044800# GND GND efet w=22800 l=7200
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M2090 diff_548400_2109600# diff_1944000_1496400# diff_1903200_2103600# GND efet w=7200 l=7200
+ ad=0 pd=0 as=2.6928e+08 ps=76800 
M2091 GND diff_1980000_2245200# diff_2005200_2265600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2092 diff_2052000_2259600# diff_2041200_2246400# GND GND efet w=24600 l=7800
+ ad=2.3184e+08 pd=72000 as=0 ps=0 
M2093 diff_664800_2251200# diff_2046000_1444800# diff_2052000_2259600# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2094 diff_2005200_2157600# diff_1994400_1460400# diff_664800_2186400# GND efet w=20400 l=7200
+ ad=2.5488e+08 pd=74400 as=0 ps=0 
M2095 GND diff_1980000_2190000# diff_2005200_2157600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2096 diff_2052000_2160000# diff_2041200_2187600# GND GND efet w=22800 l=7800
+ ad=2.2464e+08 pd=69600 as=0 ps=0 
M2097 GND diff_2118000_2386800# diff_2143200_2407200# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2098 diff_2455200_2494800# diff_2414400_2601600# GND GND efet w=25200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2099 o2 diff_2414400_2601600# GND GND efet w=196800 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2100 Vdd diff_2224800_1584000# diff_664800_2392800# GND efet w=14400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2101 Vdd diff_1892400_663600# diff_548400_2392800# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2102 diff_2374800_2434800# diff_2374800_2434800# diff_2374800_2434800# GND efet w=1800 l=3600
+ ad=9.8064e+08 pd=168000 as=0 ps=0 
M2103 diff_2374800_2434800# diff_2374800_2434800# diff_2374800_2434800# GND efet w=2400 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2104 diff_2374800_2434800# Vdd Vdd GND efet w=10800 l=19200
+ ad=0 pd=0 as=0 ps=0 
M2105 GND diff_2414400_2601600# diff_2374800_2434800# GND efet w=49800 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2106 Vdd diff_1892400_663600# diff_548400_2319600# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2107 diff_2143200_2298000# diff_2133600_1458000# diff_664800_2328000# GND efet w=21600 l=7200
+ ad=2.6208e+08 pd=76800 as=0 ps=0 
M2108 GND diff_2118000_2330400# diff_2143200_2298000# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2109 Vdd diff_2224800_1584000# diff_664800_2328000# GND efet w=14400 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2110 diff_2143200_2265600# diff_2133600_1458000# diff_664800_2251200# GND efet w=20400 l=7200
+ ad=2.52e+08 pd=76800 as=0 ps=0 
M2111 diff_548400_2252400# diff_2082000_1496400# diff_2041200_2246400# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6064e+08 ps=74400 
M2112 diff_2118000_2245200# diff_2110800_1458000# diff_548400_2252400# GND efet w=8400 l=7200
+ ad=2.5776e+08 pd=74400 as=0 ps=0 
M2113 diff_548400_2178000# diff_2082000_1496400# diff_2041200_2187600# GND efet w=7200 l=7200
+ ad=0 pd=0 as=2.6208e+08 ps=74400 
M2114 diff_2118000_2190000# diff_2110800_1458000# diff_548400_2178000# GND efet w=7200 l=7200
+ ad=2.5632e+08 pd=76800 as=0 ps=0 
M2115 diff_664800_2186400# diff_2046000_1444800# diff_2052000_2160000# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2116 diff_2005200_2124000# diff_1994400_1460400# diff_664800_2109600# GND efet w=21600 l=7200
+ ad=2.592e+08 pd=74400 as=0 ps=0 
M2117 diff_1980000_2104800# diff_1972800_1458000# diff_548400_2109600# GND efet w=7200 l=7200
+ ad=2.6496e+08 pd=79200 as=0 ps=0 
M2118 diff_548400_2036400# diff_1944000_1496400# diff_1903200_2044800# GND efet w=9600 l=7200
+ ad=0 pd=0 as=2.7216e+08 ps=76800 
M2119 diff_1980000_2047200# diff_1972800_1458000# diff_548400_2036400# GND efet w=8400 l=7200
+ ad=2.5776e+08 pd=74400 as=0 ps=0 
M2120 diff_664800_2044800# diff_1908000_1442400# diff_1914000_2018400# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2121 diff_1867200_1982400# diff_1856400_1458000# diff_664800_1966800# GND efet w=20400 l=7200
+ ad=2.6208e+08 pd=76800 as=0 ps=0 
M2122 diff_548400_1968000# diff_1806000_1496400# diff_1766400_1960800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.592e+08 ps=81600 
M2123 diff_1843200_1962000# diff_1834800_1458000# diff_548400_1968000# GND efet w=8400 l=7200
+ ad=2.4768e+08 pd=79200 as=0 ps=0 
M2124 diff_548400_1893600# diff_1806000_1496400# diff_1765200_1904400# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.5488e+08 ps=79200 
M2125 diff_1843200_1905600# diff_1834800_1458000# diff_548400_1893600# GND efet w=10200 l=7800
+ ad=2.5488e+08 pd=79200 as=0 ps=0 
M2126 diff_664800_1902000# diff_1770000_1443600# diff_1776000_1875600# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2127 diff_1730400_1838400# diff_1719600_1458000# diff_664800_1825200# GND efet w=21600 l=8400
+ ad=2.4192e+08 pd=74400 as=0 ps=0 
M2128 diff_548400_1826400# diff_1668000_1497600# diff_1628400_1819200# GND efet w=9600 l=7200
+ ad=0 pd=0 as=2.5632e+08 ps=74400 
M2129 diff_1705200_1819200# diff_1696800_1458000# diff_548400_1826400# GND efet w=9600 l=7200
+ ad=2.592e+08 pd=76800 as=0 ps=0 
M2130 GND diff_1705200_1819200# diff_1730400_1838400# GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2131 diff_1776000_1833600# diff_1765200_1822800# GND GND efet w=24000 l=7200
+ ad=2.4192e+08 pd=74400 as=0 ps=0 
M2132 diff_664800_1825200# diff_1770000_1443600# diff_1776000_1833600# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2133 diff_548400_1752000# diff_1668000_1497600# diff_1628400_1760400# GND efet w=7200 l=7800
+ ad=0 pd=0 as=2.5344e+08 ps=76800 
M2134 diff_1705200_1764000# diff_1696800_1458000# diff_548400_1752000# GND efet w=7800 l=7800
+ ad=2.5632e+08 pd=76800 as=0 ps=0 
M2135 diff_1592400_1730400# diff_1581600_1458000# diff_664800_1760400# GND efet w=21600 l=7200
+ ad=2.376e+08 pd=74400 as=0 ps=0 
M2136 GND diff_1567200_1764000# diff_1592400_1730400# GND efet w=22800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2137 diff_1638000_1734000# diff_1628400_1760400# GND GND efet w=22800 l=7200
+ ad=2.448e+08 pd=81600 as=0 ps=0 
M2138 diff_664800_1760400# diff_1633200_1442400# diff_1638000_1734000# GND efet w=24600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2139 diff_1592400_1696800# diff_1581600_1458000# diff_664800_1683600# GND efet w=20400 l=7200
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M2140 diff_548400_1684800# diff_1531200_1458000# diff_1490400_1677600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6352e+08 ps=74400 
M2141 diff_1567200_1677600# diff_1558800_1458000# diff_548400_1684800# GND efet w=8400 l=7200
+ ad=2.664e+08 pd=74400 as=0 ps=0 
M2142 diff_548400_1610400# diff_1531200_1458000# diff_1490400_1620000# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.6496e+08 ps=79200 
M2143 diff_1567200_1621200# diff_1558800_1458000# diff_548400_1610400# GND efet w=8400 l=7200
+ ad=2.52e+08 pd=74400 as=0 ps=0 
M2144 diff_664800_1620000# diff_1495200_1443600# diff_1501200_1592400# GND efet w=21000 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2145 diff_1454400_1556400# diff_1443600_1458000# diff_664800_1543200# GND efet w=24000 l=8400
+ ad=2.5488e+08 pd=79200 as=0 ps=0 
M2146 diff_548400_1543200# diff_1393200_1496400# diff_1353600_1537200# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.664e+08 ps=74400 
M2147 diff_1430400_1536000# diff_1422000_1458000# diff_548400_1543200# GND efet w=8400 l=7200
+ ad=2.5344e+08 pd=72000 as=0 ps=0 
M2148 GND diff_1430400_1536000# diff_1454400_1556400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2149 diff_1501200_1551600# diff_1490400_1537200# GND GND efet w=21600 l=8400
+ ad=2.3184e+08 pd=76800 as=0 ps=0 
M2150 diff_664800_1543200# diff_1495200_1443600# diff_1501200_1551600# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2151 GND diff_1567200_1677600# diff_1592400_1696800# GND efet w=22800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2152 diff_1638000_1692000# diff_1628400_1677600# GND GND efet w=22800 l=7200
+ ad=2.3616e+08 pd=74400 as=0 ps=0 
M2153 diff_664800_1683600# diff_1633200_1442400# diff_1638000_1692000# GND efet w=20400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2154 diff_1730400_1730400# diff_1719600_1458000# diff_664800_1760400# GND efet w=21600 l=8400
+ ad=2.2032e+08 pd=74400 as=0 ps=0 
M2155 GND diff_1705200_1764000# diff_1730400_1730400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2156 diff_1776000_1734000# diff_1765200_1762800# GND GND efet w=22800 l=7200
+ ad=2.376e+08 pd=74400 as=0 ps=0 
M2157 GND diff_1843200_1962000# diff_1867200_1982400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2158 diff_1914000_1976400# diff_1903200_1962000# GND GND efet w=22800 l=7200
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M2159 diff_664800_1966800# diff_1908000_1442400# diff_1914000_1976400# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2160 diff_1867200_1872000# diff_1856400_1458000# diff_664800_1902000# GND efet w=21600 l=7200
+ ad=2.6928e+08 pd=76800 as=0 ps=0 
M2161 GND diff_1843200_1905600# diff_1867200_1872000# GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2162 diff_1914000_1875600# diff_1903200_1903200# GND GND efet w=24000 l=7200
+ ad=2.448e+08 pd=74400 as=0 ps=0 
M2163 GND diff_1980000_2104800# diff_2005200_2124000# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2164 diff_2052000_2119200# diff_2041200_2103600# GND GND efet w=25800 l=7800
+ ad=2.3184e+08 pd=72000 as=0 ps=0 
M2165 diff_664800_2109600# diff_2046000_1444800# diff_2052000_2119200# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2166 diff_2005200_2014800# diff_1994400_1460400# diff_664800_2044800# GND efet w=21600 l=7200
+ ad=2.6208e+08 pd=76800 as=0 ps=0 
M2167 GND diff_1980000_2047200# diff_2005200_2014800# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2168 diff_2052000_2018400# diff_2041200_2044800# GND GND efet w=23400 l=7800
+ ad=2.3184e+08 pd=72000 as=0 ps=0 
M2169 GND diff_2118000_2245200# diff_2143200_2265600# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2170 Vdd diff_2224800_1584000# diff_664800_2251200# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2171 Vdd diff_1892400_663600# diff_548400_2252400# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2172 Vdd diff_1892400_663600# diff_548400_2178000# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2173 GND diff_2118000_2190000# diff_2143200_2157600# GND efet w=22200 l=7800
+ ad=0 pd=0 as=2.52e+08 ps=74400 
M2174 diff_2143200_2157600# diff_2133600_1458000# diff_664800_2186400# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2175 Vdd diff_2224800_1584000# diff_664800_2186400# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2176 diff_2416800_1954800# Vdd Vdd GND efet w=10800 l=19200
+ ad=1.31616e+09 pd=261600 as=0 ps=0 
M2177 diff_2325600_2148000# clk2 diff_231600_1357200# GND efet w=19200 l=7200
+ ad=2.6928e+08 pd=76800 as=0 ps=0 
M2178 diff_2143200_2124000# diff_2133600_1458000# diff_664800_2109600# GND efet w=21600 l=7200
+ ad=2.6064e+08 pd=74400 as=0 ps=0 
M2179 diff_548400_2109600# diff_2082000_1496400# diff_2041200_2103600# GND efet w=7200 l=7200
+ ad=0 pd=0 as=2.592e+08 ps=74400 
M2180 diff_2118000_2104800# diff_2110800_1458000# diff_548400_2109600# GND efet w=7200 l=7200
+ ad=2.592e+08 pd=76800 as=0 ps=0 
M2181 diff_548400_2036400# diff_2082000_1496400# diff_2041200_2044800# GND efet w=8400 l=8400
+ ad=0 pd=0 as=2.592e+08 ps=74400 
M2182 diff_2118000_2048400# diff_2110800_1458000# diff_548400_2036400# GND efet w=7200 l=7200
+ ad=2.6064e+08 pd=76800 as=0 ps=0 
M2183 diff_664800_2044800# diff_2046000_1444800# diff_2052000_2018400# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2184 diff_2005200_1982400# diff_1994400_1460400# diff_664800_1966800# GND efet w=20400 l=7200
+ ad=2.592e+08 pd=74400 as=0 ps=0 
M2185 diff_548400_1968000# diff_1944000_1496400# diff_1903200_1962000# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.5632e+08 ps=76800 
M2186 diff_1980000_1962000# diff_1972800_1458000# diff_548400_1968000# GND efet w=8400 l=7200
+ ad=2.592e+08 pd=76800 as=0 ps=0 
M2187 diff_548400_1893600# diff_1944000_1496400# diff_1903200_1903200# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.664e+08 ps=76800 
M2188 diff_1980000_1905600# diff_1972800_1458000# diff_548400_1893600# GND efet w=8400 l=7200
+ ad=2.6208e+08 pd=79200 as=0 ps=0 
M2189 diff_664800_1902000# diff_1908000_1442400# diff_1914000_1875600# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2190 diff_1867200_1839600# diff_1856400_1458000# diff_664800_1825200# GND efet w=21600 l=7200
+ ad=2.6352e+08 pd=74400 as=0 ps=0 
M2191 diff_548400_1826400# diff_1806000_1496400# diff_1765200_1822800# GND efet w=9600 l=7200
+ ad=0 pd=0 as=2.6496e+08 ps=79200 
M2192 diff_1843200_1819200# diff_1834800_1458000# diff_548400_1826400# GND efet w=11400 l=7800
+ ad=2.5776e+08 pd=76800 as=0 ps=0 
M2193 diff_548400_1752000# diff_1806000_1496400# diff_1765200_1762800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.7072e+08 ps=76800 
M2194 diff_1843200_1762800# diff_1834800_1458000# diff_548400_1752000# GND efet w=8400 l=8400
+ ad=2.6208e+08 pd=76800 as=0 ps=0 
M2195 diff_664800_1760400# diff_1770000_1443600# diff_1776000_1734000# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2196 diff_1730400_1696800# diff_1719600_1458000# diff_664800_1683600# GND efet w=20400 l=8400
+ ad=2.3616e+08 pd=74400 as=0 ps=0 
M2197 diff_664800_1683600# diff_1770000_1443600# diff_1776000_1692000# GND efet w=21600 l=8400
+ ad=0 pd=0 as=2.376e+08 ps=72000 
M2198 diff_548400_1684800# diff_1668000_1497600# diff_1628400_1677600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.5344e+08 ps=76800 
M2199 diff_1705200_1677600# diff_1696800_1458000# diff_548400_1684800# GND efet w=8400 l=7200
+ ad=2.5488e+08 pd=74400 as=0 ps=0 
M2200 diff_1592400_1588800# diff_1581600_1458000# diff_664800_1620000# GND efet w=21000 l=7800
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M2201 GND diff_1567200_1621200# diff_1592400_1588800# GND efet w=22800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2202 diff_1638000_1592400# diff_1628400_1620000# GND GND efet w=22800 l=7200
+ ad=2.3904e+08 pd=74400 as=0 ps=0 
M2203 GND diff_1705200_1677600# diff_1730400_1696800# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2204 diff_1776000_1692000# diff_1765200_1678800# GND GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2205 diff_548400_1610400# diff_1668000_1497600# diff_1628400_1620000# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.5056e+08 ps=74400 
M2206 diff_1705200_1621200# diff_1696800_1458000# diff_548400_1610400# GND efet w=8400 l=7200
+ ad=2.4336e+08 pd=76800 as=0 ps=0 
M2207 diff_664800_1620000# diff_1633200_1442400# diff_1638000_1592400# GND efet w=22200 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2208 diff_1592400_1555200# diff_1581600_1458000# diff_664800_1543200# GND efet w=20400 l=7200
+ ad=2.3472e+08 pd=74400 as=0 ps=0 
M2209 diff_664800_1543200# diff_1633200_1442400# diff_1638000_1550400# GND efet w=21000 l=7800
+ ad=0 pd=0 as=2.3904e+08 ps=76800 
M2210 diff_548400_1543200# diff_1531200_1458000# diff_1490400_1537200# GND efet w=9600 l=7200
+ ad=0 pd=0 as=2.7216e+08 ps=79200 
M2211 diff_1567200_1536000# diff_1558800_1458000# diff_548400_1543200# GND efet w=9600 l=7200
+ ad=2.6784e+08 pd=74400 as=0 ps=0 
M2212 GND diff_1567200_1536000# diff_1592400_1555200# GND efet w=22800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2213 diff_1638000_1550400# diff_1628400_1537200# GND GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2214 diff_1730400_1588800# diff_1719600_1458000# diff_664800_1620000# GND efet w=21000 l=9000
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M2215 GND diff_1705200_1621200# diff_1730400_1588800# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2216 diff_1776000_1592400# diff_1765200_1621200# GND GND efet w=22800 l=7200
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M2217 GND diff_1843200_1819200# diff_1867200_1839600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2218 diff_1914000_1834800# diff_1903200_1820400# GND GND efet w=22800 l=7200
+ ad=2.3616e+08 pd=72000 as=0 ps=0 
M2219 diff_664800_1825200# diff_1908000_1442400# diff_1914000_1834800# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2220 diff_1867200_1730400# diff_1856400_1458000# diff_664800_1760400# GND efet w=21600 l=7200
+ ad=2.6352e+08 pd=76800 as=0 ps=0 
M2221 GND diff_1843200_1762800# diff_1867200_1730400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2222 diff_1914000_1734000# diff_1903200_1761600# GND GND efet w=22800 l=7200
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M2223 GND diff_1980000_1962000# diff_2005200_1982400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2224 diff_2052000_1976400# diff_2041200_1962000# GND GND efet w=22800 l=7200
+ ad=2.3328e+08 pd=74400 as=0 ps=0 
M2225 diff_664800_1966800# diff_2046000_1444800# diff_2052000_1976400# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2226 diff_2005200_1873200# diff_1994400_1460400# diff_664800_1902000# GND efet w=20400 l=7200
+ ad=2.6208e+08 pd=74400 as=0 ps=0 
M2227 GND diff_1980000_1905600# diff_2005200_1873200# GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2228 diff_2052000_1875600# diff_2041200_1903200# GND GND efet w=22800 l=7200
+ ad=2.2464e+08 pd=69600 as=0 ps=0 
M2229 GND diff_2118000_2104800# diff_2143200_2124000# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2230 diff_2344800_2140800# diff_2074800_2772000# diff_2325600_2148000# GND efet w=19200 l=7200
+ ad=1.69488e+09 pd=336000 as=0 ps=0 
M2231 Vdd diff_2224800_1584000# diff_664800_2109600# GND efet w=15600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2232 GND diff_2074800_2772000# diff_2425200_2089200# GND efet w=14400 l=6600
+ ad=0 pd=0 as=3.4704e+08 ps=79200 
M2233 GND diff_2077200_2900400# diff_2344800_2140800# GND efet w=27600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2234 Vdd diff_1892400_663600# diff_548400_2109600# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2235 diff_2425200_2089200# Vdd Vdd GND efet w=9000 l=58200
+ ad=0 pd=0 as=0 ps=0 
M2236 Vdd Vdd Vdd GND efet w=6000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2237 Vdd diff_1892400_663600# diff_548400_2036400# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2238 diff_2344800_2140800# diff_2425200_2089200# diff_2455200_2066400# GND efet w=14400 l=6000
+ ad=0 pd=0 as=6.5952e+08 ps=146400 
M2239 diff_2416800_1954800# diff_2344800_2140800# GND GND efet w=111600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2240 Vdd Vdd Vdd GND efet w=4800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2241 diff_2455200_2066400# Vdd Vdd GND efet w=9600 l=30600
+ ad=0 pd=0 as=0 ps=0 
M2242 diff_2143200_2014800# diff_2133600_1458000# diff_664800_2044800# GND efet w=21600 l=7200
+ ad=2.6208e+08 pd=76800 as=0 ps=0 
M2243 GND diff_2118000_2048400# diff_2143200_2014800# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2244 Vdd diff_2224800_1584000# diff_664800_2044800# GND efet w=15600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2245 diff_2143200_1982400# diff_2133600_1458000# diff_664800_1966800# GND efet w=20400 l=7200
+ ad=2.592e+08 pd=76800 as=0 ps=0 
M2246 diff_548400_1968000# diff_2082000_1496400# diff_2041200_1962000# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.52e+08 ps=74400 
M2247 diff_2118000_1962000# diff_2110800_1458000# diff_548400_1968000# GND efet w=8400 l=7200
+ ad=2.52e+08 pd=79200 as=0 ps=0 
M2248 diff_548400_1893600# diff_2082000_1496400# diff_2041200_1903200# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.5632e+08 ps=74400 
M2249 diff_2118000_1905600# diff_2110800_1458000# diff_548400_1893600# GND efet w=8400 l=7200
+ ad=2.5344e+08 pd=76800 as=0 ps=0 
M2250 diff_664800_1902000# diff_2046000_1444800# diff_2052000_1875600# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2251 diff_2005200_1839600# diff_1994400_1460400# diff_664800_1825200# GND efet w=21600 l=7200
+ ad=2.6064e+08 pd=74400 as=0 ps=0 
M2252 diff_548400_1826400# diff_1944000_1496400# diff_1903200_1820400# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.664e+08 ps=74400 
M2253 diff_1980000_1820400# diff_1972800_1458000# diff_548400_1826400# GND efet w=9600 l=7200
+ ad=2.4768e+08 pd=76800 as=0 ps=0 
M2254 diff_548400_1752000# diff_1944000_1496400# diff_1903200_1761600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6208e+08 ps=74400 
M2255 diff_1980000_1764000# diff_1972800_1458000# diff_548400_1752000# GND efet w=8400 l=7200
+ ad=2.5632e+08 pd=76800 as=0 ps=0 
M2256 diff_664800_1760400# diff_1908000_1442400# diff_1914000_1734000# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2257 diff_1867200_1698000# diff_1856400_1458000# diff_664800_1683600# GND efet w=20400 l=7200
+ ad=2.6208e+08 pd=76800 as=0 ps=0 
M2258 diff_548400_1684800# diff_1806000_1496400# diff_1765200_1678800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.664e+08 ps=74400 
M2259 diff_1843200_1677600# diff_1834800_1458000# diff_548400_1684800# GND efet w=8400 l=8400
+ ad=2.5632e+08 pd=76800 as=0 ps=0 
M2260 diff_548400_1610400# diff_1806000_1496400# diff_1765200_1621200# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6496e+08 ps=74400 
M2261 diff_1843200_1621200# diff_1834800_1458000# diff_548400_1610400# GND efet w=8400 l=8400
+ ad=2.4912e+08 pd=79200 as=0 ps=0 
M2262 diff_664800_1620000# diff_1770000_1443600# diff_1776000_1592400# GND efet w=21000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2263 diff_1730400_1555200# diff_1719600_1458000# diff_664800_1543200# GND efet w=20400 l=8400
+ ad=2.3616e+08 pd=74400 as=0 ps=0 
M2264 diff_664800_1543200# diff_1770000_1443600# diff_1776000_1550400# GND efet w=20400 l=8400
+ ad=0 pd=0 as=2.376e+08 ps=72000 
M2265 diff_548400_1543200# diff_1668000_1497600# diff_1628400_1537200# GND efet w=9600 l=7200
+ ad=0 pd=0 as=2.5488e+08 ps=74400 
M2266 diff_1705200_1536000# diff_1696800_1458000# diff_548400_1543200# GND efet w=9600 l=7200
+ ad=2.5488e+08 pd=74400 as=0 ps=0 
M2267 GND diff_1705200_1536000# diff_1730400_1555200# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2268 diff_1776000_1550400# diff_1765200_1538400# GND GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2269 GND diff_1843200_1677600# diff_1867200_1698000# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2270 diff_1914000_1692000# diff_1903200_1678800# GND GND efet w=25200 l=8400
+ ad=2.376e+08 pd=72000 as=0 ps=0 
M2271 diff_664800_1683600# diff_1908000_1442400# diff_1914000_1692000# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2272 diff_1867200_1588800# diff_1856400_1458000# diff_664800_1620000# GND efet w=21000 l=7800
+ ad=2.6064e+08 pd=74400 as=0 ps=0 
M2273 GND diff_1843200_1621200# diff_1867200_1588800# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2274 diff_1914000_1592400# diff_1903200_1620000# GND GND efet w=23400 l=7800
+ ad=2.3472e+08 pd=72000 as=0 ps=0 
M2275 GND diff_1980000_1820400# diff_2005200_1839600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2276 diff_2052000_1834800# diff_2041200_1820400# GND GND efet w=22800 l=7200
+ ad=2.3184e+08 pd=72000 as=0 ps=0 
M2277 diff_664800_1825200# diff_2046000_1444800# diff_2052000_1834800# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2278 diff_2005200_1730400# diff_1994400_1460400# diff_664800_1760400# GND efet w=21600 l=7200
+ ad=2.6208e+08 pd=76800 as=0 ps=0 
M2279 GND diff_1980000_1764000# diff_2005200_1730400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2280 diff_2052000_1734000# diff_2041200_1761600# GND GND efet w=25200 l=7800
+ ad=2.3184e+08 pd=72000 as=0 ps=0 
M2281 GND diff_2118000_1962000# diff_2143200_1982400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2282 o3 diff_2374800_2004000# Vdd GND efet w=206400 l=7200
+ ad=-2.58647e+08 pd=684000 as=0 ps=0 
M2283 diff_2455200_2066400# diff_2416800_1954800# GND GND efet w=27600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2284 o3 diff_2416800_1954800# GND GND efet w=193800 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2285 Vdd diff_2224800_1584000# diff_664800_1966800# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2286 Vdd diff_1892400_663600# diff_548400_1968000# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2287 diff_2374800_2004000# diff_2374800_2004000# diff_2374800_2004000# GND efet w=1800 l=3000
+ ad=9.8496e+08 pd=172800 as=0 ps=0 
M2288 diff_2374800_2004000# Vdd Vdd GND efet w=12000 l=18600
+ ad=0 pd=0 as=0 ps=0 
M2289 diff_2374800_2004000# diff_2374800_2004000# diff_2374800_2004000# GND efet w=2400 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2290 diff_2374800_2004000# diff_2416800_1954800# GND GND efet w=51000 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2291 Vdd diff_1892400_663600# diff_548400_1893600# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2292 diff_2143200_1873200# diff_2133600_1458000# diff_664800_1902000# GND efet w=20400 l=7200
+ ad=2.592e+08 pd=74400 as=0 ps=0 
M2293 GND diff_2118000_1905600# diff_2143200_1873200# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2294 Vdd diff_2224800_1584000# diff_664800_1902000# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2295 diff_2143200_1839600# diff_2133600_1458000# diff_664800_1825200# GND efet w=21000 l=7800
+ ad=2.6064e+08 pd=74400 as=0 ps=0 
M2296 diff_548400_1826400# diff_2082000_1496400# diff_2041200_1820400# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6208e+08 ps=74400 
M2297 diff_2118000_1820400# diff_2110800_1458000# diff_548400_1826400# GND efet w=8400 l=7200
+ ad=2.6784e+08 pd=79200 as=0 ps=0 
M2298 diff_548400_1752000# diff_2082000_1496400# diff_2041200_1761600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6784e+08 ps=76800 
M2299 diff_2118000_1764000# diff_2110800_1458000# diff_548400_1752000# GND efet w=8400 l=7200
+ ad=2.5632e+08 pd=76800 as=0 ps=0 
M2300 diff_664800_1760400# diff_2046000_1444800# diff_2052000_1734000# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2301 diff_2005200_1698000# diff_1994400_1460400# diff_664800_1683600# GND efet w=20400 l=7200
+ ad=2.592e+08 pd=76800 as=0 ps=0 
M2302 diff_548400_1684800# diff_1944000_1496400# diff_1903200_1678800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6496e+08 ps=74400 
M2303 diff_1980000_1677600# diff_1972800_1458000# diff_548400_1684800# GND efet w=8400 l=7200
+ ad=2.6496e+08 pd=79200 as=0 ps=0 
M2304 diff_548400_1610400# diff_1944000_1496400# diff_1903200_1620000# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6208e+08 ps=74400 
M2305 diff_1980000_1621200# diff_1972800_1458000# diff_548400_1610400# GND efet w=8400 l=7200
+ ad=2.5776e+08 pd=76800 as=0 ps=0 
M2306 diff_664800_1620000# diff_1908000_1442400# diff_1914000_1592400# GND efet w=21000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2307 diff_1867200_1556400# diff_1856400_1458000# diff_664800_1543200# GND efet w=20400 l=7200
+ ad=2.6064e+08 pd=76800 as=0 ps=0 
M2308 diff_548400_1543200# diff_1806000_1496400# diff_1765200_1538400# GND efet w=9600 l=7200
+ ad=0 pd=0 as=2.6784e+08 ps=74400 
M2309 diff_1843200_1536000# diff_1834800_1458000# diff_548400_1543200# GND efet w=10800 l=8400
+ ad=2.5488e+08 pd=72000 as=0 ps=0 
M2310 GND diff_1843200_1536000# diff_1867200_1556400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2311 diff_1914000_1550400# diff_1903200_1537200# GND GND efet w=22800 l=8400
+ ad=2.3328e+08 pd=72000 as=0 ps=0 
M2312 diff_664800_1543200# diff_1908000_1442400# diff_1914000_1550400# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2313 GND diff_1980000_1677600# diff_2005200_1698000# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2314 diff_2052000_1692000# diff_2041200_1678800# GND GND efet w=23400 l=7800
+ ad=2.304e+08 pd=72000 as=0 ps=0 
M2315 diff_664800_1683600# diff_2046000_1444800# diff_2052000_1692000# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2316 diff_2005200_1588800# diff_1994400_1460400# diff_664800_1620000# GND efet w=21000 l=7800
+ ad=2.592e+08 pd=74400 as=0 ps=0 
M2317 GND diff_1980000_1621200# diff_2005200_1588800# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2318 diff_2052000_1592400# diff_2041200_1620000# GND GND efet w=22800 l=8400
+ ad=2.3184e+08 pd=72000 as=0 ps=0 
M2319 GND diff_2118000_1820400# diff_2143200_1839600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2320 Vdd diff_2224800_1584000# diff_664800_1825200# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2321 Vdd diff_1892400_663600# diff_548400_1826400# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2322 Vdd diff_1892400_663600# diff_548400_1752000# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2323 diff_2143200_1730400# diff_2133600_1458000# diff_664800_1760400# GND efet w=21600 l=7200
+ ad=2.664e+08 pd=76800 as=0 ps=0 
M2324 GND diff_2118000_1764000# diff_2143200_1730400# GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2325 Vdd diff_2224800_1584000# diff_664800_1760400# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2326 GND diff_1792800_176400# diff_2077200_2900400# GND efet w=52800 l=6000
+ ad=0 pd=0 as=7.4736e+08 ps=148800 
M2327 diff_2143200_1698000# diff_2133600_1458000# diff_664800_1683600# GND efet w=21600 l=7200
+ ad=2.592e+08 pd=74400 as=0 ps=0 
M2328 diff_548400_1684800# diff_2082000_1496400# diff_2041200_1678800# GND efet w=9600 l=7200
+ ad=0 pd=0 as=2.6064e+08 ps=76800 
M2329 diff_2118000_1677600# diff_2110800_1458000# diff_548400_1684800# GND efet w=8400 l=7200
+ ad=2.6496e+08 pd=79200 as=0 ps=0 
M2330 diff_548400_1610400# diff_2082000_1496400# diff_2041200_1620000# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6208e+08 ps=76800 
M2331 diff_2118000_1621200# diff_2110800_1458000# diff_548400_1610400# GND efet w=8400 l=7200
+ ad=2.6496e+08 pd=74400 as=0 ps=0 
M2332 diff_664800_1620000# diff_2046000_1444800# diff_2052000_1592400# GND efet w=21000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2333 diff_2005200_1556400# diff_1994400_1460400# diff_664800_1543200# GND efet w=20400 l=7200
+ ad=2.4912e+08 pd=72000 as=0 ps=0 
M2334 diff_548400_1543200# diff_1944000_1496400# diff_1903200_1537200# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.6784e+08 ps=74400 
M2335 diff_1980000_1537200# diff_1972800_1458000# diff_548400_1543200# GND efet w=8400 l=7200
+ ad=2.6352e+08 pd=74400 as=0 ps=0 
M2336 GND diff_1980000_1537200# diff_2005200_1556400# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2337 diff_2052000_1551600# diff_2041200_1537200# GND GND efet w=21600 l=8400
+ ad=2.232e+08 pd=69600 as=0 ps=0 
M2338 diff_664800_1543200# diff_2046000_1444800# diff_2052000_1551600# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2339 GND diff_2118000_1677600# diff_2143200_1698000# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2340 Vdd diff_2224800_1584000# diff_664800_1683600# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2341 Vdd diff_1892400_663600# diff_548400_1684800# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2342 diff_2077200_2900400# Vdd Vdd GND efet w=10800 l=18600
+ ad=0 pd=0 as=0 ps=0 
M2343 Vdd diff_1892400_663600# diff_548400_1610400# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2344 diff_2224800_1584000# diff_2282400_1605600# diff_2224800_1584000# GND efet w=30600 l=31800
+ ad=1.47888e+09 pd=264000 as=0 ps=0 
M2345 diff_2143200_1588800# diff_2133600_1458000# diff_664800_1620000# GND efet w=21600 l=7200
+ ad=2.5632e+08 pd=74400 as=0 ps=0 
M2346 GND diff_2118000_1621200# diff_2143200_1588800# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2347 Vdd diff_2224800_1584000# diff_664800_1620000# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2348 diff_2282400_1605600# Vdd Vdd GND efet w=8400 l=7200
+ ad=2.6064e+08 pd=81600 as=0 ps=0 
M2349 diff_2282400_1605600# diff_2282400_1605600# diff_2282400_1605600# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2350 diff_2282400_1605600# diff_2282400_1605600# diff_2282400_1605600# GND efet w=2400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2351 GND diff_2342400_1538400# diff_2224800_1584000# GND efet w=74400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2352 diff_2224800_1584000# diff_2282400_1605600# Vdd GND efet w=10800 l=12000
+ ad=0 pd=0 as=0 ps=0 
M2353 diff_2224800_1584000# diff_2224800_1584000# diff_2224800_1584000# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2354 diff_2224800_1584000# diff_2224800_1584000# diff_2224800_1584000# GND efet w=4200 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2355 diff_2143200_1556400# diff_2133600_1458000# diff_664800_1543200# GND efet w=21600 l=7200
+ ad=2.5632e+08 pd=74400 as=0 ps=0 
M2356 diff_548400_1543200# diff_2082000_1496400# diff_2041200_1537200# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.4768e+08 ps=74400 
M2357 diff_2118000_1537200# diff_2110800_1458000# diff_548400_1543200# GND efet w=7200 l=8400
+ ad=2.6064e+08 pd=74400 as=0 ps=0 
M2358 GND diff_2118000_1537200# diff_2143200_1556400# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2359 Vdd diff_2224800_1584000# diff_664800_1543200# GND efet w=13800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2360 diff_2342400_1538400# Vdd Vdd GND efet w=10800 l=19200
+ ad=9.5184e+08 pd=172800 as=0 ps=0 
M2361 Vdd diff_1892400_663600# diff_548400_1543200# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2362 diff_2342400_1538400# clk1 diff_2346000_1502400# GND efet w=73200 l=7200
+ ad=0 pd=0 as=1.29024e+09 ps=266400 
M2363 GND diff_2340000_1480800# diff_2346000_1502400# GND efet w=114000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2364 GND diff_798000_1424400# diff_807600_1443600# GND efet w=18000 l=8400
+ ad=0 pd=0 as=5.4144e+08 ps=120000 
M2365 GND diff_798000_1424400# diff_843600_1497600# GND efet w=12000 l=8400
+ ad=0 pd=0 as=2.016e+08 ps=57600 
M2366 GND diff_867600_1476000# diff_872400_1458000# GND efet w=12000 l=8400
+ ad=0 pd=0 as=2.016e+08 ps=57600 
M2367 GND diff_867600_1476000# diff_894000_1458000# GND efet w=18000 l=8400
+ ad=0 pd=0 as=4.9536e+08 ps=117600 
M2368 Vdd Vdd diff_436800_1612800# GND efet w=10800 l=38400
+ ad=0 pd=0 as=1.09296e+09 ps=268800 
M2369 Vdd Vdd diff_331200_1510800# GND efet w=10800 l=42000
+ ad=0 pd=0 as=1.54368e+09 ps=348000 
M2370 diff_327600_1404000# diff_327600_1404000# diff_327600_1404000# GND efet w=3600 l=3600
+ ad=1.32912e+09 pd=280800 as=0 ps=0 
M2371 Vdd Vdd diff_327600_1404000# GND efet w=10800 l=37200
+ ad=0 pd=0 as=0 ps=0 
M2372 diff_327600_1404000# diff_327600_1404000# diff_327600_1404000# GND efet w=1800 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2373 diff_426000_1591200# diff_714000_876000# Vdd GND efet w=38400 l=7200
+ ad=-1.70585e+09 pd=439200 as=0 ps=0 
M2374 GND diff_732000_1375200# diff_426000_1591200# GND efet w=38400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2375 diff_820800_1420800# diff_810000_1159200# diff_807600_1443600# GND efet w=31800 l=10200
+ ad=5.82865e+08 pd=2.2896e+06 as=0 ps=0 
M2376 diff_843600_1497600# diff_810000_1159200# diff_844800_1435200# GND efet w=12600 l=7800
+ ad=0 pd=0 as=2.45905e+08 ps=2.0064e+06 
M2377 diff_872400_1458000# diff_867600_1452000# diff_844800_1435200# GND efet w=12600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2378 diff_894000_1458000# diff_867600_1452000# diff_820800_1420800# GND efet w=31800 l=10200
+ ad=0 pd=0 as=0 ps=0 
M2379 diff_326400_2457600# diff_326400_2457600# diff_326400_2457600# GND efet w=4200 l=4200
+ ad=1.11312e+09 pd=288000 as=0 ps=0 
M2380 Vdd Vdd diff_326400_2457600# GND efet w=10800 l=38400
+ ad=0 pd=0 as=0 ps=0 
M2381 diff_326400_2457600# diff_326400_2457600# diff_326400_2457600# GND efet w=3600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2382 GND diff_163200_1244400# diff_231600_1357200# GND efet w=39000 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2383 diff_732000_1375200# Vdd Vdd GND efet w=8400 l=38400
+ ad=4.8816e+08 pd=108000 as=0 ps=0 
M2384 GND diff_937200_1422000# diff_945600_1442400# GND efet w=18000 l=8400
+ ad=0 pd=0 as=5.1264e+08 ps=117600 
M2385 GND diff_937200_1422000# diff_981600_1458000# GND efet w=13200 l=8400
+ ad=0 pd=0 as=2.2176e+08 ps=60000 
M2386 GND diff_1005600_1476000# diff_1009200_1458000# GND efet w=13200 l=8400
+ ad=0 pd=0 as=2.016e+08 ps=57600 
M2387 GND diff_1005600_1476000# diff_1032000_1458000# GND efet w=16800 l=8400
+ ad=0 pd=0 as=4.9104e+08 ps=117600 
M2388 diff_820800_1420800# diff_946800_1120800# diff_945600_1442400# GND efet w=31800 l=10200
+ ad=0 pd=0 as=0 ps=0 
M2389 diff_981600_1458000# diff_946800_1120800# diff_844800_1435200# GND efet w=14400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2390 diff_1009200_1458000# diff_1005600_1450800# diff_844800_1435200# GND efet w=12600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2391 diff_1032000_1458000# diff_1005600_1450800# diff_820800_1420800# GND efet w=31200 l=10800
+ ad=0 pd=0 as=0 ps=0 
M2392 GND diff_1075200_1389600# diff_1082400_1443600# GND efet w=18000 l=8400
+ ad=0 pd=0 as=5.3568e+08 ps=122400 
M2393 GND diff_1075200_1389600# diff_1118400_1497600# GND efet w=12000 l=8400
+ ad=0 pd=0 as=2.016e+08 ps=57600 
M2394 GND diff_1142400_1476000# diff_1147200_1458000# GND efet w=12000 l=8400
+ ad=0 pd=0 as=2.016e+08 ps=57600 
M2395 GND diff_1142400_1476000# diff_1168800_1458000# GND efet w=18000 l=8400
+ ad=0 pd=0 as=5.1984e+08 ps=120000 
M2396 diff_820800_1420800# diff_1084800_1160400# diff_1082400_1443600# GND efet w=34200 l=10200
+ ad=0 pd=0 as=0 ps=0 
M2397 diff_1118400_1497600# diff_1084800_1160400# diff_844800_1435200# GND efet w=12600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2398 diff_1147200_1458000# diff_1142400_1450800# diff_844800_1435200# GND efet w=12600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2399 diff_1168800_1458000# diff_1142400_1450800# diff_820800_1420800# GND efet w=31800 l=10200
+ ad=0 pd=0 as=0 ps=0 
M2400 GND diff_1212000_1422000# diff_1220400_1442400# GND efet w=16800 l=8400
+ ad=0 pd=0 as=5.0544e+08 ps=117600 
M2401 GND diff_1212000_1422000# diff_1256400_1458000# GND efet w=13200 l=8400
+ ad=0 pd=0 as=2.2176e+08 ps=60000 
M2402 GND diff_1280400_1476000# diff_1284000_1458000# GND efet w=13200 l=8400
+ ad=0 pd=0 as=2.2176e+08 ps=60000 
M2403 GND diff_1280400_1476000# diff_1306800_1458000# GND efet w=16800 l=8400
+ ad=0 pd=0 as=5.0112e+08 ps=117600 
M2404 diff_820800_1420800# diff_1221600_1159200# diff_1220400_1442400# GND efet w=30600 l=10200
+ ad=0 pd=0 as=0 ps=0 
M2405 diff_1256400_1458000# diff_1221600_1159200# diff_844800_1435200# GND efet w=13800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2406 diff_1284000_1458000# diff_1280400_1450800# diff_844800_1435200# GND efet w=15000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2407 diff_1306800_1458000# diff_1280400_1450800# diff_820800_1420800# GND efet w=31200 l=10800
+ ad=0 pd=0 as=0 ps=0 
M2408 GND diff_1350000_1389600# diff_1357200_1444800# GND efet w=18000 l=8400
+ ad=0 pd=0 as=5.1984e+08 ps=120000 
M2409 GND diff_1350000_1389600# diff_1393200_1496400# GND efet w=12000 l=8400
+ ad=0 pd=0 as=2.016e+08 ps=57600 
M2410 GND diff_1417200_1476000# diff_1422000_1458000# GND efet w=12000 l=8400
+ ad=0 pd=0 as=2.016e+08 ps=57600 
M2411 GND diff_1417200_1476000# diff_1443600_1458000# GND efet w=18000 l=8400
+ ad=0 pd=0 as=5.2272e+08 ps=120000 
M2412 diff_820800_1420800# diff_1359600_1159200# diff_1357200_1444800# GND efet w=33000 l=10200
+ ad=0 pd=0 as=0 ps=0 
M2413 diff_1393200_1496400# diff_1359600_1159200# diff_844800_1435200# GND efet w=12600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2414 diff_1422000_1458000# diff_1417200_1450800# diff_844800_1435200# GND efet w=12600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2415 diff_1443600_1458000# diff_1417200_1450800# diff_820800_1420800# GND efet w=31800 l=10200
+ ad=0 pd=0 as=0 ps=0 
M2416 GND diff_1486800_1422000# diff_1495200_1443600# GND efet w=18000 l=8400
+ ad=0 pd=0 as=5.04e+08 ps=120000 
M2417 GND diff_1486800_1422000# diff_1531200_1458000# GND efet w=13200 l=7800
+ ad=0 pd=0 as=2.2176e+08 ps=60000 
M2418 GND diff_1555200_1476000# diff_1558800_1458000# GND efet w=12600 l=8400
+ ad=0 pd=0 as=2.2176e+08 ps=60000 
M2419 GND diff_1555200_1476000# diff_1581600_1458000# GND efet w=18000 l=8400
+ ad=0 pd=0 as=4.9968e+08 ps=117600 
M2420 diff_820800_1420800# diff_1497600_1159200# diff_1495200_1443600# GND efet w=31800 l=10200
+ ad=0 pd=0 as=0 ps=0 
M2421 diff_1531200_1458000# diff_1497600_1159200# diff_844800_1435200# GND efet w=13800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2422 diff_1558800_1458000# diff_1555200_1450800# diff_844800_1435200# GND efet w=13800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2423 diff_1581600_1458000# diff_1555200_1450800# diff_820800_1420800# GND efet w=32400 l=10800
+ ad=0 pd=0 as=0 ps=0 
M2424 GND diff_1624800_1396800# diff_1633200_1442400# GND efet w=18000 l=8400
+ ad=0 pd=0 as=5.0112e+08 ps=117600 
M2425 GND diff_1624800_1396800# diff_1668000_1497600# GND efet w=12600 l=7800
+ ad=0 pd=0 as=2.016e+08 ps=57600 
M2426 GND diff_1692000_1476000# diff_1696800_1458000# GND efet w=12000 l=8400
+ ad=0 pd=0 as=2.016e+08 ps=57600 
M2427 diff_1719600_1458000# diff_1692000_1476000# GND GND efet w=16800 l=8400
+ ad=5.0256e+08 pd=117600 as=0 ps=0 
M2428 diff_820800_1420800# diff_1634400_1160400# diff_1633200_1442400# GND efet w=33000 l=10200
+ ad=0 pd=0 as=0 ps=0 
M2429 diff_1668000_1497600# diff_1634400_1160400# diff_844800_1435200# GND efet w=12600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2430 diff_1696800_1458000# diff_1692000_1450800# diff_844800_1435200# GND efet w=12600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2431 diff_1719600_1458000# diff_1692000_1450800# diff_820800_1420800# GND efet w=31800 l=10200
+ ad=0 pd=0 as=0 ps=0 
M2432 GND diff_1761600_1422000# diff_1770000_1443600# GND efet w=18000 l=8400
+ ad=0 pd=0 as=5.2128e+08 ps=120000 
M2433 GND diff_1761600_1422000# diff_1806000_1496400# GND efet w=12000 l=7800
+ ad=0 pd=0 as=2.016e+08 ps=57600 
M2434 GND diff_1830000_1476000# diff_1834800_1458000# GND efet w=12000 l=8400
+ ad=0 pd=0 as=2.016e+08 ps=57600 
M2435 GND diff_1830000_1476000# diff_1856400_1458000# GND efet w=19200 l=8400
+ ad=0 pd=0 as=5.256e+08 ps=122400 
M2436 diff_820800_1420800# diff_1759200_1120800# diff_1770000_1443600# GND efet w=33000 l=10200
+ ad=0 pd=0 as=0 ps=0 
M2437 diff_1806000_1496400# diff_1759200_1120800# diff_844800_1435200# GND efet w=12600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2438 diff_1834800_1458000# diff_1820400_1143600# diff_844800_1435200# GND efet w=12600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2439 diff_1856400_1458000# diff_1820400_1143600# diff_820800_1420800# GND efet w=33000 l=10200
+ ad=0 pd=0 as=0 ps=0 
M2440 GND diff_1899600_1422000# diff_1908000_1442400# GND efet w=19800 l=7800
+ ad=0 pd=0 as=5.1264e+08 ps=127200 
M2441 GND diff_1899600_1422000# diff_1944000_1496400# GND efet w=12000 l=7200
+ ad=0 pd=0 as=2.16e+08 ps=60000 
M2442 GND diff_1968000_1476000# diff_1972800_1458000# GND efet w=13200 l=7200
+ ad=0 pd=0 as=2.1312e+08 ps=62400 
M2443 diff_1994400_1460400# diff_1968000_1476000# GND GND efet w=17400 l=7800
+ ad=5.2992e+08 pd=122400 as=0 ps=0 
M2444 diff_820800_1420800# diff_1892400_1160400# diff_1908000_1442400# GND efet w=31200 l=10800
+ ad=0 pd=0 as=0 ps=0 
M2445 diff_1944000_1496400# diff_1892400_1160400# diff_844800_1435200# GND efet w=12000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2446 diff_1972800_1458000# diff_1965600_1276800# diff_844800_1435200# GND efet w=12600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2447 diff_1994400_1460400# diff_1965600_1276800# diff_820800_1420800# GND efet w=31200 l=10200
+ ad=0 pd=0 as=0 ps=0 
M2448 GND diff_2037600_1422000# diff_2046000_1444800# GND efet w=19800 l=7200
+ ad=0 pd=0 as=5.2416e+08 ps=124800 
M2449 GND diff_2037600_1422000# diff_2082000_1496400# GND efet w=12000 l=7200
+ ad=0 pd=0 as=2.16e+08 ps=60000 
M2450 GND diff_2106000_1476000# diff_2110800_1458000# GND efet w=12000 l=7200
+ ad=0 pd=0 as=2.16e+08 ps=60000 
M2451 diff_2133600_1458000# diff_2106000_1476000# GND GND efet w=16800 l=7200
+ ad=5.2128e+08 pd=120000 as=0 ps=0 
M2452 diff_2340000_1480800# Vdd Vdd GND efet w=10800 l=27600
+ ad=9.216e+08 pd=211200 as=0 ps=0 
M2453 diff_2340000_1480800# diff_2340000_1480800# diff_2340000_1480800# GND efet w=2400 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2454 diff_2340000_1480800# diff_2340000_1480800# diff_2340000_1480800# GND efet w=2400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2455 diff_820800_1420800# diff_2011200_1227600# diff_2046000_1444800# GND efet w=33000 l=10200
+ ad=0 pd=0 as=0 ps=0 
M2456 diff_2082000_1496400# diff_2011200_1227600# diff_844800_1435200# GND efet w=12000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2457 diff_2110800_1458000# diff_2053200_1180800# diff_844800_1435200# GND efet w=12000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2458 diff_2133600_1458000# diff_2053200_1180800# diff_820800_1420800# GND efet w=31200 l=9600
+ ad=0 pd=0 as=0 ps=0 
M2459 diff_798000_1424400# diff_798000_1424400# diff_798000_1424400# GND efet w=4800 l=7200
+ ad=5.3712e+08 pd=146400 as=0 ps=0 
M2460 diff_798000_1424400# diff_798000_1424400# diff_798000_1424400# GND efet w=6000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2461 GND diff_810000_1159200# diff_798000_1424400# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2462 diff_867600_1476000# diff_867600_1452000# GND GND efet w=14400 l=7200
+ ad=5.04e+08 pd=141600 as=0 ps=0 
M2463 diff_867600_1476000# diff_867600_1476000# diff_867600_1476000# GND efet w=4800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2464 diff_867600_1476000# diff_867600_1476000# diff_867600_1476000# GND efet w=6000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2465 Vdd Vdd diff_798000_1424400# GND efet w=7200 l=38400
+ ad=0 pd=0 as=0 ps=0 
M2466 GND diff_714000_876000# diff_732000_1375200# GND efet w=19200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2467 d3 GND GND GND efet w=103200 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2468 diff_231600_1357200# diff_170400_1274400# Vdd GND efet w=38400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2469 diff_810000_1159200# diff_810000_1159200# diff_810000_1159200# GND efet w=3000 l=3000
+ ad=1.89216e+09 pd=470400 as=0 ps=0 
M2470 diff_331200_1510800# diff_516000_1338000# GND GND efet w=25200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2471 diff_326400_2457600# diff_516000_1338000# GND GND efet w=25200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2472 diff_170400_1274400# diff_163200_1244400# GND GND efet w=22800 l=7200
+ ad=1.4112e+09 pd=276000 as=0 ps=0 
M2473 diff_170400_1274400# diff_170400_1274400# diff_170400_1274400# GND efet w=2400 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2474 diff_170400_1274400# diff_170400_1274400# diff_170400_1274400# GND efet w=1800 l=5400
+ ad=0 pd=0 as=0 ps=0 
M2475 Vdd Vdd diff_170400_1274400# GND efet w=8400 l=36600
+ ad=0 pd=0 as=0 ps=0 
M2476 diff_810000_1159200# diff_810000_1159200# diff_810000_1159200# GND efet w=2400 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2477 diff_937200_1422000# diff_937200_1422000# diff_937200_1422000# GND efet w=4800 l=6000
+ ad=5.2992e+08 pd=141600 as=0 ps=0 
M2478 diff_937200_1422000# diff_937200_1422000# diff_937200_1422000# GND efet w=5400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2479 GND diff_946800_1120800# diff_937200_1422000# GND efet w=14400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2480 diff_1005600_1476000# diff_1005600_1450800# GND GND efet w=16800 l=7200
+ ad=5.1552e+08 pd=146400 as=0 ps=0 
M2481 diff_1005600_1476000# diff_1005600_1476000# diff_1005600_1476000# GND efet w=4800 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2482 diff_1005600_1476000# diff_1005600_1476000# diff_1005600_1476000# GND efet w=5400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2483 Vdd Vdd diff_867600_1476000# GND efet w=9000 l=50400
+ ad=0 pd=0 as=0 ps=0 
M2484 diff_937200_1422000# Vdd Vdd GND efet w=9000 l=45600
+ ad=0 pd=0 as=0 ps=0 
M2485 diff_867600_1452000# diff_867600_1452000# diff_867600_1452000# GND efet w=2400 l=3600
+ ad=1.95984e+09 pd=456000 as=0 ps=0 
M2486 diff_867600_1452000# diff_867600_1452000# diff_867600_1452000# GND efet w=3600 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2487 diff_946800_1120800# diff_946800_1120800# diff_946800_1120800# GND efet w=3000 l=3000
+ ad=1.76976e+09 pd=494400 as=0 ps=0 
M2488 diff_946800_1120800# diff_946800_1120800# diff_946800_1120800# GND efet w=2400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2489 diff_1075200_1389600# diff_1075200_1389600# diff_1075200_1389600# GND efet w=4800 l=7200
+ ad=5.4e+08 pd=146400 as=0 ps=0 
M2490 diff_1075200_1389600# diff_1075200_1389600# diff_1075200_1389600# GND efet w=6000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2491 GND diff_1084800_1160400# diff_1075200_1389600# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2492 diff_1142400_1476000# diff_1142400_1450800# GND GND efet w=14400 l=7200
+ ad=5.1984e+08 pd=144000 as=0 ps=0 
M2493 diff_1142400_1476000# diff_1142400_1476000# diff_1142400_1476000# GND efet w=4800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2494 diff_1212000_1422000# diff_1212000_1422000# diff_1212000_1422000# GND efet w=4800 l=7200
+ ad=5.2272e+08 pd=141600 as=0 ps=0 
M2495 diff_1142400_1476000# diff_1142400_1476000# diff_1142400_1476000# GND efet w=6000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2496 Vdd Vdd diff_1005600_1476000# GND efet w=9000 l=48000
+ ad=0 pd=0 as=0 ps=0 
M2497 diff_1075200_1389600# Vdd Vdd GND efet w=9000 l=48000
+ ad=0 pd=0 as=0 ps=0 
M2498 diff_1005600_1450800# diff_1005600_1450800# diff_1005600_1450800# GND efet w=2400 l=3000
+ ad=1.89216e+09 pd=453600 as=0 ps=0 
M2499 diff_1005600_1450800# diff_1005600_1450800# diff_1005600_1450800# GND efet w=4200 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2500 diff_1084800_1160400# diff_1084800_1160400# diff_1084800_1160400# GND efet w=3600 l=3600
+ ad=1.87488e+09 pd=470400 as=0 ps=0 
M2501 diff_1084800_1160400# diff_1084800_1160400# diff_1084800_1160400# GND efet w=2400 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2502 GND diff_1221600_1159200# diff_1212000_1422000# GND efet w=15600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2503 diff_1212000_1422000# diff_1212000_1422000# diff_1212000_1422000# GND efet w=5400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2504 diff_1280400_1476000# diff_1280400_1450800# GND GND efet w=14400 l=7200
+ ad=5.2128e+08 pd=144000 as=0 ps=0 
M2505 diff_1280400_1476000# diff_1280400_1476000# diff_1280400_1476000# GND efet w=4800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2506 diff_1280400_1476000# diff_1280400_1476000# diff_1280400_1476000# GND efet w=6000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2507 diff_1142400_1476000# Vdd Vdd GND efet w=10200 l=46800
+ ad=0 pd=0 as=0 ps=0 
M2508 diff_1212000_1422000# Vdd Vdd GND efet w=10200 l=47400
+ ad=0 pd=0 as=0 ps=0 
M2509 diff_1142400_1450800# diff_1142400_1450800# diff_1142400_1450800# GND efet w=2400 l=3600
+ ad=1.91952e+09 pd=444000 as=0 ps=0 
M2510 diff_1142400_1450800# diff_1142400_1450800# diff_1142400_1450800# GND efet w=4200 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2511 diff_1221600_1159200# diff_1221600_1159200# diff_1221600_1159200# GND efet w=3000 l=3000
+ ad=1.86192e+09 pd=472800 as=0 ps=0 
M2512 diff_1221600_1159200# diff_1221600_1159200# diff_1221600_1159200# GND efet w=3000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2513 diff_1350000_1389600# diff_1350000_1389600# diff_1350000_1389600# GND efet w=5400 l=6600
+ ad=5.328e+08 pd=151200 as=0 ps=0 
M2514 GND diff_1359600_1159200# diff_1350000_1389600# GND efet w=17400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2515 diff_1417200_1476000# diff_1417200_1450800# GND GND efet w=16800 l=7800
+ ad=5.256e+08 pd=141600 as=0 ps=0 
M2516 diff_1417200_1476000# diff_1417200_1476000# diff_1417200_1476000# GND efet w=4800 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2517 diff_1350000_1389600# diff_1350000_1389600# diff_1350000_1389600# GND efet w=5400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2518 diff_1417200_1476000# diff_1417200_1476000# diff_1417200_1476000# GND efet w=5400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2519 Vdd Vdd diff_1280400_1476000# GND efet w=9000 l=46800
+ ad=0 pd=0 as=0 ps=0 
M2520 diff_1350000_1389600# Vdd Vdd GND efet w=9000 l=45600
+ ad=0 pd=0 as=0 ps=0 
M2521 diff_1280400_1450800# diff_1280400_1450800# diff_1280400_1450800# GND efet w=2400 l=3000
+ ad=1.87632e+09 pd=448800 as=0 ps=0 
M2522 diff_1280400_1450800# diff_1280400_1450800# diff_1280400_1450800# GND efet w=4200 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2523 diff_1359600_1159200# diff_1359600_1159200# diff_1359600_1159200# GND efet w=2400 l=3600
+ ad=1.87632e+09 pd=465600 as=0 ps=0 
M2524 diff_1359600_1159200# diff_1359600_1159200# diff_1359600_1159200# GND efet w=2400 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2525 diff_1486800_1422000# diff_1486800_1422000# diff_1486800_1422000# GND efet w=4800 l=7200
+ ad=5.184e+08 pd=144000 as=0 ps=0 
M2526 GND diff_1497600_1159200# diff_1486800_1422000# GND efet w=15600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2527 diff_1555200_1476000# diff_1555200_1450800# GND GND efet w=15600 l=7200
+ ad=5.1984e+08 pd=144000 as=0 ps=0 
M2528 diff_1486800_1422000# diff_1486800_1422000# diff_1486800_1422000# GND efet w=6000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2529 diff_1555200_1476000# diff_1555200_1476000# diff_1555200_1476000# GND efet w=4800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2530 diff_1624800_1396800# diff_1624800_1396800# diff_1624800_1396800# GND efet w=4800 l=7200
+ ad=5.2848e+08 pd=146400 as=0 ps=0 
M2531 diff_1555200_1476000# diff_1555200_1476000# diff_1555200_1476000# GND efet w=5400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2532 diff_1624800_1396800# diff_1624800_1396800# diff_1624800_1396800# GND efet w=5400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2533 GND diff_1634400_1160400# diff_1624800_1396800# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2534 diff_1692000_1476000# diff_1692000_1450800# GND GND efet w=14400 l=7200
+ ad=5.2128e+08 pd=144000 as=0 ps=0 
M2535 diff_1692000_1476000# diff_1692000_1476000# diff_1692000_1476000# GND efet w=4800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2536 diff_1692000_1476000# diff_1692000_1476000# diff_1692000_1476000# GND efet w=6000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2537 Vdd Vdd diff_1417200_1476000# GND efet w=8400 l=47400
+ ad=0 pd=0 as=0 ps=0 
M2538 diff_1486800_1422000# Vdd Vdd GND efet w=9000 l=48600
+ ad=0 pd=0 as=0 ps=0 
M2539 diff_1417200_1450800# diff_1417200_1450800# diff_1417200_1450800# GND efet w=2400 l=3000
+ ad=1.93248e+09 pd=444000 as=0 ps=0 
M2540 diff_1417200_1450800# diff_1417200_1450800# diff_1417200_1450800# GND efet w=3600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2541 diff_1497600_1159200# diff_1497600_1159200# diff_1497600_1159200# GND efet w=3000 l=3000
+ ad=1.71504e+09 pd=424800 as=0 ps=0 
M2542 diff_1497600_1159200# diff_1497600_1159200# diff_1497600_1159200# GND efet w=2400 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2543 Vdd Vdd diff_1555200_1476000# GND efet w=9000 l=47400
+ ad=0 pd=0 as=0 ps=0 
M2544 diff_1624800_1396800# Vdd Vdd GND efet w=7800 l=46800
+ ad=0 pd=0 as=0 ps=0 
M2545 diff_1555200_1450800# diff_1555200_1450800# diff_1555200_1450800# GND efet w=2400 l=3000
+ ad=1.94112e+09 pd=523200 as=0 ps=0 
M2546 diff_1555200_1450800# diff_1555200_1450800# diff_1555200_1450800# GND efet w=3600 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2547 diff_1634400_1160400# diff_1634400_1160400# diff_1634400_1160400# GND efet w=3000 l=3000
+ ad=1.89792e+09 pd=477600 as=0 ps=0 
M2548 diff_1634400_1160400# diff_1634400_1160400# diff_1634400_1160400# GND efet w=2400 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2549 diff_1761600_1422000# diff_1761600_1422000# diff_1761600_1422000# GND efet w=4800 l=6000
+ ad=5.2848e+08 pd=141600 as=0 ps=0 
M2550 diff_1761600_1422000# diff_1761600_1422000# diff_1761600_1422000# GND efet w=5400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2551 GND diff_1759200_1120800# diff_1761600_1422000# GND efet w=14400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2552 diff_1830000_1476000# diff_1820400_1143600# GND GND efet w=16200 l=7800
+ ad=5.2992e+08 pd=141600 as=0 ps=0 
M2553 diff_1830000_1476000# diff_1830000_1476000# diff_1830000_1476000# GND efet w=4800 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2554 diff_1830000_1476000# diff_1830000_1476000# diff_1830000_1476000# GND efet w=5400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2555 Vdd Vdd diff_1692000_1476000# GND efet w=9000 l=46800
+ ad=0 pd=0 as=0 ps=0 
M2556 diff_1761600_1422000# Vdd Vdd GND efet w=8400 l=46200
+ ad=0 pd=0 as=0 ps=0 
M2557 diff_1692000_1450800# diff_1692000_1450800# diff_1692000_1450800# GND efet w=1800 l=4200
+ ad=2.12688e+09 pd=530400 as=0 ps=0 
M2558 diff_1692000_1450800# diff_1692000_1450800# diff_1692000_1450800# GND efet w=3600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2559 diff_1759200_1120800# diff_1759200_1120800# diff_1759200_1120800# GND efet w=3600 l=4800
+ ad=-2.08169e+09 pd=559200 as=0 ps=0 
M2560 diff_1759200_1120800# diff_1759200_1120800# diff_1759200_1120800# GND efet w=1800 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2561 diff_1899600_1422000# diff_1899600_1422000# diff_1899600_1422000# GND efet w=4800 l=7200
+ ad=5.4e+08 pd=146400 as=0 ps=0 
M2562 diff_1899600_1422000# diff_1899600_1422000# diff_1899600_1422000# GND efet w=6000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2563 GND diff_1892400_1160400# diff_1899600_1422000# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2564 diff_1968000_1476000# diff_1965600_1276800# GND GND efet w=14400 l=7200
+ ad=5.2272e+08 pd=144000 as=0 ps=0 
M2565 diff_1968000_1476000# diff_1968000_1476000# diff_1968000_1476000# GND efet w=4800 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2566 diff_2037600_1422000# diff_2037600_1422000# diff_2037600_1422000# GND efet w=4800 l=7200
+ ad=5.2272e+08 pd=144000 as=0 ps=0 
M2567 diff_1968000_1476000# diff_1968000_1476000# diff_1968000_1476000# GND efet w=5400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2568 Vdd Vdd diff_1830000_1476000# GND efet w=9000 l=47400
+ ad=0 pd=0 as=0 ps=0 
M2569 diff_1899600_1422000# Vdd Vdd GND efet w=9000 l=46800
+ ad=0 pd=0 as=0 ps=0 
M2570 diff_1820400_1143600# diff_1820400_1143600# diff_1820400_1143600# GND efet w=1800 l=2400
+ ad=-1.93625e+09 pd=609600 as=0 ps=0 
M2571 diff_1820400_1143600# diff_1820400_1143600# diff_1820400_1143600# GND efet w=3600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2572 diff_810000_1159200# diff_824400_1339200# GND GND efet w=15600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2573 diff_867600_1452000# diff_824400_1339200# GND GND efet w=16800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2574 diff_946800_1120800# diff_824400_1339200# GND GND efet w=16200 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2575 diff_1005600_1450800# diff_824400_1339200# GND GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2576 diff_1084800_1160400# diff_824400_1339200# GND GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2577 diff_1142400_1450800# diff_824400_1339200# GND GND efet w=16200 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2578 diff_1221600_1159200# diff_824400_1339200# GND GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2579 diff_1280400_1450800# diff_824400_1339200# GND GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2580 diff_1359600_1159200# diff_1302000_1048800# GND GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2581 diff_1417200_1450800# diff_1302000_1048800# GND GND efet w=16200 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2582 diff_1497600_1159200# diff_1302000_1048800# GND GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2583 diff_1555200_1450800# diff_1302000_1048800# GND GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2584 diff_1634400_1160400# diff_1302000_1048800# GND GND efet w=16800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2585 diff_1692000_1450800# diff_1302000_1048800# GND GND efet w=15600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2586 diff_1759200_1120800# diff_1302000_1048800# GND GND efet w=16800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2587 diff_1820400_1143600# diff_1302000_1048800# GND GND efet w=15600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2588 diff_2037600_1422000# diff_2037600_1422000# diff_2037600_1422000# GND efet w=6000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2589 GND diff_2011200_1227600# diff_2037600_1422000# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2590 diff_2340000_1480800# diff_268800_446400# diff_2349600_1450800# GND efet w=69000 l=6600
+ ad=0 pd=0 as=9.72e+08 ps=201600 
M2591 diff_2349600_1450800# diff_783600_224400# GND GND efet w=72000 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2592 diff_2106000_1476000# diff_2106000_1476000# diff_2106000_1476000# GND efet w=1200 l=2400
+ ad=6.048e+08 pd=194400 as=0 ps=0 
M2593 Vdd Vdd diff_1968000_1476000# GND efet w=7800 l=46200
+ ad=0 pd=0 as=0 ps=0 
M2594 diff_2037600_1422000# Vdd Vdd GND efet w=9000 l=46800
+ ad=0 pd=0 as=0 ps=0 
M2595 diff_2106000_1476000# diff_2106000_1476000# diff_2106000_1476000# GND efet w=2400 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2596 diff_820800_1420800# diff_2310000_1364400# Vdd GND efet w=38400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2597 diff_2106000_1476000# diff_2053200_1180800# GND GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2598 Vdd Vdd diff_2106000_1476000# GND efet w=6600 l=45000
+ ad=0 pd=0 as=0 ps=0 
M2599 GND diff_2335200_1249200# diff_820800_1420800# GND efet w=43800 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2600 GND diff_2335200_1249200# diff_2310000_1364400# GND efet w=40800 l=7200
+ ad=0 pd=0 as=1.5552e+09 ps=384000 
M2601 GND diff_516000_1311600# diff_327600_1404000# GND efet w=25200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2602 GND diff_516000_1311600# diff_436800_1612800# GND efet w=25200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2603 diff_523200_1467600# diff_219600_942000# Vdd GND efet w=29400 l=7200
+ ad=1.49328e+09 pd=256800 as=0 ps=0 
M2604 GND diff_732000_1252800# diff_523200_1467600# GND efet w=27600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2605 GND diff_822000_1320000# diff_810000_1159200# GND efet w=16800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2606 diff_867600_1452000# diff_822000_1320000# GND GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2607 GND diff_822000_1320000# diff_946800_1120800# GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2608 GND diff_822000_1320000# diff_1005600_1450800# GND efet w=17400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2609 GND diff_822000_1320000# diff_1359600_1159200# GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2610 diff_1417200_1450800# diff_822000_1320000# GND GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2611 GND diff_822000_1320000# diff_1497600_1159200# GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2612 diff_1555200_1450800# diff_822000_1320000# GND GND efet w=16200 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2613 diff_2053200_1180800# diff_2076000_1311600# diff_2053200_1180800# GND efet w=84000 l=3600
+ ad=2.01888e+09 pd=576000 as=0 ps=0 
M2614 diff_1084800_1160400# diff_1096800_1296000# GND GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2615 diff_1142400_1450800# diff_1096800_1296000# GND GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2616 diff_1221600_1159200# diff_1096800_1296000# GND GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2617 diff_1280400_1450800# diff_1096800_1296000# GND GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2618 diff_1634400_1160400# diff_1096800_1296000# GND GND efet w=16200 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2619 diff_1692000_1450800# diff_1096800_1296000# GND GND efet w=17400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2620 diff_1759200_1120800# diff_1096800_1296000# GND GND efet w=15600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2621 diff_1820400_1143600# diff_1096800_1296000# GND GND efet w=15600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2622 Vdd diff_2076000_1311600# diff_2053200_1180800# GND efet w=8400 l=36000
+ ad=0 pd=0 as=0 ps=0 
M2623 diff_2076000_1311600# diff_2076000_1311600# diff_2076000_1311600# GND efet w=1200 l=3600
+ ad=2.4912e+08 pd=79200 as=0 ps=0 
M2624 diff_2076000_1311600# diff_2076000_1311600# diff_2076000_1311600# GND efet w=2400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2625 Vdd Vdd diff_2076000_1311600# GND efet w=8400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2626 diff_2310000_1364400# diff_2305200_1270800# Vdd GND efet w=9600 l=19200
+ ad=0 pd=0 as=0 ps=0 
M2627 diff_1892400_1160400# diff_1902000_1294800# GND GND efet w=20400 l=7800
+ ad=1.83888e+09 pd=388800 as=0 ps=0 
M2628 diff_327600_1404000# diff_516000_1267200# GND GND efet w=25200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2629 diff_326400_2457600# diff_516000_1267200# GND GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2630 diff_170400_1274400# diff_132000_2799600# GND GND efet w=36000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2631 diff_163200_1244400# diff_163200_1244400# diff_163200_1244400# GND efet w=2400 l=7200
+ ad=1.20384e+09 pd=288000 as=0 ps=0 
M2632 diff_163200_1244400# diff_163200_1244400# diff_163200_1244400# GND efet w=2400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2633 diff_163200_1244400# d3 GND GND efet w=55200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2634 diff_732000_1252800# Vdd Vdd GND efet w=8400 l=39000
+ ad=3.7584e+08 pd=91200 as=0 ps=0 
M2635 diff_810000_1159200# diff_822000_1273200# GND GND efet w=17400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2636 diff_867600_1452000# diff_822000_1273200# GND GND efet w=15600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2637 GND diff_822000_1273200# diff_1084800_1160400# GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2638 GND diff_219600_942000# diff_732000_1252800# GND efet w=19800 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2639 diff_1142400_1450800# diff_822000_1273200# GND GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2640 diff_2053200_1180800# diff_1902000_1294800# GND GND efet w=19200 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2641 diff_2310000_1364400# diff_2305200_1270800# diff_2310000_1364400# GND efet w=54000 l=10800
+ ad=0 pd=0 as=0 ps=0 
M2642 GND diff_516000_1240800# diff_331200_1510800# GND efet w=25200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2643 GND diff_516000_1240800# diff_436800_1612800# GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2644 diff_1359600_1159200# diff_822000_1273200# GND GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2645 diff_1417200_1450800# diff_822000_1273200# GND GND efet w=17400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2646 GND diff_822000_1273200# diff_1634400_1160400# GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2647 diff_1692000_1450800# diff_822000_1273200# GND GND efet w=17400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2648 diff_2305200_1270800# diff_2305200_1270800# diff_2305200_1270800# GND efet w=3000 l=3000
+ ad=2.4624e+08 pd=79200 as=0 ps=0 
M2649 diff_2305200_1270800# diff_2305200_1270800# diff_2305200_1270800# GND efet w=1800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2650 diff_1965600_1276800# diff_1960800_1270800# GND GND efet w=31200 l=7200
+ ad=1.81008e+09 pd=484800 as=0 ps=0 
M2651 GND diff_1960800_1270800# diff_2011200_1227600# GND efet w=32400 l=7200
+ ad=0 pd=0 as=2.09808e+09 ps=501600 
M2652 diff_2305200_1270800# Vdd Vdd GND efet w=9000 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2653 GND diff_840000_1020000# diff_946800_1120800# GND efet w=15600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2654 GND diff_840000_1020000# diff_1005600_1450800# GND efet w=16800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2655 diff_1221600_1159200# diff_840000_1020000# GND GND efet w=16200 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2656 diff_1280400_1450800# diff_840000_1020000# GND GND efet w=16200 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2657 GND diff_840000_1020000# diff_1497600_1159200# GND efet w=16800 l=9600
+ ad=0 pd=0 as=0 ps=0 
M2658 diff_1555200_1450800# diff_840000_1020000# GND GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2659 diff_1759200_1120800# diff_840000_1020000# GND GND efet w=16200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2660 diff_1820400_1143600# diff_840000_1020000# GND GND efet w=15600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2661 GND diff_132000_2799600# diff_163200_1244400# GND efet w=36000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2662 diff_810000_1159200# diff_822000_1227600# GND GND efet w=15600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2663 diff_1084800_1160400# diff_822000_1227600# GND GND efet w=17400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2664 diff_946800_1120800# diff_822000_1227600# GND GND efet w=15600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2665 GND diff_822000_1227600# diff_1221600_1159200# GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2666 GND diff_1974000_1245600# diff_1965600_1276800# GND efet w=19200 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2667 GND diff_1974000_1245600# diff_2053200_1180800# GND efet w=19200 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2668 diff_2335200_1249200# Vdd Vdd GND efet w=10800 l=19200
+ ad=8.856e+08 pd=182400 as=0 ps=0 
M2669 diff_1359600_1159200# diff_822000_1227600# GND GND efet w=15600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2670 diff_1497600_1159200# diff_822000_1227600# GND GND efet w=18600 l=9600
+ ad=0 pd=0 as=0 ps=0 
M2671 diff_1634400_1160400# diff_822000_1227600# GND GND efet w=19200 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2672 Vdd Vdd Vdd GND efet w=1200 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2673 Vdd Vdd Vdd GND efet w=4200 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2674 Vdd Vdd diff_163200_1244400# GND efet w=9000 l=36600
+ ad=0 pd=0 as=0 ps=0 
M2675 diff_1005600_1450800# diff_883200_1207200# GND GND efet w=17400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2676 diff_1142400_1450800# diff_883200_1207200# GND GND efet w=18000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2677 GND diff_822000_1227600# diff_1759200_1120800# GND efet w=16200 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2678 diff_2335200_1249200# clk2 diff_2338800_1209600# GND efet w=72000 l=7200
+ ad=0 pd=0 as=1.40112e+09 ps=261600 
M2679 GND diff_2308800_1185600# diff_2338800_1209600# GND efet w=112800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2680 diff_1892400_1160400# diff_1888800_1220400# GND GND efet w=32400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2681 diff_2011200_1227600# diff_1888800_1220400# GND GND efet w=32400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2682 diff_1555200_1450800# diff_883200_1207200# GND GND efet w=16800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2683 GND diff_883200_1207200# diff_867600_1452000# GND efet w=15600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2684 GND diff_883200_1207200# diff_1280400_1450800# GND efet w=15600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2685 GND diff_883200_1207200# diff_1417200_1450800# GND efet w=16200 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2686 diff_1692000_1450800# diff_883200_1207200# GND GND efet w=16200 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2687 diff_1820400_1143600# diff_883200_1207200# GND GND efet w=15600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2688 diff_87600_2288400# diff_219600_1101600# GND GND efet w=66000 l=7200
+ ad=1.4256e+09 pd=175200 as=0 ps=0 
M2689 Vdd diff_248400_1088400# diff_87600_2288400# GND efet w=69600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2690 diff_516000_1311600# diff_516000_1338000# GND GND efet w=19200 l=7200
+ ad=8.2656e+08 pd=144000 as=0 ps=0 
M2691 Vdd Vdd diff_516000_1311600# GND efet w=11400 l=47400
+ ad=0 pd=0 as=0 ps=0 
M2692 diff_516000_1311600# diff_566400_924000# diff_574800_1088400# GND efet w=8400 l=7200
+ ad=0 pd=0 as=6.6528e+08 ps=163200 
M2693 diff_810000_1159200# diff_808800_1118400# diff_810000_1159200# GND efet w=32400 l=48000
+ ad=0 pd=0 as=0 ps=0 
M2694 diff_219600_1101600# diff_219600_1101600# diff_219600_1101600# GND efet w=2400 l=7200
+ ad=1.9872e+08 pd=62400 as=0 ps=0 
M2695 diff_219600_1101600# diff_219600_1101600# diff_219600_1101600# GND efet w=1200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2696 diff_248400_1088400# diff_248400_1088400# diff_248400_1088400# GND efet w=2400 l=5400
+ ad=2.088e+08 pd=67200 as=0 ps=0 
M2697 diff_248400_1088400# diff_248400_1088400# diff_248400_1088400# GND efet w=2400 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2698 diff_349200_1096800# diff_202800_511200# Vdd GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2699 diff_516000_1338000# diff_574800_1088400# GND GND efet w=32400 l=7200
+ ad=1.14336e+09 pd=230400 as=0 ps=0 
M2700 Vdd Vdd diff_516000_1338000# GND efet w=10800 l=46800
+ ad=0 pd=0 as=0 ps=0 
M2701 diff_867600_1452000# diff_870000_1102800# diff_867600_1452000# GND efet w=31200 l=49200
+ ad=0 pd=0 as=0 ps=0 
M2702 diff_219600_1101600# diff_222000_1082400# diff_224400_1065600# GND efet w=15000 l=6600
+ ad=0 pd=0 as=1.08288e+09 ps=211200 
M2703 diff_248400_1088400# diff_222000_1082400# diff_219600_991200# GND efet w=14400 l=8400
+ ad=0 pd=0 as=8.1648e+08 ps=182400 
M2704 diff_574800_1088400# diff_561600_1051200# diff_349200_1096800# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2705 diff_574800_1088400# diff_574800_1088400# diff_574800_1088400# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2706 diff_574800_1088400# diff_574800_1088400# diff_574800_1088400# GND efet w=1800 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2707 diff_808800_1118400# diff_808800_1118400# diff_808800_1118400# GND efet w=3000 l=3000
+ ad=1.9296e+08 pd=69600 as=0 ps=0 
M2708 diff_808800_1118400# diff_808800_1118400# diff_808800_1118400# GND efet w=1800 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2709 diff_810000_1159200# diff_808800_1118400# Vdd GND efet w=8400 l=37200
+ ad=0 pd=0 as=0 ps=0 
M2710 diff_867600_1452000# diff_870000_1102800# Vdd GND efet w=8400 l=37200
+ ad=0 pd=0 as=0 ps=0 
M2711 diff_870000_1102800# diff_870000_1102800# diff_870000_1102800# GND efet w=3000 l=3000
+ ad=1.9584e+08 pd=69600 as=0 ps=0 
M2712 diff_808800_1118400# Vdd Vdd GND efet w=7200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2713 diff_224400_1065600# diff_219600_991200# GND GND efet w=50400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2714 diff_252000_2766000# diff_202800_511200# Vdd GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2715 diff_574800_1065600# diff_561600_1051200# diff_252000_2766000# GND efet w=13200 l=7200
+ ad=6.2784e+08 pd=163200 as=0 ps=0 
M2716 diff_574800_1065600# diff_574800_1065600# diff_574800_1065600# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2717 diff_574800_1065600# diff_574800_1065600# diff_574800_1065600# GND efet w=2400 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2718 diff_870000_1102800# diff_870000_1102800# diff_870000_1102800# GND efet w=1800 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2719 diff_870000_1102800# Vdd Vdd GND efet w=8400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2720 Vdd Vdd diff_840000_1020000# GND efet w=10200 l=28800
+ ad=0 pd=0 as=-2.04137e+09 ps=633600 
M2721 Vdd Vdd diff_224400_1065600# GND efet w=10800 l=19200
+ ad=0 pd=0 as=0 ps=0 
M2722 diff_230400_2126400# diff_202800_511200# Vdd GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2723 diff_516000_1267200# diff_574800_1065600# GND GND efet w=32400 l=7200
+ ad=1.14336e+09 pd=225600 as=0 ps=0 
M2724 Vdd Vdd diff_516000_1267200# GND efet w=10800 l=46800
+ ad=0 pd=0 as=0 ps=0 
M2725 GND diff_824400_1027200# diff_840000_1020000# GND efet w=49800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2726 diff_946800_1120800# diff_948000_1117200# diff_946800_1120800# GND efet w=51000 l=27600
+ ad=0 pd=0 as=0 ps=0 
M2727 diff_1005600_1450800# diff_1008000_1102800# diff_1005600_1450800# GND efet w=30600 l=47400
+ ad=0 pd=0 as=0 ps=0 
M2728 diff_948000_1117200# diff_948000_1117200# diff_948000_1117200# GND efet w=3000 l=3000
+ ad=2.0304e+08 pd=76800 as=0 ps=0 
M2729 diff_948000_1117200# diff_948000_1117200# diff_948000_1117200# GND efet w=2400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2730 diff_946800_1120800# diff_948000_1117200# Vdd GND efet w=8400 l=37200
+ ad=0 pd=0 as=0 ps=0 
M2731 diff_1005600_1450800# diff_1008000_1102800# Vdd GND efet w=8400 l=37200
+ ad=0 pd=0 as=0 ps=0 
M2732 diff_1008000_1102800# diff_1008000_1102800# diff_1008000_1102800# GND efet w=3000 l=3000
+ ad=2.0592e+08 pd=76800 as=0 ps=0 
M2733 diff_1008000_1102800# diff_1008000_1102800# diff_1008000_1102800# GND efet w=2400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2734 diff_948000_1117200# Vdd Vdd GND efet w=9000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2735 diff_1008000_1102800# Vdd Vdd GND efet w=8400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2736 diff_822000_1273200# Vdd Vdd GND efet w=8400 l=31200
+ ad=1.49472e+09 pd=415200 as=0 ps=0 
M2737 diff_1084800_1160400# diff_1083600_1118400# diff_1084800_1160400# GND efet w=30600 l=48000
+ ad=0 pd=0 as=0 ps=0 
M2738 diff_1142400_1450800# diff_1144800_1102800# diff_1142400_1450800# GND efet w=31200 l=46800
+ ad=0 pd=0 as=0 ps=0 
M2739 diff_1083600_1118400# diff_1083600_1118400# diff_1083600_1118400# GND efet w=3000 l=3000
+ ad=1.9008e+08 pd=72000 as=0 ps=0 
M2740 diff_1083600_1118400# diff_1083600_1118400# diff_1083600_1118400# GND efet w=1800 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2741 diff_1084800_1160400# diff_1083600_1118400# Vdd GND efet w=8400 l=37200
+ ad=0 pd=0 as=0 ps=0 
M2742 diff_1142400_1450800# diff_1144800_1102800# Vdd GND efet w=8400 l=37200
+ ad=0 pd=0 as=0 ps=0 
M2743 diff_1144800_1102800# diff_1144800_1102800# diff_1144800_1102800# GND efet w=3000 l=3000
+ ad=1.872e+08 pd=69600 as=0 ps=0 
M2744 diff_1083600_1118400# Vdd Vdd GND efet w=8400 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2745 diff_1144800_1102800# diff_1144800_1102800# diff_1144800_1102800# GND efet w=1800 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2746 diff_1144800_1102800# Vdd Vdd GND efet w=9000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2747 diff_1221600_1159200# diff_1221600_1120800# diff_1221600_1159200# GND efet w=32400 l=33600
+ ad=0 pd=0 as=0 ps=0 
M2748 diff_1280400_1450800# diff_1281600_1104000# diff_1280400_1450800# GND efet w=31800 l=27600
+ ad=0 pd=0 as=0 ps=0 
M2749 diff_1359600_1159200# diff_1358400_1116000# diff_1359600_1159200# GND efet w=31800 l=46800
+ ad=0 pd=0 as=0 ps=0 
M2750 diff_1221600_1120800# diff_1221600_1120800# diff_1221600_1120800# GND efet w=3000 l=3000
+ ad=1.9728e+08 pd=72000 as=0 ps=0 
M2751 diff_1221600_1120800# diff_1221600_1120800# diff_1221600_1120800# GND efet w=1800 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2752 diff_1221600_1159200# diff_1221600_1120800# Vdd GND efet w=8400 l=37200
+ ad=0 pd=0 as=0 ps=0 
M2753 diff_1280400_1450800# diff_1281600_1104000# Vdd GND efet w=8400 l=37200
+ ad=0 pd=0 as=0 ps=0 
M2754 diff_1281600_1104000# diff_1281600_1104000# diff_1281600_1104000# GND efet w=3000 l=3000
+ ad=2.0304e+08 pd=72000 as=0 ps=0 
M2755 diff_1281600_1104000# diff_1281600_1104000# diff_1281600_1104000# GND efet w=1800 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2756 diff_1221600_1120800# Vdd Vdd GND efet w=8400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2757 diff_1281600_1104000# Vdd Vdd GND efet w=8400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2758 diff_1417200_1450800# diff_1419600_1102800# diff_1417200_1450800# GND efet w=31800 l=47400
+ ad=0 pd=0 as=0 ps=0 
M2759 diff_1358400_1116000# diff_1358400_1116000# diff_1358400_1116000# GND efet w=2400 l=3600
+ ad=1.8576e+08 pd=67200 as=0 ps=0 
M2760 diff_1358400_1116000# diff_1358400_1116000# diff_1358400_1116000# GND efet w=1800 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2761 diff_1359600_1159200# diff_1358400_1116000# Vdd GND efet w=8400 l=37200
+ ad=0 pd=0 as=0 ps=0 
M2762 diff_1417200_1450800# diff_1419600_1102800# Vdd GND efet w=8400 l=37200
+ ad=0 pd=0 as=0 ps=0 
M2763 GND diff_1696800_1017600# diff_1892400_1160400# GND efet w=19200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2764 GND diff_1696800_1017600# diff_1965600_1276800# GND efet w=19200 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2765 GND diff_1696800_1017600# diff_2011200_1227600# GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2766 GND diff_1696800_1017600# diff_2053200_1180800# GND efet w=19200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2767 diff_1497600_1159200# diff_1496400_1116000# diff_1497600_1159200# GND efet w=31800 l=46800
+ ad=0 pd=0 as=0 ps=0 
M2768 diff_1555200_1450800# diff_1556400_1104000# diff_1555200_1450800# GND efet w=49200 l=27600
+ ad=0 pd=0 as=0 ps=0 
M2769 diff_1419600_1102800# diff_1419600_1102800# diff_1419600_1102800# GND efet w=3000 l=3000
+ ad=1.872e+08 pd=67200 as=0 ps=0 
M2770 diff_1358400_1116000# Vdd Vdd GND efet w=7800 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2771 Vdd Vdd diff_219600_991200# GND efet w=10200 l=19800
+ ad=0 pd=0 as=0 ps=0 
M2772 diff_219600_991200# diff_219600_942000# GND GND efet w=51600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2773 diff_231600_1357200# diff_202800_511200# Vdd GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2774 Vdd Vdd diff_516000_1240800# GND efet w=9600 l=46800
+ ad=0 pd=0 as=1.02672e+09 ps=254400 
M2775 GND diff_840000_1020000# diff_822000_1273200# GND efet w=26400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2776 diff_824400_1339200# diff_1126800_975600# GND GND efet w=38400 l=8400
+ ad=1.57536e+09 pd=403200 as=0 ps=0 
M2777 Vdd Vdd diff_824400_1339200# GND efet w=8400 l=30000
+ ad=0 pd=0 as=0 ps=0 
M2778 diff_1302000_1048800# Vdd Vdd GND efet w=8400 l=31200
+ ad=1.49328e+09 pd=429600 as=0 ps=0 
M2779 diff_1419600_1102800# diff_1419600_1102800# diff_1419600_1102800# GND efet w=1800 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2780 diff_1419600_1102800# Vdd Vdd GND efet w=8400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2781 diff_1496400_1116000# diff_1496400_1116000# diff_1496400_1116000# GND efet w=3000 l=3000
+ ad=2.0736e+08 pd=74400 as=0 ps=0 
M2782 diff_1496400_1116000# diff_1496400_1116000# diff_1496400_1116000# GND efet w=2400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2783 diff_1497600_1159200# diff_1496400_1116000# Vdd GND efet w=8400 l=37200
+ ad=0 pd=0 as=0 ps=0 
M2784 diff_1555200_1450800# diff_1556400_1104000# Vdd GND efet w=8400 l=37200
+ ad=0 pd=0 as=0 ps=0 
M2785 diff_1556400_1104000# diff_1556400_1104000# diff_1556400_1104000# GND efet w=1800 l=4200
+ ad=2.0592e+08 pd=74400 as=0 ps=0 
M2786 diff_1496400_1116000# Vdd Vdd GND efet w=9600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2787 diff_1556400_1104000# diff_1556400_1104000# diff_1556400_1104000# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2788 diff_1556400_1104000# Vdd Vdd GND efet w=9600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2789 diff_1302000_1048800# diff_824400_1339200# GND GND efet w=25200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2790 diff_1096800_1296000# diff_1401600_975600# GND GND efet w=38400 l=8400
+ ad=1.59408e+09 pd=424800 as=0 ps=0 
M2791 Vdd Vdd diff_1096800_1296000# GND efet w=8400 l=31200
+ ad=0 pd=0 as=0 ps=0 
M2792 diff_822000_1320000# Vdd Vdd GND efet w=7800 l=30600
+ ad=1.3896e+09 pd=400800 as=0 ps=0 
M2793 diff_1634400_1160400# diff_1633200_1118400# diff_1634400_1160400# GND efet w=30600 l=48000
+ ad=0 pd=0 as=0 ps=0 
M2794 diff_1692000_1450800# diff_1694400_1102800# diff_1692000_1450800# GND efet w=48600 l=24600
+ ad=0 pd=0 as=0 ps=0 
M2795 diff_1633200_1118400# diff_1633200_1118400# diff_1633200_1118400# GND efet w=2400 l=3600
+ ad=1.8864e+08 pd=67200 as=0 ps=0 
M2796 diff_1633200_1118400# diff_1633200_1118400# diff_1633200_1118400# GND efet w=1800 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2797 diff_1634400_1160400# diff_1633200_1118400# Vdd GND efet w=8400 l=37200
+ ad=0 pd=0 as=0 ps=0 
M2798 diff_1692000_1450800# diff_1694400_1102800# Vdd GND efet w=8400 l=37200
+ ad=0 pd=0 as=0 ps=0 
M2799 diff_1694400_1102800# diff_1694400_1102800# diff_1694400_1102800# GND efet w=2400 l=3000
+ ad=2.016e+08 pd=74400 as=0 ps=0 
M2800 diff_1633200_1118400# Vdd Vdd GND efet w=8400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2801 diff_1694400_1102800# diff_1694400_1102800# diff_1694400_1102800# GND efet w=3000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2802 diff_1759200_1120800# diff_1766400_1093200# diff_1759200_1120800# GND efet w=48000 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2803 diff_1820400_1143600# diff_1819200_1102800# diff_1820400_1143600# GND efet w=48600 l=24600
+ ad=0 pd=0 as=0 ps=0 
M2804 diff_1766400_1093200# diff_1766400_1093200# diff_1766400_1093200# GND efet w=2400 l=3600
+ ad=2.2176e+08 pd=74400 as=0 ps=0 
M2805 diff_1766400_1093200# diff_1766400_1093200# diff_1766400_1093200# GND efet w=2400 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2806 diff_1759200_1120800# diff_1766400_1093200# Vdd GND efet w=8400 l=37200
+ ad=0 pd=0 as=0 ps=0 
M2807 diff_1820400_1143600# diff_1819200_1102800# Vdd GND efet w=8400 l=37200
+ ad=0 pd=0 as=0 ps=0 
M2808 diff_1819200_1102800# diff_1819200_1102800# diff_1819200_1102800# GND efet w=2400 l=3000
+ ad=2.0304e+08 pd=74400 as=0 ps=0 
M2809 diff_1694400_1102800# Vdd Vdd GND efet w=9000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2810 Vdd Vdd Vdd GND efet w=3600 l=9600
+ ad=0 pd=0 as=0 ps=0 
M2811 Vdd Vdd Vdd GND efet w=3600 l=9600
+ ad=0 pd=0 as=0 ps=0 
M2812 Vdd Vdd Vdd GND efet w=6600 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2813 Vdd Vdd Vdd GND efet w=3600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2814 Vdd Vdd diff_822000_1227600# GND efet w=9600 l=31200
+ ad=0 pd=0 as=5.112e+08 ps=148800 
M2815 diff_822000_1320000# diff_1096800_1296000# GND GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2816 diff_1766400_1093200# Vdd Vdd GND efet w=8400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2817 diff_1819200_1102800# diff_1819200_1102800# diff_1819200_1102800# GND efet w=3000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2818 diff_1819200_1102800# Vdd Vdd GND efet w=9000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2819 Vdd Vdd Vdd GND efet w=1800 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2820 Vdd Vdd Vdd GND efet w=3000 l=9000
+ ad=0 pd=0 as=0 ps=0 
M2821 Vdd Vdd Vdd GND efet w=1800 l=5400
+ ad=0 pd=0 as=0 ps=0 
M2822 Vdd Vdd Vdd GND efet w=6600 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2823 diff_822000_1227600# diff_822000_1227600# diff_822000_1227600# GND efet w=2400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2824 diff_822000_1227600# diff_822000_1227600# diff_822000_1227600# GND efet w=3000 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2825 Vdd Vdd diff_883200_1207200# GND efet w=8400 l=30000
+ ad=0 pd=0 as=4.7808e+08 ps=141600 
M2826 diff_1892400_1160400# diff_1890000_1120800# diff_1892400_1160400# GND efet w=31200 l=49200
+ ad=0 pd=0 as=0 ps=0 
M2827 diff_1890000_1120800# diff_1890000_1120800# diff_1890000_1120800# GND efet w=3000 l=3000
+ ad=1.9872e+08 pd=74400 as=0 ps=0 
M2828 diff_1890000_1120800# diff_1890000_1120800# diff_1890000_1120800# GND efet w=3000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2829 diff_1892400_1160400# diff_1890000_1120800# Vdd GND efet w=8400 l=37200
+ ad=0 pd=0 as=0 ps=0 
M2830 diff_1890000_1120800# Vdd Vdd GND efet w=8400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2831 diff_2308800_1185600# Vdd Vdd GND efet w=10800 l=27600
+ ad=5.1552e+08 pd=112800 as=0 ps=0 
M2832 GND diff_2328000_1167600# diff_2308800_1185600# GND efet w=39000 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2833 diff_1965600_1276800# diff_1970400_1102800# diff_1965600_1276800# GND efet w=53400 l=25800
+ ad=0 pd=0 as=0 ps=0 
M2834 diff_1965600_1276800# diff_1970400_1102800# Vdd GND efet w=8400 l=38400
+ ad=0 pd=0 as=0 ps=0 
M2835 diff_2011200_1227600# diff_2020800_1093200# diff_2011200_1227600# GND efet w=50400 l=28200
+ ad=0 pd=0 as=0 ps=0 
M2836 diff_2328000_1167600# diff_2328000_1167600# diff_2328000_1167600# GND efet w=1200 l=4800
+ ad=5.7024e+08 pd=110400 as=0 ps=0 
M2837 diff_1970400_1102800# diff_1970400_1102800# diff_1970400_1102800# GND efet w=2400 l=3600
+ ad=1.8288e+08 pd=69600 as=0 ps=0 
M2838 diff_1970400_1102800# diff_1970400_1102800# diff_1970400_1102800# GND efet w=2400 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2839 diff_1696800_1017600# Vdd Vdd GND efet w=9000 l=31800
+ ad=8.568e+08 pd=208800 as=0 ps=0 
M2840 diff_883200_1207200# diff_883200_1207200# diff_883200_1207200# GND efet w=1800 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2841 diff_883200_1207200# diff_883200_1207200# diff_883200_1207200# GND efet w=2400 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2842 diff_2020800_1093200# diff_2020800_1093200# diff_2020800_1093200# GND efet w=2400 l=3600
+ ad=1.872e+08 pd=67200 as=0 ps=0 
M2843 diff_2020800_1093200# diff_2020800_1093200# diff_2020800_1093200# GND efet w=1800 l=5400
+ ad=0 pd=0 as=0 ps=0 
M2844 diff_2011200_1227600# diff_2020800_1093200# Vdd GND efet w=8400 l=37200
+ ad=0 pd=0 as=0 ps=0 
M2845 diff_1970400_1102800# Vdd Vdd GND efet w=7200 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2846 diff_2020800_1093200# Vdd Vdd GND efet w=7200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2847 Vdd Vdd Vdd GND efet w=6600 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2848 Vdd Vdd Vdd GND efet w=3000 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2849 Vdd Vdd Vdd GND efet w=6600 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2850 diff_1974000_1245600# diff_1974000_1245600# diff_1974000_1245600# GND efet w=3600 l=6000
+ ad=1.00368e+09 pd=196800 as=0 ps=0 
M2851 Vdd Vdd Vdd GND efet w=3600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2852 Vdd Vdd diff_1974000_1245600# GND efet w=8400 l=36000
+ ad=0 pd=0 as=0 ps=0 
M2853 diff_1974000_1245600# diff_1888800_1220400# GND GND efet w=42000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2854 diff_1974000_1245600# diff_1974000_1245600# diff_1974000_1245600# GND efet w=2400 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2855 diff_1696800_1017600# diff_1696800_1017600# diff_1696800_1017600# GND efet w=1800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2856 diff_1696800_1017600# diff_1696800_1017600# diff_1696800_1017600# GND efet w=3000 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2857 diff_1902000_1294800# Vdd Vdd GND efet w=9000 l=36600
+ ad=6.4944e+08 pd=141600 as=0 ps=0 
M2858 diff_1902000_1294800# diff_1902000_1294800# diff_1902000_1294800# GND efet w=3600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2859 diff_1902000_1294800# diff_1902000_1294800# diff_1902000_1294800# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2860 diff_1696800_1017600# diff_1879200_1021200# GND GND efet w=46800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2861 diff_574800_1065600# diff_566400_924000# diff_516000_1240800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2862 diff_516000_1240800# diff_516000_1267200# GND GND efet w=19200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2863 diff_822000_1227600# diff_1696800_1017600# diff_1700400_1006800# GND efet w=49200 l=7200
+ ad=0 pd=0 as=4.7232e+08 ps=117600 
M2864 diff_883200_1207200# diff_1696800_1017600# diff_1778400_1006800# GND efet w=49200 l=7200
+ ad=0 pd=0 as=6.2928e+08 ps=160800 
M2865 GND diff_1960800_1270800# diff_1902000_1294800# GND efet w=37200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2866 diff_2328000_1167600# diff_2328000_1167600# diff_2328000_1167600# GND efet w=3600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2867 diff_2328000_1167600# Vdd Vdd GND efet w=9000 l=58200
+ ad=0 pd=0 as=0 ps=0 
M2868 diff_2395200_1130400# diff_1792800_176400# diff_2328000_1167600# GND efet w=26400 l=7200
+ ad=8.928e+08 pd=184800 as=0 ps=0 
M2869 diff_2395200_1130400# diff_880800_992400# GND GND efet w=27600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2870 GND diff_848400_968400# diff_2395200_1130400# GND efet w=30000 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2871 diff_268800_446400# clk1 diff_2436000_1012800# GND efet w=15000 l=6600
+ ad=1.08576e+09 pd=237600 as=2.5488e+08 ps=64800 
M2872 diff_1773600_999600# diff_1773600_999600# diff_1773600_999600# GND efet w=1800 l=3600
+ ad=8.5968e+08 pd=201600 as=0 ps=0 
M2873 diff_1879200_1021200# diff_1879200_1021200# diff_1879200_1021200# GND efet w=1800 l=4200
+ ad=8.928e+08 pd=201600 as=0 ps=0 
M2874 diff_1888800_1220400# diff_1888800_1220400# diff_1888800_1220400# GND efet w=1800 l=4200
+ ad=8.4672e+08 pd=194400 as=0 ps=0 
M2875 diff_1773600_999600# diff_1773600_999600# diff_1773600_999600# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2876 diff_1879200_1021200# diff_1879200_1021200# diff_1879200_1021200# GND efet w=2400 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2877 diff_1888800_1220400# diff_1888800_1220400# diff_1888800_1220400# GND efet w=2400 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2878 diff_880800_946800# diff_880800_992400# diff_824400_1027200# GND efet w=13200 l=7200
+ ad=1.56528e+09 pd=309600 as=8.2512e+08 ps=168000 
M2879 diff_1126800_975600# diff_880800_992400# diff_1155600_936000# GND efet w=14400 l=7200
+ ad=1.0224e+09 pd=208800 as=1.4616e+09 ps=312000 
M2880 diff_1700400_1006800# diff_883200_1207200# GND GND efet w=51000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2881 diff_1401600_975600# diff_880800_992400# diff_1430400_934800# GND efet w=13200 l=7200
+ ad=9.7056e+08 pd=206400 as=1.44288e+09 ps=307200 
M2882 diff_1778400_1006800# diff_1773600_999600# GND GND efet w=75600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2883 diff_824400_1027200# diff_848400_968400# diff_768000_823200# GND efet w=13200 l=7200
+ ad=0 pd=0 as=1.30032e+09 ps=333600 
M2884 diff_561600_1051200# diff_566400_924000# GND GND efet w=14400 l=7200
+ ad=4.32e+08 pd=108000 as=0 ps=0 
M2885 Vdd Vdd diff_561600_1051200# GND efet w=8400 l=58800
+ ad=0 pd=0 as=0 ps=0 
M2886 diff_1126800_975600# diff_848400_968400# diff_1042800_823200# GND efet w=13200 l=7200
+ ad=0 pd=0 as=1.31328e+09 ps=345600 
M2887 diff_1773600_999600# diff_880800_992400# diff_1784400_810000# GND efet w=14400 l=7200
+ ad=0 pd=0 as=1.5552e+09 ps=319200 
M2888 GND diff_2436000_1012800# diff_848400_968400# GND efet w=52800 l=6000
+ ad=0 pd=0 as=1.7496e+09 ps=362400 
M2889 diff_1960800_1270800# diff_1960800_1270800# diff_1960800_1270800# GND efet w=3600 l=8400
+ ad=1.044e+09 pd=220800 as=0 ps=0 
M2890 diff_1879200_1021200# diff_880800_992400# diff_1692000_622800# GND efet w=13200 l=7200
+ ad=0 pd=0 as=1.26e+09 ps=292800 
M2891 diff_1401600_975600# diff_848400_968400# diff_1323600_825600# GND efet w=13800 l=7200
+ ad=0 pd=0 as=8.856e+08 ps=256800 
M2892 diff_1042800_823200# diff_1042800_823200# diff_1042800_823200# GND efet w=3000 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2893 diff_1042800_823200# diff_1042800_823200# diff_1042800_823200# GND efet w=1200 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2894 Vdd Vdd diff_237600_862800# GND efet w=8400 l=9600
+ ad=0 pd=0 as=1.7568e+08 ps=64800 
M2895 diff_237600_862800# diff_237600_862800# diff_237600_862800# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2896 diff_237600_862800# diff_237600_862800# diff_237600_862800# GND efet w=1800 l=5400
+ ad=0 pd=0 as=0 ps=0 
M2897 Vdd diff_237600_862800# diff_222000_1082400# GND efet w=9600 l=9600
+ ad=0 pd=0 as=1.44432e+09 ps=252000 
M2898 diff_222000_1082400# diff_237600_862800# diff_222000_1082400# GND efet w=36600 l=27000
+ ad=0 pd=0 as=0 ps=0 
M2899 diff_1155600_936000# diff_1155600_936000# diff_1155600_936000# GND efet w=2400 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2900 diff_1155600_936000# diff_1155600_936000# diff_1155600_936000# GND efet w=1200 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2901 diff_1773600_999600# diff_848400_968400# diff_1598400_825600# GND efet w=13200 l=7200
+ ad=0 pd=0 as=9.2016e+08 ps=261600 
M2902 diff_1323600_825600# diff_1323600_825600# diff_1323600_825600# GND efet w=3000 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2903 diff_1323600_825600# diff_1323600_825600# diff_1323600_825600# GND efet w=1200 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2904 diff_222000_1082400# clk2 GND GND efet w=51000 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2905 Vdd Vdd diff_768000_823200# GND efet w=10800 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2906 diff_764400_816000# Vdd Vdd GND efet w=7200 l=45600
+ ad=7.3152e+08 pd=189600 as=0 ps=0 
M2907 diff_768000_823200# diff_764400_816000# GND GND efet w=33600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2908 diff_764400_816000# diff_764400_816000# diff_764400_816000# GND efet w=2400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2909 diff_764400_816000# diff_764400_816000# diff_764400_816000# GND efet w=1800 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2910 Vdd Vdd diff_838800_780000# GND efet w=8400 l=57600
+ ad=0 pd=0 as=6.2928e+08 ps=151200 
M2911 diff_775200_784800# Vdd Vdd GND efet w=7200 l=45600
+ ad=7.5888e+08 pd=180000 as=0 ps=0 
M2912 diff_775200_784800# diff_775200_784800# diff_775200_784800# GND efet w=2400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2913 diff_775200_784800# diff_775200_784800# diff_775200_784800# GND efet w=2400 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2914 GND diff_775200_784800# diff_838800_780000# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2915 GND diff_386400_644400# diff_543600_736800# GND efet w=14400 l=7200
+ ad=0 pd=0 as=8.136e+08 ps=211200 
M2916 GND diff_775200_784800# diff_764400_816000# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2917 diff_543600_736800# diff_543600_736800# diff_543600_736800# GND efet w=6600 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2918 diff_543600_736800# diff_543600_736800# diff_543600_736800# GND efet w=3600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2919 diff_768000_823200# diff_768000_823200# diff_768000_823200# GND efet w=3000 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2920 diff_768000_823200# diff_768000_823200# diff_768000_823200# GND efet w=2400 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2921 diff_838800_780000# diff_386400_644400# diff_764400_708000# GND efet w=15000 l=7800
+ ad=0 pd=0 as=4.464e+08 ps=91200 
M2922 Vdd Vdd diff_880800_946800# GND efet w=10800 l=37200
+ ad=0 pd=0 as=0 ps=0 
M2923 Vdd Vdd diff_991200_742800# GND efet w=8400 l=57600
+ ad=0 pd=0 as=4.9248e+08 ps=146400 
M2924 Vdd Vdd diff_1042800_823200# GND efet w=11400 l=24600
+ ad=0 pd=0 as=0 ps=0 
M2925 diff_880800_946800# diff_880800_946800# diff_880800_946800# GND efet w=1800 l=5400
+ ad=0 pd=0 as=0 ps=0 
M2926 GND diff_764400_816000# diff_775200_784800# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2927 diff_880800_946800# diff_880800_946800# diff_880800_946800# GND efet w=3600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2928 diff_991200_742800# diff_991200_742800# diff_991200_742800# GND efet w=1800 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2929 diff_991200_742800# diff_991200_742800# diff_991200_742800# GND efet w=3000 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2930 diff_768000_823200# diff_386400_644400# diff_862800_740400# GND efet w=14400 l=7200
+ ad=0 pd=0 as=4.4784e+08 ps=91200 
M2931 diff_764400_816000# diff_543600_736800# diff_754800_711600# GND efet w=30600 l=7800
+ ad=0 pd=0 as=6.8832e+08 ps=168000 
M2932 diff_378000_734400# clk2 sync GND efet w=8400 l=7200
+ ad=2.7936e+08 pd=79200 as=6.67927e+07 ps=1.0056e+06 
M2933 diff_378000_734400# diff_378000_734400# diff_378000_734400# GND efet w=2400 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2934 diff_378000_734400# diff_378000_734400# diff_378000_734400# GND efet w=1800 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2935 diff_396000_693600# diff_378000_734400# GND GND efet w=31200 l=7200
+ ad=6.2496e+08 pd=132000 as=0 ps=0 
M2936 Vdd Vdd diff_396000_693600# GND efet w=8400 l=57600
+ ad=0 pd=0 as=0 ps=0 
M2937 diff_543600_736800# Vdd Vdd GND efet w=9600 l=58800
+ ad=0 pd=0 as=0 ps=0 
M2938 GND diff_544800_702000# diff_543600_736800# GND efet w=13800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2939 GND diff_764400_708000# diff_754800_711600# GND efet w=51000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2940 diff_544800_702000# diff_544800_702000# diff_544800_702000# GND efet w=3000 l=3000
+ ad=4.8816e+08 pd=129600 as=0 ps=0 
M2941 diff_544800_702000# diff_544800_702000# diff_544800_702000# GND efet w=3000 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2942 diff_379200_640800# clk1 diff_396000_693600# GND efet w=9000 l=7800
+ ad=3.4848e+08 pd=91200 as=0 ps=0 
M2943 diff_544800_702000# Vdd Vdd GND efet w=6600 l=54600
+ ad=0 pd=0 as=0 ps=0 
M2944 diff_386400_644400# diff_379200_640800# GND GND efet w=20400 l=7200
+ ad=4.3488e+08 pd=108000 as=0 ps=0 
M2945 diff_544800_702000# diff_396000_693600# GND GND efet w=12000 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2946 Vdd Vdd diff_386400_644400# GND efet w=8400 l=41400
+ ad=0 pd=0 as=0 ps=0 
M2947 diff_386400_644400# clk2 diff_354000_610800# GND efet w=9000 l=6600
+ ad=0 pd=0 as=2.3184e+08 ps=67200 
M2948 GND diff_354000_610800# diff_356400_602400# GND efet w=15000 l=6600
+ ad=0 pd=0 as=6.2064e+08 ps=151200 
M2949 diff_880800_946800# diff_950400_691200# diff_966000_679200# GND efet w=13200 l=8400
+ ad=0 pd=0 as=1.07136e+09 ps=247200 
M2950 diff_775200_784800# diff_543600_736800# diff_904800_746400# GND efet w=27600 l=7200
+ ad=0 pd=0 as=7.8912e+08 ps=180000 
M2951 diff_904800_746400# diff_862800_740400# GND GND efet w=51600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2952 GND diff_991200_742800# diff_880800_946800# GND efet w=25200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2953 diff_1039200_816000# Vdd Vdd GND efet w=7200 l=45600
+ ad=7.5744e+08 pd=194400 as=0 ps=0 
M2954 diff_1042800_823200# diff_1039200_816000# GND GND efet w=33600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2955 diff_1039200_816000# diff_1039200_816000# diff_1039200_816000# GND efet w=2400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2956 diff_1039200_816000# diff_1039200_816000# diff_1039200_816000# GND efet w=2400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2957 Vdd Vdd diff_1113600_780000# GND efet w=8400 l=57600
+ ad=0 pd=0 as=6.048e+08 ps=151200 
M2958 diff_1050000_784800# Vdd Vdd GND efet w=7800 l=45000
+ ad=7.416e+08 pd=177600 as=0 ps=0 
M2959 diff_1050000_784800# diff_1050000_784800# diff_1050000_784800# GND efet w=1800 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2960 diff_1050000_784800# diff_1050000_784800# diff_1050000_784800# GND efet w=2400 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2961 GND diff_1050000_784800# diff_1113600_780000# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2962 GND diff_1050000_784800# diff_1039200_816000# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2963 diff_1042800_823200# diff_1042800_823200# diff_1042800_823200# GND efet w=2400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2964 diff_1042800_823200# diff_1042800_823200# diff_1042800_823200# GND efet w=2400 l=5400
+ ad=0 pd=0 as=0 ps=0 
M2965 diff_1113600_780000# diff_764400_816000# diff_1039200_708000# GND efet w=15000 l=9000
+ ad=0 pd=0 as=4.4064e+08 ps=91200 
M2966 diff_1430400_934800# diff_1430400_934800# diff_1430400_934800# GND efet w=2400 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2967 diff_1598400_825600# diff_1598400_825600# diff_1598400_825600# GND efet w=4200 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2968 diff_1784400_810000# diff_1784400_810000# diff_1784400_810000# GND efet w=2400 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2969 diff_1430400_934800# diff_1430400_934800# diff_1430400_934800# GND efet w=1200 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2970 diff_1598400_825600# diff_1598400_825600# diff_1598400_825600# GND efet w=1800 l=1800
+ ad=0 pd=0 as=0 ps=0 
M2971 diff_1888800_1220400# diff_880800_992400# diff_1489200_434400# GND efet w=14400 l=7200
+ ad=0 pd=0 as=1.2024e+09 ps=283200 
M2972 Vdd Vdd Vdd GND efet w=1800 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2973 diff_1960800_1270800# diff_1960800_1270800# diff_1960800_1270800# GND efet w=5400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2974 diff_1879200_1021200# diff_848400_968400# diff_1873200_825600# GND efet w=14400 l=7200
+ ad=0 pd=0 as=9.9216e+08 ps=273600 
M2975 diff_1888800_1220400# diff_848400_968400# diff_1042800_823200# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2976 diff_1784400_810000# diff_1784400_810000# diff_1784400_810000# GND efet w=1200 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2977 diff_1873200_825600# diff_1873200_825600# diff_1873200_825600# GND efet w=4200 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2978 diff_1692000_622800# diff_1692000_622800# diff_1692000_622800# GND efet w=3000 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2979 diff_1873200_825600# diff_1873200_825600# diff_1873200_825600# GND efet w=1200 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2980 diff_1692000_622800# diff_1692000_622800# diff_1692000_622800# GND efet w=1200 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2981 Vdd Vdd Vdd GND efet w=3600 l=5400
+ ad=0 pd=0 as=0 ps=0 
M2982 diff_848400_968400# Vdd Vdd GND efet w=10800 l=19200
+ ad=0 pd=0 as=0 ps=0 
M2983 diff_1960800_1270800# diff_880800_992400# diff_1585200_432000# GND efet w=13200 l=7200
+ ad=0 pd=0 as=1.2168e+09 ps=290400 
M2984 diff_1489200_434400# diff_1489200_434400# diff_1489200_434400# GND efet w=2400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2985 diff_1960800_1270800# diff_848400_968400# diff_768000_823200# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2986 diff_1155600_936000# Vdd Vdd GND efet w=10200 l=37800
+ ad=0 pd=0 as=0 ps=0 
M2987 Vdd Vdd diff_1266000_742800# GND efet w=8400 l=57600
+ ad=0 pd=0 as=4.9248e+08 ps=146400 
M2988 Vdd Vdd diff_1323600_825600# GND efet w=10800 l=37200
+ ad=0 pd=0 as=0 ps=0 
M2989 diff_1315200_762000# Vdd Vdd GND efet w=7200 l=50400
+ ad=7.4592e+08 pd=199200 as=0 ps=0 
M2990 diff_1155600_936000# diff_1155600_936000# diff_1155600_936000# GND efet w=1800 l=5400
+ ad=0 pd=0 as=0 ps=0 
M2991 GND diff_1039200_816000# diff_1050000_784800# GND efet w=15000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2992 diff_1155600_936000# diff_1155600_936000# diff_1155600_936000# GND efet w=3600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2993 diff_1266000_742800# diff_1266000_742800# diff_1266000_742800# GND efet w=1800 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2994 diff_1266000_742800# diff_1266000_742800# diff_1266000_742800# GND efet w=3000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2995 diff_1042800_823200# diff_764400_816000# diff_1137600_742800# GND efet w=15600 l=7200
+ ad=0 pd=0 as=4.4496e+08 ps=91200 
M2996 diff_1039200_816000# diff_775200_784800# diff_1027200_728400# GND efet w=29400 l=7200
+ ad=0 pd=0 as=8.0928e+08 ps=184800 
M2997 diff_966000_679200# diff_966000_679200# diff_966000_679200# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2998 diff_966000_679200# diff_966000_679200# diff_966000_679200# GND efet w=1800 l=1800
+ ad=0 pd=0 as=0 ps=0 
M2999 diff_991200_742800# diff_966000_679200# GND GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3000 GND diff_1039200_708000# diff_1027200_728400# GND efet w=58200 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3001 diff_1155600_936000# diff_950400_691200# diff_1240800_674400# GND efet w=13200 l=7800
+ ad=0 pd=0 as=1.11024e+09 ps=256800 
M3002 diff_1050000_784800# diff_775200_784800# diff_1179600_747600# GND efet w=27600 l=7200
+ ad=0 pd=0 as=7.92e+08 ps=177600 
M3003 GND diff_1137600_742800# diff_1179600_747600# GND efet w=51000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3004 GND diff_1266000_742800# diff_1155600_936000# GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3005 diff_1323600_825600# diff_1315200_762000# GND GND efet w=25200 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3006 diff_1315200_762000# diff_1315200_762000# diff_1315200_762000# GND efet w=1200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3007 diff_1315200_762000# diff_1315200_762000# diff_1315200_762000# GND efet w=3000 l=4800
+ ad=0 pd=0 as=0 ps=0 
M3008 Vdd Vdd diff_1389600_780000# GND efet w=8400 l=57600
+ ad=0 pd=0 as=5.5728e+08 ps=141600 
M3009 diff_1324800_784800# Vdd Vdd GND efet w=7200 l=45600
+ ad=7.4016e+08 pd=180000 as=0 ps=0 
M3010 diff_1324800_784800# diff_1324800_784800# diff_1324800_784800# GND efet w=1200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3011 diff_1324800_784800# diff_1324800_784800# diff_1324800_784800# GND efet w=2400 l=4800
+ ad=0 pd=0 as=0 ps=0 
M3012 GND diff_1324800_784800# diff_1389600_780000# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3013 GND diff_1324800_784800# diff_1315200_762000# GND efet w=14400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M3014 diff_1323600_825600# diff_1323600_825600# diff_1323600_825600# GND efet w=2400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3015 diff_1323600_825600# diff_1323600_825600# diff_1323600_825600# GND efet w=2400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3016 diff_1489200_434400# diff_1489200_434400# diff_1489200_434400# GND efet w=1200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3017 diff_848400_968400# diff_848400_968400# diff_848400_968400# GND efet w=1800 l=5400
+ ad=0 pd=0 as=0 ps=0 
M3018 diff_848400_968400# diff_848400_968400# diff_848400_968400# GND efet w=3600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3019 diff_1585200_432000# diff_1585200_432000# diff_1585200_432000# GND efet w=2400 l=4800
+ ad=0 pd=0 as=0 ps=0 
M3020 diff_848400_968400# clk2 diff_2436000_927600# GND efet w=14400 l=7200
+ ad=0 pd=0 as=2.5632e+08 ps=64800 
M3021 diff_1585200_432000# diff_1585200_432000# diff_1585200_432000# GND efet w=1200 l=4800
+ ad=0 pd=0 as=0 ps=0 
M3022 Vdd Vdd diff_1430400_934800# GND efet w=9600 l=37200
+ ad=0 pd=0 as=0 ps=0 
M3023 Vdd Vdd diff_1540800_742800# GND efet w=8400 l=57600
+ ad=0 pd=0 as=5.904e+08 ps=151200 
M3024 Vdd Vdd diff_1598400_825600# GND efet w=9600 l=37200
+ ad=0 pd=0 as=0 ps=0 
M3025 diff_1590000_762000# Vdd Vdd GND efet w=7200 l=45600
+ ad=7.3728e+08 pd=196800 as=0 ps=0 
M3026 GND diff_2436000_927600# diff_2187600_633600# GND efet w=25800 l=7200
+ ad=0 pd=0 as=-1.32569e+09 ps=820800 
M3027 diff_1430400_934800# diff_1430400_934800# diff_1430400_934800# GND efet w=1800 l=5400
+ ad=0 pd=0 as=0 ps=0 
M3028 GND diff_1315200_762000# diff_1324800_784800# GND efet w=15000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3029 diff_1430400_934800# diff_1430400_934800# diff_1430400_934800# GND efet w=3600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3030 diff_1540800_742800# diff_1540800_742800# diff_1540800_742800# GND efet w=1800 l=6600
+ ad=0 pd=0 as=0 ps=0 
M3031 diff_1540800_742800# diff_1540800_742800# diff_1540800_742800# GND efet w=3000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3032 diff_1389600_780000# diff_1039200_816000# diff_1314000_708000# GND efet w=13200 l=8400
+ ad=0 pd=0 as=4.3056e+08 ps=96000 
M3033 diff_1323600_825600# diff_1039200_816000# diff_1412400_741600# GND efet w=14400 l=8400
+ ad=0 pd=0 as=4.464e+08 ps=91200 
M3034 diff_1240800_674400# diff_1240800_674400# diff_1240800_674400# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3035 diff_1315200_762000# diff_1050000_784800# diff_1303200_711600# GND efet w=31800 l=7800
+ ad=0 pd=0 as=7.8768e+08 ps=184800 
M3036 diff_1240800_674400# diff_1240800_674400# diff_1240800_674400# GND efet w=1800 l=1800
+ ad=0 pd=0 as=0 ps=0 
M3037 diff_1266000_742800# diff_1240800_674400# GND GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3038 GND diff_1314000_708000# diff_1303200_711600# GND efet w=58800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3039 diff_1430400_934800# diff_950400_691200# diff_1512000_679200# GND efet w=13200 l=7800
+ ad=0 pd=0 as=1.0512e+09 ps=247200 
M3040 diff_1324800_784800# diff_1050000_784800# diff_1454400_751200# GND efet w=27600 l=8400
+ ad=0 pd=0 as=7.6752e+08 ps=180000 
M3041 diff_1454400_751200# diff_1412400_741600# GND GND efet w=50400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3042 GND diff_1540800_742800# diff_1430400_934800# GND efet w=24000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3043 GND diff_1590000_762000# diff_1598400_825600# GND efet w=24000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3044 diff_1590000_762000# diff_1590000_762000# diff_1590000_762000# GND efet w=1200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3045 diff_1590000_762000# diff_1590000_762000# diff_1590000_762000# GND efet w=2400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3046 Vdd Vdd diff_1664400_780000# GND efet w=8400 l=57600
+ ad=0 pd=0 as=5.688e+08 ps=144000 
M3047 diff_1599600_784800# Vdd Vdd GND efet w=7200 l=45600
+ ad=7.2288e+08 pd=175200 as=0 ps=0 
M3048 diff_1599600_784800# diff_1599600_784800# diff_1599600_784800# GND efet w=1800 l=6600
+ ad=0 pd=0 as=0 ps=0 
M3049 diff_1599600_784800# diff_1599600_784800# diff_1599600_784800# GND efet w=2400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3050 GND diff_1599600_784800# diff_1664400_780000# GND efet w=13800 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3051 GND diff_1599600_784800# diff_1590000_762000# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3052 diff_1598400_825600# diff_1598400_825600# diff_1598400_825600# GND efet w=2400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3053 diff_1598400_825600# diff_1598400_825600# diff_1598400_825600# GND efet w=2400 l=5400
+ ad=0 pd=0 as=0 ps=0 
M3054 diff_1664400_780000# diff_1315200_762000# diff_1588800_708000# GND efet w=13800 l=7800
+ ad=0 pd=0 as=4.1184e+08 ps=88800 
M3055 Vdd Vdd diff_1784400_810000# GND efet w=9600 l=38400
+ ad=0 pd=0 as=0 ps=0 
M3056 Vdd Vdd diff_1816800_742800# GND efet w=8400 l=57600
+ ad=0 pd=0 as=5.76e+08 ps=144000 
M3057 Vdd Vdd diff_1873200_825600# GND efet w=10800 l=37200
+ ad=0 pd=0 as=0 ps=0 
M3058 diff_1866000_762000# Vdd Vdd GND efet w=6600 l=46200
+ ad=7.3152e+08 pd=201600 as=0 ps=0 
M3059 diff_1784400_810000# diff_1784400_810000# diff_1784400_810000# GND efet w=1800 l=5400
+ ad=0 pd=0 as=0 ps=0 
M3060 diff_1784400_810000# diff_1784400_810000# diff_1784400_810000# GND efet w=3000 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3061 GND diff_1590000_762000# diff_1599600_784800# GND efet w=13800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3062 diff_1816800_742800# diff_1816800_742800# diff_1816800_742800# GND efet w=1200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3063 diff_1816800_742800# diff_1816800_742800# diff_1816800_742800# GND efet w=2400 l=4800
+ ad=0 pd=0 as=0 ps=0 
M3064 GND diff_1816800_742800# diff_1784400_810000# GND efet w=28200 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3065 diff_1598400_825600# diff_1315200_762000# diff_1688400_740400# GND efet w=13200 l=7200
+ ad=0 pd=0 as=4.1184e+08 ps=88800 
M3066 diff_1590000_762000# diff_1324800_784800# diff_1578000_711600# GND efet w=29400 l=7800
+ ad=0 pd=0 as=7.848e+08 ps=177600 
M3067 diff_1512000_679200# diff_1512000_679200# diff_1512000_679200# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3068 diff_1512000_679200# diff_1512000_679200# diff_1512000_679200# GND efet w=1800 l=1800
+ ad=0 pd=0 as=0 ps=0 
M3069 diff_966000_679200# diff_962400_673200# diff_349200_1096800# GND efet w=13200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3070 diff_1240800_674400# diff_962400_673200# diff_252000_2766000# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3071 Vdd Vdd diff_356400_602400# GND efet w=8400 l=58800
+ ad=0 pd=0 as=0 ps=0 
M3072 GND GND diff_554400_535200# GND efet w=38400 l=7800
+ ad=0 pd=0 as=1.67328e+09 ps=400800 
M3073 diff_356400_602400# clk1 diff_354000_553200# GND efet w=9000 l=6600
+ ad=0 pd=0 as=2.4624e+08 ps=91200 
M3074 GND diff_231600_1357200# diff_554400_535200# GND efet w=85200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3075 diff_354000_553200# diff_354000_553200# diff_354000_553200# GND efet w=4200 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3076 GND diff_354000_553200# diff_356400_542400# GND efet w=14400 l=6600
+ ad=0 pd=0 as=6.6672e+08 ps=158400 
M3077 diff_354000_553200# diff_354000_553200# diff_354000_553200# GND efet w=3000 l=4800
+ ad=0 pd=0 as=0 ps=0 
M3078 diff_554400_499200# Vdd diff_554400_535200# GND efet w=41400 l=7800
+ ad=-2.07449e+09 pd=501600 as=0 ps=0 
M3079 Vdd Vdd diff_356400_542400# GND efet w=8400 l=57600
+ ad=0 pd=0 as=0 ps=0 
M3080 GND diff_230400_2126400# diff_632400_480000# GND efet w=88800 l=8400
+ ad=0 pd=0 as=-1.83689e+09 ps=496800 
M3081 diff_604800_403200# diff_230400_2126400# GND GND efet w=46800 l=8400
+ ad=9.3024e+08 pd=232800 as=0 ps=0 
M3082 diff_554400_535200# diff_550800_528000# diff_554400_499200# GND efet w=54000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3083 clk1 GND GND GND efet w=105600 l=6000
+ ad=-5.42327e+08 pd=638400 as=0 ps=0 
M3084 GND diff_285600_456000# diff_268800_446400# GND efet w=50400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3085 diff_356400_542400# clk2 diff_352800_493200# GND efet w=8400 l=6000
+ ad=0 pd=0 as=2.5344e+08 ps=91200 
M3086 diff_352800_493200# diff_352800_493200# diff_352800_493200# GND efet w=3600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3087 GND diff_352800_493200# diff_356400_482400# GND efet w=14400 l=6600
+ ad=0 pd=0 as=6.0336e+08 ps=146400 
M3088 GND diff_231600_1357200# diff_550800_528000# GND efet w=40800 l=8400
+ ad=0 pd=0 as=4.968e+08 ps=120000 
M3089 diff_566400_924000# diff_566400_924000# diff_566400_924000# GND efet w=4200 l=4200
+ ad=-1.44089e+09 pd=844800 as=0 ps=0 
M3090 diff_566400_924000# diff_566400_924000# diff_566400_924000# GND efet w=3000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3091 diff_744000_516000# diff_733200_441600# GND GND efet w=14400 l=7200
+ ad=6.048e+08 pd=144000 as=0 ps=0 
M3092 diff_352800_493200# diff_352800_493200# diff_352800_493200# GND efet w=3000 l=4800
+ ad=0 pd=0 as=0 ps=0 
M3093 GND diff_307200_476400# diff_310800_465600# GND efet w=34800 l=6000
+ ad=0 pd=0 as=7.7184e+08 ps=170400 
M3094 Vdd Vdd diff_356400_482400# GND efet w=8400 l=57600
+ ad=0 pd=0 as=0 ps=0 
M3095 diff_550800_528000# Vdd Vdd GND efet w=10800 l=38400
+ ad=0 pd=0 as=0 ps=0 
M3096 GND p0 diff_632400_480000# GND efet w=41400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3097 GND p0 diff_656400_399600# GND efet w=14400 l=7200
+ ad=0 pd=0 as=5.4288e+08 ps=148800 
M3098 diff_729600_462000# diff_566400_924000# diff_744000_516000# GND efet w=13800 l=7800
+ ad=5.7168e+08 pd=148800 as=0 ps=0 
M3099 GND diff_566400_924000# diff_776400_445200# GND efet w=13800 l=9000
+ ad=0 pd=0 as=5.1984e+08 ps=132000 
M3100 diff_356400_482400# clk1 diff_307200_476400# GND efet w=15000 l=6600
+ ad=0 pd=0 as=2.232e+08 ps=60000 
M3101 diff_285600_456000# diff_285600_456000# diff_285600_456000# GND efet w=2400 l=7200
+ ad=2.4192e+08 pd=76800 as=0 ps=0 
M3102 diff_268800_446400# Vdd Vdd GND efet w=9600 l=18000
+ ad=0 pd=0 as=0 ps=0 
M3103 diff_285600_456000# diff_285600_456000# diff_285600_456000# GND efet w=3600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3104 diff_310800_465600# clk2 diff_285600_456000# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3105 diff_632400_480000# diff_604800_403200# diff_554400_499200# GND efet w=55200 l=8400
+ ad=0 pd=0 as=0 ps=0 
M3106 diff_310800_465600# Vdd Vdd GND efet w=10200 l=27000
+ ad=0 pd=0 as=0 ps=0 
M3107 diff_656400_399600# diff_656400_399600# diff_656400_399600# GND efet w=3600 l=4800
+ ad=0 pd=0 as=0 ps=0 
M3108 diff_733200_441600# diff_729600_462000# GND GND efet w=24600 l=7800
+ ad=3.4704e+08 pd=84000 as=0 ps=0 
M3109 diff_656400_399600# diff_656400_399600# diff_656400_399600# GND efet w=3000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3110 diff_776400_445200# diff_776400_445200# diff_776400_445200# GND efet w=3000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3111 diff_810000_472800# diff_776400_445200# diff_554400_499200# GND efet w=13200 l=8400
+ ad=4.4496e+08 pd=120000 as=0 ps=0 
M3112 diff_554400_499200# diff_656400_399600# diff_632400_480000# GND efet w=54000 l=8400
+ ad=0 pd=0 as=0 ps=0 
M3113 Vdd Vdd diff_338400_282000# GND efet w=9000 l=6600
+ ad=0 pd=0 as=2.5632e+08 ps=84000 
M3114 diff_202800_511200# diff_338400_282000# diff_202800_511200# GND efet w=52200 l=10800
+ ad=1.5192e+09 pd=367200 as=0 ps=0 
M3115 diff_338400_282000# diff_338400_282000# diff_338400_282000# GND efet w=3000 l=5400
+ ad=0 pd=0 as=0 ps=0 
M3116 diff_338400_282000# diff_338400_282000# diff_338400_282000# GND efet w=1200 l=4800
+ ad=0 pd=0 as=0 ps=0 
M3117 diff_202800_511200# diff_338400_282000# Vdd GND efet w=12000 l=20400
+ ad=0 pd=0 as=0 ps=0 
M3118 Vdd Vdd diff_366000_230400# GND efet w=8400 l=57600
+ ad=0 pd=0 as=3.9456e+08 ps=93600 
M3119 Vdd diff_477600_328800# diff_132000_2799600# GND efet w=20400 l=6600
+ ad=0 pd=0 as=-5.66807e+08 ps=945600 
M3120 diff_132000_2799600# diff_460800_272400# GND GND efet w=19200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3121 diff_366000_230400# clk1 diff_414000_259200# GND efet w=27600 l=8400
+ ad=0 pd=0 as=4.32e+08 ps=96000 
M3122 diff_202800_511200# diff_366000_230400# GND GND efet w=44400 l=6600
+ ad=0 pd=0 as=0 ps=0 
M3123 diff_414000_259200# diff_410400_252000# GND GND efet w=26400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3124 Vdd Vdd diff_460800_272400# GND efet w=8400 l=57600
+ ad=0 pd=0 as=3.9456e+08 ps=91200 
M3125 diff_604800_403200# Vdd Vdd GND efet w=9600 l=31200
+ ad=0 pd=0 as=0 ps=0 
M3126 Vdd Vdd diff_554400_499200# GND efet w=10800 l=39600
+ ad=0 pd=0 as=0 ps=0 
M3127 diff_656400_399600# Vdd Vdd GND efet w=8400 l=58200
+ ad=0 pd=0 as=0 ps=0 
M3128 diff_776400_445200# diff_776400_445200# diff_776400_445200# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3129 diff_1540800_742800# diff_1512000_679200# GND GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3130 GND diff_1588800_708000# diff_1578000_711600# GND efet w=57000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3131 diff_1784400_810000# diff_950400_691200# diff_1790400_692400# GND efet w=14400 l=7800
+ ad=0 pd=0 as=1.03392e+09 ps=232800 
M3132 diff_1599600_784800# diff_1324800_784800# diff_1730400_746400# GND efet w=26400 l=7200
+ ad=0 pd=0 as=7.2144e+08 ps=175200 
M3133 diff_1730400_746400# diff_1688400_740400# GND GND efet w=50400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3134 diff_1873200_825600# diff_1866000_762000# GND GND efet w=25200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3135 diff_1866000_762000# diff_1866000_762000# diff_1866000_762000# GND efet w=1800 l=6600
+ ad=0 pd=0 as=0 ps=0 
M3136 diff_1866000_762000# diff_1866000_762000# diff_1866000_762000# GND efet w=3000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3137 Vdd Vdd diff_1940400_778800# GND efet w=8400 l=57600
+ ad=0 pd=0 as=5.5584e+08 ps=141600 
M3138 diff_1874400_784800# Vdd Vdd GND efet w=7200 l=51000
+ ad=7.6752e+08 pd=189600 as=0 ps=0 
M3139 diff_1874400_784800# diff_1874400_784800# diff_1874400_784800# GND efet w=1200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3140 diff_1874400_784800# diff_1874400_784800# diff_1874400_784800# GND efet w=3000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3141 GND diff_1874400_784800# diff_1940400_778800# GND efet w=13200 l=8400
+ ad=0 pd=0 as=0 ps=0 
M3142 GND diff_1874400_784800# diff_1866000_762000# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3143 diff_1873200_825600# diff_1873200_825600# diff_1873200_825600# GND efet w=1800 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3144 diff_1873200_825600# diff_1873200_825600# diff_1873200_825600# GND efet w=3000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3145 GND diff_1866000_762000# diff_1874400_784800# GND efet w=14400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3146 diff_1940400_778800# diff_1590000_762000# diff_1864800_708000# GND efet w=13800 l=7800
+ ad=0 pd=0 as=4.1616e+08 ps=91200 
M3147 diff_1873200_825600# diff_1590000_762000# diff_1963200_744000# GND efet w=14400 l=7200
+ ad=0 pd=0 as=4.4352e+08 ps=91200 
M3148 diff_1866000_762000# diff_1599600_784800# diff_1852800_734400# GND efet w=26400 l=7200
+ ad=0 pd=0 as=8.0496e+08 ps=180000 
M3149 diff_1790400_692400# diff_1790400_692400# diff_1790400_692400# GND efet w=3600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3150 diff_1790400_692400# diff_1790400_692400# diff_1790400_692400# GND efet w=2400 l=2400
+ ad=0 pd=0 as=0 ps=0 
M3151 diff_1816800_742800# diff_1790400_692400# GND GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3152 GND diff_1864800_708000# diff_1852800_734400# GND efet w=57600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3153 diff_1874400_784800# diff_1599600_784800# diff_2006400_746400# GND efet w=26400 l=7200
+ ad=0 pd=0 as=7.2576e+08 ps=180000 
M3154 GND diff_1963200_744000# diff_2006400_746400# GND efet w=52800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3155 diff_1790400_692400# diff_962400_673200# diff_231600_1357200# GND efet w=17400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3156 GND diff_1887600_699600# diff_1892400_663600# GND efet w=64800 l=7200
+ ad=0 pd=0 as=-1.86713e+09 ps=580800 
M3157 diff_1512000_679200# diff_962400_673200# diff_230400_2126400# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3158 diff_1892400_663600# diff_1887600_652800# diff_1892400_663600# GND efet w=43200 l=21600
+ ad=0 pd=0 as=0 ps=0 
M3159 diff_1640400_600000# Vdd Vdd GND efet w=11400 l=34800
+ ad=6.9696e+08 pd=148800 as=0 ps=0 
M3160 diff_1892400_663600# diff_1887600_652800# Vdd GND efet w=10200 l=11400
+ ad=0 pd=0 as=0 ps=0 
M3161 GND diff_733200_441600# diff_850800_457200# GND efet w=34800 l=7200
+ ad=0 pd=0 as=9.5184e+08 ps=208800 
M3162 diff_1086000_459600# diff_810000_472800# GND GND efet w=24000 l=7200
+ ad=8.2944e+08 pd=216000 as=0 ps=0 
M3163 Vdd Vdd diff_1692000_622800# GND efet w=10800 l=19200
+ ad=0 pd=0 as=0 ps=0 
M3164 diff_1887600_652800# diff_1887600_652800# diff_1887600_652800# GND efet w=1200 l=4800
+ ad=2.2032e+08 pd=74400 as=0 ps=0 
M3165 diff_1887600_652800# diff_1887600_652800# diff_1887600_652800# GND efet w=3000 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3166 diff_1737600_447600# Vdd Vdd GND efet w=10800 l=38400
+ ad=1.1232e+09 pd=292800 as=0 ps=0 
M3167 Vdd Vdd diff_1790400_450000# GND efet w=10200 l=37800
+ ad=0 pd=0 as=1.44288e+09 ps=362400 
M3168 diff_1588800_609600# diff_850800_457200# diff_230400_2126400# GND efet w=13200 l=7200
+ ad=2.0736e+08 pd=60000 as=0 ps=0 
M3169 diff_1640400_600000# diff_1640400_600000# diff_1640400_600000# GND efet w=1800 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3170 diff_1692000_622800# diff_1640400_600000# GND GND efet w=58200 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3171 diff_1692000_622800# diff_1692000_622800# diff_1692000_622800# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3172 diff_1737600_447600# diff_1692000_622800# GND GND efet w=32400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3173 diff_1692000_622800# diff_1692000_622800# diff_1692000_622800# GND efet w=2400 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3174 diff_1640400_600000# diff_1640400_600000# diff_1640400_600000# GND efet w=1800 l=1800
+ ad=0 pd=0 as=0 ps=0 
M3175 diff_252000_2766000# diff_850800_457200# diff_1424400_518400# GND efet w=13200 l=7200
+ ad=0 pd=0 as=2.5344e+08 ps=64800 
M3176 diff_349200_1096800# diff_850800_457200# diff_1483200_518400# GND efet w=13200 l=7200
+ ad=0 pd=0 as=2.5344e+08 ps=64800 
M3177 GND diff_386400_644400# diff_810000_472800# GND efet w=15000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3178 diff_1086000_459600# diff_1086000_459600# diff_1086000_459600# GND efet w=6600 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3179 diff_1086000_459600# diff_980400_405600# GND GND efet w=14400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M3180 GND clk2 diff_1171200_489600# GND efet w=22800 l=8400
+ ad=0 pd=0 as=3.0672e+08 ps=81600 
M3181 diff_1086000_459600# diff_1086000_459600# diff_1086000_459600# GND efet w=4200 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3182 GND diff_1086000_459600# diff_1118400_457200# GND efet w=13800 l=7800
+ ad=0 pd=0 as=2.592e+08 ps=69600 
M3183 diff_1171200_489600# diff_661200_249600# diff_1171200_472800# GND efet w=30600 l=7800
+ ad=0 pd=0 as=2.5344e+08 ps=79200 
M3184 diff_1171200_472800# diff_1118400_457200# diff_1171200_454800# GND efet w=30000 l=8400
+ ad=0 pd=0 as=7.1424e+08 ps=156000 
M3185 diff_733200_441600# Vdd Vdd GND efet w=8400 l=57600
+ ad=0 pd=0 as=0 ps=0 
M3186 diff_744000_516000# Vdd Vdd GND efet w=8400 l=57000
+ ad=0 pd=0 as=0 ps=0 
M3187 diff_776400_445200# Vdd Vdd GND efet w=8400 l=57600
+ ad=0 pd=0 as=0 ps=0 
M3188 diff_554400_499200# diff_776400_445200# diff_729600_462000# GND efet w=14400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M3189 GND diff_873600_433200# diff_850800_457200# GND efet w=33600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3190 diff_951600_416400# clk2 diff_566400_924000# GND efet w=31200 l=8400
+ ad=4.1904e+08 pd=100800 as=0 ps=0 
M3191 diff_850800_457200# Vdd Vdd GND efet w=9600 l=28800
+ ad=0 pd=0 as=0 ps=0 
M3192 diff_566400_924000# Vdd Vdd GND efet w=8400 l=57600
+ ad=0 pd=0 as=0 ps=0 
M3193 diff_460800_272400# diff_477600_328800# GND GND efet w=14400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M3194 Vdd Vdd diff_477600_328800# GND efet w=8400 l=57600
+ ad=0 pd=0 as=9.6768e+08 ps=192000 
M3195 diff_549600_303600# Vdd Vdd GND efet w=7200 l=55200
+ ad=2.952e+08 pd=81600 as=0 ps=0 
M3196 Vdd Vdd diff_588000_249600# GND efet w=7200 l=45600
+ ad=0 pd=0 as=8.8848e+08 ps=175200 
M3197 diff_627600_302400# diff_410400_252000# Vdd GND efet w=13800 l=7800
+ ad=2.7792e+08 pd=74400 as=0 ps=0 
M3198 diff_627600_302400# clk1 diff_612000_230400# GND efet w=8400 l=7200
+ ad=0 pd=0 as=6.3072e+08 ps=144000 
M3199 GND diff_697200_285600# diff_549600_303600# GND efet w=12600 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3200 diff_612000_230400# diff_612000_230400# diff_612000_230400# GND efet w=4200 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3201 diff_612000_230400# diff_612000_230400# diff_612000_230400# GND efet w=2400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3202 diff_588000_249600# diff_588000_249600# diff_588000_249600# GND efet w=4200 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3203 GND diff_612000_230400# diff_588000_249600# GND efet w=42600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3204 diff_588000_249600# diff_588000_249600# diff_588000_249600# GND efet w=1800 l=9600
+ ad=0 pd=0 as=0 ps=0 
M3205 GND diff_661200_249600# diff_612000_230400# GND efet w=16200 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3206 diff_970800_408000# diff_962400_302400# diff_951600_416400# GND efet w=40200 l=9000
+ ad=3.9168e+08 pd=100800 as=0 ps=0 
M3207 GND diff_980400_405600# diff_970800_408000# GND efet w=40800 l=8400
+ ad=0 pd=0 as=0 ps=0 
M3208 diff_1086000_459600# Vdd Vdd GND efet w=8400 l=60000
+ ad=0 pd=0 as=0 ps=0 
M3209 Vdd Vdd diff_410400_252000# GND efet w=9600 l=37800
+ ad=0 pd=0 as=6.0624e+08 ps=129600 
M3210 diff_1040400_404400# diff_980400_405600# diff_873600_433200# GND efet w=31200 l=8400
+ ad=2.9952e+08 pd=81600 as=5.0976e+08 ps=112800 
M3211 diff_1057200_405600# diff_1050000_252000# diff_1040400_404400# GND efet w=30600 l=7800
+ ad=2.7648e+08 pd=81600 as=0 ps=0 
M3212 GND clk2 diff_1057200_405600# GND efet w=23400 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3213 diff_873600_433200# Vdd Vdd GND efet w=8400 l=74400
+ ad=0 pd=0 as=0 ps=0 
M3214 GND diff_783600_224400# diff_410400_252000# GND efet w=22200 l=10200
+ ad=0 pd=0 as=0 ps=0 
M3215 diff_477600_328800# diff_549600_303600# GND GND efet w=15600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3216 GND diff_588000_249600# diff_477600_328800# GND efet w=15600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3217 clk2 GND GND GND efet w=105600 l=8400
+ ad=1.02727e+09 pd=914400 as=0 ps=0 
M3218 diff_1118400_457200# Vdd Vdd GND efet w=8400 l=58800
+ ad=0 pd=0 as=0 ps=0 
M3219 Vdd Vdd diff_1171200_454800# GND efet w=8400 l=73200
+ ad=0 pd=0 as=0 ps=0 
M3220 diff_962400_673200# diff_1171200_454800# GND GND efet w=34800 l=8400
+ ad=6.0192e+08 pd=156000 as=0 ps=0 
M3221 diff_950400_691200# diff_950400_691200# diff_950400_691200# GND efet w=1800 l=5400
+ ad=8.9424e+08 pd=244800 as=0 ps=0 
M3222 diff_950400_691200# diff_950400_691200# diff_950400_691200# GND efet w=3600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3223 diff_950400_691200# diff_962400_673200# GND GND efet w=43200 l=8400
+ ad=0 pd=0 as=0 ps=0 
M3224 diff_1640400_600000# diff_1588800_609600# GND GND efet w=40800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3225 Vdd Vdd Vdd GND efet w=2400 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3226 Vdd Vdd Vdd GND efet w=1800 l=1800
+ ad=0 pd=0 as=0 ps=0 
M3227 Vdd diff_2124000_754800# diff_844800_1435200# GND efet w=22200 l=6600
+ ad=0 pd=0 as=0 ps=0 
M3228 Vdd Vdd Vdd GND efet w=1200 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3229 diff_2187600_633600# Vdd Vdd GND efet w=10800 l=37200
+ ad=0 pd=0 as=0 ps=0 
M3230 Vdd Vdd Vdd GND efet w=3000 l=4800
+ ad=0 pd=0 as=0 ps=0 
M3231 Vdd Vdd diff_2170800_822000# GND efet w=10800 l=27600
+ ad=0 pd=0 as=7.7184e+08 ps=180000 
M3232 diff_2187600_633600# clk1 diff_2418000_853200# GND efet w=14400 l=7200
+ ad=0 pd=0 as=2.4768e+08 ps=67200 
M3233 GND diff_2418000_853200# diff_1050000_252000# GND efet w=51000 l=6600
+ ad=0 pd=0 as=-2.10041e+09 ps=595200 
M3234 Vdd Vdd diff_2122800_788400# GND efet w=8400 l=7200
+ ad=0 pd=0 as=2.16e+08 ps=76800 
M3235 diff_844800_1435200# diff_2170800_822000# GND GND efet w=20400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3236 diff_2170800_822000# diff_2170800_822000# diff_2170800_822000# GND efet w=2400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3237 diff_2122800_788400# diff_2122800_788400# diff_2122800_788400# GND efet w=2400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3238 diff_2122800_788400# diff_2122800_788400# diff_2122800_788400# GND efet w=3000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3239 diff_2196000_756000# clk2 diff_2170800_822000# GND efet w=52200 l=6600
+ ad=1.30032e+09 pd=254400 as=0 ps=0 
M3240 diff_2170800_822000# diff_2170800_822000# diff_2170800_822000# GND efet w=1800 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3241 GND diff_2170800_822000# diff_2124000_754800# GND efet w=22800 l=7200
+ ad=0 pd=0 as=1.21104e+09 ps=336000 
M3242 Vdd diff_2122800_788400# diff_2124000_754800# GND efet w=9600 l=26400
+ ad=0 pd=0 as=0 ps=0 
M3243 Vdd Vdd Vdd GND efet w=2400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3244 Vdd Vdd Vdd GND efet w=3600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3245 diff_1050000_252000# Vdd Vdd GND efet w=10800 l=19200
+ ad=0 pd=0 as=0 ps=0 
M3246 GND diff_1050000_252000# diff_2196000_756000# GND efet w=72000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3247 diff_1050000_252000# diff_1050000_252000# diff_1050000_252000# GND efet w=1800 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3248 diff_1050000_252000# diff_1050000_252000# diff_1050000_252000# GND efet w=3600 l=4800
+ ad=0 pd=0 as=0 ps=0 
M3249 diff_1050000_252000# clk2 diff_2414400_778800# GND efet w=14400 l=6600
+ ad=0 pd=0 as=2.5488e+08 ps=64800 
M3250 diff_2124000_754800# diff_2122800_788400# diff_2124000_754800# GND efet w=53400 l=18600
+ ad=0 pd=0 as=0 ps=0 
M3251 GND diff_2414400_778800# diff_783600_224400# GND efet w=52200 l=6600
+ ad=0 pd=0 as=1.06992e+09 ps=230400 
M3252 Vdd Vdd Vdd GND efet w=1800 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3253 diff_2196000_756000# diff_714000_876000# GND GND efet w=46800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3254 GND diff_2106000_673200# diff_2121600_654000# GND efet w=102000 l=7200
+ ad=0 pd=0 as=1.49472e+09 ps=324000 
M3255 Vdd Vdd Vdd GND efet w=3000 l=8400
+ ad=0 pd=0 as=0 ps=0 
M3256 diff_783600_224400# Vdd Vdd GND efet w=10800 l=19200
+ ad=0 pd=0 as=0 ps=0 
M3257 diff_783600_224400# clk1 diff_2396400_704400# GND efet w=14400 l=7200
+ ad=0 pd=0 as=2.4912e+08 ps=67200 
M3258 diff_2192400_640800# diff_2035200_427200# GND GND efet w=80400 l=7200
+ ad=1.91664e+09 pd=374400 as=0 ps=0 
M3259 Vdd Vdd Vdd GND efet w=1800 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3260 GND diff_2396400_704400# diff_880800_992400# GND efet w=50400 l=7200
+ ad=0 pd=0 as=1.02672e+09 ps=220800 
M3261 Vdd Vdd Vdd GND efet w=3000 l=5400
+ ad=0 pd=0 as=0 ps=0 
M3262 diff_880800_992400# Vdd Vdd GND efet w=10800 l=19200
+ ad=0 pd=0 as=0 ps=0 
M3263 diff_2192400_640800# diff_1903200_402000# GND GND efet w=79200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3264 diff_1887600_699600# clk1 diff_2121600_654000# GND efet w=76800 l=7200
+ ad=8.8848e+08 pd=182400 as=0 ps=0 
M3265 diff_1887600_652800# Vdd Vdd GND efet w=8400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3266 diff_1790400_450000# diff_1692000_622800# GND GND efet w=30600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3267 Vdd Vdd Vdd GND efet w=4200 l=10200
+ ad=0 pd=0 as=0 ps=0 
M3268 Vdd Vdd Vdd GND efet w=6600 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3269 GND diff_1489200_434400# diff_1790400_450000# GND efet w=30600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3270 diff_1737600_447600# diff_1435200_441600# GND GND efet w=31800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3271 diff_2007600_577200# Vdd Vdd GND efet w=7800 l=7800
+ ad=2.448e+08 pd=74400 as=0 ps=0 
M3272 diff_2007600_577200# diff_2007600_577200# diff_2007600_577200# GND efet w=1200 l=4800
+ ad=0 pd=0 as=0 ps=0 
M3273 diff_2007600_577200# diff_2007600_577200# diff_2007600_577200# GND efet w=1800 l=5400
+ ad=0 pd=0 as=0 ps=0 
M3274 diff_219600_942000# diff_2007600_577200# diff_219600_942000# GND efet w=68400 l=22800
+ ad=-1.53527e+08 pd=1.0848e+06 as=0 ps=0 
M3275 diff_1887600_699600# Vdd Vdd GND efet w=9600 l=19200
+ ad=0 pd=0 as=0 ps=0 
M3276 diff_2192400_640800# diff_2187600_633600# diff_2106000_673200# GND efet w=66600 l=7800
+ ad=0 pd=0 as=7.3008e+08 ps=153600 
M3277 diff_714000_876000# diff_2082000_540000# diff_714000_876000# GND efet w=66600 l=33000
+ ad=-7.62647e+08 pd=931200 as=0 ps=0 
M3278 diff_219600_942000# diff_2007600_577200# Vdd GND efet w=9600 l=10800
+ ad=0 pd=0 as=0 ps=0 
M3279 GND diff_1585200_432000# diff_1737600_447600# GND efet w=24000 l=9600
+ ad=0 pd=0 as=0 ps=0 
M3280 GND diff_386400_644400# diff_1338000_466800# GND efet w=13800 l=7800
+ ad=0 pd=0 as=2.6928e+08 ps=67200 
M3281 diff_962400_673200# diff_962400_673200# diff_962400_673200# GND efet w=2400 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3282 diff_962400_673200# diff_962400_673200# diff_962400_673200# GND efet w=1800 l=5400
+ ad=0 pd=0 as=0 ps=0 
M3283 GND diff_1269600_462000# diff_950400_691200# GND efet w=36000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3284 diff_1608000_514800# diff_850800_457200# diff_231600_1357200# GND efet w=13200 l=7200
+ ad=2.0448e+08 pd=74400 as=0 ps=0 
M3285 diff_1608000_514800# diff_1608000_514800# diff_1608000_514800# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3286 diff_1608000_514800# diff_1608000_514800# diff_1608000_514800# GND efet w=3000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3287 diff_1338000_466800# diff_850800_457200# Vdd GND efet w=14400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3288 diff_962400_673200# Vdd Vdd GND efet w=10200 l=29400
+ ad=0 pd=0 as=0 ps=0 
M3289 diff_1384800_436800# diff_1338000_466800# GND GND efet w=63000 l=7800
+ ad=6.8688e+08 pd=160800 as=0 ps=0 
M3290 diff_950400_691200# Vdd Vdd GND efet w=10800 l=31200
+ ad=0 pd=0 as=0 ps=0 
M3291 diff_1269600_462000# diff_783600_224400# GND GND efet w=37800 l=10200
+ ad=3.4704e+08 pd=86400 as=0 ps=0 
M3292 diff_1435200_441600# diff_1424400_518400# GND GND efet w=49200 l=7200
+ ad=7.6464e+08 pd=170400 as=0 ps=0 
M3293 diff_1435200_441600# diff_1435200_441600# diff_1435200_441600# GND efet w=3600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3294 diff_1435200_441600# diff_1435200_441600# diff_1435200_441600# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3295 diff_1489200_434400# diff_1435200_441600# GND GND efet w=32400 l=8400
+ ad=0 pd=0 as=0 ps=0 
M3296 GND diff_1515600_435600# diff_1790400_450000# GND efet w=30600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3297 diff_1790400_450000# diff_1608000_514800# GND GND efet w=51000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3298 GND diff_1384800_436800# diff_1790400_450000# GND efet w=24600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3299 Vdd Vdd diff_2082000_540000# GND efet w=7800 l=7800
+ ad=0 pd=0 as=2.3904e+08 ps=79200 
M3300 diff_2106000_673200# Vdd Vdd GND efet w=10200 l=28200
+ ad=0 pd=0 as=0 ps=0 
M3301 diff_880800_992400# clk2 diff_2401200_631200# GND efet w=14400 l=6000
+ ad=0 pd=0 as=2.5344e+08 ps=64800 
M3302 GND diff_2401200_631200# diff_2035200_427200# GND efet w=41400 l=6600
+ ad=0 pd=0 as=-1.65047e+08 ps=1.1544e+06 
M3303 Vdd Vdd Vdd GND efet w=1800 l=2400
+ ad=0 pd=0 as=0 ps=0 
M3304 Vdd Vdd Vdd GND efet w=2400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3305 diff_2035200_427200# Vdd Vdd GND efet w=11400 l=28200
+ ad=0 pd=0 as=0 ps=0 
M3306 diff_2082000_540000# diff_2082000_540000# diff_2082000_540000# GND efet w=1200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3307 diff_2082000_540000# diff_2082000_540000# diff_2082000_540000# GND efet w=2400 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3308 Vdd Vdd Vdd GND efet w=5400 l=10200
+ ad=0 pd=0 as=0 ps=0 
M3309 Vdd Vdd Vdd GND efet w=3000 l=10200
+ ad=0 pd=0 as=0 ps=0 
M3310 diff_2035200_427200# clk1 diff_2378400_554400# GND efet w=13800 l=6000
+ ad=0 pd=0 as=2.2608e+08 ps=62400 
M3311 Vdd Vdd diff_2074800_2772000# GND efet w=10200 l=19200
+ ad=0 pd=0 as=-8.33207e+08 ps=835200 
M3312 Vdd diff_2082000_540000# diff_714000_876000# GND efet w=9600 l=19200
+ ad=0 pd=0 as=0 ps=0 
M3313 diff_219600_942000# diff_1974000_518400# GND GND efet w=75600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3314 diff_714000_876000# diff_1974000_518400# GND GND efet w=46200 l=6600
+ ad=0 pd=0 as=0 ps=0 
M3315 Vdd Vdd diff_2071200_496800# GND efet w=9600 l=27600
+ ad=0 pd=0 as=6.048e+08 ps=146400 
M3316 GND diff_2378400_554400# diff_962400_302400# GND efet w=53400 l=6600
+ ad=0 pd=0 as=-1.57481e+09 ps=655200 
M3317 Vdd Vdd Vdd GND efet w=3000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3318 Vdd Vdd Vdd GND efet w=3600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3319 diff_962400_302400# Vdd Vdd GND efet w=10800 l=19200
+ ad=0 pd=0 as=0 ps=0 
M3320 diff_2074800_2772000# diff_1974000_518400# GND GND efet w=57600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3321 diff_1792800_498000# diff_1608000_514800# GND GND efet w=49200 l=7200
+ ad=1.60704e+09 pd=388800 as=0 ps=0 
M3322 GND diff_1870800_396000# diff_219600_942000# GND efet w=72000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3323 GND diff_2071200_496800# diff_714000_876000# GND efet w=43200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3324 diff_1489200_434400# diff_1489200_434400# diff_1489200_434400# GND efet w=2400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3325 GND diff_1483200_518400# diff_1515600_435600# GND efet w=45000 l=7800
+ ad=0 pd=0 as=8.6832e+08 ps=201600 
M3326 Vdd Vdd diff_1269600_462000# GND efet w=10200 l=30600
+ ad=0 pd=0 as=0 ps=0 
M3327 diff_1384800_436800# Vdd Vdd GND efet w=9600 l=28800
+ ad=0 pd=0 as=0 ps=0 
M3328 diff_1489200_434400# diff_1489200_434400# diff_1489200_434400# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3329 diff_1515600_435600# diff_1515600_435600# diff_1515600_435600# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3330 diff_1435200_441600# Vdd Vdd GND efet w=9600 l=38400
+ ad=0 pd=0 as=0 ps=0 
M3331 diff_1585200_432000# diff_1515600_435600# GND GND efet w=33600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M3332 GND diff_1608000_514800# diff_1626000_416400# GND efet w=45600 l=7200
+ ad=0 pd=0 as=7.2e+08 ps=172800 
M3333 diff_1585200_432000# diff_1585200_432000# diff_1585200_432000# GND efet w=1800 l=5400
+ ad=0 pd=0 as=0 ps=0 
M3334 diff_1515600_435600# diff_1515600_435600# diff_1515600_435600# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3335 diff_1585200_432000# diff_1585200_432000# diff_1585200_432000# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3336 diff_697200_285600# diff_1626000_416400# GND GND efet w=25200 l=7200
+ ad=1.13472e+09 pd=278400 as=0 ps=0 
M3337 GND diff_1384800_436800# diff_697200_285600# GND efet w=33000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3338 diff_697200_285600# diff_1737600_447600# GND GND efet w=25200 l=8400
+ ad=0 pd=0 as=0 ps=0 
M3339 GND diff_1384800_436800# diff_1792800_498000# GND efet w=31200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3340 diff_1792800_498000# diff_1790400_450000# GND GND efet w=31800 l=10200
+ ad=0 pd=0 as=0 ps=0 
M3341 diff_697200_285600# diff_697200_285600# diff_697200_285600# GND efet w=2400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3342 diff_1626000_416400# diff_1626000_416400# diff_1626000_416400# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3343 diff_697200_285600# diff_697200_285600# diff_697200_285600# GND efet w=2400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3344 diff_1489200_434400# Vdd Vdd GND efet w=10800 l=28800
+ ad=0 pd=0 as=0 ps=0 
M3345 diff_1626000_416400# diff_1626000_416400# diff_1626000_416400# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3346 diff_1585200_432000# Vdd Vdd GND efet w=10200 l=31200
+ ad=0 pd=0 as=0 ps=0 
M3347 Vdd Vdd diff_1626000_416400# GND efet w=10800 l=39600
+ ad=0 pd=0 as=0 ps=0 
M3348 Vdd Vdd diff_1515600_435600# GND efet w=9600 l=39600
+ ad=0 pd=0 as=0 ps=0 
M3349 diff_697200_285600# Vdd Vdd GND efet w=9600 l=38400
+ ad=0 pd=0 as=0 ps=0 
M3350 GND diff_2071200_496800# diff_2074800_2772000# GND efet w=54000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3351 diff_1974000_518400# diff_1792800_176400# GND GND efet w=31200 l=7200
+ ad=6.336e+08 pd=158400 as=0 ps=0 
M3352 GND diff_2035200_427200# diff_219600_942000# GND efet w=59400 l=11400
+ ad=0 pd=0 as=0 ps=0 
M3353 diff_714000_876000# diff_1903200_402000# GND GND efet w=44400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3354 GND diff_1737600_447600# diff_1792800_498000# GND efet w=25800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3355 GND diff_1792800_498000# diff_1903200_402000# GND efet w=21600 l=7200
+ ad=0 pd=0 as=4.7232e+08 ps=100800 
M3356 GND diff_962400_302400# diff_2071200_496800# GND efet w=38400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3357 diff_2074800_2772000# diff_1951200_409200# GND GND efet w=57000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3358 GND diff_1790400_450000# diff_1951200_409200# GND efet w=21600 l=7200
+ ad=0 pd=0 as=4.0608e+08 ps=98400 
M3359 diff_1792800_498000# Vdd Vdd GND efet w=9600 l=37200
+ ad=0 pd=0 as=0 ps=0 
M3360 diff_1870800_396000# diff_697200_285600# GND GND efet w=20400 l=8400
+ ad=5.0544e+08 pd=96000 as=0 ps=0 
M3361 Vdd Vdd diff_1870800_396000# GND efet w=10800 l=50400
+ ad=0 pd=0 as=0 ps=0 
M3362 Vdd Vdd diff_1903200_402000# GND efet w=10800 l=46800
+ ad=0 pd=0 as=0 ps=0 
M3363 diff_1951200_409200# Vdd Vdd GND efet w=10800 l=46800
+ ad=0 pd=0 as=0 ps=0 
M3364 diff_1974000_518400# Vdd Vdd GND efet w=7200 l=23400
+ ad=0 pd=0 as=0 ps=0 
M3365 diff_962400_302400# clk2 diff_2383200_470400# GND efet w=14400 l=6000
+ ad=0 pd=0 as=2.4048e+08 ps=62400 
M3366 Vdd Vdd Vdd GND efet w=1800 l=2400
+ ad=0 pd=0 as=0 ps=0 
M3367 diff_2359200_448800# Vdd Vdd GND efet w=11400 l=55800
+ ad=7.0848e+08 pd=163200 as=0 ps=0 
M3368 GND diff_2383200_470400# diff_2359200_448800# GND efet w=18000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3369 Vdd Vdd Vdd GND efet w=3000 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3370 diff_2378400_421200# clk1 diff_2359200_448800# GND efet w=13200 l=7200
+ ad=2.2176e+08 pd=60000 as=0 ps=0 
M3371 GND diff_2378400_421200# diff_661200_249600# GND efet w=51000 l=6600
+ ad=0 pd=0 as=8.3664e+08 ps=175200 
M3372 Vdd Vdd Vdd GND efet w=1800 l=1800
+ ad=0 pd=0 as=0 ps=0 
M3373 Vdd Vdd Vdd GND efet w=3000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3374 Vdd Vdd Vdd GND efet w=2400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3375 Vdd Vdd Vdd GND efet w=1200 l=1800
+ ad=0 pd=0 as=0 ps=0 
M3376 diff_1792800_176400# Vdd Vdd GND efet w=10800 l=19200
+ ad=-1.66697e+09 pd=554400 as=0 ps=0 
M3377 diff_661200_249600# Vdd Vdd GND efet w=10800 l=19800
+ ad=0 pd=0 as=0 ps=0 
M3378 Vdd Vdd diff_980400_405600# GND efet w=10800 l=27600
+ ad=0 pd=0 as=7.56e+08 ps=175200 
M3379 Vdd Vdd diff_2143200_162000# GND efet w=13200 l=45000
+ ad=0 pd=0 as=8.6976e+08 ps=194400 
M3380 diff_1792800_176400# reset GND GND efet w=126000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3381 sync GND GND GND efet w=105600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M3382 reset GND GND GND efet w=108000 l=8400
+ ad=-7.61207e+08 pd=772800 as=0 ps=0 
M3383 GND GND p0 GND efet w=105600 l=8400
+ ad=0 pd=0 as=-1.18169e+09 ps=748800 
M3384 diff_2143200_162000# diff_2143200_162000# diff_2143200_162000# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3385 diff_2143200_162000# diff_2143200_162000# diff_2143200_162000# GND efet w=1800 l=5400
+ ad=0 pd=0 as=0 ps=0 
M3386 diff_980400_405600# diff_2143200_162000# GND GND efet w=38400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3387 GND cm diff_2143200_162000# GND efet w=50400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3388 cm GND GND GND efet w=106200 l=7800
+ ad=-9.18167e+08 pd=777600 as=0 ps=0 
C0 metal_2412000_40800# gnd! 43.2fF ;**FLOATING
C1 metal_2356800_49200# gnd! 46.1fF ;**FLOATING
C2 metal_2301600_51600# gnd! 48.2fF ;**FLOATING
C3 metal_2246400_62400# gnd! 42.4fF ;**FLOATING
C4 metal_696000_55200# gnd! 6.8fF ;**FLOATING
C5 metal_675600_63600# gnd! 3.8fF ;**FLOATING
C6 metal_660000_76800# gnd! 10.7fF ;**FLOATING
C7 metal_674400_76800# gnd! 26.5fF ;**FLOATING
C8 metal_717600_111600# gnd! 75.9fF ;**FLOATING
C9 metal_156000_162000# gnd! 8.7fF ;**FLOATING
C10 metal_2354400_2950800# gnd! 54.0fF ;**FLOATING
C11 diff_2143200_162000# gnd! 133.4fF
C12 cm gnd! 631.9fF
C13 reset gnd! 831.6fF
C14 diff_2378400_421200# gnd! 73.6fF
C15 diff_2359200_448800# gnd! 87.0fF
C16 diff_2383200_470400# gnd! 63.2fF
C17 diff_1951200_409200# gnd! 186.0fF
C18 diff_1626000_416400# gnd! 139.4fF
C19 diff_1870800_396000# gnd! 167.8fF
C20 diff_1792800_498000# gnd! 307.7fF
C21 diff_2071200_496800# gnd! 140.2fF
C22 diff_1974000_518400# gnd! 192.1fF
C23 diff_2378400_554400# gnd! 70.5fF
C24 diff_2401200_631200# gnd! 68.0fF
C25 diff_1338000_466800# gnd! 103.6fF
C26 diff_1269600_462000# gnd! 97.5fF
C27 diff_1384800_436800# gnd! 343.5fF
C28 diff_1608000_514800# gnd! 211.7fF
C29 diff_1515600_435600# gnd! 281.0fF
C30 diff_2082000_540000# gnd! 127.9fF
C31 diff_1435200_441600# gnd! 278.3fF
C32 diff_2007600_577200# gnd! 120.2fF
C33 diff_1903200_402000# gnd! 324.5fF
C34 diff_2396400_704400# gnd! 74.3fF
C35 diff_2035200_427200# gnd! 844.3fF
C36 diff_2192400_640800# gnd! 254.1fF
C37 diff_2121600_654000# gnd! 181.9fF
C38 diff_2106000_673200# gnd! 178.8fF
C39 diff_2414400_778800# gnd! 73.0fF
C40 diff_2196000_756000# gnd! 185.5fF
C41 diff_2122800_788400# gnd! 122.6fF
C42 diff_2170800_822000# gnd! 135.6fF
C43 diff_2418000_853200# gnd! 72.3fF
C44 diff_2124000_754800# gnd! 242.1fF
C45 diff_1790400_450000# gnd! 371.6fF
C46 diff_1483200_518400# gnd! 93.8fF
C47 diff_1057200_405600# gnd! 35.8fF
C48 diff_1040400_404400# gnd! 38.1fF
C49 diff_1050000_252000# gnd! 440.7fF
C50 diff_970800_408000# gnd! 49.2fF
C51 diff_951600_416400# gnd! 51.9fF
C52 diff_588000_249600# gnd! 133.8fF
C53 diff_612000_230400# gnd! 112.4fF
C54 diff_697200_285600# gnd! 554.6fF
C55 diff_627600_302400# gnd! 35.2fF
C56 diff_163200_169200# gnd! 13.7fF ;**FLOATING
C57 diff_158400_180000# gnd! 18.5fF ;**FLOATING
C58 diff_154800_187200# gnd! 100.7fF ;**FLOATING
C59 diff_549600_303600# gnd! 141.2fF
C60 diff_962400_302400# gnd! 838.0fF
C61 diff_873600_433200# gnd! 139.5fF
C62 diff_1171200_472800# gnd! 33.3fF
C63 diff_661200_249600# gnd! 453.6fF
C64 diff_1118400_457200# gnd! 83.7fF
C65 diff_1171200_489600# gnd! 38.8fF
C66 diff_1171200_454800# gnd! 132.4fF
C67 diff_980400_405600# gnd! 568.8fF
C68 diff_1424400_518400# gnd! 80.2fF
C69 diff_1737600_447600# gnd! 271.8fF
C70 diff_1588800_609600# gnd! 74.5fF
C71 diff_1640400_600000# gnd! 122.0fF
C72 diff_1086000_459600# gnd! 136.2fF
C73 diff_850800_457200# gnd! 568.3fF
C74 diff_1887600_652800# gnd! 109.6fF
C75 diff_1887600_699600# gnd! 228.3fF
C76 diff_2006400_746400# gnd! 90.6fF
C77 diff_1963200_744000# gnd! 102.7fF
C78 diff_1852800_734400# gnd! 98.5fF
C79 diff_1864800_708000# gnd! 104.3fF
C80 diff_1940400_778800# gnd! 98.6fF
C81 diff_1874400_784800# gnd! 209.8fF
C82 diff_1866000_762000# gnd! 249.3fF
C83 diff_1730400_746400# gnd! 89.7fF
C84 diff_1790400_692400# gnd! 153.6fF
C85 diff_1688400_740400# gnd! 99.6fF
C86 diff_410400_252000# gnd! 251.1fF
C87 diff_414000_259200# gnd! 52.8fF
C88 diff_366000_230400# gnd! 105.5fF
C89 diff_460800_272400# gnd! 103.9fF
C90 diff_477600_328800# gnd! 198.5fF
C91 diff_338400_282000# gnd! 118.1fF
C92 diff_810000_472800# gnd! 188.2fF
C93 diff_776400_445200# gnd! 106.3fF
C94 diff_656400_399600# gnd! 112.9fF
C95 diff_729600_462000# gnd! 131.5fF
C96 p0 gnd! 1186.4fF
C97 diff_310800_465600# gnd! 94.1fF
C98 diff_307200_476400# gnd! 72.3fF
C99 diff_356400_482400# gnd! 75.0fF
C100 diff_744000_516000# gnd! 138.1fF
C101 diff_352800_493200# gnd! 54.6fF
C102 diff_285600_456000# gnd! 68.6fF
C103 diff_550800_528000# gnd! 122.2fF
C104 diff_604800_403200# gnd! 222.7fF
C105 diff_733200_441600# gnd! 200.9fF
C106 diff_632400_480000# gnd! 325.1fF
C107 diff_356400_542400# gnd! 82.5fF
C108 diff_554400_499200# gnd! 469.2fF
C109 diff_354000_553200# gnd! 54.2fF
C110 diff_554400_535200# gnd! 207.4fF
C111 diff_356400_602400# gnd! 77.2fF
C112 diff_962400_673200# gnd! 539.1fF
C113 diff_1588800_708000# gnd! 106.2fF
C114 diff_1578000_711600# gnd! 96.2fF
C115 diff_1816800_742800# gnd! 126.7fF
C116 diff_1664400_780000# gnd! 97.9fF
C117 diff_1599600_784800# gnd! 382.4fF
C118 diff_1590000_762000# gnd! 379.1fF
C119 diff_1512000_679200# gnd! 157.6fF
C120 diff_1454400_751200# gnd! 94.6fF
C121 diff_1412400_741600# gnd! 107.0fF
C122 diff_1303200_711600# gnd! 97.2fF
C123 diff_1314000_708000# gnd! 109.5fF
C124 diff_1540800_742800# gnd! 127.9fF
C125 diff_2187600_633600# gnd! 475.4fF
C126 diff_2436000_927600# gnd! 64.6fF
C127 diff_1389600_780000# gnd! 96.5fF
C128 diff_1324800_784800# gnd! 388.1fF
C129 diff_1315200_762000# gnd! 378.9fF
C130 diff_1240800_674400# gnd! 164.9fF
C131 diff_1179600_747600# gnd! 97.0fF
C132 diff_1137600_742800# gnd! 106.7fF
C133 diff_1039200_708000# gnd! 113.6fF
C134 diff_1027200_728400# gnd! 99.4fF
C135 diff_1266000_742800# gnd! 118.0fF
C136 diff_1585200_432000# gnd! 375.4fF
C137 diff_1489200_434400# gnd! 590.6fF
C138 diff_1873200_825600# gnd! 295.9fF
C139 diff_1692000_622800# gnd! 452.7fF
C140 diff_1113600_780000# gnd! 102.6fF
C141 diff_1050000_784800# gnd! 389.2fF
C142 diff_1039200_816000# gnd! 384.7fF
C143 diff_966000_679200# gnd! 159.8fF
C144 diff_904800_746400# gnd! 96.9fF
C145 diff_862800_740400# gnd! 107.1fF
C146 diff_354000_610800# gnd! 59.0fF
C147 diff_379200_640800# gnd! 79.5fF
C148 diff_764400_708000# gnd! 108.3fF
C149 diff_544800_702000# gnd! 96.8fF
C150 diff_378000_734400# gnd! 62.1fF
C151 sync gnd! 1378.5fF
C152 diff_754800_711600# gnd! 85.6fF
C153 diff_950400_691200# gnd! 711.5fF
C154 diff_991200_742800# gnd! 118.0fF
C155 diff_396000_693600# gnd! 213.1fF
C156 diff_543600_736800# gnd! 294.3fF
C157 diff_838800_780000# gnd! 105.3fF
C158 diff_775200_784800# gnd! 387.2fF
C159 diff_764400_816000# gnd! 380.0fF
C160 diff_386400_644400# gnd! 703.2fF
C161 diff_1598400_825600# gnd! 384.4fF
C162 diff_1323600_825600# gnd! 255.6fF
C163 diff_3600_802800# gnd! 1186.8fF ;**FLOATING
C164 diff_237600_862800# gnd! 107.9fF
C165 diff_1784400_810000# gnd! 358.3fF
C166 diff_1430400_934800# gnd! 288.6fF
C167 diff_1042800_823200# gnd! 580.4fF
C168 diff_768000_823200# gnd! 359.5fF
C169 diff_1155600_936000# gnd! 281.8fF
C170 diff_880800_946800# gnd! 291.8fF
C171 diff_2436000_1012800# gnd! 70.8fF
C172 diff_1778400_1006800# gnd! 79.0fF
C173 diff_1700400_1006800# gnd! 59.0fF
C174 diff_1773600_999600# gnd! 215.2fF
C175 diff_2395200_1130400# gnd! 131.3fF
C176 diff_1879200_1021200# gnd! 209.2fF
C177 diff_848400_968400# gnd! 1058.8fF
C178 diff_2020800_1093200# gnd! 146.1fF
C179 diff_880800_992400# gnd! 903.8fF
C180 diff_1970400_1102800# gnd! 138.2fF
C181 diff_1890000_1120800# gnd! 149.1fF
C182 diff_1819200_1102800# gnd! 132.1fF
C183 diff_1766400_1093200# gnd! 133.2fF
C184 diff_1694400_1102800# gnd! 132.4fF
C185 diff_1633200_1118400# gnd! 147.8fF
C186 diff_1401600_975600# gnd! 167.5fF
C187 diff_1556400_1104000# gnd! 144.5fF
C188 diff_1496400_1116000# gnd! 148.7fF
C189 diff_2328000_1167600# gnd! 106.3fF
C190 diff_1696800_1017600# gnd! 339.4fF
C191 diff_1419600_1102800# gnd! 146.6fF
C192 diff_1358400_1116000# gnd! 148.3fF
C193 diff_1281600_1104000# gnd! 143.7fF
C194 diff_1221600_1120800# gnd! 146.6fF
C195 diff_1126800_975600# gnd! 178.3fF
C196 diff_1144800_1102800# gnd! 146.5fF
C197 diff_1083600_1118400# gnd! 149.4fF
C198 diff_1008000_1102800# gnd! 145.4fF
C199 diff_948000_1117200# gnd! 145.9fF
C200 diff_824400_1027200# gnd! 152.7fF
C201 diff_574800_1065600# gnd! 142.1fF
C202 diff_219600_991200# gnd! 184.9fF
C203 diff_224400_1065600# gnd! 146.3fF
C204 diff_561600_1051200# gnd! 125.5fF
C205 diff_870000_1102800# gnd! 149.8fF
C206 diff_202800_511200# gnd! 653.3fF
C207 diff_808800_1118400# gnd! 148.6fF
C208 diff_574800_1088400# gnd! 139.9fF
C209 diff_566400_924000# gnd! 801.8fF
C210 diff_248400_1088400# gnd! 67.8fF
C211 diff_219600_1101600# gnd! 70.1fF
C212 diff_1888800_1220400# gnd! 389.5fF
C213 diff_2338800_1209600# gnd! 166.3fF
C214 diff_883200_1207200# gnd! 589.5fF
C215 diff_822000_1227600# gnd! 613.9fF
C216 diff_1974000_1245600# gnd! 277.6fF
C217 diff_2308800_1185600# gnd! 149.6fF
C218 diff_840000_1020000# gnd! 796.0fF
C219 diff_516000_1240800# gnd! 164.5fF
C220 diff_1960800_1270800# gnd! 342.1fF
C221 diff_822000_1273200# gnd! 650.4fF
C222 diff_516000_1267200# gnd! 197.5fF
C223 diff_1902000_1294800# gnd! 285.8fF
C224 diff_2305200_1270800# gnd! 119.9fF
C225 diff_1096800_1296000# gnd! 631.6fF
C226 diff_2076000_1311600# gnd! 142.9fF
C227 diff_822000_1320000# gnd! 615.4fF
C228 diff_516000_1311600# gnd! 207.3fF
C229 diff_732000_1252800# gnd! 95.1fF
C230 diff_219600_942000# gnd! 1358.8fF
C231 diff_2335200_1249200# gnd! 194.7fF
C232 diff_2310000_1364400# gnd! 254.4fF
C233 diff_783600_224400# gnd! 931.0fF
C234 diff_2349600_1450800# gnd! 117.4fF
C235 diff_268800_446400# gnd! 877.0fF
C236 diff_824400_1339200# gnd! 538.3fF
C237 diff_1302000_1048800# gnd! 469.0fF
C238 diff_516000_1338000# gnd! 309.5fF
C239 diff_170400_1274400# gnd! 239.3fF
C240 diff_2053200_1180800# gnd! 412.1fF
C241 diff_2011200_1227600# gnd! 413.2fF
C242 diff_2106000_1476000# gnd! 127.9fF
C243 diff_1965600_1276800# gnd! 359.4fF
C244 diff_1892400_1160400# gnd! 363.0fF
C245 diff_2037600_1422000# gnd! 128.2fF
C246 diff_1968000_1476000# gnd! 125.8fF
C247 diff_1820400_1143600# gnd! 424.5fF
C248 diff_1759200_1120800# gnd! 404.2fF
C249 diff_1899600_1422000# gnd! 133.6fF
C250 diff_1830000_1476000# gnd! 128.6fF
C251 diff_1692000_1450800# gnd! 383.5fF
C252 diff_1634400_1160400# gnd! 364.5fF
C253 diff_1761600_1422000# gnd! 132.6fF
C254 diff_1692000_1476000# gnd! 132.7fF
C255 diff_1555200_1450800# gnd! 367.4fF
C256 diff_1497600_1159200# gnd! 338.7fF
C257 diff_1624800_1396800# gnd! 130.0fF
C258 diff_1555200_1476000# gnd! 129.6fF
C259 diff_1417200_1450800# gnd! 361.8fF
C260 diff_1359600_1159200# gnd! 363.0fF
C261 diff_1486800_1422000# gnd! 133.1fF
C262 diff_1417200_1476000# gnd! 132.5fF
C263 diff_1350000_1389600# gnd! 131.0fF
C264 diff_1280400_1450800# gnd! 353.5fF
C265 diff_1221600_1159200# gnd! 360.8fF
C266 diff_1280400_1476000# gnd! 132.6fF
C267 diff_1142400_1450800# gnd! 359.3fF
C268 diff_1084800_1160400# gnd! 361.9fF
C269 diff_1212000_1422000# gnd! 133.3fF
C270 diff_1142400_1476000# gnd! 132.7fF
C271 diff_1005600_1450800# gnd! 357.2fF
C272 diff_946800_1120800# gnd! 355.8fF
C273 diff_1075200_1389600# gnd! 133.2fF
C274 diff_1005600_1476000# gnd! 128.7fF
C275 diff_163200_1244400# gnd! 246.9fF
C276 diff_820800_1420800# gnd! 1693.1fF
C277 diff_844800_1435200# gnd! 1426.5fF
C278 diff_867600_1452000# gnd! 360.4fF
C279 diff_810000_1159200# gnd! 361.8fF
C280 diff_732000_1375200# gnd! 108.3fF
C281 diff_714000_876000# gnd! 1355.1fF
C282 diff_937200_1422000# gnd! 133.1fF
C283 diff_867600_1476000# gnd! 131.1fF
C284 diff_798000_1424400# gnd! 137.8fF
C285 diff_2346000_1502400# gnd! 155.7fF
C286 diff_2340000_1480800# gnd! 190.5fF
C287 clk1 gnd! 1830.0fF
C288 diff_2143200_1556400# gnd! 33.1fF
C289 diff_2342400_1538400# gnd! 178.6fF
C290 diff_2118000_1537200# gnd! 69.6fF
C291 diff_2143200_1588800# gnd! 33.1fF
C292 diff_2282400_1605600# gnd! 115.1fF
C293 diff_2052000_1551600# gnd! 29.3fF
C294 diff_2041200_1537200# gnd! 70.1fF
C295 diff_1980000_1537200# gnd! 69.0fF
C296 diff_2005200_1556400# gnd! 32.1fF
C297 diff_2118000_1621200# gnd! 68.7fF
C298 diff_2118000_1677600# gnd! 69.5fF
C299 diff_2143200_1698000# gnd! 33.4fF
C300 diff_1792800_176400# gnd! 880.5fF
C301 diff_2143200_1730400# gnd! 34.2fF
C302 diff_2052000_1592400# gnd! 30.4fF
C303 diff_2005200_1588800# gnd! 33.4fF
C304 diff_2041200_1620000# gnd! 70.4fF
C305 diff_1914000_1550400# gnd! 30.5fF
C306 diff_1903200_1537200# gnd! 72.4fF
C307 diff_1843200_1536000# gnd! 69.7fF
C308 diff_1867200_1556400# gnd! 33.6fF
C309 diff_1980000_1621200# gnd! 68.5fF
C310 diff_2052000_1692000# gnd! 30.2fF
C311 diff_2041200_1678800# gnd! 70.1fF
C312 diff_1980000_1677600# gnd! 69.7fF
C313 diff_2005200_1698000# gnd! 33.6fF
C314 diff_2118000_1764000# gnd! 69.2fF
C315 diff_2118000_1820400# gnd! 70.3fF
C316 diff_2143200_1839600# gnd! 33.5fF
C317 diff_2143200_1873200# gnd! 33.4fF
C318 o3 gnd! 497.5fF
C319 diff_2052000_1734000# gnd! 30.4fF
C320 diff_2005200_1730400# gnd! 33.9fF
C321 diff_2041200_1761600# gnd! 72.0fF
C322 diff_1914000_1592400# gnd! 30.7fF
C323 diff_1867200_1588800# gnd! 33.5fF
C324 diff_1903200_1620000# gnd! 70.1fF
C325 diff_1776000_1550400# gnd! 30.8fF
C326 diff_1765200_1538400# gnd! 71.5fF
C327 diff_1730400_1555200# gnd! 30.9fF
C328 diff_1705200_1536000# gnd! 69.8fF
C329 diff_1843200_1621200# gnd! 68.0fF
C330 diff_1914000_1692000# gnd! 30.8fF
C331 diff_1903200_1678800# gnd! 70.3fF
C332 diff_1843200_1677600# gnd! 68.5fF
C333 diff_1867200_1698000# gnd! 33.9fF
C334 diff_1980000_1764000# gnd! 69.7fF
C335 diff_2052000_1834800# gnd! 30.4fF
C336 diff_2005200_1839600# gnd! 33.5fF
C337 diff_2041200_1820400# gnd! 69.9fF
C338 diff_1980000_1820400# gnd! 68.5fF
C339 diff_2118000_1905600# gnd! 67.5fF
C340 diff_2118000_1962000# gnd! 68.1fF
C341 diff_2143200_1982400# gnd! 33.6fF
C342 diff_2374800_2004000# gnd! 222.4fF
C343 diff_2455200_2066400# gnd! 80.5fF
C344 diff_2425200_2089200# gnd! 70.7fF
C345 diff_2143200_2014800# gnd! 33.9fF
C346 diff_2052000_1875600# gnd! 29.4fF
C347 diff_2005200_1873200# gnd! 33.6fF
C348 diff_2041200_1903200# gnd! 68.5fF
C349 diff_1914000_1734000# gnd! 30.7fF
C350 diff_1867200_1730400# gnd! 34.0fF
C351 diff_1903200_1761600# gnd! 70.3fF
C352 diff_1776000_1592400# gnd! 30.8fF
C353 diff_1730400_1588800# gnd! 30.8fF
C354 diff_1765200_1621200# gnd! 69.3fF
C355 diff_1638000_1550400# gnd! 31.2fF
C356 diff_1592400_1555200# gnd! 30.8fF
C357 diff_1628400_1537200# gnd! 69.8fF
C358 diff_1567200_1536000# gnd! 72.7fF
C359 diff_1705200_1621200# gnd! 66.8fF
C360 diff_1638000_1592400# gnd! 31.3fF
C361 diff_1592400_1588800# gnd! 30.8fF
C362 diff_1628400_1620000# gnd! 68.1fF
C363 diff_1776000_1692000# gnd! 30.8fF
C364 diff_1765200_1678800# gnd! 69.1fF
C365 diff_1705200_1677600# gnd! 67.9fF
C366 diff_1730400_1696800# gnd! 30.9fF
C367 diff_1843200_1762800# gnd! 70.4fF
C368 diff_1914000_1834800# gnd! 30.8fF
C369 diff_1843200_1819200# gnd! 69.7fF
C370 diff_1867200_1839600# gnd! 33.8fF
C371 diff_1903200_1820400# gnd! 70.1fF
C372 diff_1980000_1905600# gnd! 69.4fF
C373 diff_2052000_1976400# gnd! 30.6fF
C374 diff_2041200_1962000# gnd! 68.3fF
C375 diff_2005200_1982400# gnd! 33.4fF
C376 diff_1980000_1962000# gnd! 68.8fF
C377 diff_2118000_2048400# gnd! 68.4fF
C378 diff_2143200_2124000# gnd! 33.5fF
C379 diff_2344800_2140800# gnd! 310.7fF
C380 diff_2325600_2148000# gnd! 34.6fF
C381 diff_2118000_2104800# gnd! 69.1fF
C382 diff_2416800_1954800# gnd! 394.4fF
C383 diff_2143200_2157600# gnd! 32.6fF
C384 diff_2052000_2018400# gnd! 30.4fF
C385 diff_2005200_2014800# gnd! 33.9fF
C386 diff_2041200_2044800# gnd! 68.9fF
C387 diff_1914000_1875600# gnd! 31.8fF
C388 diff_1867200_1872000# gnd! 34.6fF
C389 diff_1903200_1903200# gnd! 70.0fF
C390 diff_1776000_1734000# gnd! 31.2fF
C391 diff_1730400_1730400# gnd! 29.5fF
C392 diff_1765200_1762800# gnd! 71.1fF
C393 diff_1501200_1551600# gnd! 30.9fF
C394 diff_1490400_1537200# gnd! 73.6fF
C395 diff_1454400_1556400# gnd! 33.3fF
C396 diff_1430400_1536000# gnd! 69.6fF
C397 diff_1567200_1621200# gnd! 70.0fF
C398 diff_1638000_1692000# gnd! 30.9fF
C399 diff_1628400_1677600# gnd! 68.3fF
C400 diff_1592400_1696800# gnd! 30.6fF
C401 diff_1567200_1677600# gnd! 71.2fF
C402 diff_1638000_1734000# gnd! 32.6fF
C403 diff_1705200_1764000# gnd! 69.3fF
C404 diff_1592400_1730400# gnd! 31.2fF
C405 diff_1628400_1760400# gnd! 69.5fF
C406 diff_1776000_1833600# gnd! 31.5fF
C407 diff_1765200_1822800# gnd! 70.6fF
C408 diff_1705200_1819200# gnd! 69.2fF
C409 diff_1730400_1838400# gnd! 31.5fF
C410 diff_1843200_1905600# gnd! 68.8fF
C411 diff_1914000_1976400# gnd! 30.6fF
C412 diff_1903200_1962000# gnd! 68.8fF
C413 diff_1843200_1962000# gnd! 68.3fF
C414 diff_1867200_1982400# gnd! 33.9fF
C415 diff_1980000_2047200# gnd! 68.2fF
C416 diff_2052000_2119200# gnd! 30.4fF
C417 diff_2005200_2124000# gnd! 33.4fF
C418 diff_2041200_2103600# gnd! 69.9fF
C419 diff_1980000_2104800# gnd! 70.2fF
C420 diff_2118000_2190000# gnd! 67.9fF
C421 diff_2118000_2245200# gnd! 68.5fF
C422 diff_2143200_2265600# gnd! 32.9fF
C423 diff_2143200_2298000# gnd! 33.9fF
C424 diff_2052000_2160000# gnd! 29.4fF
C425 diff_2005200_2157600# gnd! 32.9fF
C426 diff_2041200_2187600# gnd! 70.1fF
C427 diff_1914000_2018400# gnd! 30.7fF
C428 diff_1867200_2014800# gnd! 33.9fF
C429 diff_1903200_2044800# gnd! 70.4fF
C430 diff_1776000_1875600# gnd! 31.9fF
C431 diff_1730400_1872000# gnd! 31.8fF
C432 diff_1765200_1904400# gnd! 68.4fF
C433 diff_1501200_1592400# gnd! 30.5fF
C434 diff_1454400_1588800# gnd! 33.6fF
C435 diff_1490400_1620000# gnd! 72.0fF
C436 diff_1363200_1551600# gnd! 30.4fF
C437 diff_1353600_1537200# gnd! 71.2fF
C438 diff_1292400_1536000# gnd! 71.8fF
C439 diff_1317600_1555200# gnd! 30.9fF
C440 diff_1430400_1621200# gnd! 69.2fF
C441 diff_1501200_1692000# gnd! 30.8fF
C442 diff_1490400_1677600# gnd! 70.7fF
C443 diff_1430400_1677600# gnd! 67.9fF
C444 diff_1454400_1696800# gnd! 33.5fF
C445 diff_1567200_1764000# gnd! 72.5fF
C446 diff_1638000_1833600# gnd! 34.2fF
C447 diff_1628400_1819200# gnd! 69.0fF
C448 diff_1567200_1819200# gnd! 71.6fF
C449 diff_1592400_1838400# gnd! 31.4fF
C450 diff_1705200_1904400# gnd! 69.4fF
C451 diff_1776000_1976400# gnd! 31.1fF
C452 diff_1766400_1960800# gnd! 69.4fF
C453 diff_1705200_1962000# gnd! 66.5fF
C454 diff_1730400_1981200# gnd! 31.2fF
C455 diff_1843200_2047200# gnd! 69.0fF
C456 diff_1914000_2119200# gnd! 30.7fF
C457 diff_1903200_2103600# gnd! 70.0fF
C458 diff_1843200_2103600# gnd! 68.9fF
C459 diff_1867200_2124000# gnd! 33.5fF
C460 diff_1980000_2190000# gnd! 68.8fF
C461 diff_2052000_2259600# gnd! 30.3fF
C462 diff_2041200_2246400# gnd! 70.3fF
C463 diff_2005200_2265600# gnd! 33.6fF
C464 diff_1980000_2245200# gnd! 69.6fF
C465 diff_2118000_2330400# gnd! 68.0fF
C466 diff_2118000_2386800# gnd! 68.1fF
C467 diff_2143200_2407200# gnd! 33.6fF
C468 o2 gnd! 617.9fF
C469 diff_2374800_2434800# gnd! 218.7fF
C470 diff_2143200_2439600# gnd! 33.5fF
C471 diff_2455200_2494800# gnd! 77.6fF
C472 diff_2424000_2518800# gnd! 75.6fF
C473 diff_2052000_2301600# gnd! 30.4fF
C474 diff_2005200_2298000# gnd! 33.9fF
C475 diff_2041200_2329200# gnd! 69.5fF
C476 diff_1914000_2160000# gnd! 30.4fF
C477 diff_1867200_2156400# gnd! 33.5fF
C478 diff_1903200_2187600# gnd! 69.2fF
C479 diff_1730400_2014800# gnd! 29.1fF
C480 diff_1776000_2018400# gnd! 31.2fF
C481 diff_1766400_2044800# gnd! 69.8fF
C482 diff_1638000_1875600# gnd! 34.7fF
C483 diff_1592400_1872000# gnd! 31.9fF
C484 diff_1628400_1903200# gnd! 67.6fF
C485 diff_1501200_1734000# gnd! 30.5fF
C486 diff_1454400_1730400# gnd! 33.6fF
C487 diff_1490400_1761600# gnd! 71.7fF
C488 diff_1363200_1592400# gnd! 30.5fF
C489 diff_1317600_1588800# gnd! 30.8fF
C490 diff_1353600_1620000# gnd! 70.7fF
C491 diff_1363200_1692000# gnd! 30.8fF
C492 diff_1353600_1677600# gnd! 69.5fF
C493 diff_1226400_1550400# gnd! 31.4fF
C494 diff_1215600_1537200# gnd! 72.8fF
C495 diff_1180800_1554000# gnd! 31.4fF
C496 diff_1155600_1536000# gnd! 70.1fF
C497 diff_1292400_1621200# gnd! 71.2fF
C498 diff_1292400_1677600# gnd! 69.1fF
C499 diff_1317600_1696800# gnd! 31.1fF
C500 diff_1430400_1764000# gnd! 69.0fF
C501 diff_1363200_1734000# gnd! 30.7fF
C502 diff_1317600_1730400# gnd! 31.2fF
C503 diff_1353600_1760400# gnd! 70.3fF
C504 diff_1501200_1834800# gnd! 30.8fF
C505 diff_1490400_1819200# gnd! 70.9fF
C506 diff_1430400_1819200# gnd! 70.0fF
C507 diff_1454400_1839600# gnd! 33.6fF
C508 diff_1567200_1904400# gnd! 71.7fF
C509 diff_1638000_1976400# gnd! 33.3fF
C510 diff_1628400_1962000# gnd! 66.7fF
C511 diff_1592400_1981200# gnd! 30.6fF
C512 diff_1567200_1962000# gnd! 71.3fF
C513 diff_1705200_2047200# gnd! 67.8fF
C514 diff_1776000_2118000# gnd! 31.4fF
C515 diff_1765200_2109600# gnd! 69.3fF
C516 diff_1705200_2103600# gnd! 67.6fF
C517 diff_1730400_2122800# gnd! 31.7fF
C518 diff_1843200_2188800# gnd! 68.2fF
C519 diff_1914000_2259600# gnd! 30.9fF
C520 diff_1903200_2246400# gnd! 70.9fF
C521 diff_1842000_2251200# gnd! 69.9fF
C522 diff_1867200_2265600# gnd! 33.4fF
C523 diff_1980000_2330400# gnd! 68.6fF
C524 diff_2052000_2402400# gnd! 29.2fF
C525 diff_2041200_2386800# gnd! 69.8fF
C526 diff_1980000_2386800# gnd! 68.9fF
C527 diff_2005200_2407200# gnd! 32.9fF
C528 diff_2118000_2472000# gnd! 67.2fF
C529 diff_2118000_2528400# gnd! 68.3fF
C530 diff_2143200_2548800# gnd! 27.5fF
C531 diff_2344800_2570400# gnd! 307.1fF
C532 diff_2325600_2576400# gnd! 34.9fF
C533 diff_2414400_2601600# gnd! 388.5fF
C534 diff_2224800_1584000# gnd! 794.2fF
C535 diff_2143200_2581200# gnd! 34.5fF
C536 diff_2050800_2456400# gnd! 31.2fF
C537 diff_2005200_2439600# gnd! 33.7fF
C538 diff_2041200_2470800# gnd! 68.8fF
C539 diff_1914000_2301600# gnd! 30.7fF
C540 diff_1867200_2298000# gnd! 34.0fF
C541 diff_1903200_2329200# gnd! 69.5fF
C542 diff_1776000_2160000# gnd! 30.8fF
C543 diff_1729200_2158800# gnd! 31.6fF
C544 diff_1765200_2188800# gnd! 68.8fF
C545 diff_1638000_2018400# gnd! 34.0fF
C546 diff_1592400_2014800# gnd! 31.2fF
C547 diff_1628400_2044800# gnd! 68.2fF
C548 diff_1501200_1875600# gnd! 31.6fF
C549 diff_1454400_1872000# gnd! 34.9fF
C550 diff_1490400_1903200# gnd! 70.6fF
C551 diff_1226400_1592400# gnd! 30.7fF
C552 diff_1180800_1588800# gnd! 30.6fF
C553 diff_1215600_1620000# gnd! 72.4fF
C554 diff_1088400_1550400# gnd! 32.6fF
C555 diff_1042800_1555200# gnd! 31.7fF
C556 diff_1078800_1537200# gnd! 71.6fF
C557 diff_1018800_1528800# gnd! 71.9fF
C558 diff_1155600_1621200# gnd! 69.7fF
C559 diff_1088400_1592400# gnd! 30.7fF
C560 diff_1042800_1588800# gnd! 30.8fF
C561 diff_1078800_1620000# gnd! 70.9fF
C562 diff_1226400_1692000# gnd! 31.4fF
C563 diff_1215600_1677600# gnd! 70.8fF
C564 diff_1155600_1677600# gnd! 68.8fF
C565 diff_1180800_1694400# gnd! 30.9fF
C566 diff_1292400_1764000# gnd! 69.0fF
C567 diff_1363200_1834800# gnd! 30.8fF
C568 diff_1353600_1819200# gnd! 70.4fF
C569 diff_1292400_1820400# gnd! 70.7fF
C570 diff_1317600_1838400# gnd! 30.8fF
C571 diff_1430400_1904400# gnd! 69.1fF
C572 diff_1363200_1875600# gnd! 31.9fF
C573 diff_1317600_1872000# gnd! 29.8fF
C574 diff_1353600_1903200# gnd! 69.7fF
C575 diff_1501200_1976400# gnd! 30.6fF
C576 diff_1490400_1962000# gnd! 70.1fF
C577 diff_1454400_1981200# gnd! 33.6fF
C578 diff_1430400_1960800# gnd! 70.4fF
C579 diff_1567200_2047200# gnd! 70.7fF
C580 diff_1638000_2119200# gnd! 32.3fF
C581 diff_1628400_2103600# gnd! 68.4fF
C582 diff_1567200_2103600# gnd! 71.0fF
C583 diff_1592400_2122800# gnd! 30.8fF
C584 diff_1592400_2156400# gnd! 30.7fF
C585 diff_1638000_2160000# gnd! 31.1fF
C586 diff_1705200_2188800# gnd! 67.1fF
C587 diff_1628400_2187600# gnd! 67.7fF
C588 diff_1776000_2259600# gnd! 30.7fF
C589 diff_1765200_2246400# gnd! 69.5fF
C590 diff_1705200_2245200# gnd! 69.9fF
C591 diff_1729200_2264400# gnd! 33.0fF
C592 diff_1842000_2334000# gnd! 67.9fF
C593 diff_1914000_2401200# gnd! 30.9fF
C594 diff_1903200_2386800# gnd! 69.0fF
C595 diff_1842000_2389200# gnd! 68.8fF
C596 diff_1867200_2407200# gnd! 33.5fF
C597 diff_1980000_2472000# gnd! 68.3fF
C598 diff_2052000_2542800# gnd! 31.1fF
C599 diff_2041200_2528400# gnd! 69.7fF
C600 diff_1980000_2528400# gnd! 68.6fF
C601 diff_2005200_2548800# gnd! 33.7fF
C602 diff_2133600_1458000# gnd! 494.7fF
C603 diff_2110800_1458000# gnd! 457.6fF
C604 diff_2082000_1496400# gnd! 461.4fF
C605 diff_2052000_2584800# gnd! 30.4fF
C606 diff_2005200_2581200# gnd! 33.7fF
C607 diff_2046000_1444800# gnd! 494.3fF
C608 diff_2118000_2614800# gnd! 66.7fF
C609 diff_2041200_2612400# gnd! 67.4fF
C610 diff_1994400_1460400# gnd! 496.0fF
C611 diff_1914000_2443200# gnd! 30.7fF
C612 diff_1867200_2439600# gnd! 34.0fF
C613 diff_1903200_2470800# gnd! 68.7fF
C614 diff_1776000_2301600# gnd! 31.0fF
C615 diff_1729200_2298000# gnd! 33.5fF
C616 diff_1765200_2329200# gnd! 68.6fF
C617 diff_1501200_2018400# gnd! 30.5fF
C618 diff_1454400_2014800# gnd! 33.5fF
C619 diff_1490400_2044800# gnd! 71.2fF
C620 diff_1180800_1730400# gnd! 30.7fF
C621 diff_1226400_1734000# gnd! 31.2fF
C622 diff_1215600_1761600# gnd! 71.5fF
C623 diff_951600_1550400# gnd! 31.6fF
C624 diff_906000_1551600# gnd! 31.6fF
C625 diff_940800_1537200# gnd! 72.0fF
C626 diff_880800_1536000# gnd! 69.3fF
C627 diff_1018800_1621200# gnd! 71.4fF
C628 diff_1088400_1692000# gnd! 31.9fF
C629 diff_1078800_1677600# gnd! 69.3fF
C630 diff_1017600_1677600# gnd! 70.6fF
C631 diff_1042800_1696800# gnd! 31.9fF
C632 diff_1155600_1762800# gnd! 69.3fF
C633 diff_1088400_1734000# gnd! 31.4fF
C634 diff_1042800_1730400# gnd! 31.2fF
C635 diff_1078800_1761600# gnd! 70.8fF
C636 diff_1226400_1834800# gnd! 30.5fF
C637 diff_1155600_1819200# gnd! 69.6fF
C638 diff_1180800_1837200# gnd! 30.7fF
C639 diff_1215600_1819200# gnd! 71.7fF
C640 diff_1292400_1904400# gnd! 72.2fF
C641 diff_1226400_1875600# gnd! 31.5fF
C642 diff_1180800_1872000# gnd! 31.8fF
C643 diff_1215600_1903200# gnd! 71.9fF
C644 diff_1363200_1976400# gnd! 31.1fF
C645 diff_1353600_1962000# gnd! 70.8fF
C646 diff_1292400_1962000# gnd! 70.9fF
C647 diff_1317600_1981200# gnd! 31.3fF
C648 diff_1430400_2048400# gnd! 69.0fF
C649 diff_1363200_2018400# gnd! 30.7fF
C650 diff_1317600_2014800# gnd! 31.2fF
C651 diff_1353600_2044800# gnd! 69.8fF
C652 diff_1501200_2119200# gnd! 30.5fF
C653 diff_1490400_2103600# gnd! 71.5fF
C654 diff_1454400_2124000# gnd! 33.4fF
C655 diff_1430400_2104800# gnd! 69.6fF
C656 diff_1567200_2188800# gnd! 70.6fF
C657 diff_1638000_2259600# gnd! 31.2fF
C658 diff_1628400_2245200# gnd! 68.8fF
C659 diff_1567200_2245200# gnd! 70.4fF
C660 diff_1592400_2264400# gnd! 30.9fF
C661 diff_1705200_2330400# gnd! 66.2fF
C662 diff_1776000_2401200# gnd! 31.1fF
C663 diff_1765200_2388000# gnd! 70.1fF
C664 diff_1705200_2386800# gnd! 68.6fF
C665 diff_1729200_2407200# gnd! 33.7fF
C666 diff_1842000_2472000# gnd! 68.0fF
C667 diff_1914000_2542800# gnd! 31.2fF
C668 diff_1903200_2529600# gnd! 68.6fF
C669 diff_1843200_2528400# gnd! 68.2fF
C670 diff_1867200_2547600# gnd! 34.2fF
C671 diff_1972800_1458000# gnd! 461.8fF
C672 diff_1914000_2584800# gnd! 31.2fF
C673 diff_1867200_2581200# gnd! 33.9fF
C674 diff_1944000_1496400# gnd! 458.2fF
C675 diff_1980000_2614800# gnd! 68.1fF
C676 diff_1903200_2612400# gnd! 67.8fF
C677 diff_1908000_1442400# gnd! 493.2fF
C678 diff_1776000_2443200# gnd! 30.8fF
C679 diff_1729200_2439600# gnd! 33.6fF
C680 diff_1765200_2470800# gnd! 68.7fF
C681 diff_1638000_2301600# gnd! 30.8fF
C682 diff_1592400_2298000# gnd! 30.7fF
C683 diff_1628400_2328000# gnd! 67.0fF
C684 diff_1454400_2156400# gnd! 33.5fF
C685 diff_1501200_2160000# gnd! 30.9fF
C686 diff_1490400_2187600# gnd! 69.1fF
C687 diff_951600_1592400# gnd! 30.7fF
C688 diff_906000_1588800# gnd! 30.6fF
C689 diff_940800_1620000# gnd! 71.9fF
C690 diff_487200_1521600# gnd! 137.3fF
C691 diff_506400_1542000# gnd! 245.4fF
C692 diff_664800_1543200# gnd! 1396.2fF
C693 diff_814800_1551600# gnd! 30.7fF
C694 diff_804000_1537200# gnd! 72.6fF
C695 diff_880800_1621200# gnd! 69.2fF
C696 diff_951600_1692000# gnd! 31.8fF
C697 diff_940800_1677600# gnd! 69.7fF
C698 diff_880800_1677600# gnd! 67.7fF
C699 diff_906000_1693200# gnd! 31.0fF
C700 diff_1017600_1764000# gnd! 72.4fF
C701 diff_1088400_1834800# gnd! 30.8fF
C702 diff_1078800_1819200# gnd! 70.0fF
C703 diff_1017600_1820400# gnd! 70.7fF
C704 diff_1042800_1838400# gnd! 30.8fF
C705 diff_1155600_1904400# gnd! 67.7fF
C706 diff_1088400_1875600# gnd! 32.2fF
C707 diff_1042800_1872000# gnd! 31.9fF
C708 diff_1078800_1903200# gnd! 69.5fF
C709 diff_1226400_1976400# gnd! 31.1fF
C710 diff_1215600_1962000# gnd! 70.9fF
C711 diff_1180800_1980000# gnd! 30.7fF
C712 diff_1155600_1962000# gnd! 69.4fF
C713 diff_1292400_2047200# gnd! 69.7fF
C714 diff_1363200_2119200# gnd! 30.7fF
C715 diff_1353600_2103600# gnd! 69.7fF
C716 diff_1292400_2104800# gnd! 69.9fF
C717 diff_1317600_2122800# gnd! 30.7fF
C718 diff_1430400_2188800# gnd! 67.8fF
C719 diff_1363200_2160000# gnd! 30.5fF
C720 diff_1317600_2156400# gnd! 30.9fF
C721 diff_1353600_2187600# gnd! 68.7fF
C722 diff_1501200_2259600# gnd! 30.8fF
C723 diff_1490400_2246400# gnd! 69.8fF
C724 diff_1454400_2264400# gnd! 33.5fF
C725 diff_1430400_2245200# gnd! 68.4fF
C726 diff_1567200_2330400# gnd! 69.1fF
C727 diff_1638000_2401200# gnd! 30.9fF
C728 diff_1628400_2386800# gnd! 68.0fF
C729 diff_1567200_2386800# gnd! 68.7fF
C730 diff_1592400_2406000# gnd! 31.2fF
C731 diff_1705200_2472000# gnd! 67.0fF
C732 diff_1776000_2542800# gnd! 31.2fF
C733 diff_1765200_2529600# gnd! 69.0fF
C734 diff_1705200_2528400# gnd! 68.0fF
C735 diff_1729200_2547600# gnd! 34.2fF
C736 diff_1834800_1458000# gnd! 500.4fF
C737 diff_1806000_1496400# gnd! 456.1fF
C738 diff_1770000_1443600# gnd! 493.2fF
C739 diff_1776000_2584800# gnd! 31.2fF
C740 diff_1729200_2588400# gnd! 32.9fF
C741 diff_1856400_1458000# gnd! 494.7fF
C742 diff_1842000_2622000# gnd! 67.0fF
C743 diff_1765200_2612400# gnd! 68.0fF
C744 diff_1892400_663600# gnd! 1209.0fF
C745 diff_1638000_2443200# gnd! 30.8fF
C746 diff_1592400_2439600# gnd! 30.8fF
C747 diff_1628400_2470800# gnd! 67.4fF
C748 diff_1501200_2301600# gnd! 30.8fF
C749 diff_1454400_2298000# gnd! 33.4fF
C750 diff_1490400_2329200# gnd! 70.1fF
C751 diff_1180800_2014800# gnd! 30.6fF
C752 diff_1226400_2018400# gnd! 31.1fF
C753 diff_1215600_2044800# gnd! 71.7fF
C754 diff_951600_1734000# gnd! 31.8fF
C755 diff_906000_1730400# gnd! 31.0fF
C756 diff_940800_1761600# gnd! 71.7fF
C757 diff_813600_1597200# gnd! 31.3fF
C758 diff_548400_1543200# gnd! 714.9fF
C759 diff_568800_1560000# gnd! 197.4fF
C760 diff_804000_1620000# gnd! 71.9fF
C761 diff_664800_1620000# gnd! 1400.7fF
C762 diff_568800_1599600# gnd! 192.5fF
C763 diff_548400_1610400# gnd! 848.4fF
C764 diff_440400_1596000# gnd! 67.9fF
C765 diff_506400_1618800# gnd! 240.7fF
C766 diff_487200_1641600# gnd! 139.7fF
C767 diff_162000_1520400# gnd! 115.0fF
C768 diff_162000_1621200# gnd! 113.8fF
C769 diff_506400_1683600# gnd! 238.3fF
C770 diff_664800_1683600# gnd! 1257.2fF
C771 diff_813600_1692000# gnd! 34.4fF
C772 diff_804000_1677600# gnd! 69.3fF
C773 diff_880800_1762800# gnd! 69.2fF
C774 diff_951600_1834800# gnd! 30.8fF
C775 diff_940800_1819200# gnd! 71.2fF
C776 diff_880800_1820400# gnd! 69.4fF
C777 diff_906000_1836000# gnd! 30.5fF
C778 diff_1017600_1905600# gnd! 69.7fF
C779 diff_1088400_1976400# gnd! 32.2fF
C780 diff_1078800_1960800# gnd! 71.3fF
C781 diff_1017600_1962000# gnd! 71.7fF
C782 diff_1042800_1981200# gnd! 31.8fF
C783 diff_1155600_2048400# gnd! 68.1fF
C784 diff_1088400_2018400# gnd! 30.7fF
C785 diff_1042800_2014800# gnd! 31.2fF
C786 diff_1078800_2044800# gnd! 69.8fF
C787 diff_1226400_2119200# gnd! 30.5fF
C788 diff_1215600_2103600# gnd! 70.8fF
C789 diff_1155600_2103600# gnd! 68.4fF
C790 diff_1180800_2120400# gnd! 30.5fF
C791 diff_1292400_2188800# gnd! 68.9fF
C792 diff_1363200_2259600# gnd! 30.8fF
C793 diff_1353600_2245200# gnd! 70.4fF
C794 diff_1317600_2264400# gnd! 31.1fF
C795 diff_1292400_2245200# gnd! 69.6fF
C796 diff_1430400_2330400# gnd! 68.1fF
C797 diff_1500000_2420400# gnd! 31.0fF
C798 diff_1490400_2386800# gnd! 69.1fF
C799 diff_1454400_2406000# gnd! 33.4fF
C800 diff_1430400_2386800# gnd! 67.7fF
C801 diff_1567200_2472000# gnd! 67.3fF
C802 diff_1638000_2542800# gnd! 31.2fF
C803 diff_1628400_2528400# gnd! 67.4fF
C804 diff_1567200_2528400# gnd! 69.0fF
C805 diff_1592400_2547600# gnd! 30.7fF
C806 diff_1719600_1458000# gnd! 532.1fF
C807 diff_1696800_1458000# gnd! 456.4fF
C808 diff_1668000_1497600# gnd! 456.5fF
C809 diff_1638000_2584800# gnd! 30.8fF
C810 diff_1592400_2581200# gnd! 30.7fF
C811 diff_1633200_1442400# gnd! 504.8fF
C812 diff_1705200_2613600# gnd! 66.5fF
C813 diff_1628400_2611200# gnd! 67.2fF
C814 diff_1581600_1458000# gnd! 491.3fF
C815 diff_1501200_2443200# gnd! 30.7fF
C816 diff_1454400_2439600# gnd! 33.4fF
C817 diff_1490400_2470800# gnd! 68.3fF
C818 diff_1363200_2301600# gnd! 30.5fF
C819 diff_1317600_2298000# gnd! 31.2fF
C820 diff_1353600_2328000# gnd! 69.1fF
C821 diff_1363200_2401200# gnd! 31.2fF
C822 diff_1353600_2386800# gnd! 68.9fF
C823 diff_1180800_2156400# gnd! 30.6fF
C824 diff_1226400_2160000# gnd! 30.9fF
C825 diff_1215600_2187600# gnd! 70.2fF
C826 diff_951600_1875600# gnd! 31.5fF
C827 diff_906000_1872000# gnd! 31.8fF
C828 diff_940800_1903200# gnd! 70.7fF
C829 diff_813600_1734000# gnd! 34.7fF
C830 diff_804000_1760400# gnd! 70.9fF
C831 diff_548400_1684800# gnd! 833.5fF
C832 diff_568800_1701600# gnd! 189.2fF
C833 diff_423600_1570800# gnd! 288.0fF
C834 diff_487200_1690800# gnd! 156.1fF
C835 diff_664800_1760400# gnd! 1424.5fF
C836 diff_568800_1741200# gnd! 190.9fF
C837 diff_548400_1752000# gnd! 832.4fF
C838 diff_436800_1612800# gnd! 432.9fF
C839 diff_88800_1684800# gnd! 250.8fF
C840 diff_506400_1747200# gnd! 247.3fF
C841 diff_487200_1740000# gnd! 161.9fF
C842 diff_487200_1801200# gnd! 145.6fF
C843 diff_506400_1825200# gnd! 241.5fF
C844 diff_813600_1834800# gnd! 33.5fF
C845 diff_804000_1819200# gnd! 70.7fF
C846 diff_664800_1825200# gnd! 1408.6fF
C847 diff_548400_1826400# gnd! 1087.9fF
C848 diff_568800_1843200# gnd! 201.3fF
C849 diff_880800_1904400# gnd! 68.0fF
C850 diff_940800_1962000# gnd! 71.5fF
C851 diff_951600_1976400# gnd! 31.7fF
C852 diff_880800_1962000# gnd! 69.0fF
C853 diff_906000_1977600# gnd! 31.4fF
C854 diff_1017600_2048400# gnd! 69.8fF
C855 diff_1088400_2119200# gnd! 30.7fF
C856 diff_1078800_2103600# gnd! 69.6fF
C857 diff_1017600_2103600# gnd! 70.5fF
C858 diff_1042800_2122800# gnd! 30.6fF
C859 diff_1155600_2188800# gnd! 66.4fF
C860 diff_1226400_2259600# gnd! 30.8fF
C861 diff_1215600_2246400# gnd! 70.8fF
C862 diff_1155600_2245200# gnd! 69.1fF
C863 diff_1179600_2268000# gnd! 33.2fF
C864 diff_1292400_2330400# gnd! 68.5fF
C865 diff_1292400_2386800# gnd! 68.8fF
C866 diff_1317600_2406000# gnd! 31.5fF
C867 diff_1430400_2472000# gnd! 67.5fF
C868 diff_1501200_2542800# gnd! 30.7fF
C869 diff_1454400_2547600# gnd! 33.5fF
C870 diff_1430400_2528400# gnd! 68.1fF
C871 diff_1490400_2528400# gnd! 68.5fF
C872 diff_1558800_1458000# gnd! 458.0fF
C873 diff_1531200_1458000# gnd! 481.6fF
C874 diff_1495200_1443600# gnd! 491.7fF
C875 diff_1501200_2584800# gnd! 30.7fF
C876 diff_1454400_2581200# gnd! 33.8fF
C877 diff_1567200_2613600# gnd! 68.4fF
C878 diff_1490400_2612400# gnd! 68.9fF
C879 diff_1363200_2443200# gnd! 30.7fF
C880 diff_1317600_2439600# gnd! 30.8fF
C881 diff_1353600_2469600# gnd! 68.9fF
C882 diff_1226400_2301600# gnd! 30.7fF
C883 diff_1179600_2298000# gnd! 34.3fF
C884 diff_1215600_2329200# gnd! 70.2fF
C885 diff_1088400_2160000# gnd! 30.5fF
C886 diff_1042800_2156400# gnd! 30.7fF
C887 diff_1078800_2187600# gnd! 71.1fF
C888 diff_951600_2018400# gnd! 31.2fF
C889 diff_906000_2014800# gnd! 30.9fF
C890 diff_940800_2044800# gnd! 69.6fF
C891 diff_813600_1876800# gnd! 33.6fF
C892 diff_804000_1903200# gnd! 69.1fF
C893 diff_664800_1902000# gnd! 1267.1fF
C894 diff_568800_1882800# gnd! 203.1fF
C895 diff_440400_1879200# gnd! 67.1fF
C896 diff_548400_1893600# gnd! 878.1fF
C897 diff_506400_1902000# gnd! 240.4fF
C898 diff_487200_1924800# gnd! 146.6fF
C899 diff_69600_1911600# gnd! 901.3fF
C900 d3 gnd! 2592.0fF
C901 diff_68400_1594800# gnd! 835.6fF
C902 diff_506400_1968000# gnd! 237.0fF
C903 diff_664800_1966800# gnd! 1379.3fF
C904 diff_813600_1976400# gnd! 34.8fF
C905 diff_804000_1962000# gnd! 69.6fF
C906 diff_548400_1968000# gnd! 974.9fF
C907 diff_568800_1984800# gnd! 191.0fF
C908 diff_880800_2047200# gnd! 68.0fF
C909 diff_951600_2119200# gnd! 30.8fF
C910 diff_940800_2103600# gnd! 72.1fF
C911 diff_880800_2104800# gnd! 68.4fF
C912 diff_904800_2138400# gnd! 31.8fF
C913 diff_1017600_2188800# gnd! 70.7fF
C914 diff_1088400_2259600# gnd! 31.8fF
C915 diff_1078800_2245200# gnd! 71.3fF
C916 diff_1017600_2245200# gnd! 72.0fF
C917 diff_1042800_2263200# gnd! 31.4fF
C918 diff_1155600_2330400# gnd! 68.1fF
C919 diff_1088400_2300400# gnd! 31.2fF
C920 diff_1042800_2298000# gnd! 31.2fF
C921 diff_1078800_2328000# gnd! 69.5fF
C922 diff_1226400_2401200# gnd! 31.3fF
C923 diff_1215600_2386800# gnd! 70.0fF
C924 diff_1179600_2406000# gnd! 34.0fF
C925 diff_1155600_2386800# gnd! 67.8fF
C926 diff_1292400_2472000# gnd! 68.5fF
C927 diff_1363200_2542800# gnd! 30.7fF
C928 diff_1353600_2528400# gnd! 68.7fF
C929 diff_1292400_2528400# gnd! 68.3fF
C930 diff_1317600_2547600# gnd! 31.2fF
C931 diff_1443600_1458000# gnd! 495.8fF
C932 diff_1430400_2613600# gnd! 67.8fF
C933 diff_1422000_1458000# gnd! 483.6fF
C934 diff_1363200_2584800# gnd! 30.7fF
C935 diff_1317600_2581200# gnd! 31.2fF
C936 diff_1393200_1496400# gnd! 456.6fF
C937 diff_1353600_2611200# gnd! 68.4fF
C938 diff_1357200_1444800# gnd! 529.2fF
C939 diff_1226400_2443200# gnd! 30.7fF
C940 diff_1179600_2439600# gnd! 33.6fF
C941 diff_1215600_2470800# gnd! 68.6fF
C942 diff_951600_2160000# gnd! 30.9fF
C943 diff_904800_2156400# gnd! 32.0fF
C944 diff_813600_2018400# gnd! 34.2fF
C945 diff_804000_2044800# gnd! 70.1fF
C946 diff_487200_1975200# gnd! 155.1fF
C947 diff_423600_1854000# gnd! 287.2fF
C948 diff_664800_2044800# gnd! 1406.8fF
C949 diff_568800_2025600# gnd! 192.8fF
C950 diff_548400_2036400# gnd! 958.5fF
C951 diff_506400_2037600# gnd! 241.7fF
C952 diff_331200_1510800# gnd! 656.8fF
C953 diff_487200_2029200# gnd! 155.7fF
C954 diff_487200_2085600# gnd! 143.7fF
C955 diff_506400_2109600# gnd! 241.4fF
C956 diff_664800_2109600# gnd! 1442.8fF
C957 diff_813600_2119200# gnd! 33.5fF
C958 diff_804000_2103600# gnd! 70.3fF
C959 diff_813600_2160000# gnd! 33.5fF
C960 diff_548400_2109600# gnd! 828.2fF
C961 diff_568800_2127600# gnd! 194.9fF
C962 diff_940800_2187600# gnd! 71.6fF
C963 diff_880800_2188800# gnd! 68.0fF
C964 diff_804000_2187600# gnd! 68.8fF
C965 diff_951600_2259600# gnd! 31.5fF
C966 diff_940800_2246400# gnd! 72.2fF
C967 diff_880800_2245200# gnd! 69.0fF
C968 diff_904800_2264400# gnd! 33.8fF
C969 diff_1017600_2330400# gnd! 68.7fF
C970 diff_1017600_2386800# gnd! 68.3fF
C971 diff_1088400_2401200# gnd! 31.8fF
C972 diff_1078800_2386800# gnd! 69.2fF
C973 diff_1042800_2404800# gnd! 31.7fF
C974 diff_1155600_2472000# gnd! 67.0fF
C975 diff_1155600_2528400# gnd! 67.2fF
C976 diff_1179600_2547600# gnd! 33.9fF
C977 diff_1226400_2542800# gnd! 31.2fF
C978 diff_1215600_2528400# gnd! 69.0fF
C979 diff_1284000_1458000# gnd! 458.1fF
C980 diff_1256400_1458000# gnd! 495.8fF
C981 diff_1220400_1442400# gnd! 491.4fF
C982 diff_1179600_2581200# gnd! 33.9fF
C983 diff_1226400_2584800# gnd! 31.2fF
C984 diff_1306800_1458000# gnd! 491.7fF
C985 diff_1292400_2613600# gnd! 66.8fF
C986 diff_1215600_2611200# gnd! 69.5fF
C987 diff_1168800_1458000# gnd! 537.9fF
C988 diff_1088400_2443200# gnd! 30.7fF
C989 diff_1042800_2439600# gnd! 30.8fF
C990 diff_1078800_2469600# gnd! 69.1fF
C991 diff_951600_2301600# gnd! 30.8fF
C992 diff_904800_2298000# gnd! 34.2fF
C993 diff_940800_2329200# gnd! 70.4fF
C994 diff_664800_2186400# gnd! 1420.9fF
C995 diff_170400_2043600# gnd! 248.6fF
C996 diff_163200_2012400# gnd! 245.7fF
C997 diff_568800_2167200# gnd! 201.6fF
C998 diff_548400_2178000# gnd! 700.3fF
C999 diff_440400_2163600# gnd! 65.2fF
C1000 diff_506400_2186400# gnd! 241.4fF
C1001 diff_487200_2209200# gnd! 143.1fF
C1002 diff_506400_2251200# gnd! 237.4fF
C1003 diff_664800_2251200# gnd! 1270.8fF
C1004 diff_813600_2259600# gnd! 31.6fF
C1005 diff_804000_2245200# gnd! 69.4fF
C1006 diff_813600_2301600# gnd! 30.5fF
C1007 diff_880800_2330400# gnd! 68.3fF
C1008 diff_804000_2328000# gnd! 69.3fF
C1009 diff_950400_2408400# gnd! 33.7fF
C1010 diff_940800_2386800# gnd! 70.3fF
C1011 diff_880800_2386800# gnd! 68.5fF
C1012 diff_904800_2406000# gnd! 34.6fF
C1013 diff_1017600_2472000# gnd! 68.6fF
C1014 diff_1088400_2542800# gnd! 31.0fF
C1015 diff_1077600_2532000# gnd! 69.3fF
C1016 diff_1017600_2528400# gnd! 68.8fF
C1017 diff_1042800_2546400# gnd! 31.2fF
C1018 diff_1088400_2584800# gnd! 31.0fF
C1019 diff_1147200_1458000# gnd! 472.9fF
C1020 diff_1118400_1497600# gnd! 459.0fF
C1021 diff_1082400_1443600# gnd! 555.8fF
C1022 diff_1155600_2613600# gnd! 67.2fF
C1023 diff_1078800_2611200# gnd! 68.6fF
C1024 diff_1042800_2581200# gnd! 31.2fF
C1025 diff_950400_2443200# gnd! 33.4fF
C1026 diff_904800_2439600# gnd! 33.8fF
C1027 diff_940800_2470800# gnd! 67.6fF
C1028 diff_548400_2252400# gnd! 953.9fF
C1029 diff_567600_2274000# gnd! 192.8fF
C1030 diff_487200_2258400# gnd! 155.4fF
C1031 diff_423600_2138400# gnd! 281.6fF
C1032 diff_664800_2328000# gnd! 1303.6fF
C1033 diff_567600_2308800# gnd! 191.4fF
C1034 diff_548400_2319600# gnd! 823.0fF
C1035 diff_506400_2320800# gnd! 240.9fF
C1036 diff_162000_2286000# gnd! 114.9fF
C1037 diff_327600_1404000# gnd! 480.7fF
C1038 diff_487200_2312400# gnd! 158.2fF
C1039 diff_487200_2368800# gnd! 141.3fF
C1040 diff_231600_1357200# gnd! 2539.8fF
C1041 diff_506400_2392800# gnd! 242.8fF
C1042 diff_664800_2392800# gnd! 1271.3fF
C1043 diff_813600_2401200# gnd! 32.0fF
C1044 diff_804000_2386800# gnd! 69.8fF
C1045 diff_880800_2472000# gnd! 67.7fF
C1046 diff_813600_2443200# gnd! 30.4fF
C1047 diff_548400_2392800# gnd! 824.7fF
C1048 diff_567600_2410800# gnd! 198.5fF
C1049 diff_804000_2469600# gnd! 67.6fF
C1050 diff_950400_2565600# gnd! 32.0fF
C1051 diff_940800_2528400# gnd! 71.3fF
C1052 diff_904800_2547600# gnd! 34.5fF
C1053 diff_880800_2528400# gnd! 67.2fF
C1054 diff_1009200_1458000# gnd! 465.5fF
C1055 diff_981600_1458000# gnd! 486.7fF
C1056 diff_945600_1442400# gnd! 492.4fF
C1057 diff_951600_2584800# gnd! 31.2fF
C1058 diff_904800_2581200# gnd! 34.2fF
C1059 diff_1032000_1458000# gnd! 491.0fF
C1060 diff_1017600_2613600# gnd! 67.8fF
C1061 diff_940800_2611200# gnd! 70.2fF
C1062 diff_894000_1458000# gnd! 526.1fF
C1063 diff_162000_2388000# gnd! 112.5fF
C1064 diff_663600_2470800# gnd! 1319.4fF
C1065 diff_567600_2450400# gnd! 198.5fF
C1066 diff_548400_2460000# gnd! 821.4fF
C1067 diff_440400_2446800# gnd! 70.2fF
C1068 diff_506400_2467200# gnd! 244.9fF
C1069 diff_487200_2491200# gnd! 142.5fF
C1070 diff_87600_2492400# gnd! 246.6fF
C1071 diff_506400_2533200# gnd! 248.0fF
C1072 diff_664800_2534400# gnd! 1253.0fF
C1073 diff_813600_2542800# gnd! 31.5fF
C1074 diff_804000_2528400# gnd! 68.9fF
C1075 diff_813600_2584800# gnd! 31.1fF
C1076 diff_872400_1458000# gnd! 459.6fF
C1077 diff_843600_1497600# gnd! 493.2fF
C1078 diff_807600_1443600# gnd! 515.3fF
C1079 diff_880800_2613600# gnd! 68.0fF
C1080 diff_804000_2611200# gnd! 68.4fF
C1081 diff_548400_2534400# gnd! 866.1fF
C1082 diff_567600_2553600# gnd! 197.2fF
C1083 diff_487200_2554800# gnd! 158.5fF
C1084 diff_230400_2126400# gnd! 2163.8fF
C1085 diff_423600_2420400# gnd! 281.0fF
C1086 diff_663600_2611200# gnd! 1408.6fF
C1087 diff_567600_2590800# gnd! 195.2fF
C1088 diff_426000_1591200# gnd! 1113.8fF
C1089 diff_548400_2601600# gnd! 793.5fF
C1090 diff_506400_2604000# gnd! 250.9fF
C1091 diff_487200_2602800# gnd! 143.8fF
C1092 diff_523200_1467600# gnd! 737.8fF
C1093 diff_326400_2457600# gnd! 585.7fF
C1094 diff_2325600_2644800# gnd! 40.3fF
C1095 diff_2424000_2713200# gnd! 71.3fF
C1096 diff_2346000_2652000# gnd! 299.9fF
C1097 diff_2454000_2737200# gnd! 80.5fF
C1098 clk2 gnd! 2556.7fF
C1099 diff_2104800_2774400# gnd! 36.7fF
C1100 diff_69600_2534400# gnd! 903.5fF
C1101 d2 gnd! 2745.3fF
C1102 diff_68400_2361600# gnd! 833.1fF
C1103 o1 gnd! 687.0fF
C1104 diff_2373600_2752800# gnd! 235.8fF
C1105 diff_2415600_2852400# gnd! 405.3fF
C1106 diff_2074800_2772000# gnd! 1042.6fF
C1107 diff_222000_1082400# gnd! 529.2fF
C1108 diff_349200_1096800# gnd! 2225.8fF
C1109 diff_2050800_2889600# gnd! 66.3fF
C1110 diff_2016000_2904000# gnd! 70.4fF
C1111 diff_1923600_2864400# gnd! 218.2fF
C1112 diff_2077200_2900400# gnd! 522.7fF
C1113 o0 gnd! 757.7fF
C1114 diff_1358400_2856000# gnd! 113.6fF
C1115 diff_1261200_2857200# gnd! 116.5fF
C1116 diff_1009200_2812800# gnd! 245.1fF
C1117 diff_943200_2844000# gnd! 258.0fF
C1118 diff_1429200_2878800# gnd! 225.6fF
C1119 diff_1262400_2888400# gnd! 909.5fF
C1120 diff_1330800_2899200# gnd! 817.1fF
C1121 diff_252000_2766000# gnd! 2722.9fF
C1122 diff_386400_2857200# gnd! 116.3fF
C1123 Vdd gnd! 37125.4fF
C1124 diff_132000_2799600# gnd! 1242.2fF
C1125 diff_165600_2822400# gnd! 244.5fF
C1126 diff_97200_2845200# gnd! 261.9fF
C1127 diff_289200_2857200# gnd! 119.2fF
C1128 diff_457200_2878800# gnd! 244.2fF
C1129 diff_87600_2288400# gnd! 1447.8fF
C1130 diff_289200_2884800# gnd! 907.9fF
C1131 diff_358800_2898000# gnd! 830.3fF
C1132 diff_1916400_2860800# gnd! 411.9fF
C1133 d0 gnd! 2674.9fF
C1134 d1 gnd! 2657.9fF
C1135 diff_2017200_2959200# gnd! 288.6fF
