`include "common.h"

module chip_6502(
  input eclk, ereset,
  output ab0,
  output ab1,
  output ab2,
  output ab3,
  output ab4,
  output ab5,
  output ab6,
  output ab7,
  output ab8,
  output ab9,
  output ab10,
  output ab11,
  output ab12,
  output ab13,
  output ab14,
  output ab15,
  input db0_i,
  output db0_o,
  output db0_t,
  input db1_i,
  output db1_o,
  output db1_t,
  input db2_i,
  output db2_o,
  output db2_t,
  input db3_i,
  output db3_o,
  output db3_t,
  input db4_i,
  output db4_o,
  output db4_t,
  input db5_i,
  output db5_o,
  output db5_t,
  input db6_i,
  output db6_o,
  output db6_t,
  input db7_i,
  output db7_o,
  output db7_t,
  input res,
  output rw,
  output sync,
  input so,
  input clk0,
  output clk1out,
  output clk2out,
  input rdy,
  input nmi,
  input irq
);

  wire signed [`W-1:0] n_1247_port_13, n_1247_port_0, n_1247_v;
  wire signed [`W-1:0] _ABL7_port_3, _ABL7_port_1, _ABL7_v;
  wire signed [`W-1:0] _ABL6_port_3, _ABL6_port_1, _ABL6_v;
  wire signed [`W-1:0] _ABL5_port_3, _ABL5_port_0, _ABL5_v;
  wire signed [`W-1:0] _ABL3_port_3, _ABL3_port_0, _ABL3_v;
  wire signed [`W-1:0] _ABL2_port_2, _ABL2_port_3, _ABL2_v;
  wire signed [`W-1:0] _ABL1_port_2, _ABL1_port_3, _ABL1_v;
  wire signed [`W-1:0] _ABL0_port_2, _ABL0_port_3, _ABL0_v;
  wire signed [`W-1:0] dpc5_SADL_port_0, dpc5_SADL_port_7, dpc5_SADL_v;
  wire signed [`W-1:0] n_465_port_2, n_465_port_0, n_465_port_1, n_465_v;
  wire signed [`W-1:0] rw_port_0, rw_port_1, rw_v;
  wire signed [`W-1:0] idl7_port_2, idl7_port_0, idl7_port_1, idl7_v;
  wire signed [`W-1:0] idl6_port_2, idl6_port_0, idl6_port_1, idl6_v;
  wire signed [`W-1:0] idl5_port_2, idl5_port_0, idl5_port_1, idl5_v;
  wire signed [`W-1:0] idl4_port_2, idl4_port_0, idl4_port_1, idl4_v;
  wire signed [`W-1:0] idl3_port_2, idl3_port_0, idl3_port_1, idl3_v;
  wire signed [`W-1:0] idl2_port_2, idl2_port_0, idl2_port_1, idl2_v;
  wire signed [`W-1:0] idl1_port_2, idl1_port_0, idl1_port_1, idl1_v;
  wire signed [`W-1:0] idl0_port_2, idl0_port_0, idl0_port_1, idl0_v;
  wire signed [`W-1:0] n_733_port_2, n_733_port_3, n_733_port_0, n_733_port_1, n_733_v;
  wire signed [`W-1:0] dpc20_ADDSB06_port_0, dpc20_ADDSB06_port_5, dpc20_ADDSB06_v;
  wire signed [`W-1:0] n_1389_port_2, n_1389_port_3, n_1389_port_0, n_1389_port_1, n_1389_port_4, n_1389_v;
  wire signed [`W-1:0] n_1387_port_2, n_1387_port_3, n_1387_port_0, n_1387_port_1, n_1387_v;
  wire signed [`W-1:0] n_1383_port_2, n_1383_port_0, n_1383_port_1, n_1383_v;
  wire signed [`W-1:0] x6_port_0, x6_port_1, x6_v;
  wire signed [`W-1:0] irq_port_2, irq_v;
  wire signed [`W-1:0] n_1267_port_2, n_1267_port_3, n_1267_port_0, n_1267_v;
  wire signed [`W-1:0] n_7_port_2, n_7_port_4, n_7_v;
  wire signed [`W-1:0] n_3_port_2, n_3_port_3, n_3_port_0, n_3_port_1, n_3_port_4, n_3_v;
  wire signed [`W-1:0] aluanandb0_port_9, aluanandb0_port_3, aluanandb0_port_5, aluanandb0_v;
  wire signed [`W-1:0] aluanandb1_port_0, aluanandb1_port_1, aluanandb1_port_4, aluanandb1_port_5, aluanandb1_v;
  wire signed [`W-1:0] dasb6_port_3, dasb6_port_0, dasb6_port_5, dasb6_v;
  wire signed [`W-1:0] dasb5_port_3, dasb5_port_1, dasb5_port_5, dasb5_v;
  wire signed [`W-1:0] dasb3_port_3, dasb3_port_1, dasb3_port_5, dasb3_v;
  wire signed [`W-1:0] dasb2_port_3, dasb2_port_1, dasb2_port_5, dasb2_v;
  wire signed [`W-1:0] dasb1_port_3, dasb1_port_0, dasb1_port_5, dasb1_v;
  wire signed [`W-1:0] alu4_port_2, alu4_port_3, alu4_port_0, alu4_port_1, alu4_v;
  wire signed [`W-1:0] alu5_port_3, alu5_port_0, alu5_port_1, alu5_port_4, alu5_v;
  wire signed [`W-1:0] alu6_port_2, alu6_port_0, alu6_port_1, alu6_port_4, alu6_v;
  wire signed [`W-1:0] alu7_port_2, alu7_port_3, alu7_port_0, alu7_port_1, alu7_v;
  wire signed [`W-1:0] alu0_port_2, alu0_port_3, alu0_port_0, alu0_port_1, alu0_v;
  wire signed [`W-1:0] alu1_port_3, alu1_port_0, alu1_port_1, alu1_port_4, alu1_v;
  wire signed [`W-1:0] alu2_port_3, alu2_port_0, alu2_port_1, alu2_port_4, alu2_v;
  wire signed [`W-1:0] alu3_port_2, alu3_port_3, alu3_port_0, alu3_port_1, alu3_v;
  wire signed [`W-1:0] _ABL4_port_3, _ABL4_port_1, _ABL4_v;
  wire signed [`W-1:0] n_488_port_2, n_488_port_3, n_488_port_0, n_488_port_1, n_488_port_4, n_488_v;
  wire signed [`W-1:0] n_481_port_2, n_481_port_3, n_481_port_0, n_481_port_1, n_481_port_4, n_481_v;
  wire signed [`W-1:0] n_326_port_2, n_326_port_3, n_326_port_0, n_326_port_1, n_326_port_4, n_326_v;
  wire signed [`W-1:0] n_1105_port_2, n_1105_port_0, n_1105_v;
  wire signed [`W-1:0] n_1100_port_2, n_1100_port_3, n_1100_port_0, n_1100_v;
  wire signed [`W-1:0] dpc6_SBS_port_11, dpc6_SBS_port_12, dpc6_SBS_v;
  wire signed [`W-1:0] n_831_port_2, n_831_port_3, n_831_port_0, n_831_port_1, n_831_port_4, n_831_v;
  wire signed [`W-1:0] s3_port_0, s3_port_1, s3_v;
  wire signed [`W-1:0] s2_port_0, s2_port_1, s2_v;
  wire signed [`W-1:0] s1_port_0, s1_port_1, s1_v;
  wire signed [`W-1:0] s0_port_0, s0_port_1, s0_v;
  wire signed [`W-1:0] s7_port_2, s7_port_0, s7_v;
  wire signed [`W-1:0] s6_port_0, s6_port_1, s6_v;
  wire signed [`W-1:0] s5_port_0, s5_port_1, s5_v;
  wire signed [`W-1:0] s4_port_0, s4_port_1, s4_v;
  wire signed [`W-1:0] so_port_2, so_port_3, so_v;
  wire signed [`W-1:0] dpc15_ANDS_port_9, dpc15_ANDS_port_0, dpc15_ANDS_v;
  wire signed [`W-1:0] dpc27_SBADH_port_9, dpc27_SBADH_port_0, dpc27_SBADH_v;
  wire signed [`W-1:0] n_649_port_0, n_649_port_7, n_649_port_5, n_649_v;
  wire signed [`W-1:0] n_138_port_2, n_138_port_0, n_138_port_1, n_138_v;
  wire signed [`W-1:0] n_642_port_3, n_642_port_0, n_642_port_1, n_642_v;
  wire signed [`W-1:0] n_643_port_3, n_643_port_4, n_643_v;
  wire signed [`W-1:0] n_1632_port_7, n_1632_port_4, n_1632_port_5, n_1632_v;
  wire signed [`W-1:0] n_583_port_2, n_583_port_0, n_583_port_1, n_583_v;
  wire signed [`W-1:0] notir0_port_0, notir0_port_1, notir0_port_28, notir0_v;
  wire signed [`W-1:0] notir1_port_21, notir1_port_23, notir1_port_22, notir1_v;
  wire signed [`W-1:0] notir2_port_19, notir2_port_0, notir2_port_20, notir2_v;
  wire signed [`W-1:0] notir3_port_51, notir3_port_0, notir3_port_1, notir3_v;
  wire signed [`W-1:0] notir4_port_25, notir4_port_24, notir4_port_26, notir4_v;
  wire signed [`W-1:0] notir5_port_36, notir5_port_37, notir5_port_0, notir5_v;
  wire signed [`W-1:0] notir6_port_39, notir6_port_0, notir6_port_1, notir6_v;
  wire signed [`W-1:0] notir7_port_33, notir7_port_34, notir7_port_35, notir7_v;
  wire signed [`W-1:0] n_119_port_3, n_119_port_0, n_119_v;
  wire signed [`W-1:0] cp1_port_75, cp1_port_50, cp1_v;
  wire signed [`W-1:0] a3_port_0, a3_port_1, a3_v;
  wire signed [`W-1:0] a6_port_2, a6_port_0, a6_v;
  wire signed [`W-1:0] n_1479_port_0, n_1479_port_1, n_1479_v;
  wire signed [`W-1:0] sync_port_0, sync_port_1, sync_v;
  wire signed [`W-1:0] n_1325_port_2, n_1325_port_4, n_1325_v;
  wire signed [`W-1:0] n_1496_port_2, n_1496_port_3, n_1496_port_0, n_1496_port_1, n_1496_port_4, n_1496_v;
  wire signed [`W-1:0] n_564_port_2, n_564_port_3, n_564_port_0, n_564_port_1, n_564_v;
  wire signed [`W-1:0] __AxBxC_6_port_3, __AxBxC_6_port_1, __AxBxC_6_port_5, __AxBxC_6_v;
  wire signed [`W-1:0] __AxBxC_7_port_3, __AxBxC_7_port_0, __AxBxC_7_port_5, __AxBxC_7_v;
  wire signed [`W-1:0] __AxBxC_4_port_2, __AxBxC_4_port_3, __AxBxC_4_port_5, __AxBxC_4_v;
  wire signed [`W-1:0] __AxBxC_5_port_3, __AxBxC_5_port_1, __AxBxC_5_port_5, __AxBxC_5_v;
  wire signed [`W-1:0] __AxBxC_2_port_3, __AxBxC_2_port_1, __AxBxC_2_port_5, __AxBxC_2_v;
  wire signed [`W-1:0] __AxBxC_3_port_3, __AxBxC_3_port_1, __AxBxC_3_port_5, __AxBxC_3_v;
  wire signed [`W-1:0] __AxBxC_0_port_2, __AxBxC_0_port_3, __AxBxC_0_port_5, __AxBxC_0_v;
  wire signed [`W-1:0] __AxBxC_1_port_3, __AxBxC_1_port_1, __AxBxC_1_port_5, __AxBxC_1_v;
  wire signed [`W-1:0] n_304_port_2, n_304_port_3, n_304_port_0, n_304_port_1, n_304_port_4, n_304_v;
  wire signed [`W-1:0] ab12_port_0, ab12_port_1, ab12_v;
  wire signed [`W-1:0] ab13_port_0, ab13_port_1, ab13_v;
  wire signed [`W-1:0] ab10_port_0, ab10_port_1, ab10_v;
  wire signed [`W-1:0] ab11_port_0, ab11_port_1, ab11_v;
  wire signed [`W-1:0] ab14_port_0, ab14_port_1, ab14_v;
  wire signed [`W-1:0] ab15_port_0, ab15_port_1, ab15_v;
  wire signed [`W-1:0] n_72_port_2, n_72_port_3, n_72_port_0, n_72_port_1, n_72_port_4, n_72_v;
  wire signed [`W-1:0] n_177_port_2, n_177_port_0, n_177_port_1, n_177_v;
  wire signed [`W-1:0] n_794_port_1, n_794_port_4, n_794_v;
  wire signed [`W-1:0] n_798_port_1, n_798_port_4, n_798_v;
  wire signed [`W-1:0] n_1301_port_2, n_1301_port_3, n_1301_port_0, n_1301_port_1, n_1301_port_4, n_1301_v;
  wire signed [`W-1:0] n_1300_port_2, n_1300_port_3, n_1300_v;
  wire signed [`W-1:0] n_1309_port_2, n_1309_port_3, n_1309_port_1, n_1309_v;
  wire signed [`W-1:0] n_330_port_7, n_330_port_4, n_330_v;
  wire signed [`W-1:0] n_332_port_2, n_332_port_3, n_332_port_0, n_332_port_1, n_332_port_4, n_332_v;
  wire signed [`W-1:0] n_1169_port_2, n_1169_port_3, n_1169_port_0, n_1169_port_1, n_1169_v;
  wire signed [`W-1:0] n_541_port_3, n_541_port_1, n_541_v;
  wire signed [`W-1:0] n_322_port_2, n_322_port_1, n_322_v;
  wire signed [`W-1:0] dpc24_ACSB_port_1, dpc24_ACSB_port_12, dpc24_ACSB_v;
  wire signed [`W-1:0] rdy_port_2, rdy_port_3, rdy_v;
  wire signed [`W-1:0] n_520_port_0, n_520_port_4, n_520_v;
  wire signed [`W-1:0] dpc21_ADDADL_port_9, dpc21_ADDADL_port_0, dpc21_ADDADL_v;
  wire signed [`W-1:0] n_1592_port_2, n_1592_port_3, n_1592_port_0, n_1592_port_1, n_1592_port_4, n_1592_v;
  wire signed [`W-1:0] n_37_port_3, n_37_port_4, n_37_v;
  wire signed [`W-1:0] db1_port_1, db1_port_4, db1_port_5, db1_v;
  wire signed [`W-1:0] db0_port_1, db0_port_4, db0_port_5, db0_v;
  wire signed [`W-1:0] db3_port_2, db3_port_3, db3_port_5, db3_v;
  wire signed [`W-1:0] db2_port_2, db2_port_3, db2_port_5, db2_v;
  wire signed [`W-1:0] db5_port_0, db5_port_4, db5_port_5, db5_v;
  wire signed [`W-1:0] db4_port_3, db4_port_0, db4_port_5, db4_v;
  wire signed [`W-1:0] db7_port_3, db7_port_1, db7_port_5, db7_v;
  wire signed [`W-1:0] db6_port_0, db6_port_4, db6_port_5, db6_v;
  wire signed [`W-1:0] clk1out_port_0, clk1out_port_1, clk1out_v;
  wire signed [`W-1:0] n_1647_port_2, n_1647_port_3, n_1647_port_0, n_1647_port_1, n_1647_port_4, n_1647_v;
  wire signed [`W-1:0] n_1641_port_2, n_1641_port_3, n_1641_port_1, n_1641_v;
  wire signed [`W-1:0] n_1491_port_2, n_1491_port_3, n_1491_port_0, n_1491_port_1, n_1491_v;
  wire signed [`W-1:0] n_206_port_3, n_206_port_0, n_206_port_5, n_206_v;
  wire signed [`W-1:0] clock1_port_40, clock1_port_68, clock1_v;
  wire signed [`W-1:0] n_1344_port_2, n_1344_port_3, n_1344_port_0, n_1344_port_1, n_1344_port_4, n_1344_v;
  wire signed [`W-1:0] n_1084_port_0, n_1084_port_6, n_1084_port_5, n_1084_v;
  wire signed [`W-1:0] n_1083_port_1, n_1083_port_7, n_1083_port_4, n_1083_v;
  wire signed [`W-1:0] n_1661_port_2, n_1661_port_3, n_1661_port_0, n_1661_port_1, n_1661_v;
  wire signed [`W-1:0] n_1668_port_2, n_1668_port_3, n_1668_port_0, n_1668_v;
  wire signed [`W-1:0] dpc32_PCHADH_port_0, dpc32_PCHADH_port_1, dpc32_PCHADH_v;
  wire signed [`W-1:0] idb1_port_8, idb1_port_9, idb1_port_3, idb1_port_0, idb1_port_7, idb1_port_4, idb1_port_5, idb1_port_10, idb1_v;
  wire signed [`W-1:0] idb0_port_8, idb0_port_2, idb0_port_1, idb0_port_6, idb0_port_7, idb0_port_4, idb0_port_5, idb0_port_10, idb0_v;
  wire signed [`W-1:0] idb3_port_8, idb3_port_9, idb3_port_3, idb3_port_0, idb3_port_1, idb3_port_6, idb3_port_5, idb3_port_10, idb3_v;
  wire signed [`W-1:0] idb2_port_9, idb2_port_3, idb2_port_0, idb2_port_1, idb2_port_6, idb2_port_4, idb2_port_5, idb2_port_10, idb2_v;
  wire signed [`W-1:0] idb5_port_8, idb5_port_9, idb5_port_2, idb5_port_6, idb5_port_7, idb5_port_4, idb5_port_5, idb5_v;
  wire signed [`W-1:0] idb4_port_8, idb4_port_9, idb4_port_0, idb4_port_6, idb4_port_7, idb4_port_4, idb4_port_5, idb4_port_10, idb4_v;
  wire signed [`W-1:0] idb7_port_8, idb7_port_9, idb7_port_2, idb7_port_3, idb7_port_0, idb7_port_7, idb7_port_4, idb7_port_10, idb7_v;
  wire signed [`W-1:0] idb6_port_9, idb6_port_3, idb6_port_0, idb6_port_6, idb6_port_7, idb6_port_5, idb6_port_10, idb6_port_11, idb6_v;
  wire signed [`W-1:0] n_1417_port_2, n_1417_port_0, n_1417_v;
  wire signed [`W-1:0] n_381_port_2, n_381_port_3, n_381_port_1, n_381_v;
  wire signed [`W-1:0] n_927_port_3, n_927_port_1, n_927_v;
  wire signed [`W-1:0] n_928_port_2, n_928_port_3, n_928_port_1, n_928_v;
  wire signed [`W-1:0] alub2_port_0, alub2_port_1, alub2_port_4, alub2_v;
  wire signed [`W-1:0] pch7_port_2, pch7_port_1, pch7_v;
  wire signed [`W-1:0] pch6_port_2, pch6_port_0, pch6_v;
  wire signed [`W-1:0] pch5_port_2, pch5_port_0, pch5_v;
  wire signed [`W-1:0] pch4_port_2, pch4_port_1, pch4_v;
  wire signed [`W-1:0] pch3_port_2, pch3_port_1, pch3_v;
  wire signed [`W-1:0] pch2_port_0, pch2_port_1, pch2_v;
  wire signed [`W-1:0] pch1_port_2, pch1_port_1, pch1_v;
  wire signed [`W-1:0] pch0_port_2, pch0_port_1, pch0_v;
  wire signed [`W-1:0] dpc13_ORS_port_8, dpc13_ORS_port_5, dpc13_ORS_v;
  wire signed [`W-1:0] n_1063_port_2, n_1063_port_7, n_1063_port_4, n_1063_port_5, n_1063_v;
  wire signed [`W-1:0] n_1608_port_2, n_1608_port_1, n_1608_v;
  wire signed [`W-1:0] n_1609_port_3, n_1609_port_0, n_1609_v;
  wire signed [`W-1:0] n_1605_port_3, n_1605_port_0, n_1605_port_5, n_1605_v;
  wire signed [`W-1:0] n_719_port_2, n_719_port_3, n_719_port_0, n_719_port_1, n_719_v;
  wire signed [`W-1:0] n_242_port_2, n_242_port_3, n_242_port_0, n_242_port_1, n_242_v;
  wire signed [`W-1:0] dasb7_port_3, dasb7_port_1, dasb7_port_5, dasb7_v;
  wire signed [`W-1:0] n_1296_port_2, n_1296_port_0, n_1296_v;
  wire signed [`W-1:0] dpc7_SS_port_7, dpc7_SS_port_12, dpc7_SS_v;
  wire signed [`W-1:0] n_1041_port_0, n_1041_port_1, n_1041_v;
  wire signed [`W-1:0] n_1046_port_2, n_1046_port_3, n_1046_port_0, n_1046_v;
  wire signed [`W-1:0] n_1620_port_3, n_1620_port_0, n_1620_v;
  wire signed [`W-1:0] n_1621_port_2, n_1621_port_0, n_1621_port_1, n_1621_v;
  wire signed [`W-1:0] n_227_port_2, n_227_port_3, n_227_port_0, n_227_v;
  wire signed [`W-1:0] x2_port_0, x2_port_1, x2_v;
  wire signed [`W-1:0] x3_port_0, x3_port_1, x3_v;
  wire signed [`W-1:0] x0_port_0, x0_port_1, x0_v;
  wire signed [`W-1:0] x1_port_0, x1_port_1, x1_v;
  wire signed [`W-1:0] x7_port_2, x7_port_1, x7_v;
  wire signed [`W-1:0] x4_port_0, x4_port_1, x4_v;
  wire signed [`W-1:0] x5_port_2, x5_port_1, x5_v;
  wire signed [`W-1:0] n_1458_port_2, n_1458_port_3, n_1458_port_0, n_1458_port_1, n_1458_port_4, n_1458_v;
  wire signed [`W-1:0] n_694_port_2, n_694_port_3, n_694_port_0, n_694_port_1, n_694_port_4, n_694_v;
  wire signed [`W-1:0] n_963_port_2, n_963_port_1, n_963_v;
  wire signed [`W-1:0] pcl3_port_2, pcl3_port_1, pcl3_v;
  wire signed [`W-1:0] pcl2_port_2, pcl2_port_1, pcl2_v;
  wire signed [`W-1:0] pcl1_port_2, pcl1_port_1, pcl1_v;
  wire signed [`W-1:0] pcl0_port_2, pcl0_port_1, pcl0_v;
  wire signed [`W-1:0] pcl7_port_2, pcl7_port_1, pcl7_v;
  wire signed [`W-1:0] pcl6_port_2, pcl6_port_1, pcl6_v;
  wire signed [`W-1:0] pcl5_port_2, pcl5_port_1, pcl5_v;
  wire signed [`W-1:0] pcl4_port_2, pcl4_port_1, pcl4_v;
  wire signed [`W-1:0] dpc0_YSB_port_3, dpc0_YSB_port_12, dpc0_YSB_v;
  wire signed [`W-1:0] alua6_port_0, alua6_port_1, alua6_v;
  wire signed [`W-1:0] alua7_port_3, alua7_port_0, alua7_v;
  wire signed [`W-1:0] alua4_port_0, alua4_port_1, alua4_v;
  wire signed [`W-1:0] alua5_port_0, alua5_port_1, alua5_v;
  wire signed [`W-1:0] alua2_port_0, alua2_port_1, alua2_v;
  wire signed [`W-1:0] alua3_port_0, alua3_port_1, alua3_v;
  wire signed [`W-1:0] alua0_port_0, alua0_port_1, alua0_v;
  wire signed [`W-1:0] alua1_port_2, alua1_port_3, alua1_v;
  wire signed [`W-1:0] nmi_port_2, nmi_v;
  wire signed [`W-1:0] dpc41_DL_ADL_port_9, dpc41_DL_ADL_port_0, dpc41_DL_ADL_v;
  wire signed [`W-1:0] n_208_port_2, n_208_port_3, n_208_port_0, n_208_port_1, n_208_port_4, n_208_v;
  wire signed [`W-1:0] n_209_port_2, n_209_port_3, n_209_port_0, n_209_port_1, n_209_port_4, n_209_v;
  wire signed [`W-1:0] dpc37_PCLDB_port_0, dpc37_PCLDB_port_4, dpc37_PCLDB_v;
  wire signed [`W-1:0] dpc12_0ADD_port_9, dpc12_0ADD_port_12, dpc12_0ADD_v;
  wire signed [`W-1:0] dpc4_SSB_port_9, dpc4_SSB_port_0, dpc4_SSB_v;
  wire signed [`W-1:0] n_417_port_0, n_417_port_1, n_417_v;
  wire signed [`W-1:0] y1_port_2, y1_port_0, y1_v;
  wire signed [`W-1:0] y0_port_2, y0_port_0, y0_v;
  wire signed [`W-1:0] y3_port_2, y3_port_0, y3_v;
  wire signed [`W-1:0] y2_port_2, y2_port_0, y2_v;
  wire signed [`W-1:0] y5_port_0, y5_port_1, y5_v;
  wire signed [`W-1:0] y4_port_2, y4_port_0, y4_v;
  wire signed [`W-1:0] y7_port_0, y7_port_1, y7_v;
  wire signed [`W-1:0] y6_port_0, y6_port_1, y6_v;
  wire signed [`W-1:0] dpc11_SBADD_port_9, dpc11_SBADD_port_12, dpc11_SBADD_v;
  wire signed [`W-1:0] dpc10_ADLADD_port_5, dpc10_ADLADD_port_12, dpc10_ADLADD_v;
  wire signed [`W-1:0] dpc29_0ADH17_port_2, dpc29_0ADH17_port_1, dpc29_0ADH17_v;
  wire signed [`W-1:0] dpc26_ACDB_port_0, dpc26_ACDB_port_12, dpc26_ACDB_v;
  wire signed [`W-1:0] n_430_port_2, n_430_port_3, n_430_port_1, n_430_v;
  wire signed [`W-1:0] n_436_port_2, n_436_port_3, n_436_port_0, n_436_port_1, n_436_v;
  wire signed [`W-1:0] n_404_port_2, n_404_port_6, n_404_port_5, n_404_v;
  wire signed [`W-1:0] n_1654_port_2, n_1654_port_3, n_1654_port_0, n_1654_port_1, n_1654_port_4, n_1654_v;
  wire signed [`W-1:0] n_635_port_3, n_635_port_0, n_635_port_1, n_635_v;
  wire signed [`W-1:0] n_634_port_0, n_634_port_1, n_634_v;
  wire signed [`W-1:0] n_633_port_0, n_633_v;
  wire signed [`W-1:0] n_458_port_2, n_458_port_0, n_458_port_1, n_458_v;
  wire signed [`W-1:0] n_1519_port_2, n_1519_port_3, n_1519_port_0, n_1519_v;
  wire signed [`W-1:0] dpc16_EORS_port_8, dpc16_EORS_port_9, dpc16_EORS_v;
  wire signed [`W-1:0] n_1722_port_2, n_1722_port_3, n_1722_port_0, n_1722_port_1, n_1722_port_4, n_1722_v;
  wire signed [`W-1:0] n_618_port_2, n_618_port_3, n_618_port_0, n_618_port_1, n_618_port_4, n_618_v;
  wire signed [`W-1:0] n_612_port_0, n_612_port_4, n_612_v;
  wire signed [`W-1:0] n_884_port_2, n_884_port_0, n_884_port_1, n_884_v;
  wire signed [`W-1:0] Pout0_port_2, Pout0_port_0, Pout0_port_1, Pout0_v;
  wire signed [`W-1:0] n_1545_port_2, n_1545_port_1, n_1545_v;
  wire signed [`W-1:0] dpc19_ADDSB7_port_2, dpc19_ADDSB7_port_0, dpc19_ADDSB7_v;
  wire signed [`W-1:0] n_477_port_3, n_477_port_1, n_477_port_4, n_477_port_5, n_477_v;
  wire signed [`W-1:0] n_475_port_2, n_475_port_0, n_475_v;
  wire signed [`W-1:0] n_471_port_3, n_471_port_4, n_471_v;
  wire signed [`W-1:0] n_478_port_2, n_478_port_0, n_478_port_1, n_478_v;
  wire signed [`W-1:0] p6_port_2, p6_port_0, p6_port_1, p6_v;
  wire signed [`W-1:0] p7_port_2, p7_port_0, p7_port_1, p7_v;
  wire signed [`W-1:0] n_1531_port_2, n_1531_port_3, n_1531_port_0, n_1531_port_1, n_1531_v;
  wire signed [`W-1:0] n_1398_port_8, n_1398_port_1, n_1398_port_6, n_1398_v;
  wire signed [`W-1:0] n_280_port_2, n_280_port_3, n_280_port_0, n_280_port_1, n_280_port_4, n_280_v;
  wire signed [`W-1:0] n_135_port_2, n_135_port_1, n_135_v;
  wire signed [`W-1:0] n_869_port_2, n_869_port_3, n_869_port_1, n_869_v;
  wire signed [`W-1:0] n_866_v;
  wire signed [`W-1:0] n_350_port_3, n_350_port_1, n_350_port_4, n_350_port_5, n_350_v;
  wire signed [`W-1:0] dpc17_SUMS_port_0, dpc17_SUMS_port_1, dpc17_SUMS_v;
  wire signed [`W-1:0] n_1251_port_2, n_1251_port_3, n_1251_port_0, n_1251_port_1, n_1251_v;
  wire signed [`W-1:0] n_1709_port_2, n_1709_port_3, n_1709_port_0, n_1709_port_1, n_1709_v;
  wire signed [`W-1:0] dpc3_SBX_port_9, dpc3_SBX_port_12, dpc3_SBX_v;
  wire signed [`W-1:0] dpc31_PCHPCH_port_11, dpc31_PCHPCH_port_12, dpc31_PCHPCH_v;
  wire signed [`W-1:0] n_676_port_2, n_676_port_3, n_676_port_0, n_676_v;
  wire signed [`W-1:0] Pout1_port_2, Pout1_port_0, Pout1_port_1, Pout1_v;
  wire signed [`W-1:0] Pout3_port_2, Pout3_port_3, Pout3_port_4, Pout3_v;
  wire signed [`W-1:0] Pout2_port_2, Pout2_port_0, Pout2_port_1, Pout2_v;
  wire signed [`W-1:0] n_494_port_2, n_494_port_3, n_494_port_1, n_494_v;
  wire signed [`W-1:0] n_806_v;
  wire signed [`W-1:0] n_807_port_3, n_807_port_5, n_807_v;
  wire signed [`W-1:0] n_659_port_2, n_659_port_3, n_659_port_1, n_659_v;
  wire signed [`W-1:0] n_658_port_2, n_658_port_3, n_658_port_0, n_658_port_1, n_658_v;
  wire signed [`W-1:0] n_652_port_2, n_652_port_3, n_652_port_0, n_652_port_1, n_652_port_4, n_652_v;
  wire signed [`W-1:0] n_123_port_2, n_123_port_3, n_123_port_0, n_123_v;
  wire signed [`W-1:0] n_826_port_2, n_826_port_1, n_826_v;
  wire signed [`W-1:0] n_351_port_2, n_351_port_0, n_351_port_1, n_351_v;
  wire signed [`W-1:0] dpc9_DBADD_port_1, dpc9_DBADD_port_12, dpc9_DBADD_v;
  wire signed [`W-1:0] n_359_port_2, n_359_port_0, n_359_port_1, n_359_v;
  wire signed [`W-1:0] dpc33_PCHDB_port_0, dpc33_PCHDB_port_1, dpc33_PCHDB_v;
  wire signed [`W-1:0] dpc8_nDBADD_port_6, dpc8_nDBADD_port_12, dpc8_nDBADD_v;
  wire signed [`W-1:0] n_102_port_2, n_102_port_0, n_102_v;
  wire signed [`W-1:0] dpc39_PCLPCL_port_11, dpc39_PCLPCL_port_12, dpc39_PCLPCL_v;
  wire signed [`W-1:0] ADH_ABH_port_7, ADH_ABH_port_4, ADH_ABH_v;
  wire signed [`W-1:0] dpc25_SBDB_port_9, dpc25_SBDB_port_0, dpc25_SBDB_v;
  wire signed [`W-1:0] dpc23_SBAC_port_11, dpc23_SBAC_port_12, dpc23_SBAC_v;
  wire signed [`W-1:0] n_1152_port_2, n_1152_port_0, n_1152_v;
  wire signed [`W-1:0] n_373_port_0, n_373_port_4, n_373_v;
  wire signed [`W-1:0] ab0_port_0, ab0_port_1, ab0_v;
  wire signed [`W-1:0] ab1_port_0, ab1_port_1, ab1_v;
  wire signed [`W-1:0] ab2_port_0, ab2_port_1, ab2_v;
  wire signed [`W-1:0] ab3_port_0, ab3_port_1, ab3_v;
  wire signed [`W-1:0] ab4_port_0, ab4_port_1, ab4_v;
  wire signed [`W-1:0] ab5_port_0, ab5_port_1, ab5_v;
  wire signed [`W-1:0] ab6_port_0, ab6_port_1, ab6_v;
  wire signed [`W-1:0] ab7_port_0, ab7_port_1, ab7_v;
  wire signed [`W-1:0] ab8_port_0, ab8_port_1, ab8_v;
  wire signed [`W-1:0] ab9_port_0, ab9_port_1, ab9_v;
  wire signed [`W-1:0] n_87_port_2, n_87_port_3, n_87_port_0, n_87_port_1, n_87_v;
  wire signed [`W-1:0] n_86_port_2, n_86_port_3, n_86_port_0, n_86_v;
  wire signed [`W-1:0] n_168_port_2, n_168_port_3, n_168_port_0, n_168_v;
  wire signed [`W-1:0] sb2_port_8, sb2_port_9, sb2_port_2, sb2_port_3, sb2_port_0, sb2_port_1, sb2_port_6, sb2_port_7, sb2_port_4, sb2_port_10, sb2_port_11, sb2_port_12, sb2_v;
  wire signed [`W-1:0] sb3_port_8, sb3_port_9, sb3_port_2, sb3_port_3, sb3_port_0, sb3_port_1, sb3_port_6, sb3_port_7, sb3_port_4, sb3_port_5, sb3_port_10, sb3_port_11, sb3_v;
  wire signed [`W-1:0] sb0_port_8, sb0_port_9, sb0_port_2, sb0_port_3, sb0_port_0, sb0_port_1, sb0_port_6, sb0_port_7, sb0_port_4, sb0_port_5, sb0_port_10, sb0_port_11, sb0_port_12, sb0_v;
  wire signed [`W-1:0] sb1_port_8, sb1_port_9, sb1_port_2, sb1_port_0, sb1_port_1, sb1_port_6, sb1_port_7, sb1_port_4, sb1_port_5, sb1_port_10, sb1_port_11, sb1_port_12, sb1_v;
  wire signed [`W-1:0] sb6_port_8, sb6_port_9, sb6_port_2, sb6_port_3, sb6_port_0, sb6_port_1, sb6_port_6, sb6_port_7, sb6_port_4, sb6_port_10, sb6_port_11, sb6_port_12, sb6_v;
  wire signed [`W-1:0] sb7_port_8, sb7_port_9, sb7_port_2, sb7_port_3, sb7_port_0, sb7_port_1, sb7_port_6, sb7_port_7, sb7_port_4, sb7_port_5, sb7_port_10, sb7_port_11, sb7_v;
  wire signed [`W-1:0] sb4_port_8, sb4_port_9, sb4_port_2, sb4_port_3, sb4_port_0, sb4_port_1, sb4_port_6, sb4_port_7, sb4_port_4, sb4_port_5, sb4_port_10, sb4_port_11, sb4_port_12, sb4_v;
  wire signed [`W-1:0] sb5_port_8, sb5_port_2, sb5_port_3, sb5_port_0, sb5_port_1, sb5_port_6, sb5_port_7, sb5_port_4, sb5_port_5, sb5_port_10, sb5_port_11, sb5_port_12, sb5_v;
  wire signed [`W-1:0] __AxB_6_port_2, __AxB_6_port_6, __AxB_6_port_11, __AxB_6_v;
  wire signed [`W-1:0] __AxB_4_port_0, __AxB_4_port_6, __AxB_4_port_4, __AxB_4_v;
  wire signed [`W-1:0] __AxB_2_port_0, __AxB_2_port_7, __AxB_2_port_4, __AxB_2_v;
  wire signed [`W-1:0] __AxB_0_port_2, __AxB_0_port_6, __AxB_0_port_4, __AxB_0_v;
  wire signed [`W-1:0] n_1318_port_2, n_1318_port_3, n_1318_port_7, n_1318_port_5, n_1318_v;
  wire signed [`W-1:0] dpc2_XSB_port_2, dpc2_XSB_port_12, dpc2_XSB_v;
  wire signed [`W-1:0] n_578_port_2, n_578_port_3, n_578_port_0, n_578_port_1, n_578_v;
  wire signed [`W-1:0] n_571_port_2, n_571_port_3, n_571_port_1, n_571_v;
  wire signed [`W-1:0] n_310_port_3, n_310_port_0, n_310_v;
  wire signed [`W-1:0] dpc14_SRS_port_2, dpc14_SRS_port_1, dpc14_SRS_v;
  wire signed [`W-1:0] n_66_port_2, n_66_port_3, n_66_port_1, n_66_v;
  wire signed [`W-1:0] n_147_port_3, n_147_port_4, n_147_v;
  wire signed [`W-1:0] n_146_port_2, n_146_port_3, n_146_port_0, n_146_port_1, n_146_port_4, n_146_v;
  wire signed [`W-1:0] n_141_port_2, n_141_port_3, n_141_port_0, n_141_port_1, n_141_port_4, n_141_v;
  wire signed [`W-1:0] ADL_ABL_port_0, ADL_ABL_port_5, ADL_ABL_v;
  wire signed [`W-1:0] n_1724_port_2, n_1724_port_3, n_1724_port_0, n_1724_port_1, n_1724_v;
  wire signed [`W-1:0] n_1191_port_2, n_1191_port_0, n_1191_v;
  wire signed [`W-1:0] n_883_port_2, n_883_port_3, n_883_port_1, n_883_v;
  wire signed [`W-1:0] n_880_port_2, n_880_port_3, n_880_port_0, n_880_v;
  wire signed [`W-1:0] n_336_port_3, n_336_port_1, n_336_port_6, n_336_port_7, n_336_v;
  wire signed [`W-1:0] n_43_port_11, n_43_port_13, n_43_v;
  wire signed [`W-1:0] n_42_port_0, n_42_port_4, n_42_v;
  wire signed [`W-1:0] res_port_2, res_v;
  wire signed [`W-1:0] adl7_port_2, adl7_port_3, adl7_port_0, adl7_port_6, adl7_port_7, adl7_port_4, adl7_port_5, adl7_v;
  wire signed [`W-1:0] adl6_port_2, adl6_port_3, adl6_port_1, adl6_port_6, adl6_port_7, adl6_port_4, adl6_port_5, adl6_v;
  wire signed [`W-1:0] adl5_port_2, adl5_port_3, adl5_port_0, adl5_port_1, adl5_port_7, adl5_port_4, adl5_port_5, adl5_v;
  wire signed [`W-1:0] adl4_port_3, adl4_port_0, adl4_port_1, adl4_port_6, adl4_port_7, adl4_port_4, adl4_port_5, adl4_v;
  wire signed [`W-1:0] adl3_port_2, adl3_port_3, adl3_port_0, adl3_port_1, adl3_port_6, adl3_port_7, adl3_port_4, adl3_v;
  wire signed [`W-1:0] adl2_port_8, adl2_port_2, adl2_port_3, adl2_port_0, adl2_port_1, adl2_port_6, adl2_port_4, adl2_port_5, adl2_v;
  wire signed [`W-1:0] adl1_port_8, adl1_port_2, adl1_port_3, adl1_port_0, adl1_port_1, adl1_port_7, adl1_port_4, adl1_port_5, adl1_v;
  wire signed [`W-1:0] adl0_port_8, adl0_port_3, adl0_port_0, adl0_port_1, adl0_port_6, adl0_port_7, adl0_port_4, adl0_port_5, adl0_v;
  wire signed [`W-1:0] n_1014_port_2, n_1014_port_3, n_1014_port_0, n_1014_port_1, n_1014_v;
  wire signed [`W-1:0] dpc40_ADLPCL_port_0, dpc40_ADLPCL_port_12, dpc40_ADLPCL_v;
  wire signed [`W-1:0] n_929_port_2, n_929_port_3, n_929_port_0, n_929_port_1, n_929_port_4, n_929_v;
  wire signed [`W-1:0] n_1424_port_2, n_1424_port_3, n_1424_port_0, n_1424_port_1, n_1424_v;
  wire signed [`W-1:0] notaluoutmux0_port_2, notaluoutmux0_port_3, notaluoutmux0_port_0, notaluoutmux0_port_1, notaluoutmux0_port_5, notaluoutmux0_v;
  wire signed [`W-1:0] notaluoutmux1_port_2, notaluoutmux1_port_0, notaluoutmux1_port_1, notaluoutmux1_port_4, notaluoutmux1_port_5, notaluoutmux1_v;
  wire signed [`W-1:0] dpc30_ADHPCH_port_10, dpc30_ADHPCH_port_12, dpc30_ADHPCH_v;
  wire signed [`W-1:0] dpc43_DL_DB_port_9, dpc43_DL_DB_port_0, dpc43_DL_DB_v;
  wire signed [`W-1:0] n_27_port_2, n_27_port_3, n_27_port_0, n_27_port_1, n_27_port_4, n_27_v;
  wire signed [`W-1:0] aluanorb0_port_1, aluanorb0_port_6, aluanorb0_port_7, aluanorb0_v;
  wire signed [`W-1:0] n_1694_port_2, n_1694_port_3, n_1694_port_0, n_1694_port_1, n_1694_v;
  wire signed [`W-1:0] a1_port_0, a1_port_1, a1_v;
  wire signed [`W-1:0] a0_port_0, a0_port_1, a0_v;
  wire signed [`W-1:0] a2_port_2, a2_port_1, a2_v;
  wire signed [`W-1:0] a5_port_2, a5_port_0, a5_v;
  wire signed [`W-1:0] a4_port_2, a4_port_0, a4_v;
  wire signed [`W-1:0] a7_port_2, a7_port_1, a7_v;
  wire signed [`W-1:0] n_277_port_2, n_277_port_3, n_277_port_1, n_277_port_4, n_277_port_5, n_277_v;
  wire signed [`W-1:0] n_518_port_2, n_518_port_3, n_518_port_0, n_518_port_1, n_518_v;
  wire signed [`W-1:0] n_1467_port_0, n_1467_port_1, n_1467_v;
  wire signed [`W-1:0] n_1095_port_2, n_1095_port_3, n_1095_port_0, n_1095_port_1, n_1095_v;
  wire signed [`W-1:0] n_1094_port_2, n_1094_port_3, n_1094_port_1, n_1094_v;
  wire signed [`W-1:0] n_1675_port_3, n_1675_port_0, n_1675_v;
  wire signed [`W-1:0] adh3_port_2, adh3_port_3, adh3_port_0, adh3_port_6, adh3_port_4, adh3_port_5, adh3_v;
  wire signed [`W-1:0] adh2_port_3, adh2_port_0, adh2_port_1, adh2_port_6, adh2_port_4, adh2_port_5, adh2_v;
  wire signed [`W-1:0] adh1_port_2, adh1_port_0, adh1_port_1, adh1_port_6, adh1_port_4, adh1_port_5, adh1_v;
  wire signed [`W-1:0] adh0_port_2, adh0_port_3, adh0_port_0, adh0_port_1, adh0_port_6, adh0_port_4, adh0_v;
  wire signed [`W-1:0] adh7_port_2, adh7_port_3, adh7_port_0, adh7_port_1, adh7_port_4, adh7_port_5, adh7_v;
  wire signed [`W-1:0] adh6_port_3, adh6_port_0, adh6_port_1, adh6_port_6, adh6_port_4, adh6_port_5, adh6_v;
  wire signed [`W-1:0] adh5_port_2, adh5_port_3, adh5_port_0, adh5_port_1, adh5_port_4, adh5_port_5, adh5_v;
  wire signed [`W-1:0] adh4_port_2, adh4_port_0, adh4_port_1, adh4_port_6, adh4_port_4, adh4_port_5, adh4_v;
  wire signed [`W-1:0] n_254_port_2, n_254_port_3, n_254_port_1, n_254_v;
  wire signed [`W-1:0] n_1469_port_2, n_1469_port_0, n_1469_port_1, n_1469_v;
  wire signed [`W-1:0] n_935_port_2, n_935_port_3, n_935_port_1, n_935_v;
  wire signed [`W-1:0] NMIP_port_7, NMIP_port_4, NMIP_v;
  wire signed [`W-1:0] n_1076_port_0, n_1076_port_4, n_1076_v;
  wire signed [`W-1:0] n_1071_port_2, n_1071_port_3, n_1071_port_0, n_1071_port_4, n_1071_port_5, n_1071_v;
  wire signed [`W-1:0] n_1072_port_2, n_1072_port_4, n_1072_v;
  wire signed [`W-1:0] n_1140_port_2, n_1140_port_1, n_1140_v;
  wire signed [`W-1:0] n_1147_port_2, n_1147_port_3, n_1147_port_0, n_1147_port_1, n_1147_v;
  wire signed [`W-1:0] aluanorb1_port_7, aluanorb1_port_4, aluanorb1_port_5, aluanorb1_v;
  wire signed [`W-1:0] n_723_port_2, n_723_port_3, n_723_port_0, n_723_port_1, n_723_port_4, n_723_v;
  wire signed [`W-1:0] n_722_port_2, n_722_port_0, n_722_port_1, n_722_port_4, n_722_port_5, n_722_v;
  wire signed [`W-1:0] n_721_port_2, n_721_port_3, n_721_port_0, n_721_port_1, n_721_port_4, n_721_v;
  wire signed [`W-1:0] dpc1_SBY_port_3, dpc1_SBY_port_12, dpc1_SBY_v;
  wire signed [`W-1:0] cclk_port_236, cclk_port_28, cclk_v;
  wire signed [`W-1:0] RnWstretched_port_23, RnWstretched_port_22, RnWstretched_v;
  wire signed [`W-1:0] n_1059_port_0, n_1059_v;
  wire signed [`W-1:0] n_1633_port_2, n_1633_port_0, n_1633_v;
  wire signed [`W-1:0] n_1639_port_2, n_1639_port_0, n_1639_v;
  wire signed [`W-1:0] n_740_port_2, n_740_port_3, n_740_port_0, n_740_port_1, n_740_port_4, n_740_v;
  wire signed [`W-1:0] n_212_port_2, n_212_port_3, n_212_port_1, n_212_v;
  wire signed [`W-1:0] n_210_port_3, n_210_port_0, n_210_port_1, n_210_v;
  wire signed [`W-1:0] notRdy0_port_3, notRdy0_port_4, notRdy0_v;
  wire signed [`W-1:0] n_624_port_2, n_624_port_0, n_624_port_1, n_624_v;
  wire signed [`W-1:0] clk2out_port_0, clk2out_port_1, clk2out_v;
  wire signed [`W-1:0] n_681_port_8, n_681_port_3, n_681_port_1, n_681_port_6, n_681_v;
  wire signed [`W-1:0] n_976_port_2, n_976_port_3, n_976_port_0, n_976_port_1, n_976_port_4, n_976_v;
  wire signed [`W-1:0] n_975_port_3, n_975_port_6, n_975_v;
  wire signed [`W-1:0] n_1618_port_2, n_1618_port_3, n_1618_port_0, n_1618_port_1, n_1618_port_4, n_1618_v;
  wire signed [`W-1:0] alub3_port_2, alub3_port_3, alub3_port_4, alub3_v;
  wire signed [`W-1:0] alub1_port_0, alub1_port_1, alub1_port_4, alub1_v;
  wire signed [`W-1:0] alub0_port_2, alub0_port_3, alub0_port_4, alub0_v;
  wire signed [`W-1:0] alub7_port_3, alub7_port_0, alub7_port_4, alub7_v;
  wire signed [`W-1:0] alub6_port_2, alub6_port_3, alub6_port_4, alub6_v;
  wire signed [`W-1:0] alub5_port_2, alub5_port_3, alub5_port_4, alub5_v;
  wire signed [`W-1:0] alub4_port_3, alub4_port_0, alub4_port_4, alub4_v;
  wire signed [`W-1:0] dpc42_DL_ADH_port_8, dpc42_DL_ADH_port_9, dpc42_DL_ADH_v;
  wire signed [`W-1:0] n_767_port_2, n_767_port_3, n_767_port_0, n_767_port_1, n_767_v;
  wire signed [`W-1:0] n_953_port_2, n_953_port_0, n_953_port_1, n_953_v;
  wire signed [`W-1:0] n_409_port_3, n_409_port_0, n_409_port_5, n_409_v;
  wire signed [`W-1:0] n_1548_port_2, n_1548_port_3, n_1548_port_1, n_1548_v;
  wire signed [`W-1:0] n_1016_port_2, n_1016_port_3, n_1016_port_1, n_1016_v;
  wire signed [`W-1:0] p4_port_2, p4_port_0, p4_port_1, p4_v;
  wire signed [`W-1:0] n_171_port_3, n_171_port_0, n_171_port_1, n_171_v;
  wire signed [`W-1:0] clk0_port_3, clk0_v;
  wire signed [`W-1:0] n_1206_port_2, n_1206_port_3, n_1206_port_0, n_1206_port_1, n_1206_port_4, n_1206_v;
  wire signed [`W-1:0] _ABH3_port_3, _ABH3_port_1, _ABH3_v;
  wire signed [`W-1:0] _ABH2_port_2, _ABH2_port_3, _ABH2_v;
  wire signed [`W-1:0] _ABH1_port_3, _ABH1_port_0, _ABH1_v;
  wire signed [`W-1:0] _ABH0_port_2, _ABH0_port_3, _ABH0_v;
  wire signed [`W-1:0] _ABH7_port_2, _ABH7_port_3, _ABH7_v;
  wire signed [`W-1:0] _ABH6_port_2, _ABH6_port_3, _ABH6_v;
  wire signed [`W-1:0] _ABH5_port_2, _ABH5_port_3, _ABH5_v;
  wire signed [`W-1:0] _ABH4_port_2, _ABH4_port_3, _ABH4_v;
  wire signed [`W-1:0] n_1507_port_2, n_1507_port_3, n_1507_port_1, n_1507_v;
  wire signed [`W-1:0] n_423_port_2, n_423_port_0, n_423_port_1, n_423_v;
  wire signed [`W-1:0] n_1254_port_2, n_1254_port_0, n_1254_port_1, n_1254_v;
  wire signed [`W-1:0] dpc18__DAA_port_2, dpc18__DAA_port_1, dpc18__DAA_v;
  wire signed [`W-1:0] dpc38_PCLADL_port_9, dpc38_PCLADL_port_0, dpc38_PCLADL_v;
  wire signed [`W-1:0] n_1691_port_8, n_1691_port_1, n_1691_port_7, n_1691_v;
  wire signed [`W-1:0] n_1696_port_0, n_1696_port_1, n_1696_v;
  wire signed [`W-1:0] n_855_port_2, n_855_port_0, n_855_v;
  wire signed [`W-1:0] n_854_port_6, n_854_port_4, n_854_v;
  wire signed [`W-1:0] n_994_port_2, n_994_port_3, n_994_port_1, n_994_v;
  wire signed [`W-1:0] n_998_port_2, n_998_port_3, n_998_port_0, n_998_port_1, n_998_port_4, n_998_v;
  wire signed [`W-1:0] n_999_port_2, n_999_port_3, n_999_port_1, n_999_v;
  wire signed [`W-1:0] n_1501_port_1, n_1501_port_4, n_1501_v;
  wire signed [`W-1:0] n_298_port_3, n_298_port_4, n_298_v;
  wire signed [`W-1:0] n_297_port_3, n_297_port_5, n_297_v;
  wire signed [`W-1:0] n_296_port_3, n_296_port_0, n_296_port_1, n_296_port_4, n_296_port_5, n_296_v;
  wire signed [`W-1:0] n_871_port_2, n_871_port_3, n_871_port_0, n_871_port_1, n_871_v;

  wire pipedpc28_v;
  wire dor5_v;
  wire dor4_v;
  wire dor7_v;
  wire dor6_v;
  wire dor1_v;
  wire dor0_v;
  wire dor3_v;
  wire dor2_v;
  wire _DBZ_v;
  wire _DBE_v;
  wire n_1714_v;
  wire n_1715_v;
  wire n_1716_v;
  wire n_1717_v;
  wire n_1244_v;
  wire n_1245_v;
  wire n_1718_v;
  wire n_1719_v;
  wire n_604_v;
  wire n_600_v;
  wire n_602_v;
  wire n_603_v;
  wire n_608_v;
  wire n_609_v;
  wire pd6_clearIR_v;
  wire n_460_v;
  wire n_462_v;
  wire n_466_v;
  wire n_467_v;
  wire n_468_v;
  wire n_469_v;
  wire op_T4_brk_v;
  wire n_1162_v;
  wire n_1161_v;
  wire x_op_T3_plp_pla_v;
  wire n_1529_v;
  wire n_1528_v;
  wire n_1523_v;
  wire n_1521_v;
  wire n_1527_v;
  wire n_1526_v;
  wire n_1386_v;
  wire n_1380_v;
  wire n_819_v;
  wire n_818_v;
  wire n_811_v;
  wire n_810_v;
  wire n_813_v;
  wire n_812_v;
  wire n_815_v;
  wire ir0_v;
  wire ir1_v;
  wire ir2_v;
  wire ir3_v;
  wire ir4_v;
  wire ir5_v;
  wire ir6_v;
  wire ir7_v;
  wire n_599_v;
  wire n_1260_v;
  wire op_T__inx_v;
  wire n_9_v;
  wire n_5_v;
  wire n_6_v;
  wire n_1240_v;
  wire n_1711_v;
  wire n_1712_v;
  wire op_T0_php_pha_v;
  wire n_662_v;
  wire n_663_v;
  wire n_666_v;
  wire n_664_v;
  wire n_484_v;
  wire n_485_v;
  wire n_480_v;
  wire PD_xxx010x1_v;
  wire op_shift_v;
  wire op_xy_v;
  wire op_T0_cld_sed_v;
  wire n_327_v;
  wire _AxB_0__C0in_v;
  wire n_321_v;
  wire n_320_v;
  wire n_1107_v;
  wire n_1106_v;
  wire n_1101_v;
  wire n_1109_v;
  wire pd4_clearIR_v;
  wire op_ror_v;
  wire n_345_v;
  wire n_347_v;
  wire n_340_v;
  wire n_830_v;
  wire n_839_v;
  wire n_838_v;
  wire op_T0_ldy_mem_v;
  wire D1x1_v;
  wire n_1585_v;
  wire n_1586_v;
  wire _TWOCYCLE_v;
  wire pd3_clearIR_v;
  wire n_1450_v;
  wire n_139_v;
  wire n_641_v;
  wire n_132_v;
  wire n_645_v;
  wire n_646_v;
  wire n_647_v;
  wire n_1635_v;
  wire _AxB_6__C56_v;
  wire pd0_clearIR_v;
  wire op_T0_shift_a_v;
  wire __AxB7__C67_v;
  wire n_1439_v;
  wire _VEC_v;
  wire n_1129_v;
  wire n_1126_v;
  wire n_1124_v;
  wire n_1121_v;
  wire n_1120_v;
  wire n_587_v;
  wire n_586_v;
  wire n_582_v;
  wire n_588_v;
  wire op_rmw_v;
  wire n_360_v;
  wire n_366_v;
  wire n_368_v;
  wire op_jmp_v;
  wire C12_v;
  wire n_1433_v;
  wire op_shift_right_v;
  wire op_EORS_v;
  wire x_op_T__adc_sbc_v;
  wire n_1631_v;
  wire n_94_v;
  wire n_95_v;
  wire n_93_v;
  wire n_90_v;
  wire n_91_v;
  wire op_lsr_ror_dec_inc_v;
  wire n_110_v;
  wire n_111_v;
  wire n_118_v;
  wire n_696_v;
  wire n_698_v;
  wire n_1199_v;
  wire n_930_v;
  wire DA_AxB2_v;
  wire pipeVectorA2_v;
  wire n_745_v;
  wire n_1499_v;
  wire n_1495_v;
  wire n_1492_v;
  wire n_1323_v;
  wire n_1141_v;
  wire n_568_v;
  wire n_565_v;
  wire n_567_v;
  wire n_566_v;
  wire n_562_v;
  wire n_300_v;
  wire n_307_v;
  wire n_306_v;
  wire aluaorb0_v;
  wire x_op_T0_tya_v;
  wire x_op_T4_ind_y_v;
  wire pclp0_v;
  wire pclp1_v;
  wire pclp2_v;
  wire pclp3_v;
  wire pclp4_v;
  wire pclp5_v;
  wire pclp6_v;
  wire pclp7_v;
  wire op_T3_branch_v;
  wire n_79_v;
  wire n_75_v;
  wire n_70_v;
  wire n_71_v;
  wire n_1252_v;
  wire n_1705_v;
  wire n_1256_v;
  wire op_T0_tya_v;
  wire n_172_v;
  wire n_176_v;
  wire n_796_v;
  wire n_797_v;
  wire n_795_v;
  wire n_790_v;
  wire n_799_v;
  wire pd7_v;
  wire pd6_v;
  wire pd5_v;
  wire pd4_v;
  wire pd3_v;
  wire pd2_v;
  wire pd1_v;
  wire pd0_v;
  wire n_1305_v;
  wire n_1304_v;
  wire n_1303_v;
  wire n_1166_v;
  wire n_339_v;
  wire PD_1xx000x0_v;
  wire n_548_v;
  wire op_T2_brk_v;
  wire n_543_v;
  wire n_544_v;
  wire C56_v;
  wire n_890_v;
  wire n_323_v;
  wire n_897_v;
  wire n_896_v;
  wire n_329_v;
  wire pipeUNK31_v;
  wire xx_op_T5_jsr_v;
  wire PD_xxxx10x0_v;
  wire n_1028_v;
  wire n_50_v;
  wire n_55_v;
  wire n_152_v;
  wire n_154_v;
  wire n_1347_v;
  wire op_ORS_v;
  wire n_1346_v;
  wire _AxB_2__C12_v;
  wire n_1360_v;
  wire n_1364_v;
  wire n_1369_v;
  wire n_1368_v;
  wire clearIR_v;
  wire op_T__cpx_cpy_imm_zp_v;
  wire n_1187_v;
  wire n_1181_v;
  wire n_1180_v;
  wire op_T5_mem_ind_idx_v;
  wire n_521_v;
  wire n_523_v;
  wire n_525_v;
  wire n_526_v;
  wire C78_v;
  wire n_31_v;
  wire n_34_v;
  wire n_35_v;
  wire n_36_v;
  wire pchp4_v;
  wire pchp5_v;
  wire pchp6_v;
  wire pchp7_v;
  wire pchp0_v;
  wire pchp1_v;
  wire pchp2_v;
  wire pchp3_v;
  wire _WR_v;
  wire n_1642_v;
  wire n_1643_v;
  wire n_1640_v;
  wire n_1649_v;
  wire _op_branch_bit6_v;
  wire _op_branch_bit7_v;
  wire n_1184_v;
  wire op_rol_ror_v;
  wire n_201_v;
  wire clock2_v;
  wire n_1434_v;
  wire n_1341_v;
  wire op_asl_rol_v;
  wire short_circuit_idx_add_v;
  wire n_509_v;
  wire n_507_v;
  wire n_506_v;
  wire n_504_v;
  wire n_503_v;
  wire n_501_v;
  wire x_op_T0_bit_v;
  wire n_18_v;
  wire n_16_v;
  wire n_17_v;
  wire n_14_v;
  wire n_15_v;
  wire n_10_v;
  wire n_11_v;
  wire n_1085_v;
  wire n_1087_v;
  wire n_1081_v;
  wire n_1082_v;
  wire n_1089_v;
  wire n_1269_v;
  wire dpc35_PCHC_v;
  wire n_1265_v;
  wire n_1662_v;
  wire n_1262_v;
  wire op_T2_abs_y_v;
  wire n_267_v;
  wire n_264_v;
  wire n_265_v;
  wire n_262_v;
  wire n_260_v;
  wire n_261_v;
  wire n_269_v;
  wire n_8_v;
  wire op_T3_mem_abs_v;
  wire op_T2_ADL_ADD_v;
  wire n_1416_v;
  wire n_1413_v;
  wire n_1412_v;
  wire n_1411_v;
  wire n_383_v;
  wire n_385_v;
  wire n_384_v;
  wire n_386_v;
  wire n_389_v;
  wire n_388_v;
  wire op_T__shift_a_v;
  wire n_920_v;
  wire n_923_v;
  wire n_1039_v;
  wire op_T3_mem_zp_idx_v;
  wire notalucin_v;
  wire n_1069_v;
  wire n_1067_v;
  wire n_1065_v;
  wire n_1061_v;
  wire op_T0_tay_v;
  wire op_T0_tax_v;
  wire n_1606_v;
  wire op_T0_brk_rti_v;
  wire n_249_v;
  wire n_718_v;
  wire n_717_v;
  wire n_715_v;
  wire n_241_v;
  wire n_243_v;
  wire notidl0_v;
  wire op_T5_rti_rts_v;
  wire pipeT3out_v;
  wire n_669_v;
  wire _C23_v;
  wire nnT2BR_v;
  wire n_1472_v;
  wire n_1474_v;
  wire n_1477_v;
  wire op_T4_ind_y_v;
  wire n_1295_v;
  wire n_1291_v;
  wire n_1290_v;
  wire n_1293_v;
  wire op_T__iny_dey_v;
  wire n_902_v;
  wire n_906_v;
  wire n_905_v;
  wire n_1356_v;
  wire n_1423_v;
  wire pipeUNK18_v;
  wire pipeUNK16_v;
  wire pipeUNK17_v;
  wire pipeUNK14_v;
  wire pipeUNK15_v;
  wire pipeUNK12_v;
  wire pipeUNK13_v;
  wire pipeUNK11_v;
  wire n_38_v;
  wire n_1599_v;
  wire n_1043_v;
  wire n_1596_v;
  wire n_1045_v;
  wire n_1595_v;
  wire n_1624_v;
  wire n_1625_v;
  wire n_1629_v;
  wire n_228_v;
  wire n_223_v;
  wire n_220_v;
  wire n_221_v;
  wire n_226_v;
  wire n_224_v;
  wire n_225_v;
  wire op_T4_abs_idx_v;
  wire op_implied_v;
  wire n_735_v;
  wire n_730_v;
  wire n_732_v;
  wire dpc22__DSA_v;
  wire n_739_v;
  wire op_T__dex_v;
  wire n_415_v;
  wire _C01_v;
  wire op_T0_sbc_v;
  wire n_410_v;
  wire n_1452_v;
  wire n_1457_v;
  wire n_1455_v;
  wire DA_AB2_v;
  wire n_692_v;
  wire n_695_v;
  wire n_969_v;
  wire n_968_v;
  wire n_961_v;
  wire n_962_v;
  wire n_964_v;
  wire n_966_v;
  wire irline3_v;
  wire pipeUNK34_v;
  wire pipeUNK35_v;
  wire pipeUNK36_v;
  wire pipeUNK37_v;
  wire pipeUNK30_v;
  wire pipeUNK32_v;
  wire pipeUNK33_v;
  wire pipeUNK39_v;
  wire n_1020_v;
  wire n_1026_v;
  wire n_1027_v;
  wire n_1024_v;
  wire n_1025_v;
  wire n_1271_v;
  wire op_T2_branch_v;
  wire n_200_v;
  wire n_753_v;
  wire n_756_v;
  wire n_757_v;
  wire n_754_v;
  wire n_207_v;
  wire n_759_v;
  wire _C67_v;
  wire __AxB3__C23_v;
  wire pipephi2Reset0_v;
  wire pd5_clearIR_v;
  wire n_134_v;
  wire n_947_v;
  wire n_946_v;
  wire n_944_v;
  wire op_T0_cpy_iny_v;
  wire n_419_v;
  wire n_1007_v;
  wire n_1002_v;
  wire abh5_v;
  wire abh4_v;
  wire abh7_v;
  wire abh6_v;
  wire abh1_v;
  wire abh0_v;
  wire abh3_v;
  wire abh2_v;
  wire n_1552_v;
  wire alucin_v;
  wire x_op_push_pull_v;
  wire n_779_v;
  wire n_770_v;
  wire n_771_v;
  wire n_772_v;
  wire n_773_v;
  wire n_774_v;
  wire n_837_v;
  wire op_T0_bit_v;
  wire n_344_v;
  wire n_834_v;
  wire _C45_v;
  wire VEC0_v;
  wire VEC1_v;
  wire op_T4_rts_v;
  wire op_T4_rti_v;
  wire op_SRS_v;
  wire n_1343_v;
  wire n_1345_v;
  wire n_1578_v;
  wire n_1579_v;
  wire n_1573_v;
  wire n_1574_v;
  wire DC78_v;
  wire op_sta_cmp_v;
  wire op_SUMS_v;
  wire n_1688_v;
  wire pipeT2out_v;
  wire n_954_v;
  wire n_400_v;
  wire op_T4_brk_jsr_v;
  wire n_1219_v;
  wire n_1215_v;
  wire n_1214_v;
  wire n_1211_v;
  wire n_1213_v;
  wire n_1655_v;
  wire pd2_clearIR_v;
  wire n_1657_v;
  wire n_1650_v;
  wire n_182_v;
  wire n_180_v;
  wire n_184_v;
  wire n_637_v;
  wire n_636_v;
  wire n_631_v;
  wire n_630_v;
  wire n_632_v;
  wire n_459_v;
  wire n_988_v;
  wire n_983_v;
  wire n_982_v;
  wire n_981_v;
  wire n_987_v;
  wire n_986_v;
  wire n_457_v;
  wire op_T0_lda_v;
  wire abl1_v;
  wire abl0_v;
  wire abl4_v;
  wire pipe_WR_phi2_v;
  wire op_T3_plp_pla_v;
  wire n_1517_v;
  wire n_1518_v;
  wire DC78_phi2_v;
  wire n_279_v;
  wire n_846_v;
  wire n_847_v;
  wire n_844_v;
  wire n_845_v;
  wire n_842_v;
  wire op_T3_jmp_v;
  wire n_849_v;
  wire __AxB5__C45_v;
  wire n_1231_v;
  wire n_1230_v;
  wire n_1238_v;
  wire op_branch_done_v;
  wire aluvout_v;
  wire n_613_v;
  wire n_611_v;
  wire n_610_v;
  wire n_617_v;
  wire n_616_v;
  wire n_1137_v;
  wire n_620_v;
  wire n_1010_v;
  wire n_1017_v;
  wire n_1542_v;
  wire n_476_v;
  wire n_474_v;
  wire n_473_v;
  wire n_472_v;
  wire n_470_v;
  wire n_479_v;
  wire brk_done_v;
  wire p2_v;
  wire p3_v;
  wire op_T0_txa_v;
  wire p0_v;
  wire DC34_v;
  wire op_T2_stack_v;
  wire n_1534_v;
  wire n_1533_v;
  wire n_1391_v;
  wire n_1392_v;
  wire n_1395_v;
  wire n_1399_v;
  wire n_288_v;
  wire n_282_v;
  wire n_284_v;
  wire n_644_v;
  wire n_133_v;
  wire n_130_v;
  wire n_865_v;
  wire n_867_v;
  wire n_861_v;
  wire n_862_v;
  wire pipeT4out_v;
  wire pipeT_SYNC_v;
  wire _op_branch_done_v;
  wire op_T0_acc_v;
  wire BRtaken_v;
  wire n_1253_v;
  wire n_1257_v;
  wire n_1258_v;
  wire n_1708_v;
  wire op_T2_php_v;
  wire op_T2_pha_v;
  wire n_671_v;
  wire n_670_v;
  wire n_673_v;
  wire n_675_v;
  wire n_674_v;
  wire n_678_v;
  wire n_499_v;
  wire n_496_v;
  wire n_491_v;
  wire n_490_v;
  wire pd7_clearIR_v;
  wire n_1401_v;
  wire n_1404_v;
  wire op_T4_jmp_v;
  wire n_19_v;
  wire n_1117_v;
  wire n_1115_v;
  wire n_1113_v;
  wire n_1110_v;
  wire n_1111_v;
  wire n_803_v;
  wire n_800_v;
  wire n_805_v;
  wire n_432_v;
  wire n_1272_v;
  wire n_1277_v;
  wire n_1276_v;
  wire n_1275_v;
  wire n_1274_v;
  wire n_1660_v;
  wire op_inc_nop_v;
  wire n_128_v;
  wire n_127_v;
  wire n_126_v;
  wire n_653_v;
  wire n_122_v;
  wire op_T0_shift_right_a_v;
  wire op_T0_adc_sbc_v;
  wire op_push_pull_v;
  wire pipe_VEC_v;
  wire n_266_v;
  wire n_1130_v;
  wire n_1132_v;
  wire n_1133_v;
  wire n_1135_v;
  wire n_1138_v;
  wire op_T2_mem_zp_v;
  wire n_355_v;
  wire n_824_v;
  wire n_358_v;
  wire INTG_v;
  wire n_755_v;
  wire op_T2_ind_v;
  wire op_rti_rts_v;
  wire notdor1_v;
  wire notdor0_v;
  wire notdor3_v;
  wire notdor2_v;
  wire notdor5_v;
  wire notdor4_v;
  wire notdor7_v;
  wire notdor6_v;
  wire n_1570_v;
  wire n_109_v;
  wire n_108_v;
  wire n_101_v;
  wire n_105_v;
  wire n_104_v;
  wire n_1575_v;
  wire n_581_v;
  wire Reset0_v;
  wire n_1541_v;
  wire n_1484_v;
  wire x_op_jmp_v;
  wire n_1338_v;
  wire n_1339_v;
  wire n_1488_v;
  wire n_1335_v;
  wire n_1333_v;
  wire n_1159_v;
  wire n_1157_v;
  wire n_1154_v;
  wire _t2_v;
  wire _t3_v;
  wire n_595_v;
  wire n_597_v;
  wire _t4_v;
  wire _t5_v;
  wire nots3_v;
  wire nots2_v;
  wire nots1_v;
  wire nots0_v;
  wire nots7_v;
  wire nots6_v;
  wire nots5_v;
  wire nots4_v;
  wire n_1682_v;
  wire n_378_v;
  wire n_1683_v;
  wire n_374_v;
  wire n_372_v;
  wire x_op_T0_txa_v;
  wire C01_v;
  wire op_store_v;
  wire n_1687_v;
  wire n_80_v;
  wire n_83_v;
  wire n_88_v;
  wire n_1684_v;
  wire n_161_v;
  wire n_160_v;
  wire n_163_v;
  wire n_169_v;
  wire n_785_v;
  wire n_781_v;
  wire n_783_v;
  wire n_782_v;
  wire n_789_v;
  wire n_1319_v;
  wire n_1312_v;
  wire n_1315_v;
  wire n_1316_v;
  wire n_1175_v;
  wire n_1177_v;
  wire n_1170_v;
  wire n_1178_v;
  wire n_1179_v;
  wire n_572_v;
  wire n_570_v;
  wire n_318_v;
  wire n_319_v;
  wire n_312_v;
  wire n_311_v;
  wire n_317_v;
  wire PD_n_0xx0xx0x_v;
  wire C23_v;
  wire PD_0xx0xx0x_v;
  wire op_T0_dex_v;
  wire C78_phi2_v;
  wire op_T__ora_and_eor_adc_v;
  wire op_T2_ind_x_v;
  wire op_T2_ind_y_v;
  wire op_plp_pla_v;
  wire op_T0_txs_v;
  wire n_69_v;
  wire n_62_v;
  wire n_61_v;
  wire n_149_v;
  wire _op_set_C_v;
  wire op_T5_rti_v;
  wire op_T5_ind_y_v;
  wire op_T5_ind_x_v;
  wire op_T3_jsr_v;
  wire op_T5_brk_v;
  wire n_1371_v;
  wire n_1376_v;
  wire n_1377_v;
  wire n_1374_v;
  wire n_1375_v;
  wire n_1379_v;
  wire n_1194_v;
  wire n_1195_v;
  wire n_1192_v;
  wire n_1190_v;
  wire n_708_v;
  wire n_556_v;
  wire n_550_v;
  wire n_551_v;
  wire n_553_v;
  wire n_559_v;
  wire C45_v;
  wire x_op_T3_ind_y_v;
  wire op_T__asl_rol_a_v;
  wire n_882_v;
  wire n_334_v;
  wire n_335_v;
  wire n_885_v;
  wire n_888_v;
  wire n_889_v;
  wire _AxB_4__C34_v;
  wire dpc28_0ADH0_v;
  wire fetch_v;
  wire op_ANDS_v;
  wire n_47_v;
  wire n_46_v;
  wire op_T__cpx_cpy_abs_v;
  wire n_1153_v;
  wire n_0_ADL1_v;
  wire n_0_ADL0_v;
  wire n_0_ADL2_v;
  wire op_T3_abs_idx_v;
  wire op_jsr_v;
  wire n_590_v;
  wire n_593_v;
  wire n_598_v;
  wire n_1255_v;
  wire n_1358_v;
  wire n_1427_v;
  wire n_1357_v;
  wire n_533_v;
  wire n_531_v;
  wire n_538_v;
  wire C67_v;
  wire C1x5Reset_v;
  wire op_T__adc_sbc_v;
  wire op_T0_cmp_v;
  wire pipeBRtaken_v;
  wire n_1218_v;
  wire pipeUNK41_v;
  wire pipeUNK40_v;
  wire pipeUNK42_v;
  wire n_23_v;
  wire n_21_v;
  wire n_20_v;
  wire n_25_v;
  wire n_24_v;
  wire n_29_v;
  wire n_1693_v;
  wire pipephi2Reset0x_v;
  wire n_275_v;
  wire n_270_v;
  wire n_272_v;
  wire n_278_v;
  wire n_1486_v;
  wire n_638_v;
  wire n_1408_v;
  wire n_1409_v;
  wire n_188_v;
  wire n_1400_v;
  wire n_1402_v;
  wire op_T0_ora_v;
  wire n_519_v;
  wire n_510_v;
  wire n_512_v;
  wire n_513_v;
  wire n_515_v;
  wire n_1463_v;
  wire n_453_v;
  wire n_980_v;
  wire n_1464_v;
  wire alucout_v;
  wire op_brk_rti_v;
  wire DBZ_v;
  wire pipeVectorA0_v;
  wire pipeVectorA1_v;
  wire n_1602_v;
  wire pipeT5out_v;
  wire n_1600_v;
  wire n_1093_v;
  wire n_1091_v;
  wire n_1090_v;
  wire n_1097_v;
  wire n_1099_v;
  wire n_1679_v;
  wire n_1677_v;
  wire n_1676_v;
  wire n_1674_v;
  wire n_1673_v;
  wire op_T5_rts_v;
  wire n_253_v;
  wire n_251_v;
  wire n_709_v;
  wire n_256_v;
  wire n_255_v;
  wire n_700_v;
  wire n_1462_v;
  wire n_714_v;
  wire n_1286_v;
  wire n_1281_v;
  wire n_1289_v;
  wire A_B7_v;
  wire A_B5_v;
  wire A_B3_v;
  wire A_B1_v;
  wire n_392_v;
  wire n_393_v;
  wire n_390_v;
  wire n_396_v;
  wire n_397_v;
  wire n_398_v;
  wire n_1497_v;
  wire n_936_v;
  wire n_937_v;
  wire n_933_v;
  wire n_931_v;
  wire op_T2_php_pha_v;
  wire ONEBYTE_v;
  wire pipeUNK09_v;
  wire pipeUNK08_v;
  wire pipeUNK05_v;
  wire pipeUNK04_v;
  wire pipeUNK07_v;
  wire pipeUNK06_v;
  wire pipeUNK01_v;
  wire pipeUNK03_v;
  wire pipeUNK02_v;
  wire n_1075_v;
  wire n_1070_v;
  wire n_1073_v;
  wire n_1149_v;
  wire abl2_v;
  wire abl5_v;
  wire abl6_v;
  wire n_1619_v;
  wire notaluvout_v;
  wire n_1614_v;
  wire n_1145_v;
  wire dpc34_PCLC_v;
  wire H1x1_v;
  wire n_238_v;
  wire n_728_v;
  wire n_720_v;
  wire n_726_v;
  wire op_T2_abs_v;
  wire op_T0_plp_v;
  wire op_T0_pla_v;
  wire op_T2_jmp_abs_v;
  wire pipe_T0_v;
  wire _C34_v;
  wire DA_C01_v;
  wire n_1448_v;
  wire n_1449_v;
  wire n_1446_v;
  wire n_1447_v;
  wire n_1440_v;
  wire n_1441_v;
  wire notRnWprepad_v;
  wire n_1511_v;
  wire n_918_v;
  wire n_919_v;
  wire n_916_v;
  wire n_917_v;
  wire n_913_v;
  wire op_T0_tay_ldy_not_idx_v;
  wire op_T0_v;
  wire op_T3_v;
  wire op_T2_v;
  wire op_T4_v;
  wire n_1224_v;
  wire op_T3_stack_bit_jmp_v;
  wire op_T5_jsr_v;
  wire op_T2_stack_access_v;
  wire pipeUNK23_v;
  wire pipeUNK22_v;
  wire pipeUNK21_v;
  wire pipeUNK20_v;
  wire pipeUNK27_v;
  wire pipeUNK26_v;
  wire pipeUNK29_v;
  wire pipeUNK28_v;
  wire n_1056_v;
  wire n_1055_v;
  wire n_1054_v;
  wire op_T4_mem_abs_idx_v;
  wire n_1588_v;
  wire n_1581_v;
  wire n_1580_v;
  wire n_1638_v;
  wire C34_v;
  wire _DA_ADD2_v;
  wire _DA_ADD1_v;
  wire n_743_v;
  wire n_213_v;
  wire n_747_v;
  wire n_748_v;
  wire n_218_v;
  wire notalucout_v;
  wire dpc36_IPC_v;
  wire op_T0_cpx_cpy_inx_iny_v;
  wire op_T2_zp_zp_idx_v;
  wire _C12_v;
  wire n_688_v;
  wire n_689_v;
  wire n_680_v;
  wire n_1471_v;
  wire op_T4_ind_x_v;
  wire n_979_v;
  wire n_973_v;
  wire op_T__bit_v;
  wire op_T0_iny_dey_v;
  wire n_1270_v;
  wire op_T__cmp_v;
  wire op_T0_jsr_v;
  wire n_1610_v;
  wire op_T2_abs_access_v;
  wire n_1613_v;
  wire n_1033_v;
  wire n_1034_v;
  wire n_1037_v;
  wire n_1038_v;
  wire notalu4_v;
  wire notalu5_v;
  wire notalu6_v;
  wire notalu7_v;
  wire notalu0_v;
  wire notalu1_v;
  wire notalu2_v;
  wire notalu3_v;
  wire x_op_T4_rti_v;
  wire n_769_v;
  wire n_763_v;
  wire n_762_v;
  wire n_761_v;
  wire n_760_v;
  wire notidl4_v;
  wire notidl3_v;
  wire notidl1_v;
  wire op_T3_abs_idx_ind_v;
  wire op_T2_jsr_v;
  wire DA_C45_v;
  wire n_231_v;
  wire _C78_v;
  wire n_233_v;
  wire n_232_v;
  wire n_236_v;
  wire n_951_v;
  wire n_952_v;
  wire n_402_v;
  wire n_958_v;
  wire n_959_v;
  wire n_408_v;
  wire op_T0_eor_v;
  wire pd1_clearIR_v;
  wire abl3_v;
  wire op_T0_jmp_v;
  wire n_1018_v;
  wire n_1549_v;
  wire p1_v;
  wire __AxB1__C01_v;
  wire op_T2_idx_x_xy_v;
  wire _TWOCYCLE_phi1_v;
  wire op_clv_v;
  wire op_T0_and_v;
  wire op_T0_clc_sec_v;
  wire _C56_v;
  wire n_1209_v;
  wire n_1205_v;
  wire n_1202_v;
  wire n_1500_v;
  wire notidl5_v;
  wire n_428_v;
  wire n_424_v;
  wire n_420_v;
  wire op_sty_cpy_mem_v;
  wire n_1720_v;
  wire AxB5_v;
  wire AxB7_v;
  wire AxB1_v;
  wire AxB3_v;
  wire op_T3_ind_y_v;
  wire op_T3_ind_x_v;
  wire n_1566_v;
  wire n_1565_v;
  wire n_1561_v;
  wire n_1560_v;
  wire n_1697_v;
  wire n_1699_v;
  wire x_op_T3_abs_idx_v;
  wire op_from_x_v;
  wire n_850_v;
  wire n_853_v;
  wire n_852_v;
  wire op_T0_cli_sei_v;
  wire op_T0_ldx_tax_tsx_v;
  wire n_1049_v;
  wire n_1229_v;
  wire n_1593_v;
  wire n_1221_v;
  wire n_1222_v;
  wire n_1223_v;
  wire n_1225_v;
  wire n_1044_v;
  wire n_1594_v;
  wire n_1047_v;
  wire n_198_v;
  wire n_628_v;
  wire n_629_v;
  wire n_626_v;
  wire n_196_v;
  wire n_625_v;
  wire n_190_v;
  wire n_191_v;
  wire n_192_v;
  wire n_621_v;
  wire n_442_v;
  wire n_440_v;
  wire n_441_v;
  wire n_445_v;
  wire DBNeg_v;
  wire op_T0_tsx_v;
  wire notidl7_v;
  wire notidl6_v;
  wire notidl2_v;
  wire n_995_v;
  wire n_990_v;
  wire n_992_v;
  wire n_993_v;
  wire _op_store_v;
  wire n_1505_v;
  wire n_1509_v;
  wire op_T0_cpx_inx_v;
  wire n_299_v;
  wire n_293_v;
  wire n_291_v;
  wire n_877_v;
  wire n_876_v;
  wire n_875_v;
  wire n_878_v;
  wire n_956_v;

  spice_pin_input pin_4286(nmi, nmi_v, nmi_port_2);
  spice_pin_input pin_4287(irq, irq_v, irq_port_2);
  spice_pin_input pin_4285(rdy, rdy_v, rdy_port_3);
  spice_pin_input pin_4282(clk0, clk0_v, clk0_port_3);
  spice_pin_input pin_4281(so, so_v, so_port_3);
  spice_pin_input pin_4278(res, res_v, res_port_2);

  spice_pin_output pin_4284(clk2out, clk2out_v);
  spice_pin_output pin_4283(clk1out, clk1out_v);
  spice_pin_output pin_4280(sync, sync_v);
  spice_pin_output pin_4268(ab14, ab14_v);
  spice_pin_output pin_4264(ab10, ab10_v);
  spice_pin_output pin_4266(ab12, ab12_v);
  spice_pin_output pin_4260(ab6, ab6_v);
  spice_pin_output pin_4261(ab7, ab7_v);
  spice_pin_output pin_4262(ab8, ab8_v);
  spice_pin_output pin_4263(ab9, ab9_v);
  spice_pin_output pin_4269(ab15, ab15_v);
  spice_pin_output pin_4265(ab11, ab11_v);
  spice_pin_output pin_4267(ab13, ab13_v);
  spice_pin_output pin_4279(rw, rw_v);
  spice_pin_output pin_4255(ab1, ab1_v);
  spice_pin_output pin_4254(ab0, ab0_v);
  spice_pin_output pin_4257(ab3, ab3_v);
  spice_pin_output pin_4256(ab2, ab2_v);
  spice_pin_output pin_4259(ab5, ab5_v);
  spice_pin_output pin_4258(ab4, ab4_v);

  spice_pin_bidirectional pin_4277(db7_i, db7_o, db7_t, db7_v, db7_port_5);
  spice_pin_bidirectional pin_4276(db6_i, db6_o, db6_t, db6_v, db6_port_5);
  spice_pin_bidirectional pin_4275(db5_i, db5_o, db5_t, db5_v, db5_port_5);
  spice_pin_bidirectional pin_4274(db4_i, db4_o, db4_t, db4_v, db4_port_5);
  spice_pin_bidirectional pin_4273(db3_i, db3_o, db3_t, db3_v, db3_port_5);
  spice_pin_bidirectional pin_4272(db2_i, db2_o, db2_t, db2_v, db2_port_5);
  spice_pin_bidirectional pin_4271(db1_i, db1_o, db1_t, db1_v, db1_port_5);
  spice_pin_bidirectional pin_4270(db0_i, db0_o, db0_t, db0_v, db0_port_5);

  spice_transistor_nmos_gnd g_4387((dor3_v|~RnWstretched_v[`W-1]), n_643_v, n_643_port_4);
  spice_transistor_nmos t3178(~dpc39_PCLPCL_v[`W-1], pcl0_v, n_488_v, pcl0_port_1, n_488_port_3);
  spice_transistor_nmos t3179(~dpc39_PCLPCL_v[`W-1], pcl3_v, n_723_v, pcl3_port_1, n_723_port_3);
  spice_transistor_nmos t3174(~dpc39_PCLPCL_v[`W-1], pcl4_v, n_208_v, pcl4_port_1, n_208_port_3);
  spice_transistor_nmos t3175(~dpc39_PCLPCL_v[`W-1], pcl7_v, n_1647_v, pcl7_port_2, n_1647_port_3);
  spice_transistor_nmos t3176(~dpc39_PCLPCL_v[`W-1], pcl6_v, n_1458_v, pcl6_port_1, n_1458_port_3);
  spice_transistor_nmos t3177(~dpc39_PCLPCL_v[`W-1], pcl1_v, n_976_v, pcl1_port_1, n_976_port_2);
  spice_transistor_nmos t3173(~dpc39_PCLPCL_v[`W-1], pcl5_v, n_72_v, pcl5_port_1, n_72_port_3);
  spice_transistor_nmos t989(~dpc37_PCLDB_v[`W-1], idb0_v, n_488_v, idb0_port_6, n_488_port_1);
  spice_transistor_nmos_gnd t1539(n_1552_v, dpc14_SRS_v, dpc14_SRS_port_2);
  spice_transistor_nmos_gnd g_4605((~cclk_v[`W-1]|n_602_v|~n_1247_v[`W-1]), dpc2_XSB_v, dpc2_XSB_port_12);
  spice_transistor_nmos_gnd g_4600((n_1613_v|~RnWstretched_v[`W-1]), n_42_v, n_42_port_4);
  spice_transistor_nmos_gnd g_4601((~alua0_v[`W-1]|~alub0_v[`W-1]), aluanorb0_v, aluanorb0_port_7);
  spice_transistor_nmos_gnd t3365(~adl5_v[`W-1], n_1094_v, n_1094_port_1);
  spice_transistor_nmos_vdd t167(dor5_v, n_373_v, n_373_port_0);
  spice_transistor_nmos_vdd t166(~n_1296_v[`W-1], ab11_v, ab11_port_0);
  spice_transistor_nmos t1571(~cclk_v[`W-1], n_658_v, y4_v, n_658_port_0, y4_port_2);
  spice_transistor_nmos t2363(~dpc24_ACSB_v[`W-1], sb0_v, n_146_v, sb0_port_10, n_146_port_2);
  spice_transistor_nmos t2366(~dpc24_ACSB_v[`W-1], sb3_v, n_1654_v, sb3_port_10, n_1654_port_3);
  spice_transistor_nmos t2367(~dpc24_ACSB_v[`W-1], sb4_v, n_1344_v, sb4_port_11, n_1344_port_1);
  spice_transistor_nmos t2364(~dpc24_ACSB_v[`W-1], sb1_v, n_929_v, sb1_port_9, n_929_port_3);
  spice_transistor_nmos t2365(~dpc24_ACSB_v[`W-1], n_1618_v, sb2_v, n_1618_port_1, sb2_port_9);
  spice_transistor_nmos t2368(~dpc24_ACSB_v[`W-1], sb5_v, n_831_v, sb5_port_8, n_831_port_2);
  spice_transistor_nmos t2369(~dpc24_ACSB_v[`W-1], n_326_v, sb6_v, n_326_port_3, sb6_port_11);
  spice_transistor_nmos_vdd t570(n_772_v, dpc17_SUMS_v, dpc17_SUMS_port_1);
  spice_transistor_nmos_gnd t572(pclp2_v, n_481_v, n_481_port_0);
  spice_transistor_nmos_vdd t578(dor2_v, n_520_v, n_520_port_0);
  spice_transistor_nmos_gnd t2189(n_890_v, n_1694_v, n_1694_port_1);
  spice_transistor_nmos_gnd t1983(n_1033_v, dpc21_ADDADL_v, dpc21_ADDADL_port_9);
  spice_transistor_nmos t1183(~cclk_v[`W-1], x1_v, n_1709_v, x1_port_0, n_1709_port_0);
  spice_transistor_nmos_gnd t1180(abl1_v, n_66_v, n_66_port_1);
  spice_transistor_nmos_gnd t1184(n_0_ADL1_v, adl1_v, adl1_port_1);
  spice_transistor_nmos t2197(~dpc27_SBADH_v[`W-1], adh4_v, sb4_v, adh4_port_4, sb4_port_9);
  spice_transistor_nmos t372(~dpc10_ADLADD_v[`W-1], adl0_v, alub0_v, adl0_port_1, alub0_port_2);
  spice_transistor_nmos t374(~dpc4_SSB_v[`W-1], n_694_v, sb1_v, n_694_port_1, sb1_port_2);
  spice_transistor_nmos_gnd t375(~n_869_v[`W-1], ab13_v, ab13_port_1);
  spice_transistor_nmos_vdd t2523(n_747_v, clk1out_v, clk1out_port_1);
  spice_transistor_nmos t2526(~dpc38_PCLADL_v[`W-1], n_72_v, adl5_v, n_72_port_2, adl5_port_4);
  spice_transistor_nmos t2527(~dpc38_PCLADL_v[`W-1], adl6_v, n_1458_v, adl6_port_4, n_1458_port_1);
  spice_transistor_nmos_gnd g_4832((~alua5_v[`W-1]&~alub5_v[`W-1]), n_477_v, n_477_port_5);
  spice_transistor_nmos g_4839((~cp1_v[`W-1]&fetch_v), n_1641_v, n_119_v, n_1641_port_3, n_119_port_3);
  spice_transistor_nmos t3118(~dpc2_XSB_v[`W-1], n_1694_v, sb2_v, n_1694_port_2, sb2_port_10);
  spice_transistor_nmos t3119(~dpc2_XSB_v[`W-1], n_242_v, sb3_v, n_242_port_2, sb3_port_11);
  spice_transistor_nmos t3116(~dpc2_XSB_v[`W-1], n_1724_v, sb6_v, n_1724_port_2, sb6_port_12);
  spice_transistor_nmos_gnd t3117(n_1256_v, dpc15_ANDS_v, dpc15_ANDS_port_9);
  spice_transistor_nmos t3115(~dpc2_XSB_v[`W-1], n_578_v, sb5_v, n_578_port_1, sb5_port_10);
  spice_transistor_nmos_gnd t2645(notidl3_v, idl3_v, idl3_port_0);
  spice_transistor_nmos_gnd t2640(notalu5_v, alu5_v, alu5_port_3);
  spice_transistor_nmos t963(~dpc6_SBS_v[`W-1], sb0_v, s0_v, sb0_port_3, s0_port_1);
  spice_transistor_nmos t962(~cclk_v[`W-1], n_1694_v, x2_v, n_1694_port_0, x2_port_0);
  spice_transistor_nmos_vdd t961(~cclk_v[`W-1], idb3_v, idb3_port_1);
  spice_transistor_nmos_gnd t1046(pchp2_v, n_1496_v, n_1496_port_0);
  spice_transistor_nmos t1047(~cclk_v[`W-1], n_1251_v, y7_v, n_1251_port_0, y7_port_0);
  spice_transistor_nmos_gnd t1040(~adh1_v[`W-1], n_1267_v, n_1267_port_0);
  spice_transistor_nmos_gnd t1519(pchp6_v, n_652_v, n_652_port_0);
  spice_transistor_nmos_gnd t1048(~adl4_v[`W-1], n_1519_v, n_1519_port_0);
  spice_transistor_nmos_gnd g_4620((~n_1247_v[`W-1]|n_956_v|~cclk_v[`W-1]), dpc12_0ADD_v, dpc12_0ADD_port_12);
  spice_transistor_nmos_gnd g_4626((~RnWstretched_v[`W-1]|n_1463_v), n_1076_v, n_1076_port_4);
  spice_transistor_nmos_gnd g_4627((~n_1247_v[`W-1]|n_228_v|~cclk_v[`W-1]), dpc30_ADHPCH_v, dpc30_ADHPCH_port_12);
  spice_transistor_nmos_gnd t3438(n_906_v, dpc19_ADDSB7_v, dpc19_ADDSB7_port_2);
  spice_transistor_nmos t1533(~dpc3_SBX_v[`W-1], x7_v, sb7_v, x7_port_1, sb7_port_2);
  spice_transistor_nmos t3347(~dpc11_SBADD_v[`W-1], sb7_v, alua7_v, sb7_port_10, alua7_port_3);
  spice_transistor_nmos t3342(~cp1_v[`W-1], n_1095_v, idl4_v, n_1095_port_3, idl4_port_1);
  spice_transistor_nmos_vdd t3340(~cclk_v[`W-1], sb5_v, sb5_port_12);
  spice_transistor_nmos_vdd t1536(~n_520_v[`W-1], db2_v, db2_port_3);
  spice_transistor_nmos_vdd t149(n_154_v, dpc20_ADDSB06_v, dpc20_ADDSB06_port_0);
  spice_transistor_nmos_gnd t147(~idb0_v[`W-1], n_624_v, n_624_port_0);
  spice_transistor_nmos_gnd t146(AxB3_v, n_884_v, n_884_port_0);
  spice_transistor_nmos t142(~cp1_v[`W-1], n_1424_v, idl2_v, n_1424_port_0, idl2_port_1);
  spice_transistor_nmos_gnd t2252(abh2_v, n_994_v, n_994_port_1);
  spice_transistor_nmos_vdd t2250(abh2_v, n_1545_v, n_1545_port_1);
  spice_transistor_nmos_gnd t551(~n_1417_v[`W-1], clk1out_v, clk1out_port_0);
  spice_transistor_nmos t2254(~dpc27_SBADH_v[`W-1], sb1_v, adh1_v, sb1_port_8, adh1_port_4);
  spice_transistor_nmos_gnd t2255(~dpc12_0ADD_v[`W-1], alua2_v, alua2_port_1);
  spice_transistor_nmos_gnd t312(n_445_v, sync_v, sync_port_0);
  spice_transistor_nmos g_4819((~cp1_v[`W-1]&~ADH_ABH_v[`W-1]), n_1668_v, _ABH0_v, n_1668_port_3, _ABH0_port_3);
  spice_transistor_nmos_vdd t3132(n_531_v, dpc13_ORS_v, dpc13_ORS_port_8);
  spice_transistor_nmos_vdd t3133(dor7_v, n_298_v, n_298_port_3);
  spice_transistor_nmos t3134(~cclk_v[`W-1], _ABH4_v, n_999_v, _ABH4_port_2, n_999_port_3);
  spice_transistor_nmos_gnd t3137(notidl5_v, idl5_v, idl5_port_1);
  spice_transistor_nmos_gnd t1280(pd5_clearIR_v, n_928_v, n_928_port_1);
  spice_transistor_nmos t941(~dpc16_EORS_v[`W-1], n_1469_v, n_277_v, n_1469_port_0, n_277_port_1);
  spice_transistor_nmos t940(~dpc16_EORS_v[`W-1], __AxB_4_v, n_296_v, __AxB_4_port_0, n_296_port_0);
  spice_transistor_nmos t943(~dpc16_EORS_v[`W-1], n_304_v, n_177_v, n_304_port_1, n_177_port_1);
  spice_transistor_nmos t942(~dpc16_EORS_v[`W-1], __AxB_6_v, n_722_v, __AxB_6_port_2, n_722_port_1);
  spice_transistor_nmos_gnd t2889(ir4_v, notir4_v, notir4_port_25);
  spice_transistor_nmos t2883(n_771_v, n_430_v, n_465_v, n_430_port_3, n_465_port_1);
  spice_transistor_nmos_gnd g_4640((~cclk_v[`W-1]|~n_1247_v[`W-1]|n_708_v), dpc11_SBADD_v, dpc11_SBADD_port_12);
  spice_transistor_nmos_gnd g_4641((~cclk_v[`W-1]|n_441_v|~n_1247_v[`W-1]), dpc1_SBY_v, dpc1_SBY_port_12);
  spice_transistor_nmos t1476(~cclk_v[`W-1], n_676_v, _ABH1_v, n_676_port_0, _ABH1_port_0);
  spice_transistor_nmos_vdd t1471(n_91_v, dpc15_ANDS_v, dpc15_ANDS_port_0);
  spice_transistor_nmos_gnd t1126(n_1025_v, n_564_v, n_564_port_1);
  spice_transistor_nmos t128(~dpc4_SSB_v[`W-1], n_1389_v, sb2_v, n_1389_port_0, sb2_port_1);
  spice_transistor_nmos_gnd t121(pclp7_v, n_1647_v, n_1647_port_0);
  spice_transistor_nmos t127(~dpc4_SSB_v[`W-1], n_998_v, sb3_v, n_998_port_0, sb3_port_1);
  spice_transistor_nmos_gnd t1496(~n_1105_v[`W-1], cp1_v, cp1_port_50);
  spice_transistor_nmos t1723(~dpc5_SADL_v[`W-1], adl3_v, n_998_v, adl3_port_3, n_998_port_3);
  spice_transistor_nmos t1722(~dpc5_SADL_v[`W-1], adl4_v, n_3_v, adl4_port_4, n_3_port_3);
  spice_transistor_nmos t1721(~dpc5_SADL_v[`W-1], adl5_v, n_280_v, adl5_port_3, n_280_port_3);
  spice_transistor_nmos t1727(~dpc5_SADL_v[`W-1], n_721_v, adl7_v, n_721_port_3, adl7_port_2);
  spice_transistor_nmos t1724(~dpc5_SADL_v[`W-1], adl2_v, n_1389_v, adl2_port_3, n_1389_port_2);
  spice_transistor_nmos_gnd t338(pclp0_v, n_488_v, n_488_port_0);
  spice_transistor_nmos_vdd t333(dor1_v, n_798_v, n_798_port_1);
  spice_transistor_nmos_gnd g_4789((aluaorb0_v&~aluanandb0_v[`W-1]), __AxB_0_v, __AxB_0_port_6);
  spice_transistor_nmos g_4785((~cp1_v[`W-1]&~ADL_ABL_v[`W-1]), n_1016_v, _ABL1_v, n_1016_port_3, _ABL1_port_3);
  spice_transistor_nmos g_4783((~ADL_ABL_v[`W-1]&~cp1_v[`W-1]), _ABL3_v, n_1507_v, _ABL3_port_3, n_1507_port_3);
  spice_transistor_nmos_gnd g_4878(((n_36_v&n_320_v)|n_735_v), dasb1_v, dasb1_port_5);
  spice_transistor_nmos_vdd t2066(n_1028_v, RnWstretched_v, RnWstretched_port_23);
  spice_transistor_nmos t1228(~cclk_v[`W-1], n_1592_v, a7_v, n_1592_port_0, a7_port_1);
  spice_transistor_nmos_gnd t692(n_567_v, n_171_v, n_171_port_0);
  spice_transistor_nmos_vdd t694(n_567_v, n_322_v, n_322_port_1);
  spice_transistor_nmos t696(~cclk_v[`W-1], n_1620_v, notir3_v, n_1620_port_0, notir3_port_1);
  spice_transistor_nmos_gnd t2605(n_1660_v, n_855_v, n_855_port_2);
  spice_transistor_nmos_vdd t2606(n_1660_v, n_1100_v, n_1100_port_3);
  spice_transistor_nmos_gnd t1009(ir2_v, notir2_v, notir2_port_0);
  spice_transistor_nmos_gnd g_4669((dor6_v|~RnWstretched_v[`W-1]), n_471_v, n_471_port_4);
  spice_transistor_nmos_gnd g_4664((n_1720_v|~RnWstretched_v[`W-1]), n_373_v, n_373_port_4);
  spice_transistor_nmos_gnd g_4665((~n_1247_v[`W-1]|n_255_v|~cclk_v[`W-1]), dpc31_PCHPCH_v, dpc31_PCHPCH_port_12);
  spice_transistor_nmos_vdd t104(~n_963_v[`W-1], ab14_v, ab14_port_0);
  spice_transistor_nmos_vdd t109(abh3_v, n_1296_v, n_1296_port_0);
  spice_transistor_nmos t2476(~dpc31_PCHPCH_v[`W-1], pch7_v, n_1206_v, pch7_port_2, n_1206_port_1);
  spice_transistor_nmos t2477(~dpc31_PCHPCH_v[`W-1], pch4_v, n_27_v, pch4_port_2, n_27_port_1);
  spice_transistor_nmos t2475(~dpc31_PCHPCH_v[`W-1], pch6_v, n_652_v, pch6_port_2, n_652_port_1);
  spice_transistor_nmos t2478(~dpc31_PCHPCH_v[`W-1], pch5_v, n_1301_v, pch5_port_2, n_1301_port_1);
  spice_transistor_nmos t2479(~dpc31_PCHPCH_v[`W-1], pch2_v, n_1496_v, pch2_port_1, n_1496_port_1);
  spice_transistor_nmos_vdd t1(~n_1608_v[`W-1], ab13_v, ab13_port_0);
  spice_transistor_nmos_vdd t1922(~n_1152_v[`W-1], ab2_v, ab2_port_0);
  spice_transistor_nmos_vdd t481(n_670_v, n_1417_v, n_1417_port_0);
  spice_transistor_nmos_gnd t482(~n_994_v[`W-1], ab10_v, ab10_port_1);
  spice_transistor_nmos_gnd t489(n_1439_v, n_518_v, n_518_port_1);
  spice_transistor_nmos_vdd t1749(n_1596_v, dpc27_SBADH_v, dpc27_SBADH_port_0);
  spice_transistor_nmos_vdd t1746(n_966_v, dpc29_0ADH17_v, dpc29_0ADH17_port_2);
  spice_transistor_nmos g_4857((~ADH_ABH_v[`W-1]&~cp1_v[`W-1]), _ABH6_v, n_880_v, _ABH6_port_3, n_880_port_3);
  spice_transistor_nmos g_4858((~ADH_ABH_v[`W-1]&~cp1_v[`W-1]), _ABH3_v, n_883_v, _ABH3_port_3, n_883_port_3);
  spice_transistor_nmos t83(H1x1_v, idb2_v, Pout2_v, idb2_port_0, Pout2_port_0);
  spice_transistor_nmos t2257(~dpc0_YSB_v[`W-1], n_1251_v, sb7_v, n_1251_port_1, sb7_port_8);
  spice_transistor_nmos t2745(~dpc37_PCLDB_v[`W-1], n_723_v, idb3_v, n_723_port_2, idb3_port_9);
  spice_transistor_nmos t2746(~dpc37_PCLDB_v[`W-1], n_976_v, idb1_v, n_976_port_1, idb1_port_8);
  spice_transistor_nmos_vdd t2598(~cclk_v[`W-1], idb6_v, idb6_port_9);
  spice_transistor_nmos t2592(~dpc13_ORS_v[`W-1], n_404_v, n_296_v, n_404_port_2, n_296_port_5);
  spice_transistor_nmos_vdd t2622(n_1153_v, n_659_v, n_659_port_2);
  spice_transistor_nmos_gnd t2621(n_1153_v, n_1639_v, n_1639_port_2);
  spice_transistor_nmos_gnd t905(~n_635_v[`W-1], ab14_v, ab14_port_1);
  spice_transistor_nmos t1985(~dpc1_SBY_v[`W-1], y3_v, sb3_v, y3_port_2, sb3_port_8);
  spice_transistor_nmos t1984(~dpc40_ADLPCL_v[`W-1], pcl7_v, adl7_v, pcl7_port_1, adl7_port_4);
  spice_transistor_nmos_gnd t1327(n_1484_v, n_1491_v, n_1491_port_1);
  spice_transistor_nmos_gnd t1024(~n_471_v[`W-1], db6_v, db6_port_0);
  spice_transistor_nmos t1505(~dpc0_YSB_v[`W-1], n_1491_v, sb2_v, n_1491_port_2, sb2_port_3);
  spice_transistor_nmos_gnd t2459(abh7_v, n_659_v, n_659_port_1);
  spice_transistor_nmos t2450(~dpc30_ADHPCH_v[`W-1], pch1_v, adh1_v, pch1_port_1, adh1_port_5);
  spice_transistor_nmos t2453(~dpc30_ADHPCH_v[`W-1], pch0_v, adh0_v, pch0_port_1, adh0_port_4);
  spice_transistor_nmos_gnd t2455(abh1_v, n_676_v, n_676_port_2);
  spice_transistor_nmos_vdd t2457(abh7_v, n_1639_v, n_1639_port_0);
  spice_transistor_nmos_vdd t1182(abl1_v, n_1479_v, n_1479_port_0);
  spice_transistor_nmos_gnd t3057(~n_1467_v[`W-1], cclk_v, cclk_port_236);
  spice_transistor_nmos_vdd t3055(n_1364_v, dpc16_EORS_v, dpc16_EORS_port_9);
  spice_transistor_nmos_vdd t3504(~cclk_v[`W-1], idb4_v, idb4_port_10);
  spice_transistor_nmos_vdd t3501(n_951_v, n_642_v, n_642_port_3);
  spice_transistor_nmos_gnd t3500(n_951_v, n_1152_v, n_1152_port_2);
  spice_transistor_nmos_vdd t3502(~cclk_v[`W-1], sb2_v, sb2_port_12);
  spice_transistor_nmos_vdd t2902(n_830_v, dpc23_SBAC_v, dpc23_SBAC_port_11);
  spice_transistor_nmos_vdd t1760(~cclk_v[`W-1], idb2_v, idb2_port_4);
  spice_transistor_nmos_gnd g_4302((~n_1247_v[`W-1]|n_1047_v|~cclk_v[`W-1]), dpc23_SBAC_v, dpc23_SBAC_port_12);
  spice_transistor_nmos_gnd t3196(~idb7_v[`W-1], n_423_v, n_423_port_1);
  spice_transistor_nmos t3195(~dpc4_SSB_v[`W-1], n_332_v, sb0_v, n_332_port_3, sb0_port_12);
  spice_transistor_nmos_vdd t2028(~cclk_v[`W-1], adh7_v, adh7_port_2);
  spice_transistor_nmos t521(~dpc21_ADDADL_v[`W-1], adl3_v, alu3_v, adl3_port_0, alu3_port_0);
  spice_transistor_nmos t520(~cp1_v[`W-1], n_87_v, idl1_v, n_87_port_1, idl1_port_0);
  spice_transistor_nmos t1599(~dpc1_SBY_v[`W-1], y2_v, sb2_v, y2_port_2, sb2_port_6);
  spice_transistor_nmos t1590(~dpc14_SRS_v[`W-1], aluanandb1_v, notaluoutmux0_v, aluanandb1_port_0, notaluoutmux0_port_2);
  spice_transistor_nmos t1591(~dpc14_SRS_v[`W-1], notaluoutmux1_v, n_681_v, notaluoutmux1_port_2, n_681_port_1);
  spice_transistor_nmos t1592(~dpc14_SRS_v[`W-1], n_350_v, n_740_v, n_350_port_1, n_740_port_3);
  spice_transistor_nmos t1593(~dpc14_SRS_v[`W-1], n_1071_v, n_1063_v, n_1071_port_4, n_1063_port_2);
  spice_transistor_nmos t1594(~dpc14_SRS_v[`W-1], n_296_v, n_477_v, n_296_port_3, n_477_port_1);
  spice_transistor_nmos t1595(~dpc14_SRS_v[`W-1], n_277_v, n_336_v, n_277_port_3, n_336_port_1);
  spice_transistor_nmos t1596(~dpc14_SRS_v[`W-1], n_722_v, n_1318_v, n_722_port_4, n_1318_port_2);
  spice_transistor_nmos_gnd t1980(~adh4_v[`W-1], n_212_v, n_212_port_1);
  spice_transistor_nmos t588(~dpc43_DL_DB_v[`W-1], idb3_v, n_1661_v, idb3_port_0, n_1661_port_1);
  spice_transistor_nmos t585(~dpc43_DL_DB_v[`W-1], idb0_v, n_719_v, idb0_port_5, n_719_port_2);
  spice_transistor_nmos_gnd t1640(n_1521_v, n_242_v, n_242_port_1);
  spice_transistor_nmos t1641(~dpc1_SBY_v[`W-1], y1_v, sb1_v, y1_port_2, sb1_port_5);
  spice_transistor_nmos_gnd t3038(~n_147_v[`W-1], db4_v, db4_port_3);
  spice_transistor_nmos_gnd t3030(n_90_v, p6_v, p6_port_1);
  spice_transistor_nmos_vdd t3035(n_769_v, n_1072_v, n_1072_port_2);
  spice_transistor_nmos t1961(~dpc5_SADL_v[`W-1], adl0_v, n_332_v, adl0_port_4, n_332_port_1);
  spice_transistor_nmos t1964(~cclk_v[`W-1], n_1300_v, notir2_v, n_1300_port_2, notir2_port_19);
  spice_transistor_nmos_gnd t1969(pclp3_v, n_723_v, n_723_port_0);
  spice_transistor_nmos t3373(~dpc40_ADLPCL_v[`W-1], pcl1_v, adl1_v, pcl1_port_2, adl1_port_8);
  spice_transistor_nmos t3375(~dpc40_ADLPCL_v[`W-1], pcl3_v, adl3_v, pcl3_port_2, adl3_port_7);
  spice_transistor_nmos t1782(~dpc1_SBY_v[`W-1], y7_v, sb7_v, y7_port_1, sb7_port_4);
  spice_transistor_nmos g_4728((~cp1_v[`W-1]&fetch_v), n_1605_v, n_541_v, n_1605_port_5, n_541_port_3);
  spice_transistor_nmos g_4726((~ADH_ABH_v[`W-1]&~cp1_v[`W-1]), _ABH7_v, n_494_v, _ABH7_port_3, n_494_port_3);
  spice_transistor_nmos g_4723((~ADH_ABH_v[`W-1]&~cp1_v[`W-1]), _ABH2_v, n_168_v, _ABH2_port_3, n_168_port_3);
  spice_transistor_nmos_gnd g_4891(((_C67_v&AxB7_v)|__AxB7__C67_v), __AxBxC_7_v, __AxBxC_7_port_5);
  spice_transistor_nmos_gnd g_4890((_AxB_0__C0in_v|(n_105_v&~__AxB_0_v[`W-1])), __AxBxC_0_v, __AxBxC_0_port_5);
  spice_transistor_nmos_gnd g_4899(((AxB1_v&_C01_v)|__AxB1__C01_v), __AxBxC_1_v, __AxBxC_1_port_5);
  spice_transistor_nmos t49(~dpc11_SBADD_v[`W-1], alua4_v, sb4_v, alua4_port_0, sb4_port_1);
  spice_transistor_nmos t48(~dpc11_SBADD_v[`W-1], alua3_v, sb3_v, alua3_port_0, sb3_port_0);
  spice_transistor_nmos_gnd t42(pd0_clearIR_v, n_409_v, n_409_port_0);
  spice_transistor_nmos t47(~dpc11_SBADD_v[`W-1], sb2_v, alua2_v, sb2_port_0, alua2_port_0);
  spice_transistor_nmos t46(~dpc11_SBADD_v[`W-1], sb1_v, alua1_v, sb1_port_0, alua1_port_2);
  spice_transistor_nmos t45(~cclk_v[`W-1], y1_v, n_767_v, y1_port_0, n_767_port_0);
  spice_transistor_nmos_gnd t44(notalu4_v, alu4_v, alu4_port_0);
  spice_transistor_nmos t3203(~dpc10_ADLADD_v[`W-1], adl6_v, alub6_v, adl6_port_6, alub6_port_4);
  spice_transistor_nmos t3206(~dpc10_ADLADD_v[`W-1], adl1_v, alub1_v, adl1_port_7, alub1_port_4);
  spice_transistor_nmos t3207(~dpc10_ADLADD_v[`W-1], adl4_v, alub4_v, adl4_port_6, alub4_port_4);
  spice_transistor_nmos t3204(~dpc10_ADLADD_v[`W-1], adl7_v, alub7_v, adl7_port_6, alub7_port_4);
  spice_transistor_nmos t3208(~dpc10_ADLADD_v[`W-1], alub5_v, adl5_v, alub5_port_4, adl5_port_5);
  spice_transistor_nmos t283(~dpc7_SS_v[`W-1], n_618_v, s6_v, n_618_port_1, s6_port_1);
  spice_transistor_nmos t286(~dpc7_SS_v[`W-1], n_998_v, s3_v, n_998_port_1, s3_port_1);
  spice_transistor_nmos t287(~dpc7_SS_v[`W-1], n_1389_v, s2_v, n_1389_port_1, s2_port_1);
  spice_transistor_nmos t284(~dpc7_SS_v[`W-1], n_280_v, s5_v, n_280_port_0, s5_port_1);
  spice_transistor_nmos t285(~dpc7_SS_v[`W-1], n_3_v, s4_v, n_3_port_1, s4_port_1);
  spice_transistor_nmos t288(~dpc7_SS_v[`W-1], n_694_v, s1_v, n_694_port_0, s1_port_1);
  spice_transistor_nmos_gnd t289(~adh3_v[`W-1], n_883_v, n_883_port_1);
  spice_transistor_nmos t2009(~cclk_v[`W-1], n_541_v, notir7_v, n_541_port_1, notir7_port_34);
  spice_transistor_nmos_gnd t2008(n_1067_v, ADH_ABH_v, ADH_ABH_port_7);
  spice_transistor_nmos t2551(~dpc32_PCHADH_v[`W-1], adh3_v, n_141_v, adh3_port_6, n_141_port_2);
  spice_transistor_nmos t2550(~dpc32_PCHADH_v[`W-1], adh4_v, n_27_v, adh4_port_6, n_27_port_2);
  spice_transistor_nmos t2553(~dpc32_PCHADH_v[`W-1], adh1_v, n_209_v, adh1_port_6, n_209_port_1);
  spice_transistor_nmos t2552(~dpc32_PCHADH_v[`W-1], adh2_v, n_1496_v, adh2_port_6, n_1496_port_2);
  spice_transistor_nmos_gnd t1217(~adl0_v[`W-1], n_123_v, n_123_port_0);
  spice_transistor_nmos t637(~cclk_v[`W-1], y2_v, n_1491_v, y2_port_0, n_1491_port_0);
  spice_transistor_nmos t1208(~dpc20_ADDSB06_v[`W-1], alu6_v, sb6_v, alu6_port_2, sb6_port_6);
  spice_transistor_nmos t1209(~dpc20_ADDSB06_v[`W-1], alu5_v, sb5_v, alu5_port_1, sb5_port_3);
  spice_transistor_nmos_gnd t2357(~n_659_v[`W-1], ab15_v, ab15_port_0);
  spice_transistor_nmos_vdd t2353(~n_298_v[`W-1], db7_v, db7_port_3);
  spice_transistor_nmos_vdd t3016(n_1034_v, n_994_v, n_994_port_3);
  spice_transistor_nmos_gnd t3015(n_1034_v, n_1545_v, n_1545_port_2);
  spice_transistor_nmos_gnd t1947(n_849_v, dpc33_PCHDB_v, dpc33_PCHDB_port_1);
  spice_transistor_nmos_vdd t2942(n_617_v, n_676_v, n_676_port_3);
  spice_transistor_nmos_vdd t2768(n_1026_v, n_171_v, n_171_port_3);
  spice_transistor_nmos_vdd t1410(n_321_v, dpc33_PCHDB_v, dpc33_PCHDB_port_0);
  spice_transistor_nmos_gnd g_4709((~alub3_v[`W-1]&~alua3_v[`W-1]), n_350_v, n_350_port_5);
  spice_transistor_nmos_gnd t64(notalu6_v, alu6_v, alu6_port_0);
  spice_transistor_nmos_gnd t67(notidl2_v, idl2_v, idl2_port_0);
  spice_transistor_nmos t3225(~dpc2_XSB_v[`W-1], n_1709_v, sb1_v, n_1709_port_2, sb1_port_12);
  spice_transistor_nmos t3489(~dpc13_ORS_v[`W-1], aluanorb1_v, notaluoutmux1_v, aluanorb1_port_4, notaluoutmux1_port_5);
  spice_transistor_nmos_vdd t2572(~n_1639_v[`W-1], ab15_v, ab15_port_1);
  spice_transistor_nmos_vdd t2570(n_1541_v, dpc10_ADLADD_v, dpc10_ADLADD_port_5);
  spice_transistor_nmos t2683(~dpc9_DBADD_v[`W-1], alub7_v, idb7_v, alub7_port_0, idb7_port_8);
  spice_transistor_nmos t2684(~dpc9_DBADD_v[`W-1], alub6_v, idb6_v, alub6_port_2, idb6_port_10);
  spice_transistor_nmos t1883(~cclk_v[`W-1], _ABL7_v, n_171_v, _ABL7_port_1, n_171_port_1);
  spice_transistor_nmos_vdd t1880(n_1295_v, dpc25_SBDB_v, dpc25_SBDB_port_9);
  spice_transistor_nmos_gnd t1887(~n_643_v[`W-1], db3_v, db3_port_3);
  spice_transistor_nmos_vdd t2643(n_625_v, dpc3_SBX_v, dpc3_SBX_port_9);
  spice_transistor_nmos_gnd t1082(~dpc12_0ADD_v[`W-1], alua6_v, alua6_port_1);
  spice_transistor_nmos_gnd t1083(~dpc12_0ADD_v[`W-1], alua5_v, alua5_port_1);
  spice_transistor_nmos_gnd t1080(~dpc12_0ADD_v[`W-1], alua1_v, alua1_port_3);
  spice_transistor_nmos_gnd t1081(~dpc12_0ADD_v[`W-1], alua4_v, alua4_port_1);
  spice_transistor_nmos_gnd t1089(~n_37_v[`W-1], db2_v, db2_port_2);
  spice_transistor_nmos_vdd t1991(n_23_v, n_1501_v, n_1501_port_1);
  spice_transistor_nmos_vdd t1516(abh0_v, n_826_v, n_826_port_1);
  spice_transistor_nmos_gnd t1628(pd6_clearIR_v, n_1309_v, n_1309_port_1);
  spice_transistor_nmos_gnd t185(notidl6_v, idl6_v, idl6_port_0);
  spice_transistor_nmos_gnd g_4918(((~__AxB_6_v[`W-1]&C56_v)|_AxB_6__C56_v), __AxBxC_6_v, __AxBxC_6_port_5);
  spice_transistor_nmos_gnd g_4913((~n_975_v[`W-1]|(n_312_v&~cclk_v[`W-1])), n_854_v, n_854_port_6);
  spice_transistor_nmos_gnd g_4916(((n_753_v&n_1135_v)|n_1629_v), dasb5_v, dasb5_port_5);
  spice_transistor_nmos_gnd g_4915(((AxB5_v&_C45_v)|__AxB5__C45_v), __AxBxC_5_v, __AxBxC_5_port_5);
  spice_transistor_nmos t2218(~dpc15_ANDS_v[`W-1], n_336_v, n_722_v, n_336_port_3, n_722_port_5);
  spice_transistor_nmos t2219(~dpc15_ANDS_v[`W-1], n_304_v, n_1318_v, n_304_port_4, n_1318_port_3);
  spice_transistor_nmos t2216(~dpc15_ANDS_v[`W-1], n_1063_v, n_296_v, n_1063_port_4, n_296_port_4);
  spice_transistor_nmos t2217(~dpc15_ANDS_v[`W-1], n_277_v, n_477_v, n_277_port_4, n_477_port_3);
  spice_transistor_nmos t2214(~dpc15_ANDS_v[`W-1], n_681_v, n_740_v, n_681_port_3, n_740_port_4);
  spice_transistor_nmos t2747(~dpc37_PCLDB_v[`W-1], idb7_v, n_1647_v, idb7_port_9, n_1647_port_2);
  spice_transistor_nmos t2212(~dpc15_ANDS_v[`W-1], aluanandb0_v, notaluoutmux0_v, aluanandb0_port_3, notaluoutmux0_port_5);
  spice_transistor_nmos t2213(~dpc15_ANDS_v[`W-1], aluanandb1_v, notaluoutmux1_v, aluanandb1_port_1, notaluoutmux1_port_4);
  spice_transistor_nmos_gnd t2511(~idb3_v[`W-1], n_1621_v, n_1621_port_1);
  spice_transistor_nmos_gnd t896(abh6_v, n_635_v, n_635_port_1);
  spice_transistor_nmos_vdd t894(abh6_v, n_963_v, n_963_port_2);
  spice_transistor_nmos_gnd t1608(n_334_v, Pout2_v, Pout2_port_1);
  spice_transistor_nmos t2554(~dpc32_PCHADH_v[`W-1], adh0_v, n_1722_v, adh0_port_6, n_1722_port_2);
  spice_transistor_nmos t2557(~cclk_v[`W-1], _ABH0_v, n_381_v, _ABH0_port_2, n_381_port_2);
  spice_transistor_nmos_vdd t2000(~n_1633_v[`W-1], ab5_v, ab5_port_1);
  spice_transistor_nmos_gnd g_4937((~n_297_v[`W-1]|(n_284_v&~cclk_v[`W-1])), NMIP_v, NMIP_port_7);
  spice_transistor_nmos_gnd g_4932(((~__AxB_2_v[`W-1]&C12_v)|_AxB_2__C12_v), __AxBxC_2_v, __AxBxC_2_port_5);
  spice_transistor_nmos t2235(~dpc26_ACDB_v[`W-1], n_146_v, idb0_v, n_146_port_1, idb0_port_8);
  spice_transistor_nmos t2236(~dpc26_ACDB_v[`W-1], n_929_v, idb1_v, n_929_port_2, idb1_port_5);
  spice_transistor_nmos t2237(~dpc26_ACDB_v[`W-1], n_1618_v, idb2_v, n_1618_port_0, idb2_port_6);
  spice_transistor_nmos t2238(~dpc26_ACDB_v[`W-1], n_1654_v, idb3_v, n_1654_port_2, idb3_port_6);
  spice_transistor_nmos t2239(~dpc26_ACDB_v[`W-1], idb4_v, n_1344_v, idb4_port_6, n_1344_port_0);
  spice_transistor_nmos t2728(~dpc9_DBADD_v[`W-1], alub5_v, idb5_v, alub5_port_2, idb5_port_8);
  spice_transistor_nmos t2729(~dpc9_DBADD_v[`W-1], alub4_v, idb4_v, alub4_port_3, idb4_port_8);
  spice_transistor_nmos t2726(~dpc9_DBADD_v[`W-1], alub3_v, idb3_v, alub3_port_3, idb3_port_8);
  spice_transistor_nmos t2727(~dpc9_DBADD_v[`W-1], idb2_v, alub2_v, idb2_port_9, alub2_port_4);
  spice_transistor_nmos t2724(~cp1_v[`W-1], n_1147_v, idl7_v, n_1147_port_3, idl7_port_1);
  spice_transistor_nmos t2725(~dpc9_DBADD_v[`W-1], alub1_v, idb1_v, alub1_port_1, idb1_port_7);
  spice_transistor_nmos_gnd t422(~n_135_v[`W-1], clk2out_v, clk2out_port_1);
  spice_transistor_nmos_vdd t426(~cclk_v[`W-1], adh4_v, adh4_port_2);
  spice_transistor_nmos_vdd t427(~cclk_v[`W-1], adl5_v, adl5_port_0);
  spice_transistor_nmos_gnd g_4335((~cclk_v[`W-1]|n_71_v|~n_1247_v[`W-1]), dpc7_SS_v, dpc7_SS_port_12);
  spice_transistor_nmos g_4746((~ADL_ABL_v[`W-1]&~cp1_v[`W-1]), _ABL0_v, n_123_v, _ABL0_port_3, n_123_port_3);
  spice_transistor_nmos t226(~dpc7_SS_v[`W-1], n_332_v, s0_v, n_332_port_0, s0_port_0);
  spice_transistor_nmos_vdd t227(~cclk_v[`W-1], idb0_v, idb0_port_1);
  spice_transistor_nmos_gnd t25(abl0_v, n_1100_v, n_1100_port_0);
  spice_transistor_nmos_vdd t27(abl0_v, n_855_v, n_855_port_0);
  spice_transistor_nmos_gnd t2537(n_0_ADL2_v, adl2_v, adl2_port_6);
  spice_transistor_nmos t2535(~cclk_v[`W-1], n_635_v, _ABH6_v, n_635_port_3, _ABH6_port_2);
  spice_transistor_nmos t2532(~dpc38_PCLADL_v[`W-1], n_723_v, adl3_v, n_723_port_1, adl3_port_4);
  spice_transistor_nmos t2531(~dpc38_PCLADL_v[`W-1], adl2_v, n_481_v, adl2_port_5, n_481_port_2);
  spice_transistor_nmos t2530(~dpc38_PCLADL_v[`W-1], n_976_v, adl1_v, n_976_port_0, adl1_port_5);
  spice_transistor_nmos_gnd t2777(n_842_v, n_1479_v, n_1479_port_1);
  spice_transistor_nmos t1848(~dpc23_SBAC_v[`W-1], dasb7_v, a7_v, dasb7_port_1, a7_port_2);
  spice_transistor_nmos t1846(~dpc23_SBAC_v[`W-1], dasb5_v, a5_v, dasb5_port_1, a5_port_2);
  spice_transistor_nmos t1847(~dpc23_SBAC_v[`W-1], dasb6_v, a6_v, dasb6_port_0, a6_port_2);
  spice_transistor_nmos t1844(~dpc23_SBAC_v[`W-1], dasb3_v, a3_v, dasb3_port_1, a3_port_1);
  spice_transistor_nmos t1845(~dpc23_SBAC_v[`W-1], sb4_v, a4_v, sb4_port_7, a4_port_0);
  spice_transistor_nmos t1842(~dpc23_SBAC_v[`W-1], dasb1_v, a1_v, dasb1_port_0, a1_port_1);
  spice_transistor_nmos t1843(~dpc23_SBAC_v[`W-1], a2_v, dasb2_v, a2_port_1, dasb2_port_1);
  spice_transistor_nmos t1841(~dpc23_SBAC_v[`W-1], sb0_v, a0_v, sb0_port_5, a0_port_1);
  spice_transistor_nmos_gnd g_4483((n_964_v|n_732_v), clock1_v, clock1_port_68);
  spice_transistor_nmos_gnd g_4489((n_769_v|~RnWstretched_v[`W-1]), n_1325_v, n_1325_port_4);
  spice_transistor_nmos_gnd t2437(~n_1696_v[`W-1], rw_v, rw_port_1);
  spice_transistor_nmos_gnd t440(n_400_v, n_102_v, n_102_port_0);
  spice_transistor_nmos_vdd t441(n_400_v, n_1696_v, n_1696_port_0);
  spice_transistor_nmos_gnd t442(n_834_v, n_1696_v, n_1696_port_1);
  spice_transistor_nmos_vdd t446(~n_1545_v[`W-1], ab10_v, ab10_port_0);
  spice_transistor_nmos_vdd t2873(n_1315_v, n_381_v, n_381_port_3);
  spice_transistor_nmos_vdd t1477(n_17_v, clock1_v, clock1_port_40);
  spice_transistor_nmos_gnd t205(~n_999_v[`W-1], ab12_v, ab12_port_0);
  spice_transistor_nmos_vdd t3399(~n_1479_v[`W-1], ab1_v, ab1_port_1);
  spice_transistor_nmos t3391(~dpc6_SBS_v[`W-1], s7_v, sb7_v, s7_port_2, sb7_port_11);
  spice_transistor_nmos_gnd t3392(~n_642_v[`W-1], ab2_v, ab2_port_1);
  spice_transistor_nmos_gnd t1865(n_1194_v, Pout3_v, Pout3_port_2);
  spice_transistor_nmos t1860(~dpc25_SBDB_v[`W-1], idb5_v, sb5_v, idb5_port_4, sb5_port_6);
  spice_transistor_nmos t1861(~dpc25_SBDB_v[`W-1], idb6_v, sb6_v, idb6_port_5, sb6_port_8);
  spice_transistor_nmos t1862(~dpc25_SBDB_v[`W-1], sb7_v, idb7_v, sb7_port_5, idb7_port_4);
  spice_transistor_nmos_gnd t1397(notalu1_v, alu1_v, alu1_port_1);
  spice_transistor_nmos t589(~dpc43_DL_DB_v[`W-1], idb4_v, n_1095_v, idb4_port_0, n_1095_port_1);
  spice_transistor_nmos t587(~dpc43_DL_DB_v[`W-1], idb2_v, n_1424_v, idb2_port_1, n_1424_port_2);
  spice_transistor_nmos t586(~dpc43_DL_DB_v[`W-1], idb1_v, n_87_v, idb1_port_0, n_87_port_2);
  spice_transistor_nmos_gnd g_4465((~RnWstretched_v[`W-1]|n_23_v), n_298_v, n_298_port_4);
  spice_transistor_nmos t2278(~cclk_v[`W-1], n_927_v, notir4_v, n_927_port_1, notir4_port_24);
  spice_transistor_nmos_vdd t2270(~cclk_v[`W-1], idb5_v, idb5_port_6);
  spice_transistor_nmos_gnd t2276(pclp4_v, n_208_v, n_208_port_0);
  spice_transistor_nmos_vdd t466(n_35_v, dpc7_SS_v, dpc7_SS_port_7);
  spice_transistor_nmos_vdd t460(abl3_v, n_1041_v, n_1041_port_0);
  spice_transistor_nmos t268(H1x1_v, idb0_v, Pout0_v, idb0_port_2, Pout0_port_0);
  spice_transistor_nmos g_4694((~ADL_ABL_v[`W-1]&~cp1_v[`W-1]), _ABL5_v, n_1094_v, _ABL5_port_3, n_1094_port_3);
  spice_transistor_nmos_gnd t1706(ir1_v, notir1_v, notir1_port_21);
  spice_transistor_nmos g_4690((~ADL_ABL_v[`W-1]&~cp1_v[`W-1]), _ABL6_v, n_1548_v, _ABL6_port_3, n_1548_port_3);
  spice_transistor_nmos g_4693((~ADL_ABL_v[`W-1]&~cp1_v[`W-1]), _ABL7_v, n_1046_v, _ABL7_port_3, n_1046_port_3);
  spice_transistor_nmos g_4692((~ADL_ABL_v[`W-1]&~cp1_v[`W-1]), _ABL4_v, n_1519_v, _ABL4_port_3, n_1519_port_3);
  spice_transistor_nmos_vdd t1701(~n_475_v[`W-1], ab12_v, ab12_port_1);
  spice_transistor_nmos_gnd t1709(n_1399_v, n_1105_v, n_1105_port_2);
  spice_transistor_nmos_vdd t3407(n_355_v, dpc4_SSB_v, dpc4_SSB_port_9);
  spice_transistor_nmos_vdd t877(n_692_v, dpc1_SBY_v, dpc1_SBY_port_3);
  spice_transistor_nmos_vdd t870(n_291_v, dpc41_DL_ADL_v, dpc41_DL_ADL_port_0);
  spice_transistor_nmos t2130(H1x1_v, p6_v, idb6_v, p6_port_0, idb6_port_6);
  spice_transistor_nmos_vdd t1118(~cclk_v[`W-1], sb3_v, sb3_port_3);
  spice_transistor_nmos t1110(~dpc17_SUMS_v[`W-1], __AxBxC_4_v, n_296_v, __AxBxC_4_port_2, n_296_port_1);
  spice_transistor_nmos t1111(~dpc17_SUMS_v[`W-1], __AxBxC_5_v, n_277_v, __AxBxC_5_port_1, n_277_port_2);
  spice_transistor_nmos t1112(~dpc17_SUMS_v[`W-1], n_722_v, __AxBxC_6_v, n_722_port_2, __AxBxC_6_port_1);
  spice_transistor_nmos t1113(~dpc17_SUMS_v[`W-1], n_304_v, __AxBxC_7_v, n_304_port_2, __AxBxC_7_port_0);
  spice_transistor_nmos_gnd g_4509((~n_1247_v[`W-1]|n_1043_v|~cclk_v[`W-1]), dpc40_ADLPCL_v, dpc40_ADLPCL_port_12);
  spice_transistor_nmos_gnd t2012(n_1323_v, dpc37_PCLDB_v, dpc37_PCLDB_port_4);
  spice_transistor_nmos_gnd t2013(pchp7_v, n_1206_v, n_1206_port_0);
  spice_transistor_nmos t1507(~cclk_v[`W-1], n_146_v, a0_v, n_146_port_0, a0_port_0);
  spice_transistor_nmos_gnd t3351(~adh7_v[`W-1], n_494_v, n_494_port_1);
  spice_transistor_nmos_gnd t3357(n_184_v, n_1531_v, n_1531_port_2);
  spice_transistor_nmos_gnd g_4818((~alub1_v[`W-1]&~alua1_v[`W-1]), aluanandb1_v, aluanandb1_port_5);
  spice_transistor_nmos_gnd t1566(n_128_v, n_1592_v, n_1592_port_1);
  spice_transistor_nmos_gnd t1561(~n_210_v[`W-1], ab5_v, ab5_port_0);
  spice_transistor_nmos t248(~dpc6_SBS_v[`W-1], s5_v, sb5_v, s5_port_0, sb5_port_1);
  spice_transistor_nmos t249(~dpc6_SBS_v[`W-1], s6_v, sb6_v, s6_port_0, sb6_port_3);
  spice_transistor_nmos t241(~cclk_v[`W-1], n_326_v, a6_v, n_326_port_0, a6_port_0);
  spice_transistor_nmos_gnd t2767(n_1026_v, n_322_v, n_322_port_2);
  spice_transistor_nmos_vdd t2764(n_611_v, dpc31_PCHPCH_v, dpc31_PCHPCH_port_11);
  spice_transistor_nmos t2762(~cp1_v[`W-1], n_1661_v, idl3_v, n_1661_port_3, idl3_port_1);
  spice_transistor_nmos_gnd t2760(pd4_clearIR_v, n_227_v, n_227_port_0);
  spice_transistor_nmos t1829(~cclk_v[`W-1], n_119_v, notir1_v, n_119_port_0, notir1_port_22);
  spice_transistor_nmos t2482(~dpc31_PCHPCH_v[`W-1], pch1_v, n_209_v, pch1_port_2, n_209_port_0);
  spice_transistor_nmos t2481(~dpc31_PCHPCH_v[`W-1], pch0_v, n_1722_v, pch0_port_2, n_1722_port_1);
  spice_transistor_nmos t2480(~dpc31_PCHPCH_v[`W-1], pch3_v, n_141_v, pch3_port_2, n_141_port_1);
  spice_transistor_nmos_gnd t2487(~dpc29_0ADH17_v[`W-1], adh5_v, adh5_port_3);
  spice_transistor_nmos_gnd t2486(~dpc29_0ADH17_v[`W-1], adh2_v, adh2_port_5);
  spice_transistor_nmos_gnd t2485(~dpc29_0ADH17_v[`W-1], adh3_v, adh3_port_5);
  spice_transistor_nmos t2334(~dpc37_PCLDB_v[`W-1], idb4_v, n_208_v, idb4_port_7, n_208_port_1);
  spice_transistor_nmos_gnd t2488(~dpc29_0ADH17_v[`W-1], adh4_v, adh4_port_5);
  spice_transistor_nmos t1350(~cclk_v[`W-1], _ABL0_v, n_1100_v, _ABL0_port_2, n_1100_port_2);
  spice_transistor_nmos_vdd t2153(n_1534_v, dpc8_nDBADD_v, dpc8_nDBADD_port_6);
  spice_transistor_nmos_vdd t2157(~n_417_v[`W-1], sync_v, sync_port_1);
  spice_transistor_nmos_gnd g_4528((~RnWstretched_v[`W-1]|dor0_v), n_1072_v, n_1072_port_4);
  spice_transistor_nmos_gnd g_4425((dor4_v|~RnWstretched_v[`W-1]), n_147_v, n_147_port_4);
  spice_transistor_nmos_vdd t1686(n_476_v, dpc12_0ADD_v, dpc12_0ADD_port_9);
  spice_transistor_nmos_gnd t1682(n_1471_v, p4_v, p4_port_0);
  spice_transistor_nmos_vdd t382(~n_1076_v[`W-1], db4_v, db4_port_0);
  spice_transistor_nmos t385(~dpc4_SSB_v[`W-1], n_280_v, sb5_v, n_280_port_1, sb5_port_2);
  spice_transistor_nmos_gnd t3147(abl4_v, n_86_v, n_86_port_3);
  spice_transistor_nmos t3142(~dpc0_YSB_v[`W-1], n_767_v, sb1_v, n_767_port_2, sb1_port_11);
  spice_transistor_nmos_vdd t3149(abl4_v, n_634_v, n_634_port_1);
  spice_transistor_nmos_vdd t2818(dor6_v, n_7_v, n_7_port_2);
  spice_transistor_nmos_gnd t2819(n_0_ADL0_v, adl0_v, adl0_port_7);
  spice_transistor_nmos_vdd t1548(~cclk_v[`W-1], sb7_v, sb7_port_3);
  spice_transistor_nmos_gnd t3332(pd1_clearIR_v, n_1641_v, n_1641_port_1);
  spice_transistor_nmos_gnd t2669(~n_206_v[`W-1], n_465_v, n_465_port_0);
  spice_transistor_nmos_gnd g_4544((n_225_v|~n_1247_v[`W-1]|~cclk_v[`W-1]), dpc9_DBADD_v, dpc9_DBADD_port_12);
  spice_transistor_nmos_gnd t1379(pchp5_v, n_1301_v, n_1301_port_0);
  spice_transistor_nmos_gnd g_4400((n_466_v|~RnWstretched_v[`W-1]), n_7_v, n_7_port_4);
  spice_transistor_nmos_gnd t1388(notalu0_v, alu0_v, alu0_port_1);
  spice_transistor_nmos t2785(~cclk_v[`W-1], _ABL4_v, n_86_v, _ABL4_port_1, n_86_port_2);
  spice_transistor_nmos_gnd g_4396((n_491_v|~cclk_v[`W-1]|~n_1247_v[`W-1]), dpc10_ADLADD_v, dpc10_ADLADD_port_12);
  spice_transistor_nmos_gnd t3163(n_617_v, n_1140_v, n_1140_port_2);
  spice_transistor_nmos_gnd t992(abh5_v, n_869_v, n_869_port_1);
  spice_transistor_nmos t993(~dpc37_PCLDB_v[`W-1], idb2_v, n_481_v, idb2_port_3, n_481_port_1);
  spice_transistor_nmos_vdd t990(abh5_v, n_1608_v, n_1608_port_1);
  spice_transistor_nmos t1529(~dpc3_SBX_v[`W-1], x5_v, sb5_v, x5_port_1, sb5_port_4);
  spice_transistor_nmos t1528(~dpc3_SBX_v[`W-1], sb6_v, x6_v, sb6_port_7, x6_port_1);
  spice_transistor_nmos_vdd t1521(n_1677_v, n_999_v, n_999_port_1);
  spice_transistor_nmos_gnd t1520(n_1677_v, n_475_v, n_475_port_0);
  spice_transistor_nmos t1525(~dpc3_SBX_v[`W-1], x2_v, sb2_v, x2_port_1, sb2_port_4);
  spice_transistor_nmos t1524(~dpc3_SBX_v[`W-1], x3_v, sb3_v, x3_port_1, sb3_port_6);
  spice_transistor_nmos_vdd t1527(n_582_v, ADH_ABH_v, ADH_ABH_port_4);
  spice_transistor_nmos_vdd t1344(n_1715_v, n_1105_v, n_1105_port_0);
  spice_transistor_nmos t3316(~cclk_v[`W-1], y0_v, n_564_v, y0_port_2, n_564_port_2);
  spice_transistor_nmos t3317(~cclk_v[`W-1], n_659_v, _ABH7_v, n_659_port_3, _ABH7_port_2);
  spice_transistor_nmos_vdd t3313(n_1463_v, n_147_v, n_147_port_3);
  spice_transistor_nmos_vdd t176(n_714_v, dpc19_ADDSB7_v, dpc19_ADDSB7_port_0);
  spice_transistor_nmos t170(~cclk_v[`W-1], _ABL5_v, n_210_v, _ABL5_port_0, n_210_port_0);
  spice_transistor_nmos t2371(~dpc5_SADL_v[`W-1], adl1_v, n_694_v, adl1_port_4, n_694_port_3);
  spice_transistor_nmos t2370(~dpc24_ACSB_v[`W-1], n_1592_v, sb7_v, n_1592_port_3, sb7_port_9);
  spice_transistor_nmos_gnd t2373(pchp0_v, n_1722_v, n_1722_port_0);
  spice_transistor_nmos t2372(~cclk_v[`W-1], _ABL2_v, n_642_v, _ABL2_port_2, n_642_port_1);
  spice_transistor_nmos_gnd t507(~n_1100_v[`W-1], ab0_v, ab0_port_0);
  spice_transistor_nmos_gnd t501(n_1676_v, n_634_v, n_634_port_0);
  spice_transistor_nmos t503(~cclk_v[`W-1], notir0_v, n_310_v, notir0_port_1, n_310_port_0);
  spice_transistor_nmos_vdd t502(n_1676_v, n_86_v, n_86_port_0);
  spice_transistor_nmos t2199(~dpc27_SBADH_v[`W-1], adh2_v, sb2_v, adh2_port_4, sb2_port_8);
  spice_transistor_nmos t2198(~dpc27_SBADH_v[`W-1], adh3_v, sb3_v, adh3_port_3, sb3_port_9);
  spice_transistor_nmos_gnd t2195(~cp1_v[`W-1], n_1247_v, n_1247_port_13);
  spice_transistor_nmos t2191(~dpc27_SBADH_v[`W-1], sb6_v, adh6_v, sb6_port_9, adh6_port_3);
  spice_transistor_nmos t2190(~dpc27_SBADH_v[`W-1], adh7_v, sb7_v, adh7_port_3, sb7_port_7);
  spice_transistor_nmos t2193(~dpc27_SBADH_v[`W-1], adh0_v, sb0_v, adh0_port_2, sb0_port_9);
  spice_transistor_nmos t2192(~dpc1_SBY_v[`W-1], y0_v, sb0_v, y0_port_0, sb0_port_8);
  spice_transistor_nmos_gnd g_4563((~alub5_v[`W-1]|~alua5_v[`W-1]), n_1632_v, n_1632_port_7);
  spice_transistor_nmos t1315(~cclk_v[`W-1], _ABL3_v, n_138_v, _ABL3_port_0, n_138_port_2);
  spice_transistor_nmos t1165(~dpc8_nDBADD_v[`W-1], alub2_v, n_458_v, alub2_port_0, n_458_port_1);
  spice_transistor_nmos t1164(~dpc8_nDBADD_v[`W-1], alub4_v, n_478_v, alub4_port_0, n_478_port_0);
  spice_transistor_nmos_gnd t349(ir0_v, notir0_v, notir0_port_0);
  spice_transistor_nmos_vdd t345(n_525_v, dpc26_ACDB_v, dpc26_ACDB_port_0);
  spice_transistor_nmos_gnd t343(n_1305_v, dpc17_SUMS_v, dpc17_SUMS_port_0);
  spice_transistor_nmos_gnd g_4825((~alua7_v[`W-1]&~alub7_v[`W-1]), n_1318_v, n_1318_port_7);
  spice_transistor_nmos_gnd g_4823((~n_681_v[`W-1]&n_110_v), __AxB_2_v, __AxB_2_port_7);
  spice_transistor_nmos g_4821((~cp1_v[`W-1]&fetch_v), n_227_v, n_927_v, n_227_port_3, n_927_port_3);
  spice_transistor_nmos_gnd t3103(~n_1254_v[`W-1], ab6_v, ab6_port_1);
  spice_transistor_nmos t1508(~dpc0_YSB_v[`W-1], sb3_v, n_1531_v, sb3_port_5, n_1531_port_0);
  spice_transistor_nmos_gnd g_4615((~alua1_v[`W-1]|~alub1_v[`W-1]), aluanorb1_v, aluanorb1_port_7);
  spice_transistor_nmos_gnd g_4614((~cclk_v[`W-1]|n_662_v|~n_1247_v[`W-1]), dpc3_SBX_v, dpc3_SBX_port_12);
  spice_transistor_nmos t3376(~dpc40_ADLPCL_v[`W-1], adl2_v, pcl2_v, adl2_port_8, pcl2_port_2);
  spice_transistor_nmos t3377(~dpc40_ADLPCL_v[`W-1], pcl5_v, adl5_v, pcl5_port_2, adl5_port_7);
  spice_transistor_nmos t3374(~dpc40_ADLPCL_v[`W-1], adl0_v, pcl0_v, adl0_port_8, pcl0_port_2);
  spice_transistor_nmos t3378(~dpc40_ADLPCL_v[`W-1], adl4_v, pcl4_v, adl4_port_7, pcl4_port_2);
  spice_transistor_nmos t3379(~dpc40_ADLPCL_v[`W-1], adl6_v, pcl6_v, adl6_port_7, pcl6_port_2);
  spice_transistor_nmos_vdd t154(~n_798_v[`W-1], db1_v, db1_port_1);
  spice_transistor_nmos_gnd t158(~adl6_v[`W-1], n_1548_v, n_1548_port_1);
  spice_transistor_nmos_gnd t1404(nots3_v, n_998_v, n_998_port_2);
  spice_transistor_nmos_gnd t2424(n_1255_v, dpc13_ORS_v, dpc13_ORS_port_5);
  spice_transistor_nmos_gnd g_4589((n_282_v|~cclk_v[`W-1]|~n_1247_v[`W-1]), dpc6_SBS_v, dpc6_SBS_port_12);
  spice_transistor_nmos_gnd g_4584((~alub4_v[`W-1]|~alua4_v[`W-1]), n_404_v, n_404_port_6);
  spice_transistor_nmos t1338(~dpc3_SBX_v[`W-1], x1_v, sb1_v, x1_port_1, sb1_port_4);
  spice_transistor_nmos_gnd t1999(n_1129_v, n_1467_v, n_1467_port_1);
  spice_transistor_nmos t1331(~cclk_v[`W-1], n_831_v, a5_v, n_831_port_0, a5_port_0);
  spice_transistor_nmos t1333(H1x1_v, Pout1_v, idb1_v, Pout1_port_0, idb1_port_3);
  spice_transistor_nmos_gnd t1334(n_172_v, n_1633_v, n_1633_port_0);
  spice_transistor_nmos_vdd t1335(n_172_v, n_210_v, n_210_port_1);
  spice_transistor_nmos_vdd t367(n_424_v, notRdy0_v, notRdy0_port_3);
  spice_transistor_nmos_vdd t362(n_1129_v, cclk_v, cclk_port_28);
  spice_transistor_nmos_gnd t369(n_198_v, notRdy0_v, notRdy0_port_4);
  spice_transistor_nmos_gnd g_4800((~alua2_v[`W-1]&~alub2_v[`W-1]), n_681_v, n_681_port_8);
  spice_transistor_nmos g_4803((~ADH_ABH_v[`W-1]&~cp1_v[`W-1]), _ABH5_v, n_254_v, _ABH5_port_3, n_254_port_3);
  spice_transistor_nmos_gnd g_4808((n_803_v&~n_336_v[`W-1]), __AxB_6_v, __AxB_6_port_11);
  spice_transistor_nmos_gnd g_4809((~alub0_v[`W-1]&~alua0_v[`W-1]), aluanandb0_v, aluanandb0_port_9);
  spice_transistor_nmos_gnd t3125(ir5_v, notir5_v, notir5_port_36);
  spice_transistor_nmos_gnd t3123(n_1719_v, n_831_v, n_831_port_3);
  spice_transistor_nmos_vdd t3122(n_224_v, n_37_v, n_37_port_3);
  spice_transistor_nmos t3120(~dpc2_XSB_v[`W-1], n_436_v, sb4_v, n_436_port_2, sb4_port_12);
  spice_transistor_nmos_vdd t2651(dor0_v, n_1325_v, n_1325_port_2);
  spice_transistor_nmos_gnd t2658(~n_359_v[`W-1], ab11_v, ab11_port_1);
  spice_transistor_nmos_gnd t1078(~dpc12_0ADD_v[`W-1], alua0_v, alua0_port_1);
  spice_transistor_nmos_gnd t1627(n_747_v, n_1417_v, n_1417_port_2);
  spice_transistor_nmos t1621(~cclk_v[`W-1], n_1254_v, _ABL6_v, n_1254_port_1, _ABL6_port_1);
  spice_transistor_nmos_vdd t3352(~cclk_v[`W-1], adh6_v, adh6_port_6);
  spice_transistor_nmos_vdd t3353(~cclk_v[`W-1], adl7_v, adl7_port_7);
  spice_transistor_nmos_gnd t3355(pclp1_v, n_976_v, n_976_port_3);
  spice_transistor_nmos_vdd t935(n_1593_v, dpc14_SRS_v, dpc14_SRS_port_1);
  spice_transistor_nmos_vdd t130(n_1369_v, dpc38_PCLADL_v, dpc38_PCLADL_port_0);
  spice_transistor_nmos t132(~dpc4_SSB_v[`W-1], n_721_v, sb7_v, n_721_port_0, sb7_port_0);
  spice_transistor_nmos t133(~dpc4_SSB_v[`W-1], n_618_v, sb6_v, n_618_port_0, sb6_port_2);
  spice_transistor_nmos_vdd t135(n_818_v, dpc40_ADLPCL_v, dpc40_ADLPCL_port_0);
  spice_transistor_nmos t136(~dpc4_SSB_v[`W-1], n_3_v, sb4_v, n_3_port_0, sb4_port_3);
  spice_transistor_nmos_gnd t2674(abl5_v, n_210_v, n_210_port_3);
  spice_transistor_nmos_vdd t2676(abl5_v, n_1633_v, n_1633_port_2);
  spice_transistor_nmos_gnd t540(n_1635_v, dpc29_0ADH17_v, dpc29_0ADH17_port_1);
  spice_transistor_nmos t546(~dpc13_ORS_v[`W-1], n_649_v, n_1071_v, n_649_port_0, n_1071_port_0);
  spice_transistor_nmos_vdd t1712(~n_1325_v[`W-1], db0_v, db0_port_1);
  spice_transistor_nmos_gnd t301(~n_612_v[`W-1], db5_v, db5_port_0);
  spice_transistor_nmos_gnd t300(n_730_v, n_1724_v, n_1724_port_0);
  spice_transistor_nmos_gnd t309(n_445_v, n_417_v, n_417_port_0);
  spice_transistor_nmos g_4791((~ADL_ABL_v[`W-1]&~cp1_v[`W-1]), _ABL2_v, n_935_v, _ABL2_port_3, n_935_port_3);
  spice_transistor_nmos_gnd g_4792((n_918_v&~n_1063_v[`W-1]), __AxB_4_v, __AxB_4_port_6);
  spice_transistor_nmos g_4862((~cp1_v[`W-1]&fetch_v), n_1309_v, n_1675_v, n_1309_port_3, n_1675_port_3);
  spice_transistor_nmos g_4860((~cp1_v[`W-1]&~ADH_ABH_v[`W-1]), n_212_v, _ABH4_v, n_212_port_3, _ABH4_port_3);
  spice_transistor_nmos g_4861((~cp1_v[`W-1]&fetch_v), n_928_v, n_1609_v, n_928_port_3, n_1609_port_3);
  spice_transistor_nmos g_4865((~cp1_v[`W-1]&fetch_v), n_571_v, n_1300_v, n_571_port_3, n_1300_port_3);
  spice_transistor_nmos_gnd t2090(n_981_v, n_733_v, n_733_port_0);
  spice_transistor_nmos t2091(~cclk_v[`W-1], _ABL1_v, n_66_v, _ABL1_port_2, n_66_port_2);
  spice_transistor_nmos_vdd t2092(abh4_v, n_475_v, n_475_port_2);
  spice_transistor_nmos_gnd t2094(abh4_v, n_999_v, n_999_port_2);
  spice_transistor_nmos t1273(n_1446_v, n_430_v, n_206_v, n_430_port_1, n_206_port_3);
  spice_transistor_nmos t936(~dpc16_EORS_v[`W-1], __AxB_0_v, notaluoutmux0_v, __AxB_0_port_2, notaluoutmux0_port_0);
  spice_transistor_nmos t937(~dpc16_EORS_v[`W-1], notaluoutmux1_v, n_953_v, notaluoutmux1_port_0, n_953_port_0);
  spice_transistor_nmos t938(~dpc16_EORS_v[`W-1], __AxB_2_v, n_740_v, __AxB_2_port_0, n_740_port_1);
  spice_transistor_nmos t939(~dpc16_EORS_v[`W-1], n_884_v, n_1071_v, n_884_port_1, n_1071_port_2);
  spice_transistor_nmos_gnd t2678(~cp1_v[`W-1], n_43_v, n_43_port_13);
  spice_transistor_nmos_gnd t2890(pchp1_v, n_209_v, n_209_port_2);
  spice_transistor_nmos t2895(~dpc20_ADDSB06_v[`W-1], alu1_v, sb1_v, alu1_port_3, sb1_port_10);
  spice_transistor_nmos t2897(~dpc20_ADDSB06_v[`W-1], alu0_v, sb0_v, alu0_port_2, sb0_port_11);
  spice_transistor_nmos t1010(~cclk_v[`W-1], n_1675_v, notir6_v, n_1675_port_0, notir6_port_1);
  spice_transistor_nmos t1015(~cclk_v[`W-1], n_929_v, a1_v, n_929_port_0, a1_port_0);
  spice_transistor_nmos_gnd t2339(nots0_v, n_332_v, n_332_port_2);
  spice_transistor_nmos_vdd t2336(~cclk_v[`W-1], adh3_v, adh3_port_4);
  spice_transistor_nmos_gnd t112(~dpc12_0ADD_v[`W-1], alua3_v, alua3_port_1);
  spice_transistor_nmos_gnd t111(abh3_v, n_359_v, n_359_port_0);
  spice_transistor_nmos_gnd t2461(AxB5_v, n_1469_v, n_1469_port_1);
  spice_transistor_nmos_gnd t2469(n_709_v, dpc18__DAA_v, dpc18__DAA_port_2);
  spice_transistor_nmos_vdd t2468(n_133_v, dpc2_XSB_v, dpc2_XSB_port_2);
  spice_transistor_nmos_gnd t2565(abl6_v, n_1254_v, n_1254_port_2);
  spice_transistor_nmos_vdd t2567(abl6_v, n_1191_v, n_1191_port_2);
  spice_transistor_nmos_vdd t2560(~n_1041_v[`W-1], ab3_v, ab3_port_0);
  spice_transistor_nmos_vdd t2280(n_628_v, dpc24_ACSB_v, dpc24_ACSB_port_1);
  spice_transistor_nmos t1484(~dpc41_DL_ADL_v[`W-1], adl2_v, n_1424_v, adl2_port_2, n_1424_port_3);
  spice_transistor_nmos_vdd t1739(~cclk_v[`W-1], sb1_v, sb1_port_6);
  spice_transistor_nmos_gnd t1735(notidl7_v, idl7_v, idl7_port_0);
  spice_transistor_nmos t329(~dpc0_YSB_v[`W-1], n_564_v, sb0_v, n_564_port_0, sb0_port_1);
  spice_transistor_nmos t321(~dpc21_ADDADL_v[`W-1], alu2_v, adl2_v, alu2_port_0, adl2_port_0);
  spice_transistor_nmos t323(~dpc21_ADDADL_v[`W-1], adl0_v, alu0_v, adl0_port_0, alu0_port_0);
  spice_transistor_nmos t322(~dpc21_ADDADL_v[`W-1], adl1_v, alu1_v, adl1_port_0, alu1_port_0);
  spice_transistor_nmos g_4840((~cp1_v[`W-1]&fetch_v), n_409_v, n_310_v, n_409_port_5, n_310_port_3);
  spice_transistor_nmos_gnd t2076(abh0_v, n_381_v, n_381_port_1);
  spice_transistor_nmos_gnd t1253(n_31_v, Pout0_v, Pout0_port_1);
  spice_transistor_nmos_vdd t1254(dor3_v, n_42_v, n_42_port_0);
  spice_transistor_nmos_vdd t918(n_1195_v, n_1254_v, n_1254_port_0);
  spice_transistor_nmos_gnd t917(n_1195_v, n_1191_v, n_1191_port_0);
  spice_transistor_nmos_gnd t914(nots7_v, n_721_v, n_721_port_2);
  spice_transistor_nmos_gnd t2613(n_1315_v, n_826_v, n_826_port_2);
  spice_transistor_nmos_gnd t2611(n_556_v, n_1344_v, n_1344_port_2);
  spice_transistor_nmos t2616(~cclk_v[`W-1], n_733_v, y5_v, n_733_port_2, y5_port_1);
  spice_transistor_nmos_vdd t1035(n_358_v, n_1467_v, n_1467_port_0);
  spice_transistor_nmos_gnd t2677(n_419_v, n_1618_v, n_1618_port_2);
  spice_transistor_nmos_gnd g_4677((~alub3_v[`W-1]|~alua3_v[`W-1]), n_649_v, n_649_port_7);
  spice_transistor_nmos_gnd g_4676((~alub6_v[`W-1]|~alua6_v[`W-1]), n_1084_v, n_1084_port_6);
  spice_transistor_nmos_gnd g_4674((~RnWstretched_v[`W-1]|dor1_v), n_794_v, n_794_port_4);
  spice_transistor_nmos t2215(~dpc15_ANDS_v[`W-1], n_350_v, n_1071_v, n_350_port_3, n_1071_port_5);
  spice_transistor_nmos_gnd t2442(dpc28_0ADH0_v, adh0_v, adh0_port_3);
  spice_transistor_nmos_gnd t3066(n_1462_v, dpc38_PCLADL_v, dpc38_PCLADL_port_9);
  spice_transistor_nmos_gnd t3064(~adl2_v[`W-1], n_935_v, n_935_port_1);
  spice_transistor_nmos_gnd t3065(n_5_v, n_146_v, n_146_port_3);
  spice_transistor_nmos t2919(~cclk_v[`W-1], _ABH5_v, n_869_v, _ABH5_port_2, n_869_port_3);
  spice_transistor_nmos t2918(~dpc33_PCHDB_v[`W-1], idb7_v, n_1206_v, idb7_port_10, n_1206_port_3);
  spice_transistor_nmos t2915(~dpc33_PCHDB_v[`W-1], n_27_v, idb4_v, n_27_port_3, idb4_port_9);
  spice_transistor_nmos t2914(~dpc33_PCHDB_v[`W-1], n_141_v, idb3_v, n_141_port_3, idb3_port_10);
  spice_transistor_nmos t2917(~dpc33_PCHDB_v[`W-1], idb6_v, n_652_v, idb6_port_11, n_652_port_3);
  spice_transistor_nmos t2916(~dpc33_PCHDB_v[`W-1], n_1301_v, idb5_v, n_1301_port_3, idb5_port_9);
  spice_transistor_nmos t2911(~dpc33_PCHDB_v[`W-1], n_1722_v, idb0_v, n_1722_port_3, idb0_port_10);
  spice_transistor_nmos t2913(~dpc33_PCHDB_v[`W-1], idb2_v, n_1496_v, idb2_port_10, n_1496_port_3);
  spice_transistor_nmos t2912(~dpc33_PCHDB_v[`W-1], idb1_v, n_209_v, idb1_port_9, n_209_port_3);
  spice_transistor_nmos_gnd t1939(n_318_v, Pout1_v, Pout1_port_1);
  spice_transistor_nmos_vdd t1934(n_466_v, n_471_v, n_471_port_3);
  spice_transistor_nmos_gnd t495(pd3_clearIR_v, n_1083_v, n_1083_port_1);
  spice_transistor_nmos_gnd t491(~adh6_v[`W-1], n_880_v, n_880_port_0);
  spice_transistor_nmos t490(~dpc7_SS_v[`W-1], s7_v, n_721_v, s7_port_0, n_721_port_1);
  spice_transistor_nmos t499(~dpc13_ORS_v[`W-1], n_722_v, n_1084_v, n_722_port_0, n_1084_port_0);
  spice_transistor_nmos t1752(~cp1_v[`W-1], n_1014_v, idl6_v, n_1014_port_3, idl6_port_1);
  spice_transistor_nmos_vdd t1750(~cclk_v[`W-1], adl2_v, adl2_port_4);
  spice_transistor_nmos_vdd t1757(~n_373_v[`W-1], db5_v, db5_port_4);
  spice_transistor_nmos_gnd t92(~n_381_v[`W-1], ab8_v, ab8_port_1);
  spice_transistor_nmos t3181(~dpc27_SBADH_v[`W-1], adh5_v, sb5_v, adh5_port_5, sb5_port_11);
  spice_transistor_nmos t3180(~dpc39_PCLPCL_v[`W-1], pcl2_v, n_481_v, pcl2_port_1, n_481_port_3);
  spice_transistor_nmos_gnd t3183(~adh5_v[`W-1], n_254_v, n_254_port_1);
  spice_transistor_nmos t3182(~dpc5_SADL_v[`W-1], n_618_v, adl6_v, n_618_port_2, adl6_port_5);
  spice_transistor_nmos_gnd t3188(notidl1_v, idl1_v, idl1_port_1);
  spice_transistor_nmos_vdd t702(abl2_v, n_1152_v, n_1152_port_0);
  spice_transistor_nmos_gnd t700(abl2_v, n_642_v, n_642_port_0);
  spice_transistor_nmos_gnd t709(~idb6_v[`W-1], n_351_v, n_351_port_0);
  spice_transistor_nmos_gnd t708(AxB7_v, n_177_v, n_177_port_0);
  spice_transistor_nmos_vdd t2586(n_1423_v, n_869_v, n_869_port_2);
  spice_transistor_nmos_gnd t2585(n_1423_v, n_1608_v, n_1608_port_2);
  spice_transistor_nmos_gnd t2635(n_1157_v, dpc41_DL_ADL_v, dpc41_DL_ADL_port_9);
  spice_transistor_nmos t1615(~cclk_v[`W-1], n_436_v, x4_v, n_436_port_1, x4_port_1);
  spice_transistor_nmos_gnd t1619(n_1045_v, p7_v, p7_port_1);
  spice_transistor_nmos_vdd t1587(~cclk_v[`W-1], sb0_v, sb0_port_4);
  spice_transistor_nmos t924(~cclk_v[`W-1], n_359_v, _ABH3_v, n_359_port_1, _ABH3_port_1);
  spice_transistor_nmos_vdd t1911(~cclk_v[`W-1], adh2_v, adh2_port_3);
  spice_transistor_nmos_gnd t1919(n_127_v, n_135_v, n_135_port_2);
  spice_transistor_nmos_vdd t1774(n_161_v, dpc0_YSB_v, dpc0_YSB_port_3);
  spice_transistor_nmos t1779(~dpc1_SBY_v[`W-1], y5_v, sb5_v, y5_port_0, sb5_port_5);
  spice_transistor_nmos_gnd g_4888((_AxB_4__C34_v|(~__AxB_4_v[`W-1]&C34_v)), __AxBxC_4_v, __AxBxC_4_port_5);
  spice_transistor_nmos_gnd g_4887(((n_1580_v&n_613_v)|n_1159_v), dasb2_v, dasb2_port_5);
  spice_transistor_nmos t3210(~dpc10_ADLADD_v[`W-1], adl3_v, alub3_v, adl3_port_6, alub3_port_4);
  spice_transistor_nmos t3216(~cclk_v[`W-1], n_1618_v, a2_v, n_1618_port_3, a2_port_2);
  spice_transistor_nmos t1485(~dpc41_DL_ADL_v[`W-1], adl0_v, n_719_v, adl0_port_3, n_719_port_3);
  spice_transistor_nmos t1482(~dpc41_DL_ADL_v[`W-1], adl4_v, n_1095_v, adl4_port_3, n_1095_port_2);
  spice_transistor_nmos t1483(~dpc41_DL_ADL_v[`W-1], adl1_v, n_87_v, adl1_port_2, n_87_port_3);
  spice_transistor_nmos t1481(~dpc41_DL_ADL_v[`W-1], adl3_v, n_1661_v, adl3_port_2, n_1661_port_2);
  spice_transistor_nmos_gnd t2033(pd2_clearIR_v, n_571_v, n_571_port_1);
  spice_transistor_nmos_gnd t2037(notidl4_v, idl4_v, idl4_port_0);
  spice_transistor_nmos t1211(~dpc20_ADDSB06_v[`W-1], alu3_v, sb3_v, alu3_port_1, sb3_port_4);
  spice_transistor_nmos t1210(~dpc20_ADDSB06_v[`W-1], sb4_v, alu4_v, sb4_port_5, alu4_port_2);
  spice_transistor_nmos_vdd t2326(n_1566_v, dpc43_DL_DB_v, dpc43_DL_DB_port_9);
  spice_transistor_nmos_gnd t2490(~dpc29_0ADH17_v[`W-1], adh7_v, adh7_port_4);
  spice_transistor_nmos_gnd t2491(~dpc29_0ADH17_v[`W-1], adh6_v, adh6_port_4);
  spice_transistor_nmos t2320(~dpc37_PCLDB_v[`W-1], n_72_v, idb5_v, n_72_port_1, idb5_port_7);
  spice_transistor_nmos_gnd t1731(pchp3_v, n_141_v, n_141_port_0);
  spice_transistor_nmos_gnd g_4944(((~cclk_v[`W-1]&n_538_v)|~n_807_v[`W-1]), n_330_v, n_330_port_7);
  spice_transistor_nmos_gnd g_4940((n_479_v|(n_739_v&n_61_v)), dasb6_v, dasb6_port_5);
  spice_transistor_nmos_gnd g_4943(((_C23_v&AxB3_v)|__AxB3__C23_v), __AxBxC_3_v, __AxBxC_3_port_5);
  spice_transistor_nmos_vdd t2516(n_1613_v, n_643_v, n_643_port_3);
  spice_transistor_nmos_gnd t791(notalu2_v, alu2_v, alu2_port_1);
  spice_transistor_nmos_gnd t3021(~adl1_v[`W-1], n_1016_v, n_1016_port_1);
  spice_transistor_nmos_vdd t2779(abh1_v, n_1140_v, n_1140_port_1);
  spice_transistor_nmos_vdd t2778(n_842_v, n_66_v, n_66_port_3);
  spice_transistor_nmos_gnd t1792(~n_1501_v[`W-1], db7_v, db7_port_1);
  spice_transistor_nmos g_4711((~cp1_v[`W-1]&fetch_v), n_1083_v, n_1620_v, n_1083_port_7, n_1620_port_3);
  spice_transistor_nmos g_4717((~ADH_ABH_v[`W-1]&~cp1_v[`W-1]), _ABH1_v, n_1267_v, _ABH1_port_3, n_1267_port_3);
  spice_transistor_nmos_gnd t52(n_593_v, dpc4_SSB_v, dpc4_SSB_port_0);
  spice_transistor_nmos t53(~dpc11_SBADD_v[`W-1], alua0_v, sb0_v, alua0_port_0, sb0_port_0);
  spice_transistor_nmos t55(~dpc11_SBADD_v[`W-1], alua5_v, sb5_v, alua5_port_0, sb5_port_0);
  spice_transistor_nmos t56(~dpc11_SBADD_v[`W-1], alua6_v, sb6_v, alua6_port_0, sb6_port_0);
  spice_transistor_nmos_gnd t3235(n_1640_v, n_1251_v, n_1251_port_2);
  spice_transistor_nmos t3233(~cclk_v[`W-1], a4_v, n_1344_v, a4_port_2, n_1344_port_3);
  spice_transistor_nmos_vdd t299(~cclk_v[`W-1], adh0_v, adh0_port_1);
  spice_transistor_nmos_gnd t297(pd7_clearIR_v, n_1605_v, n_1605_port_0);
  spice_transistor_nmos t296(~cp1_v[`W-1], n_719_v, idl0_v, n_719_port_1, idl0_port_0);
  spice_transistor_nmos_gnd t293(n_1413_v, dpc32_PCHADH_v, dpc32_PCHADH_port_0);
  spice_transistor_nmos_vdd t3492(n_6_v, dpc6_SBS_v, dpc6_SBS_port_11);
  spice_transistor_nmos_gnd t3495(~idb1_v[`W-1], n_583_v, n_583_port_1);
  spice_transistor_nmos_vdd t2019(~n_855_v[`W-1], ab0_v, ab0_port_1);
  spice_transistor_nmos t2548(~dpc32_PCHADH_v[`W-1], adh6_v, n_652_v, adh6_port_5, n_652_port_2);
  spice_transistor_nmos t2549(~dpc32_PCHADH_v[`W-1], adh5_v, n_1301_v, adh5_port_4, n_1301_port_2);
  spice_transistor_nmos t2547(~dpc32_PCHADH_v[`W-1], adh7_v, n_1206_v, adh7_port_5, n_1206_port_2);
  spice_transistor_nmos_vdd t2544(n_839_v, n_43_v, n_43_port_11);
  spice_transistor_nmos_gnd t2543(~adl3_v[`W-1], n_1507_v, n_1507_port_1);
  spice_transistor_nmos_vdd t1894(~n_102_v[`W-1], rw_v, rw_port_0);
  spice_transistor_nmos t2733(~cclk_v[`W-1], _ABH2_v, n_994_v, _ABH2_port_2, n_994_port_2);
  spice_transistor_nmos_vdd t2227(n_1499_v, dpc18__DAA_v, dpc18__DAA_port_1);
  spice_transistor_nmos_vdd t196(n_1720_v, n_612_v, n_612_port_0);
  spice_transistor_nmos_vdd t197(dor4_v, n_1076_v, n_1076_port_0);
  spice_transistor_nmos_gnd t190(ir3_v, notir3_v, notir3_port_0);
  spice_transistor_nmos t191(~cclk_v[`W-1], n_1609_v, notir5_v, n_1609_port_0, notir5_port_0);
  spice_transistor_nmos t1958(~dpc13_ORS_v[`W-1], aluanorb0_v, notaluoutmux0_v, aluanorb0_port_1, notaluoutmux0_port_3);
  spice_transistor_nmos_gnd t1959(n_947_v, n_1654_v, n_1654_port_1);
  spice_transistor_nmos_vdd t1956(n_1230_v, dpc11_SBADD_v, dpc11_SBADD_port_9);
  spice_transistor_nmos t1957(~dpc13_ORS_v[`W-1], n_304_v, n_1398_v, n_304_port_3, n_1398_port_1);
  spice_transistor_nmos_gnd g_4341((~RnWstretched_v[`W-1]|dor2_v), n_37_v, n_37_port_4);
  spice_transistor_nmos_vdd t2752(n_21_v, dpc30_ADHPCH_v, dpc30_ADHPCH_port_10);
  spice_transistor_nmos_gnd t2209(n_75_v, dpc20_ADDSB06_v, dpc20_ADDSB06_port_5);
  spice_transistor_nmos_vdd t2208(n_834_v, n_102_v, n_102_port_2);
  spice_transistor_nmos_gnd t2754(notalu7_v, alu7_v, alu7_port_2);
  spice_transistor_nmos_gnd t1408(nots1_v, n_694_v, n_694_port_2);
  spice_transistor_nmos_gnd t1402(ir7_v, notir7_v, notir7_port_33);
  spice_transistor_nmos_gnd g_4773((~alua6_v[`W-1]&~alub6_v[`W-1]), n_336_v, n_336_port_7);
  spice_transistor_nmos t72(~dpc1_SBY_v[`W-1], y6_v, sb6_v, y6_port_1, sb6_port_1);
  spice_transistor_nmos_vdd t76(n_127_v, clk2out_v, clk2out_port_0);
  spice_transistor_nmos t77(~dpc1_SBY_v[`W-1], y4_v, sb4_v, y4_port_0, sb4_port_2);
  spice_transistor_nmos_vdd t75(~dpc14_SRS_v[`W-1], n_304_v, n_304_port_0);
  spice_transistor_nmos_vdd t4(~n_826_v[`W-1], ab8_v, ab8_port_0);
  spice_transistor_nmos_gnd t880(~idb2_v[`W-1], n_458_v, n_458_port_0);
  spice_transistor_nmos_gnd t881(pchp4_v, n_27_v, n_27_port_0);
  spice_transistor_nmos_vdd t1602(~cclk_v[`W-1], idb7_v, idb7_port_3);
  spice_transistor_nmos_gnd g_4908(((n_852_v&n_1205_v)|n_260_v), dasb7_v, dasb7_port_5);
  spice_transistor_nmos_gnd g_4907((~n_330_v[`W-1]|(~cclk_v[`W-1]&n_1599_v)), n_807_v, n_807_port_5);
  spice_transistor_nmos_gnd g_4906(((n_1392_v&~cclk_v[`W-1])|~NMIP_v[`W-1]), n_297_v, n_297_port_5);
  spice_transistor_nmos_vdd t3442(~n_7_v[`W-1], db6_v, db6_port_4);
  spice_transistor_nmos_vdd t3331(~cclk_v[`W-1], idb1_v, idb1_port_10);
  spice_transistor_nmos_gnd t2738(n_1441_v, dpc42_DL_ADH_v, dpc42_DL_ADH_port_8);
  spice_transistor_nmos_gnd t2228(n_1549_v, n_929_v, n_929_port_1);
  spice_transistor_nmos t2731(~cclk_v[`W-1], x5_v, n_578_v, x5_port_2, n_578_port_0);
  spice_transistor_nmos_vdd t2222(~n_1191_v[`W-1], ab6_v, ab6_port_0);
  spice_transistor_nmos_vdd t2221(~cclk_v[`W-1], adl1_v, adl1_port_3);
  spice_transistor_nmos_vdd t2736(~cclk_v[`W-1], adl0_v, adl0_port_6);
  spice_transistor_nmos_gnd t418(~idb5_v[`W-1], n_1383_v, n_1383_port_0);
  spice_transistor_nmos_vdd t416(~cclk_v[`W-1], sb6_v, sb6_port_4);
  spice_transistor_nmos t415(~dpc30_ADHPCH_v[`W-1], pch6_v, adh6_v, pch6_port_0, adh6_port_1);
  spice_transistor_nmos t414(~dpc30_ADHPCH_v[`W-1], pch7_v, adh7_v, pch7_port_1, adh7_port_1);
  spice_transistor_nmos t413(~dpc30_ADHPCH_v[`W-1], pch4_v, adh4_v, pch4_port_1, adh4_port_1);
  spice_transistor_nmos t412(~dpc30_ADHPCH_v[`W-1], pch5_v, adh5_v, pch5_port_0, adh5_port_1);
  spice_transistor_nmos t411(~dpc30_ADHPCH_v[`W-1], pch2_v, adh2_v, pch2_port_0, adh2_port_1);
  spice_transistor_nmos t410(~dpc30_ADHPCH_v[`W-1], pch3_v, adh3_v, pch3_port_1, adh3_port_2);
  spice_transistor_nmos_gnd g_4759((~alub4_v[`W-1]&~alua4_v[`W-1]), n_1063_v, n_1063_port_7);
  spice_transistor_nmos_vdd t15(~n_1140_v[`W-1], ab9_v, ab9_port_0);
  spice_transistor_nmos_vdd t11(n_38_v, n_1247_v, n_1247_port_0);
  spice_transistor_nmos t1859(~dpc25_SBDB_v[`W-1], idb4_v, sb4_v, idb4_port_4, sb4_port_8);
  spice_transistor_nmos t1858(~dpc25_SBDB_v[`W-1], sb3_v, idb3_v, sb3_port_7, idb3_port_3);
  spice_transistor_nmos t1855(~dpc25_SBDB_v[`W-1], sb0_v, idb0_v, sb0_port_6, idb0_port_7);
  spice_transistor_nmos t1857(~dpc25_SBDB_v[`W-1], idb2_v, sb2_v, idb2_port_5, sb2_port_7);
  spice_transistor_nmos t1856(~dpc25_SBDB_v[`W-1], sb1_v, idb1_v, sb1_port_7, idb1_port_4);
  spice_transistor_nmos_gnd t1850(n_251_v, RnWstretched_v, RnWstretched_port_22);
  spice_transistor_nmos t1677(~dpc41_DL_ADL_v[`W-1], adl5_v, n_1387_v, adl5_port_2, n_1387_port_2);
  spice_transistor_nmos_gnd g_4923(((~cclk_v[`W-1]&n_995_v)|~n_854_v[`W-1]), n_975_v, n_975_port_6);
  spice_transistor_nmos_gnd g_4921(((n_432_v&n_345_v)|n_1097_v), dasb3_v, dasb3_port_5);
  spice_transistor_nmos t2503(~dpc8_nDBADD_v[`W-1], alub1_v, n_583_v, alub1_port_0, n_583_port_0);
  spice_transistor_nmos t528(~dpc21_ADDADL_v[`W-1], adl6_v, alu6_v, adl6_port_1, alu6_port_1);
  spice_transistor_nmos t527(~dpc21_ADDADL_v[`W-1], adl5_v, alu5_v, adl5_port_1, alu5_port_0);
  spice_transistor_nmos_gnd t2501(~adh0_v[`W-1], n_1668_v, n_1668_port_0);
  spice_transistor_nmos t526(~dpc21_ADDADL_v[`W-1], alu7_v, adl7_v, alu7_port_0, adl7_port_0);
  spice_transistor_nmos t2504(~dpc8_nDBADD_v[`W-1], alub3_v, n_1621_v, alub3_port_2, n_1621_port_0);
  spice_transistor_nmos t522(~dpc21_ADDADL_v[`W-1], adl4_v, alu4_v, adl4_port_1, alu4_port_1);
  spice_transistor_nmos_vdd t2179(n_1399_v, cp1_v, cp1_port_75);
  spice_transistor_nmos t2241(~dpc26_ACDB_v[`W-1], n_326_v, idb6_v, n_326_port_2, idb6_port_7);
  spice_transistor_nmos t2240(~dpc26_ACDB_v[`W-1], n_831_v, idb5_v, n_831_port_1, idb5_port_5);
  spice_transistor_nmos_vdd t435(n_1523_v, n_635_v, n_635_port_0);
  spice_transistor_nmos_gnd t434(n_1523_v, n_963_v, n_963_port_1);
  spice_transistor_nmos_vdd t437(n_1260_v, dpc32_PCHADH_v, dpc32_PCHADH_port_1);
  spice_transistor_nmos t432(~dpc2_XSB_v[`W-1], n_1169_v, sb0_v, n_1169_port_0, sb0_port_2);
  spice_transistor_nmos_vdd t439(n_220_v, ADL_ABL_v, ADL_ABL_port_0);
  spice_transistor_nmos t2863(~cclk_v[`W-1], n_633_v, n_1059_v, n_633_port_0, n_1059_port_0);
  spice_transistor_nmos t238(~dpc42_DL_ADH_v[`W-1], adh7_v, n_1147_v, adh7_port_0, n_1147_port_0);
  spice_transistor_nmos t237(~dpc42_DL_ADH_v[`W-1], adh6_v, n_1014_v, adh6_port_0, n_1014_port_0);
  spice_transistor_nmos t236(~dpc42_DL_ADH_v[`W-1], adh5_v, n_1387_v, adh5_port_0, n_1387_port_0);
  spice_transistor_nmos t235(~dpc42_DL_ADH_v[`W-1], adh4_v, n_1095_v, adh4_port_0, n_1095_port_0);
  spice_transistor_nmos t234(~dpc42_DL_ADH_v[`W-1], adh3_v, n_1661_v, adh3_port_0, n_1661_port_0);
  spice_transistor_nmos t233(~dpc42_DL_ADH_v[`W-1], adh2_v, n_1424_v, adh2_port_0, n_1424_port_1);
  spice_transistor_nmos t232(~dpc42_DL_ADH_v[`W-1], adh1_v, n_87_v, adh1_port_0, n_87_port_0);
  spice_transistor_nmos t231(~dpc42_DL_ADH_v[`W-1], adh0_v, n_719_v, adh0_port_0, n_719_port_0);
  spice_transistor_nmos_vdd t36(~cclk_v[`W-1], sb4_v, sb4_port_0);
  spice_transistor_nmos t34(~cclk_v[`W-1], n_518_v, y6_v, n_518_port_0, y6_port_0);
  spice_transistor_nmos t2528(~dpc38_PCLADL_v[`W-1], n_1647_v, adl7_v, n_1647_port_1, adl7_port_5);
  spice_transistor_nmos t2529(~dpc38_PCLADL_v[`W-1], adl0_v, n_488_v, adl0_port_5, n_488_port_2);
  spice_transistor_nmos_gnd t3382(n_1271_v, dpc27_SBADH_v, dpc27_SBADH_port_9);
  spice_transistor_nmos_gnd t3439(n_1017_v, n_578_v, n_578_port_2);
  spice_transistor_nmos t3384(~dpc20_ADDSB06_v[`W-1], alu2_v, sb2_v, alu2_port_3, sb2_port_11);
  spice_transistor_nmos_vdd t3434(n_1270_v, dpc39_PCLPCL_v, dpc39_PCLPCL_port_11);
  spice_transistor_nmos_gnd t3388(nots6_v, n_618_v, n_618_port_3);
  spice_transistor_nmos t1876(~dpc41_DL_ADL_v[`W-1], n_1147_v, adl7_v, n_1147_port_2, adl7_port_3);
  spice_transistor_nmos_gnd t1385(n_1356_v, n_326_v, n_326_port_1);
  spice_transistor_nmos t1384(~dpc37_PCLDB_v[`W-1], n_1458_v, idb6_v, n_1458_port_0, idb6_port_3);
  spice_transistor_nmos t592(~dpc43_DL_DB_v[`W-1], idb7_v, n_1147_v, idb7_port_2, n_1147_port_1);
  spice_transistor_nmos t590(~dpc43_DL_DB_v[`W-1], idb5_v, n_1387_v, idb5_port_2, n_1387_port_1);
  spice_transistor_nmos t591(~dpc43_DL_DB_v[`W-1], idb6_v, n_1014_v, idb6_port_0, n_1014_port_1);
  spice_transistor_nmos_vdd t594(~n_322_v[`W-1], ab7_v, ab7_port_0);
  spice_transistor_nmos_gnd t1120(pclp5_v, n_72_v, n_72_port_0);
  spice_transistor_nmos_gnd t1123(n_485_v, n_436_v, n_436_port_0);
  spice_transistor_nmos_gnd t1650(n_987_v, n_1169_v, n_1169_port_1);
  spice_transistor_nmos t82(H1x1_v, p7_v, idb7_v, p7_port_0, idb7_port_0);
  spice_transistor_nmos t2263(~dpc0_YSB_v[`W-1], n_733_v, sb5_v, n_733_port_1, sb5_port_7);
  spice_transistor_nmos t2262(~dpc0_YSB_v[`W-1], n_518_v, sb6_v, n_518_port_2, sb6_port_10);
  spice_transistor_nmos t2260(~dpc0_YSB_v[`W-1], n_658_v, sb4_v, n_658_port_1, sb4_port_10);
  spice_transistor_nmos t450(~dpc9_DBADD_v[`W-1], alub0_v, idb0_v, alub0_port_3, idb0_port_4);
  spice_transistor_nmos_vdd t456(~cclk_v[`W-1], adh1_v, adh1_port_2);
  spice_transistor_nmos t455(~dpc2_XSB_v[`W-1], n_871_v, sb7_v, n_871_port_0, sb7_port_1);
  spice_transistor_nmos_gnd t458(abl3_v, n_138_v, n_138_port_0);
  spice_transistor_nmos_gnd t215(alucout_v, n_206_v, n_206_port_0);
  spice_transistor_nmos_vdd t218(n_241_v, dpc21_ADDADL_v, dpc21_ADDADL_port_0);
  spice_transistor_nmos_gnd t3410(~n_794_v[`W-1], db1_v, db1_port_4);
  spice_transistor_nmos_vdd t1679(~n_42_v[`W-1], db3_v, db3_port_2);
  spice_transistor_nmos_gnd t2040(n_196_v, dpc5_SADL_v, dpc5_SADL_port_7);
  spice_transistor_nmos t2595(~dpc13_ORS_v[`W-1], n_1632_v, n_277_v, n_1632_port_4, n_277_port_5);
  spice_transistor_nmos t1676(~dpc41_DL_ADL_v[`W-1], adl6_v, n_1014_v, adl6_port_2, n_1014_port_2);
  spice_transistor_nmos_gnd t2107(n_1138_v, n_767_v, n_767_port_1);
  spice_transistor_nmos_gnd t2101(~n_171_v[`W-1], ab7_v, ab7_port_1);
  spice_transistor_nmos_gnd t860(~adl7_v[`W-1], n_1046_v, n_1046_port_0);
  spice_transistor_nmos t2108(~cp1_v[`W-1], n_1387_v, idl5_v, n_1387_port_3, idl5_port_0);
  spice_transistor_nmos t1103(~cclk_v[`W-1], n_1724_v, x6_v, n_1724_port_1, x6_port_0);
  spice_transistor_nmos_vdd t1101(~cclk_v[`W-1], adl3_v, adl3_port_1);
  spice_transistor_nmos t1107(~dpc17_SUMS_v[`W-1], __AxBxC_1_v, notaluoutmux1_v, __AxBxC_1_port_1, notaluoutmux1_port_1);
  spice_transistor_nmos t1106(~dpc17_SUMS_v[`W-1], __AxBxC_0_v, notaluoutmux0_v, __AxBxC_0_port_2, notaluoutmux0_port_1);
  spice_transistor_nmos_gnd t1105(n_1238_v, dpc25_SBDB_v, dpc25_SBDB_port_0);
  spice_transistor_nmos t1109(~dpc17_SUMS_v[`W-1], __AxBxC_3_v, n_1071_v, __AxBxC_3_port_1, n_1071_port_3);
  spice_transistor_nmos t1108(~dpc17_SUMS_v[`W-1], __AxBxC_2_v, n_740_v, __AxBxC_2_port_1, n_740_port_2);
  spice_transistor_nmos_gnd g_4517((~RnWstretched_v[`W-1]|n_224_v), n_520_v, n_520_port_4);
  spice_transistor_nmos_gnd g_4515((~cclk_v[`W-1]|n_1518_v|~n_1247_v[`W-1]), dpc39_PCLPCL_v, dpc39_PCLPCL_port_12);
  spice_transistor_nmos_gnd t477(n_1240_v, dpc43_DL_DB_v, dpc43_DL_DB_port_0);
  spice_transistor_nmos_vdd t276(n_631_v, dpc37_PCLDB_v, dpc37_PCLDB_port_0);
  spice_transistor_nmos_vdd t279(~cclk_v[`W-1], adl4_v, adl4_port_0);
  spice_transistor_nmos t2525(~dpc38_PCLADL_v[`W-1], adl4_v, n_208_v, adl4_port_5, n_208_port_2);
  spice_transistor_nmos_gnd t3473(~n_1072_v[`W-1], db0_v, db0_port_4);
  spice_transistor_nmos_gnd t1341(~dpc12_0ADD_v[`W-1], alua7_v, alua7_port_0);
  spice_transistor_nmos t2129(H1x1_v, Pout3_v, idb3_v, Pout3_port_3, idb3_port_5);
  spice_transistor_nmos t2127(H1x1_v, p4_v, idb4_v, p4_port_1, idb4_port_5);
  spice_transistor_nmos t2123(~dpc3_SBX_v[`W-1], x0_v, sb0_v, x0_port_0, sb0_port_7);
  spice_transistor_nmos_vdd t1169(n_519_v, n_135_v, n_135_port_1);
  spice_transistor_nmos_vdd t1699(n_543_v, dpc5_SADL_v, dpc5_SADL_port_0);
  spice_transistor_nmos t1160(~dpc8_nDBADD_v[`W-1], alub0_v, n_624_v, alub0_port_4, n_624_port_1);
  spice_transistor_nmos_gnd g_4533((n_288_v|~RnWstretched_v[`W-1]), n_798_v, n_798_port_4);
  spice_transistor_nmos_gnd g_4455((~cclk_v[`W-1]|~n_1247_v[`W-1]|n_969_v), dpc0_YSB_v, dpc0_YSB_port_12);
  spice_transistor_nmos_gnd g_4452((~n_1247_v[`W-1]|n_763_v|~cclk_v[`W-1]), dpc8_nDBADD_v, dpc8_nDBADD_port_12);
  spice_transistor_nmos_gnd t512(nots4_v, n_3_v, n_3_port_2);
  spice_transistor_nmos_gnd t398(~dpc29_0ADH17_v[`W-1], adh1_v, adh1_port_1);
  spice_transistor_nmos_gnd t393(nots5_v, n_280_v, n_280_port_2);
  spice_transistor_nmos t394(~cclk_v[`W-1], n_1654_v, a3_v, n_1654_port_0, a3_port_0);
  spice_transistor_nmos_vdd t397(n_317_v, n_417_v, n_417_port_1);
  spice_transistor_nmos t2804(~cclk_v[`W-1], n_871_v, x7_v, n_871_port_1, x7_port_2);
  spice_transistor_nmos t2800(~dpc8_nDBADD_v[`W-1], alub7_v, n_423_v, alub7_port_3, n_423_port_0);
  spice_transistor_nmos t1576(~cclk_v[`W-1], y3_v, n_1531_v, y3_port_0, n_1531_port_1);
  spice_transistor_nmos t259(~cclk_v[`W-1], n_242_v, x3_v, n_242_port_0, x3_port_0);
  spice_transistor_nmos t251(~dpc6_SBS_v[`W-1], sb4_v, s4_v, sb4_port_4, s4_port_0);
  spice_transistor_nmos t250(~dpc6_SBS_v[`W-1], s3_v, sb3_v, s3_port_0, sb3_port_2);
  spice_transistor_nmos t253(~dpc6_SBS_v[`W-1], s2_v, sb2_v, s2_port_0, sb2_port_2);
  spice_transistor_nmos t252(~dpc6_SBS_v[`W-1], s1_v, sb1_v, s1_port_0, sb1_port_1);
  spice_transistor_nmos t1523(~dpc3_SBX_v[`W-1], sb4_v, x4_v, sb4_port_6, x4_port_0);
  spice_transistor_nmos_vdd t3458(~n_634_v[`W-1], ab4_v, ab4_port_1);
  spice_transistor_nmos_gnd t3321(notalu3_v, alu3_v, alu3_port_2);
  spice_transistor_nmos_vdd t3323(n_1277_v, dpc42_DL_ADH_v, dpc42_DL_ADH_port_9);
  spice_transistor_nmos_gnd t3450(~n_138_v[`W-1], ab3_v, ab3_port_1);
  spice_transistor_nmos_gnd t1369(notidl0_v, idl0_v, idl0_port_1);
  spice_transistor_nmos_gnd t1365(~idb4_v[`W-1], n_478_v, n_478_port_1);
  spice_transistor_nmos t2242(~dpc26_ACDB_v[`W-1], n_1592_v, idb7_v, n_1592_port_2, idb7_port_7);
  spice_transistor_nmos t538(~dpc13_ORS_v[`W-1], n_740_v, n_1691_v, n_740_port_0, n_1691_port_1);
  spice_transistor_nmos_gnd t534(n_990_v, n_1041_v, n_1041_port_1);
  spice_transistor_nmos_vdd t535(n_990_v, n_138_v, n_138_port_1);
  spice_transistor_nmos_vdd t2148(~cclk_v[`W-1], adh5_v, adh5_port_2);
  spice_transistor_nmos_vdd t2149(~cclk_v[`W-1], adl6_v, adl6_port_3);
  spice_transistor_nmos_gnd t2143(n_108_v, dpc16_EORS_v, dpc16_EORS_port_8);
  spice_transistor_nmos t2146(~cclk_v[`W-1], n_1169_v, x0_v, n_1169_port_2, x0_port_1);
  spice_transistor_nmos_gnd t2145(n_850_v, n_430_v, n_430_port_2);
  spice_transistor_nmos_gnd g_4558((~alua2_v[`W-1]|~alub2_v[`W-1]), n_1691_v, n_1691_port_8);
  spice_transistor_nmos_gnd g_4550((~RnWstretched_v[`W-1]|dor5_v), n_612_v, n_612_port_4);
  spice_transistor_nmos_gnd g_4554((~cclk_v[`W-1]|~n_1247_v[`W-1]|n_800_v), dpc26_ACDB_v, dpc26_ACDB_port_12);
  spice_transistor_nmos_gnd g_4555((~cclk_v[`W-1]|~n_1247_v[`W-1]|n_1335_v), dpc24_ACSB_v, dpc24_ACSB_port_12);
  spice_transistor_nmos_gnd g_4434((~alub7_v[`W-1]|~alua7_v[`W-1]), n_1398_v, n_1398_port_8);
  spice_transistor_nmos_vdd t1515(n_288_v, n_794_v, n_794_port_1);
  spice_transistor_nmos t2799(~dpc8_nDBADD_v[`W-1], alub6_v, n_351_v, alub6_port_3, n_351_port_1);
  spice_transistor_nmos t2798(~dpc8_nDBADD_v[`W-1], alub5_v, n_1383_v, alub5_port_3, n_1383_port_1);
  spice_transistor_nmos_gnd t2797(n_565_v, n_658_v, n_658_port_2);
  spice_transistor_nmos_gnd t3157(pclp6_v, n_1458_v, n_1458_port_2);
  spice_transistor_nmos_gnd t3153(n_130_v, ADL_ABL_v, ADL_ABL_port_5);
  spice_transistor_nmos_gnd t3150(n_1434_v, n_1709_v, n_1709_port_1);
  spice_transistor_nmos_gnd t3151(nots2_v, n_1389_v, n_1389_port_3);
  spice_transistor_nmos_gnd t1554(~n_86_v[`W-1], ab4_v, ab4_port_0);
  spice_transistor_nmos_gnd t2056(~n_676_v[`W-1], ab9_v, ab9_port_1);
  spice_transistor_nmos_gnd t2050(n_1346_v, n_1296_v, n_1296_port_2);
  spice_transistor_nmos_vdd t2051(n_1346_v, n_359_v, n_359_port_2);
  spice_transistor_nmos t2053(~dpc19_ADDSB7_v[`W-1], alu7_v, sb7_v, alu7_port_1, sb7_port_6);
  spice_transistor_nmos_gnd t3309(n_1561_v, n_871_v, n_871_port_2);
  spice_transistor_nmos_gnd t3056(AxB1_v, n_953_v, n_953_port_1);
  spice_transistor_nmos_gnd t518(ir6_v, notir6_v, notir6_port_0);
  spice_transistor_nmos_vdd t517(n_1223_v, dpc9_DBADD_v, dpc9_DBADD_port_1);
  spice_transistor_nmos_gnd g_4572((dor7_v|~RnWstretched_v[`W-1]), n_1501_v, n_1501_port_4);
  spice_transistor_nmos_gnd t1307(~adh2_v[`W-1], n_168_v, n_168_port_0);
  spice_transistor_nmos t1308(~dpc10_ADLADD_v[`W-1], adl2_v, alub2_v, adl2_port_1, alub2_port_1);
  spice_transistor_nmos_gnd t350(~n_66_v[`W-1], ab1_v, ab1_port_0);

  spice_pullup pullup_3283(rdy_v, rdy_port_2);
  spice_pullup pullup_4089(Pout2_v, Pout2_port_2);
  spice_pullup pullup_4084(alu3_v, alu3_port_3);
  spice_pullup pullup_3349(n_208_v, n_208_port_4);
  spice_pullup pullup_3347(n_206_v, n_206_port_5);
  spice_pullup pullup_3350(n_209_v, n_209_port_4);
  spice_pullup pullup_3605(n_624_v, n_624_port_2);
  spice_pullup pullup_3401(n_280_v, n_280_port_4);
  spice_pullup pullup_3361(n_227_v, n_227_port_2);
  spice_pullup pullup_4235(n_1694_v, n_1694_port_3);
  spice_pullup pullup_4234(n_1691_v, n_1691_port_7);
  spice_pullup pullup_3791(n_935_v, n_935_port_2);
  spice_pullup pullup_3420(__AxB_4_v, __AxB_4_port_4);
  spice_pullup pullup_3882(n_1084_v, n_1084_port_5);
  spice_pullup pullup_3881(n_1083_v, n_1083_port_4);
  spice_pullup pullup_3940(notir2_v, notir2_port_20);
  spice_pullup pullup_3487(n_423_v, n_423_port_2);
  spice_pullup pullup_3325(n_168_v, n_168_port_2);
  spice_pullup pullup_3341(notir0_v, notir0_port_28);
  spice_pullup pullup_4119(dasb3_v, dasb3_port_3);
  spice_pullup pullup_4116(n_1469_v, n_1469_port_2);
  spice_pullup pullup_3909(notir3_v, notir3_port_51);
  spice_pullup pullup_3906(p4_v, p4_port_2);
  spice_pullup pullup_3904(idl6_v, idl6_port_2);
  spice_pullup pullup_3481(n_409_v, n_409_port_3);
  spice_pullup pullup_3480(n_404_v, n_404_port_5);
  spice_pullup pullup_4132(n_1496_v, n_1496_port_4);
  spice_pullup pullup_4130(dasb7_v, dasb7_port_3);
  spice_pullup pullup_4139(n_1507_v, n_1507_port_2);
  spice_pullup pullup_3714(n_807_v, n_807_port_3);
  spice_pullup pullup_4151(n_1531_v, n_1531_port_3);
  spice_pullup pullup_4158(n_1548_v, n_1548_port_2);
  spice_pullup pullup_3389(dasb5_v, dasb5_port_3);
  spice_pullup pullup_3380(n_254_v, n_254_port_2);
  spice_pullup pullup_3528(n_488_v, n_488_port_4);
  spice_pullup pullup_3520(n_478_v, n_478_port_2);
  spice_pullup pullup_3523(n_481_v, n_481_port_4);
  spice_pullup pullup_3526(__AxBxC_5_v, __AxBxC_5_port_3);
  spice_pullup pullup_3735(aluanandb1_v, aluanandb1_port_4);
  spice_pullup pullup_3503(dasb2_v, dasb2_port_3);
  spice_pullup pullup_3506(n_458_v, n_458_port_2);
  spice_pullup pullup_3509(idl3_v, idl3_port_2);
  spice_pullup pullup_3754(alu1_v, alu1_port_4);
  spice_pullup pullup_3753(n_871_v, n_871_port_3);
  spice_pullup pullup_3752(idl1_v, idl1_port_2);
  spice_pullup pullup_4194(n_1618_v, n_1618_port_4);
  spice_pullup pullup_4196(n_1621_v, n_1621_port_2);
  spice_pullup pullup_4030(notir7_v, notir7_port_35);
  spice_pullup pullup_3989(n_1251_v, n_1251_port_3);
  spice_pullup pullup_4200(aluanandb0_v, aluanandb0_port_5);
  spice_pullup pullup_4203(n_1632_v, n_1632_port_5);
  spice_pullup pullup_3859(n_1046_v, n_1046_port_2);
  spice_pullup pullup_3548(n_518_v, n_518_port_3);
  spice_pullup pullup_3237(n_3_v, n_3_port_4);
  spice_pullup pullup_4019(idl4_v, idl4_port_2);
  spice_pullup pullup_4015(n_1301_v, n_1301_port_4);
  spice_pullup pullup_4226(so_v, so_port_2);
  spice_pullup pullup_4224(n_1668_v, n_1668_port_2);
  spice_pullup pullup_4075(n_1398_v, n_1398_port_6);
  spice_pullup pullup_4073(notir5_v, notir5_port_37);
  spice_pullup pullup_4070(n_1389_v, n_1389_port_4);
  spice_pullup pullup_3594(alu4_v, alu4_port_3);
  spice_pullup pullup_3663(n_723_v, n_723_port_4);
  spice_pullup pullup_3662(n_721_v, n_721_port_4);
  spice_pullup pullup_4240(n_1709_v, n_1709_port_3);
  spice_pullup pullup_3582(n_583_v, n_583_port_2);
  spice_pullup pullup_3274(n_72_v, n_72_port_4);
  spice_pullup pullup_3277(p6_v, p6_port_2);
  spice_pullup pullup_4055(p7_v, p7_port_2);
  spice_pullup pullup_3870(idl2_v, idl2_port_2);
  spice_pullup pullup_3646(n_694_v, n_694_port_4);
  spice_pullup pullup_3640(Pout0_v, Pout0_port_2);
  spice_pullup pullup_3351(n_212_v, n_212_port_2);
  spice_pullup pullup_3254(n_27_v, n_27_port_4);
  spice_pullup pullup_3253(notir4_v, notir4_port_26);
  spice_pullup pullup_3250(__AxBxC_2_v, __AxBxC_2_port_3);
  spice_pullup pullup_3424(alu5_v, alu5_port_4);
  spice_pullup pullup_3815(n_975_v, n_975_port_3);
  spice_pullup pullup_3816(n_976_v, n_976_port_4);
  spice_pullup pullup_3624(n_658_v, n_658_port_3);
  spice_pullup pullup_3623(n_652_v, n_652_port_4);
  spice_pullup pullup_3622(__AxBxC_4_v, __AxBxC_4_port_3);
  spice_pullup pullup_3621(n_649_v, n_649_port_5);
  spice_pullup pullup_3837(n_1016_v, n_1016_port_2);
  spice_pullup pullup_3835(dasb1_v, dasb1_port_3);
  spice_pullup pullup_3830(n_998_v, n_998_port_4);
  spice_pullup pullup_3602(n_618_v, n_618_port_4);
  spice_pullup pullup_3299(n_123_v, n_123_port_2);
  spice_pullup pullup_3370(idl5_v, idl5_port_2);
  spice_pullup pullup_3372(n_242_v, n_242_port_3);
  spice_pullup pullup_3412(n_297_v, n_297_port_3);
  spice_pullup pullup_3436(alu6_v, alu6_port_4);
  spice_pullup pullup_3437(n_332_v, n_332_port_4);
  spice_pullup pullup_3314(n_146_v, n_146_port_4);
  spice_pullup pullup_3312(aluanorb0_v, aluanorb0_port_6);
  spice_pullup pullup_3310(n_141_v, n_141_port_4);
  spice_pullup pullup_3318(aluanorb1_v, aluanorb1_port_5);
  spice_pullup pullup_3956(n_1206_v, n_1206_port_4);
  spice_pullup pullup_3950(__AxBxC_6_v, __AxBxC_6_port_3);
  spice_pullup pullup_3784(n_928_v, n_928_port_2);
  spice_pullup pullup_3785(n_929_v, n_929_port_4);
  spice_pullup pullup_3431(n_326_v, n_326_port_4);
  spice_pullup pullup_3435(n_330_v, n_330_port_4);
  spice_pullup pullup_3891(n_1094_v, n_1094_port_2);
  spice_pullup pullup_3330(n_177_v, n_177_port_2);
  spice_pullup pullup_3931(n_1169_v, n_1169_port_3);
  spice_pullup pullup_3450(n_351_v, n_351_port_2);
  spice_pullup pullup_3459(__AxBxC_0_v, __AxBxC_0_port_3);
  spice_pullup pullup_4109(__AxB_6_v, __AxB_6_port_6);
  spice_pullup pullup_4108(n_1458_v, n_1458_port_4);
  spice_pullup pullup_4101(Pout1_v, Pout1_port_2);
  spice_pullup pullup_3687(alu7_v, alu7_port_3);
  spice_pullup pullup_3688(n_767_v, n_767_port_3);
  spice_pullup pullup_3473(idl7_v, idl7_port_2);
  spice_pullup pullup_3441(n_336_v, n_336_port_6);
  spice_pullup pullup_3449(n_350_v, n_350_port_4);
  spice_pullup pullup_3494(n_436_v, n_436_port_3);
  spice_pullup pullup_3495(Pout3_v, Pout3_port_4);
  spice_pullup pullup_4144(n_1519_v, n_1519_port_2);
  spice_pullup pullup_4149(__AxB_0_v, __AxB_0_port_4);
  spice_pullup pullup_3397(__AxBxC_3_v, __AxBxC_3_port_3);
  spice_pullup pullup_3533(n_494_v, n_494_port_2);
  spice_pullup pullup_3759(n_880_v, n_880_port_2);
  spice_pullup pullup_3519(n_477_v, n_477_port_4);
  spice_pullup pullup_3510(n_465_v, n_465_port_2);
  spice_pullup pullup_3729(n_831_v, n_831_port_4);
  spice_pullup pullup_4180(n_1592_v, n_1592_port_4);
  spice_pullup pullup_4185(idl0_v, idl0_port_2);
  spice_pullup pullup_4189(n_1605_v, n_1605_port_3);
  spice_pullup pullup_3576(n_571_v, n_571_port_2);
  spice_pullup pullup_3570(n_564_v, n_564_port_3);
  spice_pullup pullup_3579(n_578_v, n_578_port_3);
  spice_pullup pullup_3999(n_1267_v, n_1267_port_2);
  spice_pullup pullup_3746(n_854_v, n_854_port_4);
  spice_pullup pullup_4213(n_1647_v, n_1647_port_4);
  spice_pullup pullup_3555(__AxBxC_7_v, __AxBxC_7_port_3);
  spice_pullup pullup_4028(n_1318_v, n_1318_port_5);
  spice_pullup pullup_4021(n_1309_v, n_1309_port_2);
  spice_pullup pullup_3767(notir6_v, notir6_port_39);
  spice_pullup pullup_3762(n_884_v, n_884_port_2);
  spice_pullup pullup_3761(n_883_v, n_883_port_2);
  spice_pullup pullup_4216(n_1654_v, n_1654_port_4);
  spice_pullup pullup_3848(NMIP_v, NMIP_port_4);
  spice_pullup pullup_4253(n_1724_v, n_1724_port_3);
  spice_pullup pullup_4252(n_1722_v, n_1722_port_4);
  spice_pullup pullup_4066(n_1383_v, n_1383_port_2);
  spice_pullup pullup_4128(n_1491_v, n_1491_port_3);
  spice_pullup pullup_3868(n_1063_v, n_1063_port_5);
  spice_pullup pullup_3670(n_733_v, n_733_port_3);
  spice_pullup pullup_4042(n_1344_v, n_1344_port_4);
  spice_pullup pullup_3801(n_953_v, n_953_port_2);
  spice_pullup pullup_3809(__AxBxC_1_v, __AxBxC_1_port_3);
  spice_pullup pullup_3652(notir1_v, notir1_port_23);
  spice_pullup pullup_3651(__AxB_2_v, __AxB_2_port_4);
  spice_pullup pullup_4206(alu2_v, alu2_port_4);
  spice_pullup pullup_4209(n_1641_v, n_1641_port_2);
  spice_pullup pullup_3636(dasb6_v, dasb6_port_3);
  spice_pullup pullup_3637(n_681_v, n_681_port_6);
  spice_pullup pullup_3478(alu0_v, alu0_port_3);

  spice_latch latch_5130(eclk,ereset, ~cclk_v[`W-1], op_EORS_v, n_982_v);
  spice_latch latch_5131(eclk,ereset, ~cclk_v[`W-1], n_1110_v, pipeUNK01_v);
  spice_latch latch_5132(eclk,ereset, ~cp1_v[`W-1], n_533_v, n_599_v);
  spice_latch latch_5133(eclk,ereset, ~cp1_v[`W-1], n_920_v, n_785_v);
  spice_latch latch_5134(eclk,ereset, ~cclk_v[`W-1], VEC1_v, n_1452_v);
  spice_latch latch_5135(eclk,ereset, ~cclk_v[`W-1], n_896_v, notidl3_v);
  spice_latch latch_5138(eclk,ereset, ~cclk_v[`W-1], n_1187_v, nots6_v);
  spice_latch latch_5109(eclk,ereset, ~cclk_v[`W-1], ~n_722_v[`W-1], notalu6_v);
  spice_latch latch_5107(eclk,ereset, ~cp1_v[`W-1], n_566_v, p1_v);
  spice_latch latch_5106(eclk,ereset, ~cp1_v[`W-1], notRnWprepad_v, n_1579_v);
  spice_latch latch_5045(eclk,ereset, ~cp1_v[`W-1], n_1215_v, n_223_v);
  spice_latch latch_5047(eclk,ereset, ~cp1_v[`W-1], n_931_v, n_1674_v);
  spice_latch latch_4972(eclk,ereset, ~cclk_v[`W-1], n_862_v, pipeUNK11_v);
  spice_latch latch_5088(eclk,ereset, ~cp1_v[`W-1], n_1497_v, n_653_v);
  spice_latch latch_5089(eclk,ereset, ~cclk_v[`W-1], n_616_v, n_460_v);
  spice_latch latch_5084(eclk,ereset, ~cclk_v[`W-1], n_1281_v, pd3_v);
  spice_latch latch_5085(eclk,ereset, ~cclk_v[`W-1], n_1588_v, pd5_v);
  spice_latch latch_5086(eclk,ereset, ~cclk_v[`W-1], n_1075_v, pd4_v);
  spice_latch latch_5087(eclk,ereset, ~cclk_v[`W-1], n_1638_v, notidl6_v);
  spice_latch latch_5080(eclk,ereset, ~cclk_v[`W-1], ~notaluoutmux0_v[`W-1], notalu0_v);
  spice_latch latch_5081(eclk,ereset, ~cclk_v[`W-1], ~n_296_v[`W-1], notalu4_v);
  spice_latch latch_5082(eclk,ereset, ~cclk_v[`W-1], n_340_v, pipeUNK12_v);
  spice_latch latch_5083(eclk,ereset, ~cp1_v[`W-1], notRnWprepad_v, n_759_v);
  spice_latch latch_5136(eclk,ereset, ~cp1_v[`W-1], n_720_v, n_1338_v);
  spice_latch latch_5137(eclk,ereset, ~cclk_v[`W-1], n_1229_v, pchp0_v);
  spice_latch latch_5139(eclk,ereset, ~cp1_v[`W-1], n_1082_v, p0_v);
  spice_latch latch_5054(eclk,ereset, ~cp1_v[`W-1], n_1376_v, notdor2_v);
  spice_latch latch_4959(eclk,ereset, ~cclk_v[`W-1], n_1194_v, pipeUNK04_v);
  spice_latch latch_4958(eclk,ereset, ~cclk_v[`W-1], n_1106_v, n_1404_v);
  spice_latch latch_4955(eclk,ereset, ~cp1_v[`W-1], n_1275_v, n_1581_v);
  spice_latch latch_4954(eclk,ereset, ~cclk_v[`W-1], n_718_v, notidl0_v);
  spice_latch latch_4957(eclk,ereset, ~cclk_v[`W-1], n_1391_v, pipeUNK15_v);
  spice_latch latch_4956(eclk,ereset, ~cp1_v[`W-1], D1x1_v, n_1472_v);
  spice_latch latch_4951(eclk,ereset, ~cclk_v[`W-1], n_548_v, nots7_v);
  spice_latch latch_4950(eclk,ereset, ~cclk_v[`W-1], n_695_v, n_1341_v);
  spice_latch latch_4953(eclk,ereset, ~cclk_v[`W-1], ~n_740_v[`W-1], notalu2_v);
  spice_latch latch_4952(eclk,ereset, ~cclk_v[`W-1], n_795_v, n_360_v);
  spice_latch latch_4977(eclk,ereset, ~cclk_v[`W-1], n_182_v, n_265_v);
  spice_latch latch_4976(eclk,ereset, ~cp1_v[`W-1], ~notRdy0_v[`W-1], n_902_v);
  spice_latch latch_4975(eclk,ereset, ~cp1_v[`W-1], n_789_v, notdor7_v);
  spice_latch latch_4974(eclk,ereset, ~cclk_v[`W-1], n_213_v, notidl1_v);
  spice_latch latch_4971(eclk,ereset, ~cp1_v[`W-1], n_299_v, n_1625_v);
  spice_latch latch_4970(eclk,ereset, ~cp1_v[`W-1], n_1687_v, notdor0_v);
  spice_latch latch_5022(eclk,ereset, ~cp1_v[`W-1], n_845_v, p2_v);
  spice_latch latch_5023(eclk,ereset, ~cclk_v[`W-1], n_318_v, pipeUNK14_v);
  spice_latch latch_5020(eclk,ereset, ~cclk_v[`W-1], notaluvout_v, n_408_v);
  spice_latch latch_5021(eclk,ereset, ~cclk_v[`W-1], n_462_v, n_878_v);
  spice_latch latch_5026(eclk,ereset, ~cclk_v[`W-1], C78_v, C78_phi2_v);
  spice_latch latch_5027(eclk,ereset, ~cclk_v[`W-1], n_1090_v, n_1683_v);
  spice_latch latch_5024(eclk,ereset, ~cclk_v[`W-1], n_188_v, pipeT4out_v);
  spice_latch latch_5025(eclk,ereset, ~cp1_v[`W-1], n_1087_v, n_1132_v);
  spice_latch latch_5028(eclk,ereset, ~cclk_v[`W-1], n_586_v, pipeBRtaken_v);
  spice_latch latch_5029(eclk,ereset, ~cclk_v[`W-1], n_983_v, nots0_v);
  spice_latch latch_5123(eclk,ereset, ~cclk_v[`W-1], n_1175_v, pipeUNK28_v);
  spice_latch latch_5122(eclk,ereset, ~cclk_v[`W-1], n_1085_v, pipeUNK23_v);
  spice_latch latch_5129(eclk,ereset, ~cclk_v[`W-1], n_484_v, pclp7_v);
  spice_latch latch_5128(eclk,ereset, ~cp1_v[`W-1], n_916_v, n_1409_v);
  spice_latch latch_5004(eclk,ereset, ~cclk_v[`W-1], _WR_v, pipe_WR_phi2_v);
  spice_latch latch_5005(eclk,ereset, ~cp1_v[`W-1], n_1375_v, n_95_v);
  spice_latch latch_5006(eclk,ereset, ~cp1_v[`W-1], n_1089_v, n_1529_v);
  spice_latch latch_5007(eclk,ereset, ~cclk_v[`W-1], n_1631_v, pclp3_v);
  spice_latch latch_5000(eclk,ereset, ~cclk_v[`W-1], n_875_v, n_469_v);
  spice_latch latch_5001(eclk,ereset, ~cp1_v[`W-1], n_913_v, n_1274_v);
  spice_latch latch_5002(eclk,ereset, ~cclk_v[`W-1], n_1688_v, n_680_v);
  spice_latch latch_5003(eclk,ereset, ~cclk_v[`W-1], VEC0_v, n_1126_v);
  spice_latch latch_5008(eclk,ereset, ~cp1_v[`W-1], brk_done_v, n_1291_v);
  spice_latch latch_5009(eclk,ereset, ~cp1_v[`W-1], n_428_v, n_644_v);
  spice_latch latch_5068(eclk,ereset, ~cclk_v[`W-1], n_1705_v, n_1020_v);
  spice_latch latch_5069(eclk,ereset, ~cclk_v[`W-1], n_944_v, pipeUNK37_v);
  spice_latch latch_5066(eclk,ereset, ~cp1_v[`W-1], INTG_v, n_50_v);
  spice_latch latch_5067(eclk,ereset, ~cclk_v[`W-1], n_396_v, n_796_v);
  spice_latch latch_5064(eclk,ereset, ~cclk_v[`W-1], op_ORS_v, n_88_v);
  spice_latch latch_5065(eclk,ereset, ~cclk_v[`W-1], n_629_v, n_760_v);
  spice_latch latch_5062(eclk,ereset, ~cclk_v[`W-1], n_515_v, n_1411_v);
  spice_latch latch_5063(eclk,ereset, ~cclk_v[`W-1], n_1211_v, n_897_v);
  spice_latch latch_5060(eclk,ereset, ~cclk_v[`W-1], n_504_v, pipeUNK41_v);
  spice_latch latch_5061(eclk,ereset, ~cclk_v[`W-1], op_ANDS_v, n_1574_v);
  spice_latch latch_5071(eclk,ereset, ~cclk_v[`W-1], n_17_v, pipe_T0_v);
  spice_latch latch_5040(eclk,ereset, ~cclk_v[`W-1], n_62_v, pd7_v);
  spice_latch latch_5041(eclk,ereset, ~cp1_v[`W-1], n_1290_v, n_698_v);
  spice_latch latch_5042(eclk,ereset, ~cclk_v[`W-1], n_374_v, pd6_v);
  spice_latch latch_5043(eclk,ereset, ~cp1_v[`W-1], n_1718_v, n_671_v);
  spice_latch latch_5044(eclk,ereset, ~cp1_v[`W-1], ~notRdy0_v[`W-1], n_1679_v);
  spice_latch latch_5046(eclk,ereset, ~cclk_v[`W-1], n_440_v, pipeUNK39_v);
  spice_latch latch_5048(eclk,ereset, ~cp1_v[`W-1], n_1526_v, n_1450_v);
  spice_latch latch_5049(eclk,ereset, ~cclk_v[`W-1], n_604_v, n_1477_v);
  spice_latch latch_5118(eclk,ereset, ~cclk_v[`W-1], n_80_v, n_1333_v);
  spice_latch latch_4973(eclk,ereset, ~cclk_v[`W-1], n_862_v, pipeT_SYNC_v);
  spice_latch latch_4979(eclk,ereset, ~cclk_v[`W-1], op_T__bit_v, n_1673_v);
  spice_latch latch_4978(eclk,ereset, ~cclk_v[`W-1], n_490_v, notidl4_v);
  spice_latch latch_5141(eclk,ereset, ~cclk_v[`W-1], n_844_v, n_459_v);
  spice_latch latch_5140(eclk,ereset, ~cclk_v[`W-1], n_1486_v, n_126_v);
  spice_latch latch_5143(eclk,ereset, ~cclk_v[`W-1], n_1575_v, pipeT2out_v);
  spice_latch latch_5142(eclk,ereset, ~cclk_v[`W-1], n_474_v, n_15_v);
  spice_latch latch_5145(eclk,ereset, ~cp1_v[`W-1], n_1339_v, n_597_v);
  spice_latch latch_5144(eclk,ereset, ~cclk_v[`W-1], n_973_v, nots4_v);
  spice_latch latch_5149(eclk,ereset, ~cclk_v[`W-1], n_29_v, pipeUNK22_v);
  spice_latch latch_5157(eclk,ereset, ~cp1_v[`W-1], n_1650_v, n_94_v);
  spice_latch latch_4989(eclk,ereset, ~cp1_v[`W-1], n_1178_v, n_590_v);
  spice_latch latch_4980(eclk,ereset, ~cclk_v[`W-1], n_513_v, pipeUNK06_v);
  spice_latch latch_4981(eclk,ereset, ~cp1_v[`W-1], ~n_854_v[`W-1], n_1395_v);
  spice_latch latch_4986(eclk,ereset, ~cclk_v[`W-1], nnT2BR_v, n_1269_v);
  spice_latch latch_4984(eclk,ereset, ~cclk_v[`W-1], n_20_v, n_993_v);
  spice_latch latch_4985(eclk,ereset, ~cclk_v[`W-1], n_1101_v, n_190_v);
  spice_latch latch_5169(eclk,ereset, ~cclk_v[`W-1], n_588_v, notidl7_v);
  spice_latch latch_5168(eclk,ereset, ~cp1_v[`W-1], n_1180_v, n_1533_v);
  spice_latch latch_5163(eclk,ereset, ~cclk_v[`W-1], n_958_v, n_865_v);
  spice_latch latch_5162(eclk,ereset, ~cclk_v[`W-1], n_889_v, pipeUNK42_v);
  spice_latch latch_5161(eclk,ereset, ~cclk_v[`W-1], n_90_v, pipeUNK05_v);
  spice_latch latch_5160(eclk,ereset, ~cp1_v[`W-1], n_472_v, n_1606_v);
  spice_latch latch_5167(eclk,ereset, ~cclk_v[`W-1], n_1455_v, n_1505_v);
  spice_latch latch_5166(eclk,ereset, ~cclk_v[`W-1], n_1037_v, n_266_v);
  spice_latch latch_5165(eclk,ereset, ~cclk_v[`W-1], n_1649_v, n_1027_v);
  spice_latch latch_5164(eclk,ereset, ~cclk_v[`W-1], Reset0_v, pipephi2Reset0_v);
  spice_latch latch_5105(eclk,ereset, ~cclk_v[`W-1], _op_set_C_v, pipeUNK08_v);
  spice_latch latch_5104(eclk,ereset, ~cclk_v[`W-1], n_678_v, pipeT3out_v);
  spice_latch latch_5101(eclk,ereset, ~cclk_v[`W-1], n_1225_v, n_1121_v);
  spice_latch latch_5100(eclk,ereset, ~cclk_v[`W-1], n_1402_v, pchp2_v);
  spice_latch latch_5103(eclk,ereset, ~cclk_v[`W-1], n_1024_v, n_1699_v);
  spice_latch latch_5102(eclk,ereset, ~cclk_v[`W-1], ~n_277_v[`W-1], notalu5_v);
  spice_latch latch_5152(eclk,ereset, ~cclk_v[`W-1], x_op_T__adc_sbc_v, pipeUNK03_v);
  spice_latch latch_5153(eclk,ereset, ~cclk_v[`W-1], DC78_v, DC78_phi2_v);
  spice_latch latch_5150(eclk,ereset, ~cclk_v[`W-1], n_14_v, pipeUNK20_v);
  spice_latch latch_5151(eclk,ereset, ~cclk_v[`W-1], n_696_v, n_610_v);
  spice_latch latch_5154(eclk,ereset, ~cclk_v[`W-1], n_207_v, n_1061_v);
  spice_latch latch_5155(eclk,ereset, ~cclk_v[`W-1], n_31_v, pipeUNK16_v);
  spice_latch latch_5127(eclk,ereset, ~cclk_v[`W-1], n_1319_v, pd1_v);
  spice_latch latch_5126(eclk,ereset, ~cclk_v[`W-1], n_93_v, pd0_v);
  spice_latch latch_5125(eclk,ereset, ~cclk_v[`W-1], op_SRS_v, pipeUNK27_v);
  spice_latch latch_5124(eclk,ereset, ~cclk_v[`W-1], n_160_v, n_1049_v);
  spice_latch latch_5121(eclk,ereset, ~cclk_v[`W-1], n_378_v, pipeT5out_v);
  spice_latch latch_5120(eclk,ereset, ~cp1_v[`W-1], n_1215_v, n_1528_v);
  spice_latch latch_5146(eclk,ereset, ~cp1_v[`W-1], notRnWprepad_v, n_402_v);
  spice_latch latch_5148(eclk,ereset, ~cclk_v[`W-1], n_1717_v, n_1113_v);
  spice_latch latch_5093(eclk,ereset, ~cclk_v[`W-1], n_1069_v, n_1177_v);
  spice_latch latch_5092(eclk,ereset, ~cclk_v[`W-1], n_1045_v, pipeUNK13_v);
  spice_latch latch_5091(eclk,ereset, ~cclk_v[`W-1], n_728_v, pipeVectorA0_v);
  spice_latch latch_5090(eclk,ereset, ~cp1_v[`W-1], n_109_v, n_1161_v);
  spice_latch latch_5097(eclk,ereset, ~cclk_v[`W-1], n_1711_v, nots1_v);
  spice_latch latch_5096(eclk,ereset, ~cclk_v[`W-1], n_1586_v, n_621_v);
  spice_latch latch_5095(eclk,ereset, ~cclk_v[`W-1], n_1225_v, pipedpc28_v);
  spice_latch latch_5094(eclk,ereset, ~cclk_v[`W-1], Reset0_v, pipephi2Reset0x_v);
  spice_latch latch_5099(eclk,ereset, ~cclk_v[`W-1], n_1073_v, pclp5_v);
  spice_latch latch_5098(eclk,ereset, ~cclk_v[`W-1], n_1358_v, n_521_v);
  spice_latch latch_4948(eclk,ereset, ~cp1_v[`W-1], n_645_v, n_562_v);
  spice_latch latch_4949(eclk,ereset, ~cp1_v[`W-1], n_262_v, n_1447_v);
  spice_latch latch_4947(eclk,ereset, ~cclk_v[`W-1], n_11_v, n_55_v);
  spice_latch latch_4960(eclk,ereset, ~cclk_v[`W-1], n_385_v, pipeUNK30_v);
  spice_latch latch_4961(eclk,ereset, ~cclk_v[`W-1], n_442_v, n_509_v);
  spice_latch latch_4962(eclk,ereset, ~cp1_v[`W-1], n_1368_v, n_1149_v);
  spice_latch latch_4963(eclk,ereset, ~cclk_v[`W-1], n_1179_v, n_393_v);
  spice_latch latch_4964(eclk,ereset, ~cp1_v[`W-1], ~n_430_v[`W-1], n_1570_v);
  spice_latch latch_4965(eclk,ereset, ~cclk_v[`W-1], _VEC_v, pipe_VEC_v);
  spice_latch latch_4966(eclk,ereset, ~cclk_v[`W-1], n_261_v, pipeUNK36_v);
  spice_latch latch_4967(eclk,ereset, ~cp1_v[`W-1], n_959_v, n_323_v);
  spice_latch latch_4968(eclk,ereset, ~cclk_v[`W-1], n_176_v, n_598_v);
  spice_latch latch_4969(eclk,ereset, ~cclk_v[`W-1], n_169_v, pipeUNK29_v);
  spice_latch latch_5031(eclk,ereset, ~cp1_v[`W-1], n_1495_v, p3_v);
  spice_latch latch_5030(eclk,ereset, ~cclk_v[`W-1], n_272_v, n_1162_v);
  spice_latch latch_5033(eclk,ereset, ~cclk_v[`W-1], n_1500_v, n_526_v);
  spice_latch latch_5032(eclk,ereset, ~cclk_v[`W-1], n_191_v, pipeUNK40_v);
  spice_latch latch_5035(eclk,ereset, ~cclk_v[`W-1], n_264_v, n_1693_v);
  spice_latch latch_5034(eclk,ereset, ~cclk_v[`W-1], n_264_v, n_799_v);
  spice_latch latch_5037(eclk,ereset, ~cclk_v[`W-1], n_824_v, n_398_v);
  spice_latch latch_5036(eclk,ereset, ~cclk_v[`W-1], n_334_v, pipeUNK17_v);
  spice_latch latch_5039(eclk,ereset, ~cclk_v[`W-1], n_111_v, pd2_v);
  spice_latch latch_5038(eclk,ereset, ~cclk_v[`W-1], n_1065_v, n_1124_v);
  spice_latch latch_5019(eclk,ereset, ~cclk_v[`W-1], n_779_v, n_805_v);
  spice_latch latch_5018(eclk,ereset, ~cp1_v[`W-1], n_1141_v, n_101_v);
  spice_latch latch_5013(eclk,ereset, ~cclk_v[`W-1], n_1374_v, n_1252_v);
  spice_latch latch_5012(eclk,ereset, ~cclk_v[`W-1], n_1347_v, n_1527_v);
  spice_latch latch_5011(eclk,ereset, ~cp1_v[`W-1], n_1380_v, n_666_v);
  spice_latch latch_5010(eclk,ereset, ~cp1_v[`W-1], n_1474_v, notdor1_v);
  spice_latch latch_5017(eclk,ereset, ~cclk_v[`W-1], n_132_v, pipeUNK26_v);
  spice_latch latch_5016(eclk,ereset, ~cclk_v[`W-1], n_1209_v, n_663_v);
  spice_latch latch_5015(eclk,ereset, ~cp1_v[`W-1], n_1181_v, n_69_v);
  spice_latch latch_5014(eclk,ereset, ~cclk_v[`W-1], n_1594_v, n_688_v);
  spice_latch latch_4982(eclk,ereset, ~cp1_v[`W-1], n_468_v, n_18_v);
  spice_latch latch_4983(eclk,ereset, ~cp1_v[`W-1], n_1039_v, n_24_v);
  spice_latch latch_4987(eclk,ereset, ~cclk_v[`W-1], n_327_v, pipeUNK09_v);
  spice_latch latch_5079(eclk,ereset, ~cclk_v[`W-1], ~n_1071_v[`W-1], notalu3_v);
  spice_latch latch_5078(eclk,ereset, ~cclk_v[`W-1], n_473_v, pipeUNK33_v);
  spice_latch latch_5075(eclk,ereset, ~cclk_v[`W-1], n_1199_v, notidl2_v);
  spice_latch latch_5074(eclk,ereset, ~cclk_v[`W-1], n_1081_v, pipeUNK32_v);
  spice_latch latch_5077(eclk,ereset, ~cclk_v[`W-1], n_389_v, pipeUNK31_v);
  spice_latch latch_5076(eclk,ereset, ~cclk_v[`W-1], n_824_v, pipeUNK34_v);
  spice_latch latch_5070(eclk,ereset, ~cp1_v[`W-1], n_1684_v, notdor6_v);
  spice_latch latch_5073(eclk,ereset, ~cclk_v[`W-1], ~notaluoutmux1_v[`W-1], notalu1_v);
  spice_latch latch_5072(eclk,ereset, ~cp1_v[`W-1], _TWOCYCLE_v, _TWOCYCLE_phi1_v);
  spice_latch latch_5108(eclk,ereset, ~cclk_v[`W-1], n_306_v, n_581_v);
  spice_latch latch_5057(eclk,ereset, ~cp1_v[`W-1], n_797_v, notdor4_v);
  spice_latch latch_5056(eclk,ereset, ~cclk_v[`W-1], n_1117_v, pipeVectorA1_v);
  spice_latch latch_5055(eclk,ereset, ~cclk_v[`W-1], n_34_v, nots3_v);
  spice_latch latch_5053(eclk,ereset, ~cclk_v[`W-1], n_952_v, n_1509_v);
  spice_latch latch_5052(eclk,ereset, ~cp1_v[`W-1], n_961_v, notdor5_v);
  spice_latch latch_5051(eclk,ereset, ~cp1_v[`W-1], ~notRdy0_v[`W-1], n_1276_v);
  spice_latch latch_5050(eclk,ereset, ~cclk_v[`W-1], n_501_v, pipeUNK35_v);
  spice_latch latch_5059(eclk,ereset, ~cp1_v[`W-1], n_1091_v, n_1360_v);
  spice_latch latch_5058(eclk,ereset, ~cclk_v[`W-1], n_700_v, n_1565_v);
  spice_latch latch_5156(eclk,ereset, ~cclk_v[`W-1], n_506_v, n_1602_v);
  spice_latch latch_5158(eclk,ereset, ~cp1_v[`W-1], ~notRdy0_v[`W-1], n_1272_v);
  spice_latch latch_5159(eclk,ereset, ~cp1_v[`W-1], n_1093_v, n_226_v);
  spice_latch latch_5147(eclk,ereset, ~cclk_v[`W-1], n_568_v, notidl5_v);
  spice_latch latch_5119(eclk,ereset, ~cclk_v[`W-1], n_1657_v, pchp4_v);
  spice_latch latch_5112(eclk,ereset, ~cp1_v[`W-1], n_626_v, n_756_v);
  spice_latch latch_5113(eclk,ereset, ~cclk_v[`W-1], n_104_v, n_1221_v);
  spice_latch latch_5170(eclk,ereset, ~cp1_v[`W-1], ~notRdy0_v[`W-1], n_1624_v);
  spice_latch latch_5171(eclk,ereset, ~cp1_v[`W-1], ~n_330_v[`W-1], n_675_v);
  spice_latch latch_5172(eclk,ereset, ~cclk_v[`W-1], n_1712_v, pipeVectorA2_v);
  spice_latch latch_5173(eclk,ereset, ~cclk_v[`W-1], n_496_v, nots5_v);
  spice_latch latch_4999(eclk,ereset, ~cclk_v[`W-1], op_SUMS_v, n_415_v);
  spice_latch latch_4998(eclk,ereset, ~cclk_v[`W-1], op_SRS_v, n_968_v);
  spice_latch latch_4991(eclk,ereset, ~cclk_v[`W-1], n_632_v, n_339_v);
  spice_latch latch_4990(eclk,ereset, ~cclk_v[`W-1], n_1192_v, pchp6_v);
  spice_latch latch_4993(eclk,ereset, ~cclk_v[`W-1], n_1379_v, pipeUNK07_v);
  spice_latch latch_4992(eclk,ereset, ~cclk_v[`W-1], n_1190_v, nots2_v);
  spice_latch latch_4995(eclk,ereset, ~cclk_v[`W-1], n_1130_v, n_512_v);
  spice_latch latch_4994(eclk,ereset, ~cclk_v[`W-1], n_1099_v, pclp1_v);
  spice_latch latch_4997(eclk,ereset, ~cclk_v[`W-1], n_774_v, pipeUNK02_v);
  spice_latch latch_4996(eclk,ereset, ~cclk_v[`W-1], n_674_v, n_745_v);
  spice_latch latch_5116(eclk,ereset, ~cclk_v[`W-1], n_19_v, pipeUNK18_v);
  spice_latch latch_5117(eclk,ereset, ~cclk_v[`W-1], ~n_304_v[`W-1], notalu7_v);
  spice_latch latch_5114(eclk,ereset, ~cp1_v[`W-1], n_420_v, n_47_v);
  spice_latch latch_5115(eclk,ereset, ~cclk_v[`W-1], n_1231_v, pipeUNK21_v);
  spice_latch latch_5110(eclk,ereset, ~cclk_v[`W-1], n_608_v, n_559_v);
  spice_latch latch_5111(eclk,ereset, ~cp1_v[`W-1], n_457_v, notdor3_v);

  assign n_318_v = ~(p1_v);
  assign op_T2_jmp_abs_v = ~((ir5_v|irline3_v|ir7_v|ir4_v|_t2_v|~notir2_v[`W-1]|~notir6_v[`W-1]|~notir3_v[`W-1]));
  assign n_937_v = ~(~pcl0_v[`W-1]);
  assign n_936_v = ~(~aluanandb1_v[`W-1]);
  assign op_SRS_v = ~(n_366_v);
  assign n_947_v = ~(~a3_v[`W-1]);
  assign n_946_v = ~((n_844_v&n_616_v));
  assign n_944_v = ~((n_1449_v|n_759_v));
  assign aluvout_v = ~(n_408_v);
  assign n_319_v = ~((DA_C01_v&n_936_v));
  assign op_T0_cmp_v = ~((~clock1_v[`W-1]|~notir0_v[`W-1]|~notir6_v[`W-1]|~notir7_v[`W-1]|ir5_v));
  assign n_19_v = ~((n_770_v|n_1708_v));
  assign n_432_v = ~(~sb3_v[`W-1]);
  assign n_428_v = ~(((pipeT3out_v&~notRdy0_v[`W-1])|(n_16_v&pipeT2out_v)));
  assign op_T3_plp_pla_v = ~((_t3_v|~notir3_v[`W-1]|ir7_v|~notir5_v[`W-1]|ir2_v|irline3_v|ir4_v));
  assign n_1488_v = ~(n_278_v);
  assign n_335_v = ~((_op_store_v|n_347_v));
  assign VEC1_v = ~(n_698_v);
  assign n_824_v = ~((op_T2_brk_v|op_T3_jsr_v));
  assign n_815_v = ~(pipeVectorA2_v);
  assign n_813_v = ~((n_1258_v|n_440_v));
  assign n_818_v = ~((n_265_v|~n_43_v[`W-1]));
  assign op_T5_brk_v = ~((ir4_v|ir7_v|ir3_v|ir2_v|ir5_v|irline3_v|_t5_v|ir6_v));
  assign op_T__adc_sbc_v = ~((clock2_v|~notir5_v[`W-1]|~notir0_v[`W-1]|~notir6_v[`W-1]));
  assign n_819_v = ~((pipephi2Reset0_v|pipeUNK23_v));
  assign n_1594_v = ~((n_779_v&n_604_v));
  assign n_1214_v = ~(pipeUNK11_v);
  assign n_1215_v = ~((brk_done_v|n_238_v|short_circuit_idx_add_v));
  assign n_1224_v = ~(~idb0_v[`W-1]);
  assign n_1213_v = ~((n_609_v|n_453_v));
  assign n_238_v = ~(pipeUNK35_v);
  assign n_1223_v = ~((n_688_v|~n_43_v[`W-1]));
  assign n_232_v = ~(~pcl6_v[`W-1]);
  assign abl5_v = ~(~_ABL5_v[`W-1]);
  assign n_231_v = ~(PD_xxxx10x0_v);
  assign n_979_v = ~(n_905_v);
  assign n_966_v = ~(n_1683_v);
  assign nnT2BR_v = ~(n_636_v);
  assign n_969_v = ~(n_161_v);
  assign n_321_v = ~(n_398_v);
  assign n_320_v = ~(~sb1_v[`W-1]);
  assign n_317_v = ~(n_445_v);
  assign n_973_v = ~(~s4_v[`W-1]);
  assign _t2_v = ~(n_1575_v);
  assign n_980_v = ~(op_T3_jmp_v);
  assign op_T2_ind_v = ~((_t2_v|ir2_v|~notir0_v[`W-1]|ir3_v));
  assign op_T2_abs_access_v = ~((~notir3_v[`W-1]|_t2_v|op_push_pull_v));
  assign n_278_v = ~(~pch6_v[`W-1]);
  assign op_T0_jsr_v = ~((ir3_v|irline3_v|ir6_v|~notir5_v[`W-1]|ir2_v|~clock1_v[`W-1]|ir4_v|ir7_v));
  assign n_272_v = ~((n_646_v|nnT2BR_v|op_T2_abs_access_v|op_T5_rts_v|n_862_v|n_236_v));
  assign n_269_v = ~((n_1038_v|AxB7_v));
  assign n_264_v = ~((n_1312_v|n_1149_v));
  assign n_267_v = ~((n_544_v|n_785_v|n_1175_v));
  assign n_218_v = ~(n_368_v);
  assign n_0_ADL0_v = ~(pipeVectorA0_v);
  assign n_291_v = ~(n_1121_v);
  assign n_288_v = ~((dor1_v|~RnWstretched_v[`W-1]));
  assign n_636_v = ~(op_T2_branch_v);
  assign op_T2_ADL_ADD_v = ~((_t2_v|ir3_v));
  assign n_213_v = ~(~db1_v[`W-1]);
  assign DA_C01_v = ~(((notalucin_v&~aluanandb0_v[`W-1])|~aluanorb0_v[`W-1]));
  assign n_282_v = ~(n_6_v);
  assign op_T4_mem_abs_idx_v = ~((~notir4_v[`W-1]|_t4_v|~notir3_v[`W-1]));
  assign n_453_v = ~(~pch7_v[`W-1]);
  assign x_op_T4_ind_y_v = ~((~notir4_v[`W-1]|ir2_v|_t4_v|~notir0_v[`W-1]|ir3_v));
  assign n_462_v = ~(n_1338_v);
  assign n_457_v = ~(~idb3_v[`W-1]);
  assign n_877_v = ~((n_506_v|n_933_v));
  assign n_1720_v = ~((dor5_v|~RnWstretched_v[`W-1]));
  assign n_875_v = ~(((n_523_v&n_499_v)|n_743_v));
  assign n_876_v = ~(n_867_v);
  assign n_867_v = ~((_DA_ADD2_v|_DA_ADD1_v));
  assign n_626_v = ~(((DBNeg_v&n_1269_v)|(pipeUNK01_v&n_1401_v)));
  assign n_625_v = ~((~n_43_v[`W-1]|n_459_v));
  assign n_221_v = ~(n_1579_v);
  assign n_617_v = ~(abh1_v);
  assign n_628_v = ~((n_55_v|~cclk_v[`W-1]));
  assign n_224_v = ~((~RnWstretched_v[`W-1]|dor2_v));
  assign n_220_v = ~(n_190_v);
  assign op_T2_mem_zp_v = ~((ir4_v|ir3_v|_t2_v|~notir2_v[`W-1]));
  assign n_616_v = ~((op_T__iny_dey_v|op_T0_tay_ldy_not_idx_v|op_T0_ldy_mem_v));
  assign n_620_v = ~((n_307_v|n_1433_v|n_1371_v|n_1293_v));
  assign n_1339_v = ~(n_799_v);
  assign n_556_v = ~(~a4_v[`W-1]);
  assign _AxB_0__C0in_v = ~((n_105_v|~__AxB_0_v[`W-1]));
  assign n_548_v = ~(~s7_v[`W-1]);
  assign op_shift_v = ~((~notir1_v[`W-1]|ir7_v|ir6_v));
  assign n_544_v = ~(op_ror_v);
  assign n_543_v = ~(n_339_v);
  assign n_553_v = ~((n_1662_v|n_781_v));
  assign _C78_v = ~((n_748_v|(C67_v&A_B7_v)));
  assign op_T0_cpx_cpy_inx_iny_v = ~((~notir7_v[`W-1]|~notir6_v[`W-1]|~clock1_v[`W-1]|irline3_v|ir4_v));
  assign n_236_v = ~(n_1708_v);
  assign n_961_v = ~(~idb5_v[`W-1]);
  assign n_962_v = ~(n_1585_v);
  assign n_1427_v = ~((n_236_v|nnT2BR_v));
  assign n_1423_v = ~(abh5_v);
  assign n_1433_v = ~((n_201_v|_op_branch_bit6_v|n_90_v));
  assign n_1343_v = ~((~notRdy0_v[`W-1]|n_152_v));
  assign n_1345_v = ~((dpc36_IPC_v|n_937_v));
  assign n_1347_v = ~((n_782_v|n_862_v|op_T0_shift_a_v|n_550_v|nnT2BR_v|n_979_v));
  assign n_1346_v = ~(abh3_v);
  assign n_1408_v = ~((n_1044_v&(op_T0_adc_sbc_v|op_rol_ror_v)));
  assign n_1413_v = ~(n_1260_v);
  assign n_1412_v = ~(n_1455_v);
  assign op_T0_lda_v = ~((ir6_v|~notir5_v[`W-1]|~notir7_v[`W-1]|~notir0_v[`W-1]|~clock1_v[`W-1]));
  assign n_397_v = ~(op_T0_lda_v);
  assign n_104_v = ~((nnT2BR_v|n_847_v|n_440_v|op_T4_jmp_v|n_275_v));
  assign n_105_v = ~(notalucin_v);
  assign op_T2_ind_x_v = ~((ir3_v|ir2_v|ir4_v|~notir0_v[`W-1]|_t2_v));
  assign n_1416_v = ~(~idb6_v[`W-1]);
  assign pd7_clearIR_v = ~((pd7_v|clearIR_v));
  assign n_981_v = ~(~y5_v[`W-1]);
  assign n_664_v = ~(op_implied_v);
  assign n_662_v = ~(n_625_v);
  assign op_T3_branch_v = ~((~notir4_v[`W-1]|ir2_v|ir3_v|irline3_v|_t3_v));
  assign n_647_v = ~(~n_477_v[`W-1]);
  assign pd5_clearIR_v = ~((clearIR_v|pd5_v));
  assign op_T0_ldy_mem_v = ~((~clock1_v[`W-1]|~notir7_v[`W-1]|~notir2_v[`W-1]|irline3_v|ir6_v|~notir5_v[`W-1]));
  assign n_420_v = ~(n_865_v);
  assign n_424_v = ~(n_198_v);
  assign n_1440_v = ~(~notRdy0_v[`W-1]);
  assign n_913_v = ~(n_1699_v);
  assign n_906_v = ~(n_1333_v);
  assign n_905_v = ~((n_440_v&op_shift_v));
  assign abl3_v = ~(~_ABL3_v[`W-1]);
  assign _t5_v = ~(n_378_v);
  assign op_T3_mem_zp_idx_v = ~((ir3_v|_t3_v|~notir2_v[`W-1]|~notir4_v[`W-1]));
  assign AxB7_v = ~((n_748_v|~n_1398_v[`W-1]));
  assign n_1240_v = ~(n_1566_v);
  assign op_T2_branch_v = ~((irline3_v|ir3_v|ir2_v|~notir4_v[`W-1]|_t2_v));
  assign n_1238_v = ~(n_1295_v);
  assign x_op_T0_bit_v = ~((ir7_v|ir4_v|~clock1_v[`W-1]|~notir2_v[`W-1]|irline3_v|ir6_v|~notir5_v[`W-1]));
  assign op_T0_brk_rti_v = ~((irline3_v|ir5_v|ir3_v|ir7_v|ir4_v|~clock1_v[`W-1]|ir2_v));
  assign _C56_v = ~((n_647_v|(A_B5_v&C45_v)));
  assign op_T__iny_dey_v = ~((ir4_v|~notir7_v[`W-1]|irline3_v|~notir3_v[`W-1]|ir5_v|clock2_v|ir2_v));
  assign n_154_v = ~(n_512_v);
  assign n_152_v = ~((n_630_v|op_T2_v|n_1002_v|n_952_v));
  assign DC78_v = ~((((n_269_v|n_570_v)&(~__AxB_6_v[`W-1]|n_757_v))|~dpc18__DAA_v[`W-1]));
  assign n_334_v = ~((brk_done_v|p2_v));
  assign op_T__cmp_v = ~((ir5_v|~notir6_v[`W-1]|clock2_v|~notir7_v[`W-1]|~notir0_v[`W-1]));
  assign op_T0_bit_v = ~((ir6_v|irline3_v|~clock1_v[`W-1]|~notir5_v[`W-1]|ir4_v|~notir2_v[`W-1]|ir7_v));
  assign n_299_v = ~(((pipeUNK05_v&n_1614_v)|(n_1416_v&n_1111_v)|n_587_v|(n_1245_v&pipeUNK03_v)));
  assign n_300_v = ~((op_T2_jsr_v|brk_done_v|n_389_v|op_rti_rts_v|x_op_T3_ind_y_v|op_T4_ind_x_v));
  assign n_149_v = ~(~alu6_v[`W-1]);
  assign n_368_v = ~((op_T5_rti_rts_v|xx_op_T5_jsr_v|x_op_T3_plp_pla_v|op_T4_jmp_v|op_T2_jmp_abs_v|op_T2_php_pha_v));
  assign n_1595_v = ~(n_754_v);
  assign n_519_v = ~(~clk0_v[`W-1]);
  assign n_5_v = ~(~a0_v[`W-1]);
  assign op_T0_tay_v = ~((~notir3_v[`W-1]|~clock1_v[`W-1]|~notir7_v[`W-1]|irline3_v|ir2_v|ir6_v|~notir5_v[`W-1]|ir4_v));
  assign H1x1_v = ~(pipeUNK15_v);
  assign n_515_v = ~(((n_783_v&n_1542_v)|n_1253_v));
  assign n_513_v = ~((n_885_v|op_T__bit_v|n_954_v));
  assign op_store_v = ~((~notir7_v[`W-1]|ir5_v|ir6_v));
  assign DA_AxB2_v = ~((DA_AB2_v|~n_1691_v[`W-1]));
  assign n_510_v = ~((op_rmw_v|n_347_v|x_op_jmp_v));
  assign n_507_v = ~(n_1049_v);
  assign n_846_v = ~(_op_branch_bit6_v);
  assign n_845_v = ~(((n_1573_v&n_781_v)|(pipeUNK17_v&n_553_v)|(n_270_v&n_1662_v)));
  assign n_839_v = ~(~cp1_v[`W-1]);
  assign n_838_v = ~(n_581_v);
  assign n_837_v = ~(op_T0_eor_v);
  assign n_834_v = ~(n_402_v);
  assign n_844_v = ~((op_T__inx_v|op_T__dex_v|op_T0_ldx_tax_tsx_v));
  assign n_842_v = ~(abl1_v);
  assign n_1588_v = ~(~db5_v[`W-1]);
  assign n_1586_v = ~(op_T0_tsx_v);
  assign op_ANDS_v = ~(n_669_v);
  assign n_249_v = ~(~pcl3_v[`W-1]);
  assign n_241_v = ~(n_745_v);
  assign n_243_v = ~(~idb1_v[`W-1]);
  assign A_B5_v = ~(~n_1632_v[`W-1]);
  assign _op_set_C_v = ~(((op_asl_rol_v&n_1258_v)|(op_T__cmp_v|op_T__asl_rol_a_v|op_T__cpx_cpy_abs_v|x_op_T__adc_sbc_v|op_T__cpx_cpy_imm_zp_v)));
  assign op_T0_txs_v = ~((~clock1_v[`W-1]|~notir3_v[`W-1]|ir2_v|ir5_v|~notir7_v[`W-1]|ir6_v|~notir1_v[`W-1]|~notir4_v[`W-1]));
  assign op_ror_v = ~((~notir5_v[`W-1]|~notir1_v[`W-1]|ir7_v|~notir6_v[`W-1]));
  assign n_251_v = ~((_DBE_v|n_221_v));
  assign op_T4_rti_v = ~((ir5_v|ir7_v|~notir6_v[`W-1]|ir4_v|irline3_v|_t4_v|ir2_v|ir3_v));
  assign n_1225_v = ~((op_T2_ind_v|op_T2_zp_zp_idx_v));
  assign n_1231_v = ~(n_1409_v);
  assign op_T3_stack_bit_jmp_v = ~((irline3_v|_t3_v|ir7_v|ir4_v));
  assign PD_xxxx10x0_v = ~((~n_1083_v[`W-1]|pd0_clearIR_v|pd2_clearIR_v));
  assign n_1026_v = ~(n_567_v);
  assign n_1028_v = ~(n_251_v);
  assign op_branch_done_v = ~((ir3_v|n_603_v|irline3_v|~notir4_v[`W-1]|~clock1_v[`W-1]|ir2_v));
  assign n_1025_v = ~(~y0_v[`W-1]);
  assign op_T3_ind_y_v = ~((ir2_v|~notir4_v[`W-1]|~notir0_v[`W-1]|ir3_v|_t3_v));
  assign op_T3_mem_abs_v = ~((ir4_v|~notir3_v[`W-1]|_t3_v|~notir2_v[`W-1]));
  assign n_608_v = ~(n_1272_v);
  assign VEC0_v = ~((~notRdy0_v[`W-1]|n_689_v));
  assign pclp2_v = ~(n_1411_v);
  assign op_T0_shift_right_a_v = ~((ir2_v|~notir6_v[`W-1]|ir4_v|~notir1_v[`W-1]|~clock1_v[`W-1]|~notir3_v[`W-1]|ir7_v));
  assign n_1371_v = ~((n_201_v|n_846_v|n_1045_v));
  assign DC34_v = ~((~dpc18__DAA_v[`W-1]|((n_319_v|~n_1691_v[`W-1])&(n_1610_v|n_388_v))));
  assign n_1070_v = ~(~pch1_v[`W-1]);
  assign n_1069_v = ~((n_1274_v|n_1024_v));
  assign n_1075_v = ~(~db4_v[`W-1]);
  assign n_1067_v = ~(n_582_v);
  assign n_1073_v = ~((n_344_v&(n_392_v|n_410_v)));
  assign clearIR_v = ~((fetch_v&D1x1_v));
  assign op_T0_v = ~(~clock1_v[`W-1]);
  assign n_1271_v = ~(n_1596_v);
  assign n_1657_v = ~(((dpc35_PCHC_v|n_83_v)&n_523_v));
  assign op_T0_cpx_inx_v = ~((ir4_v|~notir5_v[`W-1]|~notir6_v[`W-1]|irline3_v|~clock1_v[`W-1]|~notir7_v[`W-1]));
  assign n_1655_v = ~(n_1211_v);
  assign n_1705_v = ~((n_467_v|n_630_v));
  assign n_1708_v = ~(op_T3_branch_v);
  assign n_1688_v = ~(n_1304_v);
  assign n_1270_v = ~((n_509_v|~n_43_v[`W-1]));
  assign _DBZ_v = ~(DBZ_v);
  assign abl2_v = ~(~_ABL2_v[`W-1]);
  assign op_T0_and_v = ~((~notir5_v[`W-1]|~notir0_v[`W-1]|ir6_v|~clock1_v[`W-1]|ir7_v));
  assign n_1497_v = ~(pipeUNK41_v);
  assign n_1495_v = ~(((n_781_v&n_1600_v)|(n_1492_v&n_270_v)|(n_1457_v&pipeUNK04_v)));
  assign _C01_v = ~(C01_v);
  assign n_440_v = ~(n_24_v);
  assign n_1499_v = ~(n_1450_v);
  assign n_1500_v = ~(((dpc36_IPC_v&n_937_v)|n_1345_v));
  assign op_T4_brk_jsr_v = ~((ir4_v|irline3_v|ir6_v|ir2_v|_t4_v|ir3_v|ir7_v));
  assign n_803_v = ~(~n_1084_v[`W-1]);
  assign n_931_v = ~(n_415_v);
  assign n_327_v = ~((op_T0_plp_v|x_op_T4_rti_v));
  assign DBNeg_v = ~(~idb7_v[`W-1]);
  assign n_933_v = ~((n_572_v&n_1262_v));
  assign n_923_v = ~(~pch3_v[`W-1]);
  assign C1x5Reset_v = ~(n_717_v);
  assign n_674_v = ~(n_25_v);
  assign n_673_v = ~((~Pout3_v[`W-1]&op_T0_adc_sbc_v));
  assign n_678_v = ~((n_1357_v|n_644_v));
  assign n_670_v = ~(n_519_v);
  assign n_669_v = ~((op_T0_and_v|op_T0_bit_v));
  assign n_1697_v = ~(n_664_v);
  assign n_992_v = ~(n_595_v);
  assign n_1684_v = ~(~idb6_v[`W-1]);
  assign n_1687_v = ~(~idb0_v[`W-1]);
  assign Reset0_v = ~(n_1395_v);
  assign _AxB_4__C34_v = ~((~__AxB_4_v[`W-1]|C34_v));
  assign op_T0_dex_v = ~((~notir1_v[`W-1]|~clock1_v[`W-1]|~notir6_v[`W-1]|ir2_v|~notir7_v[`W-1]|ir4_v|~notir3_v[`W-1]|ir5_v));
  assign n_75_v = ~(n_154_v);
  assign n_588_v = ~(~db7_v[`W-1]);
  assign n_587_v = ~(pipeUNK12_v);
  assign n_593_v = ~(n_355_v);
  assign _C67_v = ~(C67_v);
  assign n_582_v = ~(n_610_v);
  assign op_T3_jsr_v = ~((ir2_v|irline3_v|~notir5_v[`W-1]|ir6_v|ir4_v|ir3_v|ir7_v|_t3_v));
  assign n_6_v = ~((n_521_v|~n_43_v[`W-1]));
  assign n_8_v = ~(n_551_v);
  assign n_748_v = ~(~n_1318_v[`W-1]);
  assign n_747_v = ~(n_670_v);
  assign n_20_v = ~(((n_344_v&n_232_v)|n_1316_v));
  assign n_21_v = ~((n_1162_v|~n_43_v[`W-1]));
  assign n_739_v = ~(((n_761_v&n_1257_v)|(n_1056_v&n_811_v)));
  assign DBZ_v = ~((~idb4_v[`W-1]|~idb6_v[`W-1]|~idb1_v[`W-1]|~idb5_v[`W-1]|~idb0_v[`W-1]|~idb2_v[`W-1]|~idb7_v[`W-1]|~idb3_v[`W-1]));
  assign n_260_v = ~((n_852_v|n_1205_v));
  assign n_261_v = ~((x_op_T4_ind_y_v|x_op_T3_abs_idx_v));
  assign BRtaken_v = ~(((n_270_v&n_620_v)|n_1115_v));
  assign n_1526_v = ~(n_680_v);
  assign n_1534_v = ~((n_805_v|~n_43_v[`W-1]));
  assign op_from_x_v = ~((~notir7_v[`W-1]|ir6_v|~notir1_v[`W-1]|ir5_v));
  assign n_1549_v = ~(~a1_v[`W-1]);
  assign n_262_v = ~(((pipeUNK29_v&n_1714_v)|(n_1511_v&pipeUNK28_v)));
  assign op_T2_idx_x_xy_v = ~((~notir2_v[`W-1]|~notir4_v[`W-1]|_t2_v));
  assign op_jsr_v = ~((ir4_v|ir2_v|ir7_v|ir6_v|~notir5_v[`W-1]|irline3_v|ir3_v));
  assign n_717_v = ~((pipephi2Reset0x_v|n_1132_v));
  assign n_715_v = ~(n_641_v);
  assign op_T2_jsr_v = ~((ir7_v|ir3_v|_t2_v|~notir5_v[`W-1]|irline3_v|ir6_v|ir4_v|ir2_v));
  assign n_709_v = ~(n_1499_v);
  assign _C34_v = ~(((A_B3_v&C23_v)|(n_988_v|DC34_v)));
  assign n_1434_v = ~(~x1_v[`W-1]);
  assign abh0_v = ~(~_ABH0_v[`W-1]);
  assign x_op_T3_plp_pla_v = ~((ir7_v|ir2_v|~notir3_v[`W-1]|~notir5_v[`W-1]|_t3_v|irline3_v|ir4_v));
  assign n_1640_v = ~(~y7_v[`W-1]);
  assign op_T3_ind_x_v = ~((ir4_v|~notir0_v[`W-1]|ir3_v|_t3_v|ir2_v));
  assign dor0_v = ~(notdor0_v);
  assign n_83_v = ~(n_1400_v);
  assign op_T0_cpy_iny_v = ~((~notir6_v[`W-1]|ir4_v|ir5_v|irline3_v|~clock1_v[`W-1]|~notir7_v[`W-1]));
  assign n_728_v = ~(VEC0_v);
  assign n_730_v = ~(~x6_v[`W-1]);
  assign dpc22__DSA_v = ~(n_599_v);
  assign n_726_v = ~((op_T5_rts_v|x_op_T4_ind_y_v|op_T3_abs_idx_ind_v|op_T5_ind_x_v));
  assign pclp6_v = ~(n_993_v);
  assign n_732_v = ~(((n_1528_v&_TWOCYCLE_phi1_v)|n_1161_v));
  assign n_718_v = ~(~db0_v[`W-1]);
  assign n_720_v = ~((pipeUNK34_v|~notRdy0_v[`W-1]));
  assign n_1719_v = ~(~a5_v[`W-1]);
  assign n_1718_v = ~(~notRdy0_v[`W-1]);
  assign n_1380_v = ~((n_1154_v|n_819_v));
  assign n_1379_v = ~(x_op_T0_bit_v);
  assign n_1377_v = ~(op_rti_rts_v);
  assign n_1376_v = ~(~idb2_v[`W-1]);
  assign n_1464_v = ~((op_T5_rti_v|op_T0_php_pha_v|op_T4_rts_v|op_T3_plp_pla_v|op_T5_brk_v|op_T0_jsr_v));
  assign n_385_v = ~((n_1377_v|n_604_v));
  assign n_1386_v = ~((n_715_v&n_1316_v));
  assign op_T5_mem_ind_idx_v = ~((~notir0_v[`W-1]|_t5_v|ir2_v|ir3_v));
  assign n_1055_v = ~((n_771_v|n_1708_v));
  assign n_1065_v = ~(op_T0_cli_sei_v);
  assign n_384_v = ~((n_1412_v|op_ANDS_v|n_1258_v|n_946_v));
  assign n_383_v = ~(op_T2_jsr_v);
  assign op_T0_iny_dey_v = ~((~notir7_v[`W-1]|ir2_v|~clock1_v[`W-1]|ir4_v|ir5_v|irline3_v|~notir3_v[`W-1]));
  assign dpc36_IPC_v = ~((n_1472_v&(n_1570_v|n_1581_v)));
  assign n_378_v = ~((n_18_v|n_1357_v));
  assign abl1_v = ~(~_ABL1_v[`W-1]);
  assign n_374_v = ~(~db6_v[`W-1]);
  assign n_372_v = ~(~notRdy0_v[`W-1]);
  assign n_631_v = ~(n_878_v);
  assign n_386_v = ~(~pcl5_v[`W-1]);
  assign notaluvout_v = ~(((~n_1398_v[`W-1]&C67_v)|n_637_v));
  assign n_533_v = ~(pipeUNK22_v);
  assign n_1319_v = ~(~db1_v[`W-1]);
  assign n_531_v = ~(n_95_v);
  assign pchp7_v = ~(n_663_v);
  assign xx_op_T5_jsr_v = ~((~notir5_v[`W-1]|ir7_v|_t5_v|ir6_v|ir2_v|ir3_v|irline3_v|ir4_v));
  assign n_525_v = ~((n_266_v|~cclk_v[`W-1]));
  assign n_1312_v = ~((n_1693_v|n_1291_v));
  assign A_B3_v = ~(~n_649_v[`W-1]);
  assign n_270_v = ~(n_503_v);
  assign n_46_v = ~((~notRdy0_v[`W-1]|n_992_v));
  assign op_lsr_ror_dec_inc_v = ~((~notir6_v[`W-1]|~notir1_v[`W-1]));
  assign n_1391_v = ~((op_T2_php_v|op_T4_brk_v));
  assign n_1392_v = ~(~nmi_v[`W-1]);
  assign op_T0_shift_a_v = ~((ir4_v|~clock1_v[`W-1]|~notir3_v[`W-1]|ir7_v|ir2_v|~notir1_v[`W-1]));
  assign n_1399_v = ~(n_1715_v);
  assign op_T3_abs_idx_v = ~((~notir3_v[`W-1]|~notir4_v[`W-1]|_t3_v));
  assign n_61_v = ~(~sb6_v[`W-1]);
  assign n_1401_v = ~(n_1269_v);
  assign n_1402_v = ~(((n_200_v|n_1202_v)&n_293_v));
  assign n_771_v = ~(n_1110_v);
  assign n_779_v = ~((n_1440_v&(op_T0_sbc_v|n_1002_v|n_1081_v)));
  assign n_781_v = ~((~notRdy0_v[`W-1]|pipeUNK09_v));
  assign _C12_v = ~((n_936_v|(C01_v&A_B1_v)));
  assign abh5_v = ~(~_ABH5_v[`W-1]);
  assign n_772_v = ~(n_1674_v);
  assign n_773_v = ~((op_T2_abs_access_v|n_646_v));
  assign n_770_v = ~(n_559_v);
  assign n_1120_v = ~(~notRdy0_v[`W-1]);
  assign n_1117_v = ~(n_70_v);
  assign alucout_v = ~(notalucout_v);
  assign n_1145_v = ~((op_T0_ora_v|~notRdy0_v[`W-1]));
  assign op_T2_stack_access_v = ~((_t2_v|ir4_v|irline3_v|ir7_v|ir2_v));
  assign n_163_v = ~(n_249_v);
  assign n_161_v = ~((~cclk_v[`W-1]|n_1113_v));
  assign op_T0_tax_v = ~((~notir5_v[`W-1]|~notir1_v[`W-1]|ir4_v|~notir7_v[`W-1]|ir2_v|~notir3_v[`W-1]|ir6_v|~clock1_v[`W-1]));
  assign op_clv_v = ~((~notir7_v[`W-1]|ir6_v|irline3_v|~notir4_v[`W-1]|~notir3_v[`W-1]|ir2_v|~notir5_v[`W-1]));
  assign n_1159_v = ~((n_613_v|n_1580_v));
  assign n_1157_v = ~(n_291_v);
  assign x_op_T__adc_sbc_v = ~((~notir5_v[`W-1]|~notir6_v[`W-1]|clock2_v|~notir0_v[`W-1]));
  assign n_91_v = ~(n_1529_v);
  assign D1x1_v = ~((INTG_v|C1x5Reset_v));
  assign n_358_v = ~(~clk0_v[`W-1]);
  assign n_1175_v = ~(n_1447_v);
  assign _op_branch_bit7_v = ~(ir7_v);
  assign n_1179_v = ~((dpc22__DSA_v|C34_v));
  assign n_1178_v = ~((pipeUNK33_v|pipeUNK30_v|pipeUNK31_v|pipeUNK32_v));
  assign n_1181_v = ~(((DBNeg_v&n_754_v)|(n_1595_v&pipeUNK13_v)));
  assign n_1180_v = ~((~notRdy0_v[`W-1]|pipe_T0_v));
  assign x_op_T0_tya_v = ~((irline3_v|~notir3_v[`W-1]|ir6_v|~notir7_v[`W-1]|ir2_v|~notir4_v[`W-1]|~clock1_v[`W-1]|ir5_v));
  assign n_1170_v = ~((n_781_v|n_755_v));
  assign n_1599_v = ~(~irq_v[`W-1]);
  assign n_1596_v = ~(n_1602_v);
  assign n_1593_v = ~(n_226_v);
  assign n_1600_v = ~(~idb3_v[`W-1]);
  assign n_570_v = ~((AxB5_v|DA_C45_v|n_122_v|n_647_v));
  assign n_568_v = ~(~db5_v[`W-1]);
  assign op_sty_cpy_mem_v = ~((ir5_v|~notir7_v[`W-1]|ir6_v|irline3_v|~notir2_v[`W-1]));
  assign n_572_v = ~(pipeUNK21_v);
  assign n_567_v = ~(~_ABL7_v[`W-1]);
  assign n_566_v = ~(((n_1170_v&pipeUNK14_v)|(n_755_v&_DBZ_v)|(n_243_v&n_781_v)));
  assign n_1187_v = ~(~s6_v[`W-1]);
  assign short_circuit_idx_add_v = ~((n_916_v|n_1137_v|pipeUNK36_v|~notRdy0_v[`W-1]));
  assign n_0_ADL2_v = ~(n_815_v);
  assign n_1184_v = ~((n_163_v&n_1253_v));
  assign n_1190_v = ~(~s2_v[`W-1]);
  assign n_1194_v = ~(p3_v);
  assign n_1195_v = ~(abl6_v);
  assign n_1192_v = ~(((n_743_v|n_1488_v)&n_609_v));
  assign n_345_v = ~(((n_8_v&n_876_v)|(n_986_v&n_600_v)));
  assign op_SUMS_v = ~((op_ANDS_v|op_EORS_v|op_SRS_v|op_ORS_v));
  assign n_1293_v = ~((_op_branch_bit7_v|_op_branch_bit6_v|n_318_v));
  assign n_306_v = ~(dpc22__DSA_v);
  assign n_1295_v = ~(n_1527_v);
  assign n_1304_v = ~((n_673_v|op_T0_sbc_v));
  assign op_T5_rts_v = ~((ir3_v|ir2_v|ir7_v|~notir6_v[`W-1]|~notir5_v[`W-1]|ir4_v|irline3_v|_t5_v));
  assign n_1305_v = ~(n_772_v);
  assign n_1290_v = ~(((VEC1_v&~notRdy0_v[`W-1])|n_1126_v));
  assign PD_1xx000x0_v = ~((pd4_clearIR_v|pd3_clearIR_v|~n_1605_v[`W-1]|pd2_clearIR_v|pd0_clearIR_v));
  assign n_1303_v = ~(((op_from_x_v&n_335_v)|(op_sty_cpy_mem_v&n_335_v)));
  assign op_T0_cli_sei_v = ~((~notir4_v[`W-1]|ir7_v|ir2_v|~notir3_v[`W-1]|~notir6_v[`W-1]|~clock1_v[`W-1]|irline3_v));
  assign dor5_v = ~(notdor5_v);
  assign n_1449_v = ~(n_958_v);
  assign n_755_v = ~(pipeUNK06_v);
  assign n_754_v = ~(((pipeUNK09_v&pipeUNK06_v)|n_1673_v));
  assign n_761_v = ~(~alu5_v[`W-1]);
  assign n_757_v = ~((DA_C45_v&n_647_v));
  assign n_763_v = ~(n_1534_v);
  assign n_762_v = ~((n_149_v|n_761_v));
  assign op_jmp_v = ~((irline3_v|~notir3_v[`W-1]|ir7_v|ir4_v|~notir6_v[`W-1]|~notir2_v[`W-1]));
  assign n_769_v = ~((dor0_v|~RnWstretched_v[`W-1]));
  assign n_609_v = ~((n_743_v&n_1488_v));
  assign n_849_v = ~(n_321_v);
  assign n_850_v = ~(pipeUNK18_v);
  assign n_1260_v = ~(n_598_v);
  assign n_1265_v = ~(~pch2_v[`W-1]);
  assign __AxB3__C23_v = ~((_C23_v|AxB3_v));
  assign n_861_v = ~(n_1452_v);
  assign n_852_v = ~(~sb7_v[`W-1]);
  assign n_853_v = ~(n_770_v);
  assign op_rti_rts_v = ~((ir2_v|irline3_v|ir7_v|~notir6_v[`W-1]|ir4_v|ir3_v));
  assign n_847_v = ~(n_300_v);
  assign op_T2_pha_v = ~((ir2_v|ir4_v|ir5_v|~notir3_v[`W-1]|irline3_v|~notir6_v[`W-1]|ir7_v|_t2_v));
  assign n_1087_v = ~((brk_done_v|n_717_v));
  assign dor4_v = ~(notdor4_v);
  assign n_1089_v = ~(n_1574_v);
  assign n_1090_v = ~((n_1222_v|op_T2_stack_access_v));
  assign n_1091_v = ~(((~notRdy0_v[`W-1]&pipeT2out_v)|(n_16_v&pipeT_SYNC_v)));
  assign n_311_v = ~(n_1010_v);
  assign n_312_v = ~(~res_v[`W-1]);
  assign n_1082_v = ~(((pipeUNK16_v&n_279_v)|(n_253_v&n_270_v)|(n_954_v&~n_206_v[`W-1])|(n_507_v&n_1224_v)));
  assign n_1085_v = ~(((n_862_v&~notRdy0_v[`W-1])|(((nnT2BR_v&BRtaken_v)|n_646_v)&n_372_v)));
  assign n_389_v = ~(n_1107_v);
  assign n_1492_v = ~(pipeUNK02_v);
  assign n_390_v = ~(n_653_v);
  assign n_388_v = ~((DA_AxB2_v|n_936_v|AxB1_v|DA_C01_v));
  assign n_392_v = ~(n_386_v);
  assign n_396_v = ~(n_1358_v);
  assign op_T0_txa_v = ~((ir4_v|~notir3_v[`W-1]|~notir1_v[`W-1]|ir6_v|~notir7_v[`W-1]|ir2_v|~clock1_v[`W-1]|ir5_v));
  assign n_400_v = ~(n_834_v);
  assign n_1486_v = ~(((n_1070_v&n_919_v)|n_200_v));
  assign n_1484_v = ~(~y2_v[`W-1]);
  assign n_790_v = ~((op_lsr_ror_dec_inc_v|op_asl_rol_v));
  assign op_push_pull_v = ~((ir7_v|irline3_v|ir4_v|~notir3_v[`W-1]|ir2_v));
  assign op_T2_v = ~(_t2_v);
  assign n_789_v = ~(~idb7_v[`W-1]);
  assign op_T__dex_v = ~((ir2_v|~notir7_v[`W-1]|ir4_v|~notir3_v[`W-1]|~notir1_v[`W-1]|clock2_v|ir5_v|~notir6_v[`W-1]));
  assign op_T0_sbc_v = ~((~notir0_v[`W-1]|~notir7_v[`W-1]|~clock1_v[`W-1]|~notir5_v[`W-1]|~notir6_v[`W-1]));
  assign n_783_v = ~(~pcl2_v[`W-1]);
  assign op_T5_rti_v = ~((_t5_v|ir3_v|ir5_v|~notir6_v[`W-1]|ir4_v|ir7_v|ir2_v|irline3_v));
  assign fetch_v = ~((~notRdy0_v[`W-1]|n_1214_v));
  assign n_782_v = ~((n_383_v&n_1303_v));
  assign op_T__cpx_cpy_abs_v = ~((~notir3_v[`W-1]|clock2_v|irline3_v|ir4_v|~notir6_v[`W-1]|~notir2_v[`W-1]|~notir7_v[`W-1]));
  assign n_951_v = ~(abl2_v);
  assign dpc34_PCLC_v = ~((n_783_v|n_937_v|n_1643_v|n_329_v|dpc36_IPC_v|n_386_v|n_641_v|n_249_v|n_232_v));
  assign n_1222_v = ~(n_1225_v);
  assign n_506_v = ~((n_192_v|n_236_v));
  assign C12_v = ~(_C12_v);
  assign n_1218_v = ~(n_1565_v);
  assign __AxB7__C67_v = ~((AxB7_v|_C67_v));
  assign AxB5_v = ~((n_647_v|~n_1632_v[`W-1]));
  assign n_1219_v = ~(op_T5_jsr_v);
  assign n_31_v = ~(p0_v);
  assign n_35_v = ~((n_796_v|~n_43_v[`W-1]));
  assign n_34_v = ~(~s3_v[`W-1]);
  assign op_T3_jmp_v = ~((irline3_v|ir7_v|~notir2_v[`W-1]|_t3_v|~notir3_v[`W-1]|ir4_v|~notir6_v[`W-1]));
  assign n_23_v = ~((dor7_v|~RnWstretched_v[`W-1]));
  assign n_25_v = ~((n_192_v|n_256_v));
  assign n_29_v = ~((~Pout3_v[`W-1]&op_T0_sbc_v));
  assign pchp5_v = ~(n_469_v);
  assign _t3_v = ~(n_678_v);
  assign n_1552_v = ~(n_1593_v);
  assign n_1517_v = ~((n_572_v|n_853_v));
  assign op_T2_abs_y_v = ~((~notir0_v[`W-1]|_t2_v|ir2_v|~notir3_v[`W-1]|~notir4_v[`W-1]));
  assign n_1523_v = ~(abh6_v);
  assign n_1521_v = ~(~x3_v[`W-1]);
  assign op_plp_pla_v = ~((ir2_v|~notir3_v[`W-1]|ir7_v|ir4_v|~notir5_v[`W-1]|irline3_v));
  assign n_1518_v = ~(n_1270_v);
  assign op_rmw_v = ~(n_790_v);
  assign n_441_v = ~(n_692_v);
  assign n_442_v = ~(n_182_v);
  assign dor3_v = ~(notdor3_v);
  assign n_466_v = ~((~RnWstretched_v[`W-1]|dor6_v));
  assign n_468_v = ~(((~notRdy0_v[`W-1]&pipeT5out_v)|(n_16_v&pipeT4out_v)));
  assign n_467_v = ~((n_470_v|n_134_v));
  assign n_1613_v = ~((dor3_v|~RnWstretched_v[`W-1]));
  assign n_472_v = ~(((pipeT4out_v&~notRdy0_v[`W-1])|(pipeT3out_v&n_16_v)));
  assign n_470_v = ~(n_646_v);
  assign n_474_v = ~(((n_1643_v&n_1184_v)|n_410_v));
  assign n_473_v = ~((n_1408_v&n_980_v));
  assign n_830_v = ~((n_1505_v|~n_43_v[`W-1]));
  assign __AxB5__C45_v = ~((_C45_v|AxB5_v));
  assign n_93_v = ~(~db0_v[`W-1]);
  assign n_90_v = ~(n_1625_v);
  assign n_80_v = ~((n_1130_v|n_267_v));
  assign op_T2_zp_zp_idx_v = ~((_t2_v|~notir2_v[`W-1]|ir3_v));
  assign op_T0_tay_ldy_not_idx_v = ~((~notir5_v[`W-1]|ir4_v|ir6_v|~notir7_v[`W-1]|~clock1_v[`W-1]|irline3_v));
  assign abh2_v = ~(~_ABH2_v[`W-1]);
  assign n_279_v = ~((n_507_v|n_954_v|n_253_v));
  assign dpc28_0ADH0_v = ~(pipedpc28_v);
  assign n_228_v = ~(n_21_v);
  assign _DA_ADD1_v = ~(~alu1_v[`W-1]);
  assign n_284_v = ~(n_1392_v);
  assign n_233_v = ~((n_761_v&n_149_v));
  assign n_225_v = ~(n_1223_v);
  assign op_T4_ind_y_v = ~((ir3_v|~notir0_v[`W-1]|_t4_v|~notir4_v[`W-1]|ir2_v));
  assign n_491_v = ~(n_1541_v);
  assign n_504_v = ~((n_1120_v&n_440_v));
  assign n_503_v = ~(~notir5_v[`W-1]);
  assign C56_v = ~(_C56_v);
  assign n_499_v = ~(~pch5_v[`W-1]);
  assign n_490_v = ~(~db4_v[`W-1]);
  assign n_501_v = ~((Reset0_v|n_819_v|n_180_v));
  assign n_496_v = ~(~s5_v[`W-1]);
  assign op_T5_ind_y_v = ~((ir3_v|~notir4_v[`W-1]|~notir0_v[`W-1]|_t5_v|ir2_v));
  assign n_862_v = ~(n_666_v);
  assign n_253_v = ~(pipeUNK42_v);
  assign A_B7_v = ~(~n_1398_v[`W-1]);
  assign n_110_v = ~(~n_1691_v[`W-1]);
  assign n_122_v = ~(~__AxB_6_v[`W-1]);
  assign n_108_v = ~(n_1364_v);
  assign n_111_v = ~(~db2_v[`W-1]);
  assign n_118_v = ~(n_334_v);
  assign n_109_v = ~(n_1380_v);
  assign pchp1_v = ~(n_126_v);
  assign op_T3_v = ~(_t3_v);
  assign n_930_v = ~((n_1276_v|n_134_v));
  assign n_347_v = ~((op_T4_mem_abs_idx_v|op_T3_mem_zp_idx_v|op_T2_mem_zp_v|op_T3_mem_abs_v|op_T5_mem_ind_idx_v));
  assign n_340_v = ~(op_clv_v);
  assign n_1585_v = ~(~cclk_v[`W-1]);
  assign n_1578_v = ~(pipe_VEC_v);
  assign pd3_clearIR_v = ~((clearIR_v|pd3_v));
  assign op_T2_stack_v = ~((irline3_v|ir4_v|ir7_v|_t2_v|ir2_v));
  assign ir3_v = ~(~n_1620_v[`W-1]);
  assign x_op_T3_abs_idx_v = ~((~notir3_v[`W-1]|~notir4_v[`W-1]|_t3_v));
  assign n_1580_v = ~(~sb2_v[`W-1]);
  assign n_1575_v = ~((n_1357_v|n_1360_v));
  assign n_445_v = ~(n_862_v);
  assign op_T5_rti_rts_v = ~((ir3_v|_t5_v|irline3_v|ir2_v|~notir6_v[`W-1]|ir7_v|ir4_v));
  assign n_629_v = ~((n_50_v|((n_646_v|nnT2BR_v)&n_480_v)));
  assign n_1002_v = ~(n_1219_v);
  assign op_implied_v = ~((~notir3_v[`W-1]|x_op_push_pull_v|ir2_v|ir0_v));
  assign _C23_v = ~(C23_v);
  assign n_1007_v = ~(dpc34_PCLC_v);
  assign n_1010_v = ~(~pch0_v[`W-1]);
  assign n_1018_v = ~(n_762_v);
  assign n_1017_v = ~(~x5_v[`W-1]);
  assign n_70_v = ~((_VEC_v|n_1054_v));
  assign n_1439_v = ~(~y6_v[`W-1]);
  assign n_551_v = ~(n_393_v);
  assign op_T0_php_pha_v = ~((ir2_v|ir4_v|ir7_v|~notir3_v[`W-1]|ir5_v|~clock1_v[`W-1]|irline3_v));
  assign n_275_v = ~((n_1697_v|n_773_v));
  assign n_1610_v = ~((AxB3_v|DA_AB2_v));
  assign op_T4_rts_v = ~((ir3_v|ir2_v|irline3_v|~notir6_v[`W-1]|_t4_v|ir4_v|~notir5_v[`W-1]|ir7_v));
  assign n_1619_v = ~((n_182_v|n_1448_v));
  assign pd0_clearIR_v = ~((pd0_v|clearIR_v));
  assign op_T0_eor_v = ~((~notir6_v[`W-1]|ir5_v|~notir0_v[`W-1]|ir7_v|~clock1_v[`W-1]));
  assign ir1_v = ~(~n_119_v[`W-1]);
  assign n_550_v = ~((n_384_v|op_ANDS_v));
  assign n_1511_v = ~(pipeUNK29_v);
  assign n_958_v = ~(~rdy_v[`W-1]);
  assign n_956_v = ~(n_476_v);
  assign n_954_v = ~(pipeUNK08_v);
  assign n_952_v = ~(n_272_v);
  assign n_964_v = ~((pipe_T0_v|n_1533_v));
  assign n_708_v = ~(n_1230_v);
  assign n_700_v = ~(~dpc18__DAA_v[`W-1]);
  assign abh1_v = ~(~_ABH1_v[`W-1]);
  assign n_714_v = ~(n_906_v);
  assign n_638_v = ~(op_T0_v);
  assign n_632_v = ~((op_T2_stack_v|(op_T0_jsr_v&n_1289_v)));
  assign op_T0_cld_sed_v = ~((~notir4_v[`W-1]|ir2_v|irline3_v|~notir3_v[`W-1]|~clock1_v[`W-1]|~notir7_v[`W-1]|~notir6_v[`W-1]));
  assign dor6_v = ~(notdor6_v);
  assign n_207_v = ~(((n_923_v&n_293_v)|n_810_v));
  assign n_645_v = ~(~NMIP_v[`W-1]);
  assign n_646_v = ~(n_17_v);
  assign AxB3_v = ~((n_988_v|~n_649_v[`W-1]));
  assign n_641_v = ~(~pcl7_v[`W-1]);
  assign n_637_v = ~((C67_v|~n_1318_v[`W-1]));
  assign n_1205_v = ~(((n_1257_v&n_233_v)|(n_1018_v&n_811_v)));
  assign op_T5_ind_x_v = ~((~notir0_v[`W-1]|ir4_v|_t5_v|ir3_v|ir2_v));
  assign n_1209_v = ~(((n_609_v&n_453_v)|n_1213_v));
  assign op_T2_ind_y_v = ~((ir2_v|~notir0_v[`W-1]|ir3_v|_t2_v|~notir4_v[`W-1]));
  assign clock2_v = ~(n_1533_v);
  assign C45_v = ~(((~n_1063_v[`W-1]&_C34_v)|~n_404_v[`W-1]));
  assign n_1211_v = ~((n_1002_v|nnT2BR_v|n_1286_v|op_T2_abs_access_v|n_862_v));
  assign n_38_v = ~(~cp1_v[`W-1]);
  assign n_1202_v = ~(n_1265_v);
  assign n_1199_v = ~(~db2_v[`W-1]);
  assign op_T__ora_and_eor_adc_v = ~((~notir0_v[`W-1]|clock2_v|ir7_v));
  assign n_1244_v = ~(op_xy_v);
  assign n_1245_v = ~(aluvout_v);
  assign op_shift_right_v = ~((~notir6_v[`W-1]|~notir1_v[`W-1]|ir7_v));
  assign ir5_v = ~(~n_1609_v[`W-1]);
  assign ir7_v = ~(~n_541_v[`W-1]);
  assign n_1335_v = ~(n_628_v);
  assign dpc35_PCHC_v = ~((n_1010_v|n_1007_v|n_923_v|n_1070_v|n_1265_v));
  assign op_T__shift_a_v = ~((~notir3_v[`W-1]|clock2_v|ir2_v|ir4_v|~notir1_v[`W-1]|ir7_v));
  assign n_1323_v = ~(n_631_v);
  assign n_480_v = ~(((n_888_v|n_118_v)&n_264_v));
  assign n_479_v = ~((n_61_v|n_739_v));
  assign n_485_v = ~(~x4_v[`W-1]);
  assign n_484_v = ~(((n_1316_v|n_715_v)&n_1386_v));
  assign n_256_v = ~((op_T5_rti_v|op_T5_rts_v|op_T5_ind_x_v|op_T0_jmp_v|op_T4_v|op_T3_v|op_T0_brk_rti_v));
  assign n_255_v = ~(n_611_v);
  assign abh7_v = ~(~_ABH7_v[`W-1]);
  assign op_T0_tya_v = ~((~notir4_v[`W-1]|~notir7_v[`W-1]|ir2_v|~clock1_v[`W-1]|ir6_v|~notir3_v[`W-1]|ir5_v|irline3_v));
  assign _op_branch_bit6_v = ~(ir6_v);
  assign op_T2_brk_v = ~((_t2_v|ir3_v|ir7_v|ir5_v|ir2_v|ir4_v|irline3_v|ir6_v));
  assign __AxB1__C01_v = ~((_C01_v|AxB1_v));
  assign n_293_v = ~((n_200_v&n_1202_v));
  assign abl4_v = ~(~_ABL4_v[`W-1]);
  assign op_T0_plp_v = ~((ir2_v|irline3_v|~notir3_v[`W-1]|ir6_v|ir7_v|ir4_v|~notir5_v[`W-1]|~clock1_v[`W-1]));
  assign pclp0_v = ~(n_526_v);
  assign op_T4_jmp_v = ~((~notir2_v[`W-1]|~notir6_v[`W-1]|irline3_v|ir4_v|~notir3_v[`W-1]|_t4_v|ir7_v));
  assign n_1229_v = ~(((dpc34_PCLC_v|n_311_v)&n_919_v));
  assign n_1230_v = ~((~n_43_v[`W-1]|n_360_v));
  assign n_918_v = ~(~n_404_v[`W-1]);
  assign n_1629_v = ~((n_753_v|n_1135_v));
  assign n_1631_v = ~(((n_163_v|n_1253_v)&n_1184_v));
  assign dor2_v = ~(notdor2_v);
  assign alucin_v = ~(n_590_v);
  assign n_917_v = ~((n_383_v|~notRdy0_v[`W-1]));
  assign n_916_v = ~(((~n_206_v[`W-1]&n_853_v)|n_1517_v));
  assign n_919_v = ~((n_311_v&dpc34_PCLC_v));
  assign n_1635_v = ~(n_966_v);
  assign n_1638_v = ~(~db6_v[`W-1]);
  assign n_1400_v = ~(~pch4_v[`W-1]);
  assign PD_xxx010x1_v = ~((pd2_clearIR_v|~n_1083_v[`W-1]|pd4_clearIR_v|~n_409_v[`W-1]));
  assign n_1446_v = ~((n_850_v|n_771_v));
  assign op_T2_php_pha_v = ~((_t2_v|ir2_v|~notir3_v[`W-1]|ir7_v|ir5_v|ir4_v|irline3_v));
  assign n_920_v = ~(pipeUNK27_v);
  assign _op_store_v = ~(op_store_v);
  assign n_604_v = ~(((op_T4_rti_v|op_T4_brk_jsr_v|op_T3_ind_x_v|op_T2_stack_v|~notRdy0_v[`W-1]|op_T3_stack_bit_jmp_v)|(op_T2_ADL_ADD_v&n_638_v)));
  assign n_36_v = ~((n_8_v|n_600_v));
  assign n_602_v = ~(n_133_v);
  assign pclp4_v = ~(n_15_v);
  assign dor7_v = ~(notdor7_v);
  assign n_62_v = ~(~db7_v[`W-1]);
  assign n_613_v = ~(((_DA_ADD1_v&n_600_v)|(n_8_v&n_1682_v)));
  assign n_611_v = ~((n_1509_v|~n_43_v[`W-1]));
  assign brk_done_v = ~((n_861_v|~notRdy0_v[`W-1]));
  assign ir2_v = ~(~n_1300_v[`W-1]);
  assign n_1115_v = ~((n_620_v|n_270_v));
  assign op_T0_clc_sec_v = ~((~notir4_v[`W-1]|irline3_v|ir6_v|ir2_v|ir7_v|~notir3_v[`W-1]|~clock1_v[`W-1]));
  assign ir4_v = ~(~n_927_v[`W-1]);
  assign n_1111_v = ~((pipeUNK07_v&pipeUNK09_v));
  assign notalucout_v = ~((C78_phi2_v|DC78_phi2_v));
  assign n_1677_v = ~(abh4_v);
  assign abh3_v = ~(~_ABH3_v[`W-1]);
  assign n_410_v = ~((n_1643_v|n_1184_v));
  assign AxB1_v = ~((n_936_v|~aluanorb1_v[`W-1]));
  assign n_419_v = ~(~a2_v[`W-1]);
  assign n_1106_v = ~(((op_from_x_v&n_335_v)|(op_T0_cpx_inx_v|op_T0_txs_v|op_T2_ind_x_v|x_op_T0_txa_v|op_T0_dex_v)|(op_T2_idx_x_xy_v&n_1244_v)));
  assign n_1101_v = ~((n_813_v&n_46_v));
  assign n_1099_v = ~((n_1542_v&(n_1166_v|n_1345_v)));
  assign n_1110_v = ~(n_756_v);
  assign n_1109_v = ~((n_1464_v|n_902_v));
  assign n_329_v = ~(~pcl1_v[`W-1]);
  assign op_inc_nop_v = ~((~notir5_v[`W-1]|~notir1_v[`W-1]|~notir6_v[`W-1]|~notir7_v[`W-1]));
  assign ir0_v = ~(~n_310_v[`W-1]);
  assign n_1093_v = ~(n_968_v);
  assign n_1107_v = ~(((n_440_v&op_inc_nop_v)|(op_T4_ind_y_v|op_T2_ind_y_v|op_plp_pla_v|op_T3_abs_idx_v|op_T3_ind_x_v)));
  assign op_T3_abs_idx_ind_v = ~((_t3_v|op_push_pull_v|~notir3_v[`W-1]));
  assign _t4_v = ~(n_188_v);
  assign DA_AB2_v = ~(~n_681_v[`W-1]);
  assign n_696_v = ~((((n_1343_v|n_877_v)&n_79_v)|n_0_ADL0_v));
  assign aluaorb0_v = ~(~aluanorb0_v[`W-1]);
  assign n_1081_v = ~(n_1560_v);
  assign _DA_ADD2_v = ~(~alu2_v[`W-1]);
  assign n_689_v = ~(op_T5_brk_v);
  assign op_asl_rol_v = ~((~notir1_v[`W-1]|ir7_v|ir6_v));
  assign n_692_v = ~((n_460_v|~n_43_v[`W-1]));
  assign n_695_v = ~((C34_v&n_700_v));
  assign C23_v = ~((~n_1691_v[`W-1]|(_C12_v&~n_681_v[`W-1])));
  assign n_1281_v = ~(~db3_v[`W-1]);
  assign C01_v = ~((~aluanorb0_v[`W-1]|(notalucin_v&~aluanandb0_v[`W-1])));
  assign n_1275_v = ~((ONEBYTE_v|~notRdy0_v[`W-1]|pipeBRtaken_v));
  assign n_1277_v = ~(n_1020_v);
  assign n_1286_v = ~((n_470_v|n_930_v));
  assign n_1289_v = ~(n_902_v);
  assign n_1033_v = ~(n_241_v);
  assign n_1024_v = ~(n_94_v);
  assign n_1541_v = ~((~n_43_v[`W-1]|n_1477_v));
  assign n_811_v = ~((alucout_v|n_838_v));
  assign n_812_v = ~((n_646_v|n_440_v));
  assign C78_v = ~(_C78_v);
  assign pd1_clearIR_v = ~((clearIR_v|pd1_v));
  assign n_810_v = ~((n_293_v|n_923_v));
  assign n_797_v = ~(~idb4_v[`W-1]);
  assign n_800_v = ~(n_525_v);
  assign x_op_T0_txa_v = ~((ir2_v|~notir7_v[`W-1]|ir4_v|ir6_v|~notir3_v[`W-1]|ir5_v|~notir1_v[`W-1]|~clock1_v[`W-1]));
  assign n_1542_v = ~((n_1166_v&n_1345_v));
  assign A_B1_v = ~(~aluanorb1_v[`W-1]);
  assign op_T0_ora_v = ~((~clock1_v[`W-1]|ir7_v|ir6_v|ir5_v|~notir0_v[`W-1]));
  assign op_T0_tsx_v = ~((~notir3_v[`W-1]|ir6_v|~notir4_v[`W-1]|~notir5_v[`W-1]|ir2_v|~clock1_v[`W-1]|~notir1_v[`W-1]|~notir7_v[`W-1]));
  assign n_0_ADL1_v = ~(pipeVectorA1_v);
  assign n_71_v = ~(n_35_v);
  assign C34_v = ~(_C34_v);
  assign n_79_v = ~(n_236_v);
  assign n_1375_v = ~(n_88_v);
  assign n_1374_v = ~((n_562_v|n_882_v));
  assign n_1358_v = ~((n_917_v|op_T0_txs_v|n_1109_v));
  assign n_1357_v = ~(n_223_v);
  assign n_1368_v = ~((n_1578_v|n_1374_v|n_645_v));
  assign n_1364_v = ~(n_101_v);
  assign n_1369_v = ~(n_897_v);
  assign INTG_v = ~((n_760_v|brk_done_v));
  assign _WR_v = ~((n_1258_v|op_T4_brk_v|n_440_v|op_T2_php_pha_v|n_335_v|n_1642_v));
  assign n_1356_v = ~(~a6_v[`W-1]);
  assign n_17_v = ~((n_732_v|n_964_v));
  assign n_16_v = ~(~notRdy0_v[`W-1]);
  assign n_14_v = ~((n_323_v|Reset0_v|n_671_v));
  assign n_11_v = ~(((op_T0_acc_v&n_397_v)|(op_T0_shift_a_v|op_T0_tay_v|op_T0_tax_v|op_ANDS_v)));
  assign n_10_v = ~((op_branch_done_v|n_1211_v|n_467_v));
  assign n_630_v = ~(n_726_v);
  assign n_201_v = ~(_op_branch_bit7_v);
  assign n_196_v = ~(n_543_v);
  assign _AxB_2__C12_v = ~((~__AxB_2_v[`W-1]|C12_v));
  assign n_200_v = ~((n_1070_v|n_919_v));
  assign n_198_v = ~(pipeUNK37_v);
  assign n_1154_v = ~((n_959_v|~notRdy0_v[`W-1]));
  assign n_1153_v = ~(abh7_v);
  assign n_1166_v = ~(n_329_v);
  assign notalucin_v = ~(alucin_v);
  assign op_T0_acc_v = ~((~clock1_v[`W-1]|~notir0_v[`W-1]));
  assign n_983_v = ~(~s0_v[`W-1]);
  assign n_987_v = ~(~x0_v[`W-1]);
  assign n_986_v = ~((_DA_ADD2_v&_DA_ADD1_v));
  assign n_990_v = ~(abl3_v);
  assign n_1614_v = ~((n_1177_v|n_1111_v|pipeUNK03_v));
  assign abh6_v = ~(~_ABH6_v[`W-1]);
  assign irline3_v = ~(n_1133_v);
  assign op_T0_ldx_tax_tsx_v = ~((ir6_v|~notir7_v[`W-1]|~notir5_v[`W-1]|~notir1_v[`W-1]|~clock1_v[`W-1]));
  assign n_988_v = ~(~n_350_v[`W-1]);
  assign n_995_v = ~(n_312_v);
  assign n_889_v = ~(op_T0_clc_sec_v);
  assign n_888_v = ~(n_675_v);
  assign n_882_v = ~((n_1252_v|n_597_v));
  assign n_885_v = ~(n_384_v);
  assign n_1315_v = ~(abh0_v);
  assign C67_v = ~(((_C56_v&~n_336_v[`W-1])|~n_1084_v[`W-1]));
  assign n_890_v = ~(~x2_v[`W-1]);
  assign n_1316_v = ~((n_344_v|n_232_v));
  assign op_EORS_v = ~(n_837_v);
  assign n_896_v = ~(~db3_v[`W-1]);
  assign n_1712_v = ~((n_264_v|C1x5Reset_v|_VEC_v));
  assign op_T0_jmp_v = ~((ir4_v|~clock1_v[`W-1]|~notir3_v[`W-1]|irline3_v|~notir6_v[`W-1]|~notir2_v[`W-1]|ir7_v));
  assign op_T__cpx_cpy_imm_zp_v = ~((ir4_v|~notir6_v[`W-1]|irline3_v|~notir7_v[`W-1]|clock2_v|ir3_v));
  assign n_1711_v = ~(~s1_v[`W-1]);
  assign n_1716_v = ~((n_510_v|op_T3_branch_v|n_218_v|n_1258_v));
  assign n_1717_v = ~(((op_T2_idx_x_xy_v&op_xy_v)|(n_335_v&op_sty_cpy_mem_v)|(op_T0_cpy_iny_v|op_T2_abs_y_v|op_T3_ind_y_v|x_op_T0_tya_v|op_T0_iny_dey_v)));
  assign n_1714_v = ~(pipeUNK26_v);
  assign n_1715_v = ~(n_358_v);
  assign n_595_v = ~((op_T4_abs_idx_v|op_T5_ind_y_v));
  assign n_586_v = ~(((BRtaken_v&nnT2BR_v)|n_1619_v));
  assign n_1047_v = ~(n_830_v);
  assign x_op_jmp_v = ~((irline3_v|~notir3_v[`W-1]|ir4_v|ir7_v|~notir2_v[`W-1]|~notir6_v[`W-1]));
  assign x_op_push_pull_v = ~((irline3_v|ir7_v|ir4_v|ir2_v|~notir3_v[`W-1]));
  assign op_T2_php_v = ~((ir6_v|ir5_v|irline3_v|ir4_v|_t2_v|ir7_v|ir2_v|~notir3_v[`W-1]));
  assign n_1054_v = ~(C1x5Reset_v);
  assign op_T2_abs_v = ~((ir4_v|_t2_v|~notir3_v[`W-1]|~notir2_v[`W-1]));
  assign n_1056_v = ~(n_761_v);
  assign _op_branch_done_v = ~(op_branch_done_v);
  assign n_753_v = ~((n_811_v|n_1257_v));
  assign n_735_v = ~((n_320_v|n_36_v));
  assign n_1463_v = ~((dor4_v|~RnWstretched_v[`W-1]));
  assign n_1462_v = ~(n_1369_v);
  assign pd6_clearIR_v = ~((clearIR_v|pd6_v));
  assign n_1474_v = ~(~idb1_v[`W-1]);
  assign op_T5_jsr_v = ~((_t5_v|ir4_v|ir6_v|ir3_v|~notir5_v[`W-1]|ir2_v|irline3_v|ir7_v));
  assign n_1471_v = ~(D1x1_v);
  assign op_rol_ror_v = ~((~notir5_v[`W-1]|ir7_v|ir6_v|~notir1_v[`W-1]));
  assign n_774_v = ~(op_T0_cld_sed_v);
  assign ONEBYTE_v = ~(n_231_v);
  assign n_1043_v = ~(n_818_v);
  assign n_1044_v = ~((n_812_v|n_31_v));
  assign _DBE_v = ~((n_962_v|~cclk_v[`W-1]));
  assign n_1037_v = ~((op_T2_pha_v|(op_sta_cmp_v&n_335_v)));
  assign n_1038_v = ~(~n_336_v[`W-1]);
  assign n_1039_v = ~((pipeUNK40_v|(pipeUNK39_v&~notRdy0_v[`W-1])));
  assign n_600_v = ~(n_1341_v);
  assign n_603_v = ~(n_47_v);
  assign n_1045_v = ~(n_69_v);
  assign n_1034_v = ~(abh2_v);
  assign n_743_v = ~((n_499_v|n_523_v));
  assign dor1_v = ~(notdor1_v);
  assign notRnWprepad_v = ~((~notRdy0_v[`W-1]|pipe_WR_phi2_v|C1x5Reset_v));
  assign n_188_v = ~((n_1357_v|n_1606_v));
  assign n_1097_v = ~((n_432_v|n_345_v));
  assign abl0_v = ~(~_ABL0_v[`W-1]);
  assign n_191_v = ~((n_347_v|~notRdy0_v[`W-1]|n_790_v));
  assign n_192_v = ~((n_595_v&_op_branch_done_v));
  assign n_180_v = ~((~notRdy0_v[`W-1]|n_1716_v));
  assign abl6_v = ~(~_ABL6_v[`W-1]);
  assign n_182_v = ~(((n_1262_v&n_236_v)|(n_646_v|op_T5_rts_v|n_1655_v)));
  assign n_184_v = ~(~y3_v[`W-1]);
  assign op_T0_adc_sbc_v = ~((~notir6_v[`W-1]|~clock1_v[`W-1]|~notir5_v[`W-1]|~notir0_v[`W-1]));
  assign n_565_v = ~(~y4_v[`W-1]);
  assign n_1255_v = ~(n_531_v);
  assign n_160_v = ~((n_781_v|op_SRS_v));
  assign n_1257_v = ~((n_1218_v|notalucout_v));
  assign n_1253_v = ~((n_783_v|n_1542_v));
  assign op_T4_ind_x_v = ~((ir3_v|ir2_v|ir4_v|~notir0_v[`W-1]|_t4_v));
  assign n_1256_v = ~(n_91_v);
  assign n_1262_v = ~(n_1679_v);
  assign n_1258_v = ~(n_390_v);
  assign n_169_v = ~((n_139_v|n_1624_v));
  assign n_172_v = ~(abl5_v);
  assign ir6_v = ~(~n_1675_v[`W-1]);
  assign _AxB_6__C56_v = ~((C56_v|~__AxB_6_v[`W-1]));
  assign n_176_v = ~((n_236_v|n_10_v));
  assign n_344_v = ~((n_410_v&n_392_v));
  assign x_op_T3_ind_y_v = ~((_t3_v|ir3_v|ir2_v|~notir4_v[`W-1]|~notir0_v[`W-1]));
  assign op_T4_v = ~(_t4_v);
  assign n_959_v = ~((~n_430_v[`W-1]|pipeUNK20_v));
  assign pd2_clearIR_v = ~((clearIR_v|pd2_v));
  assign n_307_v = ~((_op_branch_bit7_v|n_846_v|n_31_v));
  assign op_T__inx_v = ~((irline3_v|clock2_v|~notir5_v[`W-1]|~notir6_v[`W-1]|ir2_v|~notir7_v[`W-1]|~notir3_v[`W-1]|ir4_v));
  assign n_1682_v = ~(_DA_ADD1_v);
  assign n_1660_v = ~(abl0_v);
  assign op_T__asl_rol_a_v = ~((clock2_v|ir7_v|ir6_v|ir4_v|~notir3_v[`W-1]|ir2_v|~notir1_v[`W-1]));
  assign n_1676_v = ~(abl4_v);
  assign n_1662_v = ~(n_1124_v);
  assign n_1455_v = ~((op_T__adc_sbc_v|op_T0_tya_v|op_T__shift_a_v|op_T0_txa_v|op_T__ora_and_eor_adc_v|op_T0_pla_v|op_T0_lda_v));
  assign n_1457_v = ~((n_1492_v|n_781_v));
  assign n_1441_v = ~(n_1277_v);
  assign n_1448_v = ~(n_1427_v);
  assign n_355_v = ~(n_621_v);
  assign op_T4_abs_idx_v = ~((_t4_v|~notir4_v[`W-1]|~notir3_v[`W-1]));
  assign op_T4_brk_v = ~((ir4_v|ir3_v|irline3_v|_t4_v|ir2_v|ir5_v|ir6_v|ir7_v));
  assign n_366_v = ~((op_T0_shift_right_a_v|(n_440_v&op_shift_right_v)));
  assign PD_0xx0xx0x_v = ~((pd7_clearIR_v|pd1_clearIR_v|pd4_clearIR_v));
  assign n_538_v = ~(n_1599_v);
  assign pd4_clearIR_v = ~((clearIR_v|pd4_v));
  assign n_1649_v = ~((brk_done_v|n_389_v|op_T4_ind_x_v|op_jmp_v|~notRdy0_v[`W-1]|op_T2_jsr_v|n_1109_v|op_rti_rts_v|op_T2_abs_v));
  assign n_1650_v = ~(~so_v[`W-1]);
  assign n_1642_v = ~((n_462_v&n_824_v));
  assign n_1643_v = ~(~pcl4_v[`W-1]);
  assign op_T__bit_v = ~((irline3_v|~notir2_v[`W-1]|ir6_v|ir7_v|clock2_v|~notir5_v[`W-1]|ir4_v));
  assign _TWOCYCLE_v = ~(((PD_n_0xx0xx0x_v&PD_xxxx10x0_v)|(PD_1xx000x0_v|PD_xxx010x1_v)));
  assign op_ORS_v = ~(n_1145_v);
  assign n_523_v = ~((dpc35_PCHC_v&n_83_v));
  assign n_1141_v = ~(n_982_v);
  assign n_132_v = ~(n_31_v);
  assign n_133_v = ~((n_1404_v|~cclk_v[`W-1]));
  assign n_130_v = ~(n_220_v);
  assign op_T0_pla_v = ~((~notir5_v[`W-1]|ir2_v|ir7_v|~clock1_v[`W-1]|ir4_v|irline3_v|~notir3_v[`W-1]|~notir6_v[`W-1]));
  assign n_127_v = ~((~cp1_v[`W-1]|n_519_v));
  assign n_128_v = ~(~a7_v[`W-1]);
  assign pchp3_v = ~(n_1061_v);
  assign PD_n_0xx0xx0x_v = ~(PD_0xx0xx0x_v);
  assign n_134_v = ~((x_op_jmp_v|op_brk_rti_v|op_jsr_v));
  assign n_139_v = ~(op_SRS_v);
  assign op_sta_cmp_v = ~((~notir7_v[`W-1]|ir5_v|~notir0_v[`W-1]|ir6_v));
  assign n_1133_v = ~((ir1_v|ir0_v));
  assign _VEC_v = ~((VEC1_v|VEC0_v));
  assign n_1135_v = ~(~sb5_v[`W-1]);
  assign n_1137_v = ~((n_790_v&_op_store_v));
  assign abh4_v = ~(~_ABH4_v[`W-1]);
  assign DA_C45_v = ~(_C45_v);
  assign n_1129_v = ~((n_358_v|~cp1_v[`W-1]));
  assign n_1130_v = ~((n_862_v|n_1258_v|n_1002_v|n_192_v|n_1109_v));
  assign n_1138_v = ~(~y1_v[`W-1]);
  assign n_476_v = ~((~n_43_v[`W-1]|n_1027_v));
  assign x_op_T4_rti_v = ~((_t4_v|ir2_v|irline3_v|~notir6_v[`W-1]|ir5_v|ir3_v|ir7_v|ir4_v));
  assign n_1560_v = ~((n_1055_v|op_T0_cpx_cpy_inx_iny_v|op_T0_cmp_v));
  assign n_1561_v = ~(~x7_v[`W-1]);
  assign op_xy_v = ~((~notir1_v[`W-1]|ir6_v|~notir7_v[`W-1]));
  assign n_1566_v = ~(n_1221_v);
  assign n_1573_v = ~(~idb2_v[`W-1]);
  assign n_795_v = ~(n_1649_v);
  assign op_brk_rti_v = ~((irline3_v|ir7_v|ir5_v|ir2_v|ir3_v|ir4_v));
  assign _C45_v = ~(C45_v);

  spice_node_2 n_n_1247(eclk, ereset, n_1247_port_13,n_1247_port_0, n_1247_v);
  spice_node_2 n__ABL7(eclk, ereset, _ABL7_port_3,_ABL7_port_1, _ABL7_v);
  spice_node_2 n__ABL6(eclk, ereset, _ABL6_port_3,_ABL6_port_1, _ABL6_v);
  spice_node_2 n__ABL5(eclk, ereset, _ABL5_port_3,_ABL5_port_0, _ABL5_v);
  spice_node_2 n__ABL3(eclk, ereset, _ABL3_port_3,_ABL3_port_0, _ABL3_v);
  spice_node_2 n__ABL2(eclk, ereset, _ABL2_port_2,_ABL2_port_3, _ABL2_v);
  spice_node_2 n__ABL1(eclk, ereset, _ABL1_port_2,_ABL1_port_3, _ABL1_v);
  spice_node_2 n__ABL0(eclk, ereset, _ABL0_port_2,_ABL0_port_3, _ABL0_v);
  spice_node_2 n_dpc5_SADL(eclk, ereset, dpc5_SADL_port_0,dpc5_SADL_port_7, dpc5_SADL_v);
  spice_node_3 n_n_465(eclk, ereset, n_465_port_2,n_465_port_0,n_465_port_1, n_465_v);
  spice_node_2 n_rw(eclk, ereset, rw_port_0,rw_port_1, rw_v);
  spice_node_3 n_idl7(eclk, ereset, idl7_port_2,idl7_port_0,idl7_port_1, idl7_v);
  spice_node_3 n_idl6(eclk, ereset, idl6_port_2,idl6_port_0,idl6_port_1, idl6_v);
  spice_node_3 n_idl5(eclk, ereset, idl5_port_2,idl5_port_0,idl5_port_1, idl5_v);
  spice_node_3 n_idl4(eclk, ereset, idl4_port_2,idl4_port_0,idl4_port_1, idl4_v);
  spice_node_3 n_idl3(eclk, ereset, idl3_port_2,idl3_port_0,idl3_port_1, idl3_v);
  spice_node_3 n_idl2(eclk, ereset, idl2_port_2,idl2_port_0,idl2_port_1, idl2_v);
  spice_node_3 n_idl1(eclk, ereset, idl1_port_2,idl1_port_0,idl1_port_1, idl1_v);
  spice_node_3 n_idl0(eclk, ereset, idl0_port_2,idl0_port_0,idl0_port_1, idl0_v);
  spice_node_4 n_n_733(eclk, ereset, n_733_port_2,n_733_port_3,n_733_port_0,n_733_port_1, n_733_v);
  spice_node_2 n_dpc20_ADDSB06(eclk, ereset, dpc20_ADDSB06_port_0,dpc20_ADDSB06_port_5, dpc20_ADDSB06_v);
  spice_node_5 n_n_1389(eclk, ereset, n_1389_port_2,n_1389_port_3,n_1389_port_0,n_1389_port_1,n_1389_port_4, n_1389_v);
  spice_node_4 n_n_1387(eclk, ereset, n_1387_port_2,n_1387_port_3,n_1387_port_0,n_1387_port_1, n_1387_v);
  spice_node_3 n_n_1383(eclk, ereset, n_1383_port_2,n_1383_port_0,n_1383_port_1, n_1383_v);
  spice_node_2 n_x6(eclk, ereset, x6_port_0,x6_port_1, x6_v);
  spice_node_1 n_irq(eclk, ereset, irq_port_2, irq_v);
  spice_node_3 n_n_1267(eclk, ereset, n_1267_port_2,n_1267_port_3,n_1267_port_0, n_1267_v);
  spice_node_2 n_n_7(eclk, ereset, n_7_port_2,n_7_port_4, n_7_v);
  spice_node_5 n_n_3(eclk, ereset, n_3_port_2,n_3_port_3,n_3_port_0,n_3_port_1,n_3_port_4, n_3_v);
  spice_node_3 n_aluanandb0(eclk, ereset, aluanandb0_port_9,aluanandb0_port_3,aluanandb0_port_5, aluanandb0_v);
  spice_node_4 n_aluanandb1(eclk, ereset, aluanandb1_port_0,aluanandb1_port_1,aluanandb1_port_4,aluanandb1_port_5, aluanandb1_v);
  spice_node_3 n_dasb6(eclk, ereset, dasb6_port_3,dasb6_port_0,dasb6_port_5, dasb6_v);
  spice_node_3 n_dasb5(eclk, ereset, dasb5_port_3,dasb5_port_1,dasb5_port_5, dasb5_v);
  spice_node_3 n_dasb3(eclk, ereset, dasb3_port_3,dasb3_port_1,dasb3_port_5, dasb3_v);
  spice_node_3 n_dasb2(eclk, ereset, dasb2_port_3,dasb2_port_1,dasb2_port_5, dasb2_v);
  spice_node_3 n_dasb1(eclk, ereset, dasb1_port_3,dasb1_port_0,dasb1_port_5, dasb1_v);
  spice_node_4 n_alu4(eclk, ereset, alu4_port_2,alu4_port_3,alu4_port_0,alu4_port_1, alu4_v);
  spice_node_4 n_alu5(eclk, ereset, alu5_port_3,alu5_port_0,alu5_port_1,alu5_port_4, alu5_v);
  spice_node_4 n_alu6(eclk, ereset, alu6_port_2,alu6_port_0,alu6_port_1,alu6_port_4, alu6_v);
  spice_node_4 n_alu7(eclk, ereset, alu7_port_2,alu7_port_3,alu7_port_0,alu7_port_1, alu7_v);
  spice_node_4 n_alu0(eclk, ereset, alu0_port_2,alu0_port_3,alu0_port_0,alu0_port_1, alu0_v);
  spice_node_4 n_alu1(eclk, ereset, alu1_port_3,alu1_port_0,alu1_port_1,alu1_port_4, alu1_v);
  spice_node_4 n_alu2(eclk, ereset, alu2_port_3,alu2_port_0,alu2_port_1,alu2_port_4, alu2_v);
  spice_node_4 n_alu3(eclk, ereset, alu3_port_2,alu3_port_3,alu3_port_0,alu3_port_1, alu3_v);
  spice_node_2 n__ABL4(eclk, ereset, _ABL4_port_3,_ABL4_port_1, _ABL4_v);
  spice_node_5 n_n_488(eclk, ereset, n_488_port_2,n_488_port_3,n_488_port_0,n_488_port_1,n_488_port_4, n_488_v);
  spice_node_5 n_n_481(eclk, ereset, n_481_port_2,n_481_port_3,n_481_port_0,n_481_port_1,n_481_port_4, n_481_v);
  spice_node_5 n_n_326(eclk, ereset, n_326_port_2,n_326_port_3,n_326_port_0,n_326_port_1,n_326_port_4, n_326_v);
  spice_node_2 n_n_1105(eclk, ereset, n_1105_port_2,n_1105_port_0, n_1105_v);
  spice_node_3 n_n_1100(eclk, ereset, n_1100_port_2,n_1100_port_3,n_1100_port_0, n_1100_v);
  spice_node_2 n_dpc6_SBS(eclk, ereset, dpc6_SBS_port_11,dpc6_SBS_port_12, dpc6_SBS_v);
  spice_node_5 n_n_831(eclk, ereset, n_831_port_2,n_831_port_3,n_831_port_0,n_831_port_1,n_831_port_4, n_831_v);
  spice_node_2 n_s3(eclk, ereset, s3_port_0,s3_port_1, s3_v);
  spice_node_2 n_s2(eclk, ereset, s2_port_0,s2_port_1, s2_v);
  spice_node_2 n_s1(eclk, ereset, s1_port_0,s1_port_1, s1_v);
  spice_node_2 n_s0(eclk, ereset, s0_port_0,s0_port_1, s0_v);
  spice_node_2 n_s7(eclk, ereset, s7_port_2,s7_port_0, s7_v);
  spice_node_2 n_s6(eclk, ereset, s6_port_0,s6_port_1, s6_v);
  spice_node_2 n_s5(eclk, ereset, s5_port_0,s5_port_1, s5_v);
  spice_node_2 n_s4(eclk, ereset, s4_port_0,s4_port_1, s4_v);
  spice_node_2 n_so(eclk, ereset, so_port_2,so_port_3, so_v);
  spice_node_2 n_dpc15_ANDS(eclk, ereset, dpc15_ANDS_port_9,dpc15_ANDS_port_0, dpc15_ANDS_v);
  spice_node_2 n_dpc27_SBADH(eclk, ereset, dpc27_SBADH_port_9,dpc27_SBADH_port_0, dpc27_SBADH_v);
  spice_node_3 n_n_649(eclk, ereset, n_649_port_0,n_649_port_7,n_649_port_5, n_649_v);
  spice_node_3 n_n_138(eclk, ereset, n_138_port_2,n_138_port_0,n_138_port_1, n_138_v);
  spice_node_3 n_n_642(eclk, ereset, n_642_port_3,n_642_port_0,n_642_port_1, n_642_v);
  spice_node_2 n_n_643(eclk, ereset, n_643_port_3,n_643_port_4, n_643_v);
  spice_node_3 n_n_1632(eclk, ereset, n_1632_port_7,n_1632_port_4,n_1632_port_5, n_1632_v);
  spice_node_3 n_n_583(eclk, ereset, n_583_port_2,n_583_port_0,n_583_port_1, n_583_v);
  spice_node_3 n_notir0(eclk, ereset, notir0_port_0,notir0_port_1,notir0_port_28, notir0_v);
  spice_node_3 n_notir1(eclk, ereset, notir1_port_21,notir1_port_23,notir1_port_22, notir1_v);
  spice_node_3 n_notir2(eclk, ereset, notir2_port_19,notir2_port_0,notir2_port_20, notir2_v);
  spice_node_3 n_notir3(eclk, ereset, notir3_port_51,notir3_port_0,notir3_port_1, notir3_v);
  spice_node_3 n_notir4(eclk, ereset, notir4_port_25,notir4_port_24,notir4_port_26, notir4_v);
  spice_node_3 n_notir5(eclk, ereset, notir5_port_36,notir5_port_37,notir5_port_0, notir5_v);
  spice_node_3 n_notir6(eclk, ereset, notir6_port_39,notir6_port_0,notir6_port_1, notir6_v);
  spice_node_3 n_notir7(eclk, ereset, notir7_port_33,notir7_port_34,notir7_port_35, notir7_v);
  spice_node_2 n_n_119(eclk, ereset, n_119_port_3,n_119_port_0, n_119_v);
  spice_node_2 n_cp1(eclk, ereset, cp1_port_75,cp1_port_50, cp1_v);
  spice_node_2 n_a3(eclk, ereset, a3_port_0,a3_port_1, a3_v);
  spice_node_2 n_a6(eclk, ereset, a6_port_2,a6_port_0, a6_v);
  spice_node_2 n_n_1479(eclk, ereset, n_1479_port_0,n_1479_port_1, n_1479_v);
  spice_node_2 n_sync(eclk, ereset, sync_port_0,sync_port_1, sync_v);
  spice_node_2 n_n_1325(eclk, ereset, n_1325_port_2,n_1325_port_4, n_1325_v);
  spice_node_5 n_n_1496(eclk, ereset, n_1496_port_2,n_1496_port_3,n_1496_port_0,n_1496_port_1,n_1496_port_4, n_1496_v);
  spice_node_4 n_n_564(eclk, ereset, n_564_port_2,n_564_port_3,n_564_port_0,n_564_port_1, n_564_v);
  spice_node_3 n___AxBxC_6(eclk, ereset, __AxBxC_6_port_3,__AxBxC_6_port_1,__AxBxC_6_port_5, __AxBxC_6_v);
  spice_node_3 n___AxBxC_7(eclk, ereset, __AxBxC_7_port_3,__AxBxC_7_port_0,__AxBxC_7_port_5, __AxBxC_7_v);
  spice_node_3 n___AxBxC_4(eclk, ereset, __AxBxC_4_port_2,__AxBxC_4_port_3,__AxBxC_4_port_5, __AxBxC_4_v);
  spice_node_3 n___AxBxC_5(eclk, ereset, __AxBxC_5_port_3,__AxBxC_5_port_1,__AxBxC_5_port_5, __AxBxC_5_v);
  spice_node_3 n___AxBxC_2(eclk, ereset, __AxBxC_2_port_3,__AxBxC_2_port_1,__AxBxC_2_port_5, __AxBxC_2_v);
  spice_node_3 n___AxBxC_3(eclk, ereset, __AxBxC_3_port_3,__AxBxC_3_port_1,__AxBxC_3_port_5, __AxBxC_3_v);
  spice_node_3 n___AxBxC_0(eclk, ereset, __AxBxC_0_port_2,__AxBxC_0_port_3,__AxBxC_0_port_5, __AxBxC_0_v);
  spice_node_3 n___AxBxC_1(eclk, ereset, __AxBxC_1_port_3,__AxBxC_1_port_1,__AxBxC_1_port_5, __AxBxC_1_v);
  spice_node_5 n_n_304(eclk, ereset, n_304_port_2,n_304_port_3,n_304_port_0,n_304_port_1,n_304_port_4, n_304_v);
  spice_node_2 n_ab12(eclk, ereset, ab12_port_0,ab12_port_1, ab12_v);
  spice_node_2 n_ab13(eclk, ereset, ab13_port_0,ab13_port_1, ab13_v);
  spice_node_2 n_ab10(eclk, ereset, ab10_port_0,ab10_port_1, ab10_v);
  spice_node_2 n_ab11(eclk, ereset, ab11_port_0,ab11_port_1, ab11_v);
  spice_node_2 n_ab14(eclk, ereset, ab14_port_0,ab14_port_1, ab14_v);
  spice_node_2 n_ab15(eclk, ereset, ab15_port_0,ab15_port_1, ab15_v);
  spice_node_5 n_n_72(eclk, ereset, n_72_port_2,n_72_port_3,n_72_port_0,n_72_port_1,n_72_port_4, n_72_v);
  spice_node_3 n_n_177(eclk, ereset, n_177_port_2,n_177_port_0,n_177_port_1, n_177_v);
  spice_node_2 n_n_794(eclk, ereset, n_794_port_1,n_794_port_4, n_794_v);
  spice_node_2 n_n_798(eclk, ereset, n_798_port_1,n_798_port_4, n_798_v);
  spice_node_5 n_n_1301(eclk, ereset, n_1301_port_2,n_1301_port_3,n_1301_port_0,n_1301_port_1,n_1301_port_4, n_1301_v);
  spice_node_2 n_n_1300(eclk, ereset, n_1300_port_2,n_1300_port_3, n_1300_v);
  spice_node_3 n_n_1309(eclk, ereset, n_1309_port_2,n_1309_port_3,n_1309_port_1, n_1309_v);
  spice_node_2 n_n_330(eclk, ereset, n_330_port_7,n_330_port_4, n_330_v);
  spice_node_5 n_n_332(eclk, ereset, n_332_port_2,n_332_port_3,n_332_port_0,n_332_port_1,n_332_port_4, n_332_v);
  spice_node_4 n_n_1169(eclk, ereset, n_1169_port_2,n_1169_port_3,n_1169_port_0,n_1169_port_1, n_1169_v);
  spice_node_2 n_n_541(eclk, ereset, n_541_port_3,n_541_port_1, n_541_v);
  spice_node_2 n_n_322(eclk, ereset, n_322_port_2,n_322_port_1, n_322_v);
  spice_node_2 n_dpc24_ACSB(eclk, ereset, dpc24_ACSB_port_1,dpc24_ACSB_port_12, dpc24_ACSB_v);
  spice_node_2 n_rdy(eclk, ereset, rdy_port_2,rdy_port_3, rdy_v);
  spice_node_2 n_n_520(eclk, ereset, n_520_port_0,n_520_port_4, n_520_v);
  spice_node_2 n_dpc21_ADDADL(eclk, ereset, dpc21_ADDADL_port_9,dpc21_ADDADL_port_0, dpc21_ADDADL_v);
  spice_node_5 n_n_1592(eclk, ereset, n_1592_port_2,n_1592_port_3,n_1592_port_0,n_1592_port_1,n_1592_port_4, n_1592_v);
  spice_node_2 n_n_37(eclk, ereset, n_37_port_3,n_37_port_4, n_37_v);
  spice_node_3 n_db1(eclk, ereset, db1_port_1,db1_port_4,db1_port_5, db1_v);
  spice_node_3 n_db0(eclk, ereset, db0_port_1,db0_port_4,db0_port_5, db0_v);
  spice_node_3 n_db3(eclk, ereset, db3_port_2,db3_port_3,db3_port_5, db3_v);
  spice_node_3 n_db2(eclk, ereset, db2_port_2,db2_port_3,db2_port_5, db2_v);
  spice_node_3 n_db5(eclk, ereset, db5_port_0,db5_port_4,db5_port_5, db5_v);
  spice_node_3 n_db4(eclk, ereset, db4_port_3,db4_port_0,db4_port_5, db4_v);
  spice_node_3 n_db7(eclk, ereset, db7_port_3,db7_port_1,db7_port_5, db7_v);
  spice_node_3 n_db6(eclk, ereset, db6_port_0,db6_port_4,db6_port_5, db6_v);
  spice_node_2 n_clk1out(eclk, ereset, clk1out_port_0,clk1out_port_1, clk1out_v);
  spice_node_5 n_n_1647(eclk, ereset, n_1647_port_2,n_1647_port_3,n_1647_port_0,n_1647_port_1,n_1647_port_4, n_1647_v);
  spice_node_3 n_n_1641(eclk, ereset, n_1641_port_2,n_1641_port_3,n_1641_port_1, n_1641_v);
  spice_node_4 n_n_1491(eclk, ereset, n_1491_port_2,n_1491_port_3,n_1491_port_0,n_1491_port_1, n_1491_v);
  spice_node_3 n_n_206(eclk, ereset, n_206_port_3,n_206_port_0,n_206_port_5, n_206_v);
  spice_node_2 n_clock1(eclk, ereset, clock1_port_40,clock1_port_68, clock1_v);
  spice_node_5 n_n_1344(eclk, ereset, n_1344_port_2,n_1344_port_3,n_1344_port_0,n_1344_port_1,n_1344_port_4, n_1344_v);
  spice_node_3 n_n_1084(eclk, ereset, n_1084_port_0,n_1084_port_6,n_1084_port_5, n_1084_v);
  spice_node_3 n_n_1083(eclk, ereset, n_1083_port_1,n_1083_port_7,n_1083_port_4, n_1083_v);
  spice_node_4 n_n_1661(eclk, ereset, n_1661_port_2,n_1661_port_3,n_1661_port_0,n_1661_port_1, n_1661_v);
  spice_node_3 n_n_1668(eclk, ereset, n_1668_port_2,n_1668_port_3,n_1668_port_0, n_1668_v);
  spice_node_2 n_dpc32_PCHADH(eclk, ereset, dpc32_PCHADH_port_0,dpc32_PCHADH_port_1, dpc32_PCHADH_v);
  spice_node_8 n_idb1(eclk, ereset, idb1_port_8,idb1_port_9,idb1_port_3,idb1_port_0,idb1_port_7,idb1_port_4,idb1_port_5,idb1_port_10, idb1_v);
  spice_node_8 n_idb0(eclk, ereset, idb0_port_8,idb0_port_2,idb0_port_1,idb0_port_6,idb0_port_7,idb0_port_4,idb0_port_5,idb0_port_10, idb0_v);
  spice_node_8 n_idb3(eclk, ereset, idb3_port_8,idb3_port_9,idb3_port_3,idb3_port_0,idb3_port_1,idb3_port_6,idb3_port_5,idb3_port_10, idb3_v);
  spice_node_8 n_idb2(eclk, ereset, idb2_port_9,idb2_port_3,idb2_port_0,idb2_port_1,idb2_port_6,idb2_port_4,idb2_port_5,idb2_port_10, idb2_v);
  spice_node_7 n_idb5(eclk, ereset, idb5_port_8,idb5_port_9,idb5_port_2,idb5_port_6,idb5_port_7,idb5_port_4,idb5_port_5, idb5_v);
  spice_node_8 n_idb4(eclk, ereset, idb4_port_8,idb4_port_9,idb4_port_0,idb4_port_6,idb4_port_7,idb4_port_4,idb4_port_5,idb4_port_10, idb4_v);
  spice_node_8 n_idb7(eclk, ereset, idb7_port_8,idb7_port_9,idb7_port_2,idb7_port_3,idb7_port_0,idb7_port_7,idb7_port_4,idb7_port_10, idb7_v);
  spice_node_8 n_idb6(eclk, ereset, idb6_port_9,idb6_port_3,idb6_port_0,idb6_port_6,idb6_port_7,idb6_port_5,idb6_port_10,idb6_port_11, idb6_v);
  spice_node_2 n_n_1417(eclk, ereset, n_1417_port_2,n_1417_port_0, n_1417_v);
  spice_node_3 n_n_381(eclk, ereset, n_381_port_2,n_381_port_3,n_381_port_1, n_381_v);
  spice_node_2 n_n_927(eclk, ereset, n_927_port_3,n_927_port_1, n_927_v);
  spice_node_3 n_n_928(eclk, ereset, n_928_port_2,n_928_port_3,n_928_port_1, n_928_v);
  spice_node_3 n_alub2(eclk, ereset, alub2_port_0,alub2_port_1,alub2_port_4, alub2_v);
  spice_node_2 n_pch7(eclk, ereset, pch7_port_2,pch7_port_1, pch7_v);
  spice_node_2 n_pch6(eclk, ereset, pch6_port_2,pch6_port_0, pch6_v);
  spice_node_2 n_pch5(eclk, ereset, pch5_port_2,pch5_port_0, pch5_v);
  spice_node_2 n_pch4(eclk, ereset, pch4_port_2,pch4_port_1, pch4_v);
  spice_node_2 n_pch3(eclk, ereset, pch3_port_2,pch3_port_1, pch3_v);
  spice_node_2 n_pch2(eclk, ereset, pch2_port_0,pch2_port_1, pch2_v);
  spice_node_2 n_pch1(eclk, ereset, pch1_port_2,pch1_port_1, pch1_v);
  spice_node_2 n_pch0(eclk, ereset, pch0_port_2,pch0_port_1, pch0_v);
  spice_node_2 n_dpc13_ORS(eclk, ereset, dpc13_ORS_port_8,dpc13_ORS_port_5, dpc13_ORS_v);
  spice_node_4 n_n_1063(eclk, ereset, n_1063_port_2,n_1063_port_7,n_1063_port_4,n_1063_port_5, n_1063_v);
  spice_node_2 n_n_1608(eclk, ereset, n_1608_port_2,n_1608_port_1, n_1608_v);
  spice_node_2 n_n_1609(eclk, ereset, n_1609_port_3,n_1609_port_0, n_1609_v);
  spice_node_3 n_n_1605(eclk, ereset, n_1605_port_3,n_1605_port_0,n_1605_port_5, n_1605_v);
  spice_node_4 n_n_719(eclk, ereset, n_719_port_2,n_719_port_3,n_719_port_0,n_719_port_1, n_719_v);
  spice_node_4 n_n_242(eclk, ereset, n_242_port_2,n_242_port_3,n_242_port_0,n_242_port_1, n_242_v);
  spice_node_3 n_dasb7(eclk, ereset, dasb7_port_3,dasb7_port_1,dasb7_port_5, dasb7_v);
  spice_node_2 n_n_1296(eclk, ereset, n_1296_port_2,n_1296_port_0, n_1296_v);
  spice_node_2 n_dpc7_SS(eclk, ereset, dpc7_SS_port_7,dpc7_SS_port_12, dpc7_SS_v);
  spice_node_2 n_n_1041(eclk, ereset, n_1041_port_0,n_1041_port_1, n_1041_v);
  spice_node_3 n_n_1046(eclk, ereset, n_1046_port_2,n_1046_port_3,n_1046_port_0, n_1046_v);
  spice_node_2 n_n_1620(eclk, ereset, n_1620_port_3,n_1620_port_0, n_1620_v);
  spice_node_3 n_n_1621(eclk, ereset, n_1621_port_2,n_1621_port_0,n_1621_port_1, n_1621_v);
  spice_node_3 n_n_227(eclk, ereset, n_227_port_2,n_227_port_3,n_227_port_0, n_227_v);
  spice_node_2 n_x2(eclk, ereset, x2_port_0,x2_port_1, x2_v);
  spice_node_2 n_x3(eclk, ereset, x3_port_0,x3_port_1, x3_v);
  spice_node_2 n_x0(eclk, ereset, x0_port_0,x0_port_1, x0_v);
  spice_node_2 n_x1(eclk, ereset, x1_port_0,x1_port_1, x1_v);
  spice_node_2 n_x7(eclk, ereset, x7_port_2,x7_port_1, x7_v);
  spice_node_2 n_x4(eclk, ereset, x4_port_0,x4_port_1, x4_v);
  spice_node_2 n_x5(eclk, ereset, x5_port_2,x5_port_1, x5_v);
  spice_node_5 n_n_1458(eclk, ereset, n_1458_port_2,n_1458_port_3,n_1458_port_0,n_1458_port_1,n_1458_port_4, n_1458_v);
  spice_node_5 n_n_694(eclk, ereset, n_694_port_2,n_694_port_3,n_694_port_0,n_694_port_1,n_694_port_4, n_694_v);
  spice_node_2 n_n_963(eclk, ereset, n_963_port_2,n_963_port_1, n_963_v);
  spice_node_2 n_pcl3(eclk, ereset, pcl3_port_2,pcl3_port_1, pcl3_v);
  spice_node_2 n_pcl2(eclk, ereset, pcl2_port_2,pcl2_port_1, pcl2_v);
  spice_node_2 n_pcl1(eclk, ereset, pcl1_port_2,pcl1_port_1, pcl1_v);
  spice_node_2 n_pcl0(eclk, ereset, pcl0_port_2,pcl0_port_1, pcl0_v);
  spice_node_2 n_pcl7(eclk, ereset, pcl7_port_2,pcl7_port_1, pcl7_v);
  spice_node_2 n_pcl6(eclk, ereset, pcl6_port_2,pcl6_port_1, pcl6_v);
  spice_node_2 n_pcl5(eclk, ereset, pcl5_port_2,pcl5_port_1, pcl5_v);
  spice_node_2 n_pcl4(eclk, ereset, pcl4_port_2,pcl4_port_1, pcl4_v);
  spice_node_2 n_dpc0_YSB(eclk, ereset, dpc0_YSB_port_3,dpc0_YSB_port_12, dpc0_YSB_v);
  spice_node_2 n_alua6(eclk, ereset, alua6_port_0,alua6_port_1, alua6_v);
  spice_node_2 n_alua7(eclk, ereset, alua7_port_3,alua7_port_0, alua7_v);
  spice_node_2 n_alua4(eclk, ereset, alua4_port_0,alua4_port_1, alua4_v);
  spice_node_2 n_alua5(eclk, ereset, alua5_port_0,alua5_port_1, alua5_v);
  spice_node_2 n_alua2(eclk, ereset, alua2_port_0,alua2_port_1, alua2_v);
  spice_node_2 n_alua3(eclk, ereset, alua3_port_0,alua3_port_1, alua3_v);
  spice_node_2 n_alua0(eclk, ereset, alua0_port_0,alua0_port_1, alua0_v);
  spice_node_2 n_alua1(eclk, ereset, alua1_port_2,alua1_port_3, alua1_v);
  spice_node_1 n_nmi(eclk, ereset, nmi_port_2, nmi_v);
  spice_node_2 n_dpc41_DL_ADL(eclk, ereset, dpc41_DL_ADL_port_9,dpc41_DL_ADL_port_0, dpc41_DL_ADL_v);
  spice_node_5 n_n_208(eclk, ereset, n_208_port_2,n_208_port_3,n_208_port_0,n_208_port_1,n_208_port_4, n_208_v);
  spice_node_5 n_n_209(eclk, ereset, n_209_port_2,n_209_port_3,n_209_port_0,n_209_port_1,n_209_port_4, n_209_v);
  spice_node_2 n_dpc37_PCLDB(eclk, ereset, dpc37_PCLDB_port_0,dpc37_PCLDB_port_4, dpc37_PCLDB_v);
  spice_node_2 n_dpc12_0ADD(eclk, ereset, dpc12_0ADD_port_9,dpc12_0ADD_port_12, dpc12_0ADD_v);
  spice_node_2 n_dpc4_SSB(eclk, ereset, dpc4_SSB_port_9,dpc4_SSB_port_0, dpc4_SSB_v);
  spice_node_2 n_n_417(eclk, ereset, n_417_port_0,n_417_port_1, n_417_v);
  spice_node_2 n_y1(eclk, ereset, y1_port_2,y1_port_0, y1_v);
  spice_node_2 n_y0(eclk, ereset, y0_port_2,y0_port_0, y0_v);
  spice_node_2 n_y3(eclk, ereset, y3_port_2,y3_port_0, y3_v);
  spice_node_2 n_y2(eclk, ereset, y2_port_2,y2_port_0, y2_v);
  spice_node_2 n_y5(eclk, ereset, y5_port_0,y5_port_1, y5_v);
  spice_node_2 n_y4(eclk, ereset, y4_port_2,y4_port_0, y4_v);
  spice_node_2 n_y7(eclk, ereset, y7_port_0,y7_port_1, y7_v);
  spice_node_2 n_y6(eclk, ereset, y6_port_0,y6_port_1, y6_v);
  spice_node_2 n_dpc11_SBADD(eclk, ereset, dpc11_SBADD_port_9,dpc11_SBADD_port_12, dpc11_SBADD_v);
  spice_node_2 n_dpc10_ADLADD(eclk, ereset, dpc10_ADLADD_port_5,dpc10_ADLADD_port_12, dpc10_ADLADD_v);
  spice_node_2 n_dpc29_0ADH17(eclk, ereset, dpc29_0ADH17_port_2,dpc29_0ADH17_port_1, dpc29_0ADH17_v);
  spice_node_2 n_dpc26_ACDB(eclk, ereset, dpc26_ACDB_port_0,dpc26_ACDB_port_12, dpc26_ACDB_v);
  spice_node_3 n_n_430(eclk, ereset, n_430_port_2,n_430_port_3,n_430_port_1, n_430_v);
  spice_node_4 n_n_436(eclk, ereset, n_436_port_2,n_436_port_3,n_436_port_0,n_436_port_1, n_436_v);
  spice_node_3 n_n_404(eclk, ereset, n_404_port_2,n_404_port_6,n_404_port_5, n_404_v);
  spice_node_5 n_n_1654(eclk, ereset, n_1654_port_2,n_1654_port_3,n_1654_port_0,n_1654_port_1,n_1654_port_4, n_1654_v);
  spice_node_3 n_n_635(eclk, ereset, n_635_port_3,n_635_port_0,n_635_port_1, n_635_v);
  spice_node_2 n_n_634(eclk, ereset, n_634_port_0,n_634_port_1, n_634_v);
  spice_node_1 n_n_633(eclk, ereset, n_633_port_0, n_633_v);
  spice_node_3 n_n_458(eclk, ereset, n_458_port_2,n_458_port_0,n_458_port_1, n_458_v);
  spice_node_3 n_n_1519(eclk, ereset, n_1519_port_2,n_1519_port_3,n_1519_port_0, n_1519_v);
  spice_node_2 n_dpc16_EORS(eclk, ereset, dpc16_EORS_port_8,dpc16_EORS_port_9, dpc16_EORS_v);
  spice_node_5 n_n_1722(eclk, ereset, n_1722_port_2,n_1722_port_3,n_1722_port_0,n_1722_port_1,n_1722_port_4, n_1722_v);
  spice_node_5 n_n_618(eclk, ereset, n_618_port_2,n_618_port_3,n_618_port_0,n_618_port_1,n_618_port_4, n_618_v);
  spice_node_2 n_n_612(eclk, ereset, n_612_port_0,n_612_port_4, n_612_v);
  spice_node_3 n_n_884(eclk, ereset, n_884_port_2,n_884_port_0,n_884_port_1, n_884_v);
  spice_node_3 n_Pout0(eclk, ereset, Pout0_port_2,Pout0_port_0,Pout0_port_1, Pout0_v);
  spice_node_2 n_n_1545(eclk, ereset, n_1545_port_2,n_1545_port_1, n_1545_v);
  spice_node_2 n_dpc19_ADDSB7(eclk, ereset, dpc19_ADDSB7_port_2,dpc19_ADDSB7_port_0, dpc19_ADDSB7_v);
  spice_node_4 n_n_477(eclk, ereset, n_477_port_3,n_477_port_1,n_477_port_4,n_477_port_5, n_477_v);
  spice_node_2 n_n_475(eclk, ereset, n_475_port_2,n_475_port_0, n_475_v);
  spice_node_2 n_n_471(eclk, ereset, n_471_port_3,n_471_port_4, n_471_v);
  spice_node_3 n_n_478(eclk, ereset, n_478_port_2,n_478_port_0,n_478_port_1, n_478_v);
  spice_node_3 n_p6(eclk, ereset, p6_port_2,p6_port_0,p6_port_1, p6_v);
  spice_node_3 n_p7(eclk, ereset, p7_port_2,p7_port_0,p7_port_1, p7_v);
  spice_node_4 n_n_1531(eclk, ereset, n_1531_port_2,n_1531_port_3,n_1531_port_0,n_1531_port_1, n_1531_v);
  spice_node_3 n_n_1398(eclk, ereset, n_1398_port_8,n_1398_port_1,n_1398_port_6, n_1398_v);
  spice_node_5 n_n_280(eclk, ereset, n_280_port_2,n_280_port_3,n_280_port_0,n_280_port_1,n_280_port_4, n_280_v);
  spice_node_2 n_n_135(eclk, ereset, n_135_port_2,n_135_port_1, n_135_v);
  spice_node_3 n_n_869(eclk, ereset, n_869_port_2,n_869_port_3,n_869_port_1, n_869_v);
  spice_node_0 n_n_866(eclk, ereset,  n_866_v);
  spice_node_4 n_n_350(eclk, ereset, n_350_port_3,n_350_port_1,n_350_port_4,n_350_port_5, n_350_v);
  spice_node_2 n_dpc17_SUMS(eclk, ereset, dpc17_SUMS_port_0,dpc17_SUMS_port_1, dpc17_SUMS_v);
  spice_node_4 n_n_1251(eclk, ereset, n_1251_port_2,n_1251_port_3,n_1251_port_0,n_1251_port_1, n_1251_v);
  spice_node_4 n_n_1709(eclk, ereset, n_1709_port_2,n_1709_port_3,n_1709_port_0,n_1709_port_1, n_1709_v);
  spice_node_2 n_dpc3_SBX(eclk, ereset, dpc3_SBX_port_9,dpc3_SBX_port_12, dpc3_SBX_v);
  spice_node_2 n_dpc31_PCHPCH(eclk, ereset, dpc31_PCHPCH_port_11,dpc31_PCHPCH_port_12, dpc31_PCHPCH_v);
  spice_node_3 n_n_676(eclk, ereset, n_676_port_2,n_676_port_3,n_676_port_0, n_676_v);
  spice_node_3 n_Pout1(eclk, ereset, Pout1_port_2,Pout1_port_0,Pout1_port_1, Pout1_v);
  spice_node_3 n_Pout3(eclk, ereset, Pout3_port_2,Pout3_port_3,Pout3_port_4, Pout3_v);
  spice_node_3 n_Pout2(eclk, ereset, Pout2_port_2,Pout2_port_0,Pout2_port_1, Pout2_v);
  spice_node_3 n_n_494(eclk, ereset, n_494_port_2,n_494_port_3,n_494_port_1, n_494_v);
  spice_node_0 n_n_806(eclk, ereset,  n_806_v);
  spice_node_2 n_n_807(eclk, ereset, n_807_port_3,n_807_port_5, n_807_v);
  spice_node_3 n_n_659(eclk, ereset, n_659_port_2,n_659_port_3,n_659_port_1, n_659_v);
  spice_node_4 n_n_658(eclk, ereset, n_658_port_2,n_658_port_3,n_658_port_0,n_658_port_1, n_658_v);
  spice_node_5 n_n_652(eclk, ereset, n_652_port_2,n_652_port_3,n_652_port_0,n_652_port_1,n_652_port_4, n_652_v);
  spice_node_3 n_n_123(eclk, ereset, n_123_port_2,n_123_port_3,n_123_port_0, n_123_v);
  spice_node_2 n_n_826(eclk, ereset, n_826_port_2,n_826_port_1, n_826_v);
  spice_node_3 n_n_351(eclk, ereset, n_351_port_2,n_351_port_0,n_351_port_1, n_351_v);
  spice_node_2 n_dpc9_DBADD(eclk, ereset, dpc9_DBADD_port_1,dpc9_DBADD_port_12, dpc9_DBADD_v);
  spice_node_3 n_n_359(eclk, ereset, n_359_port_2,n_359_port_0,n_359_port_1, n_359_v);
  spice_node_2 n_dpc33_PCHDB(eclk, ereset, dpc33_PCHDB_port_0,dpc33_PCHDB_port_1, dpc33_PCHDB_v);
  spice_node_2 n_dpc8_nDBADD(eclk, ereset, dpc8_nDBADD_port_6,dpc8_nDBADD_port_12, dpc8_nDBADD_v);
  spice_node_2 n_n_102(eclk, ereset, n_102_port_2,n_102_port_0, n_102_v);
  spice_node_2 n_dpc39_PCLPCL(eclk, ereset, dpc39_PCLPCL_port_11,dpc39_PCLPCL_port_12, dpc39_PCLPCL_v);
  spice_node_2 n_ADH_ABH(eclk, ereset, ADH_ABH_port_7,ADH_ABH_port_4, ADH_ABH_v);
  spice_node_2 n_dpc25_SBDB(eclk, ereset, dpc25_SBDB_port_9,dpc25_SBDB_port_0, dpc25_SBDB_v);
  spice_node_2 n_dpc23_SBAC(eclk, ereset, dpc23_SBAC_port_11,dpc23_SBAC_port_12, dpc23_SBAC_v);
  spice_node_2 n_n_1152(eclk, ereset, n_1152_port_2,n_1152_port_0, n_1152_v);
  spice_node_2 n_n_373(eclk, ereset, n_373_port_0,n_373_port_4, n_373_v);
  spice_node_2 n_ab0(eclk, ereset, ab0_port_0,ab0_port_1, ab0_v);
  spice_node_2 n_ab1(eclk, ereset, ab1_port_0,ab1_port_1, ab1_v);
  spice_node_2 n_ab2(eclk, ereset, ab2_port_0,ab2_port_1, ab2_v);
  spice_node_2 n_ab3(eclk, ereset, ab3_port_0,ab3_port_1, ab3_v);
  spice_node_2 n_ab4(eclk, ereset, ab4_port_0,ab4_port_1, ab4_v);
  spice_node_2 n_ab5(eclk, ereset, ab5_port_0,ab5_port_1, ab5_v);
  spice_node_2 n_ab6(eclk, ereset, ab6_port_0,ab6_port_1, ab6_v);
  spice_node_2 n_ab7(eclk, ereset, ab7_port_0,ab7_port_1, ab7_v);
  spice_node_2 n_ab8(eclk, ereset, ab8_port_0,ab8_port_1, ab8_v);
  spice_node_2 n_ab9(eclk, ereset, ab9_port_0,ab9_port_1, ab9_v);
  spice_node_4 n_n_87(eclk, ereset, n_87_port_2,n_87_port_3,n_87_port_0,n_87_port_1, n_87_v);
  spice_node_3 n_n_86(eclk, ereset, n_86_port_2,n_86_port_3,n_86_port_0, n_86_v);
  spice_node_3 n_n_168(eclk, ereset, n_168_port_2,n_168_port_3,n_168_port_0, n_168_v);
  spice_node_12 n_sb2(eclk, ereset, sb2_port_8,sb2_port_9,sb2_port_2,sb2_port_3,sb2_port_0,sb2_port_1,sb2_port_6,sb2_port_7,sb2_port_4,sb2_port_10,sb2_port_11,sb2_port_12, sb2_v);
  spice_node_12 n_sb3(eclk, ereset, sb3_port_8,sb3_port_9,sb3_port_2,sb3_port_3,sb3_port_0,sb3_port_1,sb3_port_6,sb3_port_7,sb3_port_4,sb3_port_5,sb3_port_10,sb3_port_11, sb3_v);
  spice_node_13 n_sb0(eclk, ereset, sb0_port_8,sb0_port_9,sb0_port_2,sb0_port_3,sb0_port_0,sb0_port_1,sb0_port_6,sb0_port_7,sb0_port_4,sb0_port_5,sb0_port_10,sb0_port_11,sb0_port_12, sb0_v);
  spice_node_12 n_sb1(eclk, ereset, sb1_port_8,sb1_port_9,sb1_port_2,sb1_port_0,sb1_port_1,sb1_port_6,sb1_port_7,sb1_port_4,sb1_port_5,sb1_port_10,sb1_port_11,sb1_port_12, sb1_v);
  spice_node_12 n_sb6(eclk, ereset, sb6_port_8,sb6_port_9,sb6_port_2,sb6_port_3,sb6_port_0,sb6_port_1,sb6_port_6,sb6_port_7,sb6_port_4,sb6_port_10,sb6_port_11,sb6_port_12, sb6_v);
  spice_node_12 n_sb7(eclk, ereset, sb7_port_8,sb7_port_9,sb7_port_2,sb7_port_3,sb7_port_0,sb7_port_1,sb7_port_6,sb7_port_7,sb7_port_4,sb7_port_5,sb7_port_10,sb7_port_11, sb7_v);
  spice_node_13 n_sb4(eclk, ereset, sb4_port_8,sb4_port_9,sb4_port_2,sb4_port_3,sb4_port_0,sb4_port_1,sb4_port_6,sb4_port_7,sb4_port_4,sb4_port_5,sb4_port_10,sb4_port_11,sb4_port_12, sb4_v);
  spice_node_12 n_sb5(eclk, ereset, sb5_port_8,sb5_port_2,sb5_port_3,sb5_port_0,sb5_port_1,sb5_port_6,sb5_port_7,sb5_port_4,sb5_port_5,sb5_port_10,sb5_port_11,sb5_port_12, sb5_v);
  spice_node_3 n___AxB_6(eclk, ereset, __AxB_6_port_2,__AxB_6_port_6,__AxB_6_port_11, __AxB_6_v);
  spice_node_3 n___AxB_4(eclk, ereset, __AxB_4_port_0,__AxB_4_port_6,__AxB_4_port_4, __AxB_4_v);
  spice_node_3 n___AxB_2(eclk, ereset, __AxB_2_port_0,__AxB_2_port_7,__AxB_2_port_4, __AxB_2_v);
  spice_node_3 n___AxB_0(eclk, ereset, __AxB_0_port_2,__AxB_0_port_6,__AxB_0_port_4, __AxB_0_v);
  spice_node_4 n_n_1318(eclk, ereset, n_1318_port_2,n_1318_port_3,n_1318_port_7,n_1318_port_5, n_1318_v);
  spice_node_2 n_dpc2_XSB(eclk, ereset, dpc2_XSB_port_2,dpc2_XSB_port_12, dpc2_XSB_v);
  spice_node_4 n_n_578(eclk, ereset, n_578_port_2,n_578_port_3,n_578_port_0,n_578_port_1, n_578_v);
  spice_node_3 n_n_571(eclk, ereset, n_571_port_2,n_571_port_3,n_571_port_1, n_571_v);
  spice_node_2 n_n_310(eclk, ereset, n_310_port_3,n_310_port_0, n_310_v);
  spice_node_2 n_dpc14_SRS(eclk, ereset, dpc14_SRS_port_2,dpc14_SRS_port_1, dpc14_SRS_v);
  spice_node_3 n_n_66(eclk, ereset, n_66_port_2,n_66_port_3,n_66_port_1, n_66_v);
  spice_node_2 n_n_147(eclk, ereset, n_147_port_3,n_147_port_4, n_147_v);
  spice_node_5 n_n_146(eclk, ereset, n_146_port_2,n_146_port_3,n_146_port_0,n_146_port_1,n_146_port_4, n_146_v);
  spice_node_5 n_n_141(eclk, ereset, n_141_port_2,n_141_port_3,n_141_port_0,n_141_port_1,n_141_port_4, n_141_v);
  spice_node_2 n_ADL_ABL(eclk, ereset, ADL_ABL_port_0,ADL_ABL_port_5, ADL_ABL_v);
  spice_node_4 n_n_1724(eclk, ereset, n_1724_port_2,n_1724_port_3,n_1724_port_0,n_1724_port_1, n_1724_v);
  spice_node_2 n_n_1191(eclk, ereset, n_1191_port_2,n_1191_port_0, n_1191_v);
  spice_node_3 n_n_883(eclk, ereset, n_883_port_2,n_883_port_3,n_883_port_1, n_883_v);
  spice_node_3 n_n_880(eclk, ereset, n_880_port_2,n_880_port_3,n_880_port_0, n_880_v);
  spice_node_4 n_n_336(eclk, ereset, n_336_port_3,n_336_port_1,n_336_port_6,n_336_port_7, n_336_v);
  spice_node_2 n_n_43(eclk, ereset, n_43_port_11,n_43_port_13, n_43_v);
  spice_node_2 n_n_42(eclk, ereset, n_42_port_0,n_42_port_4, n_42_v);
  spice_node_1 n_res(eclk, ereset, res_port_2, res_v);
  spice_node_7 n_adl7(eclk, ereset, adl7_port_2,adl7_port_3,adl7_port_0,adl7_port_6,adl7_port_7,adl7_port_4,adl7_port_5, adl7_v);
  spice_node_7 n_adl6(eclk, ereset, adl6_port_2,adl6_port_3,adl6_port_1,adl6_port_6,adl6_port_7,adl6_port_4,adl6_port_5, adl6_v);
  spice_node_7 n_adl5(eclk, ereset, adl5_port_2,adl5_port_3,adl5_port_0,adl5_port_1,adl5_port_7,adl5_port_4,adl5_port_5, adl5_v);
  spice_node_7 n_adl4(eclk, ereset, adl4_port_3,adl4_port_0,adl4_port_1,adl4_port_6,adl4_port_7,adl4_port_4,adl4_port_5, adl4_v);
  spice_node_7 n_adl3(eclk, ereset, adl3_port_2,adl3_port_3,adl3_port_0,adl3_port_1,adl3_port_6,adl3_port_7,adl3_port_4, adl3_v);
  spice_node_8 n_adl2(eclk, ereset, adl2_port_8,adl2_port_2,adl2_port_3,adl2_port_0,adl2_port_1,adl2_port_6,adl2_port_4,adl2_port_5, adl2_v);
  spice_node_8 n_adl1(eclk, ereset, adl1_port_8,adl1_port_2,adl1_port_3,adl1_port_0,adl1_port_1,adl1_port_7,adl1_port_4,adl1_port_5, adl1_v);
  spice_node_8 n_adl0(eclk, ereset, adl0_port_8,adl0_port_3,adl0_port_0,adl0_port_1,adl0_port_6,adl0_port_7,adl0_port_4,adl0_port_5, adl0_v);
  spice_node_4 n_n_1014(eclk, ereset, n_1014_port_2,n_1014_port_3,n_1014_port_0,n_1014_port_1, n_1014_v);
  spice_node_2 n_dpc40_ADLPCL(eclk, ereset, dpc40_ADLPCL_port_0,dpc40_ADLPCL_port_12, dpc40_ADLPCL_v);
  spice_node_5 n_n_929(eclk, ereset, n_929_port_2,n_929_port_3,n_929_port_0,n_929_port_1,n_929_port_4, n_929_v);
  spice_node_4 n_n_1424(eclk, ereset, n_1424_port_2,n_1424_port_3,n_1424_port_0,n_1424_port_1, n_1424_v);
  spice_node_5 n_notaluoutmux0(eclk, ereset, notaluoutmux0_port_2,notaluoutmux0_port_3,notaluoutmux0_port_0,notaluoutmux0_port_1,notaluoutmux0_port_5, notaluoutmux0_v);
  spice_node_5 n_notaluoutmux1(eclk, ereset, notaluoutmux1_port_2,notaluoutmux1_port_0,notaluoutmux1_port_1,notaluoutmux1_port_4,notaluoutmux1_port_5, notaluoutmux1_v);
  spice_node_2 n_dpc30_ADHPCH(eclk, ereset, dpc30_ADHPCH_port_10,dpc30_ADHPCH_port_12, dpc30_ADHPCH_v);
  spice_node_2 n_dpc43_DL_DB(eclk, ereset, dpc43_DL_DB_port_9,dpc43_DL_DB_port_0, dpc43_DL_DB_v);
  spice_node_5 n_n_27(eclk, ereset, n_27_port_2,n_27_port_3,n_27_port_0,n_27_port_1,n_27_port_4, n_27_v);
  spice_node_3 n_aluanorb0(eclk, ereset, aluanorb0_port_1,aluanorb0_port_6,aluanorb0_port_7, aluanorb0_v);
  spice_node_4 n_n_1694(eclk, ereset, n_1694_port_2,n_1694_port_3,n_1694_port_0,n_1694_port_1, n_1694_v);
  spice_node_2 n_a1(eclk, ereset, a1_port_0,a1_port_1, a1_v);
  spice_node_2 n_a0(eclk, ereset, a0_port_0,a0_port_1, a0_v);
  spice_node_2 n_a2(eclk, ereset, a2_port_2,a2_port_1, a2_v);
  spice_node_2 n_a5(eclk, ereset, a5_port_2,a5_port_0, a5_v);
  spice_node_2 n_a4(eclk, ereset, a4_port_2,a4_port_0, a4_v);
  spice_node_2 n_a7(eclk, ereset, a7_port_2,a7_port_1, a7_v);
  spice_node_5 n_n_277(eclk, ereset, n_277_port_2,n_277_port_3,n_277_port_1,n_277_port_4,n_277_port_5, n_277_v);
  spice_node_4 n_n_518(eclk, ereset, n_518_port_2,n_518_port_3,n_518_port_0,n_518_port_1, n_518_v);
  spice_node_2 n_n_1467(eclk, ereset, n_1467_port_0,n_1467_port_1, n_1467_v);
  spice_node_4 n_n_1095(eclk, ereset, n_1095_port_2,n_1095_port_3,n_1095_port_0,n_1095_port_1, n_1095_v);
  spice_node_3 n_n_1094(eclk, ereset, n_1094_port_2,n_1094_port_3,n_1094_port_1, n_1094_v);
  spice_node_2 n_n_1675(eclk, ereset, n_1675_port_3,n_1675_port_0, n_1675_v);
  spice_node_6 n_adh3(eclk, ereset, adh3_port_2,adh3_port_3,adh3_port_0,adh3_port_6,adh3_port_4,adh3_port_5, adh3_v);
  spice_node_6 n_adh2(eclk, ereset, adh2_port_3,adh2_port_0,adh2_port_1,adh2_port_6,adh2_port_4,adh2_port_5, adh2_v);
  spice_node_6 n_adh1(eclk, ereset, adh1_port_2,adh1_port_0,adh1_port_1,adh1_port_6,adh1_port_4,adh1_port_5, adh1_v);
  spice_node_6 n_adh0(eclk, ereset, adh0_port_2,adh0_port_3,adh0_port_0,adh0_port_1,adh0_port_6,adh0_port_4, adh0_v);
  spice_node_6 n_adh7(eclk, ereset, adh7_port_2,adh7_port_3,adh7_port_0,adh7_port_1,adh7_port_4,adh7_port_5, adh7_v);
  spice_node_6 n_adh6(eclk, ereset, adh6_port_3,adh6_port_0,adh6_port_1,adh6_port_6,adh6_port_4,adh6_port_5, adh6_v);
  spice_node_6 n_adh5(eclk, ereset, adh5_port_2,adh5_port_3,adh5_port_0,adh5_port_1,adh5_port_4,adh5_port_5, adh5_v);
  spice_node_6 n_adh4(eclk, ereset, adh4_port_2,adh4_port_0,adh4_port_1,adh4_port_6,adh4_port_4,adh4_port_5, adh4_v);
  spice_node_3 n_n_254(eclk, ereset, n_254_port_2,n_254_port_3,n_254_port_1, n_254_v);
  spice_node_3 n_n_1469(eclk, ereset, n_1469_port_2,n_1469_port_0,n_1469_port_1, n_1469_v);
  spice_node_3 n_n_935(eclk, ereset, n_935_port_2,n_935_port_3,n_935_port_1, n_935_v);
  spice_node_2 n_NMIP(eclk, ereset, NMIP_port_7,NMIP_port_4, NMIP_v);
  spice_node_2 n_n_1076(eclk, ereset, n_1076_port_0,n_1076_port_4, n_1076_v);
  spice_node_5 n_n_1071(eclk, ereset, n_1071_port_2,n_1071_port_3,n_1071_port_0,n_1071_port_4,n_1071_port_5, n_1071_v);
  spice_node_2 n_n_1072(eclk, ereset, n_1072_port_2,n_1072_port_4, n_1072_v);
  spice_node_2 n_n_1140(eclk, ereset, n_1140_port_2,n_1140_port_1, n_1140_v);
  spice_node_4 n_n_1147(eclk, ereset, n_1147_port_2,n_1147_port_3,n_1147_port_0,n_1147_port_1, n_1147_v);
  spice_node_3 n_aluanorb1(eclk, ereset, aluanorb1_port_7,aluanorb1_port_4,aluanorb1_port_5, aluanorb1_v);
  spice_node_5 n_n_723(eclk, ereset, n_723_port_2,n_723_port_3,n_723_port_0,n_723_port_1,n_723_port_4, n_723_v);
  spice_node_5 n_n_722(eclk, ereset, n_722_port_2,n_722_port_0,n_722_port_1,n_722_port_4,n_722_port_5, n_722_v);
  spice_node_5 n_n_721(eclk, ereset, n_721_port_2,n_721_port_3,n_721_port_0,n_721_port_1,n_721_port_4, n_721_v);
  spice_node_2 n_dpc1_SBY(eclk, ereset, dpc1_SBY_port_3,dpc1_SBY_port_12, dpc1_SBY_v);
  spice_node_2 n_cclk(eclk, ereset, cclk_port_236,cclk_port_28, cclk_v);
  spice_node_2 n_RnWstretched(eclk, ereset, RnWstretched_port_23,RnWstretched_port_22, RnWstretched_v);
  spice_node_1 n_n_1059(eclk, ereset, n_1059_port_0, n_1059_v);
  spice_node_2 n_n_1633(eclk, ereset, n_1633_port_2,n_1633_port_0, n_1633_v);
  spice_node_2 n_n_1639(eclk, ereset, n_1639_port_2,n_1639_port_0, n_1639_v);
  spice_node_5 n_n_740(eclk, ereset, n_740_port_2,n_740_port_3,n_740_port_0,n_740_port_1,n_740_port_4, n_740_v);
  spice_node_3 n_n_212(eclk, ereset, n_212_port_2,n_212_port_3,n_212_port_1, n_212_v);
  spice_node_3 n_n_210(eclk, ereset, n_210_port_3,n_210_port_0,n_210_port_1, n_210_v);
  spice_node_2 n_notRdy0(eclk, ereset, notRdy0_port_3,notRdy0_port_4, notRdy0_v);
  spice_node_3 n_n_624(eclk, ereset, n_624_port_2,n_624_port_0,n_624_port_1, n_624_v);
  spice_node_2 n_clk2out(eclk, ereset, clk2out_port_0,clk2out_port_1, clk2out_v);
  spice_node_4 n_n_681(eclk, ereset, n_681_port_8,n_681_port_3,n_681_port_1,n_681_port_6, n_681_v);
  spice_node_5 n_n_976(eclk, ereset, n_976_port_2,n_976_port_3,n_976_port_0,n_976_port_1,n_976_port_4, n_976_v);
  spice_node_2 n_n_975(eclk, ereset, n_975_port_3,n_975_port_6, n_975_v);
  spice_node_5 n_n_1618(eclk, ereset, n_1618_port_2,n_1618_port_3,n_1618_port_0,n_1618_port_1,n_1618_port_4, n_1618_v);
  spice_node_3 n_alub3(eclk, ereset, alub3_port_2,alub3_port_3,alub3_port_4, alub3_v);
  spice_node_3 n_alub1(eclk, ereset, alub1_port_0,alub1_port_1,alub1_port_4, alub1_v);
  spice_node_3 n_alub0(eclk, ereset, alub0_port_2,alub0_port_3,alub0_port_4, alub0_v);
  spice_node_3 n_alub7(eclk, ereset, alub7_port_3,alub7_port_0,alub7_port_4, alub7_v);
  spice_node_3 n_alub6(eclk, ereset, alub6_port_2,alub6_port_3,alub6_port_4, alub6_v);
  spice_node_3 n_alub5(eclk, ereset, alub5_port_2,alub5_port_3,alub5_port_4, alub5_v);
  spice_node_3 n_alub4(eclk, ereset, alub4_port_3,alub4_port_0,alub4_port_4, alub4_v);
  spice_node_2 n_dpc42_DL_ADH(eclk, ereset, dpc42_DL_ADH_port_8,dpc42_DL_ADH_port_9, dpc42_DL_ADH_v);
  spice_node_4 n_n_767(eclk, ereset, n_767_port_2,n_767_port_3,n_767_port_0,n_767_port_1, n_767_v);
  spice_node_3 n_n_953(eclk, ereset, n_953_port_2,n_953_port_0,n_953_port_1, n_953_v);
  spice_node_3 n_n_409(eclk, ereset, n_409_port_3,n_409_port_0,n_409_port_5, n_409_v);
  spice_node_3 n_n_1548(eclk, ereset, n_1548_port_2,n_1548_port_3,n_1548_port_1, n_1548_v);
  spice_node_3 n_n_1016(eclk, ereset, n_1016_port_2,n_1016_port_3,n_1016_port_1, n_1016_v);
  spice_node_3 n_p4(eclk, ereset, p4_port_2,p4_port_0,p4_port_1, p4_v);
  spice_node_3 n_n_171(eclk, ereset, n_171_port_3,n_171_port_0,n_171_port_1, n_171_v);
  spice_node_1 n_clk0(eclk, ereset, clk0_port_3, clk0_v);
  spice_node_5 n_n_1206(eclk, ereset, n_1206_port_2,n_1206_port_3,n_1206_port_0,n_1206_port_1,n_1206_port_4, n_1206_v);
  spice_node_2 n__ABH3(eclk, ereset, _ABH3_port_3,_ABH3_port_1, _ABH3_v);
  spice_node_2 n__ABH2(eclk, ereset, _ABH2_port_2,_ABH2_port_3, _ABH2_v);
  spice_node_2 n__ABH1(eclk, ereset, _ABH1_port_3,_ABH1_port_0, _ABH1_v);
  spice_node_2 n__ABH0(eclk, ereset, _ABH0_port_2,_ABH0_port_3, _ABH0_v);
  spice_node_2 n__ABH7(eclk, ereset, _ABH7_port_2,_ABH7_port_3, _ABH7_v);
  spice_node_2 n__ABH6(eclk, ereset, _ABH6_port_2,_ABH6_port_3, _ABH6_v);
  spice_node_2 n__ABH5(eclk, ereset, _ABH5_port_2,_ABH5_port_3, _ABH5_v);
  spice_node_2 n__ABH4(eclk, ereset, _ABH4_port_2,_ABH4_port_3, _ABH4_v);
  spice_node_3 n_n_1507(eclk, ereset, n_1507_port_2,n_1507_port_3,n_1507_port_1, n_1507_v);
  spice_node_3 n_n_423(eclk, ereset, n_423_port_2,n_423_port_0,n_423_port_1, n_423_v);
  spice_node_3 n_n_1254(eclk, ereset, n_1254_port_2,n_1254_port_0,n_1254_port_1, n_1254_v);
  spice_node_2 n_dpc18__DAA(eclk, ereset, dpc18__DAA_port_2,dpc18__DAA_port_1, dpc18__DAA_v);
  spice_node_2 n_dpc38_PCLADL(eclk, ereset, dpc38_PCLADL_port_9,dpc38_PCLADL_port_0, dpc38_PCLADL_v);
  spice_node_3 n_n_1691(eclk, ereset, n_1691_port_8,n_1691_port_1,n_1691_port_7, n_1691_v);
  spice_node_2 n_n_1696(eclk, ereset, n_1696_port_0,n_1696_port_1, n_1696_v);
  spice_node_2 n_n_855(eclk, ereset, n_855_port_2,n_855_port_0, n_855_v);
  spice_node_2 n_n_854(eclk, ereset, n_854_port_6,n_854_port_4, n_854_v);
  spice_node_3 n_n_994(eclk, ereset, n_994_port_2,n_994_port_3,n_994_port_1, n_994_v);
  spice_node_5 n_n_998(eclk, ereset, n_998_port_2,n_998_port_3,n_998_port_0,n_998_port_1,n_998_port_4, n_998_v);
  spice_node_3 n_n_999(eclk, ereset, n_999_port_2,n_999_port_3,n_999_port_1, n_999_v);
  spice_node_2 n_n_1501(eclk, ereset, n_1501_port_1,n_1501_port_4, n_1501_v);
  spice_node_2 n_n_298(eclk, ereset, n_298_port_3,n_298_port_4, n_298_v);
  spice_node_2 n_n_297(eclk, ereset, n_297_port_3,n_297_port_5, n_297_v);
  spice_node_5 n_n_296(eclk, ereset, n_296_port_3,n_296_port_0,n_296_port_1,n_296_port_4,n_296_port_5, n_296_v);
  spice_node_4 n_n_871(eclk, ereset, n_871_port_2,n_871_port_3,n_871_port_0,n_871_port_1, n_871_v);

endmodule

module spice_node_0(input eclk,ereset, output signed [`W-1:0] v);
  assign v = 0;
endmodule

module spice_node_1(input eclk,ereset, input signed [`W-1:0] i0, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_2(input eclk,ereset, input signed [`W-1:0] i0,i1, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_3(input eclk,ereset, input signed [`W-1:0] i0,i1,i2, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_4(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_5(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_6(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_7(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_8(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6,i7, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6+i7;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_12(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6+i7+i8+i9+i10+i11;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_13(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6+i7+i8+i9+i10+i11+i12;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

