* top-level ngspice script

.control
  source 4004-system.spice
  tran 5ns 240us
  write 4004-spice-rawfile.raw
.endc

.end
