* SPICE3 file created from 6502.ext - technology: nmos

.option scale=0.01u

M1000 nmi GND GND GND efet w=4888 l=752
+ ad=3.9117e+07 pd=103588 as=1.82881e+09 ps=2.64888e+07 
M1001 GND nmi n_1392 GND efet w=6580 l=658
+ ad=0 pd=0 as=7.24552e+06 ps=19364 
M1002 n_1392 n_1392 Vdd GND dfet w=846 l=1128
+ ad=1.87146e+07 pd=62980 as=0 ps=0 
M1003 GND pipeT4out n_1703 GND efet w=10340 l=658
+ ad=0 pd=0 as=1.19374e+07 ps=33088 
M1004 n_468 n_16 n_1703 GND efet w=5546 l=658
+ ad=7.8287e+06 pd=28764 as=0 ps=0 
M1005 GND pipeT5out n_1615 GND efet w=10998 l=658
+ ad=0 pd=0 as=9.86981e+06 ps=29892 
M1006 n_1615 notRdy0 n_468 GND efet w=7003 l=705
+ ad=0 pd=0 as=0 ps=0 
M1007 GND pipeT4out n_395 GND efet w=11656 l=658
+ ad=0 pd=0 as=7.24552e+06 ps=22936 
M1008 n_378 n_18 GND GND efet w=6251 l=611
+ ad=1.12571e+07 pd=32712 as=0 ps=0 
M1009 Vdd n_468 n_468 GND dfet w=940 l=1598
+ ad=0 pd=0 as=3.56974e+06 ps=9776 
M1010 n_395 notRdy0 n_472 GND efet w=4559 l=611
+ ad=0 pd=0 as=9.53404e+06 ps=26696 
M1011 GND n_378 _t5 GND efet w=6909 l=611
+ ad=0 pd=0 as=8.84484e+06 ps=22372 
M1012 pipeT5out cclk n_378 GND efet w=1128 l=846
+ ad=1.68768e+06 pd=7144 as=0 ps=0 
M1013 GND n_1392 n_284 GND efet w=3478 l=658
+ ad=0 pd=0 as=4.56821e+06 ps=12972 
M1014 GND NMIP n_645 GND efet w=4089 l=611
+ ad=0 pd=0 as=7.03346e+06 ps=26132 
M1015 n_891 cclk GND GND efet w=4324 l=658
+ ad=4.17059e+06 pd=12032 as=0 ps=0 
M1016 n_468 cp1 n_18 GND efet w=1128 l=752
+ ad=0 pd=0 as=2.82752e+06 ps=9588 
M1017 pipeT4out cclk n_188 GND efet w=1128 l=752
+ ad=2.21784e+06 pd=8648 as=1.52863e+07 ps=42864 
M1018 n_472 n_16 n_1366 GND efet w=5217 l=705
+ ad=0 pd=0 as=9.78145e+06 ps=26132 
M1019 GND pipeT3out n_1366 GND efet w=10340 l=658
+ ad=0 pd=0 as=0 ps=0 
M1020 n_378 n_378 Vdd GND dfet w=940 l=1598
+ ad=8.21748e+06 pd=27072 as=0 ps=0 
M1021 GND n_1357 n_378 GND efet w=4418 l=658
+ ad=0 pd=0 as=0 ps=0 
M1022 NMIP n_284 n_891 GND efet w=4512 l=658
+ ad=8.4914e+06 pd=26320 as=0 ps=0 
M1023 n_284 n_284 Vdd GND dfet w=940 l=1128
+ ad=8.75648e+06 pd=28764 as=0 ps=0 
M1024 GND nNMIP NMIP GND efet w=2350 l=658
+ ad=0 pd=0 as=0 ps=0 
M1025 nNMIP NMIP GND GND efet w=2350 l=564
+ ad=6.4061e+06 pd=20492 as=0 ps=0 
M1026 n_346 n_1392 nNMIP GND efet w=4418 l=658
+ ad=2.07646e+06 pd=9776 as=0 ps=0 
M1027 GND cclk n_346 GND efet w=4418 l=564
+ ad=0 pd=0 as=0 ps=0 
M1028 irq GND GND GND efet w=4794 l=752
+ ad=4.11758e+07 pd=109228 as=0 ps=0 
M1029 Vdd n_472 n_472 GND dfet w=940 l=1504
+ ad=0 pd=0 as=3.44604e+06 ps=9400 
M1030 _t5 _t5 Vdd GND dfet w=940 l=564
+ ad=1.81288e+08 pd=586372 as=0 ps=0 
M1031 n_645 n_645 Vdd GND dfet w=846 l=940
+ ad=5.36434e+07 pd=188564 as=0 ps=0 
M1032 NMIP NMIP Vdd GND dfet w=658 l=1316
+ ad=1.25383e+07 pd=43992 as=0 ps=0 
M1033 nNMIP nNMIP Vdd GND dfet w=940 l=1504
+ ad=7.10414e+06 pd=20868 as=0 ps=0 
M1034 GND irq n_1599 GND efet w=5828 l=564
+ ad=0 pd=0 as=7.5106e+06 ps=19740 
M1035 n_881 cclk GND GND efet w=5029 l=611
+ ad=7.13949e+06 pd=16168 as=0 ps=0 
M1036 n_538 n_1599 GND GND efet w=3149 l=611
+ ad=5.15139e+06 pd=13724 as=0 ps=0 
M1037 GND n_807 n_330 GND efet w=2256 l=658
+ ad=0 pd=0 as=1.22909e+07 ps=30456 
M1038 n_431 n_1599 n_807 GND efet w=5499 l=611
+ ad=5.7434e+06 pd=16168 as=8.57092e+06 ps=22936 
M1039 n_1599 n_1599 Vdd GND dfet w=1034 l=1222
+ ad=1.97838e+07 pd=66176 as=0 ps=0 
M1040 n_538 n_538 Vdd GND dfet w=940 l=1128
+ ad=6.54748e+06 pd=21056 as=0 ps=0 
M1041 n_881 n_538 n_330 GND efet w=5123 l=611
+ ad=0 pd=0 as=0 ps=0 
M1042 GND n_330 n_807 GND efet w=3102 l=658
+ ad=0 pd=0 as=0 ps=0 
M1043 GND cclk n_431 GND efet w=4324 l=658
+ ad=0 pd=0 as=0 ps=0 
M1044 n_806 GND GND GND efet w=4324 l=752
+ ad=3.07493e+07 pd=25568 as=0 ps=0 
M1045 n_807 n_807 Vdd GND dfet w=846 l=1316
+ ad=6.80372e+06 pd=22936 as=0 ps=0 
M1046 GND IRQP nIRQP GND efet w=3948 l=564
+ ad=0 pd=0 as=9.75494e+06 ps=22560 
M1047 n_330 n_330 Vdd GND dfet w=940 l=1316
+ ad=5.5225e+06 pd=18424 as=0 ps=0 
M1048 IRQP cp1 n_330 GND efet w=1128 l=752
+ ad=1.2017e+06 pd=6580 as=0 ps=0 
M1049 GND IRQP nIRQP GND efet w=4512 l=658
+ ad=0 pd=0 as=0 ps=0 
M1050 nIRQP nIRQP Vdd GND dfet w=1034 l=940
+ ad=4.48427e+07 pd=164500 as=0 ps=0 
M1051 clk1out n_1417 GND GND efet w=9776 l=564
+ ad=1.08541e+08 pd=153596 as=0 ps=0 
M1052 GND n_1417 clk1out GND efet w=20774 l=564
+ ad=0 pd=0 as=0 ps=0 
M1053 clk1out n_1417 GND GND efet w=20774 l=658
+ ad=0 pd=0 as=0 ps=0 
M1054 GND n_1417 clk1out GND efet w=20774 l=564
+ ad=0 pd=0 as=0 ps=0 
M1055 clk1out n_1417 GND GND efet w=20774 l=564
+ ad=0 pd=0 as=0 ps=0 
M1056 GND n_747 n_1417 GND efet w=21291 l=705
+ ad=0 pd=0 as=3.30643e+07 ps=49256 
M1057 GND n_670 n_747 GND efet w=25991 l=705
+ ad=0 pd=0 as=3.96383e+07 ps=57528 
M1058 GND GND rdy GND efet w=4794 l=658
+ ad=0 pd=0 as=4.3049e+07 ps=117500 
M1059 GND rdy n_958 GND efet w=14006 l=752
+ ad=0 pd=0 as=1.34661e+07 ps=38540 
M1060 rdy rdy Vdd GND dfet w=940 l=1504
+ ad=2.05702e+07 pd=64108 as=0 ps=0 
M1061 n_420 n_865 GND GND efet w=5076 l=658
+ ad=7.89055e+06 pd=27824 as=0 ps=0 
M1062 n_47 cp1 n_420 GND efet w=1222 l=658
+ ad=1.35191e+06 pd=6016 as=0 ps=0 
M1063 n_1449 n_958 GND GND efet w=11139 l=611
+ ad=1.05679e+07 pd=33464 as=0 ps=0 
M1064 n_865 cclk n_958 GND efet w=1222 l=752
+ ad=1.52863e+06 pd=6016 as=0 ps=0 
M1065 GND n_47 n_603 GND efet w=4747 l=705
+ ad=0 pd=0 as=4.957e+06 ps=15228 
M1066 clk1out n_747 Vdd GND dfet w=6392 l=658
+ ad=0 pd=0 as=7.31435e+08 ps=1.00682e+07 
M1067 n_1417 n_670 Vdd GND dfet w=2350 l=752
+ ad=0 pd=0 as=0 ps=0 
M1068 Vdd n_747 n_747 GND dfet w=2444 l=752
+ ad=0 pd=0 as=2.50236e+07 ps=76704 
M1069 n_420 n_420 Vdd GND dfet w=940 l=1598
+ ad=4.1971e+06 pd=10152 as=0 ps=0 
M1070 n_958 n_958 Vdd GND dfet w=846 l=564
+ ad=1.43585e+07 pd=49632 as=0 ps=0 
M1071 n_603 n_603 Vdd GND dfet w=940 l=1598
+ ad=4.84478e+07 pd=169388 as=0 ps=0 
M1072 clk2out n_135 GND GND efet w=31208 l=658
+ ad=9.27161e+07 pd=141376 as=0 ps=0 
M1073 GND GND res GND efet w=7379 l=705
+ ad=0 pd=0 as=4.72196e+07 ps=124080 
M1074 n_312 res GND GND efet w=7379 l=611
+ ad=8.50907e+06 pd=26132 as=0 ps=0 
M1075 Vdd n_1449 n_1449 GND dfet w=1504 l=658
+ ad=0 pd=0 as=7.21901e+07 ps=281812 
M1076 GND n_312 n_995 GND efet w=3008 l=564
+ ad=0 pd=0 as=5.18673e+06 ps=14664 
M1077 n_886 cclk GND GND efet w=4418 l=564
+ ad=2.07646e+06 pd=9776 as=0 ps=0 
M1078 n_975 n_995 n_886 GND efet w=4418 l=658
+ ad=6.77721e+06 pd=18048 as=0 ps=0 
M1079 GND n_854 n_975 GND efet w=2350 l=564
+ ad=0 pd=0 as=0 ps=0 
M1080 n_854 n_975 GND GND efet w=2350 l=564
+ ad=8.66812e+06 pd=29516 as=0 ps=0 
M1081 n_742 n_312 n_854 GND efet w=4418 l=564
+ ad=2.07646e+06 pd=9776 as=0 ps=0 
M1082 GND cclk n_742 GND efet w=4418 l=658
+ ad=0 pd=0 as=0 ps=0 
M1083 GND n_1395 Reset0 GND efet w=7379 l=705
+ ad=0 pd=0 as=1.47208e+07 ps=39292 
M1084 n_1395 cp1 n_854 GND efet w=1128 l=752
+ ad=1.4226e+06 pd=5828 as=0 ps=0 
M1085 n_312 n_312 Vdd GND dfet w=940 l=1128
+ ad=1.42878e+07 pd=50572 as=0 ps=0 
M1086 n_995 n_995 Vdd GND dfet w=1034 l=1128
+ ad=1.07446e+07 pd=36284 as=0 ps=0 
M1087 n_975 n_975 Vdd GND dfet w=846 l=1316
+ ad=5.70806e+06 pd=18048 as=0 ps=0 
M1088 n_854 n_854 Vdd GND dfet w=846 l=1316
+ ad=1.2715e+07 pd=45684 as=0 ps=0 
M1089 Reset0 n_1395 GND GND efet w=6674 l=658
+ ad=0 pd=0 as=0 ps=0 
M1090 GND n_519 n_670 GND efet w=8272 l=658
+ ad=0 pd=0 as=1.85114e+07 ps=45684 
M1091 Vdd Reset0 Reset0 GND dfet w=940 l=846
+ ad=0 pd=0 as=1.25789e+08 ps=458908 
M1092 n_670 n_670 Vdd GND dfet w=2350 l=658
+ ad=3.40716e+07 pd=108476 as=0 ps=0 
M1093 GND n_519 n_670 GND efet w=7990 l=846
+ ad=0 pd=0 as=0 ps=0 
M1094 clk2out n_135 GND GND efet w=22184 l=658
+ ad=0 pd=0 as=0 ps=0 
M1095 GND n_135 clk2out GND efet w=22184 l=564
+ ad=0 pd=0 as=0 ps=0 
M1096 clk2out n_135 GND GND efet w=22184 l=752
+ ad=0 pd=0 as=0 ps=0 
M1097 Vdd n_127 clk2out GND dfet w=6298 l=658
+ ad=0 pd=0 as=0 ps=0 
M1098 n_135 n_519 Vdd GND dfet w=2256 l=658
+ ad=2.01991e+07 pd=48128 as=0 ps=0 
M1099 GND n_127 n_135 GND efet w=20915 l=611
+ ad=0 pd=0 as=0 ps=0 
M1100 n_127 cp1 GND GND efet w=11844 l=658
+ ad=2.69056e+07 pd=60912 as=0 ps=0 
M1101 GND n_519 n_127 GND efet w=21291 l=611
+ ad=0 pd=0 as=0 ps=0 
M1102 GND clk0 n_519 GND efet w=26367 l=611
+ ad=0 pd=0 as=2.4732e+07 ps=60536 
M1103 GND GND so GND efet w=4324 l=658
+ ad=0 pd=0 as=5.3714e+07 ps=137992 
M1104 clk0 GND GND GND efet w=5217 l=705
+ ad=7.53534e+07 pd=181044 as=0 ps=0 
M1105 n_127 n_127 Vdd GND dfet w=2350 l=752
+ ad=3.27109e+07 pd=106596 as=0 ps=0 
M1106 n_519 n_519 Vdd GND dfet w=2350 l=658
+ ad=5.11516e+07 pd=163936 as=0 ps=0 
M1107 n_1650 cp1 n_94 GND efet w=1128 l=752
+ ad=1.30684e+07 pd=32524 as=1.96159e+06 ps=7332 
M1108 so so Vdd GND dfet w=940 l=1504
+ ad=1.82905e+07 pd=62228 as=0 ps=0 
M1109 n_1069 n_1024 GND GND efet w=2820 l=658
+ ad=1.19993e+07 pd=31584 as=0 ps=0 
M1110 n_1069 n_1069 Vdd GND dfet w=940 l=1222
+ ad=4.0195e+07 pd=141376 as=0 ps=0 
M1111 GND n_1274 n_1069 GND efet w=5922 l=658
+ ad=0 pd=0 as=0 ps=0 
M1112 n_1024 cclk n_1699 GND efet w=1128 l=658
+ ad=1.46147e+07 pd=43428 as=1.23704e+06 ps=6956 
M1113 n_913 n_1699 GND GND efet w=4136 l=564
+ ad=6.56515e+06 pd=21808 as=0 ps=0 
M1114 GND n_94 n_1024 GND efet w=5922 l=564
+ ad=0 pd=0 as=0 ps=0 
M1115 n_913 cp1 n_1274 GND efet w=1128 l=752
+ ad=0 pd=0 as=1.94392e+06 ps=6768 
M1116 n_1024 n_1024 Vdd GND dfet w=940 l=1316
+ ad=6.19404e+06 pd=20868 as=0 ps=0 
M1117 GND so n_1650 GND efet w=11562 l=658
+ ad=0 pd=0 as=0 ps=0 
M1118 Vdd op_sty_cpy_mem op_sty_cpy_mem GND dfet w=846 l=1786
+ ad=0 pd=0 as=2.24611e+07 ps=70124 
M1119 Vdd _t4 _t4 GND dfet w=846 l=564
+ ad=0 pd=0 as=1.63386e+08 ps=576408 
M1120 n_472 cp1 n_1606 GND efet w=1128 l=752
+ ad=0 pd=0 as=1.63466e+06 ps=7520 
M1121 Vdd n_188 n_188 GND dfet w=940 l=1222
+ ad=0 pd=0 as=1.24499e+07 ps=39104 
M1122 _t4 n_188 GND GND efet w=9071 l=705
+ ad=5.3988e+06 pd=19364 as=0 ps=0 
M1123 n_188 n_1606 GND GND efet w=6956 l=564
+ ad=0 pd=0 as=0 ps=0 
M1124 Vdd op_T2_abs_y op_T2_abs_y GND dfet w=846 l=1786
+ ad=0 pd=0 as=7.02462e+06 ps=19176 
M1125 Vdd op_T3_ind_y op_T3_ind_y GND dfet w=846 l=1692
+ ad=0 pd=0 as=9.96701e+06 ps=31772 
M1126 Vdd x_op_T0_tya x_op_T0_tya GND dfet w=846 l=1786
+ ad=0 pd=0 as=7.61663e+06 ps=20304 
M1127 Vdd op_T0_iny_dey op_T0_iny_dey GND dfet w=940 l=1786
+ ad=0 pd=0 as=7.13949e+06 ps=21056 
M1128 Vdd op_xy op_xy GND dfet w=846 l=1786
+ ad=0 pd=0 as=1.79017e+07 ps=56400 
M1129 Vdd op_T0_cpy_iny op_T0_cpy_iny GND dfet w=846 l=1786
+ ad=0 pd=0 as=7.02462e+06 ps=21432 
M1130 Vdd op_T2_idx_x_xy op_T2_idx_x_xy GND dfet w=940 l=1786
+ ad=0 pd=0 as=2.07204e+07 ps=66740 
M1131 Vdd x_op_T0_txa x_op_T0_txa GND dfet w=940 l=1786
+ ad=0 pd=0 as=6.75954e+06 ps=19176 
M1132 Vdd op_T0_cpx_inx op_T0_cpx_inx GND dfet w=893 l=1739
+ ad=0 pd=0 as=6.86557e+06 ps=18988 
M1133 Vdd op_T2_ind_x op_T2_ind_x GND dfet w=940 l=1786
+ ad=0 pd=0 as=7.4134e+06 ps=21996 
M1134 Vdd op_T0_dex op_T0_dex GND dfet w=846 l=1786
+ ad=0 pd=0 as=6.86557e+06 ps=21244 
M1135 Vdd op_T0_txs op_T0_txs GND dfet w=846 l=1786
+ ad=0 pd=0 as=1.72479e+07 ps=59032 
M1136 Vdd op_from_x op_from_x GND dfet w=940 l=1786
+ ad=0 pd=0 as=2.21077e+07 ps=75952 
M1137 Vdd op_T__dex op_T__dex GND dfet w=846 l=1692
+ ad=0 pd=0 as=5.34578e+06 ps=16920 
M1138 Vdd op_T0_ldx_tax_tsx op_T0_ldx_tax_tsx GND dfet w=1034 l=1786
+ ad=0 pd=0 as=7.61663e+06 ps=24064 
M1139 Vdd op_T0_tsx op_T0_tsx GND dfet w=940 l=1786
+ ad=0 pd=0 as=1.30066e+07 ps=41924 
M1140 Vdd op_T0_ldy_mem op_T0_ldy_mem GND dfet w=846 l=1786
+ ad=0 pd=0 as=7.75801e+06 ps=22372 
M1141 Vdd op_T__inx op_T__inx GND dfet w=846 l=1786
+ ad=0 pd=0 as=6.77721e+06 ps=21056 
M1142 Vdd op_T__iny_dey op_T__iny_dey GND dfet w=846 l=1786
+ ad=0 pd=0 as=6.17636e+06 ps=19928 
M1143 Vdd op_T0_tay_ldy_not_idx op_T0_tay_ldy_not_idx GND dfet w=846 l=1786
+ ad=0 pd=0 as=7.6343e+06 ps=24064 
M1144 Vdd op_T5_brk op_T5_brk GND dfet w=940 l=1786
+ ad=0 pd=0 as=1.12659e+07 ps=33088 
M1145 Vdd op_T0_jsr op_T0_jsr GND dfet w=940 l=1786
+ ad=0 pd=0 as=1.79901e+07 ps=59596 
M1146 Vdd op_T4_rts op_T4_rts GND dfet w=940 l=1786
+ ad=0 pd=0 as=6.56515e+06 ps=18048 
M1147 Vdd op_T5_rti op_T5_rti GND dfet w=893 l=1833
+ ad=0 pd=0 as=4.21742e+07 ps=160552 
M1148 Vdd op_T0_php_pha op_T0_php_pha GND dfet w=940 l=1786
+ ad=0 pd=0 as=6.93626e+06 ps=20304 
M1149 GND n_1357 n_188 GND efet w=4559 l=611
+ ad=0 pd=0 as=0 ps=0 
M1150 GND pipeT3out n_1456 GND efet w=11985 l=705
+ ad=0 pd=0 as=6.91859e+06 ps=23124 
M1151 Vdd op_T3_plp_pla op_T3_plp_pla GND dfet w=846 l=1786
+ ad=0 pd=0 as=7.3869e+06 ps=21244 
M1152 Vdd op_T2 op_T2 GND dfet w=940 l=1786
+ ad=0 pd=0 as=4.40916e+07 ps=156604 
M1153 Vdd op_ror op_ror GND dfet w=1034 l=1786
+ ad=0 pd=0 as=1.88207e+07 ps=61664 
M1154 Vdd op_jmp op_jmp GND dfet w=846 l=1786
+ ad=0 pd=0 as=1.66647e+07 ps=55836 
M1155 Vdd op_T0_eor op_T0_eor GND dfet w=940 l=1786
+ ad=0 pd=0 as=2.35921e+07 ps=84600 
M1156 Vdd op_T0_ora op_T0_ora GND dfet w=846 l=1786
+ ad=0 pd=0 as=2.03935e+07 ps=65612 
M1157 Vdd op_T2_abs op_T2_abs GND dfet w=940 l=1786
+ ad=0 pd=0 as=1.75571e+07 ps=59032 
M1158 Vdd op_T0 op_T0 GND dfet w=846 l=1786
+ ad=0 pd=0 as=9.51637e+06 ps=28952 
M1159 Vdd op_T2_ADL_ADD op_T2_ADL_ADD GND dfet w=846 l=1786
+ ad=0 pd=0 as=1.66205e+07 ps=56588 
M1160 Vdd op_T3_stack_bit_jmp op_T3_stack_bit_jmp GND dfet w=940 l=1786
+ ad=0 pd=0 as=7.09531e+06 ps=20116 
M1161 Vdd op_T2_stack op_T2_stack GND dfet w=846 l=1786
+ ad=0 pd=0 as=1.67707e+07 ps=55460 
M1162 Vdd op_T4_rti op_T4_rti GND dfet w=940 l=1786
+ ad=0 pd=0 as=6.33541e+06 ps=18424 
M1163 Vdd op_T4_brk_jsr op_T4_brk_jsr GND dfet w=940 l=1786
+ ad=0 pd=0 as=7.33388e+06 ps=22184 
M1164 Vdd op_T4_ind_y op_T4_ind_y GND dfet w=846 l=1786
+ ad=0 pd=0 as=8.35886e+06 ps=26508 
M1165 Vdd op_T3_ind_x op_T3_ind_x GND dfet w=940 l=1786
+ ad=0 pd=0 as=1.0347e+07 ps=37788 
M1166 Vdd op_T3_abs_idx op_T3_abs_idx GND dfet w=846 l=1786
+ ad=0 pd=0 as=8.46489e+06 ps=26132 
M1167 Vdd op_T2_ind_y op_T2_ind_y GND dfet w=846 l=1692
+ ad=0 pd=0 as=9.02156e+06 ps=27448 
M1168 Vdd op_inc_nop op_inc_nop GND dfet w=846 l=1786
+ ad=0 pd=0 as=1.05944e+07 ps=29140 
M1169 Vdd op_plp_pla op_plp_pla GND dfet w=940 l=1786
+ ad=0 pd=0 as=8.35886e+06 ps=27260 
M1170 Vdd x_op_T3_ind_y x_op_T3_ind_y GND dfet w=846 l=1692
+ ad=0 pd=0 as=7.31621e+06 ps=21244 
M1171 Vdd op_T4_ind_x op_T4_ind_x GND dfet w=893 l=1833
+ ad=0 pd=0 as=1.67531e+07 ps=59032 
M1172 Vdd op_T2_jsr op_T2_jsr GND dfet w=846 l=1786
+ ad=0 pd=0 as=2.07734e+07 ps=71064 
M1173 Vdd op_rti_rts op_rti_rts GND dfet w=846 l=1786
+ ad=0 pd=0 as=2.17012e+07 ps=70876 
M1174 Vdd op_T0_cmp op_T0_cmp GND dfet w=846 l=1786
+ ad=0 pd=0 as=7.50176e+06 ps=22184 
M1175 Vdd op_T0_cpx_cpy_inx_iny op_T0_cpx_cpy_inx_iny GND dfet w=846 l=1786
+ ad=0 pd=0 as=7.91706e+06 ps=24816 
M1176 Vdd op_T0_adc_sbc op_T0_adc_sbc GND dfet w=846 l=1786
+ ad=0 pd=0 as=3.21454e+07 ps=120132 
M1177 Vdd op_T3_jmp op_T3_jmp GND dfet w=846 l=1786
+ ad=0 pd=0 as=7.40457e+06 ps=21808 
M1178 Vdd op_T0_sbc op_T0_sbc GND dfet w=846 l=1786
+ ad=0 pd=0 as=4.46395e+07 ps=158860 
M1179 Vdd op_rol_ror op_rol_ror GND dfet w=940 l=1786
+ ad=0 pd=0 as=1.00907e+07 ps=30456 
M1180 Vdd op_T5_jsr op_T5_jsr GND dfet w=940 l=1786
+ ad=0 pd=0 as=2.39721e+07 ps=87044 
M1181 op_shift op_shift Vdd GND dfet w=940 l=1786
+ ad=1.64438e+07 pd=53392 as=0 ps=0 
M1182 Vdd op_T0_tya op_T0_tya GND dfet w=846 l=1692
+ ad=0 pd=0 as=7.68732e+06 ps=21620 
M1183 Vdd op_T2_stack_access op_T2_stack_access GND dfet w=940 l=1786
+ ad=0 pd=0 as=1.4385e+07 ps=51136 
M1184 Vdd op_T__adc_sbc op_T__adc_sbc GND dfet w=940 l=1692
+ ad=0 pd=0 as=9.71076e+06 ps=31584 
M1185 Vdd op_T__ora_and_eor_adc op_T__ora_and_eor_adc GND dfet w=752 l=1786
+ ad=0 pd=0 as=1.27238e+07 ps=45684 
M1186 Vdd op_T0_txa op_T0_txa GND dfet w=846 l=1786
+ ad=0 pd=0 as=7.5106e+06 ps=20868 
M1187 Vdd op_T__shift_a op_T__shift_a GND dfet w=846 l=1692
+ ad=0 pd=0 as=7.5106e+06 ps=23124 
M1188 Vdd op_T0_lda op_T0_lda GND dfet w=940 l=1786
+ ad=0 pd=0 as=9.76378e+06 ps=28388 
M1189 Vdd op_T0_pla op_T0_pla GND dfet w=940 l=1786
+ ad=0 pd=0 as=7.33388e+06 ps=21432 
M1190 Vdd op_T0_tay op_T0_tay GND dfet w=846 l=1786
+ ad=0 pd=0 as=7.36922e+06 ps=20868 
M1191 Vdd op_T0_acc op_T0_acc GND dfet w=940 l=1692
+ ad=0 pd=0 as=8.70346e+06 ps=26132 
M1192 Vdd op_T0_tax op_T0_tax GND dfet w=846 l=1786
+ ad=0 pd=0 as=8.15563e+06 ps=22184 
M1193 Vdd op_T0_shift_a op_T0_shift_a GND dfet w=846 l=1786
+ ad=0 pd=0 as=1.86351e+07 ps=63732 
M1194 Vdd op_T0_and op_T0_and GND dfet w=846 l=1786
+ ad=0 pd=0 as=8.63277e+06 ps=24628 
M1195 Vdd op_T0_bit op_T0_bit GND dfet w=893 l=1833
+ ad=0 pd=0 as=1.01879e+07 ps=31208 
M1196 Vdd op_T5_ind_y op_T5_ind_y GND dfet w=846 l=1786
+ ad=0 pd=0 as=8.0496e+06 ps=24064 
M1197 Vdd op_T4_abs_idx op_T4_abs_idx GND dfet w=940 l=1692
+ ad=0 pd=0 as=9.96701e+06 ps=30080 
M1198 Vdd op_branch_done op_branch_done GND dfet w=846 l=1692
+ ad=0 pd=0 as=4.31462e+07 ps=153972 
M1199 Vdd op_T0_shift_right_a op_T0_shift_right_a GND dfet w=846 l=1692
+ ad=0 pd=0 as=7.98774e+06 ps=23688 
M1200 Vdd op_T2_pha op_T2_pha GND dfet w=940 l=1692
+ ad=0 pd=0 as=1.53393e+07 ps=53392 
M1201 Vdd op_T2_brk op_T2_brk GND dfet w=846 l=1786
+ ad=0 pd=0 as=6.90975e+06 ps=20116 
M1202 op_branch_done n_603 GND GND efet w=1692 l=658
+ ad=1.21495e+07 pd=33088 as=0 ps=0 
M1203 Vdd op_shift_right op_shift_right GND dfet w=846 l=1786
+ ad=0 pd=0 as=9.25129e+06 ps=28012 
M1204 Vdd op_sta_cmp op_sta_cmp GND dfet w=846 l=1692
+ ad=0 pd=0 as=2.07027e+07 ps=71440 
M1205 Vdd op_T3_jsr op_T3_jsr GND dfet w=940 l=1786
+ ad=0 pd=0 as=8.19097e+06 ps=23688 
M1206 Vdd op_T2_zp_zp_idx op_T2_zp_zp_idx GND dfet w=846 l=1786
+ ad=0 pd=0 as=1.66824e+07 ps=52452 
M1207 n_913 n_913 Vdd GND dfet w=940 l=1504
+ ad=5.0807e+06 pd=15040 as=0 ps=0 
M1208 cp1 n_1105 GND GND efet w=18612 l=658
+ ad=3.19201e+08 pd=535236 as=0 ps=0 
M1209 GND n_1105 cp1 GND efet w=18800 l=658
+ ad=0 pd=0 as=0 ps=0 
M1210 cp1 n_1105 GND GND efet w=18612 l=752
+ ad=0 pd=0 as=0 ps=0 
M1211 GND n_1105 cp1 GND efet w=18847 l=611
+ ad=0 pd=0 as=0 ps=0 
M1212 cp1 n_1105 GND GND efet w=18612 l=752
+ ad=0 pd=0 as=0 ps=0 
M1213 Vdd n_1399 cp1 GND dfet w=6392 l=658
+ ad=0 pd=0 as=0 ps=0 
M1214 n_1650 n_1650 Vdd GND dfet w=940 l=658
+ ad=2.51826e+06 pd=10152 as=0 ps=0 
M1215 n_1105 n_1715 Vdd GND dfet w=2256 l=564
+ ad=2.29471e+07 pd=51700 as=0 ps=0 
M1216 GND n_1399 n_1105 GND efet w=20868 l=658
+ ad=0 pd=0 as=0 ps=0 
M1217 n_1399 n_1715 GND GND efet w=9212 l=658
+ ad=2.06674e+07 pd=48880 as=0 ps=0 
M1218 GND n_1715 n_1399 GND efet w=17437 l=611
+ ad=0 pd=0 as=0 ps=0 
M1219 GND n_358 n_1715 GND efet w=14570 l=564
+ ad=0 pd=0 as=2.34596e+07 ps=49068 
M1220 Vdd n_1399 n_1399 GND dfet w=2350 l=658
+ ad=0 pd=0 as=2.55625e+07 ps=79524 
M1221 Vdd n_1715 n_1715 GND dfet w=2350 l=658
+ ad=0 pd=0 as=4.03894e+07 ps=135548 
M1222 GND n_1467 cclk GND efet w=23218 l=564
+ ad=0 pd=0 as=5.32449e+08 ps=894880 
M1223 cclk n_1467 GND GND efet w=23218 l=564
+ ad=0 pd=0 as=0 ps=0 
M1224 GND n_1467 cclk GND efet w=23218 l=564
+ ad=0 pd=0 as=0 ps=0 
M1225 cclk n_1467 GND GND efet w=23218 l=564
+ ad=0 pd=0 as=0 ps=0 
M1226 Vdd n_1129 cclk GND dfet w=6392 l=752
+ ad=0 pd=0 as=0 ps=0 
M1227 n_1467 n_358 Vdd GND dfet w=2350 l=564
+ ad=2.45641e+07 pd=52828 as=0 ps=0 
M1228 GND n_1129 n_1467 GND efet w=20680 l=658
+ ad=0 pd=0 as=0 ps=0 
M1229 n_1129 n_358 GND GND efet w=3666 l=564
+ ad=2.40693e+07 pd=51888 as=0 ps=0 
M1230 n_1129 cp1 GND GND efet w=10528 l=564
+ ad=0 pd=0 as=0 ps=0 
M1231 GND n_358 n_1129 GND efet w=16638 l=564
+ ad=0 pd=0 as=0 ps=0 
M1232 n_358 clk0 GND GND efet w=26696 l=658
+ ad=1.8697e+07 pd=38728 as=0 ps=0 
M1233 n_358 n_358 Vdd GND dfet w=2350 l=564
+ ad=4.22803e+07 pd=155476 as=0 ps=0 
M1234 Vdd n_1129 n_1129 GND dfet w=2350 l=658
+ ad=0 pd=0 as=3.54147e+07 ps=110168 
M1235 rw n_102 Vdd GND efet w=13066 l=658
+ ad=1.33123e+08 pd=209996 as=0 ps=0 
M1236 Vdd n_102 rw GND efet w=13066 l=564
+ ad=0 pd=0 as=0 ps=0 
M1237 GND GND clk0 GND efet w=4418 l=752
+ ad=0 pd=0 as=0 ps=0 
M1238 rw n_102 Vdd GND efet w=13019 l=611
+ ad=0 pd=0 as=0 ps=0 
M1239 Vdd n_102 rw GND efet w=12972 l=658
+ ad=0 pd=0 as=0 ps=0 
M1240 rw n_102 Vdd GND efet w=12972 l=658
+ ad=0 pd=0 as=0 ps=0 
M1241 Vdd n_102 rw GND efet w=12972 l=658
+ ad=0 pd=0 as=0 ps=0 
M1242 rw n_102 Vdd GND efet w=14617 l=611
+ ad=0 pd=0 as=0 ps=0 
M1243 n_633 cclk n_1059 GND efet w=940 l=1504
+ ad=3.6581e+06 pd=9212 as=9.90516e+06 ps=22560 
M1244 rw n_1696 GND GND efet w=14194 l=658
+ ad=0 pd=0 as=0 ps=0 
M1245 GND n_1696 rw GND efet w=14194 l=658
+ ad=0 pd=0 as=0 ps=0 
M1246 rw n_1696 GND GND efet w=14194 l=564
+ ad=0 pd=0 as=0 ps=0 
M1247 GND n_1696 rw GND efet w=14194 l=658
+ ad=0 pd=0 as=0 ps=0 
M1248 rw n_1696 GND GND efet w=20069 l=611
+ ad=0 pd=0 as=0 ps=0 
M1249 GND n_400 n_102 GND efet w=11562 l=752
+ ad=0 pd=0 as=1.06562e+07 ps=28388 
M1250 GND GND cclk GND efet w=5217 l=611
+ ad=0 pd=0 as=0 ps=0 
M1251 n_834 n_402 GND GND efet w=6674 l=658
+ ad=4.72726e+06 pd=15980 as=0 ps=0 
M1252 n_102 n_834 Vdd GND dfet w=1598 l=658
+ ad=0 pd=0 as=0 ps=0 
M1253 Vdd op_T2_abs_access op_T2_abs_access GND dfet w=846 l=1786
+ ad=0 pd=0 as=5.36345e+07 ps=186684 
M1254 Vdd op_T2_branch op_T2_branch GND dfet w=846 l=1692
+ ad=0 pd=0 as=1.41641e+07 ps=47376 
M1255 op_T2_ind op_T2_ind Vdd GND dfet w=940 l=1786
+ ad=1.07446e+07 pd=34216 as=0 ps=0 
M1256 Vdd op_T4 op_T4 GND dfet w=846 l=1786
+ ad=0 pd=0 as=7.90822e+06 ps=22372 
M1257 op_T5_rts op_T5_rts Vdd GND dfet w=940 l=1786
+ ad=5.50571e+07 pd=197400 as=0 ps=0 
M1258 Vdd op_T0_brk_rti op_T0_brk_rti GND dfet w=846 l=1786
+ ad=0 pd=0 as=8.80949e+06 ps=25004 
M1259 Vdd op_T5_ind_x op_T5_ind_x GND dfet w=846 l=1786
+ ad=0 pd=0 as=9.95817e+06 ps=29704 
M1260 Vdd op_T3 op_T3 GND dfet w=846 l=1786
+ ad=0 pd=0 as=8.05843e+06 ps=23688 
M1261 Vdd op_T0_jmp op_T0_jmp GND dfet w=846 l=1786
+ ad=0 pd=0 as=8.45605e+06 ps=25944 
M1262 Vdd x_op_T3_abs_idx x_op_T3_abs_idx GND dfet w=846 l=1786
+ ad=0 pd=0 as=7.67848e+06 ps=21056 
M1263 Vdd op_brk_rti op_brk_rti GND dfet w=846 l=1786
+ ad=0 pd=0 as=7.30737e+06 ps=20680 
M1264 Vdd op_T3_abs_idx_ind op_T3_abs_idx_ind GND dfet w=940 l=1692
+ ad=0 pd=0 as=7.37806e+06 ps=23688 
M1265 Vdd x_op_T4_ind_y x_op_T4_ind_y GND dfet w=846 l=1786
+ ad=0 pd=0 as=9.50754e+06 ps=30456 
M1266 Vdd op_T3_branch op_T3_branch GND dfet w=846 l=1692
+ ad=0 pd=0 as=1.7619e+07 ps=60536 
M1267 Vdd x_op_jmp x_op_jmp GND dfet w=940 l=1786
+ ad=0 pd=0 as=1.04265e+07 ps=31396 
M1268 Vdd diff_244212_338400# n_9 GND dfet w=940 l=1786
+ ad=0 pd=0 as=2.27969e+06 ps=6204 
M1269 Vdd op_jsr op_jsr GND dfet w=893 l=1833
+ ad=0 pd=0 as=6.58282e+06 ps=20304 
M1270 Vdd op_push_pull op_push_pull GND dfet w=846 l=1786
+ ad=0 pd=0 as=2.08618e+07 ps=77080 
M1271 Vdd op_T4_brk op_T4_brk GND dfet w=846 l=1786
+ ad=0 pd=0 as=1.45087e+07 ps=46248 
M1272 Vdd op_store op_store GND dfet w=940 l=1786
+ ad=0 pd=0 as=8.64161e+06 ps=26320 
M1273 Vdd op_T2_php_pha op_T2_php_pha GND dfet w=846 l=1786
+ ad=0 pd=0 as=1.34307e+07 ps=40984 
M1274 Vdd n_173 n_173 GND dfet w=846 l=1786
+ ad=0 pd=0 as=3.26048e+06 ps=7708 
M1275 Vdd op_T2_php op_T2_php GND dfet w=752 l=1786
+ ad=0 pd=0 as=7.74034e+06 ps=22748 
M1276 Vdd op_T4_jmp op_T4_jmp GND dfet w=940 l=1786
+ ad=0 pd=0 as=2.55625e+07 ps=89300 
M1277 Vdd xx_op_T5_jsr xx_op_T5_jsr GND dfet w=846 l=1692
+ ad=0 pd=0 as=6.65351e+06 ps=18236 
M1278 Vdd op_T2_jmp_abs op_T2_jmp_abs GND dfet w=846 l=1786
+ ad=0 pd=0 as=6.64467e+06 ps=18236 
M1279 Vdd op_T5_rti_rts op_T5_rti_rts GND dfet w=893 l=1833
+ ad=0 pd=0 as=7.30737e+06 ps=21432 
M1280 Vdd op_lsr_ror_dec_inc op_lsr_ror_dec_inc GND dfet w=846 l=1786
+ ad=0 pd=0 as=6.5033e+06 ps=17860 
M1281 Vdd x_op_T3_plp_pla x_op_T3_plp_pla GND dfet w=846 l=1786
+ ad=0 pd=0 as=6.90092e+06 ps=20680 
M1282 Vdd op_T0_cli_sei op_T0_cli_sei GND dfet w=846 l=1786
+ ad=0 pd=0 as=6.14986e+06 ps=18236 
M1283 GND _t5 op_T5_brk GND efet w=1410 l=564
+ ad=0 pd=0 as=2.0906e+07 ps=55460 
M1284 GND _t5 op_T5_rti GND efet w=1410 l=564
+ ad=0 pd=0 as=1.82375e+07 ps=48880 
M1285 op_T2_abs_access op_push_pull GND GND efet w=1316 l=564
+ ad=8.55325e+06 pd=22372 as=0 ps=0 
M1286 op_T3_abs_idx_ind op_push_pull GND GND efet w=1269 l=611
+ ad=9.57822e+06 pd=24628 as=0 ps=0 
M1287 Vdd op_asl_rol op_asl_rol GND dfet w=846 l=1786
+ ad=0 pd=0 as=1.2715e+07 ps=40796 
M1288 Vdd op_T__bit op_T__bit GND dfet w=846 l=1786
+ ad=0 pd=0 as=2.90439e+07 ps=100392 
M1289 Vdd n_1363 n_1363 GND dfet w=893 l=1833
+ ad=0 pd=0 as=3.9762e+06 ps=10340 
M1290 Vdd op_T3_mem_zp_idx op_T3_mem_zp_idx GND dfet w=940 l=1786
+ ad=0 pd=0 as=8.18214e+06 ps=22560 
M1291 Vdd op_T0_clc_sec op_T0_clc_sec GND dfet w=846 l=1786
+ ad=0 pd=0 as=1.59401e+07 ps=52076 
M1292 Vdd x_op_T0_bit x_op_T0_bit GND dfet w=846 l=1786
+ ad=0 pd=0 as=1.62582e+07 ps=53956 
M1293 Vdd x_op_T__adc_sbc x_op_T__adc_sbc GND dfet w=940 l=1786
+ ad=0 pd=0 as=3.09967e+07 ps=108100 
M1294 Vdd x_op_T4_rti x_op_T4_rti GND dfet w=846 l=1786
+ ad=0 pd=0 as=7.40457e+06 ps=20304 
M1295 Vdd op_T0_plp op_T0_plp GND dfet w=846 l=1786
+ ad=0 pd=0 as=7.09531e+06 ps=21244 
M1296 Vdd op_T__cpx_cpy_abs op_T__cpx_cpy_abs GND dfet w=846 l=1786
+ ad=0 pd=0 as=5.61086e+06 ps=16544 
M1297 Vdd op_T__cmp op_T__cmp GND dfet w=940 l=1786
+ ad=0 pd=0 as=6.5033e+06 ps=20680 
M1298 Vdd op_T__cpx_cpy_imm_zp op_T__cpx_cpy_imm_zp GND dfet w=846 l=1786
+ ad=0 pd=0 as=6.41494e+06 ps=18988 
M1299 Vdd op_T0_cld_sed op_T0_cld_sed GND dfet w=846 l=1786
+ ad=0 pd=0 as=6.44144e+06 ps=17860 
M1300 Vdd op_T3_mem_abs op_T3_mem_abs GND dfet w=846 l=1786
+ ad=0 pd=0 as=8.30584e+06 ps=22184 
M1301 Vdd op_T__asl_rol_a op_T__asl_rol_a GND dfet w=846 l=1692
+ ad=0 pd=0 as=6.90975e+06 ps=22748 
M1302 Vdd x_op_push_pull x_op_push_pull GND dfet w=940 l=1880
+ ad=0 pd=0 as=1.50654e+07 ps=54332 
M1303 Vdd nop_branch_bit6 nop_branch_bit6 GND dfet w=940 l=1880
+ ad=0 pd=0 as=4.58147e+07 ps=155852 
M1304 Vdd op_T5_mem_ind_idx op_T5_mem_ind_idx GND dfet w=846 l=1692
+ ad=0 pd=0 as=8.35002e+06 ps=23124 
M1305 Vdd nop_branch_bit7 nop_branch_bit7 GND dfet w=940 l=1410
+ ad=0 pd=0 as=4.58677e+07 ps=154912 
M1306 Vdd op_T2_mem_zp op_T2_mem_zp GND dfet w=940 l=1880
+ ad=0 pd=0 as=8.03192e+06 ps=25944 
M1307 Vdd op_T4_mem_abs_idx op_T4_mem_abs_idx GND dfet w=940 l=1786
+ ad=0 pd=0 as=8.16446e+06 ps=23500 
M1308 Vdd op_implied op_implied GND dfet w=846 l=1692
+ ad=0 pd=0 as=1.29978e+07 ps=41548 
M1309 Vdd op_clv op_clv GND dfet w=987 l=1833
+ ad=0 pd=0 as=2.3168e+07 ps=76140 
M1310 n_1696 n_400 Vdd GND dfet w=1880 l=564
+ ad=1.49593e+07 pd=35344 as=0 ps=0 
M1311 GND n_834 n_1696 GND efet w=13254 l=658
+ ad=0 pd=0 as=0 ps=0 
M1312 Vdd n_834 n_834 GND dfet w=940 l=1128
+ ad=0 pd=0 as=2.08088e+07 ps=63920 
M1313 n_400 n_400 Vdd GND dfet w=940 l=940
+ ad=1.50212e+07 pd=44368 as=0 ps=0 
M1314 n_402 cp1 notRnWprepad GND efet w=1222 l=658
+ ad=2.12064e+06 pd=7144 as=2.61015e+07 ps=65988 
M1315 GND _t5 op_T5_jsr GND efet w=1316 l=658
+ ad=0 pd=0 as=1.96248e+07 ps=53768 
M1316 GND _t5 op_T5_ind_y GND efet w=1316 l=658
+ ad=0 pd=0 as=1.11245e+07 ps=30268 
M1317 GND n_678 _t3 GND efet w=6439 l=611
+ ad=0 pd=0 as=8.50023e+06 ps=26320 
M1318 op_T4_rts _t4 GND GND efet w=1316 l=564
+ ad=2.06497e+07 pd=55084 as=0 ps=0 
M1319 op_T4_brk_jsr _t4 GND GND efet w=1316 l=564
+ ad=1.88649e+07 pd=52640 as=0 ps=0 
M1320 op_T4_rti _t4 GND GND efet w=1316 l=564
+ ad=1.82375e+07 pd=48880 as=0 ps=0 
M1321 op_T4_ind_y _t4 GND GND efet w=1316 l=564
+ ad=1.11687e+07 pd=30268 as=0 ps=0 
M1322 op_T4_ind_x _t4 GND GND efet w=1410 l=564
+ ad=1.44734e+07 pd=39480 as=0 ps=0 
M1323 GND _t5 op_T5_rts GND efet w=1316 l=564
+ ad=0 pd=0 as=2.08441e+07 ps=58280 
M1324 GND _t5 op_T5_ind_x GND efet w=1316 l=564
+ ad=0 pd=0 as=1.32098e+07 ps=35908 
M1325 GND _t5 op_T5_rti_rts GND efet w=1316 l=658
+ ad=0 pd=0 as=1.85114e+07 ps=50760 
M1326 GND _t5 xx_op_T5_jsr GND efet w=1222 l=658
+ ad=0 pd=0 as=1.95011e+07 ps=53580 
M1327 op_T4_abs_idx _t4 GND GND efet w=1316 l=564
+ ad=9.83447e+06 pd=28764 as=0 ps=0 
M1328 op_T4 _t4 GND GND efet w=1316 l=564
+ ad=4.37382e+06 pd=12032 as=0 ps=0 
M1329 x_op_T4_ind_y _t4 GND GND efet w=1222 l=564
+ ad=1.23704e+07 pd=34968 as=0 ps=0 
M1330 GND _t5 op_T5_mem_ind_idx GND efet w=1222 l=658
+ ad=0 pd=0 as=1.0886e+07 ps=29892 
M1331 GND x_op_push_pull op_implied GND efet w=1974 l=658
+ ad=0 pd=0 as=1.02586e+07 ps=25944 
M1332 GND n_834 n_400 GND efet w=3384 l=658
+ ad=0 pd=0 as=3.81715e+06 ps=13724 
M1333 Vdd notir1 notir1 GND dfet w=940 l=658
+ ad=0 pd=0 as=1.81854e+08 ps=621904 
M1334 GND ir1 n_1133 GND efet w=6110 l=658
+ ad=0 pd=0 as=1.0453e+07 ps=28012 
M1335 n_119 cclk notir1 GND efet w=1128 l=658
+ ad=4.94816e+06 pd=14852 as=6.73303e+06 ps=19552 
M1336 notir1 ir1 GND GND efet w=5922 l=658
+ ad=0 pd=0 as=0 ps=0 
M1337 op_T4_brk _t4 GND GND efet w=1316 l=564
+ ad=2.01903e+07 pd=54520 as=0 ps=0 
M1338 op_T4_jmp _t4 GND GND efet w=1316 l=564
+ ad=1.95629e+07 pd=53392 as=0 ps=0 
M1339 x_op_T4_rti _t4 GND GND efet w=1316 l=564
+ ad=1.75306e+07 pd=47752 as=0 ps=0 
M1340 op_T4_mem_abs_idx _t4 GND GND efet w=1316 l=564
+ ad=1.03028e+07 pd=28764 as=0 ps=0 
M1341 n_1456 notRdy0 n_428 GND efet w=4418 l=658
+ ad=0 pd=0 as=1.11864e+07 ps=28012 
M1342 pipeT3out cclk n_678 GND efet w=1128 l=752
+ ad=1.9881e+06 pd=7520 as=1.42613e+07 ps=39480 
M1343 _t3 _t3 Vdd GND dfet w=1034 l=658
+ ad=1.65375e+08 pd=559488 as=0 ps=0 
M1344 GND _t3 op_T3_ind_y GND efet w=1316 l=564
+ ad=0 pd=0 as=1.2609e+07 ps=35344 
M1345 GND _t3 op_T3_plp_pla GND efet w=1316 l=564
+ ad=0 pd=0 as=1.76632e+07 ps=46812 
M1346 n_428 n_16 n_1558 GND efet w=4841 l=611
+ ad=0 pd=0 as=8.75648e+06 ps=26132 
M1347 GND pipeT2out n_1558 GND efet w=10387 l=611
+ ad=0 pd=0 as=0 ps=0 
M1348 Vdd n_428 n_428 GND dfet w=846 l=1504
+ ad=0 pd=0 as=2.70382e+06 ps=7896 
M1349 Vdd n_678 n_678 GND dfet w=940 l=1128
+ ad=0 pd=0 as=9.82563e+06 ps=33088 
M1350 GND n_1357 n_678 GND efet w=3008 l=658
+ ad=0 pd=0 as=0 ps=0 
M1351 GND _t3 op_T3_stack_bit_jmp GND efet w=1316 l=564
+ ad=0 pd=0 as=1.12747e+07 ps=30456 
M1352 GND _t3 op_T3_ind_x GND efet w=1316 l=564
+ ad=0 pd=0 as=1.45175e+07 ps=40984 
M1353 GND _t3 op_T3_abs_idx GND efet w=1222 l=564
+ ad=0 pd=0 as=8.95087e+06 ps=24252 
M1354 op_T2_abs_y _t2 GND GND efet w=1316 l=564
+ ad=1.14515e+07 pd=30832 as=0 ps=0 
M1355 op_T2_idx_x_xy _t2 GND GND efet w=1316 l=564
+ ad=1.04353e+07 pd=29140 as=0 ps=0 
M1356 op_T2_ind_x _t2 GND GND efet w=1410 l=564
+ ad=1.50389e+07 pd=41360 as=0 ps=0 
M1357 op_T2 _t2 GND GND efet w=1504 l=564
+ ad=4.7626e+06 pd=12596 as=0 ps=0 
M1358 GND _t3 x_op_T3_ind_y GND efet w=1410 l=658
+ ad=0 pd=0 as=1.17961e+07 ps=31208 
M1359 GND _t3 op_T3_jmp GND efet w=1316 l=658
+ ad=0 pd=0 as=1.79636e+07 ps=48692 
M1360 GND _t3 op_T3_jsr GND efet w=1316 l=564
+ ad=0 pd=0 as=2.1498e+07 ps=59220 
M1361 op_T2_abs _t2 GND GND efet w=1410 l=564
+ ad=1.25471e+07 pd=35344 as=0 ps=0 
M1362 op_T2_ADL_ADD _t2 GND GND efet w=1410 l=564
+ ad=7.96124e+06 pd=22936 as=0 ps=0 
M1363 op_T2_stack _t2 GND GND efet w=1410 l=564
+ ad=1.48975e+07 pd=40984 as=0 ps=0 
M1364 op_T2_ind_y _t2 GND GND efet w=1410 l=564
+ ad=1.29182e+07 pd=34404 as=0 ps=0 
M1365 GND _t3 op_T3 GND efet w=1410 l=564
+ ad=0 pd=0 as=5.85827e+06 ps=15792 
M1366 GND _t3 op_T3_abs_idx_ind GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1367 GND _t3 x_op_T3_abs_idx GND efet w=1316 l=564
+ ad=0 pd=0 as=9.48986e+06 ps=25004 
M1368 GND _t3 op_T3_branch GND efet w=1316 l=564
+ ad=0 pd=0 as=1.2556e+07 ps=35532 
M1369 n_1133 n_1133 Vdd GND dfet w=846 l=752
+ ad=8.836e+06 pd=28764 as=0 ps=0 
M1370 op_T2_jsr _t2 GND GND efet w=1222 l=564
+ ad=1.97661e+07 pd=53956 as=0 ps=0 
M1371 op_T2_stack_access _t2 GND GND efet w=1316 l=564
+ ad=1.44115e+07 pd=40984 as=0 ps=0 
M1372 op_T2_pha _t2 GND GND efet w=1316 l=564
+ ad=1.73804e+07 pd=48504 as=0 ps=0 
M1373 op_T2_brk _t2 GND GND efet w=1316 l=564
+ ad=1.94304e+07 pd=53392 as=0 ps=0 
M1374 op_T2_branch _t2 GND GND efet w=1316 l=564
+ ad=1.23527e+07 pd=33464 as=0 ps=0 
M1375 op_T2_zp_zp_idx _t2 GND GND efet w=1316 l=564
+ ad=8.81833e+06 pd=24064 as=0 ps=0 
M1376 GND _t3 x_op_T3_plp_pla GND efet w=1410 l=564
+ ad=0 pd=0 as=1.69121e+07 ps=47188 
M1377 GND _t3 op_T3_mem_zp_idx GND efet w=1457 l=611
+ ad=0 pd=0 as=9.48986e+06 ps=25192 
M1378 n_678 n_644 GND GND efet w=5734 l=564
+ ad=0 pd=0 as=0 ps=0 
M1379 n_644 cp1 n_428 GND efet w=1222 l=846
+ ad=2.18249e+06 pd=9588 as=0 ps=0 
M1380 GND n_1575 _t2 GND efet w=7191 l=611
+ ad=0 pd=0 as=8.12912e+06 ps=21432 
M1381 GND pipeT2out n_12 GND efet w=11656 l=658
+ ad=0 pd=0 as=5.1779e+06 ps=20868 
M1382 n_1575 cclk pipeT2out GND efet w=1128 l=752
+ ad=9.38383e+06 pd=28200 as=2.82752e+06 ps=8648 
M1383 _t2 _t2 Vdd GND dfet w=940 l=658
+ ad=1.64102e+08 pd=582048 as=0 ps=0 
M1384 op_T2_ind _t2 GND GND efet w=1316 l=564
+ ad=1.11334e+07 pd=30268 as=0 ps=0 
M1385 op_T2_abs_access _t2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1386 GND _t3 op_T3_mem_abs GND efet w=1316 l=658
+ ad=0 pd=0 as=1.14338e+07 ps=30644 
M1387 GND ir0 op_implied GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1388 GND n_1133 irline3 GND efet w=7896 l=658
+ ad=0 pd=0 as=7.88171e+06 ps=22372 
M1389 n_1133 ir0 GND GND efet w=6627 l=517
+ ad=0 pd=0 as=0 ps=0 
M1390 ir1 ir1 Vdd GND dfet w=1034 l=1128
+ ad=1.44115e+07 pd=42864 as=0 ps=0 
M1391 GND n_119 ir1 GND efet w=7285 l=705
+ ad=0 pd=0 as=7.05113e+06 ps=22936 
M1392 n_237 fetch n_119 GND efet w=2068 l=752
+ ad=971960 pd=5076 as=0 ps=0 
M1393 n_1641 cp1 n_237 GND efet w=2068 l=658
+ ad=9.48986e+06 pd=28388 as=0 ps=0 
M1394 op_T2_php _t2 GND GND efet w=1316 l=564
+ ad=1.93773e+07 pd=52264 as=0 ps=0 
M1395 op_T2_php_pha _t2 GND GND efet w=1316 l=564
+ ad=1.57281e+07 pd=42488 as=0 ps=0 
M1396 op_T2_jmp_abs _t2 GND GND efet w=1316 l=564
+ ad=1.85909e+07 pd=49256 as=0 ps=0 
M1397 op_T2_mem_zp _t2 GND GND efet w=1410 l=564
+ ad=1.21848e+07 pd=34592 as=0 ps=0 
M1398 ir0 ir0 Vdd GND dfet w=940 l=1034
+ ad=2.62871e+07 pd=88736 as=0 ps=0 
M1399 ir0 n_310 GND GND efet w=6580 l=752
+ ad=8.72997e+06 pd=21056 as=0 ps=0 
M1400 irline3 irline3 Vdd GND dfet w=1222 l=564
+ ad=1.65702e+08 pd=589944 as=0 ps=0 
M1401 n_724 fetch n_310 GND efet w=2162 l=752
+ ad=1.01614e+06 pd=5264 as=4.55938e+06 ps=14288 
M1402 n_409 cp1 n_724 GND efet w=2162 l=658
+ ad=1.08329e+07 pd=25756 as=0 ps=0 
M1403 GND ir0 notir0 GND efet w=6204 l=658
+ ad=0 pd=0 as=8.44722e+06 ps=24252 
M1404 GND notir1 op_xy GND efet w=1316 l=564
+ ad=0 pd=0 as=9.04806e+06 ps=24440 
M1405 GND notir1 x_op_T0_txa GND efet w=1316 l=564
+ ad=0 pd=0 as=1.66028e+07 ps=43616 
M1406 GND notir1 op_T0_dex GND efet w=1316 l=564
+ ad=0 pd=0 as=1.54895e+07 ps=42488 
M1407 GND notir1 op_from_x GND efet w=1316 l=564
+ ad=0 pd=0 as=1.169e+07 ps=33840 
M1408 GND notir1 op_T0_txs GND efet w=1410 l=564
+ ad=0 pd=0 as=1.85909e+07 ps=49820 
M1409 GND notir1 op_T0_ldx_tax_tsx GND efet w=1316 l=564
+ ad=0 pd=0 as=1.25294e+07 ps=35156 
M1410 GND notir1 op_T__dex GND efet w=1410 l=564
+ ad=0 pd=0 as=1.44204e+07 ps=39480 
M1411 GND notir1 op_T0_tsx GND efet w=1504 l=564
+ ad=0 pd=0 as=1.66824e+07 ps=43804 
M1412 GND notir1 op_ror GND efet w=1316 l=564
+ ad=0 pd=0 as=1.27857e+07 ps=35532 
M1413 op_sty_cpy_mem irline3 GND GND efet w=1316 l=564
+ ad=1.15398e+07 pd=30832 as=0 ps=0 
M1414 op_T0_iny_dey irline3 GND GND efet w=1316 l=564
+ ad=1.50831e+07 pd=41360 as=0 ps=0 
M1415 x_op_T0_tya irline3 GND GND efet w=1316 l=564
+ ad=1.89621e+07 pd=49820 as=0 ps=0 
M1416 op_T0_cpy_iny irline3 GND GND efet w=1316 l=564
+ ad=1.31303e+07 pd=35720 as=0 ps=0 
M1417 op_T0_cpx_inx irline3 GND GND efet w=1316 l=564
+ ad=1.23085e+07 pd=31960 as=0 ps=0 
M1418 GND notir1 op_inc_nop GND efet w=1316 l=658
+ ad=0 pd=0 as=1.11334e+07 ps=30080 
M1419 GND notir1 op_rol_ror GND efet w=1222 l=564
+ ad=0 pd=0 as=1.1743e+07 ps=32900 
M1420 GND notir1 op_shift GND efet w=1410 l=564
+ ad=0 pd=0 as=1.00819e+07 ps=28576 
M1421 GND notir1 op_T__shift_a GND efet w=1316 l=564
+ ad=0 pd=0 as=1.52509e+07 ps=42676 
M1422 GND notir1 op_T0_txa GND efet w=1316 l=564
+ ad=0 pd=0 as=1.61699e+07 ps=43240 
M1423 op_T__inx irline3 GND GND efet w=1410 l=564
+ ad=1.76101e+07 pd=48880 as=0 ps=0 
M1424 op_T__iny_dey irline3 GND GND efet w=1316 l=564
+ ad=1.60462e+07 pd=44368 as=0 ps=0 
M1425 op_T0_ldy_mem irline3 GND GND efet w=1222 l=564
+ ad=1.18579e+07 pd=31396 as=0 ps=0 
M1426 op_T0_tay_ldy_not_idx irline3 GND GND efet w=1316 l=564
+ ad=1.31038e+07 pd=36096 as=0 ps=0 
M1427 op_T0_jsr irline3 GND GND efet w=1316 l=564
+ ad=2.00666e+07 pd=54332 as=0 ps=0 
M1428 op_T5_brk irline3 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1429 op_T0_php_pha irline3 GND GND efet w=1410 l=564
+ ad=1.76985e+07 pd=48128 as=0 ps=0 
M1430 op_T4_rts irline3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1431 op_T3_plp_pla irline3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1432 op_T5_rti irline3 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1433 op_jmp irline3 GND GND efet w=1316 l=564
+ ad=1.64526e+07 pd=43428 as=0 ps=0 
M1434 op_T2_stack irline3 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1435 op_T3_stack_bit_jmp irline3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1436 op_T4_brk_jsr irline3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1437 op_T4_rti irline3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1438 op_plp_pla irline3 GND GND efet w=1316 l=564
+ ad=1.45087e+07 pd=40608 as=0 ps=0 
M1439 GND notir1 op_T0_shift_a GND efet w=1316 l=564
+ ad=0 pd=0 as=1.51449e+07 ps=41924 
M1440 GND notir1 op_T0_tax GND efet w=1316 l=564
+ ad=0 pd=0 as=1.36781e+07 ps=36848 
M1441 GND notir1 op_T0_shift_right_a GND efet w=1316 l=564
+ ad=0 pd=0 as=1.60727e+07 ps=43052 
M1442 GND notir1 op_shift_right GND efet w=1316 l=564
+ ad=0 pd=0 as=1.05502e+07 ps=29704 
M1443 op_rti_rts irline3 GND GND efet w=1316 l=564
+ ad=1.70093e+07 pd=47188 as=0 ps=0 
M1444 op_T2_jsr irline3 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1445 op_T0_cpx_cpy_inx_iny irline3 GND GND efet w=1316 l=564
+ ad=1.27062e+07 pd=35720 as=0 ps=0 
M1446 op_T3_jmp irline3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1447 op_T5_jsr irline3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1448 op_T2_stack_access irline3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1449 op_T0_tya irline3 GND GND efet w=1316 l=564
+ ad=1.80078e+07 pd=48692 as=0 ps=0 
M1450 op_T0_pla irline3 GND GND efet w=1410 l=564
+ ad=1.74511e+07 pd=48128 as=0 ps=0 
M1451 GND notir1 op_lsr_ror_dec_inc GND efet w=1316 l=658
+ ad=0 pd=0 as=6.46795e+06 ps=17860 
M1452 GND notir1 op_asl_rol GND efet w=1316 l=658
+ ad=0 pd=0 as=9.83447e+06 ps=28576 
M1453 GND notir1 op_T__asl_rol_a GND efet w=1316 l=564
+ ad=0 pd=0 as=1.69209e+07 ps=47564 
M1454 op_T0_tay irline3 GND GND efet w=1316 l=564
+ ad=1.36163e+07 pd=36848 as=0 ps=0 
M1455 op_T0_bit irline3 GND GND efet w=1316 l=564
+ ad=1.51184e+07 pd=42112 as=0 ps=0 
M1456 op_branch_done irline3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1457 op_T2_pha irline3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1458 op_T2_brk irline3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1459 op_T3_jsr irline3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1460 op_T2_branch irline3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1461 op_T5_rts irline3 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1462 op_T0_brk_rti irline3 GND GND efet w=1316 l=564
+ ad=1.68944e+07 pd=47188 as=0 ps=0 
M1463 op_T0_jmp irline3 GND GND efet w=1316 l=564
+ ad=1.94392e+07 pd=53768 as=0 ps=0 
M1464 op_T3_branch irline3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1465 op_brk_rti irline3 GND GND efet w=1410 l=564
+ ad=1.56662e+07 pd=42300 as=0 ps=0 
M1466 op_jsr irline3 GND GND efet w=1410 l=564
+ ad=1.89002e+07 pd=52828 as=0 ps=0 
M1467 x_op_jmp irline3 GND GND efet w=1316 l=564
+ ad=1.60462e+07 pd=42864 as=0 ps=0 
M1468 op_push_pull irline3 GND GND efet w=1316 l=564
+ ad=1.22997e+07 pd=33464 as=0 ps=0 
M1469 notir0 notir0 Vdd GND dfet w=940 l=658
+ ad=1.7695e+08 pd=599344 as=0 ps=0 
M1470 op_T4_brk irline3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1471 op_T2_php irline3 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1472 op_T2_php_pha irline3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1473 op_T4_jmp irline3 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1474 op_T5_rti_rts irline3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1475 xx_op_T5_jsr irline3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1476 op_T2_jmp_abs irline3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1477 x_op_T3_plp_pla irline3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1478 op_T0_cli_sei irline3 GND GND efet w=1316 l=564
+ ad=1.5622e+07 pd=42300 as=0 ps=0 
M1479 op_T__bit irline3 GND GND efet w=1316 l=564
+ ad=1.73097e+07 pd=50008 as=0 ps=0 
M1480 op_T0_clc_sec irline3 GND GND efet w=1316 l=564
+ ad=1.67796e+07 pd=46812 as=0 ps=0 
M1481 x_op_T0_bit irline3 GND GND efet w=1316 l=564
+ ad=1.37046e+07 pd=36660 as=0 ps=0 
M1482 op_T0_plp irline3 GND GND efet w=1222 l=564
+ ad=1.68237e+07 pd=47564 as=0 ps=0 
M1483 x_op_T4_rti irline3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1484 op_T__cpx_cpy_abs irline3 GND GND efet w=1410 l=564
+ ad=1.64261e+07 pd=45684 as=0 ps=0 
M1485 op_T__cpx_cpy_imm_zp irline3 GND GND efet w=1410 l=564
+ ad=1.46413e+07 pd=39856 as=0 ps=0 
M1486 x_op_push_pull irline3 GND GND efet w=1316 l=564
+ ad=1.24499e+07 pd=34216 as=0 ps=0 
M1487 op_T0_cld_sed irline3 GND GND efet w=1316 l=564
+ ad=1.60373e+07 pd=42864 as=0 ps=0 
M1488 op_clv irline3 GND GND efet w=1222 l=564
+ ad=1.71949e+07 pd=45684 as=0 ps=0 
M1489 n_310 cclk notir0 GND efet w=1222 l=658
+ ad=0 pd=0 as=0 ps=0 
M1490 GND notir0 op_T3_ind_y GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1491 GND notir0 op_T2_abs_y GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1492 n_1575 n_1575 Vdd GND dfet w=940 l=1128
+ ad=1.00907e+07 pd=35344 as=0 ps=0 
M1493 GND notir0 op_T2_ind_x GND efet w=1410 l=658
+ ad=0 pd=0 as=0 ps=0 
M1494 GND notir0 op_T0_eor GND efet w=1410 l=564
+ ad=0 pd=0 as=1.1045e+07 ps=30080 
M1495 GND notir0 op_T0_ora GND efet w=1316 l=564
+ ad=0 pd=0 as=1.16193e+07 ps=31020 
M1496 GND notir0 op_T3_ind_x GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1497 GND notir0 op_T4_ind_y GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1498 GND notir0 op_T2_ind_y GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1499 GND notir0 op_T4_ind_x GND efet w=1363 l=611
+ ad=0 pd=0 as=0 ps=0 
M1500 GND n_1357 n_1575 GND efet w=4418 l=658
+ ad=0 pd=0 as=0 ps=0 
M1501 op_T0_jsr ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1502 op_T5_brk ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1503 op_T0_php_pha ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1504 op_T4_rts ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1505 op_T3_plp_pla ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1506 op_T5_rti ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1507 op_ror ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1508 GND notir0 x_op_T3_ind_y GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1509 GND notir0 op_T0_cmp GND efet w=1316 l=658
+ ad=0 pd=0 as=1.16812e+07 ps=31020 
M1510 GND notir0 op_T0_sbc GND efet w=1316 l=658
+ ad=0 pd=0 as=1.24588e+07 ps=35156 
M1511 GND notir0 op_T0_adc_sbc GND efet w=1316 l=658
+ ad=0 pd=0 as=9.61357e+06 ps=25192 
M1512 GND notir0 op_T__ora_and_eor_adc GND efet w=1316 l=658
+ ad=0 pd=0 as=8.33235e+06 ps=25568 
M1513 GND notir0 op_T__adc_sbc GND efet w=1316 l=658
+ ad=0 pd=0 as=1.12924e+07 ps=31396 
M1514 GND notir0 op_T0_lda GND efet w=1410 l=564
+ ad=0 pd=0 as=1.11687e+07 ps=30268 
M1515 GND notir0 op_T0_acc GND efet w=1222 l=564
+ ad=0 pd=0 as=7.90822e+06 ps=23312 
M1516 GND notir0 op_T0_and GND efet w=1316 l=564
+ ad=0 pd=0 as=9.13642e+06 ps=24628 
M1517 GND notir0 op_T5_ind_y GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1518 GND notir0 op_sta_cmp GND efet w=1222 l=564
+ ad=0 pd=0 as=1.11775e+07 ps=30268 
M1519 op_T0_eor ir7 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1520 op_jmp ir7 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1521 op_T0_ora ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1522 op_T2_stack ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1523 op_T3_stack_bit_jmp ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1524 op_T4_brk_jsr ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1525 op_T4_rti ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1526 op_plp_pla ir7 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1527 op_rti_rts ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1528 op_T2_jsr ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1529 op_rol_ror ir7 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1530 op_T3_jmp ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1531 op_shift ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1532 op_T5_jsr ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1533 op_T2_stack_access ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1534 op_T__ora_and_eor_adc ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1535 op_T__shift_a ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1536 op_T0_pla ir7 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1537 GND notir0 op_T2_ind GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1538 GND notir0 op_T5_ind_x GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1539 GND notir0 x_op_T4_ind_y GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1540 op_T0_shift_a ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1541 op_T0_bit ir7 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1542 op_T0_and ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1543 op_T2_pha ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1544 op_T0_shift_right_a ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1545 op_shift_right ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1546 op_T2_brk ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1547 op_T3_jsr ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1548 GND notir0 x_op_T__adc_sbc GND efet w=1410 l=658
+ ad=0 pd=0 as=1.96159e+07 ps=55460 
M1549 GND notir0 op_T__cmp GND efet w=1222 l=658
+ ad=0 pd=0 as=1.26532e+07 ps=36284 
M1550 GND notir0 op_T5_mem_ind_idx GND efet w=1363 l=611
+ ad=0 pd=0 as=0 ps=0 
M1551 op_T5_rts ir7 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1552 op_T0_brk_rti ir7 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1553 op_T0_jmp ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1554 op_brk_rti ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1555 op_jsr ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1556 x_op_jmp ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1557 op_push_pull ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1558 op_T4_brk ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1559 op_T2_php ir7 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1560 op_T2_php_pha ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1561 op_T4_jmp ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1562 op_T5_rti_rts ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1563 xx_op_T5_jsr ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1564 op_T2_jmp_abs ir7 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1565 x_op_T3_plp_pla ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1566 op_asl_rol ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1567 op_T0_cli_sei ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1568 op_T__bit ir7 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1569 op_T0_clc_sec ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1570 ir7 ir7 Vdd GND dfet w=940 l=564
+ ad=1.76199e+08 pd=624536 as=0 ps=0 
M1571 GND n_541 ir7 GND efet w=11374 l=564
+ ad=0 pd=0 as=1.10627e+07 ps=27824 
M1572 notir7 notir7 Vdd GND dfet w=940 l=658
+ ad=1.70473e+08 pd=576596 as=0 ps=0 
M1573 GND ir7 notir7 GND efet w=8366 l=564
+ ad=0 pd=0 as=1.58783e+07 ps=37976 
M1574 n_1183 fetch n_541 GND efet w=2068 l=752
+ ad=971960 pd=5076 as=4.13525e+06 ps=10528 
M1575 n_1605 cp1 n_1183 GND efet w=2068 l=752
+ ad=1.08506e+07 pd=25380 as=0 ps=0 
M1576 n_541 cclk notir7 GND efet w=1128 l=752
+ ad=0 pd=0 as=0 ps=0 
M1577 n_12 notRdy0 n_1091 GND efet w=4794 l=752
+ ad=0 pd=0 as=9.5959e+06 ps=22936 
M1578 x_op_T0_bit ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1579 op_T0_plp ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1580 x_op_T4_rti ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1581 op_T__asl_rol_a ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1582 x_op_push_pull ir7 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1583 nop_branch_bit7 ir7 GND GND efet w=2914 l=564
+ ad=5.85827e+06 pd=15604 as=0 ps=0 
M1584 n_1575 n_1360 GND GND efet w=6862 l=658
+ ad=0 pd=0 as=0 ps=0 
M1585 n_1091 n_16 n_363 GND efet w=4841 l=611
+ ad=0 pd=0 as=8.7388e+06 ps=24064 
M1586 n_1360 cp1 n_1091 GND efet w=1128 l=658
+ ad=1.47561e+06 pd=6956 as=0 ps=0 
M1587 GND notir7 op_sty_cpy_mem GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1588 GND notir7 op_T0_iny_dey GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1589 GND notir7 x_op_T0_tya GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1590 GND notir7 op_T0_cpy_iny GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1591 GND notir7 op_xy GND efet w=1410 l=658
+ ad=0 pd=0 as=0 ps=0 
M1592 GND notir7 x_op_T0_txa GND efet w=1410 l=658
+ ad=0 pd=0 as=0 ps=0 
M1593 GND notir7 op_T0_dex GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1594 GND notir7 op_T0_cpx_inx GND efet w=1410 l=658
+ ad=0 pd=0 as=0 ps=0 
M1595 GND notir7 op_from_x GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1596 GND notir7 op_T0_txs GND efet w=1551 l=611
+ ad=0 pd=0 as=0 ps=0 
M1597 GND notir7 op_T0_ldx_tax_tsx GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1598 GND notir7 op_T__dex GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1599 GND notir7 op_T__inx GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1600 GND notir7 op_T0_tsx GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1601 GND notir7 op_T__iny_dey GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1602 GND notir7 op_T0_ldy_mem GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1603 GND notir7 op_T0_tay_ldy_not_idx GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1604 GND pipeT_SYNC n_363 GND efet w=11280 l=564
+ ad=0 pd=0 as=0 ps=0 
M1605 Vdd n_1091 n_1091 GND dfet w=940 l=1504
+ ad=0 pd=0 as=2.88054e+06 ps=7896 
M1606 op_T0_iny_dey ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1607 op_T0_cpy_iny ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1608 op_T2_ind_x ir4 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1609 x_op_T0_txa ir4 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1610 op_T0_dex ir4 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1611 op_T0_cpx_inx ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1612 GND notir7 op_inc_nop GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1613 op_T__dex ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1614 op_T__inx ir4 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1615 op_T__iny_dey ir4 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1616 op_T0_tay_ldy_not_idx ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1617 op_T0_jsr ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1618 op_T5_brk ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1619 op_T0_php_pha ir4 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1620 op_T4_rts ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1621 op_T3_plp_pla ir4 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1622 op_T5_rti ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1623 op_jmp ir4 GND GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1624 op_T2_abs ir4 GND GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1625 op_T2_stack ir4 GND GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1626 op_T3_stack_bit_jmp ir4 GND GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1627 GND notir7 op_T0_cpx_cpy_inx_iny GND efet w=1410 l=658
+ ad=0 pd=0 as=0 ps=0 
M1628 GND notir7 op_T0_cmp GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1629 GND notir7 op_T0_sbc GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1630 GND notir7 op_T0_tya GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1631 GND notir7 op_T0_txa GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1632 GND notir7 op_T0_lda GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1633 GND notir7 op_T0_tay GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1634 GND notir7 op_T0_tax GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1635 GND notir7 op_sta_cmp GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1636 op_T4_brk_jsr ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1637 op_T4_rti ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1638 op_T3_ind_x ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1639 op_plp_pla ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1640 op_T4_ind_x ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1641 op_rti_rts ir4 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1642 op_T2_jsr ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1643 op_T0_cpx_cpy_inx_iny ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1644 op_T3_jmp ir4 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1645 op_T5_jsr ir4 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1646 op_T2_stack_access ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1647 op_T__shift_a ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1648 op_T0_txa ir4 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1649 op_T0_pla ir4 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1650 GND notir7 op_store GND efet w=1316 l=564
+ ad=0 pd=0 as=9.45452e+06 ps=26884 
M1651 n_862 cclk pipeT_SYNC GND efet w=1128 l=658
+ ad=1.61964e+07 pd=49820 as=1.67884e+06 ps=7144 
M1652 op_T0_tay ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1653 op_T0_shift_a ir4 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1654 op_T0_tax ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1655 op_T0_bit ir4 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1656 op_T2_pha ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1657 op_T0_shift_right_a ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1658 op_T2_brk ir4 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1659 op_T3_jsr ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1660 GND notir7 op_T__cmp GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1661 GND notir7 op_T__cpx_cpy_abs GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1662 GND notir7 op_T__cpx_cpy_imm_zp GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1663 GND notir7 op_T0_cld_sed GND efet w=1410 l=658
+ ad=0 pd=0 as=0 ps=0 
M1664 GND notir7 op_clv GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1665 op_T5_rts ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1666 op_T0_brk_rti ir4 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1667 op_T0_jmp ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1668 op_T5_ind_x ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1669 op_brk_rti ir4 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1670 op_jsr ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1671 x_op_jmp ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1672 op_push_pull ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1673 op_T4_brk ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1674 op_T2_php ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1675 op_T2_php_pha ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1676 op_T4_jmp ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1677 op_T5_rti_rts ir4 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1678 xx_op_T5_jsr ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1679 op_T2_jmp_abs ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1680 x_op_T3_plp_pla ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1681 op_T__bit ir4 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1682 ir4 ir4 Vdd GND dfet w=940 l=658
+ ad=1.7854e+08 pd=624724 as=0 ps=0 
M1683 GND n_927 ir4 GND efet w=11515 l=611
+ ad=0 pd=0 as=9.79912e+06 ps=26696 
M1684 x_op_T0_bit ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1685 op_T0_plp ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1686 x_op_T4_rti ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1687 op_T__cpx_cpy_abs ir4 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1688 op_T__asl_rol_a ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1689 op_T__cpx_cpy_imm_zp ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1690 x_op_push_pull ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1691 op_T3_mem_abs ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1692 op_T2_mem_zp ir4 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1693 notir4 notir4 Vdd GND dfet w=940 l=564
+ ad=1.67486e+08 pd=568136 as=0 ps=0 
M1694 GND ir4 notir4 GND efet w=8131 l=611
+ ad=0 pd=0 as=1.7619e+07 ps=38916 
M1695 n_703 fetch n_927 GND efet w=2256 l=752
+ ad=1.06032e+06 pd=5452 as=4.04689e+06 ps=10152 
M1696 n_227 cp1 n_703 GND efet w=2256 l=752
+ ad=1.14338e+07 pd=27072 as=0 ps=0 
M1697 n_927 cclk notir4 GND efet w=1128 l=658
+ ad=0 pd=0 as=0 ps=0 
M1698 GND notir4 op_T3_ind_y GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1699 GND notir4 op_T2_abs_y GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1700 GND notir4 x_op_T0_tya GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1701 GND notir4 op_T2_idx_x_xy GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1702 GND notir4 op_T0_txs GND efet w=1504 l=564
+ ad=0 pd=0 as=0 ps=0 
M1703 n_1368 NMIL GND GND efet w=4841 l=611
+ ad=1.54983e+07 pd=45684 as=0 ps=0 
M1704 GND n_562 NMIL GND efet w=6251 l=611
+ ad=0 pd=0 as=1.01349e+07 ps=30268 
M1705 NMIL NMIL Vdd GND dfet w=940 l=1316
+ ad=1.24146e+07 pd=40420 as=0 ps=0 
M1706 GND notRdy0 n_16 GND efet w=5217 l=611
+ ad=0 pd=0 as=6.88324e+06 ps=15792 
M1707 Vdd n_16 n_16 GND dfet w=940 l=940
+ ad=0 pd=0 as=2.32387e+07 ps=77080 
M1708 NMIL n_882 GND GND efet w=3290 l=658
+ ad=0 pd=0 as=0 ps=0 
M1709 n_562 cp1 n_645 GND efet w=1128 l=846
+ ad=2.26202e+06 pd=8460 as=0 ps=0 
M1710 GND n_645 n_1368 GND efet w=3384 l=658
+ ad=0 pd=0 as=0 ps=0 
M1711 n_1368 n_1578 GND GND efet w=4183 l=705
+ ad=0 pd=0 as=0 ps=0 
M1712 Vdd n_1368 n_1368 GND dfet w=940 l=940
+ ad=0 pd=0 as=2.16924e+07 ps=76892 
M1713 NMIL cclk n_1252 GND efet w=1222 l=658
+ ad=0 pd=0 as=3.02191e+06 ps=8836 
M1714 n_1578 pipenVEC GND GND efet w=5640 l=752
+ ad=4.58588e+06 pd=12032 as=0 ps=0 
M1715 Vdd n_1578 n_1578 GND dfet w=1034 l=1598
+ ad=0 pd=0 as=7.05113e+06 ps=19740 
M1716 n_882 n_1252 GND GND efet w=5123 l=705
+ ad=8.84484e+06 pd=26696 as=0 ps=0 
M1717 GND notir4 op_T0_tsx GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1718 GND notir4 op_T4_ind_y GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1719 GND notir4 op_T2_ind_y GND efet w=1410 l=658
+ ad=0 pd=0 as=0 ps=0 
M1720 GND notir4 op_T3_abs_idx GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1721 GND notir4 x_op_T3_ind_y GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1722 GND notir4 op_T0_tya GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1723 op_T3_ind_y ir3 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1724 op_T2_ind_x ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1725 op_T0_jsr ir3 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1726 op_T5_brk ir3 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1727 op_T4_rts ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1728 op_T5_rti ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1729 op_T2_ADL_ADD ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1730 op_T4_brk_jsr ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1731 op_T4_rti ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1732 op_T3_ind_x ir3 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1733 op_T4_ind_y ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1734 op_T2_ind_y ir3 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1735 op_T4_ind_x ir3 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1736 GND notir4 op_T4_abs_idx GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1737 GND notir4 op_T5_ind_y GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1738 GND notir4 op_branch_done GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1739 GND notir4 op_T2_branch GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1740 GND notir4 x_op_T4_ind_y GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1741 GND notir4 x_op_T3_abs_idx GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1742 GND notir4 op_T3_branch GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1743 x_op_T3_ind_y ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1744 op_rti_rts ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1745 op_T2_jsr ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1746 op_T5_jsr ir3 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1747 op_T5_ind_y ir3 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1748 op_branch_done ir3 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1749 op_T2_brk ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1750 op_T3_jsr ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1751 op_T2_branch ir3 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1752 op_T2_zp_zp_idx ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1753 GND notir4 op_T0_cli_sei GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1754 GND notir4 op_T0_clc_sec GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1755 GND notir4 op_T3_mem_zp_idx GND efet w=1363 l=611
+ ad=0 pd=0 as=0 ps=0 
M1756 GND notir4 op_T0_cld_sed GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1757 op_T2_ind ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1758 op_T5_rts ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1759 op_T0_brk_rti ir3 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1760 op_T5_ind_x ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1761 x_op_T4_ind_y ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1762 op_T3_branch ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1763 op_brk_rti ir3 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1764 op_jsr ir3 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1765 GND notir4 op_T4_mem_abs_idx GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1766 GND notir4 op_clv GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1767 ir3 ir3 Vdd GND dfet w=846 l=658
+ ad=1.76269e+08 pd=613820 as=0 ps=0 
M1768 op_T4_brk ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1769 op_T5_rti_rts ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1770 xx_op_T5_jsr ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1771 op_T3_mem_zp_idx ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1772 x_op_T4_rti ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1773 op_T__cpx_cpy_imm_zp ir3 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1774 op_T2_mem_zp ir3 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1775 op_T5_mem_ind_idx ir3 GND GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1776 GND n_1620 ir3 GND efet w=12032 l=658
+ ad=0 pd=0 as=1.14603e+07 ps=28388 
M1777 GND notir3 op_T2_abs_y GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1778 GND notir3 op_T0_iny_dey GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1779 GND notir3 x_op_T0_tya GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1780 GND notir3 x_op_T0_txa GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1781 GND notir3 op_T0_dex GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1782 GND notir3 op_T0_txs GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1783 GND notir3 op_T__dex GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1784 GND notir3 op_T__inx GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1785 GND notir3 op_T0_tsx GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1786 GND notir3 op_T__iny_dey GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1787 GND notir3 op_T0_php_pha GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1788 GND notir3 op_T3_plp_pla GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1789 GND notir3 op_jmp GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1790 GND notir3 op_T2_abs GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1791 GND notir3 op_T3_abs_idx GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1792 GND notir3 op_plp_pla GND efet w=1222 l=658
+ ad=0 pd=0 as=0 ps=0 
M1793 GND notir3 op_T3_jmp GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1794 GND notir3 op_T0_tya GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1795 GND notir3 op_T__shift_a GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1796 GND notir3 op_T0_txa GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1797 GND notir3 op_T0_pla GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1798 notir3 notir3 Vdd GND dfet w=846 l=658
+ ad=1.65507e+08 pd=564752 as=0 ps=0 
M1799 GND ir3 notir3 GND efet w=7990 l=658
+ ad=0 pd=0 as=1.5949e+07 ps=37788 
M1800 op_T3_ind_y ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1801 op_T2_abs_y ir2 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1802 op_T0_iny_dey ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1803 x_op_T0_tya ir2 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1804 op_T2_ind_x ir2 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1805 x_op_T0_txa ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1806 op_T0_dex ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1807 op_T0_txs ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1808 op_T__dex ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1809 op_T__inx ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1810 op_T0_tsx ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1811 op_T__iny_dey ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1812 op_T0_jsr ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1813 op_T5_brk ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1814 op_T0_php_pha ir2 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1815 op_T4_rts ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1816 op_T3_plp_pla ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1817 op_T5_rti ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1818 GND n_597 n_882 GND efet w=6674 l=658
+ ad=0 pd=0 as=0 ps=0 
M1819 n_882 n_882 Vdd GND dfet w=846 l=1598
+ ad=7.90822e+06 pd=23500 as=0 ps=0 
M1820 op_T2_stack ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1821 op_T4_brk_jsr ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1822 op_T4_rti ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1823 op_T3_ind_x ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1824 op_T4_ind_y ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1825 op_T2_ind_y ir2 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1826 op_plp_pla ir2 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1827 op_T4_ind_x ir2 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1828 GND notir3 op_T0_tay GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1829 GND notir3 op_T0_shift_a GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1830 GND notir3 op_T0_tax GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1831 GND notir3 op_T4_abs_idx GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1832 GND notir3 op_T2_pha GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1833 GND notir3 op_T0_shift_right_a GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1834 GND notir3 op_T2_abs_access GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1835 GND notir3 op_T0_jmp GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1836 GND notir3 op_T3_abs_idx_ind GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1837 GND notir3 x_op_T3_abs_idx GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1838 GND notir3 x_op_jmp GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1839 GND notir3 op_push_pull GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1840 x_op_T3_ind_y ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1841 op_rti_rts ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1842 op_T2_jsr ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1843 op_T5_jsr ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1844 op_T2_stack_access ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1845 op_T0_tya ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1846 op_T__shift_a ir2 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1847 op_T0_txa ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1848 op_T0_pla ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1849 op_T0_tay ir2 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1850 op_T0_shift_a ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1851 op_T0_tax ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1852 op_T5_ind_y ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1853 op_branch_done ir2 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1854 op_T2_pha ir2 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1855 op_T0_shift_right_a ir2 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1856 op_T2_brk ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1857 op_T3_jsr ir2 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1858 op_T2_branch ir2 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1859 GND notir3 op_T2_php GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1860 GND notir3 op_T2_php_pha GND efet w=1410 l=658
+ ad=0 pd=0 as=0 ps=0 
M1861 GND notir3 op_T4_jmp GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1862 GND notir3 op_T2_jmp_abs GND efet w=1410 l=658
+ ad=0 pd=0 as=0 ps=0 
M1863 GND notir3 x_op_T3_plp_pla GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1864 GND notir3 op_T0_cli_sei GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1865 GND notir3 op_T0_clc_sec GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1866 n_1590 fetch n_1620 GND efet w=2256 l=752
+ ad=1.06032e+06 pd=5452 as=4.24128e+06 ps=10528 
M1867 n_1083 cp1 n_1590 GND efet w=2256 l=752
+ ad=9.52521e+06 pd=25192 as=0 ps=0 
M1868 n_1620 cclk notir3 GND efet w=1034 l=658
+ ad=0 pd=0 as=0 ps=0 
M1869 GND notir3 op_T0_plp GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1870 GND notir3 op_T__cpx_cpy_abs GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1871 GND notir3 op_T__asl_rol_a GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1872 GND notir3 x_op_push_pull GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1873 GND notir3 op_T0_cld_sed GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1874 GND notir3 op_T3_mem_abs GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1875 GND notir3 op_T4_mem_abs_idx GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1876 GND notir3 op_clv GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1877 GND notir3 op_implied GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1878 op_T2_ind ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1879 op_T5_rts ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1880 op_T0_brk_rti ir2 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1881 op_T5_ind_x ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1882 x_op_T4_ind_y ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1883 op_T3_branch ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1884 op_brk_rti ir2 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1885 op_jsr ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1886 op_push_pull ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1887 op_T4_brk ir2 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1888 op_T2_php ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1889 op_T2_php_pha ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1890 op_T5_rti_rts ir2 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1891 xx_op_T5_jsr ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1892 x_op_T3_plp_pla ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1893 op_T0_cli_sei ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1894 op_T0_clc_sec ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1895 op_T0_plp ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1896 x_op_T4_rti ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1897 op_T__asl_rol_a ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1898 x_op_push_pull ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1899 op_T0_cld_sed ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1900 op_T5_mem_ind_idx ir2 GND GND efet w=1363 l=611
+ ad=0 pd=0 as=0 ps=0 
M1901 op_clv ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1902 op_implied ir2 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1903 ir2 ir2 Vdd GND dfet w=940 l=658
+ ad=1.73601e+08 pd=611000 as=0 ps=0 
M1904 GND notir2 op_sty_cpy_mem GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1905 GND notir2 op_T2_idx_x_xy GND efet w=1410 l=658
+ ad=0 pd=0 as=0 ps=0 
M1906 GND notir2 op_T0_ldy_mem GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1907 op_sty_cpy_mem ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1908 x_op_T0_tya ir6 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1909 op_xy ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1910 x_op_T0_txa ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1911 op_from_x ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1912 op_T0_txs ir6 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1913 GND notir2 op_jmp GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1914 GND notir2 op_T2_abs GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1915 GND notir2 op_T3_jmp GND efet w=1222 l=658
+ ad=0 pd=0 as=0 ps=0 
M1916 GND notir2 op_T0_bit GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1917 GND notir2 op_T2_zp_zp_idx GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1918 op_T0_ldx_tax_tsx ir6 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1919 op_T0_tsx ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1920 op_T0_ldy_mem ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1921 op_T0_tay_ldy_not_idx ir6 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1922 op_T0_jsr ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1923 op_T5_brk ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1924 op_T0_ora ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1925 op_T4_brk_jsr ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1926 op_rol_ror ir6 GND GND efet w=1363 l=611
+ ad=0 pd=0 as=0 ps=0 
M1927 op_T2_jsr ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1928 op_shift ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1929 op_T5_jsr ir6 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1930 op_T0_tya ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1931 op_T0_txa ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1932 op_T0_lda ir6 GND GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1933 op_T0_tay ir6 GND GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1934 op_T0_tax ir6 GND GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1935 op_T0_bit ir6 GND GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1936 op_T0_and ir6 GND GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1937 GND notir2 op_T0_jmp GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1938 GND notir2 x_op_jmp GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1939 GND notir2 op_T4_jmp GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1940 GND notir2 op_T2_jmp_abs GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1941 GND notir2 op_T__bit GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1942 GND notir2 op_T3_mem_zp_idx GND efet w=1363 l=611
+ ad=0 pd=0 as=0 ps=0 
M1943 op_T2_brk ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1944 op_T3_jsr ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1945 op_sta_cmp ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1946 op_jsr ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1947 GND notir2 x_op_T0_bit GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1948 GND notir2 op_T__cpx_cpy_abs GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1949 GND notir2 op_T3_mem_abs GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1950 GND notir2 op_T2_mem_zp GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1951 GND n_1300 ir2 GND efet w=11938 l=658
+ ad=0 pd=0 as=1.24941e+07 ps=28388 
M1952 op_store ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1953 op_T4_brk ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1954 op_T2_php ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1955 xx_op_T5_jsr ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1956 op_asl_rol ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1957 op_T__bit ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1958 op_T0_clc_sec ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1959 x_op_T0_bit ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1960 op_T0_plp ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1961 op_T__asl_rol_a ir6 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M1962 GND notir6 op_T0_cpy_iny GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1963 GND notir6 op_T0_dex GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1964 GND notir6 op_T0_cpx_inx GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1965 nop_branch_bit6 ir6 GND GND efet w=1316 l=564
+ ad=5.29276e+06 pd=16168 as=0 ps=0 
M1966 notir2 notir2 Vdd GND dfet w=940 l=658
+ ad=1.69077e+08 pd=570768 as=0 ps=0 
M1967 GND ir2 notir2 GND efet w=8178 l=658
+ ad=0 pd=0 as=1.68591e+07 ps=37976 
M1968 n_343 fetch n_1300 GND efet w=2162 l=752
+ ad=1.01614e+06 pd=5264 as=4.16176e+06 ps=10528 
M1969 n_571 cp1 n_343 GND efet w=2162 l=846
+ ad=1.16105e+07 pd=26696 as=0 ps=0 
M1970 n_1300 cclk notir2 GND efet w=1034 l=658
+ ad=0 pd=0 as=0 ps=0 
M1971 op_clv ir6 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1972 GND notir6 op_T__dex GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1973 GND notir6 op_T__inx GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1974 GND notir6 op_T4_rts GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1975 GND notir6 op_T5_rti GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1976 GND notir6 op_ror GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1977 pipenVEC cclk nVEC GND efet w=1034 l=752
+ ad=2.209e+06 pd=9024 as=9.58706e+06 ps=30832 
M1978 n_597 cp1 n_1339 GND efet w=1222 l=658
+ ad=1.33424e+06 pd=7144 as=7.00695e+06 ps=17108 
M1979 n_1368 cp1 n_1149 GND efet w=1222 l=658
+ ad=0 pd=0 as=1.5463e+06 ps=7332 
M1980 op_sty_cpy_mem ir5 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1981 op_T0_iny_dey ir5 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1982 x_op_T0_tya ir5 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1983 op_T0_cpy_iny ir5 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1984 x_op_T0_txa ir5 GND GND efet w=1410 l=658
+ ad=0 pd=0 as=0 ps=0 
M1985 op_T0_dex ir5 GND GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1986 op_from_x ir5 GND GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1987 op_T0_txs ir5 GND GND efet w=1363 l=611
+ ad=0 pd=0 as=0 ps=0 
M1988 GND notir6 op_T0_eor GND efet w=1410 l=658
+ ad=0 pd=0 as=0 ps=0 
M1989 GND notir6 op_jmp GND efet w=1410 l=658
+ ad=0 pd=0 as=0 ps=0 
M1990 GND notir6 op_T4_rti GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M1991 GND notir6 op_inc_nop GND efet w=1410 l=658
+ ad=0 pd=0 as=0 ps=0 
M1992 GND notir6 op_rti_rts GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1993 GND notir6 op_T0_cpx_cpy_inx_iny GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1994 GND notir6 op_T0_cmp GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1995 GND notir6 op_T0_sbc GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1996 GND notir6 op_T0_adc_sbc GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M1997 GND notir6 op_T3_jmp GND efet w=1363 l=611
+ ad=0 pd=0 as=0 ps=0 
M1998 GND notir6 op_T__adc_sbc GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M1999 GND notir6 op_T0_pla GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M2000 op_T__dex ir5 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M2001 op_T__iny_dey ir5 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2002 op_T5_brk ir5 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2003 op_T0_php_pha ir5 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2004 op_T5_rti ir5 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2005 GND notir6 op_T2_pha GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M2006 GND notir6 op_T0_shift_right_a GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2007 GND notir6 op_shift_right GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M2008 op_T0_eor ir5 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M2009 op_T0_ora ir5 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2010 op_T4_rti ir5 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2011 op_T0_cmp ir5 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2012 op_T0_tya ir5 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2013 op_T0_txa ir5 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2014 GND notir6 op_T5_rts GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2015 GND notir6 op_T0_jmp GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2016 GND notir6 x_op_jmp GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M2017 op_T2_pha ir5 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2018 op_T2_brk ir5 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2019 op_sta_cmp ir5 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2020 GND notir6 op_T4_jmp GND efet w=1410 l=658
+ ad=0 pd=0 as=0 ps=0 
M2021 GND notir6 op_T5_rti_rts GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M2022 GND notir6 op_T2_jmp_abs GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M2023 GND notir6 op_lsr_ror_dec_inc GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M2024 GND notir6 op_T0_cli_sei GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M2025 ir6 ir6 Vdd GND dfet w=940 l=658
+ ad=1.74299e+08 pd=612504 as=0 ps=0 
M2026 GND n_1675 ir6 GND efet w=12126 l=658
+ ad=0 pd=0 as=1.13454e+07 ps=28576 
M2027 GND notir6 x_op_T__adc_sbc GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2028 GND notir6 x_op_T4_rti GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2029 GND notir6 op_T__cmp GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2030 GND notir6 op_T__cpx_cpy_abs GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2031 GND notir6 op_T__cpx_cpy_imm_zp GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2032 GND notir6 op_T0_cld_sed GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M2033 op_T0_brk_rti ir5 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M2034 op_brk_rti ir5 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M2035 op_store ir5 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2036 op_T4_brk ir5 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2037 op_T2_php ir5 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M2038 op_T2_php_pha ir5 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2039 op_T2_jmp_abs ir5 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2040 notir6 notir6 Vdd GND dfet w=940 l=658
+ ad=1.67486e+08 pd=569828 as=0 ps=0 
M2041 GND ir6 notir6 GND efet w=8272 l=658
+ ad=0 pd=0 as=1.62317e+07 ps=39480 
M2042 x_op_T4_rti ir5 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2043 op_T__cmp ir5 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M2044 n_1339 n_1339 Vdd GND dfet w=940 l=1128
+ ad=2.91588e+06 pd=8648 as=0 ps=0 
M2045 GND n_799 n_1339 GND efet w=6721 l=705
+ ad=0 pd=0 as=0 ps=0 
M2046 nNMIG cclk n_1693 GND efet w=1222 l=658
+ ad=2.01019e+07 pd=50572 as=1.9881e+06 ps=7896 
M2047 n_799 cclk nNMIG GND efet w=1128 l=658
+ ad=1.7672e+06 pd=8084 as=0 ps=0 
M2048 GND notir5 op_T0_cpx_inx GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2049 GND n_1149 nNMIG GND efet w=10246 l=658
+ ad=0 pd=0 as=0 ps=0 
M2050 op_T0_cpy_iny clock1 GND GND efet w=1363 l=611
+ ad=0 pd=0 as=0 ps=0 
M2051 op_T0_iny_dey clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2052 x_op_T0_tya clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2053 GND notir5 op_T0_ldx_tax_tsx GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M2054 GND notir5 op_T__inx GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2055 GND notir5 op_T0_tsx GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2056 GND notir5 op_T0_ldy_mem GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2057 GND notir5 op_T0_tay_ldy_not_idx GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2058 GND notir5 op_T0_jsr GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M2059 GND notir5 op_T4_rts GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2060 GND notir5 op_T3_plp_pla GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M2061 GND notir5 op_ror GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M2062 x_op_T0_txa clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2063 op_T0_dex clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2064 op_T0_cpx_inx clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2065 op_T0_txs clock1 GND GND efet w=1504 l=564
+ ad=0 pd=0 as=0 ps=0 
M2066 op_T0_tay_ldy_not_idx clock1 GND GND efet w=1363 l=611
+ ad=0 pd=0 as=0 ps=0 
M2067 GND notir5 op_plp_pla GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2068 GND notir5 op_inc_nop GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2069 GND notir5 op_T2_jsr GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2070 GND notir5 op_T0_sbc GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2071 GND notir5 op_T0_adc_sbc GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2072 GND notir5 op_rol_ror GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M2073 op_T0_ldx_tax_tsx clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2074 op_T0_tsx clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2075 op_T0_ldy_mem clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2076 op_T0_jsr clock1 GND GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M2077 op_T0_php_pha clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2078 op_T0_eor clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2079 op_T0_ora clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2080 op_T0 clock1 GND GND efet w=1410 l=564
+ ad=4.86864e+06 pd=12784 as=0 ps=0 
M2081 GND notir5 op_T5_jsr GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M2082 GND notir5 op_T__adc_sbc GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M2083 GND notir5 op_T0_pla GND efet w=1363 l=611
+ ad=0 pd=0 as=0 ps=0 
M2084 GND notir5 op_T0_lda GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2085 GND notir5 op_T0_tay GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2086 GND notir5 op_T0_tax GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M2087 GND notir5 op_T0_bit GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2088 GND notir5 op_T0_and GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M2089 GND notir5 op_T3_jsr GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M2090 op_T0_cpx_cpy_inx_iny clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2091 op_T0_cmp clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2092 op_T0_sbc clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2093 op_T0_adc_sbc clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2094 op_T0_tya clock1 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M2095 op_T0_txa clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2096 op_T0_pla clock1 GND GND efet w=1269 l=611
+ ad=0 pd=0 as=0 ps=0 
M2097 op_T0_lda clock1 GND GND efet w=1410 l=658
+ ad=0 pd=0 as=0 ps=0 
M2098 op_T0_acc clock1 GND GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M2099 op_T0_tay clock1 GND GND efet w=1222 l=658
+ ad=0 pd=0 as=0 ps=0 
M2100 op_T0_shift_a clock1 GND GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M2101 op_T0_tax clock1 GND GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M2102 op_T0_bit clock1 GND GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M2103 op_T0_and clock1 GND GND efet w=1222 l=658
+ ad=0 pd=0 as=0 ps=0 
M2104 GND notir5 op_T5_rts GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2105 GND notir5 op_jsr GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2106 GND notir5 xx_op_T5_jsr GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M2107 GND notir5 x_op_T3_plp_pla GND efet w=1222 l=658
+ ad=0 pd=0 as=0 ps=0 
M2108 GND notir5 op_T__bit GND efet w=1222 l=658
+ ad=0 pd=0 as=0 ps=0 
M2109 GND notir5 x_op_T__adc_sbc GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2110 GND notir5 x_op_T0_bit GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2111 GND notir5 op_T0_plp GND efet w=1410 l=564
+ ad=0 pd=0 as=0 ps=0 
M2112 n_74 fetch n_1675 GND efet w=2162 l=752
+ ad=1.01614e+06 pd=5264 as=3.879e+06 ps=10152 
M2113 n_1309 cp1 n_74 GND efet w=2162 l=940
+ ad=1.11157e+07 pd=34404 as=0 ps=0 
M2114 n_1675 cclk notir6 GND efet w=1222 l=752
+ ad=0 pd=0 as=0 ps=0 
M2115 op_branch_done clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2116 op_T0_shift_right_a clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2117 op_T0_brk_rti clock1 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M2118 op_T0_jmp clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2119 GND notir5 op_clv GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2120 op_T0_cli_sei clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2121 op_T0_clc_sec clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2122 x_op_T0_bit clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2123 op_T0_plp clock1 GND GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M2124 ir5 ir5 Vdd GND dfet w=940 l=658
+ ad=1.75121e+08 pd=615324 as=0 ps=0 
M2125 op_T0_cld_sed clock1 GND GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2126 GND n_1609 ir5 GND efet w=11844 l=658
+ ad=0 pd=0 as=1.23174e+07 ps=28576 
M2127 GND n_1693 n_1312 GND efet w=5687 l=611
+ ad=0 pd=0 as=6.36192e+06 ps=21808 
M2128 Vdd n_1312 n_1312 GND dfet w=940 l=1504
+ ad=0 pd=0 as=1.12924e+07 ps=33276 
M2129 nNMIG nNMIG Vdd GND dfet w=940 l=752
+ ad=5.72396e+07 pd=204356 as=0 ps=0 
M2130 GND n_1312 nNMIG GND efet w=5123 l=611
+ ad=0 pd=0 as=0 ps=0 
M2131 n_1312 n_1291 GND GND efet w=5546 l=658
+ ad=0 pd=0 as=0 ps=0 
M2132 GND clock2 op_T__dex GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M2133 GND clock2 op_T__inx GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M2134 GND clock2 op_T__iny_dey GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M2135 brk_done notRdy0 GND GND efet w=8131 l=611
+ ad=1.78929e+07 pd=43240 as=0 ps=0 
M2136 n_1291 cp1 brk_done GND efet w=1222 l=752
+ ad=2.06762e+06 pd=8648 as=0 ps=0 
M2137 Vdd brk_done brk_done GND dfet w=846 l=752
+ ad=0 pd=0 as=1.1478e+08 ps=417924 
M2138 GND n_861 brk_done GND efet w=9071 l=611
+ ad=0 pd=0 as=0 ps=0 
M2139 GND n_1452 n_861 GND efet w=7144 l=658
+ ad=0 pd=0 as=9.93166e+06 ps=27824 
M2140 Vdd n_861 n_861 GND dfet w=940 l=1128
+ ad=0 pd=0 as=1.70535e+07 ps=55084 
M2141 VEC1 cclk n_1452 GND efet w=1128 l=846
+ ad=8.70346e+06 pd=27260 as=2.04995e+06 ps=8272 
M2142 n_912 VEC1 GND GND efet w=4512 l=658
+ ad=3.83482e+06 pd=12972 as=0 ps=0 
M2143 n_912 notRdy0 n_1290 GND efet w=3666 l=564
+ ad=0 pd=0 as=1.207e+07 ps=33840 
M2144 Vdd n_1290 n_1290 GND dfet w=940 l=1598
+ ad=0 pd=0 as=6.90975e+06 ps=21244 
M2145 n_1290 n_1126 GND GND efet w=4136 l=564
+ ad=0 pd=0 as=0 ps=0 
M2146 n_1717 op_T2_abs_y GND GND efet w=2820 l=658
+ ad=2.81162e+07 pd=68620 as=0 ps=0 
M2147 GND op_T0_iny_dey n_1717 GND efet w=2820 l=658
+ ad=0 pd=0 as=0 ps=0 
M2148 n_1717 x_op_T0_tya GND GND efet w=2820 l=658
+ ad=0 pd=0 as=0 ps=0 
M2149 GND op_T0_cpy_iny n_1717 GND efet w=2820 l=564
+ ad=0 pd=0 as=0 ps=0 
M2150 n_1717 op_T3_ind_y GND GND efet w=2914 l=658
+ ad=0 pd=0 as=0 ps=0 
M2151 n_1717 n_1717 Vdd GND dfet w=940 l=1410
+ ad=6.17195e+07 pd=223532 as=0 ps=0 
M2152 n_1303 n_1303 Vdd GND dfet w=940 l=1316
+ ad=2.39102e+07 pd=82720 as=0 ps=0 
M2153 n_1303 n_335 n_508 GND efet w=6909 l=611
+ ad=1.2556e+07 pd=34028 as=5.19557e+06 ps=18800 
M2154 n_508 op_from_x GND GND efet w=7708 l=564
+ ad=0 pd=0 as=0 ps=0 
M2155 n_1126 cclk VEC0 GND efet w=1128 l=752
+ ad=1.85556e+06 pd=6580 as=1.78576e+07 ps=48692 
M2156 n_1290 cp1 n_698 GND efet w=1128 l=752
+ ad=0 pd=0 as=1.50212e+06 ps=7144 
M2157 n_1397 n_335 n_1303 GND efet w=5546 l=564
+ ad=2.60662e+06 pd=12032 as=0 ps=0 
M2158 GND op_sty_cpy_mem n_1397 GND efet w=5546 l=658
+ ad=0 pd=0 as=0 ps=0 
M2159 n_1604 op_sty_cpy_mem GND GND efet w=5546 l=658
+ ad=2.60662e+06 pd=12032 as=0 ps=0 
M2160 n_1717 n_335 n_1604 GND efet w=5546 l=564
+ ad=0 pd=0 as=0 ps=0 
M2161 n_1106 op_T2_ind_x GND GND efet w=2820 l=658
+ ad=2.68438e+07 pd=65800 as=0 ps=0 
M2162 GND x_op_T0_txa n_1106 GND efet w=2820 l=564
+ ad=0 pd=0 as=0 ps=0 
M2163 n_1106 op_T0_dex GND GND efet w=2820 l=564
+ ad=0 pd=0 as=0 ps=0 
M2164 GND op_T0_cpx_inx n_1106 GND efet w=2820 l=658
+ ad=0 pd=0 as=0 ps=0 
M2165 n_1106 n_1106 Vdd GND dfet w=846 l=1316
+ ad=6.35573e+07 pd=254928 as=0 ps=0 
M2166 GND op_T0_txs n_1106 GND efet w=2820 l=564
+ ad=0 pd=0 as=0 ps=0 
M2167 Vdd n_1244 n_1244 GND dfet w=940 l=1598
+ ad=0 pd=0 as=9.90516e+06 ps=29516 
M2168 n_1351 op_T2_idx_x_xy n_1717 GND efet w=5640 l=658
+ ad=4.39149e+06 pd=13160 as=0 ps=0 
M2169 GND op_xy n_1351 GND efet w=5875 l=611
+ ad=0 pd=0 as=0 ps=0 
M2170 n_1244 op_xy GND GND efet w=3243 l=611
+ ad=3.69345e+06 pd=10716 as=0 ps=0 
M2171 GND clock2 op_T__ora_and_eor_adc GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2172 GND clock2 op_T__adc_sbc GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M2173 GND clock2 op_T__shift_a GND efet w=1363 l=611
+ ad=0 pd=0 as=0 ps=0 
M2174 n_844 op_T0_ldx_tax_tsx GND GND efet w=2726 l=564
+ ad=1.25825e+07 pd=35532 as=0 ps=0 
M2175 GND op_T__dex n_844 GND efet w=2726 l=470
+ ad=0 pd=0 as=0 ps=0 
M2176 n_844 op_T__inx GND GND efet w=2726 l=658
+ ad=0 pd=0 as=0 ps=0 
M2177 GND op_T__iny_dey n_616 GND efet w=2726 l=564
+ ad=0 pd=0 as=1.2229e+07 ps=34968 
M2178 n_616 op_T0_ldy_mem GND GND efet w=2726 l=564
+ ad=0 pd=0 as=0 ps=0 
M2179 GND op_T0_tay_ldy_not_idx n_616 GND efet w=2773 l=611
+ ad=0 pd=0 as=0 ps=0 
M2180 n_1464 op_T0_jsr GND GND efet w=2444 l=658
+ ad=1.92713e+07 pd=47376 as=0 ps=0 
M2181 GND op_T5_brk n_1464 GND efet w=2444 l=658
+ ad=0 pd=0 as=0 ps=0 
M2182 n_1464 op_T0_php_pha GND GND efet w=2444 l=658
+ ad=0 pd=0 as=0 ps=0 
M2183 GND op_T4_rts n_1464 GND efet w=2444 l=658
+ ad=0 pd=0 as=0 ps=0 
M2184 n_1464 op_T3_plp_pla GND GND efet w=2444 l=658
+ ad=0 pd=0 as=0 ps=0 
M2185 GND op_T5_rti n_1464 GND efet w=2444 l=752
+ ad=0 pd=0 as=0 ps=0 
M2186 n_844 n_844 Vdd GND dfet w=846 l=1598
+ ad=6.63142e+07 pd=261320 as=0 ps=0 
M2187 VEC0 notRdy0 GND GND efet w=3666 l=564
+ ad=0 pd=0 as=0 ps=0 
M2188 GND n_698 VEC1 GND efet w=5781 l=799
+ ad=0 pd=0 as=0 ps=0 
M2189 Vdd VEC1 VEC1 GND dfet w=1034 l=1034
+ ad=0 pd=0 as=2.51914e+07 ps=79524 
M2190 GND VEC1 nVEC GND efet w=3572 l=658
+ ad=0 pd=0 as=0 ps=0 
M2191 Vdd nVEC nVEC GND dfet w=940 l=940
+ ad=0 pd=0 as=8.06108e+07 ps=287076 
M2192 nVEC VEC0 GND GND efet w=3478 l=564
+ ad=0 pd=0 as=0 ps=0 
M2193 n_445 n_862 GND GND efet w=16262 l=564
+ ad=7.81102e+06 pd=23876 as=0 ps=0 
M2194 n_1103 n_1244 GND GND efet w=5452 l=658
+ ad=2.04995e+06 pd=11656 as=0 ps=0 
M2195 n_1106 op_T2_idx_x_xy n_1103 GND efet w=5452 l=658
+ ad=0 pd=0 as=0 ps=0 
M2196 n_734 n_335 n_1106 GND efet w=5546 l=564
+ ad=5.73456e+06 pd=13160 as=0 ps=0 
M2197 GND op_from_x n_734 GND efet w=5593 l=611
+ ad=0 pd=0 as=0 ps=0 
M2198 Vdd VEC0 VEC0 GND dfet w=940 l=1316
+ ad=0 pd=0 as=5.30602e+07 ps=196272 
M2199 Vdd n_946 n_946 GND dfet w=846 l=1222
+ ad=0 pd=0 as=1.08153e+07 ps=35344 
M2200 n_616 n_616 Vdd GND dfet w=752 l=1504
+ ad=6.91682e+07 pd=266772 as=0 ps=0 
M2201 Vdd n_1586 n_1586 GND dfet w=940 l=1504
+ ad=0 pd=0 as=6.38666e+07 ps=251168 
M2202 VEC0 n_689 GND GND efet w=3196 l=564
+ ad=0 pd=0 as=0 ps=0 
M2203 n_454 n_844 n_946 GND efet w=5640 l=658
+ ad=3.41953e+06 pd=12972 as=1.00907e+07 ps=27448 
M2204 GND n_616 n_454 GND efet w=5969 l=517
+ ad=0 pd=0 as=0 ps=0 
M2205 n_1586 op_T0_tsx GND GND efet w=2914 l=658
+ ad=5.99964e+06 pd=20304 as=0 ps=0 
M2206 n_1464 n_1464 Vdd GND dfet w=846 l=1598
+ ad=6.77721e+06 pd=19364 as=0 ps=0 
M2207 n_1109 n_1464 GND GND efet w=3290 l=658
+ ad=1.23439e+07 pd=34968 as=0 ps=0 
M2208 GND op_T5_brk n_689 GND efet w=2538 l=658
+ ad=0 pd=0 as=4.80678e+06 ps=16356 
M2209 Vdd n_1109 n_1109 GND dfet w=846 l=1222
+ ad=0 pd=0 as=3.15975e+07 ps=104904 
M2210 Vdd n_632 n_632 GND dfet w=846 l=1504
+ ad=0 pd=0 as=5.12576e+07 ps=198152 
M2211 Vdd n_1358 n_1358 GND dfet w=846 l=940
+ ad=0 pd=0 as=4.92165e+07 ps=198340 
M2212 n_689 n_689 Vdd GND dfet w=940 l=1598
+ ad=1.24499e+07 pd=40420 as=0 ps=0 
M2213 n_632 op_T2_stack GND GND efet w=3196 l=658
+ ad=9.79912e+06 pd=33088 as=0 ps=0 
M2214 Vdd n_1714 n_1714 GND dfet w=940 l=1504
+ ad=0 pd=0 as=9.86098e+06 ps=32148 
M2215 n_445 n_445 Vdd GND dfet w=1598 l=564
+ ad=8.13354e+07 pd=286700 as=0 ps=0 
M2216 n_317 n_445 GND GND efet w=4512 l=658
+ ad=4.02038e+06 pd=14100 as=0 ps=0 
M2217 n_1714 pipeUNK26 GND GND efet w=5546 l=564
+ ad=7.74034e+06 pd=18800 as=0 ps=0 
M2218 pipeUNK26 cclk n_132 GND efet w=1034 l=752
+ ad=1.15752e+06 pd=5264 as=6.24705e+06 ps=21056 
M2219 Vdd n_317 n_317 GND dfet w=940 l=940
+ ad=0 pd=0 as=1.35368e+07 ps=47564 
M2220 GND n_445 n_417 GND efet w=6909 l=705
+ ad=0 pd=0 as=1.336e+07 ps=35156 
M2221 Vdd n_317 n_417 GND dfet w=1504 l=658
+ ad=0 pd=0 as=0 ps=0 
M2222 n_417 n_445 GND GND efet w=5076 l=564
+ ad=0 pd=0 as=0 ps=0 
M2223 sync n_445 GND GND efet w=17108 l=658
+ ad=1.67866e+08 pd=229736 as=0 ps=0 
M2224 Vdd n_417 sync GND efet w=8789 l=611
+ ad=0 pd=0 as=0 ps=0 
M2225 Vdd n_417 sync GND efet w=16309 l=611
+ ad=0 pd=0 as=0 ps=0 
M2226 GND n_445 sync GND efet w=17108 l=564
+ ad=0 pd=0 as=0 ps=0 
M2227 sync n_417 Vdd GND efet w=14852 l=564
+ ad=0 pd=0 as=0 ps=0 
M2228 sync n_445 GND GND efet w=17108 l=564
+ ad=0 pd=0 as=0 ps=0 
M2229 Vdd n_417 sync GND efet w=12502 l=658
+ ad=0 pd=0 as=0 ps=0 
M2230 GND n_445 sync GND efet w=17108 l=564
+ ad=0 pd=0 as=0 ps=0 
M2231 sync n_417 Vdd GND efet w=11938 l=658
+ ad=0 pd=0 as=0 ps=0 
M2232 GND n_1447 n_1175 GND efet w=4700 l=658
+ ad=0 pd=0 as=5.50483e+06 ps=20304 
M2233 n_1175 n_1175 Vdd GND dfet w=846 l=1598
+ ad=1.21672e+07 pd=37600 as=0 ps=0 
M2234 n_1447 cp1 n_262 GND efet w=1034 l=658
+ ad=2.10297e+06 pd=8460 as=1.32452e+07 ps=35720 
M2235 Vdd n_169 n_169 GND dfet w=846 l=1692
+ ad=0 pd=0 as=3.51673e+06 ps=8272 
M2236 pipeUNK29 cclk n_169 GND efet w=1128 l=658
+ ad=1.49328e+06 pd=6768 as=7.98774e+06 ps=25756 
M2237 n_1058 n_1289 n_632 GND efet w=4794 l=658
+ ad=2.70382e+06 pd=10716 as=0 ps=0 
M2238 GND op_T0_jsr n_1058 GND efet w=4794 l=564
+ ad=0 pd=0 as=0 ps=0 
M2239 n_1358 n_1109 GND GND efet w=4935 l=611
+ ad=1.5516e+07 pd=43992 as=0 ps=0 
M2240 n_1358 op_T0_txs GND GND efet w=4230 l=564
+ ad=0 pd=0 as=0 ps=0 
M2241 GND n_917 n_1358 GND efet w=5217 l=611
+ ad=0 pd=0 as=0 ps=0 
M2242 n_267 n_267 Vdd GND dfet w=940 l=1410
+ ad=4.47102e+07 pd=173148 as=0 ps=0 
M2243 n_1175 cclk pipeUNK28 GND efet w=1034 l=752
+ ad=0 pd=0 as=1.44027e+06 ps=6768 
M2244 GND n_1175 n_267 GND efet w=4136 l=658
+ ad=0 pd=0 as=1.67884e+07 ps=43240 
M2245 n_169 n_1624 GND GND efet w=5029 l=611
+ ad=0 pd=0 as=0 ps=0 
M2246 GND n_139 n_169 GND efet w=4982 l=564
+ ad=0 pd=0 as=0 ps=0 
M2247 n_1189 pipeUNK29 GND GND efet w=9400 l=564
+ ad=6.90092e+06 pd=21056 as=0 ps=0 
M2248 n_262 n_1714 n_1189 GND efet w=7238 l=564
+ ad=0 pd=0 as=0 ps=0 
M2249 n_267 n_544 GND GND efet w=2726 l=658
+ ad=0 pd=0 as=0 ps=0 
M2250 n_917 notRdy0 GND GND efet w=2538 l=658
+ ad=6.70652e+06 pd=16544 as=0 ps=0 
M2251 GND n_383 n_917 GND efet w=2538 l=564
+ ad=0 pd=0 as=0 ps=0 
M2252 n_1624 cp1 notRdy0 GND efet w=1128 l=658
+ ad=3.2163e+06 pd=11656 as=1.94392e+07 ps=62604 
M2253 n_1598 n_1511 n_262 GND efet w=4324 l=658
+ ad=4.49752e+06 pd=14476 as=0 ps=0 
M2254 GND pipeUNK28 n_1598 GND efet w=6533 l=517
+ ad=0 pd=0 as=0 ps=0 
M2255 n_262 n_262 Vdd GND dfet w=940 l=2538
+ ad=4.69192e+06 pd=10904 as=0 ps=0 
M2256 GND n_785 n_267 GND efet w=3854 l=658
+ ad=0 pd=0 as=0 ps=0 
M2257 n_920 cp1 n_785 GND efet w=1034 l=564
+ ad=5.46948e+06 pd=17860 as=1.31656e+06 ps=5452 
M2258 GND pipeUNK29 n_1511 GND efet w=4606 l=564
+ ad=0 pd=0 as=3.73763e+06 ps=13724 
M2259 n_139 n_139 Vdd GND dfet w=940 l=1504
+ ad=1.07092e+07 pd=35908 as=0 ps=0 
M2260 n_1511 n_1511 Vdd GND dfet w=846 l=1598
+ ad=9.09224e+06 pd=27636 as=0 ps=0 
M2261 GND pipeUNK27 n_920 GND efet w=4136 l=517
+ ad=0 pd=0 as=0 ps=0 
M2262 Vdd n_917 n_917 GND dfet w=940 l=1128
+ ad=0 pd=0 as=7.21901e+06 ps=25004 
M2263 notRdy0 cp1 n_902 GND efet w=1128 l=752
+ ad=0 pd=0 as=1.31656e+06 ps=6768 
M2264 n_1109 n_902 GND GND efet w=4324 l=564
+ ad=0 pd=0 as=0 ps=0 
M2265 GND n_902 n_1109 GND efet w=3290 l=658
+ ad=0 pd=0 as=0 ps=0 
M2266 n_1289 n_1289 Vdd GND dfet w=940 l=1598
+ ad=1.57192e+07 pd=55272 as=0 ps=0 
M2267 GND n_902 n_1289 GND efet w=4935 l=611
+ ad=0 pd=0 as=6.7507e+06 ps=18988 
M2268 n_920 n_920 Vdd GND dfet w=940 l=1598
+ ad=4.05572e+06 pd=10340 as=0 ps=0 
M2269 op_SRS cclk pipeUNK27 GND efet w=1175 l=893
+ ad=6.30007e+06 pd=25380 as=1.51096e+06 ps=7332 
M2270 GND op_SRS n_139 GND efet w=3572 l=658
+ ad=0 pd=0 as=6.76838e+06 ps=18048 
M2271 Vdd n_728 n_728 GND dfet w=940 l=1504
+ ad=0 pd=0 as=1.36251e+07 ps=46812 
M2272 n_728 VEC0 GND GND efet w=2444 l=658
+ ad=5.87594e+06 pd=16356 as=0 ps=0 
M2273 sync n_445 GND GND efet w=17108 l=470
+ ad=0 pd=0 as=0 ps=0 
M2274 Vdd n_417 sync GND efet w=11938 l=564
+ ad=0 pd=0 as=0 ps=0 
M2275 sync n_417 Vdd GND efet w=11938 l=658
+ ad=0 pd=0 as=0 ps=0 
M2276 Vdd n_1712 n_1712 GND dfet w=940 l=940
+ ad=0 pd=0 as=8.31468e+06 ps=31772 
M2277 Vdd C1x5Reset C1x5Reset GND dfet w=940 l=658
+ ad=0 pd=0 as=7.56803e+07 ps=275796 
M2278 Vdd n_1087 n_1087 GND dfet w=846 l=658
+ ad=0 pd=0 as=2.66847e+06 ps=10340 
M2279 GND nVEC n_1712 GND efet w=3478 l=564
+ ad=0 pd=0 as=1.35544e+07 ps=33840 
M2280 n_1712 nNMIG GND GND efet w=3478 l=564
+ ad=0 pd=0 as=0 ps=0 
M2281 GND C1x5Reset n_1712 GND efet w=3572 l=564
+ ad=0 pd=0 as=0 ps=0 
M2282 GND n_717 C1x5Reset GND efet w=5922 l=564
+ ad=0 pd=0 as=7.71383e+06 ps=21056 
M2283 Vdd n_717 n_717 GND dfet w=846 l=1598
+ ad=0 pd=0 as=1.65852e+07 ps=59220 
M2284 Reset0 cclk pipephi2Reset0x GND efet w=1034 l=846
+ ad=0 pd=0 as=1.4226e+06 ps=6392 
M2285 n_1087 brk_done GND GND efet w=5170 l=564
+ ad=1.18491e+07 pd=26320 as=0 ps=0 
M2286 GND n_717 n_1087 GND efet w=5170 l=564
+ ad=0 pd=0 as=0 ps=0 
M2287 n_717 n_1132 GND GND efet w=4371 l=611
+ ad=6.0615e+06 pd=18988 as=0 ps=0 
M2288 GND pipephi2Reset0x n_717 GND efet w=4418 l=564
+ ad=0 pd=0 as=0 ps=0 
M2289 n_1132 cp1 n_1087 GND efet w=1034 l=658
+ ad=2.31503e+06 pd=8272 as=0 ps=0 
M2290 n_696 n_0_ADL0 GND GND efet w=3948 l=564
+ ad=1.28564e+07 pd=39292 as=0 ps=0 
M2291 n_696 n_79 n_911 GND efet w=9165 l=705
+ ad=0 pd=0 as=2.28234e+07 ps=51512 
M2292 n_728 cclk pipeVectorA0 GND efet w=1034 l=846
+ ad=0 pd=0 as=1.28122e+06 ps=6580 
M2293 n_696 n_696 Vdd GND dfet w=846 l=752
+ ad=1.50124e+07 pd=52264 as=0 ps=0 
M2294 n_70 nVEC GND GND efet w=3478 l=658
+ ad=7.46642e+06 pd=18048 as=0 ps=0 
M2295 GND n_1054 n_70 GND efet w=3478 l=658
+ ad=0 pd=0 as=0 ps=0 
M2296 n_1054 C1x5Reset GND GND efet w=3478 l=564
+ ad=6.0615e+06 pd=18236 as=0 ps=0 
M2297 n_70 n_70 Vdd GND dfet w=940 l=940
+ ad=1.01791e+07 pd=35344 as=0 ps=0 
M2298 n_1712 cclk pipeVectorA2 GND efet w=1034 l=846
+ ad=0 pd=0 as=1.23704e+06 ps=6204 
M2299 GND op_ror n_544 GND efet w=5452 l=658
+ ad=0 pd=0 as=9.04806e+06 ps=21996 
M2300 GND op_T3_stack_bit_jmp n_604 GND efet w=3243 l=611
+ ad=0 pd=0 as=2.58718e+07 ps=76892 
M2301 n_604 op_T2_stack GND GND efet w=3384 l=564
+ ad=0 pd=0 as=0 ps=0 
M2302 GND op_T0 n_638 GND efet w=3337 l=611
+ ad=0 pd=0 as=4.63006e+06 ps=13724 
M2303 n_604 op_T4_brk_jsr GND GND efet w=3525 l=611
+ ad=0 pd=0 as=0 ps=0 
M2304 GND op_T4_rti n_604 GND efet w=2820 l=564
+ ad=0 pd=0 as=0 ps=0 
M2305 n_638 n_638 Vdd GND dfet w=846 l=1504
+ ad=7.8287e+06 pd=26132 as=0 ps=0 
M2306 n_604 n_604 Vdd GND dfet w=940 l=1410
+ ad=6.77721e+07 pd=250040 as=0 ps=0 
M2307 GND op_T3_ind_x n_604 GND efet w=3337 l=517
+ ad=0 pd=0 as=0 ps=0 
M2308 n_1107 op_T3_ind_x GND GND efet w=3102 l=470
+ ad=1.60904e+07 pd=47000 as=0 ps=0 
M2309 GND op_T4_ind_y n_1107 GND efet w=3243 l=611
+ ad=0 pd=0 as=0 ps=0 
M2310 n_1107 op_T2_ind_y GND GND efet w=3149 l=611
+ ad=0 pd=0 as=0 ps=0 
M2311 GND op_T3_abs_idx n_1107 GND efet w=3149 l=611
+ ad=0 pd=0 as=0 ps=0 
M2312 n_1107 op_plp_pla GND GND efet w=3713 l=517
+ ad=0 pd=0 as=0 ps=0 
M2313 n_1649 op_jmp GND GND efet w=3196 l=564
+ ad=2.46966e+07 pd=72004 as=0 ps=0 
M2314 GND op_T2_abs n_1649 GND efet w=4371 l=611
+ ad=0 pd=0 as=0 ps=0 
M2315 n_544 n_544 Vdd GND dfet w=940 l=1222
+ ad=1.3793e+07 pd=47188 as=0 ps=0 
M2316 n_1118 op_T2_ADL_ADD GND GND efet w=5170 l=564
+ ad=2.91588e+06 pd=11468 as=0 ps=0 
M2317 n_604 n_638 n_1118 GND efet w=5170 l=564
+ ad=0 pd=0 as=0 ps=0 
M2318 Vdd n_1649 n_1649 GND dfet w=940 l=1316
+ ad=0 pd=0 as=5.13107e+07 ps=203040 
M2319 n_1555 op_inc_nop n_1107 GND efet w=4982 l=752
+ ad=2.34154e+06 pd=10904 as=0 ps=0 
M2320 GND n_440 n_1555 GND efet w=4982 l=564
+ ad=0 pd=0 as=0 ps=0 
M2321 n_300 x_op_T3_ind_y GND GND efet w=2820 l=564
+ ad=2.17277e+07 pd=65612 as=0 ps=0 
M2322 GND op_rti_rts n_300 GND efet w=3149 l=611
+ ad=0 pd=0 as=0 ps=0 
M2323 n_1000 op_T0_adc_sbc GND GND efet w=6627 l=611
+ ad=1.01261e+07 pd=32148 as=0 ps=0 
M2324 GND op_T4_ind_x n_300 GND efet w=3713 l=611
+ ad=0 pd=0 as=0 ps=0 
M2325 GND op_T2_jsr n_300 GND efet w=3760 l=564
+ ad=0 pd=0 as=0 ps=0 
M2326 n_1560 op_T0_cpx_cpy_inx_iny GND GND efet w=2444 l=564
+ ad=8.3942e+06 pd=21620 as=0 ps=0 
M2327 GND op_T0_cmp n_1560 GND efet w=2444 l=564
+ ad=0 pd=0 as=0 ps=0 
M2328 n_1560 n_1055 GND GND efet w=2679 l=611
+ ad=0 pd=0 as=0 ps=0 
M2329 Vdd n_1107 n_1107 GND dfet w=940 l=1598
+ ad=0 pd=0 as=5.37229e+06 ps=15792 
M2330 Vdd n_383 n_383 GND dfet w=940 l=1316
+ ad=0 pd=0 as=2.02433e+07 ps=65424 
M2331 n_389 n_1107 GND GND efet w=3525 l=611
+ ad=5.95546e+06 pd=17672 as=0 ps=0 
M2332 Vdd n_389 n_389 GND dfet w=940 l=1222
+ ad=0 pd=0 as=2.54654e+07 ps=89112 
M2333 n_1560 n_1560 Vdd GND dfet w=752 l=1410
+ ad=8.24399e+06 pd=28576 as=0 ps=0 
M2334 GND op_rol_ror n_1000 GND efet w=4982 l=658
+ ad=0 pd=0 as=0 ps=0 
M2335 n_980 op_T3_jmp GND GND efet w=3384 l=564
+ ad=6.26472e+06 pd=17296 as=0 ps=0 
M2336 n_300 n_300 Vdd GND dfet w=846 l=1222
+ ad=2.36716e+07 pd=96068 as=0 ps=0 
M2337 GND op_T2_jsr n_383 GND efet w=4230 l=658
+ ad=0 pd=0 as=5.2044e+06 ps=16356 
M2338 GND op_T0_ora n_1145 GND efet w=3619 l=611
+ ad=0 pd=0 as=6.37959e+06 ps=24064 
M2339 Vdd n_837 n_837 GND dfet w=940 l=1598
+ ad=0 pd=0 as=2.58806e+07 ps=91180 
M2340 n_837 op_T0_eor GND GND efet w=3807 l=611
+ ad=7.30737e+06 pd=21432 as=0 ps=0 
M2341 n_1145 n_1145 Vdd GND dfet w=940 l=1316
+ ad=1.22555e+07 pd=43616 as=0 ps=0 
M2342 GND op_rti_rts n_1649 GND efet w=4371 l=611
+ ad=0 pd=0 as=0 ps=0 
M2343 Vdd n_480 n_480 GND dfet w=940 l=940
+ ad=0 pd=0 as=1.01702e+07 ps=34404 
M2344 n_480 nNMIG n_1092 GND efet w=7473 l=611
+ ad=1.08329e+07 pd=32900 as=1.51272e+07 ps=37036 
M2345 GND nIRQP n_1092 GND efet w=6768 l=564
+ ad=0 pd=0 as=0 ps=0 
M2346 n_1092 n_118 GND GND efet w=7755 l=611
+ ad=0 pd=0 as=0 ps=0 
M2347 n_1145 notRdy0 GND GND efet w=3008 l=470
+ ad=0 pd=0 as=0 ps=0 
M2348 GND op_rti_rts n_1377 GND efet w=3619 l=611
+ ad=0 pd=0 as=3.73763e+06 ps=12408 
M2349 n_1377 n_1377 Vdd GND dfet w=846 l=1598
+ ad=9.96701e+06 pd=30080 as=0 ps=0 
M2350 n_1040 n_383 GND GND efet w=6110 l=658
+ ad=9.78145e+06 pd=26132 as=0 ps=0 
M2351 n_1649 n_389 GND GND efet w=2820 l=470
+ ad=0 pd=0 as=0 ps=0 
M2352 GND op_T4_ind_x n_1649 GND efet w=2914 l=658
+ ad=0 pd=0 as=0 ps=0 
M2353 Vdd n_385 n_385 GND dfet w=846 l=1222
+ ad=0 pd=0 as=2.70382e+06 ps=8084 
M2354 n_604 notRdy0 GND GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M2355 n_385 n_604 GND GND efet w=4841 l=611
+ ad=7.78452e+06 pd=25944 as=0 ps=0 
M2356 GND n_1377 n_385 GND efet w=4653 l=611
+ ad=0 pd=0 as=0 ps=0 
M2357 GND n_1145 op_ORS GND efet w=4183 l=611
+ ad=0 pd=0 as=4.35615e+06 ps=15604 
M2358 op_ORS op_ORS Vdd GND dfet w=752 l=846
+ ad=4.19357e+07 pd=160364 as=0 ps=0 
M2359 n_202 nnT2BR GND GND efet w=4324 l=752
+ ad=8.16446e+06 pd=24816 as=0 ps=0 
M2360 n_202 n_646 GND GND efet w=4324 l=564
+ ad=0 pd=0 as=0 ps=0 
M2361 n_629 n_480 n_202 GND efet w=4418 l=658
+ ad=1.76808e+07 pd=47188 as=0 ps=0 
M2362 Vdd n_629 n_629 GND dfet w=940 l=1504
+ ad=0 pd=0 as=1.27945e+07 ps=43428 
M2363 n_1040 n_383 GND GND efet w=2820 l=658
+ ad=0 pd=0 as=0 ps=0 
M2364 n_782 n_1303 n_1040 GND efet w=8836 l=564
+ ad=1.53835e+07 pd=37036 as=0 ps=0 
M2365 Vdd n_782 n_782 GND dfet w=846 l=658
+ ad=0 pd=0 as=4.52403e+06 ps=16732 
M2366 n_1649 notRdy0 GND GND efet w=3478 l=658
+ ad=0 pd=0 as=0 ps=0 
M2367 GND n_1109 n_1649 GND efet w=4089 l=611
+ ad=0 pd=0 as=0 ps=0 
M2368 GND brk_done n_300 GND efet w=4747 l=611
+ ad=0 pd=0 as=0 ps=0 
M2369 n_1649 brk_done GND GND efet w=2914 l=564
+ ad=0 pd=0 as=0 ps=0 
M2370 GND op_T2_jsr n_1649 GND efet w=3384 l=564
+ ad=0 pd=0 as=0 ps=0 
M2371 n_385 cclk pipeUNK30 GND efet w=1128 l=658
+ ad=0 pd=0 as=1.40492e+06 ps=6204 
M2372 Vdd n_1178 n_1178 GND dfet w=940 l=1222
+ ad=0 pd=0 as=2.92737e+07 ps=106596 
M2373 GND pipeUNK31 n_1178 GND efet w=5687 l=611
+ ad=0 pd=0 as=1.67884e+07 ps=51324 
M2374 GND pipeVectorA2 n_815 GND efet w=4841 l=705
+ ad=0 pd=0 as=6.3089e+06 ps=19176 
M2375 n_1054 n_1054 Vdd GND dfet w=940 l=846
+ ad=6.16753e+06 pd=21244 as=0 ps=0 
M2376 Vdd n_0_ADL0 n_0_ADL0 GND dfet w=940 l=1598
+ ad=0 pd=0 as=3.82157e+07 ps=132540 
M2377 GND pipeVectorA0 n_0_ADL0 GND efet w=9870 l=658
+ ad=0 pd=0 as=1.14691e+07 ps=32336 
M2378 n_1117 cclk pipeVectorA1 GND efet w=1034 l=658
+ ad=7.07764e+06 pd=22748 as=1.31656e+06 ps=6768 
M2379 n_815 n_815 Vdd GND dfet w=846 l=1504
+ ad=9.82563e+06 pd=26320 as=0 ps=0 
M2380 n_1117 n_1117 Vdd GND dfet w=940 l=846
+ ad=3.44604e+06 pd=11656 as=0 ps=0 
M2381 n_1117 n_70 GND GND efet w=4230 l=564
+ ad=0 pd=0 as=0 ps=0 
M2382 GND pipeVectorA1 n_0_ADL1 GND efet w=8836 l=658
+ ad=0 pd=0 as=9.13642e+06 ps=29704 
M2383 Vdd n_0_ADL1 n_0_ADL1 GND dfet w=846 l=1504
+ ad=0 pd=0 as=3.09348e+07 ps=116748 
M2384 Vdd n_0_ADL2 n_0_ADL2 GND dfet w=846 l=1410
+ ad=0 pd=0 as=4.12641e+07 ps=163184 
M2385 GND n_815 n_0_ADL2 GND efet w=4841 l=611
+ ad=0 pd=0 as=5.87594e+06 ps=15792 
M2386 n_696 cclk n_610 GND efet w=1175 l=987
+ ad=0 pd=0 as=1.94392e+06 ps=7520 
M2387 n_1101 cclk n_190 GND efet w=1128 l=752
+ ad=1.04442e+07 pd=31396 as=1.57281e+06 ps=5828 
M2388 n_1717 cclk n_1113 GND efet w=1128 l=846
+ ad=0 pd=0 as=1.08683e+06 ps=5452 
M2389 Vdd n_582 n_582 GND dfet w=846 l=940
+ ad=0 pd=0 as=1.16724e+07 ps=37600 
M2390 GND n_610 n_582 GND efet w=6721 l=611
+ ad=0 pd=0 as=7.54594e+06 ps=18800 
M2391 GND cp1 n_43 GND efet w=19364 l=658
+ ad=0 pd=0 as=2.23904e+07 ps=52264 
M2392 n_43 n_839 Vdd GND dfet w=3948 l=658
+ ad=0 pd=0 as=0 ps=0 
M2393 GND cp1 n_43 GND efet w=11891 l=611
+ ad=0 pd=0 as=0 ps=0 
M2394 Vdd n_220 n_220 GND dfet w=846 l=940
+ ad=0 pd=0 as=1.14691e+07 ps=36660 
M2395 GND n_190 n_220 GND efet w=6627 l=611
+ ad=0 pd=0 as=7.27203e+06 ps=18612 
M2396 n_161 n_1113 GND GND efet w=5405 l=611
+ ad=7.18367e+06 pd=20116 as=0 ps=0 
M2397 Vdd n_161 n_161 GND dfet w=940 l=1128
+ ad=0 pd=0 as=9.12759e+06 ps=30832 
M2398 n_1106 cclk n_1404 GND efet w=1128 l=940
+ ad=0 pd=0 as=1.1045e+06 ps=6204 
M2399 n_133 n_133 Vdd GND dfet w=752 l=1034
+ ad=9.69309e+06 pd=30456 as=0 ps=0 
M2400 GND n_1404 n_133 GND efet w=5687 l=517
+ ad=0 pd=0 as=7.2897e+06 ps=21620 
M2401 GND cp1 n_1247 GND efet w=9776 l=564
+ ad=0 pd=0 as=2.44227e+07 ps=63168 
M2402 testpad_5 n_1127 testpad_5 GND efet w=7896 l=6862
+ ad=4.73168e+07 pd=60348 as=0 ps=0 
M2403 testpad_1 n_1127 testpad_1 GND efet w=5969 l=6439
+ ad=2.49617e+07 pd=30832 as=0 ps=0 
M2404 testpad_2 testpad_4 testpad_5 GND efet w=940 l=564
+ ad=7.40015e+07 pd=48504 as=0 ps=0 
M2405 n_1247 cp1 GND GND efet w=19646 l=658
+ ad=0 pd=0 as=0 ps=0 
M2406 GND cp1 n_1247 GND efet w=16967 l=611
+ ad=0 pd=0 as=0 ps=0 
M2407 n_1247 n_38 Vdd GND dfet w=6016 l=658
+ ad=0 pd=0 as=0 ps=0 
M2408 n_839 n_839 Vdd GND dfet w=1222 l=658
+ ad=8.28817e+06 pd=26508 as=0 ps=0 
M2409 GND cp1 n_839 GND efet w=5922 l=658
+ ad=0 pd=0 as=5.31927e+06 ps=16168 
M2410 n_1067 n_582 GND GND efet w=2350 l=658
+ ad=2.84519e+06 pd=9588 as=0 ps=0 
M2411 n_130 n_220 GND GND efet w=2444 l=658
+ ad=3.06609e+06 pd=9776 as=0 ps=0 
M2412 GND cclk n_161 GND efet w=2350 l=564
+ ad=0 pd=0 as=0 ps=0 
M2413 n_133 cclk GND GND efet w=2350 l=564
+ ad=0 pd=0 as=0 ps=0 
M2414 n_969 n_161 GND GND efet w=2350 l=564
+ ad=3.03075e+06 pd=8460 as=0 ps=0 
M2415 n_1067 n_1067 Vdd GND dfet w=940 l=1222
+ ad=1.32098e+07 pd=44556 as=0 ps=0 
M2416 Vdd n_582 ADH_ABH GND dfet w=1128 l=752
+ ad=0 pd=0 as=1.53305e+07 ps=35532 
M2417 n_130 n_130 Vdd GND dfet w=1034 l=1316
+ ad=1.08948e+07 pd=33840 as=0 ps=0 
M2418 n_38 cp1 GND GND efet w=5170 l=564
+ ad=4.79795e+06 pd=15792 as=0 ps=0 
M2419 Vdd n_38 n_38 GND dfet w=1316 l=658
+ ad=0 pd=0 as=1.00642e+07 ps=34404 
M2420 GND n_1067 ADH_ABH GND efet w=14006 l=564
+ ad=0 pd=0 as=0 ps=0 
M2421 Vdd n_220 ADL_ABL GND dfet w=846 l=752
+ ad=0 pd=0 as=1.13278e+07 ps=28764 
M2422 Vdd n_969 n_969 GND dfet w=940 l=1128
+ ad=0 pd=0 as=1.04883e+07 ps=33652 
M2423 testpad_5 diff_22278_155664# n_1701 GND efet w=1034 l=3948
+ ad=0 pd=0 as=1.28299e+07 ps=22748 
M2424 testpad_6 diff_22278_155664# n_1701 GND efet w=940 l=564
+ ad=7.49293e+06 pd=12032 as=0 ps=0 
M2425 testpad_2 testpad_4 testpad_6 GND efet w=3572 l=564
+ ad=0 pd=0 as=0 ps=0 
M2426 GND n_130 ADL_ABL GND efet w=9165 l=611
+ ad=0 pd=0 as=0 ps=0 
M2427 Vdd n_161 dpc0_YSB GND dfet w=1034 l=752
+ ad=0 pd=0 as=1.45087e+07 ps=30268 
M2428 GND n_133 n_602 GND efet w=2350 l=658
+ ad=0 pd=0 as=3.28699e+06 ps=10152 
M2429 n_602 n_602 Vdd GND dfet w=940 l=1034
+ ad=1.00112e+07 pd=36284 as=0 ps=0 
M2430 Vdd n_133 dpc2_XSB GND dfet w=940 l=752
+ ad=0 pd=0 as=1.5516e+07 ps=34028 
M2431 dpc0_YSB n_1247 GND GND efet w=6956 l=564
+ ad=0 pd=0 as=0 ps=0 
M2432 GND n_969 dpc0_YSB GND efet w=7238 l=564
+ ad=0 pd=0 as=0 ps=0 
M2433 dpc2_XSB n_602 GND GND efet w=8648 l=564
+ ad=0 pd=0 as=0 ps=0 
M2434 GND n_1247 dpc2_XSB GND efet w=8601 l=517
+ ad=0 pd=0 as=0 ps=0 
M2435 ab0 n_1100 GND GND efet w=41642 l=658
+ ad=1.28679e+08 pd=210372 as=0 ps=0 
M2436 ab0 n_1100 GND GND efet w=33135 l=611
+ ad=0 pd=0 as=0 ps=0 
M2437 ab0 n_1100 GND GND efet w=15980 l=658
+ ad=0 pd=0 as=0 ps=0 
M2438 Vdd n_855 ab0 GND efet w=6392 l=658
+ ad=0 pd=0 as=0 ps=0 
M2439 Vdd n_855 ab0 GND efet w=22513 l=611
+ ad=0 pd=0 as=0 ps=0 
M2440 GND n_1660 n_855 GND efet w=11844 l=658
+ ad=0 pd=0 as=1.38195e+07 ps=35532 
M2441 Vdd n_855 ab0 GND efet w=22419 l=611
+ ad=0 pd=0 as=0 ps=0 
M2442 Vdd n_855 ab0 GND efet w=22560 l=658
+ ad=0 pd=0 as=0 ps=0 
M2443 n_1660 abl0 GND GND efet w=3384 l=752
+ ad=4.11758e+06 pd=13160 as=0 ps=0 
M2444 n_1660 n_1660 Vdd GND dfet w=940 l=940
+ ad=1.58341e+07 pd=50008 as=0 ps=0 
M2445 GND abl0 n_1100 GND efet w=14476 l=658
+ ad=0 pd=0 as=1.32805e+07 ps=37600 
M2446 n_855 abl0 Vdd GND dfet w=1692 l=658
+ ad=0 pd=0 as=0 ps=0 
M2447 n_1100 n_1660 Vdd GND dfet w=1974 l=658
+ ad=0 pd=0 as=0 ps=0 
M2448 n_629 n_50 GND GND efet w=3760 l=658
+ ad=0 pd=0 as=0 ps=0 
M2449 n_50 cp1 INTG GND efet w=1128 l=846
+ ad=1.24588e+06 pd=5640 as=1.22202e+07 ps=34968 
M2450 Vdd n_152 n_152 GND dfet w=846 l=1128
+ ad=0 pd=0 as=1.39344e+07 ps=49820 
M2451 n_152 n_1002 GND GND efet w=2726 l=564
+ ad=1.0992e+07 pd=26696 as=0 ps=0 
M2452 n_1178 pipeUNK30 GND GND efet w=5123 l=611
+ ad=0 pd=0 as=0 ps=0 
M2453 n_389 cclk pipeUNK31 GND efet w=1034 l=658
+ ad=0 pd=0 as=1.63466e+06 ps=7144 
M2454 n_1178 pipeUNK32 GND GND efet w=5123 l=611
+ ad=0 pd=0 as=0 ps=0 
M2455 GND pipeUNK33 n_1178 GND efet w=4700 l=564
+ ad=0 pd=0 as=0 ps=0 
M2456 n_1081 cclk pipeUNK32 GND efet w=1128 l=658
+ ad=8.9332e+06 pd=27448 as=2.46524e+06 ps=6392 
M2457 n_473 cclk pipeUNK33 GND efet w=1222 l=658
+ ad=9.18944e+06 pd=24252 as=1.82022e+06 ps=7896 
M2458 Vdd n_1081 n_1081 GND dfet w=846 l=1222
+ ad=0 pd=0 as=2.54919e+07 ps=99640 
M2459 n_1081 n_1560 GND GND efet w=3619 l=611
+ ad=0 pd=0 as=0 ps=0 
M2460 n_300 n_389 GND GND efet w=2914 l=658
+ ad=0 pd=0 as=0 ps=0 
M2461 Vdd n_1130 n_1130 GND dfet w=940 l=1222
+ ad=0 pd=0 as=4.91282e+07 ps=184616 
M2462 n_1130 n_1109 GND GND efet w=2820 l=658
+ ad=1.99252e+07 pd=59784 as=0 ps=0 
M2463 GND n_1258 n_1130 GND efet w=3948 l=564
+ ad=0 pd=0 as=0 ps=0 
M2464 n_1130 n_862 GND GND efet w=2726 l=564
+ ad=0 pd=0 as=0 ps=0 
M2465 GND n_192 n_1130 GND efet w=2632 l=658
+ ad=0 pd=0 as=0 ps=0 
M2466 n_847 n_300 GND GND efet w=3478 l=564
+ ad=6.33541e+06 pd=18988 as=0 ps=0 
M2467 GND op_T2 n_152 GND efet w=3901 l=611
+ ad=0 pd=0 as=0 ps=0 
M2468 n_256 op_T5_rti GND GND efet w=2914 l=564
+ ad=2.02786e+07 pd=63920 as=0 ps=0 
M2469 n_152 n_952 GND GND efet w=2632 l=658
+ ad=0 pd=0 as=0 ps=0 
M2470 GND n_630 n_152 GND efet w=4230 l=564
+ ad=0 pd=0 as=0 ps=0 
M2471 Vdd op_EORS op_EORS GND dfet w=940 l=1598
+ ad=0 pd=0 as=2.59425e+07 ps=86292 
M2472 op_EORS n_837 GND GND efet w=3525 l=611
+ ad=6.68002e+06 pd=18988 as=0 ps=0 
M2473 n_372 notRdy0 GND GND efet w=2726 l=658
+ ad=3.05726e+06 pd=9212 as=0 ps=0 
M2474 n_372 n_372 Vdd GND dfet w=940 l=1128
+ ad=8.72997e+06 pd=29328 as=0 ps=0 
M2475 n_847 n_847 Vdd GND dfet w=846 l=1034
+ ad=6.83906e+06 pd=22372 as=0 ps=0 
M2476 n_1408 n_1044 n_1000 GND efet w=5264 l=564
+ ad=4.17059e+06 pd=13536 as=0 ps=0 
M2477 n_980 n_980 Vdd GND dfet w=846 l=1504
+ ad=1.90593e+07 pd=65424 as=0 ps=0 
M2478 Vdd n_1408 n_1408 GND dfet w=846 l=1598
+ ad=0 pd=0 as=1.57899e+07 ps=55836 
M2479 n_104 n_847 GND GND efet w=3290 l=658
+ ad=2.78069e+07 pd=73132 as=0 ps=0 
M2480 n_1130 n_1002 GND GND efet w=3102 l=564
+ ad=0 pd=0 as=0 ps=0 
M2481 n_1365 n_862 GND GND efet w=3760 l=470
+ ad=2.12064e+06 pd=8648 as=0 ps=0 
M2482 n_1085 notRdy0 n_1365 GND efet w=3760 l=658
+ ad=1.2017e+07 pd=34216 as=0 ps=0 
M2483 n_911 n_877 GND GND efet w=2068 l=658
+ ad=0 pd=0 as=0 ps=0 
M2484 GND n_1343 n_911 GND efet w=9165 l=611
+ ad=0 pd=0 as=0 ps=0 
M2485 n_911 n_877 GND GND efet w=5734 l=564
+ ad=0 pd=0 as=0 ps=0 
M2486 n_1172 n_372 n_1085 GND efet w=5170 l=564
+ ad=1.10362e+07 pd=23312 as=0 ps=0 
M2487 n_405 BRtaken n_1172 GND efet w=5170 l=658
+ ad=4.8598e+06 pd=12220 as=0 ps=0 
M2488 GND nnT2BR n_405 GND efet w=5170 l=658
+ ad=0 pd=0 as=0 ps=0 
M2489 n_1343 n_152 GND GND efet w=2820 l=658
+ ad=5.98197e+06 pd=18424 as=0 ps=0 
M2490 GND notRdy0 n_1343 GND efet w=2820 l=564
+ ad=0 pd=0 as=0 ps=0 
M2491 Vdd n_1085 n_1085 GND dfet w=846 l=1598
+ ad=0 pd=0 as=7.50176e+06 ps=24440 
M2492 n_79 n_236 GND GND efet w=8554 l=564
+ ad=1.02498e+07 pd=28576 as=0 ps=0 
M2493 GND n_646 n_1172 GND efet w=3384 l=658
+ ad=0 pd=0 as=0 ps=0 
M2494 n_1343 n_1343 Vdd GND dfet w=752 l=1128
+ ad=8.7388e+06 pd=27260 as=0 ps=0 
M2495 n_629 cclk n_760 GND efet w=1034 l=846
+ ad=0 pd=0 as=3.27816e+06 ps=10528 
M2496 D1x1 D1x1 Vdd GND dfet w=846 l=752
+ ad=7.55301e+07 pd=290272 as=0 ps=0 
M2497 Vdd n_1594 n_1594 GND dfet w=846 l=1222
+ ad=0 pd=0 as=9.09224e+06 ps=34404 
M2498 GND n_1358 n_396 GND efet w=2726 l=658
+ ad=0 pd=0 as=4.80678e+06 ps=17672 
M2499 INTG brk_done GND GND efet w=2350 l=470
+ ad=0 pd=0 as=0 ps=0 
M2500 GND n_760 INTG GND efet w=4136 l=564
+ ad=0 pd=0 as=0 ps=0 
M2501 D1x1 C1x5Reset GND GND efet w=5875 l=517
+ ad=1.35102e+07 pd=33088 as=0 ps=0 
M2502 GND INTG D1x1 GND efet w=6016 l=658
+ ad=0 pd=0 as=0 ps=0 
M2503 n_79 n_79 Vdd GND dfet w=940 l=846
+ ad=1.28475e+07 pd=41548 as=0 ps=0 
M2504 n_656 n_779 n_1594 GND efet w=5076 l=658
+ ad=2.38572e+06 pd=11092 as=6.71536e+06 ps=24064 
M2505 GND n_604 n_656 GND efet w=5076 l=658
+ ad=0 pd=0 as=0 ps=0 
M2506 n_795 n_1649 GND GND efet w=2726 l=658
+ ad=4.67424e+06 pd=18424 as=0 ps=0 
M2507 Vdd n_795 n_795 GND dfet w=846 l=1128
+ ad=0 pd=0 as=6.24705e+06 ps=22372 
M2508 n_396 n_396 Vdd GND dfet w=940 l=1034
+ ad=4.28546e+06 pd=13348 as=0 ps=0 
M2509 n_616 cclk n_460 GND efet w=1128 l=846
+ ad=0 pd=0 as=1.23704e+06 ps=7144 
M2510 n_844 cclk n_459 GND efet w=1222 l=846
+ ad=0 pd=0 as=1.30773e+06 ps=7332 
M2511 n_1586 cclk n_621 GND efet w=1034 l=846
+ ad=0 pd=0 as=1.40492e+06 ps=7144 
M2512 n_632 cclk n_339 GND efet w=1128 l=940
+ ad=0 pd=0 as=1.36958e+06 ps=5452 
M2513 n_1358 cclk n_521 GND efet w=1222 l=940
+ ad=0 pd=0 as=1.30773e+06 ps=6580 
M2514 INTG INTG Vdd GND dfet w=940 l=1504
+ ad=2.02168e+07 pd=74636 as=0 ps=0 
M2515 n_1304 op_T0_sbc GND GND efet w=4465 l=611
+ ad=7.03346e+06 pd=17296 as=0 ps=0 
M2516 GND n_673 n_1304 GND efet w=3666 l=658
+ ad=0 pd=0 as=0 ps=0 
M2517 n_1304 n_1304 Vdd GND dfet w=987 l=1269
+ ad=1.27945e+07 pd=44744 as=0 ps=0 
M2518 n_605 n_1081 GND GND efet w=7661 l=611
+ ad=1.5622e+07 pd=49068 as=0 ps=0 
M2519 GND op_T0_sbc n_605 GND efet w=7614 l=564
+ ad=0 pd=0 as=0 ps=0 
M2520 GND clock2 op_T__bit GND efet w=1222 l=658
+ ad=0 pd=0 as=0 ps=0 
M2521 GND clock2 x_op_T__adc_sbc GND efet w=1410 l=752
+ ad=0 pd=0 as=0 ps=0 
M2522 GND clock2 op_T__cmp GND efet w=1269 l=705
+ ad=0 pd=0 as=0 ps=0 
M2523 GND clock2 op_T__cpx_cpy_abs GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M2524 GND clock2 op_T__asl_rol_a GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M2525 notir5 notir5 Vdd GND dfet w=940 l=564
+ ad=1.94913e+08 pd=674356 as=0 ps=0 
M2526 GND ir5 notir5 GND efet w=8742 l=658
+ ad=0 pd=0 as=1.85291e+07 ps=43616 
M2527 GND clock2 op_T__cpx_cpy_imm_zp GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M2528 n_1378 fetch n_1609 GND efet w=2162 l=752
+ ad=1.01614e+06 pd=5264 as=3.84366e+06 ps=10152 
M2529 n_928 cp1 n_1378 GND efet w=2162 l=940
+ ad=1.41641e+07 pd=36660 as=0 ps=0 
M2530 n_1609 cclk notir5 GND efet w=1128 l=752
+ ad=0 pd=0 as=0 ps=0 
M2531 n_1455 op_T0_tya GND GND efet w=3478 l=658
+ ad=2.24081e+07 pd=58844 as=0 ps=0 
M2532 n_1455 n_1455 Vdd GND dfet w=846 l=1598
+ ad=6.74275e+07 pd=248536 as=0 ps=0 
M2533 n_1455 op_T__shift_a GND GND efet w=3572 l=658
+ ad=0 pd=0 as=0 ps=0 
M2534 GND op_T0_txa n_1455 GND efet w=2820 l=658
+ ad=0 pd=0 as=0 ps=0 
M2535 n_1455 op_T0_pla GND GND efet w=2726 l=658
+ ad=0 pd=0 as=0 ps=0 
M2536 GND op_T0_lda n_1455 GND efet w=2726 l=658
+ ad=0 pd=0 as=0 ps=0 
M2537 n_1563 op_T0_acc GND GND efet w=4794 l=658
+ ad=2.23551e+06 pd=10528 as=0 ps=0 
M2538 n_11 n_397 n_1563 GND efet w=4794 l=658
+ ad=1.8264e+07 pd=59032 as=0 ps=0 
M2539 GND op_T0_tay n_11 GND efet w=3290 l=564
+ ad=0 pd=0 as=0 ps=0 
M2540 n_11 op_T0_shift_a GND GND efet w=3807 l=517
+ ad=0 pd=0 as=0 ps=0 
M2541 GND op_T__adc_sbc n_1455 GND efet w=3290 l=658
+ ad=0 pd=0 as=0 ps=0 
M2542 GND op_T__ora_and_eor_adc n_1455 GND efet w=2914 l=658
+ ad=0 pd=0 as=0 ps=0 
M2543 GND op_T0_lda n_397 GND efet w=3149 l=611
+ ad=0 pd=0 as=5.66388e+06 ps=16544 
M2544 GND op_T0_tax n_11 GND efet w=3948 l=658
+ ad=0 pd=0 as=0 ps=0 
M2545 n_669 op_T0_bit GND GND efet w=3948 l=658
+ ad=4.6389e+06 pd=16544 as=0 ps=0 
M2546 Vdd n_397 n_397 GND dfet w=846 l=1222
+ ad=0 pd=0 as=7.1925e+06 ps=21056 
M2547 Vdd n_1090 n_1090 GND dfet w=846 l=1128
+ ad=0 pd=0 as=4.95169e+07 ps=195708 
M2548 n_1681 n_440 n_905 GND efet w=4888 l=658
+ ad=2.41223e+06 pd=10716 as=4.94816e+06 ps=15416 
M2549 GND op_shift n_1681 GND efet w=4888 l=658
+ ad=0 pd=0 as=0 ps=0 
M2550 Vdd n_384 n_384 GND dfet w=846 l=1222
+ ad=0 pd=0 as=1.00289e+07 ps=32148 
M2551 Vdd n_1412 n_1412 GND dfet w=846 l=1128
+ ad=0 pd=0 as=5.59319e+06 ps=18612 
M2552 GND n_1222 n_1090 GND efet w=3478 l=658
+ ad=0 pd=0 as=1.24676e+07 ps=37600 
M2553 n_1090 op_T2_stack_access GND GND efet w=3666 l=658
+ ad=0 pd=0 as=0 ps=0 
M2554 n_1222 n_1225 GND GND efet w=4042 l=658
+ ad=6.42377e+06 pd=21432 as=0 ps=0 
M2555 n_905 n_905 Vdd GND dfet w=940 l=1504
+ ad=5.76107e+06 pd=16920 as=0 ps=0 
M2556 GND op_T0_and n_669 GND efet w=2820 l=658
+ ad=0 pd=0 as=0 ps=0 
M2557 n_595 op_T4_abs_idx GND GND efet w=4982 l=658
+ ad=6.71536e+06 pd=18236 as=0 ps=0 
M2558 GND op_T5_ind_y n_595 GND efet w=3525 l=611
+ ad=0 pd=0 as=0 ps=0 
M2559 nop_branch_done op_branch_done GND GND efet w=3478 l=658
+ ad=4.46218e+06 pd=15416 as=0 ps=0 
M2560 n_11 n_11 Vdd GND dfet w=893 l=1551
+ ad=6.1746e+07 pd=224848 as=0 ps=0 
M2561 n_669 n_669 Vdd GND dfet w=846 l=1504
+ ad=8.02309e+06 pd=24628 as=0 ps=0 
M2562 n_595 n_595 Vdd GND dfet w=846 l=1222
+ ad=1.25736e+07 pd=42676 as=0 ps=0 
M2563 GND n_1412 n_384 GND efet w=3243 l=611
+ ad=0 pd=0 as=2.24611e+07 ps=55460 
M2564 Vdd op_ANDS op_ANDS GND dfet w=940 l=1504
+ ad=0 pd=0 as=6.10833e+07 ps=224848 
M2565 nop_branch_done nop_branch_done Vdd GND dfet w=940 l=1504
+ ad=7.70499e+06 pd=22560 as=0 ps=0 
M2566 n_366 op_T0_shift_right_a GND GND efet w=4653 l=611
+ ad=8.34118e+06 pd=24816 as=0 ps=0 
M2567 n_1012 n_440 n_366 GND efet w=5264 l=564
+ ad=3.19863e+06 pd=12972 as=0 ps=0 
M2568 GND op_shift_right n_1012 GND efet w=5593 l=611
+ ad=0 pd=0 as=0 ps=0 
M2569 n_824 op_T2_brk GND GND efet w=3384 l=564
+ ad=1.13631e+07 pd=33652 as=0 ps=0 
M2570 GND op_T3_jsr n_824 GND efet w=3760 l=658
+ ad=0 pd=0 as=0 ps=0 
M2571 GND op_ANDS n_11 GND efet w=3666 l=564
+ ad=0 pd=0 as=0 ps=0 
M2572 Vdd n_1037 n_1037 GND dfet w=846 l=1504
+ ad=0 pd=0 as=6.03587e+07 ps=211688 
M2573 Vdd n_366 n_366 GND dfet w=940 l=1034
+ ad=0 pd=0 as=5.97314e+06 ps=20492 
M2574 n_1222 n_1222 Vdd GND dfet w=940 l=1128
+ ad=7.02462e+06 pd=21432 as=0 ps=0 
M2575 GND n_946 n_384 GND efet w=2632 l=658
+ ad=0 pd=0 as=0 ps=0 
M2576 GND n_1455 n_1412 GND efet w=4089 l=611
+ ad=0 pd=0 as=5.1779e+06 ps=14288 
M2577 n_1347 op_T0_shift_a GND GND efet w=4371 l=705
+ ad=2.61457e+07 pd=75012 as=0 ps=0 
M2578 GND n_905 n_979 GND efet w=2538 l=564
+ ad=0 pd=0 as=3.99387e+06 ps=12596 
M2579 n_979 n_979 Vdd GND dfet w=846 l=1598
+ ad=6.22054e+06 pd=18988 as=0 ps=0 
M2580 Vdd n_473 n_473 GND dfet w=846 l=1222
+ ad=0 pd=0 as=1.56927e+07 ps=62228 
M2581 n_1004 n_1408 GND GND efet w=6721 l=611
+ ad=3.4372e+06 pd=14476 as=0 ps=0 
M2582 n_473 n_980 n_1004 GND efet w=6721 l=611
+ ad=0 pd=0 as=0 ps=0 
M2583 n_1347 n_979 GND GND efet w=2726 l=658
+ ad=0 pd=0 as=0 ps=0 
M2584 GND op_T5_jsr n_1219 GND efet w=2444 l=564
+ ad=0 pd=0 as=3.5344e+06 ps=9964 
M2585 n_1347 n_782 GND GND efet w=2632 l=658
+ ad=0 pd=0 as=0 ps=0 
M2586 GND n_1219 n_1002 GND efet w=4277 l=611
+ ad=0 pd=0 as=5.69922e+06 ps=15792 
M2587 n_1219 n_1219 Vdd GND dfet w=940 l=1598
+ ad=7.3869e+06 pd=22184 as=0 ps=0 
M2588 n_1347 n_862 GND GND efet w=3384 l=658
+ ad=0 pd=0 as=0 ps=0 
M2589 n_384 n_1258 GND GND efet w=3666 l=658
+ ad=0 pd=0 as=0 ps=0 
M2590 GND n_550 n_1347 GND efet w=3337 l=611
+ ad=0 pd=0 as=0 ps=0 
M2591 n_384 op_ANDS GND GND efet w=1598 l=564
+ ad=0 pd=0 as=0 ps=0 
M2592 GND op_ANDS n_550 GND efet w=3619 l=611
+ ad=0 pd=0 as=8.87134e+06 ps=23688 
M2593 n_384 op_ANDS GND GND efet w=1880 l=658
+ ad=0 pd=0 as=0 ps=0 
M2594 n_1347 n_1347 Vdd GND dfet w=752 l=1222
+ ad=4.86864e+07 pd=180480 as=0 ps=0 
M2595 Vdd n_506 n_506 GND dfet w=752 l=1034
+ ad=0 pd=0 as=5.26979e+07 ps=190632 
M2596 GND n_669 op_ANDS GND efet w=4794 l=658
+ ad=0 pd=0 as=6.088e+06 ps=19552 
M2597 GND n_192 n_506 GND efet w=3619 l=611
+ ad=0 pd=0 as=1.00995e+07 ps=33088 
M2598 GND n_1258 n_813 GND efet w=3384 l=658
+ ad=0 pd=0 as=7.26319e+06 ps=21808 
M2599 n_1002 n_1002 Vdd GND dfet w=846 l=940
+ ad=3.05284e+07 pd=110544 as=0 ps=0 
M2600 Vdd n_673 n_673 GND dfet w=940 l=1222
+ ad=0 pd=0 as=1.00907e+07 ps=31584 
M2601 n_1053 op_T0_adc_sbc n_673 GND efet w=6251 l=611
+ ad=4.18826e+06 pd=15980 as=4.7626e+06 ps=15980 
M2602 GND n_1002 n_605 GND efet w=3431 l=611
+ ad=0 pd=0 as=0 ps=0 
M2603 n_605 n_1002 GND GND efet w=2914 l=564
+ ad=0 pd=0 as=0 ps=0 
M2604 n_779 n_1440 n_605 GND efet w=5828 l=564
+ ad=7.66081e+06 pd=23500 as=0 ps=0 
M2605 GND Pout3 n_1053 GND efet w=5546 l=564
+ ad=0 pd=0 as=0 ps=0 
M2606 Vdd n_25 n_25 GND dfet w=846 l=1128
+ ad=0 pd=0 as=3.60862e+07 ps=128028 
M2607 n_25 n_192 GND GND efet w=4183 l=611
+ ad=7.93473e+06 pd=21056 as=0 ps=0 
M2608 Vdd n_1440 n_1440 GND dfet w=846 l=1128
+ ad=0 pd=0 as=9.43685e+06 ps=31772 
M2609 n_779 n_779 Vdd GND dfet w=752 l=1410
+ ad=3.78181e+07 pd=131224 as=0 ps=0 
M2610 GND n_384 n_550 GND efet w=3008 l=658
+ ad=0 pd=0 as=0 ps=0 
M2611 n_885 n_384 GND GND efet w=4324 l=658
+ ad=4.90398e+06 pd=18424 as=0 ps=0 
M2612 n_813 n_440 GND GND efet w=3290 l=658
+ ad=0 pd=0 as=0 ps=0 
M2613 GND n_595 n_992 GND efet w=3102 l=564
+ ad=0 pd=0 as=4.85096e+06 ps=14664 
M2614 n_239 n_595 GND GND efet w=4606 l=658
+ ad=2.16482e+06 pd=10152 as=0 ps=0 
M2615 n_192 nop_branch_done n_239 GND efet w=4606 l=658
+ ad=6.85674e+06 pd=19364 as=0 ps=0 
M2616 GND n_992 n_46 GND efet w=4277 l=611
+ ad=0 pd=0 as=8.25282e+06 ps=23500 
M2617 n_813 n_813 Vdd GND dfet w=940 l=1692
+ ad=1.15398e+07 pd=31960 as=0 ps=0 
M2618 n_992 n_992 Vdd GND dfet w=940 l=1222
+ ad=7.15716e+06 pd=22560 as=0 ps=0 
M2619 Vdd n_1101 n_1101 GND dfet w=846 l=1034
+ ad=0 pd=0 as=5.18938e+07 ps=181984 
M2620 n_192 n_192 Vdd GND dfet w=846 l=1222
+ ad=4.26956e+07 pd=155100 as=0 ps=0 
M2621 Vdd n_46 n_46 GND dfet w=893 l=1645
+ ad=0 pd=0 as=1.06032e+07 ps=34968 
M2622 GND notRdy0 n_46 GND efet w=4794 l=658
+ ad=0 pd=0 as=0 ps=0 
M2623 n_550 n_550 Vdd GND dfet w=752 l=1222
+ ad=8.78298e+06 pd=29328 as=0 ps=0 
M2624 n_885 n_885 Vdd GND dfet w=846 l=1034
+ ad=4.04335e+07 pd=143632 as=0 ps=0 
M2625 n_1508 n_813 n_1101 GND efet w=8084 l=658
+ ad=7.25436e+06 pd=21432 as=0 ps=0 
M2626 GND n_334 n_118 GND efet w=4042 l=658
+ ad=0 pd=0 as=5.50483e+06 ps=15980 
M2627 n_1688 n_1304 GND GND efet w=2914 l=658
+ ad=7.66081e+06 pd=22748 as=0 ps=0 
M2628 n_118 n_118 Vdd GND dfet w=940 l=940
+ ad=9.79912e+06 pd=33276 as=0 ps=0 
M2629 n_1688 n_1688 Vdd GND dfet w=846 l=1128
+ ad=2.45022e+07 pd=86480 as=0 ps=0 
M2630 n_1440 notRdy0 GND GND efet w=3431 l=611
+ ad=2.45641e+06 pd=7896 as=0 ps=0 
M2631 n_25 n_256 GND GND efet w=2632 l=658
+ ad=0 pd=0 as=0 ps=0 
M2632 n_51 Pout3 GND GND efet w=5828 l=564
+ ad=2.73916e+06 pd=12596 as=0 ps=0 
M2633 n_29 op_T0_sbc n_51 GND efet w=5828 l=564
+ ad=1.0347e+07 pd=30080 as=0 ps=0 
M2634 Vdd n_29 n_29 GND dfet w=846 l=1316
+ ad=0 pd=0 as=4.02922e+06 ps=11656 
M2635 n_819 pipephi2Reset0 GND GND efet w=6298 l=658
+ ad=1.11334e+07 pd=23876 as=0 ps=0 
M2636 GND pipeUNK23 n_819 GND efet w=7520 l=658
+ ad=0 pd=0 as=0 ps=0 
M2637 n_334 brk_done GND GND efet w=4277 l=611
+ ad=2.04465e+07 pd=62228 as=0 ps=0 
M2638 n_533 pipeUNK22 GND GND efet w=4136 l=658
+ ad=7.13949e+06 pd=22372 as=0 ps=0 
M2639 pipeUNK22 cclk n_29 GND efet w=1222 l=752
+ ad=2.04112e+06 pd=7520 as=0 ps=0 
M2640 n_1347 nnT2BR GND GND efet w=2914 l=658
+ ad=0 pd=0 as=0 ps=0 
M2641 GND n_223 n_1357 GND efet w=12831 l=705
+ ad=0 pd=0 as=1.59313e+07 ps=36660 
M2642 n_223 cp1 n_1215 GND efet w=1128 l=752
+ ad=1.53746e+06 pd=6956 as=3.08288e+07 ps=76704 
M2643 n_1357 n_1357 Vdd GND dfet w=940 l=752
+ ad=5.39615e+07 pd=188752 as=0 ps=0 
M2644 n_104 nnT2BR GND GND efet w=4653 l=611
+ ad=0 pd=0 as=0 ps=0 
M2645 pipephi2Reset0 cclk Reset0 GND efet w=1128 l=752
+ ad=1.23704e+06 pd=5452 as=0 ps=0 
M2646 Vdd n_819 n_819 GND dfet w=846 l=940
+ ad=0 pd=0 as=4.14585e+07 ps=150776 
M2647 n_533 n_533 Vdd GND dfet w=846 l=1786
+ ad=1.46854e+07 pd=49820 as=0 ps=0 
M2648 pipeUNK23 cclk n_1085 GND efet w=1222 l=846
+ ad=1.27238e+06 pd=6204 as=0 ps=0 
M2649 n_590 cp1 n_1178 GND efet w=1128 l=658
+ ad=1.69651e+06 pd=7520 as=0 ps=0 
M2650 GND op_ANDS op_SUMS GND efet w=2632 l=658
+ ad=0 pd=0 as=1.2556e+07 ps=34216 
M2651 op_SUMS op_EORS GND GND efet w=2726 l=658
+ ad=0 pd=0 as=0 ps=0 
M2652 GND op_ORS op_SUMS GND efet w=4277 l=611
+ ad=0 pd=0 as=0 ps=0 
M2653 op_SUMS op_SUMS Vdd GND dfet w=846 l=1410
+ ad=2.68614e+06 pd=7708 as=0 ps=0 
M2654 op_ANDS cclk n_1574 GND efet w=1128 l=752
+ ad=0 pd=0 as=1.4491e+06 ps=7332 
M2655 n_796 cclk n_396 GND efet w=1175 l=893
+ ad=1.11334e+06 pd=6392 as=0 ps=0 
M2656 GND n_590 alucin GND efet w=6392 l=564
+ ad=0 pd=0 as=6.05266e+06 ps=20680 
M2657 op_SUMS op_SRS GND GND efet w=3102 l=564
+ ad=0 pd=0 as=0 ps=0 
M2658 notRdy0 cp1 n_1679 GND efet w=1128 l=658
+ ad=0 pd=0 as=1.74953e+06 ps=7332 
M2659 n_1262 n_1679 GND GND efet w=4136 l=658
+ ad=6.9451e+06 pd=19176 as=0 ps=0 
M2660 GND n_236 n_506 GND efet w=3619 l=611
+ ad=0 pd=0 as=0 ps=0 
M2661 GND n_46 n_1508 GND efet w=9071 l=611
+ ad=0 pd=0 as=0 ps=0 
M2662 GND op_T2_pha n_1037 GND efet w=3337 l=611
+ ad=0 pd=0 as=1.68326e+07 ps=47564 
M2663 n_824 n_824 Vdd GND dfet w=940 l=1410
+ ad=7.91617e+07 pd=277112 as=0 ps=0 
M2664 Vdd op_SRS op_SRS GND dfet w=846 l=1034
+ ad=0 pd=0 as=1.00377e+08 ps=378256 
M2665 op_SRS n_366 GND GND efet w=3102 l=564
+ ad=0 pd=0 as=0 ps=0 
M2666 n_1280 op_sta_cmp n_1037 GND efet w=5076 l=564
+ ad=3.49022e+06 pd=11844 as=0 ps=0 
M2667 GND n_335 n_1280 GND efet w=5311 l=611
+ ad=0 pd=0 as=0 ps=0 
M2668 n_1225 op_T2_ind GND GND efet w=4277 l=611
+ ad=1.50124e+07 pd=56212 as=0 ps=0 
M2669 n_272 op_T2_abs_access GND GND efet w=5123 l=705
+ ad=1.9722e+07 pd=69748 as=0 ps=0 
M2670 GND op_T5_rts n_272 GND efet w=3384 l=658
+ ad=0 pd=0 as=0 ps=0 
M2671 n_256 op_T4 GND GND efet w=4277 l=611
+ ad=0 pd=0 as=0 ps=0 
M2672 GND op_T3 n_256 GND efet w=3854 l=658
+ ad=0 pd=0 as=0 ps=0 
M2673 n_726 op_T5_ind_x GND GND efet w=3995 l=611
+ ad=1.38902e+07 pd=47188 as=0 ps=0 
M2674 n_256 op_T0_brk_rti GND GND efet w=4042 l=658
+ ad=0 pd=0 as=0 ps=0 
M2675 n_1225 n_1225 Vdd GND dfet w=940 l=846
+ ad=1.11466e+08 pd=402508 as=0 ps=0 
M2676 n_272 n_272 Vdd GND dfet w=846 l=1222
+ ad=7.01667e+07 pd=245528 as=0 ps=0 
M2677 GND op_T2_zp_zp_idx n_1225 GND efet w=6016 l=658
+ ad=0 pd=0 as=0 ps=0 
M2678 n_636 op_T2_branch GND GND efet w=2350 l=658
+ ad=4.55938e+06 pd=14664 as=0 ps=0 
M2679 n_256 op_T5_rts GND GND efet w=3290 l=658
+ ad=0 pd=0 as=0 ps=0 
M2680 GND op_T0_jmp n_256 GND efet w=3948 l=564
+ ad=0 pd=0 as=0 ps=0 
M2681 GND op_T3_abs_idx_ind n_726 GND efet w=3572 l=564
+ ad=0 pd=0 as=0 ps=0 
M2682 n_256 op_T5_ind_x GND GND efet w=3619 l=611
+ ad=0 pd=0 as=0 ps=0 
M2683 n_726 n_726 Vdd GND dfet w=846 l=1222
+ ad=1.18756e+07 pd=43240 as=0 ps=0 
M2684 n_256 n_256 Vdd GND dfet w=940 l=1410
+ ad=3.98062e+07 pd=153972 as=0 ps=0 
M2685 GND Reset0 n_501 GND efet w=5170 l=564
+ ad=0 pd=0 as=1.69209e+07 ps=49444 
M2686 pipeUNK34 cclk n_824 GND efet w=1034 l=752
+ ad=1.43143e+06 pd=7144 as=0 ps=0 
M2687 n_1215 brk_done GND GND efet w=15087 l=611
+ ad=0 pd=0 as=0 ps=0 
M2688 n_272 n_236 GND GND efet w=2961 l=705
+ ad=0 pd=0 as=0 ps=0 
M2689 n_720 pipeUNK34 GND GND efet w=6533 l=611
+ ad=1.52156e+07 pd=41924 as=0 ps=0 
M2690 n_636 n_636 Vdd GND dfet w=987 l=1551
+ ad=1.1045e+07 pd=37224 as=0 ps=0 
M2691 GND pipeUNK35 n_238 GND efet w=5593 l=611
+ ad=0 pd=0 as=8.58859e+06 ps=26696 
M2692 n_261 x_op_T4_ind_y GND GND efet w=3384 l=564
+ ad=5.69038e+06 pd=23124 as=0 ps=0 
M2693 GND x_op_T3_abs_idx n_261 GND efet w=3572 l=658
+ ad=0 pd=0 as=0 ps=0 
M2694 n_726 x_op_T4_ind_y GND GND efet w=3478 l=564
+ ad=0 pd=0 as=0 ps=0 
M2695 n_134 op_brk_rti GND GND efet w=3572 l=658
+ ad=9.93166e+06 pd=24064 as=0 ps=0 
M2696 GND op_jsr n_134 GND efet w=2538 l=564
+ ad=0 pd=0 as=0 ps=0 
M2697 n_261 n_261 Vdd GND dfet w=940 l=1316
+ ad=1.18579e+07 pd=43616 as=0 ps=0 
M2698 n_501 cclk pipeUNK35 GND efet w=1034 l=658
+ ad=0 pd=0 as=1.21937e+06 ps=5452 
M2699 n_726 op_T5_rts GND GND efet w=3102 l=658
+ ad=0 pd=0 as=0 ps=0 
M2700 n_238 n_238 Vdd GND dfet w=940 l=1504
+ ad=1.62052e+07 pd=53580 as=0 ps=0 
M2701 Vdd nnT2BR nnT2BR GND dfet w=987 l=987
+ ad=0 pd=0 as=7.64226e+07 ps=268276 
M2702 n_720 notRdy0 GND GND efet w=3525 l=705
+ ad=0 pd=0 as=0 ps=0 
M2703 n_272 n_862 GND GND efet w=2256 l=658
+ ad=0 pd=0 as=0 ps=0 
M2704 GND nnT2BR n_272 GND efet w=2162 l=564
+ ad=0 pd=0 as=0 ps=0 
M2705 nnT2BR n_636 GND GND efet w=3572 l=658
+ ad=1.19639e+07 pd=36848 as=0 ps=0 
M2706 n_720 n_720 Vdd GND dfet w=846 l=1222
+ ad=1.44822e+07 pd=53768 as=0 ps=0 
M2707 n_680 cclk n_1688 GND efet w=1128 l=846
+ ad=2.51826e+06 pd=10528 as=0 ps=0 
M2708 op_EORS cclk n_982 GND efet w=1034 l=658
+ ad=0 pd=0 as=1.30773e+06 ps=6768 
M2709 op_ORS cclk n_88 GND efet w=1128 l=658
+ ad=0 pd=0 as=1.4491e+06 ps=7332 
M2710 Vdd n_1089 n_1089 GND dfet w=846 l=1598
+ ad=0 pd=0 as=7.97007e+06 ps=24252 
M2711 n_1089 n_1574 GND GND efet w=5593 l=705
+ ad=6.45912e+06 pd=22184 as=0 ps=0 
M2712 Vdd n_1141 n_1141 GND dfet w=846 l=1410
+ ad=0 pd=0 as=3.83482e+06 ps=11280 
M2713 alucin alucin Vdd GND dfet w=846 l=1128
+ ad=1.14249e+07 pd=39668 as=0 ps=0 
M2714 Vdd n_1262 n_1262 GND dfet w=846 l=1598
+ ad=0 pd=0 as=1.70093e+07 ps=53956 
M2715 n_1225 cclk pipedpc28 GND efet w=1128 l=752
+ ad=0 pd=0 as=1.40492e+06 ps=6580 
M2716 n_1407 n_1262 n_933 GND efet w=5875 l=705
+ ad=4.15292e+06 pd=13536 as=7.66965e+06 ps=22372 
M2717 GND n_572 n_1407 GND efet w=6110 l=658
+ ad=0 pd=0 as=0 ps=0 
M2718 Vdd n_10 n_10 GND dfet w=846 l=1128
+ ad=0 pd=0 as=2.16129e+07 ps=82156 
M2719 n_1215 n_1215 Vdd GND dfet w=1410 l=658
+ ad=2.08971e+07 pd=80840 as=0 ps=0 
M2720 GND x_op_jmp n_134 GND efet w=3196 l=658
+ ad=0 pd=0 as=0 ps=0 
M2721 n_510 x_op_jmp GND GND efet w=3478 l=564
+ ad=1.44822e+07 pd=37788 as=0 ps=0 
M2722 GND op_store nop_store GND efet w=4606 l=658
+ ad=0 pd=0 as=6.66234e+06 ps=18612 
M2723 n_1391 op_T4_brk GND GND efet w=3666 l=658
+ ad=1.08064e+07 pd=34028 as=0 ps=0 
M2724 GND op_T2_php n_1391 GND efet w=3572 l=658
+ ad=0 pd=0 as=0 ps=0 
M2725 n_368 op_T2_php_pha GND GND efet w=2679 l=611
+ ad=1.80166e+07 pd=44932 as=0 ps=0 
M2726 GND op_T4_jmp n_368 GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M2727 n_368 op_T5_rti_rts GND GND efet w=2679 l=611
+ ad=0 pd=0 as=0 ps=0 
M2728 GND xx_op_T5_jsr n_368 GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M2729 n_368 op_T2_jmp_abs GND GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M2730 GND x_op_T3_plp_pla n_368 GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M2731 n_790 op_lsr_ror_dec_inc GND GND efet w=2538 l=658
+ ad=7.37806e+06 pd=19552 as=0 ps=0 
M2732 GND op_asl_rol n_790 GND efet w=2585 l=611
+ ad=0 pd=0 as=0 ps=0 
M2733 n_1065 op_T0_cli_sei GND GND efet w=2538 l=564
+ ad=5.93779e+06 pd=16732 as=0 ps=0 
M2734 n_134 n_134 Vdd GND dfet w=846 l=1504
+ ad=3.83659e+07 pd=150024 as=0 ps=0 
M2735 Vdd nop_store nop_store GND dfet w=940 l=1128
+ ad=0 pd=0 as=1.58253e+07 ps=55272 
M2736 GND n_726 n_630 GND efet w=5640 l=658
+ ad=0 pd=0 as=8.16446e+06 ps=24440 
M2737 Vdd short_circuit_idx_add short_circuit_idx_add GND dfet w=846 l=1034
+ ad=0 pd=0 as=1.22114e+07 ps=39856 
M2738 GND n_238 n_1215 GND efet w=16356 l=564
+ ad=0 pd=0 as=0 ps=0 
M2739 GND pipeUNK36 short_circuit_idx_add GND efet w=9588 l=658
+ ad=0 pd=0 as=1.30066e+07 ps=36472 
M2740 short_circuit_idx_add n_1137 GND GND efet w=3760 l=658
+ ad=0 pd=0 as=0 ps=0 
M2741 n_1215 short_circuit_idx_add GND GND efet w=11421 l=611
+ ad=0 pd=0 as=0 ps=0 
M2742 n_335 n_335 Vdd GND dfet w=893 l=705
+ ad=5.63914e+07 pd=204356 as=0 ps=0 
M2743 n_630 n_630 Vdd GND dfet w=940 l=940
+ ad=3.71377e+07 pd=139872 as=0 ps=0 
M2744 n_261 cclk pipeUNK36 GND efet w=1128 l=752
+ ad=0 pd=0 as=3.05726e+06 ps=7520 
M2745 short_circuit_idx_add n_916 GND GND efet w=3666 l=564
+ ad=0 pd=0 as=0 ps=0 
M2746 n_10 op_branch_done GND GND efet w=5029 l=517
+ ad=1.85733e+07 pd=56964 as=0 ps=0 
M2747 Vdd n_1211 n_1211 GND dfet w=752 l=1034
+ ad=0 pd=0 as=5.21147e+07 ps=195144 
M2748 GND op_T2_abs_access n_1211 GND efet w=4183 l=517
+ ad=0 pd=0 as=2.44492e+07 ps=73508 
M2749 n_1211 nnT2BR GND GND efet w=1786 l=752
+ ad=0 pd=0 as=0 ps=0 
M2750 GND n_1211 n_10 GND efet w=4982 l=564
+ ad=0 pd=0 as=0 ps=0 
M2751 n_1211 nnT2BR GND GND efet w=1128 l=752
+ ad=0 pd=0 as=0 ps=0 
M2752 GND n_862 n_1211 GND efet w=3337 l=611
+ ad=0 pd=0 as=0 ps=0 
M2753 GND notRdy0 short_circuit_idx_add GND efet w=3666 l=752
+ ad=0 pd=0 as=0 ps=0 
M2754 GND n_1716 n_180 GND efet w=3384 l=564
+ ad=0 pd=0 as=7.36922e+06 ps=26132 
M2755 n_720 cp1 n_1338 GND efet w=1128 l=752
+ ad=0 pd=0 as=1.2017e+06 ps=6768 
M2756 n_462 n_1338 GND GND efet w=7285 l=611
+ ad=8.58859e+06 pd=29516 as=0 ps=0 
M2757 Vdd n_462 n_462 GND dfet w=846 l=1128
+ ad=0 pd=0 as=3.92053e+07 ps=141188 
M2758 Vdd n_933 n_933 GND dfet w=846 l=1128
+ ad=0 pd=0 as=1.24146e+07 ps=40420 
M2759 n_533 cp1 n_599 GND efet w=1128 l=846
+ ad=0 pd=0 as=2.3062e+06 ps=6956 
M2760 op_SUMS cclk n_415 GND efet w=1034 l=752
+ ad=0 pd=0 as=2.43874e+06 ps=9024 
M2761 op_SRS cclk n_968 GND efet w=1128 l=752
+ ad=0 pd=0 as=1.66117e+06 ps=7332 
M2762 Vdd notalucin notalucin GND dfet w=846 l=752
+ ad=0 pd=0 as=4.09637e+07 ps=153596 
M2763 Vdd n_1375 n_1375 GND dfet w=940 l=1504
+ ad=0 pd=0 as=8.43838e+06 ps=25568 
M2764 GND n_982 n_1141 GND efet w=5969 l=611
+ ad=0 pd=0 as=9.64891e+06 ps=23312 
M2765 n_1375 n_88 GND GND efet w=4324 l=564
+ ad=5.80525e+06 pd=20868 as=0 ps=0 
M2766 notalucin alucin GND GND efet w=5969 l=705
+ ad=5.38996e+06 pd=18424 as=0 ps=0 
M2767 Vdd n_1093 n_1093 GND dfet w=846 l=1598
+ ad=0 pd=0 as=3.94969e+06 ps=9964 
M2768 n_1526 n_1526 Vdd GND dfet w=846 l=1222
+ ad=4.10874e+06 pd=14100 as=0 ps=0 
M2769 GND n_968 n_1093 GND efet w=6204 l=564
+ ad=0 pd=0 as=9.92283e+06 ps=28952 
M2770 n_931 n_415 GND GND efet w=4982 l=658
+ ad=7.87288e+06 pd=29892 as=0 ps=0 
M2771 Vdd n_931 n_931 GND dfet w=940 l=1316
+ ad=0 pd=0 as=6.60933e+06 ps=23688 
M2772 GND n_680 n_1526 GND efet w=5969 l=611
+ ad=0 pd=0 as=8.50023e+06 ps=29892 
M2773 n_1089 cp1 n_1529 GND efet w=1034 l=752
+ ad=0 pd=0 as=2.51826e+06 ps=9588 
M2774 n_1141 cp1 n_101 GND efet w=1128 l=752
+ ad=0 pd=0 as=2.67731e+06 ps=7708 
M2775 n_1375 cp1 n_95 GND efet w=1128 l=752
+ ad=0 pd=0 as=2.83636e+06 ps=7896 
M2776 n_779 cclk n_805 GND efet w=1128 l=846
+ ad=0 pd=0 as=1.21053e+06 ps=6392 
M2777 n_1594 cclk n_688 GND efet w=1128 l=846
+ ad=0 pd=0 as=1.19286e+06 ps=6392 
M2778 n_1649 cclk n_1027 GND efet w=1128 l=846
+ ad=0 pd=0 as=1.16635e+06 ps=6768 
M2779 n_795 cclk n_360 GND efet w=1128 l=846
+ ad=0 pd=0 as=1.24588e+06 ps=6768 
M2780 n_604 cclk n_1477 GND efet w=1128 l=846
+ ad=0 pd=0 as=1.43143e+06 ps=6768 
M2781 n_692 n_460 GND GND efet w=5029 l=611
+ ad=7.44875e+06 pd=21432 as=0 ps=0 
M2782 Vdd n_692 n_692 GND dfet w=846 l=1222
+ ad=0 pd=0 as=9.61357e+06 ps=31772 
M2783 n_625 n_459 GND GND efet w=4982 l=564
+ ad=7.75801e+06 pd=21620 as=0 ps=0 
M2784 Vdd n_625 n_625 GND dfet w=846 l=1222
+ ad=0 pd=0 as=9.87865e+06 ps=31960 
M2785 Vdd n_355 n_355 GND dfet w=846 l=940
+ ad=0 pd=0 as=1.00907e+07 ps=36472 
M2786 GND n_621 n_355 GND efet w=6768 l=564
+ ad=0 pd=0 as=7.70499e+06 ps=19364 
M2787 GND n_43 n_692 GND efet w=2256 l=658
+ ad=0 pd=0 as=0 ps=0 
M2788 n_441 n_692 GND GND efet w=2256 l=564
+ ad=3.23398e+06 pd=10340 as=0 ps=0 
M2789 GND n_43 n_625 GND efet w=2256 l=564
+ ad=0 pd=0 as=0 ps=0 
M2790 Vdd n_543 n_543 GND dfet w=846 l=940
+ ad=0 pd=0 as=1.03823e+07 ps=36096 
M2791 GND n_339 n_543 GND efet w=6768 l=564
+ ad=0 pd=0 as=7.8287e+06 ps=19740 
M2792 n_662 n_625 GND GND efet w=2350 l=564
+ ad=3.25165e+06 pd=9964 as=0 ps=0 
M2793 n_6 n_521 GND GND efet w=4982 l=564
+ ad=7.78452e+06 pd=22184 as=0 ps=0 
M2794 Vdd n_6 n_6 GND dfet w=940 l=1222
+ ad=0 pd=0 as=9.82563e+06 ps=32148 
M2795 n_35 n_796 GND GND efet w=4982 l=564
+ ad=7.75801e+06 pd=21432 as=0 ps=0 
M2796 Vdd n_35 n_35 GND dfet w=940 l=1222
+ ad=0 pd=0 as=9.71076e+06 ps=31960 
M2797 n_1534 n_805 GND GND efet w=4982 l=564
+ ad=8.0496e+06 pd=21620 as=0 ps=0 
M2798 Vdd n_1534 n_1534 GND dfet w=846 l=1222
+ ad=0 pd=0 as=9.96701e+06 ps=32148 
M2799 n_1223 n_688 GND GND efet w=4935 l=517
+ ad=7.94356e+06 pd=21996 as=0 ps=0 
M2800 Vdd n_1223 n_1223 GND dfet w=940 l=1222
+ ad=0 pd=0 as=9.72844e+06 ps=31960 
M2801 n_476 n_1027 GND GND efet w=4982 l=564
+ ad=7.78452e+06 pd=21620 as=0 ps=0 
M2802 Vdd n_476 n_476 GND dfet w=846 l=1222
+ ad=0 pd=0 as=9.99352e+06 ps=32148 
M2803 GND n_43 n_6 GND efet w=2444 l=564
+ ad=0 pd=0 as=0 ps=0 
M2804 n_593 n_355 GND GND efet w=2350 l=564
+ ad=3.07493e+06 pd=10152 as=0 ps=0 
M2805 n_441 n_441 Vdd GND dfet w=940 l=1316
+ ad=1.02498e+07 pd=34028 as=0 ps=0 
M2806 Vdd n_692 dpc1_SBY GND dfet w=940 l=940
+ ad=0 pd=0 as=1.57281e+07 ps=31396 
M2807 n_662 n_662 Vdd GND dfet w=940 l=1222
+ ad=1.00112e+07 pd=33276 as=0 ps=0 
M2808 n_196 n_543 GND GND efet w=2350 l=564
+ ad=3.18096e+06 pd=9776 as=0 ps=0 
M2809 Vdd n_625 dpc3_SBX GND dfet w=846 l=940
+ ad=0 pd=0 as=1.541e+07 ps=31960 
M2810 n_593 n_593 Vdd GND dfet w=846 l=1222
+ ad=1.002e+07 pd=34216 as=0 ps=0 
M2811 n_282 n_6 GND GND efet w=2350 l=564
+ ad=3.25165e+06 pd=10152 as=0 ps=0 
M2812 GND n_43 n_35 GND efet w=2350 l=658
+ ad=0 pd=0 as=0 ps=0 
M2813 Vdd n_355 dpc4_SSB GND dfet w=940 l=846
+ ad=0 pd=0 as=1.20258e+07 ps=29704 
M2814 n_196 n_196 Vdd GND dfet w=846 l=1316
+ ad=1.0347e+07 pd=34028 as=0 ps=0 
M2815 dpc1_SBY n_1247 GND GND efet w=7003 l=611
+ ad=0 pd=0 as=0 ps=0 
M2816 GND n_441 dpc1_SBY GND efet w=7238 l=564
+ ad=0 pd=0 as=0 ps=0 
M2817 dpc3_SBX n_1247 GND GND efet w=7144 l=658
+ ad=0 pd=0 as=0 ps=0 
M2818 GND n_662 dpc3_SBX GND efet w=7238 l=564
+ ad=0 pd=0 as=0 ps=0 
M2819 GND n_593 dpc4_SSB GND efet w=9212 l=564
+ ad=0 pd=0 as=0 ps=0 
M2820 Vdd n_543 dpc5_SADL GND dfet w=940 l=752
+ ad=0 pd=0 as=1.17342e+07 ps=29516 
M2821 n_71 n_35 GND GND efet w=2350 l=564
+ ad=3.45488e+06 pd=10528 as=0 ps=0 
M2822 GND n_43 n_1534 GND efet w=2350 l=564
+ ad=0 pd=0 as=0 ps=0 
M2823 n_1230 n_360 GND GND efet w=4982 l=564
+ ad=7.76684e+06 pd=21808 as=0 ps=0 
M2824 Vdd n_1230 n_1230 GND dfet w=1034 l=1222
+ ad=0 pd=0 as=9.7196e+06 ps=31772 
M2825 n_1541 n_1477 GND GND efet w=4982 l=564
+ ad=7.79335e+06 pd=21808 as=0 ps=0 
M2826 Vdd n_1541 n_1541 GND dfet w=940 l=1222
+ ad=0 pd=0 as=9.63124e+06 ps=31772 
M2827 n_91 n_1529 GND GND efet w=7191 l=611
+ ad=6.61816e+06 pd=20492 as=0 ps=0 
M2828 Vdd n_91 n_91 GND dfet w=940 l=1034
+ ad=0 pd=0 as=1.26885e+07 ps=44368 
M2829 n_282 n_282 Vdd GND dfet w=846 l=1222
+ ad=1.00024e+07 pd=33464 as=0 ps=0 
M2830 GND n_196 dpc5_SADL GND efet w=9118 l=564
+ ad=0 pd=0 as=0 ps=0 
M2831 Vdd n_6 dpc6_SBS GND dfet w=940 l=846
+ ad=0 pd=0 as=1.70623e+07 ps=35344 
M2832 n_763 n_1534 GND GND efet w=2256 l=564
+ ad=3.29583e+06 pd=10340 as=0 ps=0 
M2833 GND n_43 n_1223 GND efet w=2256 l=564
+ ad=0 pd=0 as=0 ps=0 
M2834 n_71 n_71 Vdd GND dfet w=940 l=1222
+ ad=1.00465e+07 pd=33464 as=0 ps=0 
M2835 Vdd n_35 dpc7_SS GND dfet w=940 l=940
+ ad=0 pd=0 as=1.89709e+07 ps=40044 
M2836 n_225 n_1223 GND GND efet w=2350 l=564
+ ad=3.4107e+06 pd=10340 as=0 ps=0 
M2837 GND n_43 n_476 GND efet w=2256 l=564
+ ad=0 pd=0 as=0 ps=0 
M2838 n_763 n_763 Vdd GND dfet w=940 l=1222
+ ad=9.97584e+06 pd=33464 as=0 ps=0 
M2839 Vdd n_1534 dpc8_nDBADD GND dfet w=940 l=940
+ ad=0 pd=0 as=1.62671e+07 ps=32148 
M2840 dpc6_SBS n_1247 GND GND efet w=7144 l=564
+ ad=0 pd=0 as=0 ps=0 
M2841 GND n_282 dpc6_SBS GND efet w=7332 l=564
+ ad=0 pd=0 as=0 ps=0 
M2842 n_956 n_476 GND GND efet w=2350 l=564
+ ad=3.7553e+06 pd=10528 as=0 ps=0 
M2843 GND n_43 n_1230 GND efet w=2256 l=658
+ ad=0 pd=0 as=0 ps=0 
M2844 n_225 n_225 Vdd GND dfet w=846 l=1222
+ ad=1.08594e+07 pd=33276 as=0 ps=0 
M2845 Vdd n_1223 dpc9_DBADD GND dfet w=940 l=846
+ ad=0 pd=0 as=1.60638e+07 ps=32336 
M2846 dpc7_SS n_1247 GND GND efet w=7144 l=564
+ ad=0 pd=0 as=0 ps=0 
M2847 GND n_71 dpc7_SS GND efet w=7238 l=564
+ ad=0 pd=0 as=0 ps=0 
M2848 n_708 n_1230 GND GND efet w=2350 l=564
+ ad=3.58742e+06 pd=10340 as=0 ps=0 
M2849 GND n_43 n_1541 GND efet w=2350 l=564
+ ad=0 pd=0 as=0 ps=0 
M2850 Vdd n_1364 n_1364 GND dfet w=846 l=1034
+ ad=0 pd=0 as=1.19021e+07 ps=42112 
M2851 n_956 n_956 Vdd GND dfet w=940 l=1222
+ ad=9.95817e+06 pd=33088 as=0 ps=0 
M2852 Vdd n_476 dpc12_0ADD GND dfet w=846 l=940
+ ad=0 pd=0 as=1.71683e+07 ps=36284 
M2853 dpc8_nDBADD n_1247 GND GND efet w=7144 l=658
+ ad=0 pd=0 as=0 ps=0 
M2854 GND n_763 dpc8_nDBADD GND efet w=7332 l=564
+ ad=0 pd=0 as=0 ps=0 
M2855 n_491 n_1541 GND GND efet w=2350 l=564
+ ad=3.35768e+06 pd=10152 as=0 ps=0 
M2856 GND n_91 n_1256 GND efet w=2350 l=564
+ ad=0 pd=0 as=3.61392e+06 ps=12408 
M2857 n_708 n_708 Vdd GND dfet w=846 l=1222
+ ad=1.00112e+07 pd=33276 as=0 ps=0 
M2858 Vdd n_1230 dpc11_SBADD GND dfet w=940 l=940
+ ad=0 pd=0 as=2.004e+07 ps=39856 
M2859 dpc9_DBADD n_1247 GND GND efet w=7144 l=564
+ ad=0 pd=0 as=0 ps=0 
M2860 GND n_225 dpc9_DBADD GND efet w=7285 l=611
+ ad=0 pd=0 as=0 ps=0 
M2861 n_491 n_491 Vdd GND dfet w=940 l=1222
+ ad=1.00642e+07 pd=33464 as=0 ps=0 
M2862 Vdd n_1541 dpc10_ADLADD GND dfet w=846 l=940
+ ad=0 pd=0 as=1.66912e+07 ps=30268 
M2863 dpc12_0ADD n_1247 GND GND efet w=7144 l=564
+ ad=0 pd=0 as=0 ps=0 
M2864 GND n_956 dpc12_0ADD GND efet w=7238 l=564
+ ad=0 pd=0 as=0 ps=0 
M2865 dpc11_SBADD n_1247 GND GND efet w=7144 l=658
+ ad=0 pd=0 as=0 ps=0 
M2866 GND n_708 dpc11_SBADD GND efet w=7238 l=564
+ ad=0 pd=0 as=0 ps=0 
M2867 n_1256 n_1256 Vdd GND dfet w=940 l=1316
+ ad=1.34749e+07 pd=38164 as=0 ps=0 
M2868 dpc10_ADLADD n_1247 GND GND efet w=6956 l=564
+ ad=0 pd=0 as=0 ps=0 
M2869 GND n_491 dpc10_ADLADD GND efet w=7144 l=564
+ ad=0 pd=0 as=0 ps=0 
M2870 dpc15_ANDS n_1256 GND GND efet w=11891 l=705
+ ad=9.61357e+06 pd=27072 as=0 ps=0 
M2871 Vdd n_91 dpc15_ANDS GND dfet w=846 l=752
+ ad=0 pd=0 as=0 ps=0 
M2872 GND n_101 n_1364 GND efet w=7097 l=611
+ ad=0 pd=0 as=6.51213e+06 ps=19552 
M2873 n_531 n_95 GND GND efet w=7097 l=611
+ ad=6.45028e+06 pd=19364 as=0 ps=0 
M2874 Vdd n_531 n_531 GND dfet w=846 l=940
+ ad=0 pd=0 as=1.2715e+07 ps=42488 
M2875 GND n_1364 n_108 GND efet w=2256 l=564
+ ad=0 pd=0 as=3.17212e+06 ps=10152 
M2876 GND n_531 n_1255 GND efet w=2256 l=564
+ ad=0 pd=0 as=3.19863e+06 ps=10152 
M2877 n_108 n_108 Vdd GND dfet w=940 l=1316
+ ad=1.03293e+07 pd=36096 as=0 ps=0 
M2878 Vdd n_1364 dpc16_EORS GND dfet w=846 l=846
+ ad=0 pd=0 as=8.52674e+06 ps=26508 
M2879 n_1255 n_1255 Vdd GND dfet w=846 l=1316
+ ad=1.19993e+07 pd=35908 as=0 ps=0 
M2880 adl0 n_0_ADL0 GND GND efet w=1410 l=658
+ ad=2.60927e+07 pd=71064 as=0 ps=0 
M2881 nABL0 cclk n_1100 GND efet w=1128 l=752
+ ad=2.54477e+06 pd=8460 as=0 ps=0 
M2882 n_246 ADL_ABL nABL0 GND efet w=1128 l=564
+ ad=848256 pd=3760 as=0 ps=0 
M2883 n_123 cp1 n_246 GND efet w=1128 l=658
+ ad=8.03192e+06 pd=24064 as=0 ps=0 
M2884 abl0 nABL0 GND GND efet w=8836 l=658
+ ad=7.4134e+06 pd=23312 as=0 ps=0 
M2885 abl0 abl0 Vdd GND dfet w=846 l=1316
+ ad=2.51119e+07 pd=78584 as=0 ps=0 
M2886 ab0 n_855 Vdd GND efet w=10340 l=658
+ ad=0 pd=0 as=0 ps=0 
M2887 GND n_66 ab1 GND efet w=11844 l=564
+ ad=0 pd=0 as=1.43885e+08 ps=231804 
M2888 ab1 n_66 GND GND efet w=28435 l=705
+ ad=0 pd=0 as=0 ps=0 
M2889 ab1 n_66 GND GND efet w=33417 l=611
+ ad=0 pd=0 as=0 ps=0 
M2890 ab1 n_66 GND GND efet w=16074 l=658
+ ad=0 pd=0 as=0 ps=0 
M2891 GND n_842 n_1479 GND efet w=11938 l=658
+ ad=0 pd=0 as=1.37842e+07 ps=35156 
M2892 Vdd n_1479 ab1 GND efet w=6392 l=564
+ ad=0 pd=0 as=0 ps=0 
M2893 Vdd n_1479 ab1 GND efet w=22560 l=658
+ ad=0 pd=0 as=0 ps=0 
M2894 n_842 abl1 GND GND efet w=3384 l=658
+ ad=4.00271e+06 pd=12596 as=0 ps=0 
M2895 Vdd n_1479 ab1 GND efet w=22560 l=658
+ ad=0 pd=0 as=0 ps=0 
M2896 n_842 n_842 Vdd GND dfet w=940 l=1034
+ ad=1.50919e+07 pd=50948 as=0 ps=0 
M2897 GND abl1 n_66 GND efet w=14523 l=705
+ ad=0 pd=0 as=1.31833e+07 ps=37976 
M2898 n_1479 abl1 Vdd GND dfet w=1598 l=564
+ ad=0 pd=0 as=0 ps=0 
M2899 Vdd n_1479 ab1 GND efet w=22513 l=611
+ ad=0 pd=0 as=0 ps=0 
M2900 n_66 n_842 Vdd GND dfet w=1880 l=658
+ ad=0 pd=0 as=0 ps=0 
M2901 GND adl0 n_123 GND efet w=7802 l=658
+ ad=0 pd=0 as=0 ps=0 
M2902 n_123 n_123 Vdd GND dfet w=940 l=1128
+ ad=2.73032e+06 pd=7708 as=0 ps=0 
M2903 GND n_0_ADL1 adl1 GND efet w=1504 l=752
+ ad=0 pd=0 as=2.51561e+07 ps=67680 
M2904 nABL1 cclk n_66 GND efet w=1034 l=658
+ ad=2.40339e+06 pd=8460 as=0 ps=0 
M2905 n_416 ADL_ABL nABL1 GND efet w=1034 l=564
+ ad=777568 pd=3572 as=0 ps=0 
M2906 n_1016 cp1 n_416 GND efet w=1034 l=846
+ ad=8.16446e+06 pd=24628 as=0 ps=0 
M2907 abl1 nABL1 GND GND efet w=9024 l=611
+ ad=8.28817e+06 pd=23876 as=0 ps=0 
M2908 abl1 abl1 Vdd GND dfet w=940 l=1222
+ ad=2.49087e+07 pd=78960 as=0 ps=0 
M2909 ab1 n_1479 Vdd GND efet w=10434 l=658
+ ad=0 pd=0 as=0 ps=0 
M2910 GND n_642 ab2 GND efet w=11938 l=658
+ ad=0 pd=0 as=1.47499e+08 ps=233308 
M2911 GND n_951 n_1152 GND efet w=11844 l=658
+ ad=0 pd=0 as=1.50035e+07 ps=35532 
M2912 ab2 n_642 GND GND efet w=28435 l=611
+ ad=0 pd=0 as=0 ps=0 
M2913 ab2 n_642 GND GND efet w=33370 l=658
+ ad=0 pd=0 as=0 ps=0 
M2914 ab2 n_642 GND GND efet w=16074 l=658
+ ad=0 pd=0 as=0 ps=0 
M2915 n_951 abl2 GND GND efet w=3384 l=658
+ ad=3.77297e+06 pd=12596 as=0 ps=0 
M2916 Vdd n_1152 ab2 GND efet w=6392 l=564
+ ad=0 pd=0 as=0 ps=0 
M2917 Vdd n_1152 ab2 GND efet w=22607 l=611
+ ad=0 pd=0 as=0 ps=0 
M2918 n_951 n_951 Vdd GND dfet w=940 l=1034
+ ad=1.62494e+07 pd=50760 as=0 ps=0 
M2919 GND abl2 n_642 GND efet w=14617 l=705
+ ad=0 pd=0 as=1.39255e+07 ps=39292 
M2920 n_1152 abl2 Vdd GND dfet w=1598 l=564
+ ad=0 pd=0 as=0 ps=0 
M2921 n_642 n_951 Vdd GND dfet w=1974 l=658
+ ad=0 pd=0 as=0 ps=0 
M2922 GND adl1 n_1016 GND efet w=7708 l=658
+ ad=0 pd=0 as=0 ps=0 
M2923 n_1016 n_1016 Vdd GND dfet w=940 l=940
+ ad=2.20016e+06 pd=6956 as=0 ps=0 
M2924 Vdd n_564 n_564 GND dfet w=987 l=1645
+ ad=0 pd=0 as=3.33117e+06 ps=9776 
M2925 GND noty0 n_564 GND efet w=5170 l=564
+ ad=0 pd=0 as=1.30684e+07 ps=29892 
M2926 Vdd noty0 noty0 GND dfet w=940 l=1974
+ ad=0 pd=0 as=7.58129e+06 ps=23312 
M2927 noty0 y0 GND GND efet w=3384 l=658
+ ad=4.83329e+06 pd=15604 as=0 ps=0 
M2928 y0 cclk n_564 GND efet w=1128 l=846
+ ad=2.209e+06 pd=8084 as=0 ps=0 
M2929 n_564 dpc0_YSB sb0 GND efet w=1316 l=658
+ ad=0 pd=0 as=4.08135e+07 ps=105844 
M2930 y0 dpc1_SBY sb0 GND efet w=1128 l=658
+ ad=0 pd=0 as=0 ps=0 
M2931 GND n_0_ADL2 adl2 GND efet w=1504 l=658
+ ad=0 pd=0 as=2.47673e+07 ps=66740 
M2932 Vdd n_767 n_767 GND dfet w=940 l=1598
+ ad=0 pd=0 as=2.73032e+06 ps=7708 
M2933 GND noty1 n_767 GND efet w=5170 l=658
+ ad=0 pd=0 as=1.36605e+07 ps=33276 
M2934 Vdd noty1 noty1 GND dfet w=940 l=1974
+ ad=0 pd=0 as=8.54441e+06 ps=24064 
M2935 noty1 y1 GND GND efet w=3290 l=564
+ ad=5.02768e+06 pd=15980 as=0 ps=0 
M2936 y1 cclk n_767 GND efet w=1128 l=752
+ ad=2.45641e+06 pd=9212 as=0 ps=0 
M2937 n_767 dpc0_YSB sb1 GND efet w=1316 l=658
+ ad=0 pd=0 as=3.61834e+07 ps=92308 
M2938 nABL2 cclk n_642 GND efet w=1128 l=752
+ ad=2.6508e+06 pd=8648 as=0 ps=0 
M2939 n_1636 ADL_ABL nABL2 GND efet w=1128 l=564
+ ad=848256 pd=3760 as=0 ps=0 
M2940 n_935 cp1 n_1636 GND efet w=1128 l=752
+ ad=7.6343e+06 pd=24628 as=0 ps=0 
M2941 abl2 nABL2 GND GND efet w=8836 l=611
+ ad=7.86404e+06 pd=23688 as=0 ps=0 
M2942 abl2 abl2 Vdd GND dfet w=846 l=1222
+ ad=2.50942e+07 pd=78960 as=0 ps=0 
M2943 Vdd n_1152 ab2 GND efet w=22701 l=611
+ ad=0 pd=0 as=0 ps=0 
M2944 Vdd n_1152 ab2 GND efet w=22701 l=611
+ ad=0 pd=0 as=0 ps=0 
M2945 ab2 n_1152 Vdd GND efet w=10528 l=658
+ ad=0 pd=0 as=0 ps=0 
M2946 GND n_990 n_1041 GND efet w=11844 l=658
+ ad=0 pd=0 as=1.69651e+07 ps=41172 
M2947 n_990 abl3 GND GND efet w=3290 l=752
+ ad=3.62276e+06 pd=12408 as=0 ps=0 
M2948 GND n_138 ab3 GND efet w=11938 l=658
+ ad=0 pd=0 as=1.45891e+08 ps=232368 
M2949 n_990 n_990 Vdd GND dfet w=940 l=940
+ ad=1.63554e+07 pd=50760 as=0 ps=0 
M2950 GND abl3 n_138 GND efet w=14570 l=658
+ ad=0 pd=0 as=1.41288e+07 ps=39292 
M2951 n_1041 abl3 Vdd GND dfet w=1692 l=564
+ ad=0 pd=0 as=0 ps=0 
M2952 ab3 n_138 GND GND efet w=28388 l=658
+ ad=0 pd=0 as=0 ps=0 
M2953 ab3 n_138 GND GND efet w=33417 l=705
+ ad=0 pd=0 as=0 ps=0 
M2954 ab3 n_138 GND GND efet w=16074 l=658
+ ad=0 pd=0 as=0 ps=0 
M2955 n_138 n_990 Vdd GND dfet w=2068 l=752
+ ad=0 pd=0 as=0 ps=0 
M2956 GND adl2 n_935 GND efet w=7849 l=611
+ ad=0 pd=0 as=0 ps=0 
M2957 y1 dpc1_SBY sb1 GND efet w=1034 l=752
+ ad=0 pd=0 as=0 ps=0 
M2958 Vdd n_1491 n_1491 GND dfet w=940 l=1598
+ ad=0 pd=0 as=2.73032e+06 ps=7708 
M2959 Vdd n_1169 n_1169 GND dfet w=940 l=1504
+ ad=0 pd=0 as=2.59778e+06 ps=7520 
M2960 GND notx0 n_1169 GND efet w=5170 l=658
+ ad=0 pd=0 as=1.33512e+07 ps=33088 
M2961 Vdd notx0 notx0 GND dfet w=846 l=1974
+ ad=0 pd=0 as=8.56208e+06 ps=24064 
M2962 notx0 x0 GND GND efet w=3337 l=611
+ ad=4.25012e+06 pd=15416 as=0 ps=0 
M2963 x0 cclk n_1169 GND efet w=1128 l=752
+ ad=2.35038e+06 pd=8648 as=0 ps=0 
M2964 n_1169 dpc2_XSB sb0 GND efet w=1222 l=752
+ ad=0 pd=0 as=0 ps=0 
M2965 Vdd n_332 n_332 GND dfet w=940 l=1598
+ ad=0 pd=0 as=3.26932e+06 ps=9588 
M2966 n_332 dpc5_SADL adl0 GND efet w=1504 l=658
+ ad=1.73716e+07 pd=43052 as=0 ps=0 
M2967 Vdd n_983 n_983 GND dfet w=846 l=1880
+ ad=0 pd=0 as=4.31197e+06 ps=12408 
M2968 x0 dpc3_SBX sb0 GND efet w=1034 l=752
+ ad=0 pd=0 as=0 ps=0 
M2969 Vdd n_1709 n_1709 GND dfet w=940 l=1504
+ ad=0 pd=0 as=2.59778e+06 ps=7520 
M2970 GND notx1 n_1709 GND efet w=5217 l=611
+ ad=0 pd=0 as=1.29271e+07 ps=33276 
M2971 Vdd notx1 notx1 GND dfet w=940 l=1974
+ ad=0 pd=0 as=8.42071e+06 ps=24252 
M2972 notx1 x1 GND GND efet w=3290 l=658
+ ad=4.70075e+06 pd=15792 as=0 ps=0 
M2973 x1 cclk n_1709 GND efet w=1034 l=658
+ ad=2.21784e+06 pd=8836 as=0 ps=0 
M2974 n_332 dpc4_SSB sb0 GND efet w=1598 l=752
+ ad=0 pd=0 as=0 ps=0 
M2975 GND nots0 n_332 GND efet w=4230 l=658
+ ad=0 pd=0 as=0 ps=0 
M2976 n_983 s0 GND GND efet w=3008 l=658
+ ad=7.50176e+06 pd=21620 as=0 ps=0 
M2977 n_983 cclk nots0 GND efet w=1128 l=658
+ ad=0 pd=0 as=2.86286e+06 ps=9776 
M2978 n_332 dpc7_SS s0 GND efet w=1128 l=752
+ ad=0 pd=0 as=2.94239e+06 ps=7144 
M2979 s0 dpc6_SBS sb0 GND efet w=1128 l=752
+ ad=0 pd=0 as=0 ps=0 
M2980 sb0 cclk Vdd GND efet w=2256 l=658
+ ad=0 pd=0 as=0 ps=0 
M2981 Vdd n_694 n_694 GND dfet w=940 l=1598
+ ad=0 pd=0 as=3.34001e+06 ps=9588 
M2982 n_694 dpc5_SADL adl1 GND efet w=1410 l=752
+ ad=1.67619e+07 pd=42676 as=0 ps=0 
M2983 Vdd n_1711 n_1711 GND dfet w=846 l=1880
+ ad=0 pd=0 as=4.31197e+06 ps=12408 
M2984 n_1709 dpc2_XSB sb1 GND efet w=1222 l=752
+ ad=0 pd=0 as=0 ps=0 
M2985 x1 dpc3_SBX sb1 GND efet w=1034 l=752
+ ad=0 pd=0 as=0 ps=0 
M2986 GND noty2 n_1491 GND efet w=5311 l=611
+ ad=0 pd=0 as=1.3687e+07 ps=33464 
M2987 Vdd noty2 noty2 GND dfet w=846 l=1974
+ ad=0 pd=0 as=8.5179e+06 ps=24252 
M2988 noty2 y2 GND GND efet w=3525 l=705
+ ad=4.67424e+06 pd=15416 as=0 ps=0 
M2989 y2 cclk n_1491 GND efet w=1128 l=752
+ ad=2.48292e+06 pd=9024 as=0 ps=0 
M2990 n_935 n_935 Vdd GND dfet w=846 l=1034
+ ad=2.209e+06 pd=6956 as=0 ps=0 
M2991 n_1491 dpc0_YSB sb2 GND efet w=1222 l=658
+ ad=0 pd=0 as=3.52998e+07 ps=92120 
M2992 nABL3 cclk n_138 GND efet w=1128 l=752
+ ad=2.49175e+06 pd=8648 as=0 ps=0 
M2993 n_864 ADL_ABL nABL3 GND efet w=1128 l=658
+ ad=742224 pd=3572 as=0 ps=0 
M2994 n_1507 cp1 n_864 GND efet w=1128 l=752
+ ad=9.75494e+06 pd=27072 as=0 ps=0 
M2995 abl3 nABL3 GND GND efet w=8883 l=658
+ ad=7.76684e+06 pd=23500 as=0 ps=0 
M2996 abl3 abl3 Vdd GND dfet w=940 l=1316
+ ad=2.41223e+07 pd=77456 as=0 ps=0 
M2997 Vdd n_1041 ab3 GND efet w=6486 l=564
+ ad=0 pd=0 as=0 ps=0 
M2998 GND adl3 n_1507 GND efet w=8178 l=658
+ ad=0 pd=0 as=0 ps=0 
M2999 n_1507 n_1507 Vdd GND dfet w=846 l=940
+ ad=1.94392e+06 pd=6580 as=0 ps=0 
M3000 y2 dpc1_SBY sb2 GND efet w=1128 l=752
+ ad=0 pd=0 as=0 ps=0 
M3001 Vdd n_1531 n_1531 GND dfet w=940 l=1504
+ ad=0 pd=0 as=2.68614e+06 ps=7520 
M3002 GND noty3 n_1531 GND efet w=5311 l=611
+ ad=0 pd=0 as=1.31303e+07 ps=33652 
M3003 Vdd noty3 noty3 GND dfet w=846 l=1974
+ ad=0 pd=0 as=8.5179e+06 ps=24252 
M3004 noty3 y3 GND GND efet w=3478 l=564
+ ad=4.52403e+06 pd=15416 as=0 ps=0 
M3005 y3 cclk n_1531 GND efet w=1034 l=846
+ ad=2.34154e+06 pd=9024 as=0 ps=0 
M3006 n_1531 dpc0_YSB sb3 GND efet w=1222 l=752
+ ad=0 pd=0 as=3.56179e+07 ps=92120 
M3007 y3 dpc1_SBY sb3 GND efet w=1034 l=752
+ ad=0 pd=0 as=0 ps=0 
M3008 Vdd n_1041 ab3 GND efet w=22654 l=658
+ ad=0 pd=0 as=0 ps=0 
M3009 Vdd n_1041 ab3 GND efet w=22654 l=658
+ ad=0 pd=0 as=0 ps=0 
M3010 Vdd n_1041 ab3 GND efet w=22607 l=611
+ ad=0 pd=0 as=0 ps=0 
M3011 ab3 n_1041 Vdd GND efet w=10434 l=658
+ ad=0 pd=0 as=0 ps=0 
M3012 GND n_1676 n_634 GND efet w=11844 l=658
+ ad=0 pd=0 as=1.39874e+07 ps=35344 
M3013 n_1676 abl4 GND GND efet w=3384 l=658
+ ad=4.25012e+06 pd=12596 as=0 ps=0 
M3014 n_1676 n_1676 Vdd GND dfet w=940 l=940
+ ad=1.58341e+07 pd=50948 as=0 ps=0 
M3015 GND abl4 n_86 GND efet w=14570 l=658
+ ad=0 pd=0 as=1.40934e+07 ps=39668 
M3016 n_634 abl4 Vdd GND dfet w=1692 l=564
+ ad=0 pd=0 as=0 ps=0 
M3017 n_86 n_1676 Vdd GND dfet w=2068 l=658
+ ad=0 pd=0 as=0 ps=0 
M3018 nABL4 cclk n_86 GND efet w=1128 l=752
+ ad=2.49175e+06 pd=8648 as=0 ps=0 
M3019 n_738 ADL_ABL nABL4 GND efet w=1128 l=658
+ ad=742224 pd=3572 as=0 ps=0 
M3020 n_1519 cp1 n_738 GND efet w=1128 l=752
+ ad=7.97891e+06 pd=25004 as=0 ps=0 
M3021 abl4 nABL4 GND GND efet w=8977 l=611
+ ad=7.8552e+06 pd=23876 as=0 ps=0 
M3022 abl4 abl4 Vdd GND dfet w=846 l=1316
+ ad=2.40339e+07 pd=78584 as=0 ps=0 
M3023 GND n_86 ab4 GND efet w=11844 l=658
+ ad=0 pd=0 as=1.44044e+08 ps=231804 
M3024 ab4 n_86 GND GND efet w=28294 l=658
+ ad=0 pd=0 as=0 ps=0 
M3025 ab4 n_86 GND GND efet w=33511 l=705
+ ad=0 pd=0 as=0 ps=0 
M3026 ab4 n_86 GND GND efet w=16168 l=658
+ ad=0 pd=0 as=0 ps=0 
M3027 Vdd n_634 ab4 GND efet w=6392 l=564
+ ad=0 pd=0 as=0 ps=0 
M3028 Vdd n_634 ab4 GND efet w=22419 l=705
+ ad=0 pd=0 as=0 ps=0 
M3029 Vdd n_634 ab4 GND efet w=22513 l=611
+ ad=0 pd=0 as=0 ps=0 
M3030 Vdd n_634 ab4 GND efet w=22513 l=611
+ ad=0 pd=0 as=0 ps=0 
M3031 ab4 n_634 Vdd GND efet w=10434 l=658
+ ad=0 pd=0 as=0 ps=0 
M3032 GND n_172 n_1633 GND efet w=11844 l=658
+ ad=0 pd=0 as=1.40846e+07 ps=35344 
M3033 n_172 abl5 GND GND efet w=3384 l=752
+ ad=3.62276e+06 pd=12596 as=0 ps=0 
M3034 GND n_210 ab5 GND efet w=11844 l=658
+ ad=0 pd=0 as=1.46952e+08 ps=232368 
M3035 ab5 n_210 GND GND efet w=28388 l=658
+ ad=0 pd=0 as=0 ps=0 
M3036 ab5 n_210 GND GND efet w=33652 l=658
+ ad=0 pd=0 as=0 ps=0 
M3037 ab5 n_210 GND GND efet w=16074 l=564
+ ad=0 pd=0 as=0 ps=0 
M3038 n_172 n_172 Vdd GND dfet w=1034 l=940
+ ad=1.51891e+07 pd=50760 as=0 ps=0 
M3039 GND abl5 n_210 GND efet w=14476 l=658
+ ad=0 pd=0 as=1.41995e+07 ps=37600 
M3040 n_1633 abl5 Vdd GND dfet w=1786 l=564
+ ad=0 pd=0 as=0 ps=0 
M3041 n_210 n_172 Vdd GND dfet w=1974 l=658
+ ad=0 pd=0 as=0 ps=0 
M3042 GND adl4 n_1519 GND efet w=7849 l=611
+ ad=0 pd=0 as=0 ps=0 
M3043 Vdd n_658 n_658 GND dfet w=940 l=1504
+ ad=0 pd=0 as=2.68614e+06 ps=7520 
M3044 GND noty4 n_658 GND efet w=5264 l=658
+ ad=0 pd=0 as=1.26355e+07 ps=32712 
M3045 Vdd noty4 noty4 GND dfet w=940 l=1974
+ ad=0 pd=0 as=8.6151e+06 ps=24252 
M3046 noty4 y4 GND GND efet w=3290 l=658
+ ad=4.61239e+06 pd=15604 as=0 ps=0 
M3047 y4 cclk n_658 GND efet w=1034 l=752
+ ad=2.31503e+06 pd=8460 as=0 ps=0 
M3048 n_1519 n_1519 Vdd GND dfet w=846 l=940
+ ad=1.97926e+06 pd=6768 as=0 ps=0 
M3049 n_658 dpc0_YSB sb4 GND efet w=1222 l=752
+ ad=0 pd=0 as=3.66517e+07 ps=98888 
M3050 nABL5 cclk n_210 GND efet w=1034 l=658
+ ad=2.40339e+06 pd=8460 as=0 ps=0 
M3051 n_463 ADL_ABL nABL5 GND efet w=1034 l=658
+ ad=680372 pd=3384 as=0 ps=0 
M3052 n_1094 cp1 n_463 GND efet w=1034 l=752
+ ad=8.24399e+06 pd=25192 as=0 ps=0 
M3053 abl5 nABL5 GND GND efet w=9165 l=611
+ ad=8.32351e+06 pd=23876 as=0 ps=0 
M3054 abl5 abl5 Vdd GND dfet w=940 l=1316
+ ad=2.48468e+07 pd=78584 as=0 ps=0 
M3055 Vdd n_1633 ab5 GND efet w=6486 l=564
+ ad=0 pd=0 as=0 ps=0 
M3056 Vdd n_1633 ab5 GND efet w=22654 l=658
+ ad=0 pd=0 as=0 ps=0 
M3057 Vdd n_1633 ab5 GND efet w=22560 l=658
+ ad=0 pd=0 as=0 ps=0 
M3058 Vdd n_1633 ab5 GND efet w=22513 l=611
+ ad=0 pd=0 as=0 ps=0 
M3059 ab5 n_1633 Vdd GND efet w=10434 l=658
+ ad=0 pd=0 as=0 ps=0 
M3060 GND n_1195 n_1191 GND efet w=11938 l=658
+ ad=0 pd=0 as=1.39962e+07 ps=35156 
M3061 n_1195 abl6 GND GND efet w=3384 l=658
+ ad=3.78181e+06 pd=12596 as=0 ps=0 
M3062 n_1195 n_1195 Vdd GND dfet w=940 l=1034
+ ad=1.50919e+07 pd=50948 as=0 ps=0 
M3063 GND abl6 n_1254 GND efet w=14711 l=705
+ ad=0 pd=0 as=1.33424e+07 ps=38352 
M3064 n_1191 abl6 Vdd GND dfet w=1786 l=658
+ ad=0 pd=0 as=0 ps=0 
M3065 n_1254 n_1195 Vdd GND dfet w=1880 l=658
+ ad=0 pd=0 as=0 ps=0 
M3066 GND adl5 n_1094 GND efet w=7896 l=658
+ ad=0 pd=0 as=0 ps=0 
M3067 y4 dpc1_SBY sb4 GND efet w=1128 l=752
+ ad=0 pd=0 as=0 ps=0 
M3068 Vdd n_733 n_733 GND dfet w=846 l=1598
+ ad=0 pd=0 as=2.82752e+06 ps=7708 
M3069 GND noty5 n_733 GND efet w=5358 l=658
+ ad=0 pd=0 as=1.29624e+07 ps=33088 
M3070 Vdd noty5 noty5 GND dfet w=846 l=1880
+ ad=0 pd=0 as=8.45605e+06 ps=24064 
M3071 noty5 y5 GND GND efet w=3290 l=658
+ ad=4.33848e+06 pd=15228 as=0 ps=0 
M3072 y5 cclk n_733 GND efet w=1034 l=752
+ ad=2.3327e+06 pd=8460 as=0 ps=0 
M3073 n_1094 n_1094 Vdd GND dfet w=846 l=1034
+ ad=2.35921e+06 pd=7144 as=0 ps=0 
M3074 n_733 dpc0_YSB sb5 GND efet w=1222 l=752
+ ad=0 pd=0 as=3.53793e+07 ps=92120 
M3075 y5 dpc1_SBY sb5 GND efet w=1034 l=658
+ ad=0 pd=0 as=0 ps=0 
M3076 nABL6 cclk n_1254 GND efet w=1128 l=658
+ ad=2.59778e+06 pd=8836 as=0 ps=0 
M3077 n_524 ADL_ABL nABL6 GND efet w=1128 l=658
+ ad=742224 pd=3572 as=0 ps=0 
M3078 n_1548 cp1 n_524 GND efet w=1128 l=752
+ ad=8.42071e+06 pd=24816 as=0 ps=0 
M3079 abl6 nABL6 GND GND efet w=9118 l=611
+ ad=8.08494e+06 pd=23500 as=0 ps=0 
M3080 abl6 abl6 Vdd GND dfet w=940 l=1316
+ ad=2.52091e+07 pd=78772 as=0 ps=0 
M3081 GND n_1254 ab6 GND efet w=13066 l=658
+ ad=0 pd=0 as=1.49479e+08 ps=231804 
M3082 ab6 n_1254 GND GND efet w=30550 l=658
+ ad=0 pd=0 as=0 ps=0 
M3083 ab6 n_1254 GND GND efet w=33746 l=658
+ ad=0 pd=0 as=0 ps=0 
M3084 GND n_1026 n_322 GND efet w=11797 l=611
+ ad=0 pd=0 as=1.55602e+07 ps=36660 
M3085 n_1026 abl7 GND GND efet w=3384 l=658
+ ad=3.84366e+06 pd=12596 as=0 ps=0 
M3086 Vdd n_1191 ab6 GND efet w=11656 l=658
+ ad=0 pd=0 as=0 ps=0 
M3087 ab6 n_1254 GND GND efet w=19787 l=611
+ ad=0 pd=0 as=0 ps=0 
M3088 Vdd n_1191 ab6 GND efet w=22466 l=658
+ ad=0 pd=0 as=0 ps=0 
M3089 Vdd n_1191 ab6 GND efet w=22513 l=611
+ ad=0 pd=0 as=0 ps=0 
M3090 Vdd n_1191 ab6 GND efet w=23500 l=658
+ ad=0 pd=0 as=0 ps=0 
M3091 n_1026 n_1026 Vdd GND dfet w=1034 l=940
+ ad=1.49505e+07 pd=50384 as=0 ps=0 
M3092 GND abl7 n_171 GND efet w=14617 l=705
+ ad=0 pd=0 as=1.38637e+07 ps=38916 
M3093 n_322 abl7 Vdd GND dfet w=1739 l=705
+ ad=0 pd=0 as=0 ps=0 
M3094 n_171 n_1026 Vdd GND dfet w=1880 l=658
+ ad=0 pd=0 as=0 ps=0 
M3095 GND adl6 n_1548 GND efet w=7802 l=564
+ ad=0 pd=0 as=0 ps=0 
M3096 Vdd n_518 n_518 GND dfet w=940 l=1504
+ ad=0 pd=0 as=2.68614e+06 ps=7520 
M3097 Vdd n_1694 n_1694 GND dfet w=940 l=1598
+ ad=0 pd=0 as=2.73032e+06 ps=7708 
M3098 GND notx2 n_1694 GND efet w=5311 l=611
+ ad=0 pd=0 as=1.31215e+07 ps=33464 
M3099 Vdd notx2 notx2 GND dfet w=940 l=1974
+ ad=0 pd=0 as=8.36769e+06 ps=24064 
M3100 n_694 dpc4_SSB sb1 GND efet w=1598 l=658
+ ad=0 pd=0 as=0 ps=0 
M3101 notx2 x2 GND GND efet w=3384 l=658
+ ad=4.74493e+06 pd=15604 as=0 ps=0 
M3102 x2 cclk n_1694 GND efet w=1128 l=846
+ ad=2.35038e+06 pd=9024 as=0 ps=0 
M3103 GND nots1 n_694 GND efet w=4042 l=564
+ ad=0 pd=0 as=0 ps=0 
M3104 n_1711 s1 GND GND efet w=3008 l=658
+ ad=7.7315e+06 pd=21808 as=0 ps=0 
M3105 n_1711 cclk nots1 GND efet w=1128 l=752
+ ad=0 pd=0 as=2.46524e+06 ps=9400 
M3106 n_694 dpc7_SS s1 GND efet w=1128 l=846
+ ad=0 pd=0 as=3.02191e+06 ps=7144 
M3107 s1 dpc6_SBS sb1 GND efet w=1222 l=752
+ ad=0 pd=0 as=0 ps=0 
M3108 sb1 cclk Vdd GND efet w=2256 l=658
+ ad=0 pd=0 as=0 ps=0 
M3109 Vdd n_1389 n_1389 GND dfet w=940 l=1598
+ ad=0 pd=0 as=3.28699e+06 ps=9588 
M3110 n_1389 dpc5_SADL adl2 GND efet w=1504 l=470
+ ad=1.69209e+07 pd=43428 as=0 ps=0 
M3111 Vdd n_1190 n_1190 GND dfet w=846 l=1880
+ ad=0 pd=0 as=4.25895e+06 ps=12220 
M3112 n_1694 dpc2_XSB sb2 GND efet w=1222 l=752
+ ad=0 pd=0 as=0 ps=0 
M3113 x2 dpc3_SBX sb2 GND efet w=1128 l=752
+ ad=0 pd=0 as=0 ps=0 
M3114 Vdd n_242 n_242 GND dfet w=940 l=1504
+ ad=0 pd=0 as=2.59778e+06 ps=7520 
M3115 GND notx3 n_242 GND efet w=5217 l=611
+ ad=0 pd=0 as=1.40227e+07 ps=33276 
M3116 Vdd notx3 notx3 GND dfet w=846 l=1974
+ ad=0 pd=0 as=8.36769e+06 ps=24064 
M3117 notx3 x3 GND GND efet w=3384 l=564
+ ad=4.92165e+06 pd=15792 as=0 ps=0 
M3118 x3 cclk n_242 GND efet w=1128 l=752
+ ad=2.5536e+06 pd=9024 as=0 ps=0 
M3119 n_242 dpc2_XSB sb3 GND efet w=1222 l=752
+ ad=0 pd=0 as=0 ps=0 
M3120 n_1389 dpc4_SSB sb2 GND efet w=1598 l=752
+ ad=0 pd=0 as=0 ps=0 
M3121 GND nots2 n_1389 GND efet w=4136 l=658
+ ad=0 pd=0 as=0 ps=0 
M3122 n_1190 s2 GND GND efet w=3102 l=658
+ ad=7.72266e+06 pd=21620 as=0 ps=0 
M3123 n_1190 cclk nots2 GND efet w=1128 l=752
+ ad=0 pd=0 as=2.40339e+06 ps=9400 
M3124 GND n_108 dpc16_EORS GND efet w=10481 l=517
+ ad=0 pd=0 as=0 ps=0 
M3125 dpc13_ORS n_1255 GND GND efet w=10434 l=658
+ ad=8.43838e+06 pd=24440 as=0 ps=0 
M3126 Vdd n_531 dpc13_ORS GND dfet w=846 l=846
+ ad=0 pd=0 as=0 ps=0 
M3127 GND pipedpc28 dpc28_0ADH0 GND efet w=8883 l=611
+ ad=0 pd=0 as=9.08341e+06 ps=25944 
M3128 n_877 n_506 GND GND efet w=5311 l=611
+ ad=9.82563e+06 pd=31208 as=0 ps=0 
M3129 Vdd dpc28_0ADH0 dpc28_0ADH0 GND dfet w=893 l=1551
+ ad=0 pd=0 as=3.67578e+07 ps=142880 
M3130 n_674 n_674 Vdd GND dfet w=893 l=1081
+ ad=5.92896e+06 pd=22560 as=0 ps=0 
M3131 Vdd dpc22_nDSA dpc22_nDSA GND dfet w=846 l=1128
+ ad=0 pd=0 as=5.99346e+07 ps=253988 
M3132 n_674 n_25 GND GND efet w=4747 l=611
+ ad=8.2705e+06 pd=30268 as=0 ps=0 
M3133 n_80 n_267 GND GND efet w=3572 l=658
+ ad=8.19097e+06 pd=23500 as=0 ps=0 
M3134 GND n_1130 n_80 GND efet w=4371 l=517
+ ad=0 pd=0 as=0 ps=0 
M3135 GND n_599 dpc22_nDSA GND efet w=7473 l=611
+ ad=0 pd=0 as=5.90245e+06 ps=19740 
M3136 Vdd n_80 n_80 GND dfet w=752 l=940
+ ad=0 pd=0 as=2.03228e+06 ps=6768 
M3137 n_1245 n_1245 Vdd GND dfet w=987 l=799
+ ad=2.78864e+07 pd=97948 as=0 ps=0 
M3138 n_1245 aluvout GND GND efet w=6956 l=611
+ ad=8.03192e+06 pd=23500 as=0 ps=0 
M3139 GND n_933 n_877 GND efet w=4606 l=658
+ ad=0 pd=0 as=0 ps=0 
M3140 n_1211 n_1002 GND GND efet w=3431 l=611
+ ad=0 pd=0 as=0 ps=0 
M3141 n_182 n_182 Vdd GND dfet w=940 l=1128
+ ad=3.31615e+07 pd=122952 as=0 ps=0 
M3142 GND op_T5_rts n_182 GND efet w=2726 l=564
+ ad=0 pd=0 as=2.54654e+07 ps=75012 
M3143 n_1151 n_1262 GND GND efet w=6392 l=564
+ ad=3.6581e+06 pd=14100 as=0 ps=0 
M3144 GND n_467 n_10 GND efet w=2632 l=564
+ ad=0 pd=0 as=0 ps=0 
M3145 n_182 n_236 n_1151 GND efet w=6439 l=611
+ ad=0 pd=0 as=0 ps=0 
M3146 GND n_1286 n_1211 GND efet w=4230 l=658
+ ad=0 pd=0 as=0 ps=0 
M3147 Vdd n_467 n_467 GND dfet w=846 l=1316
+ ad=0 pd=0 as=1.07446e+07 ps=36284 
M3148 GND nnT2BR n_1427 GND efet w=4324 l=658
+ ad=0 pd=0 as=1.13189e+07 ps=37600 
M3149 n_1427 n_1427 Vdd GND dfet w=846 l=1598
+ ad=1.70005e+07 pd=61288 as=0 ps=0 
M3150 n_930 n_930 Vdd GND dfet w=846 l=1598
+ ad=1.23969e+07 pd=40796 as=0 ps=0 
M3151 n_930 n_134 GND GND efet w=3196 l=564
+ ad=1.05148e+07 pd=33840 as=0 ps=0 
M3152 n_1705 n_467 GND GND efet w=3055 l=564
+ ad=1.18137e+07 pd=35532 as=0 ps=0 
M3153 n_877 n_877 Vdd GND dfet w=846 l=940
+ ad=8.3942e+06 pd=29140 as=0 ps=0 
M3154 n_1093 cp1 n_226 GND efet w=1128 l=752
+ ad=0 pd=0 as=2.47408e+06 ps=7520 
M3155 n_931 cp1 n_1674 GND efet w=1128 l=752
+ ad=0 pd=0 as=2.59778e+06 ps=7708 
M3156 n_1526 cp1 n_1450 GND efet w=1128 l=752
+ ad=0 pd=0 as=2.79218e+06 ps=10528 
M3157 n_80 cclk n_1333 GND efet w=1128 l=846
+ ad=0 pd=0 as=1.67e+06 ps=7332 
M3158 n_1130 cclk n_512 GND efet w=1175 l=893
+ ad=0 pd=0 as=1.88207e+06 ps=7708 
M3159 n_674 cclk n_745 GND efet w=1128 l=846
+ ad=0 pd=0 as=1.61699e+06 ps=5828 
M3160 Vdd n_1593 n_1593 GND dfet w=846 l=1128
+ ad=0 pd=0 as=1.31833e+07 ps=43428 
M3161 GND n_226 n_1593 GND efet w=6956 l=658
+ ad=0 pd=0 as=6.3089e+06 ps=19176 
M3162 n_772 n_1674 GND GND efet w=6909 l=611
+ ad=5.60202e+06 pd=20680 as=0 ps=0 
M3163 Vdd n_772 n_772 GND dfet w=846 l=1034
+ ad=0 pd=0 as=1.15221e+07 ps=42488 
M3164 GND n_1593 n_1552 GND efet w=2256 l=564
+ ad=0 pd=0 as=3.04842e+06 ps=9964 
M3165 GND n_772 n_1305 GND efet w=2256 l=564
+ ad=0 pd=0 as=3.33117e+06 ps=10340 
M3166 n_1552 n_1552 Vdd GND dfet w=752 l=1316
+ ad=1.23085e+07 pd=37224 as=0 ps=0 
M3167 Vdd n_1593 dpc14_SRS GND dfet w=752 l=846
+ ad=0 pd=0 as=7.6343e+06 ps=21808 
M3168 n_1305 n_1305 Vdd GND dfet w=940 l=1316
+ ad=1.2176e+07 pd=37788 as=0 ps=0 
M3169 dpc14_SRS n_1552 GND GND efet w=11327 l=611
+ ad=0 pd=0 as=0 ps=0 
M3170 dpc17_SUMS n_1305 GND GND efet w=11468 l=658
+ ad=9.65775e+06 pd=30268 as=0 ps=0 
M3171 Vdd n_772 dpc17_SUMS GND dfet w=1034 l=846
+ ad=0 pd=0 as=0 ps=0 
M3172 Vdd n_1499 n_1499 GND dfet w=846 l=1128
+ ad=0 pd=0 as=1.15752e+07 ps=42300 
M3173 GND n_1450 n_1499 GND efet w=7191 l=611
+ ad=0 pd=0 as=7.22785e+06 ps=20868 
M3174 n_906 n_1333 GND GND efet w=7144 l=564
+ ad=7.27203e+06 pd=21244 as=0 ps=0 
M3175 Vdd n_906 n_906 GND dfet w=846 l=940
+ ad=0 pd=0 as=1.72302e+07 ps=59408 
M3176 Vdd n_154 n_154 GND dfet w=846 l=1128
+ ad=0 pd=0 as=1.13896e+07 ps=41924 
M3177 n_714 n_906 GND GND efet w=4089 l=517
+ ad=4.34731e+06 pd=13348 as=0 ps=0 
M3178 GND n_1499 n_709 GND efet w=2256 l=564
+ ad=0 pd=0 as=3.11027e+06 ps=10152 
M3179 GND n_512 n_154 GND efet w=6956 l=658
+ ad=0 pd=0 as=5.85827e+06 ps=20492 
M3180 n_241 n_745 GND GND efet w=6909 l=611
+ ad=6.02615e+06 pd=19176 as=0 ps=0 
M3181 Vdd n_241 n_241 GND dfet w=752 l=940
+ ad=0 pd=0 as=1.25294e+07 ps=42300 
M3182 GND n_154 n_75 GND efet w=2350 l=564
+ ad=0 pd=0 as=3.32234e+06 ps=10528 
M3183 GND n_241 n_1033 GND efet w=2256 l=564
+ ad=0 pd=0 as=2.9689e+06 ps=9776 
M3184 n_709 n_709 Vdd GND dfet w=846 l=1316
+ ad=1.16105e+07 pd=37976 as=0 ps=0 
M3185 Vdd n_1499 dpc18_nDAA GND dfet w=846 l=846
+ ad=0 pd=0 as=1.11599e+07 ps=33088 
M3186 n_714 n_714 Vdd GND dfet w=846 l=1410
+ ad=6.22938e+06 pd=17860 as=0 ps=0 
M3187 adl0 dpc10_ADLADD alub0 GND efet w=1034 l=658
+ ad=0 pd=0 as=4.96583e+06 ps=13536 
M3188 alub0 dpc8_nDBADD n_624 GND efet w=1034 l=658
+ ad=0 pd=0 as=7.81102e+06 ps=25756 
M3189 alub0 dpc9_DBADD idb0 GND efet w=1034 l=658
+ ad=0 pd=0 as=1.87942e+07 ps=52452 
M3190 GND idb0 n_624 GND efet w=5687 l=705
+ ad=0 pd=0 as=0 ps=0 
M3191 n_624 n_624 Vdd GND dfet w=940 l=1692
+ ad=3.16329e+06 pd=8272 as=0 ps=0 
M3192 n_316 alua0 GND GND efet w=5734 l=564
+ ad=2.69498e+06 pd=12408 as=0 ps=0 
M3193 nA_B0 alub0 n_316 GND efet w=5734 l=658
+ ad=9.26896e+06 pd=27260 as=0 ps=0 
M3194 Vdd nA_B0 nA_B0 GND dfet w=987 l=2115
+ ad=0 pd=0 as=2.21519e+07 ps=72568 
M3195 naluresult0 dpc13_ORS n_A_B_0 GND efet w=1222 l=752
+ ad=1.44115e+07 pd=41736 as=9.48986e+06 ps=27072 
M3196 GND dpc12_0ADD alua0 GND efet w=1222 l=564
+ ad=0 pd=0 as=4.90398e+06 ps=13536 
M3197 alua0 dpc11_SBADD sb0 GND efet w=1128 l=752
+ ad=0 pd=0 as=0 ps=0 
M3198 adl1 dpc10_ADLADD alub1 GND efet w=1034 l=658
+ ad=0 pd=0 as=5.11604e+06 ps=13536 
M3199 alub1 dpc8_nDBADD n_583 GND efet w=1128 l=752
+ ad=0 pd=0 as=8.66812e+06 ps=26132 
M3200 alub1 dpc9_DBADD idb1 GND efet w=1128 l=658
+ ad=0 pd=0 as=1.89002e+07 ps=51888 
M3201 GND idb1 n_583 GND efet w=5781 l=705
+ ad=0 pd=0 as=0 ps=0 
M3202 n_583 n_583 Vdd GND dfet w=799 l=1645
+ ad=2.93355e+06 pd=8084 as=0 ps=0 
M3203 n_A_B_0 alua0 GND GND efet w=3008 l=564
+ ad=0 pd=0 as=0 ps=0 
M3204 GND alub0 n_A_B_0 GND efet w=3008 l=658
+ ad=0 pd=0 as=0 ps=0 
M3205 Vdd n_A_B_0 n_A_B_0 GND dfet w=940 l=2162
+ ad=0 pd=0 as=2.10032e+07 ps=71816 
M3206 n_189 alua1 GND GND efet w=5734 l=564
+ ad=3.23398e+06 pd=12596 as=0 ps=0 
M3207 nA_B1 alub1 n_189 GND efet w=5734 l=564
+ ad=9.80796e+06 pd=27824 as=0 ps=0 
M3208 Vdd nA_B1 nA_B1 GND dfet w=846 l=2068
+ ad=0 pd=0 as=8.23515e+06 ps=22748 
M3209 GND n_709 dpc18_nDAA GND efet w=11515 l=611
+ ad=0 pd=0 as=0 ps=0 
M3210 dpc19_ADDSB7 n_906 GND GND efet w=10763 l=611
+ ad=9.0569e+06 pd=29140 as=0 ps=0 
M3211 Vdd n_714 dpc19_ADDSB7 GND dfet w=940 l=846
+ ad=0 pd=0 as=0 ps=0 
M3212 n_75 n_75 Vdd GND dfet w=846 l=1316
+ ad=1.14426e+07 pd=36848 as=0 ps=0 
M3213 Vdd n_154 dpc20_ADDSB06 GND dfet w=846 l=846
+ ad=0 pd=0 as=9.79029e+06 ps=30268 
M3214 n_1033 n_1033 Vdd GND dfet w=846 l=1410
+ ad=1.17784e+07 pd=35532 as=0 ps=0 
M3215 GND n_75 dpc20_ADDSB06 GND efet w=11139 l=611
+ ad=0 pd=0 as=0 ps=0 
M3216 dpc21_ADDADL n_1033 GND GND efet w=10481 l=611
+ ad=8.89785e+06 pd=28388 as=0 ps=0 
M3217 Vdd n_241 dpc21_ADDADL GND dfet w=846 l=752
+ ad=0 pd=0 as=0 ps=0 
M3218 A_B0 A_B0 Vdd GND dfet w=940 l=1410
+ ad=7.83753e+06 pd=24628 as=0 ps=0 
M3219 Vdd n_105 n_105 GND dfet w=940 l=1504
+ ad=0 pd=0 as=1.07622e+07 ps=32336 
M3220 n_105 notalucin GND GND efet w=1692 l=564
+ ad=2.80985e+06 pd=9212 as=0 ps=0 
M3221 A_B0 n_A_B_0 GND GND efet w=1692 l=564
+ ad=2.9689e+06 pd=8648 as=0 ps=0 
M3222 n_1348 A_B0 n_AxB_0 GND efet w=3431 l=611
+ ad=1.67e+06 pd=7708 as=6.79488e+06 ps=22184 
M3223 naluresult0 dpc15_ANDS nA_B0 GND efet w=1034 l=752
+ ad=0 pd=0 as=0 ps=0 
M3224 n_AxB_0 dpc16_EORS naluresult0 GND efet w=1034 l=752
+ ad=0 pd=0 as=0 ps=0 
M3225 nA_B1 dpc14_SRS naluresult0 GND efet w=1034 l=752
+ ad=0 pd=0 as=0 ps=0 
M3226 naluresult1 dpc13_ORS n_A_B_1 GND efet w=1128 l=752
+ ad=1.66382e+07 pd=47000 as=9.375e+06 ps=26508 
M3227 GND dpc12_0ADD alua1 GND efet w=1128 l=564
+ ad=0 pd=0 as=4.97467e+06 ps=13160 
M3228 alua1 dpc11_SBADD sb1 GND efet w=1175 l=893
+ ad=0 pd=0 as=0 ps=0 
M3229 n_1389 dpc7_SS s2 GND efet w=1128 l=658
+ ad=0 pd=0 as=3.04842e+06 ps=7332 
M3230 s2 dpc6_SBS sb2 GND efet w=1128 l=752
+ ad=0 pd=0 as=0 ps=0 
M3231 sb2 cclk Vdd GND efet w=2162 l=658
+ ad=0 pd=0 as=0 ps=0 
M3232 Vdd n_998 n_998 GND dfet w=846 l=1504
+ ad=0 pd=0 as=3.20747e+06 ps=9588 
M3233 n_998 dpc5_SADL adl3 GND efet w=1410 l=611
+ ad=1.75748e+07 pd=43616 as=2.2196e+07 ps=59032 
M3234 Vdd n_34 n_34 GND dfet w=846 l=1880
+ ad=0 pd=0 as=4.25895e+06 ps=12220 
M3235 x3 dpc3_SBX sb3 GND efet w=1128 l=658
+ ad=0 pd=0 as=0 ps=0 
M3236 Vdd n_436 n_436 GND dfet w=940 l=1504
+ ad=0 pd=0 as=2.68614e+06 ps=7520 
M3237 n_998 dpc4_SSB sb3 GND efet w=1504 l=658
+ ad=0 pd=0 as=0 ps=0 
M3238 GND notx4 n_436 GND efet w=5264 l=658
+ ad=0 pd=0 as=1.28475e+07 ps=33088 
M3239 Vdd notx4 notx4 GND dfet w=940 l=1974
+ ad=0 pd=0 as=8.6151e+06 ps=24252 
M3240 notx4 x4 GND GND efet w=3290 l=564
+ ad=4.63006e+06 pd=15604 as=0 ps=0 
M3241 x4 cclk n_436 GND efet w=1034 l=752
+ ad=2.31503e+06 pd=8648 as=0 ps=0 
M3242 GND nots3 n_998 GND efet w=4136 l=564
+ ad=0 pd=0 as=0 ps=0 
M3243 n_34 s3 GND GND efet w=3196 l=564
+ ad=8.12028e+06 pd=21432 as=0 ps=0 
M3244 n_34 cclk nots3 GND efet w=1034 l=752
+ ad=0 pd=0 as=2.5536e+06 ps=9400 
M3245 n_998 dpc7_SS s3 GND efet w=1034 l=752
+ ad=0 pd=0 as=2.95122e+06 ps=7144 
M3246 s3 dpc6_SBS sb3 GND efet w=1128 l=658
+ ad=0 pd=0 as=0 ps=0 
M3247 sb3 cclk Vdd GND efet w=2115 l=611
+ ad=0 pd=0 as=0 ps=0 
M3248 Vdd n_3 n_3 GND dfet w=846 l=1598
+ ad=0 pd=0 as=3.16329e+06 ps=9400 
M3249 n_3 dpc5_SADL adl4 GND efet w=1316 l=658
+ ad=1.71683e+07 pd=42676 as=2.1498e+07 ps=57152 
M3250 Vdd n_973 n_973 GND dfet w=846 l=1974
+ ad=0 pd=0 as=4.418e+06 ps=12408 
M3251 n_436 dpc2_XSB sb4 GND efet w=1222 l=658
+ ad=0 pd=0 as=0 ps=0 
M3252 x4 dpc3_SBX sb4 GND efet w=1128 l=752
+ ad=0 pd=0 as=0 ps=0 
M3253 Vdd n_578 n_578 GND dfet w=846 l=1504
+ ad=0 pd=0 as=2.59778e+06 ps=7520 
M3254 GND notx5 n_578 GND efet w=5264 l=658
+ ad=0 pd=0 as=1.38814e+07 ps=33464 
M3255 Vdd notx5 notx5 GND dfet w=846 l=1974
+ ad=0 pd=0 as=8.52674e+06 ps=24064 
M3256 notx5 x5 GND GND efet w=3431 l=705
+ ad=4.60356e+06 pd=15792 as=0 ps=0 
M3257 x5 cclk n_578 GND efet w=1034 l=752
+ ad=2.3327e+06 pd=8648 as=0 ps=0 
M3258 n_3 dpc4_SSB sb4 GND efet w=1504 l=846
+ ad=0 pd=0 as=0 ps=0 
M3259 GND nots4 n_3 GND efet w=4136 l=564
+ ad=0 pd=0 as=0 ps=0 
M3260 n_973 s4 GND GND efet w=3196 l=564
+ ad=7.8287e+06 pd=21620 as=0 ps=0 
M3261 n_973 cclk nots4 GND efet w=1128 l=752
+ ad=0 pd=0 as=2.50059e+06 ps=9212 
M3262 n_3 dpc7_SS s4 GND efet w=1034 l=752
+ ad=0 pd=0 as=2.84519e+06 ps=6956 
M3263 s4 dpc6_SBS sb4 GND efet w=1128 l=752
+ ad=0 pd=0 as=0 ps=0 
M3264 sb4 cclk Vdd GND efet w=2162 l=658
+ ad=0 pd=0 as=0 ps=0 
M3265 Vdd n_280 n_280 GND dfet w=846 l=1504
+ ad=0 pd=0 as=3.17212e+06 ps=9588 
M3266 n_280 dpc5_SADL adl5 GND efet w=1410 l=564
+ ad=1.71507e+07 pd=42676 as=2.20105e+07 ps=58092 
M3267 Vdd n_496 n_496 GND dfet w=846 l=1880
+ ad=0 pd=0 as=4.13525e+06 ps=12032 
M3268 n_578 dpc2_XSB sb5 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M3269 x5 dpc3_SBX sb5 GND efet w=1034 l=752
+ ad=0 pd=0 as=0 ps=0 
M3270 GND noty6 n_518 GND efet w=5358 l=658
+ ad=0 pd=0 as=1.30243e+07 ps=33464 
M3271 Vdd noty6 noty6 GND dfet w=940 l=1880
+ ad=0 pd=0 as=8.45605e+06 ps=24064 
M3272 noty6 y6 GND GND efet w=3290 l=564
+ ad=4.78028e+06 pd=15792 as=0 ps=0 
M3273 y6 cclk n_518 GND efet w=1034 l=752
+ ad=2.29736e+06 pd=8648 as=0 ps=0 
M3274 n_1548 n_1548 Vdd GND dfet w=846 l=940
+ ad=2.12064e+06 pd=6956 as=0 ps=0 
M3275 n_518 dpc0_YSB sb6 GND efet w=1222 l=752
+ ad=0 pd=0 as=3.67136e+07 ps=92872 
M3276 y6 dpc1_SBY sb6 GND efet w=1034 l=658
+ ad=0 pd=0 as=0 ps=0 
M3277 nABL7 cclk n_171 GND efet w=1128 l=752
+ ad=2.59778e+06 pd=8836 as=0 ps=0 
M3278 n_577 ADL_ABL nABL7 GND efet w=1128 l=658
+ ad=742224 pd=3572 as=0 ps=0 
M3279 n_1046 cp1 n_577 GND efet w=1128 l=658
+ ad=9.1541e+06 pd=24440 as=0 ps=0 
M3280 abl7 nABL7 GND GND efet w=8930 l=611
+ ad=8.5179e+06 pd=24064 as=0 ps=0 
M3281 abl7 abl7 Vdd GND dfet w=846 l=1316
+ ad=2.44934e+07 pd=78584 as=0 ps=0 
M3282 Vdd n_1668 n_1668 GND dfet w=846 l=940
+ ad=0 pd=0 as=2.88937e+06 ps=9776 
M3283 GND adh0 n_1668 GND efet w=7238 l=658
+ ad=0 pd=0 as=9.92283e+06 ps=25380 
M3284 abh0 nABH0 GND GND efet w=6204 l=658
+ ad=4.55054e+06 pd=18424 as=0 ps=0 
M3285 GND adl7 n_1046 GND efet w=7614 l=564
+ ad=0 pd=0 as=0 ps=0 
M3286 Vdd n_1251 n_1251 GND dfet w=940 l=1504
+ ad=0 pd=0 as=2.59778e+06 ps=7520 
M3287 GND noty7 n_1251 GND efet w=5264 l=658
+ ad=0 pd=0 as=1.37577e+07 ps=32900 
M3288 Vdd noty7 noty7 GND dfet w=846 l=1880
+ ad=0 pd=0 as=8.45605e+06 ps=24064 
M3289 noty7 y7 GND GND efet w=3290 l=658
+ ad=4.69192e+06 pd=15792 as=0 ps=0 
M3290 y7 cclk n_1251 GND efet w=1034 l=752
+ ad=2.29736e+06 pd=8460 as=0 ps=0 
M3291 n_1046 n_1046 Vdd GND dfet w=940 l=1034
+ ad=2.09413e+06 pd=6768 as=0 ps=0 
M3292 n_1251 dpc0_YSB sb7 GND efet w=1316 l=752
+ ad=0 pd=0 as=3.60597e+07 ps=94000 
M3293 y7 dpc1_SBY sb7 GND efet w=1034 l=752
+ ad=0 pd=0 as=0 ps=0 
M3294 Vdd n_1724 n_1724 GND dfet w=940 l=1504
+ ad=0 pd=0 as=2.68614e+06 ps=7520 
M3295 GND notx6 n_1724 GND efet w=5264 l=658
+ ad=0 pd=0 as=1.38107e+07 ps=33088 
M3296 Vdd notx6 notx6 GND dfet w=846 l=1880
+ ad=0 pd=0 as=8.35002e+06 ps=24064 
M3297 n_280 dpc4_SSB sb5 GND efet w=1504 l=752
+ ad=0 pd=0 as=0 ps=0 
M3298 notx6 x6 GND GND efet w=3431 l=611
+ ad=5.06303e+06 pd=15980 as=0 ps=0 
M3299 x6 cclk n_1724 GND efet w=1128 l=752
+ ad=2.38572e+06 pd=8460 as=0 ps=0 
M3300 GND nots5 n_280 GND efet w=4136 l=564
+ ad=0 pd=0 as=0 ps=0 
M3301 n_496 s5 GND GND efet w=3102 l=564
+ ad=7.9524e+06 pd=21432 as=0 ps=0 
M3302 n_496 cclk nots5 GND efet w=1128 l=752
+ ad=0 pd=0 as=2.50059e+06 ps=9212 
M3303 n_280 dpc7_SS s5 GND efet w=1034 l=752
+ ad=0 pd=0 as=2.89821e+06 ps=7144 
M3304 s5 dpc6_SBS sb5 GND efet w=1128 l=658
+ ad=0 pd=0 as=0 ps=0 
M3305 sb5 cclk Vdd GND efet w=2162 l=658
+ ad=0 pd=0 as=0 ps=0 
M3306 Vdd n_618 n_618 GND dfet w=846 l=1598
+ ad=0 pd=0 as=3.16329e+06 ps=9400 
M3307 n_618 dpc5_SADL adl6 GND efet w=1410 l=470
+ ad=1.66559e+07 pd=42676 as=2.18779e+07 ps=57904 
M3308 Vdd n_1187 n_1187 GND dfet w=940 l=1880
+ ad=0 pd=0 as=4.03805e+06 ps=12220 
M3309 n_1724 dpc2_XSB sb6 GND efet w=1222 l=658
+ ad=0 pd=0 as=0 ps=0 
M3310 x6 dpc3_SBX sb6 GND efet w=1128 l=752
+ ad=0 pd=0 as=0 ps=0 
M3311 Vdd n_871 n_871 GND dfet w=940 l=1504
+ ad=0 pd=0 as=2.59778e+06 ps=7520 
M3312 GND notx7 n_871 GND efet w=5358 l=658
+ ad=0 pd=0 as=1.28034e+07 ps=33276 
M3313 Vdd notx7 notx7 GND dfet w=940 l=1880
+ ad=0 pd=0 as=8.45605e+06 ps=24064 
M3314 notx7 x7 GND GND efet w=3196 l=564
+ ad=4.75377e+06 pd=15792 as=0 ps=0 
M3315 x7 cclk n_871 GND efet w=1034 l=752
+ ad=2.3327e+06 pd=8460 as=0 ps=0 
M3316 n_871 dpc2_XSB sb7 GND efet w=1222 l=752
+ ad=0 pd=0 as=0 ps=0 
M3317 n_618 dpc4_SSB sb6 GND efet w=1598 l=846
+ ad=0 pd=0 as=0 ps=0 
M3318 GND nots6 n_618 GND efet w=4230 l=658
+ ad=0 pd=0 as=0 ps=0 
M3319 n_1187 s6 GND GND efet w=3149 l=611
+ ad=7.50176e+06 pd=21620 as=0 ps=0 
M3320 n_1187 cclk nots6 GND efet w=1034 l=752
+ ad=0 pd=0 as=2.41223e+06 ps=8836 
M3321 adl2 dpc10_ADLADD alub2 GND efet w=1175 l=799
+ ad=0 pd=0 as=5.23975e+06 ps=13912 
M3322 alub2 dpc8_nDBADD n_458 GND efet w=1128 l=658
+ ad=0 pd=0 as=8.52674e+06 ps=25944 
M3323 alub2 dpc9_DBADD idb2 GND efet w=1128 l=658
+ ad=0 pd=0 as=1.88295e+07 ps=52452 
M3324 GND idb2 n_458 GND efet w=5687 l=705
+ ad=0 pd=0 as=0 ps=0 
M3325 n_458 n_458 Vdd GND dfet w=846 l=1598
+ ad=2.93355e+06 pd=8084 as=0 ps=0 
M3326 n_A_B_1 alua1 GND GND efet w=2914 l=564
+ ad=0 pd=0 as=0 ps=0 
M3327 GND alub1 n_A_B_1 GND efet w=2914 l=658
+ ad=0 pd=0 as=0 ps=0 
M3328 Vdd n_A_B_1 n_A_B_1 GND dfet w=846 l=2162
+ ad=0 pd=0 as=1.23881e+07 ps=38728 
M3329 naluresult1 dpc15_ANDS nA_B1 GND efet w=1034 l=752
+ ad=0 pd=0 as=0 ps=0 
M3330 n_452 alua2 GND GND efet w=5734 l=658
+ ad=2.69498e+06 pd=12408 as=0 ps=0 
M3331 nA_B2 alub2 n_452 GND efet w=5734 l=658
+ ad=1.0073e+07 pd=28388 as=0 ps=0 
M3332 Vdd nA_B2 nA_B2 GND dfet w=987 l=2021
+ ad=0 pd=0 as=2.04112e+07 ps=66740 
M3333 GND nA_B0 n_1348 GND efet w=3196 l=658
+ ad=0 pd=0 as=0 ps=0 
M3334 C01 n_A_B_0 GND GND efet w=2632 l=564
+ ad=9.12759e+06 pd=24816 as=0 ps=0 
M3335 n_942 nA_B0 C01 GND efet w=5264 l=564
+ ad=4.23244e+06 pd=15228 as=0 ps=0 
M3336 GND notalucin n_942 GND efet w=6862 l=564
+ ad=0 pd=0 as=0 ps=0 
M3337 n_406 n_AxB_0 GND GND efet w=3290 l=658
+ ad=1.5463e+06 pd=7520 as=0 ps=0 
M3338 n_AxBxC_0 n_105 n_406 GND efet w=3290 l=658
+ ad=7.39573e+06 pd=20492 as=0 ps=0 
M3339 Vdd n_AxBxC_0 n_AxBxC_0 GND dfet w=846 l=1692
+ ad=0 pd=0 as=4.02922e+06 ps=9776 
M3340 GND n_134 n_467 GND efet w=2444 l=564
+ ad=0 pd=0 as=8.10261e+06 ps=19928 
M3341 GND n_236 n_1427 GND efet w=3666 l=564
+ ad=0 pd=0 as=0 ps=0 
M3342 GND n_470 n_467 GND efet w=2726 l=470
+ ad=0 pd=0 as=0 ps=0 
M3343 n_930 n_1276 GND GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M3344 n_180 n_180 Vdd GND dfet w=987 l=1175
+ ad=8.57976e+06 pd=27448 as=0 ps=0 
M3345 n_501 n_501 Vdd GND dfet w=846 l=1128
+ ad=1.57546e+07 pd=60160 as=0 ps=0 
M3346 n_501 n_180 GND GND efet w=3619 l=611
+ ad=0 pd=0 as=0 ps=0 
M3347 n_180 notRdy0 GND GND efet w=3854 l=658
+ ad=0 pd=0 as=0 ps=0 
M3348 GND op_T3_branch n_1708 GND efet w=3572 l=658
+ ad=0 pd=0 as=5.75224e+06 ps=17484 
M3349 n_1716 op_T3_branch GND GND efet w=2820 l=564
+ ad=1.52421e+07 pd=38352 as=0 ps=0 
M3350 GND n_510 n_1716 GND efet w=2914 l=564
+ ad=0 pd=0 as=0 ps=0 
M3351 n_510 n_347 GND GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M3352 GND op_rmw n_510 GND efet w=3149 l=705
+ ad=0 pd=0 as=0 ps=0 
M3353 Vdd op_rmw op_rmw GND dfet w=752 l=1222
+ ad=0 pd=0 as=5.66388e+06 ps=16732 
M3354 n_510 n_510 Vdd GND dfet w=940 l=1504
+ ad=7.07764e+06 pd=23312 as=0 ps=0 
M3355 op_rmw n_790 GND GND efet w=3478 l=658
+ ad=3.56974e+06 pd=11656 as=0 ps=0 
M3356 n_335 nop_store GND GND efet w=8272 l=564
+ ad=9.66658e+06 pd=30644 as=0 ps=0 
M3357 GND n_368 n_218 GND efet w=3572 l=658
+ ad=0 pd=0 as=7.23668e+06 ps=21808 
M3358 n_368 n_368 Vdd GND dfet w=1034 l=1504
+ ad=7.18367e+06 pd=22936 as=0 ps=0 
M3359 n_790 n_790 Vdd GND dfet w=846 l=1504
+ ad=2.58895e+07 pd=90616 as=0 ps=0 
M3360 Vdd n_218 n_218 GND dfet w=940 l=940
+ ad=0 pd=0 as=6.58282e+06 ps=24628 
M3361 GND n_347 n_335 GND efet w=8178 l=658
+ ad=0 pd=0 as=0 ps=0 
M3362 n_1708 n_1708 Vdd GND dfet w=940 l=1222
+ ad=4.18738e+07 pd=153220 as=0 ps=0 
M3363 n_1716 n_1716 Vdd GND dfet w=940 l=1222
+ ad=2.00135e+07 pd=71252 as=0 ps=0 
M3364 Vdd n_944 n_944 GND dfet w=940 l=1128
+ ad=0 pd=0 as=2.88937e+06 ps=8836 
M3365 GND n_1449 n_944 GND efet w=4700 l=658
+ ad=0 pd=0 as=1.25118e+07 ps=33652 
M3366 GND n_1708 n_236 GND efet w=6157 l=611
+ ad=0 pd=0 as=6.33541e+06 ps=16356 
M3367 n_944 cclk pipeUNK37 GND efet w=1316 l=658
+ ad=0 pd=0 as=1.37842e+06 ps=7144 
M3368 GND pipeUNK37 n_198 GND efet w=8789 l=611
+ ad=0 pd=0 as=9.21595e+06 ps=25756 
M3369 n_198 pipeUNK37 GND GND efet w=1128 l=752
+ ad=0 pd=0 as=0 ps=0 
M3370 GND n_759 n_944 GND efet w=7379 l=611
+ ad=0 pd=0 as=0 ps=0 
M3371 n_236 n_236 Vdd GND dfet w=846 l=752
+ ad=6.69592e+07 pd=235000 as=0 ps=0 
M3372 n_501 n_819 GND GND efet w=3995 l=611
+ ad=0 pd=0 as=0 ps=0 
M3373 GND op_T2_abs_access n_773 GND efet w=3008 l=564
+ ad=0 pd=0 as=6.85674e+06 ps=19552 
M3374 n_1272 cp1 notRdy0 GND efet w=1034 l=752
+ ad=3.40186e+06 pd=13160 as=0 ps=0 
M3375 n_773 n_646 GND GND efet w=4183 l=705
+ ad=0 pd=0 as=0 ps=0 
M3376 n_773 n_773 Vdd GND dfet w=846 l=1222
+ ad=9.99352e+06 pd=32148 as=0 ps=0 
M3377 Vdd n_275 n_275 GND dfet w=846 l=1034
+ ad=0 pd=0 as=6.73303e+06 ps=19928 
M3378 n_275 n_1697 GND GND efet w=4747 l=893
+ ad=6.57398e+06 pd=19176 as=0 ps=0 
M3379 notRdy0 cp1 n_1276 GND efet w=1128 l=752
+ ad=0 pd=0 as=2.3327e+06 ps=6204 
M3380 GND n_630 n_1705 GND efet w=2632 l=658
+ ad=0 pd=0 as=0 ps=0 
M3381 n_930 n_1276 GND GND efet w=1598 l=658
+ ad=0 pd=0 as=0 ps=0 
M3382 Vdd n_1655 n_1655 GND dfet w=846 l=940
+ ad=0 pd=0 as=7.2897e+06 ps=24816 
M3383 n_1655 n_1211 GND GND efet w=3478 l=564
+ ad=2.92472e+06 pd=9776 as=0 ps=0 
M3384 GND n_236 n_176 GND efet w=3901 l=611
+ ad=0 pd=0 as=8.72113e+06 ps=28200 
M3385 n_176 n_10 GND GND efet w=4136 l=564
+ ad=0 pd=0 as=0 ps=0 
M3386 GND n_646 n_272 GND efet w=2914 l=564
+ ad=0 pd=0 as=0 ps=0 
M3387 n_1278 n_824 n_1642 GND efet w=7896 l=564
+ ad=4.17059e+06 pd=16732 as=6.71536e+06 ps=19176 
M3388 GND n_462 n_1278 GND efet w=7802 l=658
+ ad=0 pd=0 as=0 ps=0 
M3389 n_1642 n_1642 Vdd GND dfet w=940 l=940
+ ad=3.91612e+07 pd=151340 as=0 ps=0 
M3390 n_182 n_1655 GND GND efet w=2538 l=564
+ ad=0 pd=0 as=0 ps=0 
M3391 n_176 n_176 Vdd GND dfet w=940 l=1034
+ ad=2.33094e+07 pd=88736 as=0 ps=0 
M3392 Vdd n_952 n_952 GND dfet w=940 l=846
+ ad=0 pd=0 as=3.35415e+07 ps=124268 
M3393 n_952 n_272 GND GND efet w=5264 l=658
+ ad=7.17483e+06 pd=23876 as=0 ps=0 
M3394 n_182 n_646 GND GND efet w=4136 l=564
+ ad=0 pd=0 as=0 ps=0 
M3395 GND n_930 n_1286 GND efet w=6204 l=564
+ ad=0 pd=0 as=9.2778e+06 ps=22372 
M3396 GND n_773 n_275 GND efet w=4089 l=611
+ ad=0 pd=0 as=0 ps=0 
M3397 GND n_1272 n_608 GND efet w=4935 l=705
+ ad=0 pd=0 as=6.15869e+06 ps=20116 
M3398 Vdd n_608 n_608 GND dfet w=846 l=1598
+ ad=0 pd=0 as=3.1898e+06 ps=8460 
M3399 n_559 cclk n_608 GND efet w=1128 l=846
+ ad=1.8909e+06 pd=8648 as=0 ps=0 
M3400 Vdd n_916 n_916 GND dfet w=846 l=846
+ ad=0 pd=0 as=2.19928e+07 ps=78772 
M3401 GND n_275 n_104 GND efet w=3666 l=752
+ ad=0 pd=0 as=0 ps=0 
M3402 n_916 n_1517 GND GND efet w=5922 l=564
+ ad=1.39167e+07 pd=35532 as=0 ps=0 
M3403 n_387 n_206 n_916 GND efet w=11327 l=611
+ ad=5.76991e+06 pd=23688 as=0 ps=0 
M3404 GND n_853 n_387 GND efet w=11327 l=611
+ ad=0 pd=0 as=0 ps=0 
M3405 notRdy0 n_198 GND GND efet w=12784 l=658
+ ad=0 pd=0 as=0 ps=0 
M3406 nWR op_T4_brk GND GND efet w=3290 l=564
+ ad=2.76213e+07 pd=68620 as=0 ps=0 
M3407 GND op_T2_php_pha nWR GND efet w=3290 l=658
+ ad=0 pd=0 as=0 ps=0 
M3408 n_191 n_790 GND GND efet w=3666 l=658
+ ad=9.52521e+06 pd=29328 as=0 ps=0 
M3409 n_1065 n_1065 Vdd GND dfet w=940 l=1504
+ ad=7.62547e+06 pd=24252 as=0 ps=0 
M3410 n_591 n_1258 GND GND efet w=7896 l=658
+ ad=4.47985e+06 pd=18424 as=0 ps=0 
M3411 nop_set_C op_asl_rol n_591 GND efet w=6392 l=564
+ ad=2.68438e+07 pd=68808 as=0 ps=0 
M3412 GND op_T3_mem_zp_idx n_347 GND efet w=3478 l=658
+ ad=0 pd=0 as=1.49593e+07 ps=42488 
M3413 nop_set_C x_op_T__adc_sbc GND GND efet w=2820 l=564
+ ad=0 pd=0 as=0 ps=0 
M3414 n_327 op_T0_plp GND GND efet w=2914 l=658
+ ad=8.34118e+06 pd=24252 as=0 ps=0 
M3415 GND x_op_T4_rti n_327 GND efet w=3572 l=658
+ ad=0 pd=0 as=0 ps=0 
M3416 nop_set_C op_T__cmp GND GND efet w=2444 l=564
+ ad=0 pd=0 as=0 ps=0 
M3417 GND op_T__cpx_cpy_abs nop_set_C GND efet w=2350 l=564
+ ad=0 pd=0 as=0 ps=0 
M3418 nop_set_C op_T__asl_rol_a GND GND efet w=3243 l=611
+ ad=0 pd=0 as=0 ps=0 
M3419 nop_set_C nop_set_C Vdd GND dfet w=940 l=1598
+ ad=8.37653e+06 pd=26132 as=0 ps=0 
M3420 GND op_T__cpx_cpy_imm_zp nop_set_C GND efet w=3525 l=611
+ ad=0 pd=0 as=0 ps=0 
M3421 n_327 n_327 Vdd GND dfet w=1034 l=1692
+ ad=7.90822e+06 pd=25004 as=0 ps=0 
M3422 GND op_T0_cld_sed n_774 GND efet w=2632 l=658
+ ad=0 pd=0 as=1.09655e+07 ps=29516 
M3423 n_347 op_T3_mem_abs GND GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M3424 GND op_T2_mem_zp n_347 GND efet w=3102 l=564
+ ad=0 pd=0 as=0 ps=0 
M3425 n_347 op_T5_mem_ind_idx GND GND efet w=3807 l=611
+ ad=0 pd=0 as=0 ps=0 
M3426 GND op_T4_mem_abs_idx n_347 GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M3427 Vdd n_1137 n_1137 GND dfet w=846 l=1222
+ ad=0 pd=0 as=6.74187e+06 ps=20304 
M3428 Vdd nWR nWR GND dfet w=846 l=1034
+ ad=0 pd=0 as=2.32387e+06 ps=6768 
M3429 GND n_218 n_1716 GND efet w=3431 l=517
+ ad=0 pd=0 as=0 ps=0 
M3430 GND n_347 n_191 GND efet w=3008 l=564
+ ad=0 pd=0 as=0 ps=0 
M3431 Vdd n_1258 n_1258 GND dfet w=940 l=564
+ ad=0 pd=0 as=3.88784e+07 ps=134420 
M3432 n_1391 n_1391 Vdd GND dfet w=1034 l=1410
+ ad=6.03676e+07 pd=233120 as=0 ps=0 
M3433 n_816 n_790 n_1137 GND efet w=4324 l=658
+ ad=3.81715e+06 pd=14852 as=6.4061e+06 ps=16732 
M3434 GND nop_store n_816 GND efet w=5311 l=611
+ ad=0 pd=0 as=0 ps=0 
M3435 n_198 n_198 Vdd GND dfet w=940 l=1034
+ ad=1.63819e+07 pd=52452 as=0 ps=0 
M3436 notRnWprepad cp1 n_759 GND efet w=1034 l=846
+ ad=0 pd=0 as=1.35191e+06 ps=7144 
M3437 Vdd n_424 notRdy0 GND dfet w=1692 l=564
+ ad=0 pd=0 as=0 ps=0 
M3438 notRnWprepad notRnWprepad Vdd GND dfet w=846 l=846
+ ad=6.03145e+07 pd=212252 as=0 ps=0 
M3439 GND n_1258 nWR GND efet w=3478 l=564
+ ad=0 pd=0 as=0 ps=0 
M3440 nWR n_335 GND GND efet w=6063 l=517
+ ad=0 pd=0 as=0 ps=0 
M3441 GND n_440 nWR GND efet w=5076 l=564
+ ad=0 pd=0 as=0 ps=0 
M3442 GND n_1642 nWR GND efet w=3431 l=611
+ ad=0 pd=0 as=0 ps=0 
M3443 GND n_1258 n_1716 GND efet w=3572 l=564
+ ad=0 pd=0 as=0 ps=0 
M3444 n_191 n_191 Vdd GND dfet w=1034 l=1034
+ ad=5.24858e+06 pd=20868 as=0 ps=0 
M3445 GND notRdy0 n_191 GND efet w=2632 l=564
+ ad=0 pd=0 as=0 ps=0 
M3446 Vdd n_1120 n_1120 GND dfet w=940 l=1034
+ ad=0 pd=0 as=5.53134e+06 ps=20304 
M3447 n_1258 n_390 GND GND efet w=6815 l=611
+ ad=6.9716e+06 pd=19176 as=0 ps=0 
M3448 n_889 op_T0_clc_sec GND GND efet w=2538 l=658
+ ad=7.81986e+06 pd=26132 as=0 ps=0 
M3449 n_347 n_347 Vdd GND dfet w=846 l=1504
+ ad=3.79595e+07 pd=131224 as=0 ps=0 
M3450 GND n_1533 clock2 GND efet w=12220 l=564
+ ad=0 pd=0 as=1.85998e+07 ps=43240 
M3451 Vdd clock2 clock2 GND dfet w=846 l=564
+ ad=0 pd=0 as=1.7983e+08 ps=575844 
M3452 n_664 n_664 Vdd GND dfet w=940 l=1504
+ ad=6.42377e+06 pd=18988 as=0 ps=0 
M3453 GND op_implied n_664 GND efet w=3807 l=611
+ ad=0 pd=0 as=5.28393e+06 ps=15416 
M3454 GND pd6_clearIR n_1309 GND efet w=6768 l=658
+ ad=0 pd=0 as=0 ps=0 
M3455 n_1309 n_1309 Vdd GND dfet w=1034 l=658
+ ad=6.29123e+06 pd=24440 as=0 ps=0 
M3456 GND notRdy0 n_1180 GND efet w=4042 l=658
+ ad=0 pd=0 as=9.77262e+06 ps=24628 
M3457 n_1533 cp1 n_1180 GND efet w=1504 l=752
+ ad=1.4491e+06 pd=8084 as=0 ps=0 
M3458 n_1180 pipenT0 GND GND efet w=4371 l=611
+ ad=0 pd=0 as=0 ps=0 
M3459 n_390 n_653 GND GND efet w=4559 l=611
+ ad=4.74493e+06 pd=12220 as=0 ps=0 
M3460 Vdd n_390 n_390 GND dfet w=846 l=1974
+ ad=0 pd=0 as=1.37223e+07 ps=41736 
M3461 n_889 n_889 Vdd GND dfet w=1128 l=1880
+ ad=4.13525e+06 pd=11844 as=0 ps=0 
M3462 Vdd n_1180 n_1180 GND dfet w=846 l=1598
+ ad=0 pd=0 as=3.84366e+06 ps=9588 
M3463 n_653 cp1 n_1497 GND efet w=1222 l=752
+ ad=1.48445e+06 pd=6768 as=8.09378e+06 ps=25568 
M3464 GND n_1533 n_964 GND efet w=5170 l=658
+ ad=0 pd=0 as=8.60626e+06 ps=20868 
M3465 n_1497 pipeUNK41 GND GND efet w=4841 l=611
+ ad=0 pd=0 as=0 ps=0 
M3466 n_191 cclk pipeUNK40 GND efet w=1222 l=846
+ ad=0 pd=0 as=1.35191e+06 ps=6016 
M3467 nWR cclk pipenWR_phi2 GND efet w=1128 l=752
+ ad=0 pd=0 as=2.48292e+06 ps=8648 
M3468 GND C1x5Reset notRnWprepad GND efet w=6627 l=611
+ ad=0 pd=0 as=0 ps=0 
M3469 Vdd n_424 n_424 GND dfet w=940 l=658
+ ad=0 pd=0 as=5.99964e+06 ps=23688 
M3470 n_424 n_198 GND GND efet w=5687 l=611
+ ad=8.44722e+06 pd=21432 as=0 ps=0 
M3471 GND Reset0 n_14 GND efet w=1880 l=658
+ ad=0 pd=0 as=1.58695e+07 ps=40608 
M3472 GND n_666 n_862 GND efet w=14194 l=564
+ ad=0 pd=0 as=0 ps=0 
M3473 notRnWprepad notRdy0 GND GND efet w=5170 l=564
+ ad=0 pd=0 as=0 ps=0 
M3474 n_14 n_14 Vdd GND dfet w=940 l=1786
+ ad=1.74423e+07 pd=65236 as=0 ps=0 
M3475 n_862 n_862 Vdd GND dfet w=846 l=752
+ ad=1.30578e+08 pd=463608 as=0 ps=0 
M3476 n_109 n_1380 GND GND efet w=8601 l=611
+ ad=1.01614e+07 pd=32712 as=0 ps=0 
M3477 notRnWprepad pipenWR_phi2 GND GND efet w=8178 l=564
+ ad=0 pd=0 as=0 ps=0 
M3478 n_104 op_T4_jmp GND GND efet w=3948 l=564
+ ad=0 pd=0 as=0 ps=0 
M3479 n_964 pipenT0 GND GND efet w=4324 l=564
+ ad=0 pd=0 as=0 ps=0 
M3480 GND n_664 n_1697 GND efet w=3008 l=658
+ ad=0 pd=0 as=6.89208e+06 ps=19176 
M3481 Vdd n_409 n_409 GND dfet w=1128 l=564
+ ad=0 pd=0 as=1.60904e+07 ps=56212 
M3482 Vdd n_1497 n_1497 GND dfet w=940 l=1504
+ ad=0 pd=0 as=5.54017e+06 ps=15980 
M3483 n_889 cclk pipeUNK42 GND efet w=1128 l=752
+ ad=0 pd=0 as=2.45641e+06 ps=6392 
M3484 pipenT0 cclk n_17 GND efet w=1128 l=752
+ ad=4.00271e+06 pd=12220 as=8.70346e+06 ps=18800 
M3485 pipeUNK41 cclk n_504 GND efet w=1128 l=752
+ ad=2.03228e+06 pd=7708 as=1.10362e+07 ps=29140 
M3486 Vdd n_964 n_964 GND dfet w=940 l=1504
+ ad=0 pd=0 as=1.31921e+07 ps=41736 
M3487 n_1697 n_1697 Vdd GND dfet w=940 l=1034
+ ad=1.29359e+07 pd=41360 as=0 ps=0 
M3488 nTWOCYCLE PD_xxx010x1 GND GND efet w=4559 l=611
+ ad=1.83259e+07 pd=50008 as=0 ps=0 
M3489 Vdd n_1641 n_1641 GND dfet w=1128 l=658
+ ad=0 pd=0 as=1.35279e+07 ps=48128 
M3490 GND pd0_clearIR n_409 GND efet w=7191 l=611
+ ad=0 pd=0 as=0 ps=0 
M3491 n_1641 pd1_clearIR GND GND efet w=7050 l=564
+ ad=0 pd=0 as=0 ps=0 
M3492 Vdd n_1605 n_1605 GND dfet w=1128 l=564
+ ad=0 pd=0 as=1.93685e+07 ps=69184 
M3493 Vdd n_227 n_227 GND dfet w=1128 l=564
+ ad=0 pd=0 as=8.62394e+06 ps=30644 
M3494 GND pd7_clearIR n_1605 GND efet w=6956 l=564
+ ad=0 pd=0 as=0 ps=0 
M3495 n_227 pd4_clearIR GND GND efet w=6815 l=611
+ ad=0 pd=0 as=0 ps=0 
M3496 clock1 n_964 GND GND efet w=7943 l=611
+ ad=1.22555e+07 pd=21056 as=0 ps=0 
M3497 GND n_964 n_17 GND efet w=3478 l=658
+ ad=0 pd=0 as=0 ps=0 
M3498 GND n_440 n_812 GND efet w=5828 l=658
+ ad=0 pd=0 as=6.8479e+06 ps=20868 
M3499 n_104 n_440 GND GND efet w=3807 l=611
+ ad=0 pd=0 as=0 ps=0 
M3500 n_812 n_646 GND GND efet w=5781 l=611
+ ad=0 pd=0 as=0 ps=0 
M3501 Vdd n_109 n_109 GND dfet w=846 l=564
+ ad=0 pd=0 as=2.81427e+07 ps=102648 
M3502 n_770 n_559 GND GND efet w=5076 l=658
+ ad=4.67424e+06 pd=15980 as=0 ps=0 
M3503 n_666 cp1 n_1380 GND efet w=1128 l=752
+ ad=1.29889e+06 pd=6392 as=1.06209e+07 ps=30080 
M3504 GND notRdy0 n_1718 GND efet w=3760 l=564
+ ad=0 pd=0 as=6.00848e+06 ps=18424 
M3505 GND notRdy0 n_1120 GND efet w=3290 l=564
+ ad=0 pd=0 as=6.42377e+06 ps=19176 
M3506 n_137 n_1120 GND GND efet w=3196 l=564
+ ad=1.80254e+06 pd=7520 as=0 ps=0 
M3507 n_504 n_440 n_137 GND efet w=3196 l=564
+ ad=0 pd=0 as=0 ps=0 
M3508 Vdd n_504 n_504 GND dfet w=940 l=1410
+ ad=0 pd=0 as=3.76414e+06 ps=10904 
M3509 n_17 n_17 Vdd GND dfet w=846 l=846
+ ad=1.41818e+07 pd=49256 as=0 ps=0 
M3510 n_1065 cclk n_1124 GND efet w=1410 l=752
+ ad=0 pd=0 as=2.51826e+06 ps=6392 
M3511 n_1039 pipeUNK40 GND GND efet w=5640 l=658
+ ad=1.00024e+07 pd=28952 as=0 ps=0 
M3512 n_2 notRdy0 n_1039 GND efet w=4982 l=564
+ ad=7.1925e+06 pd=22748 as=0 ps=0 
M3513 GND pipeUNK39 n_2 GND efet w=7990 l=658
+ ad=0 pd=0 as=0 ps=0 
M3514 n_17 n_732 GND GND efet w=3478 l=658
+ ad=0 pd=0 as=0 ps=0 
M3515 clock1 n_732 GND GND efet w=7050 l=658
+ ad=0 pd=0 as=0 ps=0 
M3516 Vdd n_17 clock1 GND dfet w=1034 l=658
+ ad=0 pd=0 as=0 ps=0 
M3517 GND PD_1xx000x0 nTWOCYCLE GND efet w=4230 l=564
+ ad=0 pd=0 as=0 ps=0 
M3518 PD_xxx010x1 PD_xxx010x1 Vdd GND dfet w=940 l=940
+ ad=9.03923e+06 pd=32712 as=0 ps=0 
M3519 n_928 n_928 Vdd GND dfet w=1128 l=564
+ ad=7.68732e+06 pd=27636 as=0 ps=0 
M3520 Vdd n_1083 n_1083 GND dfet w=1128 l=658
+ ad=0 pd=0 as=1.51449e+07 ps=57152 
M3521 Vdd n_571 n_571 GND dfet w=1222 l=564
+ ad=0 pd=0 as=8.7123e+06 ps=33652 
M3522 GND pd3_clearIR n_1083 GND efet w=7050 l=658
+ ad=0 pd=0 as=0 ps=0 
M3523 n_571 pd2_clearIR GND GND efet w=6815 l=611
+ ad=0 pd=0 as=0 ps=0 
M3524 GND pd5_clearIR n_928 GND efet w=8366 l=658
+ ad=0 pd=0 as=0 ps=0 
M3525 nTWOCYCLE PD_xxxx10x0 n_1515 GND efet w=9541 l=517
+ ad=0 pd=0 as=6.67118e+06 ps=20304 
M3526 Vdd nTWOCYCLE nTWOCYCLE GND dfet w=846 l=940
+ ad=0 pd=0 as=8.24399e+06 ps=28576 
M3527 n_646 n_17 GND GND efet w=6157 l=611
+ ad=8.82716e+06 pd=19928 as=0 ps=0 
M3528 nTWOCYCLE cp1 nTWOCYCLE_phi1 GND efet w=1316 l=658
+ ad=0 pd=0 as=1.47561e+06 ps=7896 
M3529 n_440 cclk pipeUNK39 GND efet w=1128 l=752
+ ad=1.12217e+07 pd=35908 as=1.61699e+06 ps=7144 
M3530 n_253 pipeUNK42 GND GND efet w=4230 l=658
+ ad=7.14832e+06 pd=18612 as=0 ps=0 
M3531 n_1718 n_1718 Vdd GND dfet w=846 l=1598
+ ad=1.01261e+07 pd=34968 as=0 ps=0 
M3532 n_770 n_770 Vdd GND dfet w=846 l=1598
+ ad=1.47384e+07 pd=50760 as=0 ps=0 
M3533 Vdd n_586 n_586 GND dfet w=752 l=940
+ ad=0 pd=0 as=1.17342e+07 ps=43804 
M3534 n_1330 BRtaken n_586 GND efet w=4606 l=658
+ ad=5.78758e+06 pd=16732 as=1.89179e+07 ps=63732 
M3535 n_1286 n_470 GND GND efet w=3760 l=658
+ ad=0 pd=0 as=0 ps=0 
M3536 n_470 n_646 GND GND efet w=4888 l=658
+ ad=5.3016e+06 pd=17484 as=0 ps=0 
M3537 n_1286 n_1286 Vdd GND dfet w=940 l=940
+ ad=1.94922e+07 pd=68996 as=0 ps=0 
M3538 n_1448 n_1427 GND GND efet w=3290 l=658
+ ad=3.9762e+06 pd=13724 as=0 ps=0 
M3539 n_1330 BRtaken n_586 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M3540 GND nnT2BR n_1330 GND efet w=6768 l=564
+ ad=0 pd=0 as=0 ps=0 
M3541 n_853 n_770 GND GND efet w=2068 l=658
+ ad=2.6508e+06 pd=9212 as=0 ps=0 
M3542 n_1409 cp1 n_916 GND efet w=1128 l=752
+ ad=2.16482e+06 pd=8460 as=0 ps=0 
M3543 n_853 n_853 Vdd GND dfet w=940 l=1504
+ ad=1.97838e+07 pd=62792 as=0 ps=0 
M3544 n_1380 n_1154 GND GND efet w=6110 l=658
+ ad=0 pd=0 as=0 ps=0 
M3545 GND n_819 n_1380 GND efet w=4888 l=658
+ ad=0 pd=0 as=0 ps=0 
M3546 n_781 notRdy0 GND GND efet w=1410 l=658
+ ad=1.41199e+07 pd=39292 as=0 ps=0 
M3547 n_781 notRdy0 GND GND efet w=1598 l=658
+ ad=0 pd=0 as=0 ps=0 
M3548 n_1055 n_1708 GND GND efet w=3995 l=611
+ ad=9.18944e+06 pd=31396 as=0 ps=0 
M3549 n_1380 n_1380 Vdd GND dfet w=940 l=658
+ ad=9.42801e+06 pd=33276 as=0 ps=0 
M3550 n_1154 notRdy0 GND GND efet w=5734 l=564
+ ad=9.90516e+06 pd=32336 as=0 ps=0 
M3551 n_1517 n_572 GND GND efet w=3478 l=564
+ ad=9.58706e+06 pd=27448 as=0 ps=0 
M3552 Vdd n_1517 n_1517 GND dfet w=940 l=846
+ ad=0 pd=0 as=9.12759e+06 ps=31584 
M3553 Vdd n_1231 n_1231 GND dfet w=846 l=1880
+ ad=0 pd=0 as=3.95853e+06 ps=10340 
M3554 n_470 n_470 Vdd GND dfet w=940 l=940
+ ad=1.44999e+07 pd=53956 as=0 ps=0 
M3555 n_1448 n_1448 Vdd GND dfet w=940 l=1128
+ ad=8.9332e+06 pd=30268 as=0 ps=0 
M3556 Vdd n_572 n_572 GND dfet w=940 l=1222
+ ad=0 pd=0 as=2.05437e+07 ps=70688 
M3557 n_586 n_1619 GND GND efet w=4089 l=611
+ ad=0 pd=0 as=0 ps=0 
M3558 Vdd n_442 n_442 GND dfet w=893 l=1269
+ ad=0 pd=0 as=1.47119e+07 ps=53580 
M3559 GND n_182 n_442 GND efet w=4747 l=611
+ ad=0 pd=0 as=9.375e+06 ps=31396 
M3560 n_1347 cclk n_1527 GND efet w=1128 l=846
+ ad=0 pd=0 as=1.33424e+06 ps=5640 
M3561 n_1455 cclk n_1505 GND efet w=1222 l=846
+ ad=0 pd=0 as=1.34307e+06 ps=6956 
M3562 GND pipeUNK21 n_572 GND efet w=7238 l=564
+ ad=0 pd=0 as=8.13796e+06 ps=20680 
M3563 n_1231 n_1409 GND GND efet w=3384 l=658
+ ad=7.71383e+06 pd=23312 as=0 ps=0 
M3564 Vdd n_19 n_19 GND dfet w=940 l=1504
+ ad=0 pd=0 as=3.1898e+06 ps=9212 
M3565 Vdd n_1154 n_1154 GND dfet w=752 l=658
+ ad=0 pd=0 as=6.2824e+06 ps=22184 
M3566 n_1718 cp1 n_671 GND efet w=1128 l=752
+ ad=0 pd=0 as=1.2017e+06 ps=6768 
M3567 n_812 n_812 Vdd GND dfet w=940 l=940
+ ad=6.67118e+06 pd=22936 as=0 ps=0 
M3568 n_104 n_104 Vdd GND dfet w=940 l=1034
+ ad=4.25188e+07 pd=153032 as=0 ps=0 
M3569 n_1044 n_812 GND GND efet w=4042 l=564
+ ad=1.39874e+07 pd=39480 as=0 ps=0 
M3570 Vdd n_1044 n_1044 GND dfet w=940 l=1128
+ ad=0 pd=0 as=2.42106e+07 ps=93812 
M3571 n_1039 n_1039 Vdd GND dfet w=846 l=1974
+ ad=4.00271e+06 pd=9400 as=0 ps=0 
M3572 n_1161 cp1 n_109 GND efet w=1316 l=846
+ ad=2.59778e+06 pd=8648 as=0 ps=0 
M3573 Vdd n_253 n_253 GND dfet w=940 l=1786
+ ad=0 pd=0 as=3.70847e+07 ps=128968 
M3574 GND x_op_T0_bit n_1379 GND efet w=2867 l=611
+ ad=0 pd=0 as=1.27503e+07 ps=31960 
M3575 Vdd n_646 n_646 GND dfet w=940 l=658
+ ad=0 pd=0 as=1.06209e+08 ps=395176 
M3576 GND n_1161 n_732 GND efet w=7379 l=611
+ ad=0 pd=0 as=1.61876e+07 ps=43052 
M3577 Vdd n_732 n_732 GND dfet w=1034 l=940
+ ad=0 pd=0 as=1.06562e+07 ps=34216 
M3578 PD_xxxx10x0 PD_xxxx10x0 Vdd GND dfet w=940 l=846
+ ad=1.88914e+07 pd=71440 as=0 ps=0 
M3579 n_1515 PD_n_0xx0xx0x GND GND efet w=9400 l=564
+ ad=0 pd=0 as=0 ps=0 
M3580 GND n_409 PD_xxx010x1 GND efet w=3008 l=658
+ ad=0 pd=0 as=1.46501e+07 ps=39856 
M3581 PD_xxxx10x0 pd0_clearIR GND GND efet w=3572 l=564
+ ad=1.58341e+07 pd=40796 as=0 ps=0 
M3582 GND PD_0xx0xx0x PD_n_0xx0xx0x GND efet w=6110 l=658
+ ad=0 pd=0 as=8.62394e+06 ps=24440 
M3583 PD_0xx0xx0x PD_0xx0xx0x Vdd GND dfet w=846 l=1034
+ ad=9.76378e+06 pd=33276 as=0 ps=0 
M3584 PD_n_0xx0xx0x PD_n_0xx0xx0x Vdd GND dfet w=846 l=658
+ ad=1.0073e+07 pd=37412 as=0 ps=0 
M3585 PD_1xx000x0 PD_1xx000x0 Vdd GND dfet w=940 l=940
+ ad=1.58164e+07 pd=60724 as=0 ps=0 
M3586 GND pd1_clearIR PD_0xx0xx0x GND efet w=2914 l=564
+ ad=0 pd=0 as=1.41818e+07 ps=38352 
M3587 PD_xxx010x1 pd4_clearIR GND GND efet w=4559 l=611
+ ad=0 pd=0 as=0 ps=0 
M3588 GND n_1083 PD_xxx010x1 GND efet w=4324 l=564
+ ad=0 pd=0 as=0 ps=0 
M3589 PD_1xx000x0 pd0_clearIR GND GND efet w=2914 l=564
+ ad=1.7725e+07 pd=47376 as=0 ps=0 
M3590 GND PD_xxxx10x0 n_231 GND efet w=8178 l=564
+ ad=0 pd=0 as=1.24853e+07 ps=31208 
M3591 Vdd n_231 n_231 GND dfet w=846 l=658
+ ad=0 pd=0 as=9.36616e+06 ps=35344 
M3592 n_106 nTWOCYCLE_phi1 n_732 GND efet w=14147 l=611
+ ad=8.89785e+06 pd=29516 as=0 ps=0 
M3593 n_1528 cp1 n_1215 GND efet w=1316 l=846
+ ad=1.82905e+06 pd=7708 as=0 ps=0 
M3594 n_106 n_1528 GND GND efet w=14147 l=611
+ ad=0 pd=0 as=0 ps=0 
M3595 GND pd7_clearIR PD_0xx0xx0x GND efet w=4277 l=611
+ ad=0 pd=0 as=0 ps=0 
M3596 PD_1xx000x0 n_1605 GND GND efet w=3102 l=564
+ ad=0 pd=0 as=0 ps=0 
M3597 ONEBYTE n_231 GND GND efet w=7003 l=611
+ ad=6.91859e+06 pd=23876 as=0 ps=0 
M3598 GND D1x1 n_380 GND efet w=5264 l=564
+ ad=0 pd=0 as=2.9689e+06 ps=11656 
M3599 n_1039 cp1 n_24 GND efet w=1222 l=752
+ ad=0 pd=0 as=1.74953e+06 ps=7332 
M3600 n_440 n_24 GND GND efet w=14006 l=658
+ ad=0 pd=0 as=0 ps=0 
M3601 Vdd n_440 n_440 GND dfet w=1034 l=846
+ ad=0 pd=0 as=6.32923e+07 ps=227104 
M3602 GND n_31 n_1044 GND efet w=3995 l=705
+ ad=0 pd=0 as=0 ps=0 
M3603 p2 cp1 n_845 GND efet w=1128 l=752
+ ad=1.36958e+06 pd=5452 as=1.46943e+07 ps=45120 
M3604 GND p2 n_334 GND efet w=7238 l=752
+ ad=0 pd=0 as=0 ps=0 
M3605 Vdd n_334 n_334 GND dfet w=846 l=846
+ ad=0 pd=0 as=3.98592e+07 ps=145136 
M3606 Vdd n_845 n_845 GND dfet w=940 l=1786
+ ad=0 pd=0 as=7.54594e+06 ps=25380 
M3607 Vdd n_553 n_553 GND dfet w=940 l=1504
+ ad=0 pd=0 as=7.56362e+06 ps=24628 
M3608 ONEBYTE ONEBYTE Vdd GND dfet w=940 l=658
+ ad=6.08712e+07 pd=222216 as=0 ps=0 
M3609 n_380 fetch clearIR GND efet w=5264 l=658
+ ad=0 pd=0 as=6.87441e+06 ps=17860 
M3610 Vdd clearIR clearIR GND dfet w=940 l=1128
+ ad=0 pd=0 as=3.18715e+07 ps=104152 
M3611 PD_0xx0xx0x pd4_clearIR GND GND efet w=2914 l=564
+ ad=0 pd=0 as=0 ps=0 
M3612 GND n_1083 PD_xxxx10x0 GND efet w=3760 l=564
+ ad=0 pd=0 as=0 ps=0 
M3613 GND pd2_clearIR PD_xxx010x1 GND efet w=3008 l=564
+ ad=0 pd=0 as=0 ps=0 
M3614 GND pd2_clearIR PD_xxxx10x0 GND efet w=3666 l=564
+ ad=0 pd=0 as=0 ps=0 
M3615 PD_1xx000x0 pd3_clearIR GND GND efet w=3854 l=658
+ ad=0 pd=0 as=0 ps=0 
M3616 PD_1xx000x0 pd4_clearIR GND GND efet w=3008 l=564
+ ad=0 pd=0 as=0 ps=0 
M3617 GND pd2_clearIR PD_1xx000x0 GND efet w=3008 l=564
+ ad=0 pd=0 as=0 ps=0 
M3618 GND pd3 pd3_clearIR GND efet w=7896 l=564
+ ad=0 pd=0 as=1.02674e+07 ps=28764 
M3619 pd5_clearIR pd5 GND GND efet w=8037 l=705
+ ad=9.48103e+06 pd=26696 as=0 ps=0 
M3620 GND pd0 pd0_clearIR GND efet w=7896 l=658
+ ad=0 pd=0 as=9.02156e+06 ps=28200 
M3621 pd1_clearIR pd1 GND GND efet w=7990 l=658
+ ad=9.00388e+06 pd=28012 as=0 ps=0 
M3622 n_1662 n_1124 GND GND efet w=4606 l=658
+ ad=6.25589e+06 pd=18612 as=0 ps=0 
M3623 GND clearIR pd4_clearIR GND efet w=3055 l=611
+ ad=0 pd=0 as=8.68579e+06 ps=27824 
M3624 GND notRdy0 fetch GND efet w=3572 l=564
+ ad=0 pd=0 as=7.76684e+06 ps=18800 
M3625 n_1662 n_1662 Vdd GND dfet w=846 l=2162
+ ad=1.44115e+07 pd=44556 as=0 ps=0 
M3626 GND op_T__bit n_513 GND efet w=4512 l=658
+ ad=0 pd=0 as=1.08948e+07 ps=30268 
M3627 n_1426 n_270 GND GND efet w=3572 l=658
+ ad=5.69922e+06 pd=15228 as=0 ps=0 
M3628 n_845 n_1662 n_1426 GND efet w=3760 l=564
+ ad=0 pd=0 as=0 ps=0 
M3629 n_511 n_553 n_845 GND efet w=5264 l=564
+ ad=4.52403e+06 pd=13724 as=0 ps=0 
M3630 Vdd n_1055 n_1055 GND dfet w=940 l=1222
+ ad=0 pd=0 as=4.3102e+07 ps=162432 
M3631 n_1154 n_959 GND GND efet w=4700 l=564
+ ad=0 pd=0 as=0 ps=0 
M3632 n_19 n_770 GND GND efet w=3290 l=658
+ ad=6.9451e+06 pd=17108 as=0 ps=0 
M3633 GND n_1708 n_19 GND efet w=3760 l=564
+ ad=0 pd=0 as=0 ps=0 
M3634 GND n_853 n_1517 GND efet w=4371 l=611
+ ad=0 pd=0 as=0 ps=0 
M3635 n_1055 n_771 GND GND efet w=2444 l=658
+ ad=0 pd=0 as=0 ps=0 
M3636 n_19 cclk pipeUNK18 GND efet w=1128 l=846
+ ad=0 pd=0 as=1.5463e+06 ps=6580 
M3637 n_1231 cclk pipeUNK21 GND efet w=1034 l=752
+ ad=0 pd=0 as=3.6316e+06 ps=11844 
M3638 n_14 n_671 GND GND efet w=3478 l=658
+ ad=0 pd=0 as=0 ps=0 
M3639 n_1550 n_781 GND GND efet w=3760 l=658
+ ad=3.00424e+06 pd=10528 as=0 ps=0 
M3640 n_845 n_1573 n_1550 GND efet w=4700 l=564
+ ad=0 pd=0 as=0 ps=0 
M3641 GND pipeUNK17 n_511 GND efet w=6016 l=658
+ ad=0 pd=0 as=0 ps=0 
M3642 n_14 n_323 GND GND efet w=4418 l=564
+ ad=0 pd=0 as=0 ps=0 
M3643 n_959 short_circuit_branch_add GND GND efet w=15040 l=658
+ ad=1.5357e+07 pd=46060 as=0 ps=0 
M3644 n_323 cp1 n_959 GND efet w=1128 l=752
+ ad=1.37842e+06 pd=6392 as=0 ps=0 
M3645 GND pipeUNK18 n_850 GND efet w=7285 l=611
+ ad=0 pd=0 as=6.83906e+06 ps=18612 
M3646 Vdd n_1619 n_1619 GND dfet w=940 l=1598
+ ad=0 pd=0 as=8.60626e+06 ps=29516 
M3647 n_1619 n_1448 GND GND efet w=2820 l=658
+ ad=1.05944e+07 pd=32336 as=0 ps=0 
M3648 n_1619 n_182 GND GND efet w=2820 l=658
+ ad=0 pd=0 as=0 ps=0 
M3649 n_465 n_465 Vdd GND dfet w=846 l=658
+ ad=2.07646e+06 pd=8460 as=0 ps=0 
M3650 Vdd n_1446 n_1446 GND dfet w=940 l=1222
+ ad=0 pd=0 as=4.78028e+06 ps=15228 
M3651 n_850 n_850 Vdd GND dfet w=940 l=1504
+ ad=1.22114e+07 pd=37976 as=0 ps=0 
M3652 GND pipeUNK20 n_959 GND efet w=15322 l=564
+ ad=0 pd=0 as=0 ps=0 
M3653 n_14 cclk pipeUNK20 GND efet w=1128 l=752
+ ad=0 pd=0 as=1.79371e+06 ps=7332 
M3654 pipeBRtaken cclk n_586 GND efet w=1316 l=658
+ ad=3.11911e+06 pd=9024 as=0 ps=0 
M3655 Vdd n_959 n_959 GND dfet w=752 l=752
+ ad=0 pd=0 as=5.82292e+06 ps=21244 
M3656 GND n_206 n_465 GND efet w=7097 l=611
+ ad=0 pd=0 as=1.01526e+07 ps=28388 
M3657 n_1446 n_771 GND GND efet w=4982 l=564
+ ad=8.31468e+06 pd=25192 as=0 ps=0 
M3658 GND n_850 n_1446 GND efet w=4230 l=658
+ ad=0 pd=0 as=0 ps=0 
M3659 short_circuit_branch_add cp1 n_1570 GND efet w=1222 l=752
+ ad=1.75836e+07 pd=49444 as=1.50212e+06 ps=6580 
M3660 short_circuit_branch_add n_771 n_465 GND efet w=1692 l=752
+ ad=0 pd=0 as=0 ps=0 
M3661 n_206 n_1446 short_circuit_branch_add GND efet w=1692 l=658
+ ad=1.66028e+07 pd=43804 as=0 ps=0 
M3662 short_circuit_branch_add n_850 GND GND efet w=7144 l=564
+ ad=0 pd=0 as=0 ps=0 
M3663 n_1472 cp1 D1x1 GND efet w=1316 l=658
+ ad=2.50942e+06 pd=10152 as=0 ps=0 
M3664 n_1275 pipeBRtaken GND GND efet w=9165 l=611
+ ad=1.44292e+07 pd=38540 as=0 ps=0 
M3665 Vdd n_1275 n_1275 GND dfet w=940 l=1034
+ ad=0 pd=0 as=2.35038e+06 ps=8272 
M3666 Vdd dpc36_nIPC dpc36_nIPC GND dfet w=940 l=1222
+ ad=0 pd=0 as=2.40339e+07 ps=78208 
M3667 n_1480 n_1472 GND GND efet w=15134 l=564
+ ad=2.7586e+07 pd=63168 as=0 ps=0 
M3668 dpc36_nIPC n_1570 n_1480 GND efet w=14805 l=517
+ ad=1.68768e+07 pd=45684 as=0 ps=0 
M3669 GND notRdy0 n_1275 GND efet w=4606 l=564
+ ad=0 pd=0 as=0 ps=0 
M3670 n_1705 n_1705 Vdd GND dfet w=940 l=1034
+ ad=2.3115e+07 pd=78396 as=0 ps=0 
M3671 GND ONEBYTE n_1275 GND efet w=4277 l=611
+ ad=0 pd=0 as=0 ps=0 
M3672 n_1275 cp1 n_1581 GND efet w=1222 l=658
+ ad=0 pd=0 as=1.36074e+06 ps=6768 
M3673 n_506 cclk n_1602 GND efet w=1128 l=752
+ ad=0 pd=0 as=1.41376e+06 ps=7332 
M3674 n_1683 cclk n_1090 GND efet w=1128 l=752
+ ad=1.47561e+06 pd=5640 as=0 ps=0 
M3675 n_11 cclk n_55 GND efet w=1128 l=846
+ ad=0 pd=0 as=1.41376e+06 ps=6956 
M3676 n_1037 cclk n_266 GND efet w=1081 l=893
+ ad=0 pd=0 as=1.30773e+06 ps=5828 
M3677 n_272 cclk n_1162 GND efet w=1222 l=846
+ ad=0 pd=0 as=1.31656e+06 ps=6956 
M3678 n_952 cclk n_1509 GND efet w=1128 l=752
+ ad=0 pd=0 as=1.31656e+06 ps=7144 
M3679 n_824 cclk n_398 GND efet w=1128 l=752
+ ad=0 pd=0 as=1.58164e+06 ps=5828 
M3680 Vdd n_1295 n_1295 GND dfet w=846 l=940
+ ad=0 pd=0 as=1.16812e+07 ps=37036 
M3681 GND n_1527 n_1295 GND efet w=6768 l=658
+ ad=0 pd=0 as=7.13065e+06 ps=19740 
M3682 n_830 n_1505 GND GND efet w=4888 l=658
+ ad=7.74917e+06 pd=21056 as=0 ps=0 
M3683 Vdd n_830 n_830 GND dfet w=846 l=1410
+ ad=0 pd=0 as=1.11069e+07 ps=31584 
M3684 Vdd n_1596 n_1596 GND dfet w=846 l=1034
+ ad=0 pd=0 as=1.12129e+07 ps=37412 
M3685 GND n_1602 n_1596 GND efet w=6768 l=564
+ ad=0 pd=0 as=7.32504e+06 ps=19176 
M3686 GND n_43 n_830 GND efet w=2491 l=611
+ ad=0 pd=0 as=0 ps=0 
M3687 Vdd n_966 n_966 GND dfet w=799 l=987
+ ad=0 pd=0 as=1.05148e+07 ps=36660 
M3688 GND n_1683 n_966 GND efet w=6815 l=611
+ ad=0 pd=0 as=7.35155e+06 ps=19552 
M3689 n_1238 n_1295 GND GND efet w=2256 l=658
+ ad=2.96006e+06 pd=9964 as=0 ps=0 
M3690 n_1047 n_830 GND GND efet w=2162 l=752
+ ad=2.95122e+06 pd=9400 as=0 ps=0 
M3691 n_628 n_55 GND GND efet w=5593 l=517
+ ad=7.6078e+06 pd=20868 as=0 ps=0 
M3692 Vdd n_628 n_628 GND dfet w=987 l=1269
+ ad=0 pd=0 as=8.35886e+06 ps=30268 
M3693 n_1238 n_1238 Vdd GND dfet w=846 l=1316
+ ad=1.17607e+07 pd=33464 as=0 ps=0 
M3694 n_1271 n_1596 GND GND efet w=2350 l=658
+ ad=3.26048e+06 pd=9776 as=0 ps=0 
M3695 n_462 cclk n_878 GND efet w=1222 l=846
+ ad=0 pd=0 as=1.49328e+06 ps=5828 
M3696 n_598 cclk n_176 GND efet w=1128 l=846
+ ad=1.34307e+06 pd=5640 as=0 ps=0 
M3697 n_442 cclk n_509 GND efet w=1128 l=846
+ ad=0 pd=0 as=1.27238e+06 ps=6956 
M3698 n_1211 cclk n_897 GND efet w=1128 l=940
+ ad=0 pd=0 as=1.3254e+06 ps=5452 
M3699 n_182 cclk n_265 GND efet w=1128 l=940
+ ad=0 pd=0 as=1.36958e+06 ps=6768 
M3700 Vdd n_525 n_525 GND dfet w=987 l=1175
+ ad=0 pd=0 as=9.17177e+06 ps=30268 
M3701 GND n_266 n_525 GND efet w=5405 l=517
+ ad=0 pd=0 as=8.35886e+06 ps=21244 
M3702 n_21 n_1162 GND GND efet w=5076 l=564
+ ad=7.70499e+06 pd=20868 as=0 ps=0 
M3703 Vdd n_21 n_21 GND dfet w=846 l=1222
+ ad=0 pd=0 as=1.11245e+07 ps=31960 
M3704 GND cclk n_628 GND efet w=2350 l=470
+ ad=0 pd=0 as=0 ps=0 
M3705 n_525 cclk GND GND efet w=2350 l=564
+ ad=0 pd=0 as=0 ps=0 
M3706 n_611 n_1509 GND GND efet w=5076 l=564
+ ad=7.36922e+06 pd=21244 as=0 ps=0 
M3707 Vdd n_611 n_611 GND dfet w=846 l=1316
+ ad=0 pd=0 as=1.12217e+07 ps=31772 
M3708 n_1047 n_1047 Vdd GND dfet w=940 l=1410
+ ad=1.07622e+07 pd=33840 as=0 ps=0 
M3709 n_1635 n_966 GND GND efet w=2256 l=564
+ ad=2.97773e+06 pd=9776 as=0 ps=0 
M3710 Vdd n_1295 dpc25_SBDB GND dfet w=1034 l=940
+ ad=0 pd=0 as=1.19551e+07 ps=29704 
M3711 GND n_1238 dpc25_SBDB GND efet w=8836 l=752
+ ad=0 pd=0 as=0 ps=0 
M3712 Vdd n_830 dpc23_SBAC GND dfet w=940 l=940
+ ad=0 pd=0 as=1.76455e+07 ps=37788 
M3713 n_1271 n_1271 Vdd GND dfet w=846 l=1410
+ ad=1.10362e+07 pd=33652 as=0 ps=0 
M3714 n_1335 n_628 GND GND efet w=2350 l=470
+ ad=3.24281e+06 pd=10152 as=0 ps=0 
M3715 GND n_43 n_21 GND efet w=2350 l=658
+ ad=0 pd=0 as=0 ps=0 
M3716 Vdd n_321 n_321 GND dfet w=940 l=940
+ ad=0 pd=0 as=1.05944e+07 ps=36848 
M3717 GND n_398 n_321 GND efet w=6862 l=658
+ ad=0 pd=0 as=7.00695e+06 ps=20304 
M3718 n_1635 n_1635 Vdd GND dfet w=846 l=1316
+ ad=1.08594e+07 pd=33840 as=0 ps=0 
M3719 Vdd n_1596 dpc27_SBADH GND dfet w=846 l=846
+ ad=0 pd=0 as=1.13984e+07 ps=26508 
M3720 dpc23_SBAC n_1247 GND GND efet w=7144 l=564
+ ad=0 pd=0 as=0 ps=0 
M3721 GND n_1047 dpc23_SBAC GND efet w=7238 l=658
+ ad=0 pd=0 as=0 ps=0 
M3722 GND n_1271 dpc27_SBADH GND efet w=9024 l=658
+ ad=0 pd=0 as=0 ps=0 
M3723 Vdd n_966 dpc29_0ADH17 GND dfet w=940 l=846
+ ad=0 pd=0 as=1.07534e+07 ps=24628 
M3724 n_1335 n_1335 Vdd GND dfet w=846 l=1128
+ ad=9.39267e+06 pd=33464 as=0 ps=0 
M3725 GND n_1635 dpc29_0ADH17 GND efet w=9071 l=611
+ ad=0 pd=0 as=0 ps=0 
M3726 Vdd n_628 dpc24_ACSB GND dfet w=940 l=752
+ ad=0 pd=0 as=1.57192e+07 ps=36096 
M3727 GND n_525 n_800 GND efet w=2444 l=564
+ ad=0 pd=0 as=3.44604e+06 ps=10152 
M3728 n_228 n_21 GND GND efet w=2444 l=752
+ ad=2.9689e+06 pd=9964 as=0 ps=0 
M3729 GND n_43 n_611 GND efet w=2256 l=564
+ ad=0 pd=0 as=0 ps=0 
M3730 Vdd n_631 n_631 GND dfet w=846 l=940
+ ad=0 pd=0 as=1.08771e+07 ps=37224 
M3731 GND n_878 n_631 GND efet w=6862 l=658
+ ad=0 pd=0 as=7.28086e+06 ps=20116 
M3732 n_800 n_800 Vdd GND dfet w=940 l=1128
+ ad=9.71076e+06 pd=34028 as=0 ps=0 
M3733 Vdd n_525 dpc26_ACDB GND dfet w=846 l=846
+ ad=0 pd=0 as=1.68061e+07 ps=40232 
M3734 n_255 n_611 GND GND efet w=2256 l=752
+ ad=2.79218e+06 pd=9588 as=0 ps=0 
M3735 Vdd n_1260 n_1260 GND dfet w=846 l=940
+ ad=0 pd=0 as=1.06032e+07 ps=37412 
M3736 GND n_598 n_1260 GND efet w=6862 l=658
+ ad=0 pd=0 as=6.71536e+06 ps=19740 
M3737 n_1270 n_509 GND GND efet w=5029 l=517
+ ad=8.1733e+06 pd=20868 as=0 ps=0 
M3738 Vdd n_1270 n_1270 GND dfet w=940 l=1410
+ ad=0 pd=0 as=1.01702e+07 ps=31584 
M3739 Vdd n_1369 n_1369 GND dfet w=846 l=940
+ ad=0 pd=0 as=1.12747e+07 ps=37600 
M3740 GND n_897 n_1369 GND efet w=6956 l=658
+ ad=0 pd=0 as=7.12182e+06 ps=20304 
M3741 GND n_43 n_1270 GND efet w=2538 l=752
+ ad=0 pd=0 as=0 ps=0 
M3742 n_228 n_228 Vdd GND dfet w=940 l=1410
+ ad=1.14603e+07 pd=33652 as=0 ps=0 
M3743 Vdd n_21 dpc30_ADHPCH GND dfet w=940 l=1034
+ ad=0 pd=0 as=1.66735e+07 ps=41924 
M3744 DA_C01 DA_C01 Vdd GND dfet w=940 l=1504
+ ad=1.45175e+07 pd=47188 as=0 ps=0 
M3745 naluresult0 dpc17_SUMS n_AxBxC_0 GND efet w=940 l=658
+ ad=0 pd=0 as=0 ps=0 
M3746 n_AxBxC_0 _AxB_0_nC0in GND GND efet w=2303 l=611
+ ad=0 pd=0 as=0 ps=0 
M3747 _AxB_0_nC0in n_AxB_0 GND GND efet w=1692 l=658
+ ad=5.77874e+06 pd=20868 as=0 ps=0 
M3748 n_AxB_0 n_AxB_0 Vdd GND dfet w=846 l=1598
+ ad=1.14691e+07 pd=36096 as=0 ps=0 
M3749 GND n_105 _AxB_0_nC0in GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M3750 C01 C01 Vdd GND dfet w=940 l=940
+ ad=9.88748e+06 pd=36096 as=0 ps=0 
M3751 Vdd n_936 n_936 GND dfet w=846 l=1598
+ ad=0 pd=0 as=2.14273e+07 ps=75576 
M3752 Vdd A_B1 A_B1 GND dfet w=846 l=1504
+ ad=0 pd=0 as=7.64314e+06 ps=23688 
M3753 Vdd _AxB_0_nC0in _AxB_0_nC0in GND dfet w=940 l=1504
+ ad=0 pd=0 as=8.42954e+06 ps=27636 
M3754 Vdd nC01 nC01 GND dfet w=846 l=1504
+ ad=0 pd=0 as=1.00112e+07 ps=31584 
M3755 n_936 nA_B1 GND GND efet w=1692 l=564
+ ad=6.21171e+06 pd=17672 as=0 ps=0 
M3756 nC01 C01 GND GND efet w=1692 l=564
+ ad=2.50942e+06 pd=9024 as=0 ps=0 
M3757 DA_C01 n_A_B_0 GND GND efet w=2350 l=564
+ ad=7.6078e+06 pd=20116 as=0 ps=0 
M3758 n_1707 n_936 GND GND efet w=5076 l=564
+ ad=2.86286e+06 pd=11280 as=0 ps=0 
M3759 n_319 DA_C01 n_1707 GND efet w=5076 l=564
+ ad=5.88478e+06 pd=18048 as=0 ps=0 
M3760 n_1354 nA_B0 DA_C01 GND efet w=4982 l=564
+ ad=2.34154e+06 pd=10904 as=0 ps=0 
M3761 GND notalucin n_1354 GND efet w=4982 l=658
+ ad=0 pd=0 as=0 ps=0 
M3762 GND n_A_B_1 A_B1 GND efet w=2256 l=658
+ ad=0 pd=0 as=5.07186e+06 ps=15980 
M3763 n_1510 A_B1 GND GND efet w=5076 l=564
+ ad=2.79218e+06 pd=11280 as=0 ps=0 
M3764 nC12 C01 n_1510 GND efet w=5076 l=564
+ ad=7.24552e+06 pd=21620 as=0 ps=0 
M3765 n_AxB_1 dpc16_EORS naluresult1 GND efet w=1034 l=752
+ ad=4.02038e+06 pd=12784 as=0 ps=0 
M3766 GND AxB1 n_AxB_1 GND efet w=2726 l=564
+ ad=0 pd=0 as=0 ps=0 
M3767 AxB1 n_936 GND GND efet w=1692 l=564
+ ad=4.87747e+06 pd=15416 as=0 ps=0 
M3768 GND n_A_B_1 AxB1 GND efet w=1692 l=658
+ ad=0 pd=0 as=0 ps=0 
M3769 GND n_936 nC12 GND efet w=2444 l=564
+ ad=0 pd=0 as=0 ps=0 
M3770 n_1388 AxB1 GND GND efet w=3290 l=564
+ ad=1.85556e+06 pd=7708 as=0 ps=0 
M3771 n_AxBxC_1 nC01 n_1388 GND efet w=3290 l=564
+ ad=7.46642e+06 pd=20304 as=0 ps=0 
M3772 Vdd n_AxBxC_1 n_AxBxC_1 GND dfet w=940 l=1598
+ ad=0 pd=0 as=4.17059e+06 ps=9964 
M3773 n_319 n_319 Vdd GND dfet w=846 l=1504
+ ad=2.97155e+07 pd=102272 as=0 ps=0 
M3774 n_388 n_388 Vdd GND dfet w=940 l=1222
+ ad=2.75506e+07 pd=104152 as=0 ps=0 
M3775 n_388 DA_C01 GND GND efet w=3149 l=611
+ ad=1.31921e+07 pd=35532 as=0 ps=0 
M3776 n_388 DA_AxB2 GND GND efet w=3243 l=611
+ ad=0 pd=0 as=0 ps=0 
M3777 n_AxBxC_1 n_AxB1__C01 GND GND efet w=2585 l=611
+ ad=0 pd=0 as=0 ps=0 
M3778 naluresult1 dpc17_SUMS n_AxBxC_1 GND efet w=1128 l=752
+ ad=0 pd=0 as=0 ps=0 
M3779 n_388 n_936 GND GND efet w=2538 l=564
+ ad=0 pd=0 as=0 ps=0 
M3780 GND AxB1 n_388 GND efet w=2820 l=564
+ ad=0 pd=0 as=0 ps=0 
M3781 n_AxB1__C01 AxB1 GND GND efet w=1692 l=564
+ ad=4.62123e+06 pd=15604 as=0 ps=0 
M3782 n_AxB_1 n_AxB_1 Vdd GND dfet w=846 l=1504
+ ad=3.77297e+06 pd=11280 as=0 ps=0 
M3783 AxB1 AxB1 Vdd GND dfet w=846 l=1504
+ ad=2.14361e+07 pd=75576 as=0 ps=0 
M3784 GND nC01 n_AxB1__C01 GND efet w=3290 l=658
+ ad=0 pd=0 as=0 ps=0 
M3785 Vdd nC12 nC12 GND dfet w=846 l=846
+ ad=0 pd=0 as=1.28829e+07 ps=43240 
M3786 n_AxB1__C01 n_AxB1__C01 Vdd GND dfet w=940 l=1598
+ ad=6.81256e+06 pd=21432 as=0 ps=0 
M3787 A_B2 A_B2 Vdd GND dfet w=846 l=1504
+ ad=7.8552e+06 pd=25004 as=0 ps=0 
M3788 Vdd C12 C12 GND dfet w=846 l=1504
+ ad=0 pd=0 as=9.30431e+06 ps=32336 
M3789 nA_B2 dpc14_SRS naluresult1 GND efet w=1034 l=658
+ ad=0 pd=0 as=0 ps=0 
M3790 naluresult2 dpc13_ORS n_A_B_2 GND efet w=1128 l=658
+ ad=1.46324e+07 pd=41172 as=8.95087e+06 ps=26132 
M3791 GND dpc12_0ADD alua2 GND efet w=1128 l=564
+ ad=0 pd=0 as=5.06303e+06 ps=13348 
M3792 alua2 dpc11_SBADD sb2 GND efet w=1128 l=658
+ ad=0 pd=0 as=0 ps=0 
M3793 n_A_B_2 alua2 GND GND efet w=2914 l=658
+ ad=0 pd=0 as=0 ps=0 
M3794 GND alub2 n_A_B_2 GND efet w=3008 l=564
+ ad=0 pd=0 as=0 ps=0 
M3795 Vdd n_A_B_2 n_A_B_2 GND dfet w=846 l=1974
+ ad=0 pd=0 as=3.03782e+07 ps=99828 
M3796 adl3 dpc10_ADLADD alub3 GND efet w=1034 l=658
+ ad=0 pd=0 as=5.0807e+06 ps=13536 
M3797 alub3 dpc8_nDBADD n_1621 GND efet w=1034 l=752
+ ad=0 pd=0 as=8.16446e+06 ps=26132 
M3798 alub3 dpc9_DBADD idb3 GND efet w=1128 l=564
+ ad=0 pd=0 as=1.86086e+07 ps=51700 
M3799 GND idb3 n_1621 GND efet w=5828 l=658
+ ad=0 pd=0 as=0 ps=0 
M3800 n_1621 n_1621 Vdd GND dfet w=846 l=1598
+ ad=3.03075e+06 pd=8084 as=0 ps=0 
M3801 n_313 alua3 GND GND efet w=5734 l=564
+ ad=3.23398e+06 pd=12596 as=0 ps=0 
M3802 nA_B3 alub3 n_313 GND efet w=5734 l=564
+ ad=1.05413e+07 pd=28764 as=0 ps=0 
M3803 Vdd nA_B3 nA_B3 GND dfet w=940 l=1974
+ ad=0 pd=0 as=8.7123e+06 ps=23312 
M3804 C12 nC12 GND GND efet w=1598 l=564
+ ad=2.38572e+06 pd=9024 as=0 ps=0 
M3805 A_B2 n_A_B_2 GND GND efet w=1692 l=752
+ ad=2.70382e+06 pd=8272 as=0 ps=0 
M3806 n_716 A_B2 n_AxB_2 GND efet w=3431 l=611
+ ad=1.74069e+06 pd=7896 as=7.13065e+06 ps=22184 
M3807 naluresult2 dpc15_ANDS nA_B2 GND efet w=1128 l=752
+ ad=0 pd=0 as=0 ps=0 
M3808 n_AxB_2 dpc16_EORS naluresult2 GND efet w=1128 l=658
+ ad=0 pd=0 as=0 ps=0 
M3809 GND nA_B2 n_716 GND efet w=3196 l=564
+ ad=0 pd=0 as=0 ps=0 
M3810 C23 n_A_B_2 GND GND efet w=2632 l=564
+ ad=8.80949e+06 pd=24628 as=0 ps=0 
M3811 n_433 nA_B2 C23 GND efet w=5170 l=564
+ ad=4.418e+06 pd=15228 as=0 ps=0 
M3812 GND nC12 n_433 GND efet w=6815 l=611
+ ad=0 pd=0 as=0 ps=0 
M3813 n_1572 n_AxB_2 GND GND efet w=3384 l=658
+ ad=1.90858e+06 pd=7896 as=0 ps=0 
M3814 n_AxBxC_2 C12 n_1572 GND efet w=3384 l=470
+ ad=8.53558e+06 pd=22372 as=0 ps=0 
M3815 Vdd n_AxBxC_2 n_AxBxC_2 GND dfet w=846 l=1598
+ ad=0 pd=0 as=3.99387e+06 ps=9776 
M3816 DA_AxB2 DA_AB2 GND GND efet w=3149 l=517
+ ad=1.13454e+07 pd=29516 as=0 ps=0 
M3817 n_1610 AxB3 GND GND efet w=3854 l=658
+ ad=5.33694e+06 pd=17296 as=0 ps=0 
M3818 GND DA_AB2 n_1610 GND efet w=2538 l=564
+ ad=0 pd=0 as=0 ps=0 
M3819 n_1610 n_1610 Vdd GND dfet w=940 l=1504
+ ad=2.07558e+07 pd=68620 as=0 ps=0 
M3820 naluresult2 dpc17_SUMS n_AxBxC_2 GND efet w=1034 l=658
+ ad=0 pd=0 as=0 ps=0 
M3821 n_AxBxC_2 _AxB_2_nC12 GND GND efet w=2585 l=611
+ ad=0 pd=0 as=0 ps=0 
M3822 _AxB_2_nC12 n_AxB_2 GND GND efet w=1692 l=470
+ ad=5.70806e+06 pd=19740 as=0 ps=0 
M3823 nA_B3 dpc14_SRS naluresult2 GND efet w=1034 l=658
+ ad=0 pd=0 as=0 ps=0 
M3824 naluresult3 dpc13_ORS n_A_B_3 GND efet w=1222 l=658
+ ad=1.64703e+07 pd=47000 as=9.31314e+06 ps=26508 
M3825 GND dpc12_0ADD alua3 GND efet w=1222 l=658
+ ad=0 pd=0 as=4.87747e+06 ps=13536 
M3826 alua3 dpc11_SBADD sb3 GND efet w=1128 l=658
+ ad=0 pd=0 as=0 ps=0 
M3827 adl4 dpc10_ADLADD alub4 GND efet w=1034 l=564
+ ad=0 pd=0 as=4.99234e+06 ps=13536 
M3828 alub4 dpc8_nDBADD n_478 GND efet w=1128 l=846
+ ad=0 pd=0 as=8.13796e+06 ps=25944 
M3829 alub4 dpc9_DBADD idb4 GND efet w=1175 l=799
+ ad=0 pd=0 as=1.92536e+07 ps=52828 
M3830 GND idb4 n_478 GND efet w=5828 l=658
+ ad=0 pd=0 as=0 ps=0 
M3831 n_478 n_478 Vdd GND dfet w=846 l=1598
+ ad=2.93355e+06 pd=8084 as=0 ps=0 
M3832 n_A_B_3 alua3 GND GND efet w=3008 l=564
+ ad=0 pd=0 as=0 ps=0 
M3833 GND alub3 n_A_B_3 GND efet w=2914 l=658
+ ad=0 pd=0 as=0 ps=0 
M3834 Vdd n_A_B_3 n_A_B_3 GND dfet w=940 l=2068
+ ad=0 pd=0 as=1.21053e+07 ps=39104 
M3835 n_185 alua4 GND GND efet w=5734 l=564
+ ad=3.23398e+06 pd=12596 as=0 ps=0 
M3836 nA_B4 alub4 n_185 GND efet w=5734 l=658
+ ad=9.80796e+06 pd=27824 as=0 ps=0 
M3837 Vdd nA_B4 nA_B4 GND dfet w=846 l=1974
+ ad=0 pd=0 as=1.42525e+07 ps=40796 
M3838 naluresult3 dpc15_ANDS nA_B3 GND efet w=1128 l=658
+ ad=0 pd=0 as=0 ps=0 
M3839 n_AxB_2 n_AxB_2 Vdd GND dfet w=846 l=1504
+ ad=1.05767e+07 pd=35908 as=0 ps=0 
M3840 GND C12 _AxB_2_nC12 GND efet w=2444 l=658
+ ad=0 pd=0 as=0 ps=0 
M3841 DA_AB2 nA_B2 GND GND efet w=2538 l=564
+ ad=8.56208e+06 pd=28576 as=0 ps=0 
M3842 C23 C23 Vdd GND dfet w=940 l=846
+ ad=9.89632e+06 pd=35908 as=0 ps=0 
M3843 Vdd n_988 n_988 GND dfet w=940 l=1598
+ ad=0 pd=0 as=8.30584e+06 ps=28576 
M3844 Vdd A_B3 A_B3 GND dfet w=940 l=1598
+ ad=0 pd=0 as=7.28086e+06 ps=23500 
M3845 n_988 nA_B3 GND GND efet w=1598 l=658
+ ad=6.37959e+06 pd=18424 as=0 ps=0 
M3846 Vdd _AxB_2_nC12 _AxB_2_nC12 GND dfet w=752 l=1598
+ ad=0 pd=0 as=8.5179e+06 ps=27448 
M3847 Vdd nC23 nC23 GND dfet w=940 l=1504
+ ad=0 pd=0 as=1.00907e+07 ps=31960 
M3848 DA_AB2 DA_AB2 Vdd GND dfet w=846 l=1504
+ ad=1.51891e+07 pd=55460 as=0 ps=0 
M3849 DA_AxB2 DA_AxB2 Vdd GND dfet w=940 l=1598
+ ad=7.59012e+06 pd=25192 as=0 ps=0 
M3850 DA_AxB2 n_A_B_2 GND GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M3851 nC23 C23 GND GND efet w=1692 l=564
+ ad=3.00424e+06 pd=8836 as=0 ps=0 
M3852 GND n_A_B_3 A_B3 GND efet w=2256 l=658
+ ad=0 pd=0 as=5.23975e+06 ps=18424 
M3853 n_AxB_3 dpc16_EORS naluresult3 GND efet w=1128 l=658
+ ad=4.1971e+06 pd=13160 as=0 ps=0 
M3854 GND AxB3 n_AxB_3 GND efet w=2726 l=564
+ ad=0 pd=0 as=0 ps=0 
M3855 AxB3 n_988 GND GND efet w=1692 l=564
+ ad=5.23091e+06 pd=17296 as=0 ps=0 
M3856 GND n_A_B_3 AxB3 GND efet w=1692 l=658
+ ad=0 pd=0 as=0 ps=0 
M3857 n_924 A_B3 GND GND efet w=4982 l=564
+ ad=2.80985e+06 pd=11092 as=0 ps=0 
M3858 nC34 C23 n_924 GND efet w=4982 l=564
+ ad=9.10108e+06 pd=25192 as=0 ps=0 
M3859 GND n_988 nC34 GND efet w=2444 l=564
+ ad=0 pd=0 as=0 ps=0 
M3860 n_136 AxB3 GND GND efet w=3290 l=564
+ ad=1.85556e+06 pd=7708 as=0 ps=0 
M3861 n_AxBxC_3 nC23 n_136 GND efet w=3290 l=564
+ ad=7.31621e+06 pd=19740 as=0 ps=0 
M3862 Vdd n_AxBxC_3 n_AxBxC_3 GND dfet w=940 l=1598
+ ad=0 pd=0 as=4.25895e+06 ps=9964 
M3863 n_AxBxC_3 n_AxB3__C23 GND GND efet w=2444 l=564
+ ad=0 pd=0 as=0 ps=0 
M3864 naluresult3 dpc17_SUMS n_AxBxC_3 GND efet w=1034 l=752
+ ad=0 pd=0 as=0 ps=0 
M3865 GND DC34 nC34 GND efet w=2538 l=564
+ ad=0 pd=0 as=0 ps=0 
M3866 n_AxB3__C23 AxB3 GND GND efet w=1692 l=564
+ ad=4.8598e+06 pd=15792 as=0 ps=0 
M3867 GND nC23 n_AxB3__C23 GND efet w=3243 l=611
+ ad=0 pd=0 as=0 ps=0 
M3868 n_AxB_3 n_AxB_3 Vdd GND dfet w=752 l=1598
+ ad=3.93202e+06 pd=11468 as=0 ps=0 
M3869 AxB3 AxB3 Vdd GND dfet w=846 l=1504
+ ad=3.35149e+07 pd=119756 as=0 ps=0 
M3870 nC34 nC34 Vdd GND dfet w=846 l=940
+ ad=1.19728e+07 pd=41548 as=0 ps=0 
M3871 A_B4 A_B4 Vdd GND dfet w=987 l=1457
+ ad=6.98928e+06 pd=23124 as=0 ps=0 
M3872 nA_B4 dpc14_SRS naluresult3 GND efet w=1034 l=752
+ ad=0 pd=0 as=0 ps=0 
M3873 naluresult4 dpc13_ORS n_A_B_4 GND efet w=1128 l=658
+ ad=1.44469e+07 pd=42112 as=8.72997e+06 ps=25944 
M3874 GND dpc12_0ADD alua4 GND efet w=1128 l=658
+ ad=0 pd=0 as=4.3208e+06 ps=12596 
M3875 alua4 dpc11_SBADD sb4 GND efet w=1034 l=752
+ ad=0 pd=0 as=0 ps=0 
M3876 adl5 dpc10_ADLADD alub5 GND efet w=940 l=752
+ ad=0 pd=0 as=5.01885e+06 ps=13536 
M3877 alub5 dpc8_nDBADD n_1383 GND efet w=1128 l=658
+ ad=0 pd=0 as=8.56208e+06 ps=25944 
M3878 alub5 dpc9_DBADD idb5 GND efet w=1175 l=799
+ ad=0 pd=0 as=1.5357e+07 ps=42112 
M3879 GND idb5 n_1383 GND efet w=5734 l=658
+ ad=0 pd=0 as=0 ps=0 
M3880 n_1383 n_1383 Vdd GND dfet w=752 l=1598
+ ad=2.93355e+06 pd=8084 as=0 ps=0 
M3881 n_A_B_4 alua4 GND GND efet w=2914 l=564
+ ad=0 pd=0 as=0 ps=0 
M3882 GND alub4 n_A_B_4 GND efet w=3008 l=564
+ ad=0 pd=0 as=0 ps=0 
M3883 Vdd n_A_B_4 n_A_B_4 GND dfet w=940 l=2068
+ ad=0 pd=0 as=1.45441e+07 ps=49256 
M3884 A_B4 n_A_B_4 GND GND efet w=1692 l=564
+ ad=4.93049e+06 pd=14852 as=0 ps=0 
M3885 n_AxB3__C23 n_AxB3__C23 Vdd GND dfet w=846 l=1598
+ ad=6.7507e+06 pd=21620 as=0 ps=0 
M3886 n_972 n_A_B_2 GND GND efet w=5264 l=658
+ ad=1.49417e+07 pd=40420 as=0 ps=0 
M3887 GND n_319 n_972 GND efet w=6345 l=611
+ ad=0 pd=0 as=0 ps=0 
M3888 adl0 dpc21_ADDADL alu0 GND efet w=1504 l=752
+ ad=0 pd=0 as=1.42701e+07 ps=39668 
M3889 naluresult0 cclk notalu0 GND efet w=1034 l=752
+ ad=0 pd=0 as=1.62582e+06 ps=7144 
M3890 GND notalu0 alu0 GND efet w=9400 l=564
+ ad=0 pd=0 as=0 ps=0 
M3891 alu0 dpc20_ADDSB06 sb0 GND efet w=1974 l=752
+ ad=0 pd=0 as=0 ps=0 
M3892 alu0 alu0 Vdd GND dfet w=940 l=1222
+ ad=3.13678e+06 pd=9776 as=0 ps=0 
M3893 adl1 dpc21_ADDADL alu1 GND efet w=1504 l=752
+ ad=0 pd=0 as=1.35809e+07 ps=39668 
M3894 naluresult1 cclk notalu1 GND efet w=1081 l=893
+ ad=0 pd=0 as=1.4491e+06 ps=6768 
M3895 GND notalu1 alu1 GND efet w=9588 l=658
+ ad=0 pd=0 as=0 ps=0 
M3896 alu1 dpc20_ADDSB06 sb1 GND efet w=1974 l=752
+ ad=0 pd=0 as=0 ps=0 
M3897 n_700 dpc18_nDAA GND GND efet w=2538 l=564
+ ad=7.5106e+06 pd=23876 as=0 ps=0 
M3898 n_972 n_1610 DC34 GND efet w=5546 l=658
+ ad=0 pd=0 as=9.94934e+06 ps=32712 
M3899 n_972 n_388 DC34 GND efet w=5546 l=564
+ ad=0 pd=0 as=0 ps=0 
M3900 n_700 n_700 Vdd GND dfet w=846 l=1410
+ ad=1.47296e+07 pd=49444 as=0 ps=0 
M3901 n_700 cclk n_1565 GND efet w=1128 l=752
+ ad=0 pd=0 as=1.23704e+06 ps=6392 
M3902 GND dpc18_nDAA DC34 GND efet w=3243 l=611
+ ad=0 pd=0 as=0 ps=0 
M3903 Vdd C34 C34 GND dfet w=940 l=1410
+ ad=0 pd=0 as=2.31415e+07 ps=78960 
M3904 DC34 DC34 Vdd GND dfet w=940 l=940
+ ad=9.56939e+06 pd=33464 as=0 ps=0 
M3905 n_1218 n_1565 GND GND efet w=2444 l=658
+ ad=6.45028e+06 pd=19364 as=0 ps=0 
M3906 GND n_1565 n_1218 GND efet w=2162 l=564
+ ad=0 pd=0 as=0 ps=0 
M3907 C34 nC34 GND GND efet w=1692 l=658
+ ad=2.93355e+06 pd=11280 as=0 ps=0 
M3908 naluresult4 dpc15_ANDS nA_B4 GND efet w=1034 l=658
+ ad=0 pd=0 as=0 ps=0 
M3909 n_AxB_4 dpc16_EORS naluresult4 GND efet w=1034 l=658
+ ad=7.72266e+06 pd=24064 as=0 ps=0 
M3910 n_1559 alua5 GND GND efet w=5734 l=658
+ ad=2.69498e+06 pd=12408 as=0 ps=0 
M3911 nA_B5 alub5 n_1559 GND efet w=5734 l=564
+ ad=1.03381e+07 pd=28200 as=0 ps=0 
M3912 Vdd nA_B5 nA_B5 GND dfet w=846 l=1974
+ ad=0 pd=0 as=8.56208e+06 ps=22936 
M3913 nA_B5 dpc14_SRS naluresult4 GND efet w=1034 l=658
+ ad=0 pd=0 as=0 ps=0 
M3914 naluresult5 dpc13_ORS n_A_B_5 GND efet w=1128 l=752
+ ad=1.64526e+07 pd=47376 as=8.19097e+06 ps=25756 
M3915 GND dpc12_0ADD alua5 GND efet w=1128 l=658
+ ad=0 pd=0 as=4.58588e+06 ps=12972 
M3916 alua5 dpc11_SBADD sb5 GND efet w=1034 l=752
+ ad=0 pd=0 as=0 ps=0 
M3917 n_618 dpc7_SS s6 GND efet w=1128 l=752
+ ad=0 pd=0 as=2.75683e+06 ps=6956 
M3918 s6 dpc6_SBS sb6 GND efet w=1128 l=658
+ ad=0 pd=0 as=0 ps=0 
M3919 sb6 cclk Vdd GND efet w=2068 l=564
+ ad=0 pd=0 as=0 ps=0 
M3920 Vdd n_721 n_721 GND dfet w=940 l=1598
+ ad=0 pd=0 as=3.13678e+06 ps=9400 
M3921 n_721 dpc5_SADL adl7 GND efet w=1410 l=658
+ ad=1.72037e+07 pd=42488 as=2.19575e+07 ps=58844 
M3922 Vdd n_548 n_548 GND dfet w=846 l=1880
+ ad=0 pd=0 as=4.24128e+06 ps=12220 
M3923 x7 dpc3_SBX sb7 GND efet w=1034 l=752
+ ad=0 pd=0 as=0 ps=0 
M3924 n_721 dpc4_SSB sb7 GND efet w=1504 l=752
+ ad=0 pd=0 as=0 ps=0 
M3925 GND nots7 n_721 GND efet w=4136 l=564
+ ad=0 pd=0 as=0 ps=0 
M3926 n_548 s7 GND GND efet w=3102 l=564
+ ad=7.76684e+06 pd=21808 as=0 ps=0 
M3927 n_548 cclk nots7 GND efet w=1128 l=752
+ ad=0 pd=0 as=2.50059e+06 ps=9212 
M3928 n_721 dpc7_SS s7 GND efet w=1128 l=752
+ ad=0 pd=0 as=3.11027e+06 ps=7332 
M3929 s7 dpc6_SBS sb7 GND efet w=1128 l=658
+ ad=0 pd=0 as=0 ps=0 
M3930 sb7 cclk Vdd GND efet w=2068 l=658
+ ad=0 pd=0 as=0 ps=0 
M3931 adl6 dpc10_ADLADD alub6 GND efet w=1128 l=658
+ ad=0 pd=0 as=5.26626e+06 ps=14100 
M3932 alub6 dpc8_nDBADD n_351 GND efet w=1128 l=658
+ ad=0 pd=0 as=8.59743e+06 ps=26320 
M3933 alub6 dpc9_DBADD idb6 GND efet w=1034 l=658
+ ad=0 pd=0 as=1.74423e+07 ps=50948 
M3934 GND idb6 n_351 GND efet w=5640 l=658
+ ad=0 pd=0 as=0 ps=0 
M3935 n_351 n_351 Vdd GND dfet w=846 l=1598
+ ad=3.03075e+06 pd=8084 as=0 ps=0 
M3936 n_A_B_5 alua5 GND GND efet w=3008 l=658
+ ad=0 pd=0 as=0 ps=0 
M3937 GND alub5 n_A_B_5 GND efet w=3008 l=658
+ ad=0 pd=0 as=0 ps=0 
M3938 naluresult5 dpc15_ANDS nA_B5 GND efet w=1034 l=752
+ ad=0 pd=0 as=0 ps=0 
M3939 Vdd n_A_B_5 n_A_B_5 GND dfet w=846 l=2068
+ ad=0 pd=0 as=1.26178e+07 ps=38916 
M3940 n_1483 alua6 GND GND efet w=5734 l=564
+ ad=3.23398e+06 pd=12596 as=0 ps=0 
M3941 nA_B6 alub6 n_1483 GND efet w=5734 l=564
+ ad=9.6224e+06 pd=28200 as=0 ps=0 
M3942 Vdd nA_B6 nA_B6 GND dfet w=940 l=2068
+ ad=0 pd=0 as=2.11092e+07 ps=68808 
M3943 n_1583 nA_B4 n_AxB_4 GND efet w=3102 l=658
+ ad=1.74953e+06 pd=7332 as=0 ps=0 
M3944 GND A_B4 n_1583 GND efet w=3102 l=564
+ ad=0 pd=0 as=0 ps=0 
M3945 C45 n_A_B_4 GND GND efet w=2726 l=564
+ ad=7.54594e+06 pd=20868 as=0 ps=0 
M3946 n_1310 nC34 C45 GND efet w=5123 l=611
+ ad=2.44757e+06 pd=11092 as=0 ps=0 
M3947 GND nA_B4 n_1310 GND efet w=4888 l=658
+ ad=0 pd=0 as=0 ps=0 
M3948 n_375 n_AxB_4 GND GND efet w=3290 l=658
+ ad=1.85556e+06 pd=7708 as=0 ps=0 
M3949 n_AxBxC_4 C34 n_375 GND efet w=3290 l=470
+ ad=8.0496e+06 pd=20868 as=0 ps=0 
M3950 Vdd n_AxBxC_4 n_AxBxC_4 GND dfet w=846 l=1692
+ ad=0 pd=0 as=4.30313e+06 ps=9964 
M3951 naluresult4 dpc17_SUMS n_AxBxC_4 GND efet w=1034 l=658
+ ad=0 pd=0 as=0 ps=0 
M3952 Vdd DA_C45 DA_C45 GND dfet w=846 l=1598
+ ad=0 pd=0 as=1.5896e+07 ps=53956 
M3953 n_AxBxC_4 _AxB_4_nC34 GND GND efet w=2867 l=611
+ ad=0 pd=0 as=0 ps=0 
M3954 _AxB_4_nC34 n_AxB_4 GND GND efet w=1692 l=658
+ ad=4.69192e+06 pd=16732 as=0 ps=0 
M3955 DA_C45 nC45 GND GND efet w=2538 l=564
+ ad=2.61546e+06 pd=10340 as=0 ps=0 
M3956 n_AxB_4 n_AxB_4 Vdd GND dfet w=846 l=1598
+ ad=1.0559e+07 pd=32148 as=0 ps=0 
M3957 GND C34 _AxB_4_nC34 GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M3958 C45 C45 Vdd GND dfet w=846 l=846
+ ad=1.0453e+07 pd=38164 as=0 ps=0 
M3959 Vdd n_647 n_647 GND dfet w=752 l=1598
+ ad=0 pd=0 as=1.92536e+07 ps=65800 
M3960 Vdd A_B5 A_B5 GND dfet w=846 l=1504
+ ad=0 pd=0 as=7.86404e+06 ps=23876 
M3961 n_647 nA_B5 GND GND efet w=1692 l=658
+ ad=6.60933e+06 pd=18424 as=0 ps=0 
M3962 Vdd _AxB_4_nC34 _AxB_4_nC34 GND dfet w=846 l=1504
+ ad=0 pd=0 as=8.05843e+06 ps=26320 
M3963 Vdd nC45 nC45 GND dfet w=940 l=1598
+ ad=0 pd=0 as=2.01549e+07 ps=66552 
M3964 n_1218 n_1218 Vdd GND dfet w=846 l=1598
+ ad=1.03735e+07 pd=32336 as=0 ps=0 
M3965 Vdd alucout alucout GND dfet w=1034 l=658
+ ad=0 pd=0 as=6.22673e+07 ps=227480 
M3966 Vdd n_757 n_757 GND dfet w=846 l=1504
+ ad=0 pd=0 as=2.46966e+07 ps=92684 
M3967 n_939 n_647 GND GND efet w=4982 l=564
+ ad=3.27816e+06 pd=11280 as=0 ps=0 
M3968 n_757 DA_C45 n_939 GND efet w=4982 l=564
+ ad=5.9643e+06 pd=16544 as=0 ps=0 
M3969 nC45 C45 GND GND efet w=1692 l=564
+ ad=2.64196e+06 pd=9212 as=0 ps=0 
M3970 GND n_A_B_5 A_B5 GND efet w=2209 l=705
+ ad=0 pd=0 as=4.99234e+06 ps=15980 
M3971 n_165 A_B5 GND GND efet w=5170 l=564
+ ad=2.88937e+06 pd=11468 as=0 ps=0 
M3972 nC56 C45 n_165 GND efet w=5170 l=564
+ ad=6.90975e+06 pd=21244 as=0 ps=0 
M3973 n_AxB_5 dpc16_EORS naluresult5 GND efet w=1034 l=658
+ ad=4.02922e+06 pd=13160 as=0 ps=0 
M3974 GND AxB5 n_AxB_5 GND efet w=2726 l=658
+ ad=0 pd=0 as=0 ps=0 
M3975 AxB5 n_647 GND GND efet w=1692 l=564
+ ad=5.11604e+06 pd=15416 as=0 ps=0 
M3976 GND n_A_B_5 AxB5 GND efet w=1692 l=752
+ ad=0 pd=0 as=0 ps=0 
M3977 GND n_647 nC56 GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M3978 n_547 AxB5 GND GND efet w=3290 l=564
+ ad=1.85556e+06 pd=7708 as=0 ps=0 
M3979 n_AxBxC_5 nC45 n_547 GND efet w=3290 l=564
+ ad=7.74034e+06 pd=19740 as=0 ps=0 
M3980 Vdd n_AxBxC_5 n_AxBxC_5 GND dfet w=846 l=1692
+ ad=0 pd=0 as=4.22361e+06 ps=10528 
M3981 n_1257 n_1218 GND GND efet w=3290 l=658
+ ad=9.91399e+06 pd=25192 as=0 ps=0 
M3982 alucout notalucout GND GND efet w=7144 l=564
+ ad=8.56208e+06 pd=24628 as=0 ps=0 
M3983 n_1257 notalucout GND GND efet w=3572 l=658
+ ad=0 pd=0 as=0 ps=0 
M3984 n_1257 n_1257 Vdd GND dfet w=940 l=940
+ ad=3.34354e+07 pd=132540 as=0 ps=0 
M3985 n_AxBxC_5 n_AxB5__C45 GND GND efet w=2444 l=564
+ ad=0 pd=0 as=0 ps=0 
M3986 naluresult5 dpc17_SUMS n_AxBxC_5 GND efet w=1128 l=752
+ ad=0 pd=0 as=0 ps=0 
M3987 n_AxB5__C45 AxB5 GND GND efet w=1692 l=564
+ ad=4.69192e+06 pd=15416 as=0 ps=0 
M3988 n_AxB_5 n_AxB_5 Vdd GND dfet w=846 l=1598
+ ad=3.84366e+06 pd=11468 as=0 ps=0 
M3989 AxB5 AxB5 Vdd GND dfet w=940 l=1504
+ ad=2.02433e+07 pd=66928 as=0 ps=0 
M3990 GND nC45 n_AxB5__C45 GND efet w=3384 l=658
+ ad=0 pd=0 as=0 ps=0 
M3991 Vdd nC56 nC56 GND dfet w=846 l=940
+ ad=0 pd=0 as=1.30684e+07 ps=45120 
M3992 n_570 AxB5 GND GND efet w=2444 l=564
+ ad=9.74611e+06 pd=28764 as=0 ps=0 
M3993 GND n_647 n_570 GND efet w=2444 l=564
+ ad=0 pd=0 as=0 ps=0 
M3994 n_570 DA_C45 GND GND efet w=2444 l=658
+ ad=0 pd=0 as=0 ps=0 
M3995 GND n_122 n_570 GND efet w=2444 l=564
+ ad=0 pd=0 as=0 ps=0 
M3996 A_B6 A_B6 Vdd GND dfet w=846 l=1504
+ ad=7.77568e+06 pd=23124 as=0 ps=0 
M3997 nA_B6 dpc14_SRS naluresult5 GND efet w=1034 l=658
+ ad=0 pd=0 as=0 ps=0 
M3998 naluresult6 dpc13_ORS n_A_B_6 GND efet w=1128 l=658
+ ad=1.51714e+07 pd=42300 as=8.50023e+06 ps=26132 
M3999 GND dpc12_0ADD alua6 GND efet w=1269 l=705
+ ad=0 pd=0 as=4.7626e+06 ps=12784 
M4000 alua6 dpc11_SBADD sb6 GND efet w=1128 l=752
+ ad=0 pd=0 as=0 ps=0 
M4001 adl7 dpc10_ADLADD alub7 GND efet w=940 l=752
+ ad=0 pd=0 as=5.38996e+06 ps=13912 
M4002 alub7 dpc8_nDBADD n_423 GND efet w=1128 l=752
+ ad=0 pd=0 as=8.66812e+06 ps=25756 
M4003 alub7 dpc9_DBADD idb7 GND efet w=1128 l=658
+ ad=0 pd=0 as=1.85644e+07 ps=52640 
M4004 GND idb7 n_423 GND efet w=5640 l=658
+ ad=0 pd=0 as=0 ps=0 
M4005 n_423 n_423 Vdd GND dfet w=752 l=1598
+ ad=3.11027e+06 pd=8084 as=0 ps=0 
M4006 n_A_B_6 alua6 GND GND efet w=2820 l=564
+ ad=0 pd=0 as=0 ps=0 
M4007 GND alub6 n_A_B_6 GND efet w=2820 l=658
+ ad=0 pd=0 as=0 ps=0 
M4008 Vdd n_A_B_6 n_A_B_6 GND dfet w=940 l=2068
+ ad=0 pd=0 as=1.45175e+07 ps=48504 
M4009 n_1695 alua7 GND GND efet w=5734 l=564
+ ad=3.23398e+06 pd=12596 as=0 ps=0 
M4010 nA_B7 alub7 n_1695 GND efet w=5734 l=658
+ ad=1.26443e+07 pd=37036 as=0 ps=0 
M4011 Vdd nA_B7 nA_B7 GND dfet w=940 l=1974
+ ad=0 pd=0 as=1.50919e+07 ps=49444 
M4012 A_B6 n_A_B_6 GND GND efet w=1692 l=564
+ ad=4.5417e+06 pd=15228 as=0 ps=0 
M4013 n_AxB5__C45 n_AxB5__C45 Vdd GND dfet w=940 l=1692
+ ad=6.90092e+06 pd=21432 as=0 ps=0 
M4014 n_570 n_570 Vdd GND dfet w=940 l=1222
+ ad=2.20016e+07 pd=75764 as=0 ps=0 
M4015 GND nA_B6 n_1038 GND efet w=3384 l=564
+ ad=0 pd=0 as=3.46371e+06 ps=12220 
M4016 Vdd C56 C56 GND dfet w=846 l=1504
+ ad=0 pd=0 as=1.01172e+07 ps=31020 
M4017 C56 nC56 GND GND efet w=1692 l=564
+ ad=3.4107e+06 pd=11844 as=0 ps=0 
M4018 naluresult6 dpc15_ANDS nA_B6 GND efet w=1128 l=658
+ ad=0 pd=0 as=0 ps=0 
M4019 n_AxB_6 dpc16_EORS naluresult6 GND efet w=1128 l=658
+ ad=7.31621e+06 pd=23688 as=0 ps=0 
M4020 n_482 nA_B6 n_AxB_6 GND efet w=3196 l=564
+ ad=1.80254e+06 pd=7520 as=0 ps=0 
M4021 GND A_B6 n_482 GND efet w=3196 l=658
+ ad=0 pd=0 as=0 ps=0 
M4022 C67 n_A_B_6 GND GND efet w=2632 l=564
+ ad=7.40457e+06 pd=20680 as=0 ps=0 
M4023 n_112 nC56 C67 GND efet w=5123 l=611
+ ad=2.89821e+06 pd=11280 as=0 ps=0 
M4024 GND nA_B6 n_112 GND efet w=4982 l=564
+ ad=0 pd=0 as=0 ps=0 
M4025 n_1390 n_AxB_6 GND GND efet w=3290 l=658
+ ad=1.5463e+06 pd=7520 as=0 ps=0 
M4026 n_AxBxC_6 C56 n_1390 GND efet w=3290 l=658
+ ad=7.43108e+06 pd=20492 as=0 ps=0 
M4027 Vdd n_AxBxC_6 n_AxBxC_6 GND dfet w=940 l=1598
+ ad=0 pd=0 as=4.04689e+06 ps=9964 
M4028 n_1038 n_1038 Vdd GND dfet w=940 l=1410
+ ad=7.25436e+06 pd=29328 as=0 ps=0 
M4029 naluresult6 dpc17_SUMS n_AxBxC_6 GND efet w=1034 l=658
+ ad=0 pd=0 as=0 ps=0 
M4030 n_AxBxC_6 _AxB_6_nC56 GND GND efet w=2726 l=564
+ ad=0 pd=0 as=0 ps=0 
M4031 _AxB_6_nC56 n_AxB_6 GND GND efet w=1598 l=658
+ ad=4.77144e+06 pd=16732 as=0 ps=0 
M4032 nA_B7 dpc14_SRS naluresult6 GND efet w=1034 l=658
+ ad=0 pd=0 as=0 ps=0 
M4033 naluresult7 dpc13_ORS n_A_B_7 GND efet w=1128 l=658
+ ad=1.14603e+07 pd=30644 as=8.7123e+06 ps=26320 
M4034 GND dpc12_0ADD alua7 GND efet w=1128 l=658
+ ad=0 pd=0 as=4.72726e+06 ps=13160 
M4035 alua7 dpc11_SBADD sb7 GND efet w=1034 l=846
+ ad=0 pd=0 as=0 ps=0 
M4036 n_A_B_7 alua7 GND GND efet w=2914 l=564
+ ad=0 pd=0 as=0 ps=0 
M4037 GND alub7 n_A_B_7 GND efet w=2914 l=564
+ ad=0 pd=0 as=0 ps=0 
M4038 naluresult7 dpc14_SRS Vdd GND efet w=1128 l=752
+ ad=0 pd=0 as=0 ps=0 
M4039 naluresult7 dpc15_ANDS nA_B7 GND efet w=940 l=658
+ ad=0 pd=0 as=0 ps=0 
M4040 n_AxB_6 n_AxB_6 Vdd GND dfet w=846 l=940
+ ad=1.66912e+07 pd=56212 as=0 ps=0 
M4041 C67 C67 Vdd GND dfet w=940 l=940
+ ad=2.76744e+07 pd=94376 as=0 ps=0 
M4042 GND C56 _AxB_6_nC56 GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M4043 Vdd n_748 n_748 GND dfet w=846 l=1598
+ ad=0 pd=0 as=8.80066e+06 ps=29328 
M4044 Vdd A_B7 A_B7 GND dfet w=846 l=1598
+ ad=0 pd=0 as=7.91706e+06 ps=24816 
M4045 n_748 nA_B7 GND GND efet w=1786 l=564
+ ad=6.23822e+06 pd=18048 as=0 ps=0 
M4046 Vdd n_122 n_122 GND dfet w=846 l=1504
+ ad=0 pd=0 as=1.08064e+07 ps=36660 
M4047 n_122 n_AxB_6 GND GND efet w=3337 l=611
+ ad=5.02768e+06 pd=17108 as=0 ps=0 
M4048 n_269 AxB7 GND GND efet w=2444 l=658
+ ad=5.14255e+06 pd=14664 as=0 ps=0 
M4049 GND n_1038 n_269 GND efet w=2444 l=564
+ ad=0 pd=0 as=0 ps=0 
M4050 Vdd _AxB_6_nC56 _AxB_6_nC56 GND dfet w=846 l=1504
+ ad=0 pd=0 as=7.88171e+06 ps=25944 
M4051 Vdd nC67 nC67 GND dfet w=846 l=1598
+ ad=0 pd=0 as=1.00642e+07 ps=31584 
M4052 nC67 C67 GND GND efet w=1692 l=564
+ ad=2.47408e+06 pd=9024 as=0 ps=0 
M4053 n_1030 n_757 GND GND efet w=4794 l=564
+ ad=1.62494e+07 pd=39480 as=0 ps=0 
M4054 n_269 n_269 Vdd GND dfet w=940 l=1598
+ ad=1.04972e+07 pd=34592 as=0 ps=0 
M4055 GND n_AxB_6 n_1030 GND efet w=4888 l=564
+ ad=0 pd=0 as=0 ps=0 
M4056 GND n_A_B_7 A_B7 GND efet w=2162 l=658
+ ad=0 pd=0 as=5.35462e+06 ps=18424 
M4057 n_1617 A_B7 GND GND efet w=5217 l=611
+ ad=2.60662e+06 pd=11468 as=0 ps=0 
M4058 nC78 C67 n_1617 GND efet w=5217 l=611
+ ad=7.05996e+06 pd=21244 as=0 ps=0 
M4059 n_AxB_7 dpc16_EORS naluresult7 GND efet w=1034 l=658
+ ad=4.14408e+06 pd=12596 as=0 ps=0 
M4060 Vdd n_A_B_7 n_A_B_7 GND dfet w=846 l=2068
+ ad=0 pd=0 as=2.52533e+07 ps=78020 
M4061 dpc0_YSB cclk GND GND efet w=2538 l=752
+ ad=0 pd=0 as=0 ps=0 
M4062 dpc1_SBY cclk GND GND efet w=2632 l=752
+ ad=0 pd=0 as=0 ps=0 
M4063 dpc2_XSB cclk GND GND efet w=2350 l=752
+ ad=0 pd=0 as=0 ps=0 
M4064 dpc3_SBX cclk GND GND efet w=2538 l=752
+ ad=0 pd=0 as=0 ps=0 
M4065 GND AxB7 n_AxB_7 GND efet w=2726 l=658
+ ad=0 pd=0 as=0 ps=0 
M4066 AxB7 n_748 GND GND efet w=2256 l=658
+ ad=4.97467e+06 pd=15980 as=0 ps=0 
M4067 GND n_A_B_7 AxB7 GND efet w=1598 l=658
+ ad=0 pd=0 as=0 ps=0 
M4068 GND n_748 nC78 GND efet w=2444 l=564
+ ad=0 pd=0 as=0 ps=0 
M4069 n_1013 AxB7 GND GND efet w=3290 l=658
+ ad=1.5463e+06 pd=7520 as=0 ps=0 
M4070 n_AxBxC_7 nC67 n_1013 GND efet w=3290 l=658
+ ad=7.65198e+06 pd=20492 as=0 ps=0 
M4071 Vdd n_AxBxC_7 n_AxBxC_7 GND dfet w=846 l=1504
+ ad=0 pd=0 as=3.8525e+06 ps=9776 
M4072 n_1030 n_269 DC78 GND efet w=5687 l=611
+ ad=0 pd=0 as=1.18667e+07 ps=38728 
M4073 n_1030 n_570 DC78 GND efet w=5546 l=658
+ ad=0 pd=0 as=0 ps=0 
M4074 n_AxBxC_7 n_AxB7__C67 GND GND efet w=2820 l=564
+ ad=0 pd=0 as=0 ps=0 
M4075 naluresult7 dpc17_SUMS n_AxBxC_7 GND efet w=1034 l=752
+ ad=0 pd=0 as=0 ps=0 
M4076 n_AxB_7 n_AxB_7 Vdd GND dfet w=940 l=1598
+ ad=3.91435e+06 pd=11280 as=0 ps=0 
M4077 AxB7 AxB7 Vdd GND dfet w=846 l=1504
+ ad=2.69321e+07 pd=92120 as=0 ps=0 
M4078 n_AxB7__C67 AxB7 GND GND efet w=1692 l=658
+ ad=4.37382e+06 pd=15228 as=0 ps=0 
M4079 GND nC67 n_AxB7__C67 GND efet w=3243 l=705
+ ad=0 pd=0 as=0 ps=0 
M4080 alu1 alu1 Vdd GND dfet w=846 l=1128
+ ad=7.89055e+06 pd=25568 as=0 ps=0 
M4081 dpc24_ACSB n_1247 GND GND efet w=6862 l=470
+ ad=0 pd=0 as=0 ps=0 
M4082 GND n_1335 dpc24_ACSB GND efet w=7144 l=564
+ ad=0 pd=0 as=0 ps=0 
M4083 dpc26_ACDB n_800 GND GND efet w=7144 l=564
+ ad=0 pd=0 as=0 ps=0 
M4084 n_849 n_321 GND GND efet w=2350 l=658
+ ad=3.20747e+06 pd=9964 as=0 ps=0 
M4085 Vdd n_255 n_255 GND dfet w=893 l=1457
+ ad=0 pd=0 as=1.06297e+07 ps=33276 
M4086 n_1323 n_631 GND GND efet w=2350 l=564
+ ad=3.07493e+06 pd=9964 as=0 ps=0 
M4087 Vdd n_611 dpc31_PCHPCH GND dfet w=940 l=1034
+ ad=0 pd=0 as=1.67e+07 ps=37224 
M4088 n_849 n_849 Vdd GND dfet w=846 l=1410
+ ad=1.10715e+07 pd=33652 as=0 ps=0 
M4089 n_1413 n_1260 GND GND efet w=2256 l=658
+ ad=3.12794e+06 pd=9964 as=0 ps=0 
M4090 n_1518 n_1270 GND GND efet w=2350 l=564
+ ad=3.13678e+06 pd=9776 as=0 ps=0 
M4091 n_818 n_265 GND GND efet w=5123 l=611
+ ad=7.74034e+06 pd=20680 as=0 ps=0 
M4092 Vdd n_818 n_818 GND dfet w=940 l=1316
+ ad=0 pd=0 as=1.01879e+07 ps=32336 
M4093 n_1480 n_1581 dpc36_nIPC GND efet w=14476 l=564
+ ad=0 pd=0 as=0 ps=0 
M4094 pipeUNK17 cclk n_334 GND efet w=1128 l=846
+ ad=2.05879e+06 pd=7332 as=0 ps=0 
M4095 nop_set_C cclk pipeUNK08 GND efet w=1128 l=846
+ ad=0 pd=0 as=1.50212e+06 ps=7144 
M4096 n_513 n_885 GND GND efet w=4935 l=611
+ ad=0 pd=0 as=0 ps=0 
M4097 Vdd n_513 n_513 GND dfet w=940 l=752
+ ad=0 pd=0 as=1.79371e+06 ps=6768 
M4098 n_553 n_1662 GND GND efet w=2820 l=658
+ ad=1.02056e+07 pd=28388 as=0 ps=0 
M4099 n_553 n_781 GND GND efet w=3854 l=658
+ ad=0 pd=0 as=0 ps=0 
M4100 n_954 n_954 Vdd GND dfet w=1034 l=1128
+ ad=3.70493e+07 pd=131600 as=0 ps=0 
M4101 GND n_954 n_513 GND efet w=3854 l=658
+ ad=0 pd=0 as=0 ps=0 
M4102 GND pipeUNK08 n_954 GND efet w=7849 l=611
+ ad=0 pd=0 as=9.50754e+06 ps=25380 
M4103 n_1379 cclk pipeUNK07 GND efet w=1034 l=846
+ ad=0 pd=0 as=1.05148e+06 ps=5640 
M4104 Vdd n_1379 n_1379 GND dfet w=940 l=1692
+ ad=0 pd=0 as=3.9762e+06 ps=9588 
M4105 n_327 cclk pipeUNK09 GND efet w=1410 l=752
+ ad=0 pd=0 as=1.41376e+06 ps=7332 
M4106 GND pipeUNK09 n_941 GND efet w=5875 l=611
+ ad=0 pd=0 as=4.31197e+06 ps=16168 
M4107 pipeUNK11 cclk n_862 GND efet w=1128 l=658
+ ad=1.44027e+06 pd=7144 as=0 ps=0 
M4108 Vdd fetch fetch GND dfet w=846 l=940
+ ad=0 pd=0 as=8.31468e+07 ps=263388 
M4109 n_941 pipeUNK07 n_1111 GND efet w=7191 l=611
+ ad=0 pd=0 as=9.60473e+06 ps=23500 
M4110 Vdd n_774 n_774 GND dfet w=940 l=1692
+ ad=0 pd=0 as=1.65763e+07 ps=58092 
M4111 n_513 cclk pipeUNK06 GND efet w=1128 l=752
+ ad=0 pd=0 as=1.67e+06 ps=7708 
M4112 n_754 n_754 Vdd GND dfet w=940 l=1786
+ ad=4.10609e+07 pd=137616 as=0 ps=0 
M4113 n_1225 cclk n_1121 GND efet w=1128 l=940
+ ad=0 pd=0 as=1.27238e+06 ps=6204 
M4114 n_1705 cclk n_1020 GND efet w=1128 l=940
+ ad=0 pd=0 as=1.99694e+06 ps=7520 
M4115 n_104 cclk n_1221 GND efet w=1128 l=846
+ ad=0 pd=0 as=1.99694e+06 ps=7520 
M4116 n_754 n_1673 GND GND efet w=3760 l=658
+ ad=1.12217e+07 pd=25568 as=0 ps=0 
M4117 n_1422 pipeUNK06 n_754 GND efet w=7238 l=470
+ ad=4.58588e+06 pd=17860 as=0 ps=0 
M4118 GND pipeUNK09 n_1422 GND efet w=8460 l=658
+ ad=0 pd=0 as=0 ps=0 
M4119 n_781 pipeUNK09 GND GND efet w=7285 l=611
+ ad=0 pd=0 as=0 ps=0 
M4120 Vdd n_781 n_781 GND dfet w=940 l=940
+ ad=0 pd=0 as=5.58435e+07 ps=196648 
M4121 n_1111 n_1111 Vdd GND dfet w=940 l=2162
+ ad=3.40009e+07 pd=104904 as=0 ps=0 
M4122 nnT2BR cclk n_1269 GND efet w=1222 l=752
+ ad=0 pd=0 as=1.58164e+06 ps=6956 
M4123 Vdd n_1401 n_1401 GND dfet w=940 l=1692
+ ad=0 pd=0 as=7.3869e+06 ps=24816 
M4124 fetch n_1214 GND GND efet w=3572 l=658
+ ad=0 pd=0 as=0 ps=0 
M4125 GND pipeUNK11 n_1214 GND efet w=4136 l=658
+ ad=0 pd=0 as=5.12488e+06 ps=14100 
M4126 Vdd n_1214 n_1214 GND dfet w=1081 l=1457
+ ad=0 pd=0 as=8.05843e+06 ps=26696 
M4127 pd3_clearIR clearIR GND GND efet w=2820 l=658
+ ad=0 pd=0 as=0 ps=0 
M4128 pd4_clearIR pd4 GND GND efet w=7050 l=658
+ ad=0 pd=0 as=0 ps=0 
M4129 GND clearIR pd5_clearIR GND efet w=2820 l=658
+ ad=0 pd=0 as=0 ps=0 
M4130 pd0_clearIR clearIR GND GND efet w=2820 l=564
+ ad=0 pd=0 as=0 ps=0 
M4131 GND clearIR pd1_clearIR GND efet w=2914 l=658
+ ad=0 pd=0 as=0 ps=0 
M4132 pd7_clearIR clearIR GND GND efet w=3854 l=564
+ ad=9.33965e+06 pd=28200 as=0 ps=0 
M4133 pd3_clearIR pd3_clearIR Vdd GND dfet w=940 l=940
+ ad=1.76985e+07 pd=60912 as=0 ps=0 
M4134 Vdd pd4_clearIR pd4_clearIR GND dfet w=940 l=1034
+ ad=0 pd=0 as=2.07911e+07 ps=71816 
M4135 GND pd7 pd7_clearIR GND efet w=8460 l=658
+ ad=0 pd=0 as=0 ps=0 
M4136 pd2_clearIR pd2 GND GND efet w=9494 l=658
+ ad=8.99505e+06 pd=27824 as=0 ps=0 
M4137 GND clearIR pd2_clearIR GND efet w=2914 l=564
+ ad=0 pd=0 as=0 ps=0 
M4138 pd6_clearIR clearIR GND GND efet w=2914 l=658
+ ad=8.91552e+06 pd=27448 as=0 ps=0 
M4139 GND pd6 pd6_clearIR GND efet w=8319 l=705
+ ad=0 pd=0 as=0 ps=0 
M4140 pd5_clearIR pd5_clearIR Vdd GND dfet w=940 l=1034
+ ad=2.22667e+07 pd=69372 as=0 ps=0 
M4141 pd0_clearIR pd0_clearIR Vdd GND dfet w=1034 l=846
+ ad=1.94834e+07 pd=70688 as=0 ps=0 
M4142 pd1_clearIR pd1_clearIR Vdd GND dfet w=940 l=940
+ ad=2.05084e+07 pd=72380 as=0 ps=0 
M4143 pd7_clearIR pd7_clearIR Vdd GND dfet w=940 l=940
+ ad=2.06321e+07 pd=70876 as=0 ps=0 
M4144 pd2_clearIR pd2_clearIR Vdd GND dfet w=940 l=940
+ ad=1.97661e+07 pd=70312 as=0 ps=0 
M4145 pd6_clearIR pd6_clearIR Vdd GND dfet w=1034 l=940
+ ad=2.87789e+07 pd=100204 as=0 ps=0 
M4146 pd4 cclk n_1075 GND efet w=1410 l=658
+ ad=1.99694e+06 pd=8272 as=1.27769e+07 ps=33464 
M4147 pd3 cclk n_1281 GND efet w=1504 l=846
+ ad=1.57281e+06 pd=7144 as=1.2821e+07 ps=32712 
M4148 pd5 cclk n_1588 GND efet w=1410 l=846
+ ad=1.36074e+06 pd=5828 as=1.37842e+07 ps=34216 
M4149 pd0 cclk n_93 GND efet w=1504 l=846
+ ad=1.5463e+06 pd=7332 as=1.37577e+07 ps=33840 
M4150 pd1 cclk n_1319 GND efet w=1316 l=846
+ ad=1.27238e+06 pd=5640 as=1.30419e+07 ps=32524 
M4151 pd7 cclk n_62 GND efet w=1410 l=846
+ ad=1.4491e+06 pd=6956 as=1.24941e+07 ps=33464 
M4152 pd2 cclk n_111 GND efet w=1410 l=846
+ ad=1.34307e+06 pd=5828 as=1.28741e+07 ps=31960 
M4153 pd6 cclk n_374 GND efet w=1410 l=846
+ ad=1.93508e+06 pd=7332 as=1.2715e+07 ps=35532 
M4154 GND op_clv n_340 GND efet w=4277 l=611
+ ad=0 pd=0 as=5.07186e+06 ps=14100 
M4155 n_503 notir5 GND GND efet w=3431 l=611
+ ad=4.1971e+06 pd=11280 as=0 ps=0 
M4156 n_340 n_340 Vdd GND dfet w=940 l=1504
+ ad=3.94969e+06 pd=10904 as=0 ps=0 
M4157 Vdd n_587 n_587 GND dfet w=940 l=1692
+ ad=0 pd=0 as=3.09879e+07 ps=111860 
M4158 n_340 cclk pipeUNK12 GND efet w=1128 l=752
+ ad=0 pd=0 as=1.25471e+06 ps=5828 
M4159 n_1673 cclk op_T__bit GND efet w=1128 l=752
+ ad=1.31656e+06 pd=5640 as=0 ps=0 
M4160 n_160 op_SRS GND GND efet w=3102 l=564
+ ad=9.31314e+06 pd=26508 as=0 ps=0 
M4161 GND n_781 n_160 GND efet w=2820 l=658
+ ad=0 pd=0 as=0 ps=0 
M4162 n_1049 cclk n_160 GND efet w=1222 l=752
+ ad=1.31656e+06 pd=6392 as=0 ps=0 
M4163 GND n_1049 n_507 GND efet w=5499 l=611
+ ad=0 pd=0 as=6.088e+06 ps=17672 
M4164 n_160 n_160 Vdd GND dfet w=940 l=1222
+ ad=2.8717e+06 pd=8836 as=0 ps=0 
M4165 n_507 n_507 Vdd GND dfet w=940 l=1410
+ ad=9.72844e+06 pd=31960 as=0 ps=0 
M4166 Vdd n_279 n_279 GND dfet w=846 l=1410
+ ad=0 pd=0 as=9.92283e+06 ps=33088 
M4167 n_279 n_253 GND GND efet w=3102 l=658
+ ad=9.55172e+06 pd=23688 as=0 ps=0 
M4168 n_279 n_954 GND GND efet w=2162 l=564
+ ad=0 pd=0 as=0 ps=0 
M4169 GND n_507 n_279 GND efet w=2256 l=564
+ ad=0 pd=0 as=0 ps=0 
M4170 n_1692 n_270 n_1082 GND efet w=3337 l=611
+ ad=1.70535e+06 pd=7708 as=2.18868e+07 ps=54332 
M4171 GND n_253 n_1692 GND efet w=3290 l=564
+ ad=0 pd=0 as=0 ps=0 
M4172 GND pipeUNK06 n_755 GND efet w=5734 l=658
+ ad=0 pd=0 as=6.95393e+06 ps=19176 
M4173 n_1401 n_1269 GND GND efet w=5264 l=564
+ ad=6.61816e+06 pd=19364 as=0 ps=0 
M4174 n_1249 n_1269 GND GND efet w=8460 l=658
+ ad=6.60049e+06 pd=15792 as=0 ps=0 
M4175 n_755 n_755 Vdd GND dfet w=940 l=1692
+ ad=3.87812e+07 pd=139872 as=0 ps=0 
M4176 Vdd n_771 n_771 GND dfet w=940 l=1316
+ ad=0 pd=0 as=2.23639e+07 ps=75012 
M4177 GND pipeUNK01 n_1198 GND efet w=5875 l=611
+ ad=0 pd=0 as=5.31044e+06 ps=15604 
M4178 Vdd n_503 n_503 GND dfet w=940 l=1504
+ ad=0 pd=0 as=6.64467e+06 ps=19176 
M4179 GND pipeUNK12 n_587 GND efet w=4982 l=564
+ ad=0 pd=0 as=6.8479e+06 ps=19176 
M4180 n_1198 n_1401 n_626 GND efet w=3384 l=564
+ ad=0 pd=0 as=9.39267e+06 ps=23500 
M4181 n_626 DBNeg n_1249 GND efet w=4230 l=658
+ ad=0 pd=0 as=0 ps=0 
M4182 Vdd n_1110 n_1110 GND dfet w=940 l=940
+ ad=0 pd=0 as=1.05944e+07 ps=36472 
M4183 n_626 n_626 Vdd GND dfet w=846 l=1786
+ ad=3.87017e+06 pd=10716 as=0 ps=0 
M4184 pipeUNK01 cclk n_1110 GND efet w=1128 l=846
+ ad=1.27238e+06 pd=5264 as=1.46678e+07 ps=37412 
M4185 GND n_756 n_1110 GND efet w=12596 l=658
+ ad=0 pd=0 as=0 ps=0 
M4186 n_626 cp1 n_756 GND efet w=1034 l=752
+ ad=0 pd=0 as=1.94392e+06 ps=8084 
M4187 GND n_1110 n_771 GND efet w=3290 l=752
+ ad=0 pd=0 as=6.39726e+06 ps=18612 
M4188 n_367 n_954 GND GND efet w=3337 l=611
+ ad=2.96006e+06 pd=10716 as=0 ps=0 
M4189 n_1082 n_206 n_367 GND efet w=3478 l=564
+ ad=0 pd=0 as=0 ps=0 
M4190 n_186 n_507 n_1082 GND efet w=2914 l=658
+ ad=1.36958e+06 pd=6768 as=0 ps=0 
M4191 GND n_1224 n_186 GND efet w=2914 l=658
+ ad=0 pd=0 as=0 ps=0 
M4192 Vdd n_132 n_132 GND dfet w=846 l=846
+ ad=0 pd=0 as=5.48981e+07 ps=205672 
M4193 GND n_31 n_132 GND efet w=4324 l=564
+ ad=0 pd=0 as=0 ps=0 
M4194 GND n_43 n_818 GND efet w=2256 l=564
+ ad=0 pd=0 as=0 ps=0 
M4195 Vdd n_291 n_291 GND dfet w=846 l=1034
+ ad=0 pd=0 as=1.16105e+07 ps=36848 
M4196 GND n_1121 n_291 GND efet w=7379 l=611
+ ad=0 pd=0 as=7.45758e+06 ps=18800 
M4197 n_1277 n_1020 GND GND efet w=6768 l=564
+ ad=6.92742e+06 pd=19364 as=0 ps=0 
M4198 Vdd n_1277 n_1277 GND dfet w=940 l=1034
+ ad=0 pd=0 as=1.02409e+07 ps=35908 
M4199 Vdd n_321 dpc33_PCHDB GND dfet w=752 l=846
+ ad=0 pd=0 as=1.04883e+07 ps=26132 
M4200 n_1323 n_1323 Vdd GND dfet w=846 l=1316
+ ad=1.04176e+07 pd=34028 as=0 ps=0 
M4201 GND n_1247 dpc26_ACDB GND efet w=7050 l=564
+ ad=0 pd=0 as=0 ps=0 
M4202 dpc30_ADHPCH n_1247 GND GND efet w=7238 l=752
+ ad=0 pd=0 as=0 ps=0 
M4203 GND n_228 dpc30_ADHPCH GND efet w=7379 l=705
+ ad=0 pd=0 as=0 ps=0 
M4204 dpc31_PCHPCH n_1247 GND GND efet w=7144 l=752
+ ad=0 pd=0 as=0 ps=0 
M4205 GND n_255 dpc31_PCHPCH GND efet w=7097 l=611
+ ad=0 pd=0 as=0 ps=0 
M4206 GND n_849 dpc33_PCHDB GND efet w=9118 l=658
+ ad=0 pd=0 as=0 ps=0 
M4207 Vdd n_631 dpc37_PCLDB GND dfet w=752 l=846
+ ad=0 pd=0 as=1.0886e+07 ps=25756 
M4208 n_1413 n_1413 Vdd GND dfet w=940 l=1410
+ ad=1.12836e+07 pd=33840 as=0 ps=0 
M4209 n_1462 n_1369 GND GND efet w=2350 l=564
+ ad=3.2163e+06 pd=9964 as=0 ps=0 
M4210 n_1518 n_1518 Vdd GND dfet w=940 l=1316
+ ad=1.16989e+07 pd=37224 as=0 ps=0 
M4211 n_1043 n_818 GND GND efet w=2444 l=564
+ ad=3.74646e+06 pd=10340 as=0 ps=0 
M4212 GND dpc34_PCLC n_1007 GND efet w=2068 l=564
+ ad=0 pd=0 as=3.16329e+06 ps=10716 
M4213 GND n_1323 dpc37_PCLDB GND efet w=8977 l=611
+ ad=0 pd=0 as=0 ps=0 
M4214 Vdd n_1260 dpc32_PCHADH GND dfet w=940 l=846
+ ad=0 pd=0 as=1.1098e+07 ps=28576 
M4215 GND n_1413 dpc32_PCHADH GND efet w=9212 l=658
+ ad=0 pd=0 as=0 ps=0 
M4216 Vdd n_1270 dpc39_PCLPCL GND dfet w=846 l=940
+ ad=0 pd=0 as=1.69209e+07 ps=32524 
M4217 n_1462 n_1462 Vdd GND dfet w=940 l=1316
+ ad=1.11687e+07 pd=34592 as=0 ps=0 
M4218 n_1043 n_1043 Vdd GND dfet w=940 l=1316
+ ad=1.08506e+07 pd=33088 as=0 ps=0 
M4219 Vdd n_1369 dpc38_PCLADL GND dfet w=940 l=940
+ ad=0 pd=0 as=1.05148e+07 ps=24064 
M4220 GND n_1462 dpc38_PCLADL GND efet w=9306 l=658
+ ad=0 pd=0 as=0 ps=0 
M4221 dpc39_PCLPCL n_1247 GND GND efet w=7943 l=611
+ ad=0 pd=0 as=0 ps=0 
M4222 adl2 dpc21_ADDADL alu2 GND efet w=1410 l=752
+ ad=0 pd=0 as=1.38107e+07 ps=39668 
M4223 naluresult2 cclk notalu2 GND efet w=1034 l=752
+ ad=0 pd=0 as=1.6435e+06 ps=6956 
M4224 GND notalu2 alu2 GND efet w=9494 l=564
+ ad=0 pd=0 as=0 ps=0 
M4225 alu2 dpc20_ADDSB06 sb2 GND efet w=1974 l=752
+ ad=0 pd=0 as=0 ps=0 
M4226 alu2 alu2 Vdd GND dfet w=846 l=1128
+ ad=1.13719e+07 pd=37600 as=0 ps=0 
M4227 adl3 dpc21_ADDADL alu3 GND efet w=1504 l=752
+ ad=0 pd=0 as=1.34926e+07 ps=39668 
M4228 naluresult3 cclk notalu3 GND efet w=1034 l=752
+ ad=0 pd=0 as=1.67884e+06 ps=6956 
M4229 GND notalu3 alu3 GND efet w=9447 l=611
+ ad=0 pd=0 as=0 ps=0 
M4230 alu3 dpc20_ADDSB06 sb3 GND efet w=1974 l=752
+ ad=0 pd=0 as=0 ps=0 
M4231 alu3 alu3 Vdd GND dfet w=940 l=1128
+ ad=3.16329e+06 pd=9776 as=0 ps=0 
M4232 adl4 dpc21_ADDADL alu4 GND efet w=1504 l=658
+ ad=0 pd=0 as=1.41199e+07 ps=39480 
M4233 naluresult4 cclk notalu4 GND efet w=1128 l=846
+ ad=0 pd=0 as=1.53746e+06 ps=6956 
M4234 GND notalu4 alu4 GND efet w=9259 l=611
+ ad=0 pd=0 as=0 ps=0 
M4235 alu4 dpc20_ADDSB06 sb4 GND efet w=1974 l=752
+ ad=0 pd=0 as=0 ps=0 
M4236 alu4 alu4 Vdd GND dfet w=846 l=1128
+ ad=3.16329e+06 pd=9776 as=0 ps=0 
M4237 adl5 dpc21_ADDADL alu5 GND efet w=1504 l=752
+ ad=0 pd=0 as=1.40404e+07 ps=39668 
M4238 naluresult5 cclk notalu5 GND efet w=1128 l=846
+ ad=0 pd=0 as=1.53746e+06 ps=6956 
M4239 GND notalu5 alu5 GND efet w=9306 l=658
+ ad=0 pd=0 as=0 ps=0 
M4240 Vdd notalucout notalucout GND dfet w=846 l=1504
+ ad=0 pd=0 as=3.51143e+07 ps=120696 
M4241 DC78 dpc18_nDAA GND GND efet w=2538 l=564
+ ad=0 pd=0 as=0 ps=0 
M4242 Vdd nC78 nC78 GND dfet w=940 l=846
+ ad=0 pd=0 as=1.25471e+07 ps=48316 
M4243 n_1489 n_A_B_7 GND GND efet w=5217 l=705
+ ad=4.90398e+06 pd=16168 as=0 ps=0 
M4244 dpc6_SBS cclk GND GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M4245 dpc7_SS cclk GND GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M4246 dpc8_nDBADD cclk GND GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M4247 dpc9_DBADD cclk GND GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M4248 dpc10_ADLADD cclk GND GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M4249 dpc11_SBADD cclk GND GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M4250 dpc12_0ADD cclk GND GND efet w=2444 l=752
+ ad=0 pd=0 as=0 ps=0 
M4251 n_637 nA_B7 GND GND efet w=2256 l=564
+ ad=4.57705e+06 pd=15604 as=0 ps=0 
M4252 GND C67 n_637 GND efet w=2867 l=611
+ ad=0 pd=0 as=0 ps=0 
M4253 notaluvout C67 n_1489 GND efet w=4888 l=658
+ ad=9.35732e+06 pd=31020 as=0 ps=0 
M4254 DC78 DC78 Vdd GND dfet w=846 l=1034
+ ad=5.48716e+06 pd=18236 as=0 ps=0 
M4255 n_AxB7__C67 n_AxB7__C67 Vdd GND dfet w=987 l=1551
+ ad=6.63584e+06 pd=21432 as=0 ps=0 
M4256 Vdd C78 C78 GND dfet w=846 l=752
+ ad=0 pd=0 as=2.68614e+06 ps=9776 
M4257 notalucout DC78_phi2 GND GND efet w=3948 l=564
+ ad=9.48103e+06 pd=23124 as=0 ps=0 
M4258 GND C78_phi2 notalucout GND efet w=3948 l=564
+ ad=0 pd=0 as=0 ps=0 
M4259 alu5 dpc20_ADDSB06 sb5 GND efet w=1974 l=658
+ ad=0 pd=0 as=0 ps=0 
M4260 alu5 alu5 Vdd GND dfet w=846 l=1222
+ ad=7.66081e+06 pd=22748 as=0 ps=0 
M4261 adl6 dpc21_ADDADL alu6 GND efet w=1410 l=846
+ ad=0 pd=0 as=1.38107e+07 ps=39292 
M4262 naluresult6 cclk notalu6 GND efet w=1034 l=846
+ ad=0 pd=0 as=1.57281e+06 ps=7144 
M4263 GND notalu6 alu6 GND efet w=9353 l=611
+ ad=0 pd=0 as=0 ps=0 
M4264 alu6 dpc20_ADDSB06 sb6 GND efet w=1974 l=658
+ ad=0 pd=0 as=0 ps=0 
M4265 alu6 alu6 Vdd GND dfet w=846 l=1128
+ ad=7.54594e+06 pd=24628 as=0 ps=0 
M4266 notalu7 cclk naluresult7 GND efet w=1034 l=752
+ ad=1.90858e+06 pd=7332 as=0 ps=0 
M4267 n_1556 nDA_ADD1 GND GND efet w=3196 l=658
+ ad=1.9881e+06 pd=8084 as=0 ps=0 
M4268 n_986 nDA_ADD2 n_1556 GND efet w=3478 l=658
+ ad=4.23244e+06 pd=12408 as=0 ps=0 
M4269 Vdd n_986 n_986 GND dfet w=846 l=1598
+ ad=0 pd=0 as=3.20482e+07 ps=119756 
M4270 Vdd n_1682 n_1682 GND dfet w=846 l=1598
+ ad=0 pd=0 as=7.05113e+06 ps=21244 
M4271 n_36 n_36 Vdd GND dfet w=846 l=1598
+ ad=1.70093e+07 pd=61476 as=0 ps=0 
M4272 n_36 n_8 GND GND efet w=1786 l=658
+ ad=7.61663e+06 pd=23688 as=0 ps=0 
M4273 n_867 nDA_ADD1 GND GND efet w=2538 l=658
+ ad=6.59166e+06 pd=15980 as=0 ps=0 
M4274 GND nDA_ADD2 n_867 GND efet w=3196 l=658
+ ad=0 pd=0 as=0 ps=0 
M4275 n_867 n_867 Vdd GND dfet w=940 l=1598
+ ad=1.40227e+07 pd=45120 as=0 ps=0 
M4276 Vdd nDA_ADD1 nDA_ADD1 GND dfet w=1034 l=1504
+ ad=0 pd=0 as=1.78576e+07 ps=57716 
M4277 n_1682 nDA_ADD1 GND GND efet w=1692 l=658
+ ad=3.08376e+06 pd=11280 as=0 ps=0 
M4278 n_150 n_1682 n_613 GND efet w=3478 l=564
+ ad=3.4372e+06 pd=8836 as=1.1584e+07 ps=34968 
M4279 GND n_8 n_150 GND efet w=3290 l=658
+ ad=0 pd=0 as=0 ps=0 
M4280 n_36 n_600 GND GND efet w=1974 l=658
+ ad=0 pd=0 as=0 ps=0 
M4281 n_1362 nDA_ADD1 GND GND efet w=4982 l=564
+ ad=4.1971e+06 pd=13348 as=0 ps=0 
M4282 n_613 n_600 n_1362 GND efet w=7332 l=564
+ ad=0 pd=0 as=0 ps=0 
M4283 nDA_ADD1 alu1 GND GND efet w=4324 l=658
+ ad=4.99234e+06 pd=14852 as=0 ps=0 
M4284 nDA_ADD2 alu2 GND GND efet w=4183 l=611
+ ad=3.95853e+06 pd=13724 as=0 ps=0 
M4285 GND n_867 n_876 GND efet w=1692 l=564
+ ad=0 pd=0 as=3.94969e+06 ps=12972 
M4286 nDA_ADD2 nDA_ADD2 Vdd GND dfet w=940 l=1598
+ ad=1.96601e+07 pd=63168 as=0 ps=0 
M4287 n_876 n_876 Vdd GND dfet w=846 l=1504
+ ad=1.81757e+07 pd=64108 as=0 ps=0 
M4288 Vdd n_600 n_600 GND dfet w=846 l=940
+ ad=0 pd=0 as=3.45841e+07 ps=129156 
M4289 n_600 n_1341 GND GND efet w=7426 l=658
+ ad=8.21748e+06 pd=21432 as=0 ps=0 
M4290 Vdd n_146 n_146 GND dfet w=940 l=1128
+ ad=0 pd=0 as=3.12794e+06 ps=10152 
M4291 GND n_1518 dpc39_PCLPCL GND efet w=8554 l=564
+ ad=0 pd=0 as=0 ps=0 
M4292 Vdd n_818 dpc40_ADLPCL GND dfet w=846 l=1034
+ ad=0 pd=0 as=1.51802e+07 ps=29328 
M4293 n_1566 n_1221 GND GND efet w=6580 l=564
+ ad=7.07764e+06 pd=18988 as=0 ps=0 
M4294 Vdd n_1566 n_1566 GND dfet w=940 l=1034
+ ad=0 pd=0 as=9.97584e+06 ps=37412 
M4295 GND n_334 Pout2 GND efet w=6298 l=658
+ ad=0 pd=0 as=1.05855e+07 ps=29140 
M4296 p7 n_1045 GND GND efet w=6298 l=658
+ ad=1.0347e+07 pd=28200 as=0 ps=0 
M4297 Vdd Pout2 Pout2 GND dfet w=940 l=940
+ ad=0 pd=0 as=2.45641e+06 ps=8084 
M4298 p7 p7 Vdd GND dfet w=940 l=846
+ ad=2.3327e+06 pd=8084 as=0 ps=0 
M4299 Pout2 H1x1 idb2 GND efet w=2350 l=752
+ ad=0 pd=0 as=0 ps=0 
M4300 p7 H1x1 idb7 GND efet w=2256 l=752
+ ad=0 pd=0 as=0 ps=0 
M4301 n_1007 n_1007 Vdd GND dfet w=940 l=1598
+ ad=9.72844e+06 pd=30456 as=0 ps=0 
M4302 dpc40_ADLPCL n_1247 GND GND efet w=7050 l=658
+ ad=0 pd=0 as=0 ps=0 
M4303 GND n_1043 dpc40_ADLPCL GND efet w=7238 l=658
+ ad=0 pd=0 as=0 ps=0 
M4304 dpc35_PCHC n_1007 GND GND efet w=5170 l=564
+ ad=2.56244e+07 pd=75388 as=0 ps=0 
M4305 n_1157 n_291 GND GND efet w=2350 l=564
+ ad=3.11027e+06 pd=9588 as=0 ps=0 
M4306 n_1157 n_1157 Vdd GND dfet w=940 l=1316
+ ad=1.12217e+07 pd=34968 as=0 ps=0 
M4307 n_1441 n_1441 Vdd GND dfet w=940 l=1316
+ ad=1.19639e+07 pd=37224 as=0 ps=0 
M4308 GND n_1277 n_1441 GND efet w=2350 l=564
+ ad=0 pd=0 as=4.06456e+06 ps=10904 
M4309 GND n_1566 n_1240 GND efet w=2350 l=564
+ ad=0 pd=0 as=3.16329e+06 ps=9588 
M4310 GND idb2 n_1573 GND efet w=6768 l=564
+ ad=0 pd=0 as=7.21018e+06 ps=20680 
M4311 DBNeg idb7 GND GND efet w=7896 l=564
+ ad=6.60049e+06 pd=18236 as=0 ps=0 
M4312 Vdd n_291 dpc41_DL_ADL GND dfet w=846 l=846
+ ad=0 pd=0 as=1.06297e+07 ps=23688 
M4313 Vdd n_1277 dpc42_DL_ADH GND dfet w=940 l=846
+ ad=0 pd=0 as=9.87865e+06 ps=24628 
M4314 n_1240 n_1240 Vdd GND dfet w=846 l=1316
+ ad=1.17342e+07 pd=36472 as=0 ps=0 
M4315 n_1573 n_1573 Vdd GND dfet w=846 l=1128
+ ad=3.0926e+07 pd=115244 as=0 ps=0 
M4316 DBNeg DBNeg Vdd GND dfet w=940 l=752
+ ad=5.97137e+07 pd=221088 as=0 ps=0 
M4317 GND n_90 p6 GND efet w=6204 l=564
+ ad=0 pd=0 as=1.02939e+07 ps=28200 
M4318 Pout3 n_1194 GND GND efet w=9353 l=611
+ ad=1.36339e+07 pd=34216 as=0 ps=0 
M4319 Vdd p6 p6 GND dfet w=940 l=1034
+ ad=0 pd=0 as=2.57128e+06 ps=7896 
M4320 Pout3 Pout3 Vdd GND dfet w=940 l=940
+ ad=4.38442e+07 pd=156792 as=0 ps=0 
M4321 p6 H1x1 idb6 GND efet w=2350 l=752
+ ad=0 pd=0 as=0 ps=0 
M4322 Pout3 H1x1 idb3 GND efet w=2350 l=752
+ ad=0 pd=0 as=0 ps=0 
M4323 GND idb6 n_1416 GND efet w=6909 l=611
+ ad=0 pd=0 as=7.0688e+06 ps=21056 
M4324 n_1600 idb3 GND GND efet w=6862 l=564
+ ad=7.0688e+06 pd=21244 as=0 ps=0 
M4325 n_455 n_279 GND GND efet w=5734 l=564
+ ad=3.23398e+06 pd=12596 as=0 ps=0 
M4326 n_1082 pipeUNK16 n_455 GND efet w=5734 l=564
+ ad=0 pd=0 as=0 ps=0 
M4327 n_31 p0 GND GND efet w=6157 l=611
+ ad=1.12482e+07 pd=28952 as=0 ps=0 
M4328 Vdd n_1471 n_1471 GND dfet w=940 l=1598
+ ad=0 pd=0 as=1.2821e+07 ps=39856 
M4329 p0 cp1 n_1082 GND efet w=1222 l=752
+ ad=1.70535e+06 pd=6580 as=0 ps=0 
M4330 n_31 n_31 Vdd GND dfet w=940 l=1128
+ ad=7.66258e+07 pd=269216 as=0 ps=0 
M4331 n_1471 D1x1 GND GND efet w=3807 l=611
+ ad=3.83482e+06 pd=13348 as=0 ps=0 
M4332 n_1082 n_1082 Vdd GND dfet w=940 l=1974
+ ad=4.03805e+06 pd=10340 as=0 ps=0 
M4333 n_31 cclk pipeUNK16 GND efet w=1128 l=658
+ ad=0 pd=0 as=1.44027e+06 ps=6016 
M4334 p4 n_1471 GND GND efet w=8366 l=658
+ ad=1.40316e+07 pd=36284 as=0 ps=0 
M4335 p4 p4 Vdd GND dfet w=1034 l=940
+ ad=2.49175e+06 pd=8084 as=0 ps=0 
M4336 n_270 n_503 GND GND efet w=3008 l=658
+ ad=4.2943e+06 pd=13724 as=0 ps=0 
M4337 Vdd n_270 n_270 GND dfet w=940 l=1222
+ ad=0 pd=0 as=1.05846e+08 ps=385212 
M4338 pipeUNK02 cclk n_774 GND efet w=940 l=752
+ ad=1.29006e+06 pd=6392 as=0 ps=0 
M4339 GND pipeUNK02 n_1492 GND efet w=3854 l=564
+ ad=0 pd=0 as=4.56821e+06 ps=13348 
M4340 GND db4 n_1075 GND efet w=12690 l=658
+ ad=0 pd=0 as=0 ps=0 
M4341 n_1281 db3 GND GND efet w=12972 l=564
+ ad=0 pd=0 as=0 ps=0 
M4342 n_1075 n_1075 Vdd GND dfet w=940 l=658
+ ad=1.5463e+06 pd=6016 as=0 ps=0 
M4343 GND db5 n_1588 GND efet w=13019 l=517
+ ad=0 pd=0 as=0 ps=0 
M4344 n_93 db0 GND GND efet w=13442 l=1034
+ ad=0 pd=0 as=0 ps=0 
M4345 Vdd n_1281 n_1281 GND dfet w=940 l=658
+ ad=0 pd=0 as=1.60815e+06 ps=6204 
M4346 n_1588 n_1588 Vdd GND dfet w=940 l=658
+ ad=1.5463e+06 pd=6016 as=0 ps=0 
M4347 Vdd n_1492 n_1492 GND dfet w=846 l=1692
+ ad=0 pd=0 as=2.24081e+07 ps=73884 
M4348 GND db1 n_1319 GND efet w=13019 l=705
+ ad=0 pd=0 as=0 ps=0 
M4349 n_62 db7 GND GND efet w=13066 l=564
+ ad=0 pd=0 as=0 ps=0 
M4350 Vdd n_93 n_93 GND dfet w=940 l=752
+ ad=0 pd=0 as=1.7672e+06 ps=6204 
M4351 n_1319 n_1319 Vdd GND dfet w=940 l=658
+ ad=1.5463e+06 pd=6016 as=0 ps=0 
M4352 Vdd n_62 n_62 GND dfet w=940 l=564
+ ad=0 pd=0 as=1.3254e+06 ps=5828 
M4353 n_111 n_111 Vdd GND dfet w=940 l=658
+ ad=1.5463e+06 pd=6016 as=0 ps=0 
M4354 GND db2 n_111 GND efet w=11609 l=705
+ ad=0 pd=0 as=0 ps=0 
M4355 GND db6 n_374 GND efet w=11562 l=658
+ ad=0 pd=0 as=0 ps=0 
M4356 n_374 n_374 Vdd GND dfet w=846 l=752
+ ad=1.7672e+06 pd=6204 as=0 ps=0 
M4357 pipeUNK04 cclk n_1194 GND efet w=1128 l=752
+ ad=2.72149e+06 pd=7896 as=9.29547e+06 ps=27260 
M4358 GND p3 n_1194 GND efet w=5640 l=658
+ ad=0 pd=0 as=0 ps=0 
M4359 n_1495 cp1 p3 GND efet w=1128 l=752
+ ad=1.1584e+07 pd=26696 as=1.62582e+06 ps=7520 
M4360 n_1194 n_1194 Vdd GND dfet w=940 l=1316
+ ad=2.28411e+07 pd=75764 as=0 ps=0 
M4361 n_1495 n_1495 Vdd GND dfet w=1034 l=1880
+ ad=3.35768e+06 pd=8648 as=0 ps=0 
M4362 n_1644 n_1457 n_1495 GND efet w=3102 l=564
+ ad=6.04382e+06 pd=15040 as=0 ps=0 
M4363 GND pipeUNK04 n_1644 GND efet w=6204 l=658
+ ad=0 pd=0 as=0 ps=0 
M4364 GND DBNeg n_648 GND efet w=4465 l=611
+ ad=0 pd=0 as=2.41223e+06 ps=9964 
M4365 n_648 n_754 n_1181 GND efet w=4465 l=611
+ ad=0 pd=0 as=1.10008e+07 ps=30644 
M4366 n_1069 cclk n_1177 GND efet w=1034 l=658
+ ad=0 pd=0 as=3.02191e+06 ps=10528 
M4367 GND n_587 n_299 GND efet w=1974 l=658
+ ad=0 pd=0 as=1.21318e+07 ps=32524 
M4368 x_op_T__adc_sbc cclk pipeUNK03 GND efet w=1128 l=846
+ ad=0 pd=0 as=3.14562e+06 ps=10152 
M4369 n_299 n_1245 n_1723 GND efet w=3008 l=658
+ ad=0 pd=0 as=4.99234e+06 ps=14476 
M4370 Vdd n_299 n_299 GND dfet w=940 l=1880
+ ad=0 pd=0 as=6.31774e+06 ps=18800 
M4371 n_1723 pipeUNK03 GND GND efet w=6298 l=564
+ ad=0 pd=0 as=0 ps=0 
M4372 Vdd n_1614 n_1614 GND dfet w=940 l=1692
+ ad=0 pd=0 as=9.86098e+06 ps=28576 
M4373 n_1614 n_1177 GND GND efet w=4183 l=611
+ ad=1.43673e+07 pd=41172 as=0 ps=0 
M4374 n_1595 n_754 GND GND efet w=2632 l=658
+ ad=2.75683e+06 pd=11092 as=0 ps=0 
M4375 n_1181 n_1181 Vdd GND dfet w=940 l=1880
+ ad=1.04176e+07 pd=30456 as=0 ps=0 
M4376 Vdd n_1595 n_1595 GND dfet w=940 l=1504
+ ad=0 pd=0 as=1.01437e+07 ps=31396 
M4377 n_1181 n_1595 n_793 GND efet w=2914 l=564
+ ad=0 pd=0 as=4.84213e+06 ps=14100 
M4378 n_793 pipeUNK13 GND GND efet w=6110 l=564
+ ad=0 pd=0 as=0 ps=0 
M4379 n_1614 pipeUNK03 GND GND efet w=3948 l=564
+ ad=0 pd=0 as=0 ps=0 
M4380 GND n_1111 n_1470 GND efet w=3008 l=658
+ ad=0 pd=0 as=1.69651e+06 ps=7144 
M4381 n_1546 n_781 GND GND efet w=3008 l=658
+ ad=1.69651e+06 pd=7144 as=0 ps=0 
M4382 n_1495 n_1600 n_1546 GND efet w=3008 l=564
+ ad=0 pd=0 as=0 ps=0 
M4383 n_1445 n_270 n_1495 GND efet w=3008 l=658
+ ad=1.41376e+06 pd=6956 as=0 ps=0 
M4384 GND n_1492 n_1445 GND efet w=3008 l=564
+ ad=0 pd=0 as=0 ps=0 
M4385 n_1470 n_1416 n_299 GND efet w=3008 l=658
+ ad=0 pd=0 as=0 ps=0 
M4386 GND n_1111 n_1614 GND efet w=1880 l=658
+ ad=0 pd=0 as=0 ps=0 
M4387 pipeUNK13 cclk n_1045 GND efet w=1128 l=940
+ ad=1.19286e+06 pd=6580 as=7.1925e+06 ps=23500 
M4388 n_1181 cp1 n_69 GND efet w=1222 l=846
+ ad=0 pd=0 as=1.37842e+06 ps=7520 
M4389 n_1045 n_1045 Vdd GND dfet w=1034 l=1128
+ ad=4.4286e+07 pd=149836 as=0 ps=0 
M4390 GND n_69 n_1045 GND efet w=7567 l=611
+ ad=0 pd=0 as=0 ps=0 
M4391 n_299 n_1614 n_1616 GND efet w=3008 l=752
+ ad=0 pd=0 as=4.56821e+06 ps=14288 
M4392 n_1457 n_1457 Vdd GND dfet w=1034 l=1316
+ ad=7.58129e+06 pd=24816 as=0 ps=0 
M4393 n_1457 n_781 GND GND efet w=2350 l=658
+ ad=7.77568e+06 pd=16168 as=0 ps=0 
M4394 GND n_1492 n_1457 GND efet w=2350 l=658
+ ad=0 pd=0 as=0 ps=0 
M4395 n_1616 pipeUNK05 GND GND efet w=6439 l=611
+ ad=0 pd=0 as=0 ps=0 
M4396 n_307 n_31 GND GND efet w=3572 l=658
+ ad=1.26178e+07 pd=35720 as=0 ps=0 
M4397 n_299 cp1 n_1625 GND efet w=1222 l=752
+ ad=0 pd=0 as=1.68768e+06 ps=7520 
M4398 GND nop_branch_bit7 n_307 GND efet w=3807 l=611
+ ad=0 pd=0 as=0 ps=0 
M4399 GND n_1625 n_90 GND efet w=6533 l=611
+ ad=0 pd=0 as=7.9524e+06 ps=22748 
M4400 pipeUNK05 cclk n_90 GND efet w=1222 l=752
+ ad=1.85556e+06 pd=6768 as=0 ps=0 
M4401 n_307 n_846 GND GND efet w=3901 l=611
+ ad=0 pd=0 as=0 ps=0 
M4402 GND n_31 Pout0 GND efet w=6298 l=658
+ ad=0 pd=0 as=9.71076e+06 ps=29140 
M4403 Pout1 n_318 GND GND efet w=7896 l=564
+ ad=1.09831e+07 pd=30456 as=0 ps=0 
M4404 n_1416 n_1416 Vdd GND dfet w=940 l=1128
+ ad=2.90881e+07 pd=103776 as=0 ps=0 
M4405 n_1600 n_1600 Vdd GND dfet w=940 l=1034
+ ad=1.99605e+07 pd=78208 as=0 ps=0 
M4406 GND alucout n_206 GND efet w=11891 l=611
+ ad=0 pd=0 as=0 ps=0 
M4407 p4 H1x1 idb4 GND efet w=2350 l=658
+ ad=0 pd=0 as=0 ps=0 
M4408 GND dpc36_nIPC dpc34_PCLC GND efet w=5264 l=752
+ ad=0 pd=0 as=4.01419e+07 ps=122200 
M4409 n_146 cclk a0 GND efet w=1128 l=658
+ ad=1.46236e+07 pd=37600 as=3.86133e+06 ps=12784 
M4410 a0 dpc23_SBAC sb0 GND efet w=1034 l=658
+ ad=0 pd=0 as=0 ps=0 
M4411 n_146 n_5 GND GND efet w=7520 l=564
+ ad=0 pd=0 as=0 ps=0 
M4412 n_613 n_613 Vdd GND dfet w=940 l=1504
+ ad=1.9722e+07 pd=70688 as=0 ps=0 
M4413 Vdd dasb1 dasb1 GND dfet w=846 l=1598
+ ad=0 pd=0 as=3.44604e+06 ps=9588 
M4414 GND a0 n_5 GND efet w=4136 l=564
+ ad=0 pd=0 as=6.92742e+06 ps=18048 
M4415 n_146 dpc26_ACDB idb0 GND efet w=1222 l=752
+ ad=0 pd=0 as=0 ps=0 
M4416 idb0 dpc25_SBDB sb0 GND efet w=2162 l=658
+ ad=0 pd=0 as=0 ps=0 
M4417 sb0 dpc24_ACSB n_146 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M4418 Vdd n_5 n_5 GND dfet w=940 l=1504
+ ad=0 pd=0 as=8.91552e+06 ps=27260 
M4419 n_1322 n_320 GND GND efet w=3290 l=564
+ ad=1.85556e+06 pd=7708 as=0 ps=0 
M4420 dasb1 n_36 n_1322 GND efet w=3290 l=564
+ ad=6.52097e+06 pd=17108 as=0 ps=0 
M4421 a1 dpc23_SBAC dasb1 GND efet w=1034 l=658
+ ad=4.00271e+06 pd=13160 as=0 ps=0 
M4422 GND n_735 dasb1 GND efet w=1692 l=564
+ ad=0 pd=0 as=0 ps=0 
M4423 n_735 n_320 GND GND efet w=2162 l=564
+ ad=5.03652e+06 pd=14852 as=0 ps=0 
M4424 GND n_36 n_735 GND efet w=2397 l=611
+ ad=0 pd=0 as=0 ps=0 
M4425 n_1341 cclk n_695 GND efet w=1034 l=752
+ ad=1.13984e+06 pd=5264 as=6.60049e+06 ps=21620 
M4426 Vdd n_695 n_695 GND dfet w=846 l=1410
+ ad=0 pd=0 as=5.04536e+06 ps=15980 
M4427 n_619 n_700 GND GND efet w=4418 l=564
+ ad=2.47408e+06 pd=9964 as=0 ps=0 
M4428 n_695 C34 n_619 GND efet w=4418 l=564
+ ad=0 pd=0 as=0 ps=0 
M4429 n_320 sb1 GND GND efet w=5076 l=658
+ ad=4.10874e+06 pd=13724 as=0 ps=0 
M4430 n_735 n_735 Vdd GND dfet w=846 l=1598
+ ad=7.88171e+06 pd=25004 as=0 ps=0 
M4431 Vdd n_929 n_929 GND dfet w=940 l=1128
+ ad=0 pd=0 as=2.88937e+06 ps=9024 
M4432 n_929 cclk a1 GND efet w=1128 l=752
+ ad=1.40139e+07 pd=35720 as=0 ps=0 
M4433 n_929 n_1549 GND GND efet w=7520 l=658
+ ad=0 pd=0 as=0 ps=0 
M4434 GND a1 n_1549 GND efet w=4324 l=564
+ ad=0 pd=0 as=5.92012e+06 ps=18800 
M4435 Vdd n_320 n_320 GND dfet w=846 l=1598
+ ad=0 pd=0 as=9.01272e+06 ps=29892 
M4436 Vdd dasb2 dasb2 GND dfet w=846 l=1598
+ ad=0 pd=0 as=3.44604e+06 ps=9588 
M4437 n_1656 n_1580 GND GND efet w=3713 l=611
+ ad=1.84672e+06 pd=8460 as=0 ps=0 
M4438 dasb2 n_613 n_1656 GND efet w=3478 l=564
+ ad=6.9451e+06 pd=17672 as=0 ps=0 
M4439 adh0 dpc27_SBADH sb0 GND efet w=1974 l=658
+ ad=1.45352e+07 pd=41172 as=0 ps=0 
M4440 GND dpc28_0ADH0 adh0 GND efet w=1974 l=752
+ ad=0 pd=0 as=0 ps=0 
M4441 n_929 dpc26_ACDB idb1 GND efet w=1410 l=752
+ ad=0 pd=0 as=0 ps=0 
M4442 idb1 dpc25_SBDB sb1 GND efet w=2068 l=658
+ ad=0 pd=0 as=0 ps=0 
M4443 sb1 dpc24_ACSB n_929 GND efet w=1222 l=752
+ ad=0 pd=0 as=0 ps=0 
M4444 Vdd n_1549 n_1549 GND dfet w=846 l=1504
+ ad=0 pd=0 as=9.32198e+06 ps=26696 
M4445 a2 dpc23_SBAC dasb2 GND efet w=1034 l=658
+ ad=3.82599e+06 pd=12972 as=0 ps=0 
M4446 Vdd n_1618 n_1618 GND dfet w=940 l=1222
+ ad=0 pd=0 as=2.80985e+06 ps=9212 
M4447 GND n_1159 dasb2 GND efet w=1692 l=564
+ ad=0 pd=0 as=0 ps=0 
M4448 n_1159 n_1580 GND GND efet w=1880 l=564
+ ad=4.59472e+06 pd=13348 as=0 ps=0 
M4449 GND n_613 n_1159 GND efet w=2303 l=611
+ ad=0 pd=0 as=0 ps=0 
M4450 n_1580 sb2 GND GND efet w=1410 l=470
+ ad=5.60202e+06 pd=17296 as=0 ps=0 
M4451 Vdd n_1580 n_1580 GND dfet w=752 l=1316
+ ad=0 pd=0 as=7.99658e+06 ps=26508 
M4452 n_1159 n_1159 Vdd GND dfet w=846 l=1598
+ ad=7.81986e+06 pd=23688 as=0 ps=0 
M4453 n_1580 sb2 GND GND efet w=4324 l=564
+ ad=0 pd=0 as=0 ps=0 
M4454 Vdd dasb3 dasb3 GND dfet w=940 l=1598
+ ad=0 pd=0 as=3.44604e+06 ps=9588 
M4455 n_1179 C34 GND GND efet w=2303 l=611
+ ad=1.04707e+07 pd=32524 as=0 ps=0 
M4456 GND dpc22_nDSA n_1179 GND efet w=1974 l=658
+ ad=0 pd=0 as=0 ps=0 
M4457 n_1584 n_876 GND GND efet w=4794 l=564
+ ad=2.4299e+06 pd=10528 as=0 ps=0 
M4458 n_345 n_8 n_1584 GND efet w=4700 l=658
+ ad=8.76531e+06 pd=21432 as=0 ps=0 
M4459 n_1686 n_432 GND GND efet w=3196 l=658
+ ad=1.50212e+06 pd=7332 as=0 ps=0 
M4460 dasb3 n_345 n_1686 GND efet w=3196 l=564
+ ad=6.49446e+06 pd=16168 as=0 ps=0 
M4461 n_1618 cclk a2 GND efet w=1034 l=752
+ ad=1.42525e+07 pd=36472 as=0 ps=0 
M4462 n_1618 n_419 GND GND efet w=7614 l=564
+ ad=0 pd=0 as=0 ps=0 
M4463 GND a2 n_419 GND efet w=4136 l=564
+ ad=0 pd=0 as=6.5298e+06 ps=19176 
M4464 Vdd cclk adh0 GND efet w=2162 l=658
+ ad=0 pd=0 as=0 ps=0 
M4465 GND dpc29_0ADH17 adh1 GND efet w=2162 l=752
+ ad=0 pd=0 as=1.45264e+07 ps=38352 
M4466 adh1 dpc27_SBADH sb1 GND efet w=2162 l=658
+ ad=0 pd=0 as=0 ps=0 
M4467 Vdd cclk adh1 GND efet w=2256 l=564
+ ad=0 pd=0 as=0 ps=0 
M4468 dpc35_PCHC dpc35_PCHC Vdd GND dfet w=1222 l=658
+ ad=5.06568e+07 pd=201536 as=0 ps=0 
M4469 n_311 n_311 Vdd GND dfet w=846 l=1504
+ ad=1.20258e+07 pd=39480 as=0 ps=0 
M4470 Vdd cclk adl0 GND efet w=2068 l=658
+ ad=0 pd=0 as=0 ps=0 
M4471 Vdd n_919 n_919 GND dfet w=846 l=1410
+ ad=0 pd=0 as=1.92536e+07 ps=65424 
M4472 n_1229 cclk npchp0 GND efet w=1128 l=752
+ ad=8.22632e+06 pd=21996 as=1.96159e+06 ps=7520 
M4473 pchp0 dpc31_PCHPCH pch0 GND efet w=1316 l=846
+ ad=1.32893e+07 pd=35344 as=5.21324e+06 ps=14664 
M4474 pch0 dpc30_ADHPCH adh0 GND efet w=1316 l=752
+ ad=0 pd=0 as=0 ps=0 
M4475 GND npchp0 pchp0 GND efet w=3948 l=658
+ ad=0 pd=0 as=0 ps=0 
M4476 n_856 dpc34_PCLC n_919 GND efet w=4230 l=658
+ ad=4.17943e+06 pd=11468 as=4.60356e+06 ps=13724 
M4477 GND n_311 n_856 GND efet w=4136 l=564
+ ad=0 pd=0 as=0 ps=0 
M4478 n_1010 pch0 GND GND efet w=3666 l=564
+ ad=3.68461e+06 pd=11092 as=0 ps=0 
M4479 Vdd n_1010 n_1010 GND dfet w=940 l=1880
+ ad=0 pd=0 as=9.78145e+06 ps=32336 
M4480 pchp0 dpc33_PCHDB idb0 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M4481 adh0 dpc32_PCHADH pchp0 GND efet w=1316 l=752
+ ad=0 pd=0 as=0 ps=0 
M4482 adl1 cclk Vdd GND efet w=2068 l=658
+ ad=0 pd=0 as=0 ps=0 
M4483 pchp1 dpc31_PCHPCH pch1 GND efet w=1316 l=752
+ ad=1.50654e+07 pd=40044 as=5.23091e+06 ps=14852 
M4484 pch1 dpc30_ADHPCH adh1 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M4485 n_1618 dpc26_ACDB idb2 GND efet w=1316 l=752
+ ad=0 pd=0 as=0 ps=0 
M4486 idb2 dpc25_SBDB sb2 GND efet w=2115 l=517
+ ad=0 pd=0 as=0 ps=0 
M4487 sb2 dpc24_ACSB n_1618 GND efet w=1410 l=752
+ ad=0 pd=0 as=0 ps=0 
M4488 Vdd n_419 n_419 GND dfet w=940 l=1504
+ ad=0 pd=0 as=8.86251e+06 ps=26508 
M4489 a3 dpc23_SBAC dasb3 GND efet w=1034 l=658
+ ad=4.03805e+06 pd=12784 as=0 ps=0 
M4490 Vdd n_1654 n_1654 GND dfet w=940 l=1222
+ ad=0 pd=0 as=2.80985e+06 ps=9212 
M4491 GND n_1097 dasb3 GND efet w=2350 l=564
+ ad=0 pd=0 as=0 ps=0 
M4492 n_1279 n_986 n_345 GND efet w=3666 l=564
+ ad=2.06762e+06 pd=8460 as=0 ps=0 
M4493 GND n_600 n_1279 GND efet w=3666 l=564
+ ad=0 pd=0 as=0 ps=0 
M4494 n_1097 n_432 GND GND efet w=2961 l=611
+ ad=4.93932e+06 pd=16920 as=0 ps=0 
M4495 n_1179 n_1179 Vdd GND dfet w=846 l=1410
+ ad=6.3089e+06 pd=18988 as=0 ps=0 
M4496 n_8 n_551 GND GND efet w=3478 l=564
+ ad=3.95853e+06 pd=11656 as=0 ps=0 
M4497 GND n_345 n_1097 GND efet w=3055 l=611
+ ad=0 pd=0 as=0 ps=0 
M4498 n_345 n_345 Vdd GND dfet w=940 l=1504
+ ad=8.32351e+06 pd=27260 as=0 ps=0 
M4499 n_432 sb3 GND GND efet w=1222 l=658
+ ad=7.58129e+06 pd=22748 as=0 ps=0 
M4500 n_8 n_8 Vdd GND dfet w=940 l=940
+ ad=3.7067e+07 pd=132540 as=0 ps=0 
M4501 n_1097 n_1097 Vdd GND dfet w=846 l=1504
+ ad=9.02156e+06 pd=28764 as=0 ps=0 
M4502 n_1179 cclk n_393 GND efet w=1034 l=752
+ ad=0 pd=0 as=1.01614e+06 ps=5076 
M4503 Vdd n_306 n_306 GND dfet w=940 l=1504
+ ad=0 pd=0 as=4.20594e+06 ps=11656 
M4504 n_306 cclk n_581 GND efet w=1128 l=752
+ ad=6.58282e+06 pd=21808 as=1.56397e+06 ps=6580 
M4505 GND dpc22_nDSA n_306 GND efet w=3384 l=564
+ ad=0 pd=0 as=0 ps=0 
M4506 n_432 sb3 GND GND efet w=3196 l=658
+ ad=0 pd=0 as=0 ps=0 
M4507 Vdd n_432 n_432 GND dfet w=846 l=1504
+ ad=0 pd=0 as=1.04265e+07 ps=33840 
M4508 n_1654 cclk a3 GND efet w=1128 l=658
+ ad=1.46766e+07 pd=36096 as=0 ps=0 
M4509 n_1654 n_947 GND GND efet w=7614 l=564
+ ad=0 pd=0 as=0 ps=0 
M4510 GND a3 n_947 GND efet w=4136 l=658
+ ad=0 pd=0 as=6.77721e+06 ps=19176 
M4511 adh2 dpc27_SBADH sb2 GND efet w=2068 l=752
+ ad=1.56574e+07 pd=42864 as=0 ps=0 
M4512 GND dpc29_0ADH17 adh2 GND efet w=2068 l=658
+ ad=0 pd=0 as=0 ps=0 
M4513 n_1654 dpc26_ACDB idb3 GND efet w=1316 l=752
+ ad=0 pd=0 as=0 ps=0 
M4514 idb3 dpc25_SBDB sb3 GND efet w=2068 l=564
+ ad=0 pd=0 as=0 ps=0 
M4515 sb3 dpc24_ACSB n_1654 GND efet w=1316 l=846
+ ad=0 pd=0 as=0 ps=0 
M4516 Vdd n_947 n_947 GND dfet w=940 l=1504
+ ad=0 pd=0 as=8.57976e+06 ps=26508 
M4517 GND alucout n_811 GND efet w=3854 l=564
+ ad=0 pd=0 as=8.20864e+06 ps=20868 
M4518 n_753 n_811 GND GND efet w=1128 l=564
+ ad=9.54288e+06 pd=26508 as=0 ps=0 
M4519 a4 dpc23_SBAC sb4 GND efet w=1128 l=658
+ ad=3.73763e+06 pd=12596 as=0 ps=0 
M4520 n_551 n_393 GND GND efet w=4136 l=658
+ ad=5.09837e+06 pd=17108 as=0 ps=0 
M4521 GND n_581 n_838 GND efet w=4230 l=564
+ ad=0 pd=0 as=5.92896e+06 ps=16732 
M4522 n_811 n_838 GND GND efet w=4606 l=658
+ ad=0 pd=0 as=0 ps=0 
M4523 n_753 n_811 GND GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M4524 n_753 n_1257 GND GND efet w=2914 l=564
+ ad=0 pd=0 as=0 ps=0 
M4525 n_551 n_551 Vdd GND dfet w=846 l=1410
+ ad=1.40139e+07 pd=49444 as=0 ps=0 
M4526 n_838 n_838 Vdd GND dfet w=940 l=1598
+ ad=7.71383e+06 pd=22748 as=0 ps=0 
M4527 n_811 n_811 Vdd GND dfet w=846 l=846
+ ad=3.30378e+07 pd=125396 as=0 ps=0 
M4528 Vdd n_761 n_761 GND dfet w=752 l=1504
+ ad=0 pd=0 as=2.78864e+07 ps=95316 
M4529 GND alu5 n_761 GND efet w=3478 l=752
+ ad=0 pd=0 as=5.91128e+06 ps=17296 
M4530 Vdd n_233 n_233 GND dfet w=846 l=1504
+ ad=0 pd=0 as=2.70735e+07 ps=98512 
M4531 n_233 n_761 n_970 GND efet w=4277 l=611
+ ad=6.45028e+06 pd=20116 as=3.57858e+06 ps=10716 
M4532 n_970 n_149 GND GND efet w=3572 l=564
+ ad=0 pd=0 as=0 ps=0 
M4533 n_753 n_753 Vdd GND dfet w=846 l=1504
+ ad=1.07711e+07 pd=34780 as=0 ps=0 
M4534 n_762 n_149 GND GND efet w=3384 l=564
+ ad=5.8671e+06 pd=17860 as=0 ps=0 
M4535 GND n_761 n_762 GND efet w=3384 l=658
+ ad=0 pd=0 as=0 ps=0 
M4536 adl7 dpc21_ADDADL alu7 GND efet w=1504 l=752
+ ad=0 pd=0 as=1.09831e+07 ps=32524 
M4537 GND notalu7 alu7 GND efet w=9494 l=658
+ ad=0 pd=0 as=0 ps=0 
M4538 Vdd notaluvout notaluvout GND dfet w=940 l=1504
+ ad=0 pd=0 as=5.89361e+06 ps=21244 
M4539 GND n_1315 n_826 GND efet w=10716 l=752
+ ad=0 pd=0 as=1.6055e+07 ps=37036 
M4540 GND n_617 n_1140 GND efet w=10716 l=564
+ ad=0 pd=0 as=1.65233e+07 ps=37600 
M4541 Vdd abh0 abh0 GND dfet w=846 l=1410
+ ad=0 pd=0 as=2.27174e+07 ps=73696 
M4542 GND n_171 ab7 GND efet w=10904 l=3384
+ ad=0 pd=0 as=1.71454e+08 ps=260192 
M4543 n_1668 cp1 n_705 GND efet w=1034 l=846
+ ad=0 pd=0 as=583176 ps=3196 
M4544 n_705 ADH_ABH nABH0 GND efet w=1034 l=752
+ ad=0 pd=0 as=3.35768e+06 ps=11280 
M4545 GND n_171 ab7 GND efet w=19928 l=564
+ ad=0 pd=0 as=0 ps=0 
M4546 ab7 n_171 GND GND efet w=19928 l=564
+ ad=0 pd=0 as=0 ps=0 
M4547 ab7 n_171 GND GND efet w=41125 l=611
+ ad=0 pd=0 as=0 ps=0 
M4548 n_826 abh0 Vdd GND dfet w=1692 l=658
+ ad=0 pd=0 as=0 ps=0 
M4549 Vdd n_1315 n_1315 GND dfet w=846 l=940
+ ad=0 pd=0 as=1.81315e+07 ps=57528 
M4550 Vdd n_322 ab7 GND efet w=24064 l=564
+ ad=0 pd=0 as=0 ps=0 
M4551 nABH0 cclk n_381 GND efet w=1034 l=658
+ ad=0 pd=0 as=1.13366e+07 ps=35532 
M4552 Vdd n_1315 n_381 GND dfet w=1974 l=752
+ ad=0 pd=0 as=0 ps=0 
M4553 GND abh0 n_1315 GND efet w=3384 l=658
+ ad=0 pd=0 as=4.05572e+06 ps=12220 
M4554 GND abh0 n_381 GND efet w=14570 l=658
+ ad=0 pd=0 as=0 ps=0 
M4555 GND n_381 ab8 GND efet w=1316 l=564
+ ad=0 pd=0 as=1.61496e+08 ps=216952 
M4556 GND n_381 ab8 GND efet w=3948 l=564
+ ad=0 pd=0 as=0 ps=0 
M4557 Vdd n_322 ab7 GND efet w=24816 l=658
+ ad=0 pd=0 as=0 ps=0 
M4558 Vdd n_322 ab7 GND efet w=22090 l=658
+ ad=0 pd=0 as=0 ps=0 
M4559 Vdd n_322 ab7 GND efet w=21949 l=611
+ ad=0 pd=0 as=0 ps=0 
M4560 ab8 n_381 GND GND efet w=15322 l=564
+ ad=0 pd=0 as=0 ps=0 
M4561 GND n_381 ab8 GND efet w=15322 l=658
+ ad=0 pd=0 as=0 ps=0 
M4562 ab8 n_381 GND GND efet w=15322 l=658
+ ad=0 pd=0 as=0 ps=0 
M4563 GND n_381 ab8 GND efet w=15322 l=658
+ ad=0 pd=0 as=0 ps=0 
M4564 ab8 n_381 GND GND efet w=15322 l=564
+ ad=0 pd=0 as=0 ps=0 
M4565 Vdd n_826 ab8 GND efet w=38963 l=611
+ ad=0 pd=0 as=0 ps=0 
M4566 Vdd n_826 ab8 GND efet w=29845 l=611
+ ad=0 pd=0 as=0 ps=0 
M4567 Vdd n_826 ab8 GND efet w=14946 l=658
+ ad=0 pd=0 as=0 ps=0 
M4568 ab9 n_1140 Vdd GND efet w=14946 l=564
+ ad=1.62688e+08 pd=217516 as=0 ps=0 
M4569 Vdd n_1140 ab9 GND efet w=29798 l=658
+ ad=0 pd=0 as=0 ps=0 
M4570 Vdd n_1140 ab9 GND efet w=39151 l=611
+ ad=0 pd=0 as=0 ps=0 
M4571 Vdd abh1 n_1140 GND dfet w=1692 l=752
+ ad=0 pd=0 as=0 ps=0 
M4572 n_617 abh1 GND GND efet w=4230 l=658
+ ad=3.93202e+06 pd=13536 as=0 ps=0 
M4573 Vdd n_617 n_617 GND dfet w=940 l=940
+ ad=0 pd=0 as=1.77427e+07 ps=63920 
M4574 abh1 abh1 Vdd GND dfet w=846 l=1316
+ ad=2.15687e+07 pd=62228 as=0 ps=0 
M4575 GND nABH1 abh1 GND efet w=6110 l=658
+ ad=0 pd=0 as=5.31927e+06 ps=17484 
M4576 n_637 n_637 Vdd GND dfet w=846 l=1410
+ ad=1.14868e+07 pd=42112 as=0 ps=0 
M4577 GND n_637 notaluvout GND efet w=2867 l=611
+ ad=0 pd=0 as=0 ps=0 
M4578 alu7 dpc19_ADDSB7 sb7 GND efet w=1880 l=658
+ ad=0 pd=0 as=0 ps=0 
M4579 DC78_phi2 cclk DC78 GND efet w=1128 l=752
+ ad=1.43143e+06 pd=6768 as=0 ps=0 
M4580 C78_phi2 cclk C78 GND efet w=1034 l=752
+ ad=1.28122e+06 pd=6580 as=9.52521e+06 ps=27824 
M4581 alu7 alu7 Vdd GND dfet w=940 l=1222
+ ad=3.13678e+06 pd=9776 as=0 ps=0 
M4582 n_762 n_762 Vdd GND dfet w=846 l=1504
+ ad=2.03228e+07 pd=69372 as=0 ps=0 
M4583 Vdd n_149 n_149 GND dfet w=846 l=1598
+ ad=0 pd=0 as=8.91552e+06 ps=29140 
M4584 GND alu6 n_149 GND efet w=4653 l=611
+ ad=0 pd=0 as=7.39573e+06 ps=21996 
M4585 C78 nC78 GND GND efet w=5546 l=564
+ ad=0 pd=0 as=0 ps=0 
M4586 n_408 cclk notaluvout GND efet w=1034 l=658
+ ad=1.8644e+06 pd=8084 as=0 ps=0 
M4587 GND n_408 aluvout GND efet w=12220 l=658
+ ad=0 pd=0 as=1.45264e+07 ps=37036 
M4588 n_1203 n_1135 GND GND efet w=4324 l=564
+ ad=2.5271e+06 pd=9776 as=0 ps=0 
M4589 Vdd dasb5 dasb5 GND dfet w=846 l=1598
+ ad=0 pd=0 as=3.47255e+06 ps=9588 
M4590 Vdd n_1344 n_1344 GND dfet w=940 l=1222
+ ad=0 pd=0 as=3.05726e+06 ps=9400 
M4591 n_1344 cclk a4 GND efet w=1034 l=752
+ ad=1.32452e+07 pd=36284 as=0 ps=0 
M4592 n_1344 n_556 GND GND efet w=7708 l=658
+ ad=0 pd=0 as=0 ps=0 
M4593 GND a4 n_556 GND efet w=4042 l=564
+ ad=0 pd=0 as=6.67118e+06 ps=19176 
M4594 Vdd cclk adh2 GND efet w=2068 l=658
+ ad=0 pd=0 as=0 ps=0 
M4595 adh3 dpc27_SBADH sb3 GND efet w=1974 l=658
+ ad=1.75571e+07 pd=46812 as=0 ps=0 
M4596 GND dpc29_0ADH17 adh3 GND efet w=1974 l=752
+ ad=0 pd=0 as=0 ps=0 
M4597 n_1344 dpc26_ACDB idb4 GND efet w=1316 l=752
+ ad=0 pd=0 as=0 ps=0 
M4598 idb4 dpc25_SBDB sb4 GND efet w=2068 l=470
+ ad=0 pd=0 as=0 ps=0 
M4599 sb4 dpc24_ACSB n_1344 GND efet w=1316 l=752
+ ad=0 pd=0 as=0 ps=0 
M4600 Vdd n_556 n_556 GND dfet w=846 l=1504
+ ad=0 pd=0 as=9.11875e+06 ps=26696 
M4601 dasb5 n_753 n_1203 GND efet w=3196 l=564
+ ad=5.82292e+06 pd=17296 as=0 ps=0 
M4602 a5 dpc23_SBAC dasb5 GND efet w=1034 l=658
+ ad=4.1971e+06 pd=13160 as=0 ps=0 
M4603 Vdd n_831 n_831 GND dfet w=846 l=1222
+ ad=0 pd=0 as=2.80985e+06 ps=9212 
M4604 GND n_1629 dasb5 GND efet w=1692 l=658
+ ad=0 pd=0 as=0 ps=0 
M4605 GND sb5 n_1135 GND efet w=5828 l=658
+ ad=0 pd=0 as=1.15575e+07 ps=33840 
M4606 n_1629 n_1135 GND GND efet w=1692 l=564
+ ad=5.18673e+06 pd=15416 as=0 ps=0 
M4607 GND n_753 n_1629 GND efet w=2444 l=658
+ ad=0 pd=0 as=0 ps=0 
M4608 Vdd n_1056 n_1056 GND dfet w=940 l=1504
+ ad=0 pd=0 as=8.58859e+06 ps=28012 
M4609 GND n_761 n_1056 GND efet w=2726 l=658
+ ad=0 pd=0 as=3.34884e+06 ps=11656 
M4610 n_1629 n_1629 Vdd GND dfet w=940 l=1598
+ ad=8.46489e+06 pd=25380 as=0 ps=0 
M4611 Vdd n_1135 n_1135 GND dfet w=846 l=1316
+ ad=0 pd=0 as=9.95817e+06 ps=31960 
M4612 Vdd dasb6 dasb6 GND dfet w=846 l=1598
+ ad=0 pd=0 as=3.16329e+06 ps=9776 
M4613 n_1554 n_61 GND GND efet w=3384 l=564
+ ad=1.90858e+06 pd=7896 as=0 ps=0 
M4614 dasb6 n_739 n_1554 GND efet w=3384 l=658
+ ad=5.94663e+06 pd=17860 as=0 ps=0 
M4615 n_831 cclk a5 GND efet w=1128 l=752
+ ad=1.35721e+07 pd=36096 as=0 ps=0 
M4616 n_831 n_1719 GND GND efet w=7567 l=611
+ ad=0 pd=0 as=0 ps=0 
M4617 GND a5 n_1719 GND efet w=4136 l=658
+ ad=0 pd=0 as=5.99964e+06 ps=18988 
M4618 adh4 dpc27_SBADH sb4 GND efet w=2068 l=658
+ ad=1.45264e+07 pd=37976 as=0 ps=0 
M4619 GND dpc29_0ADH17 adh4 GND efet w=2068 l=752
+ ad=0 pd=0 as=0 ps=0 
M4620 n_831 dpc26_ACDB idb5 GND efet w=1316 l=752
+ ad=0 pd=0 as=0 ps=0 
M4621 idb5 dpc25_SBDB sb5 GND efet w=1974 l=658
+ ad=0 pd=0 as=0 ps=0 
M4622 sb5 dpc24_ACSB n_831 GND efet w=1316 l=752
+ ad=0 pd=0 as=0 ps=0 
M4623 Vdd n_1719 n_1719 GND dfet w=846 l=1504
+ ad=0 pd=0 as=9.20711e+06 ps=26696 
M4624 a6 dpc23_SBAC dasb6 GND efet w=1128 l=658
+ ad=4.08223e+06 pd=13160 as=0 ps=0 
M4625 Vdd n_326 n_326 GND dfet w=940 l=1222
+ ad=0 pd=0 as=2.92472e+06 ps=9400 
M4626 n_1080 n_811 GND GND efet w=3290 l=658
+ ad=1.5463e+06 pd=7520 as=0 ps=0 
M4627 n_739 n_1056 n_1080 GND efet w=3290 l=564
+ ad=8.11145e+06 pd=22184 as=0 ps=0 
M4628 GND n_479 dasb6 GND efet w=1692 l=658
+ ad=0 pd=0 as=0 ps=0 
M4629 n_479 n_61 GND GND efet w=1880 l=564
+ ad=5.6197e+06 pd=15980 as=0 ps=0 
M4630 GND n_739 n_479 GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M4631 n_711 n_761 n_739 GND efet w=3196 l=564
+ ad=1.80254e+06 pd=7520 as=0 ps=0 
M4632 GND n_1257 n_711 GND efet w=3196 l=564
+ ad=0 pd=0 as=0 ps=0 
M4633 Vdd n_61 n_61 GND dfet w=940 l=1598
+ ad=0 pd=0 as=7.66081e+06 ps=25380 
M4634 n_739 n_739 Vdd GND dfet w=846 l=1598
+ ad=9.31314e+06 pd=29516 as=0 ps=0 
M4635 n_61 sb6 GND GND efet w=4700 l=564
+ ad=5.15139e+06 pd=16356 as=0 ps=0 
M4636 n_479 n_479 Vdd GND dfet w=940 l=1598
+ ad=8.65928e+06 pd=25944 as=0 ps=0 
M4637 Vdd dasb7 dasb7 GND dfet w=940 l=1504
+ ad=0 pd=0 as=3.13678e+06 ps=9776 
M4638 GND n_762 n_1018 GND efet w=3948 l=658
+ ad=0 pd=0 as=5.19557e+06 ps=15792 
M4639 n_100 n_1018 GND GND efet w=4465 l=611
+ ad=2.56244e+06 pd=10152 as=0 ps=0 
M4640 n_1205 n_811 n_100 GND efet w=4512 l=564
+ ad=7.66965e+06 pd=22184 as=0 ps=0 
M4641 n_1454 n_852 GND GND efet w=3384 l=658
+ ad=1.90858e+06 pd=7896 as=0 ps=0 
M4642 dasb7 n_1205 n_1454 GND efet w=3384 l=658
+ ad=6.19404e+06 pd=16920 as=0 ps=0 
M4643 n_326 cclk a6 GND efet w=1128 l=752
+ ad=1.33954e+07 pd=36472 as=0 ps=0 
M4644 n_326 n_1356 GND GND efet w=7708 l=564
+ ad=0 pd=0 as=0 ps=0 
M4645 GND a6 n_1356 GND efet w=4136 l=658
+ ad=0 pd=0 as=6.37076e+06 ps=18612 
M4646 adh5 dpc27_SBADH sb5 GND efet w=2068 l=658
+ ad=1.47296e+07 pd=40420 as=0 ps=0 
M4647 GND dpc29_0ADH17 adh5 GND efet w=2068 l=752
+ ad=0 pd=0 as=0 ps=0 
M4648 n_326 dpc26_ACDB idb6 GND efet w=1316 l=752
+ ad=0 pd=0 as=0 ps=0 
M4649 idb6 dpc25_SBDB sb6 GND efet w=2068 l=658
+ ad=0 pd=0 as=0 ps=0 
M4650 sb6 dpc24_ACSB n_326 GND efet w=1222 l=752
+ ad=0 pd=0 as=0 ps=0 
M4651 Vdd n_1356 n_1356 GND dfet w=752 l=1598
+ ad=0 pd=0 as=8.97738e+06 ps=26696 
M4652 a7 dpc23_SBAC dasb7 GND efet w=1128 l=752
+ ad=3.82599e+06 pd=12784 as=0 ps=0 
M4653 GND n_260 dasb7 GND efet w=1692 l=564
+ ad=0 pd=0 as=0 ps=0 
M4654 n_260 n_852 GND GND efet w=1786 l=658
+ ad=5.40763e+06 pd=15980 as=0 ps=0 
M4655 GND n_1205 n_260 GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M4656 n_1018 n_1018 Vdd GND dfet w=846 l=940
+ ad=6.68002e+06 pd=22372 as=0 ps=0 
M4657 n_569 n_233 n_1205 GND efet w=3384 l=658
+ ad=1.59048e+06 pd=7708 as=0 ps=0 
M4658 GND n_1257 n_569 GND efet w=3384 l=564
+ ad=0 pd=0 as=0 ps=0 
M4659 n_852 sb7 GND GND efet w=2632 l=564
+ ad=4.6389e+06 pd=14288 as=0 ps=0 
M4660 Vdd n_852 n_852 GND dfet w=940 l=1504
+ ad=0 pd=0 as=8.50023e+06 ps=25944 
M4661 n_1205 n_1205 Vdd GND dfet w=846 l=1598
+ ad=9.2778e+06 pd=27636 as=0 ps=0 
M4662 n_852 sb7 GND GND efet w=1786 l=564
+ ad=0 pd=0 as=0 ps=0 
M4663 n_260 n_260 Vdd GND dfet w=846 l=1598
+ ad=9.25129e+06 pd=26132 as=0 ps=0 
M4664 Vdd n_1592 n_1592 GND dfet w=940 l=1316
+ ad=0 pd=0 as=3.2163e+06 ps=9400 
M4665 n_1592 cclk a7 GND efet w=1034 l=658
+ ad=1.2662e+07 pd=34968 as=0 ps=0 
M4666 n_1592 n_128 GND GND efet w=7238 l=564
+ ad=0 pd=0 as=0 ps=0 
M4667 GND a7 n_128 GND efet w=4230 l=564
+ ad=0 pd=0 as=6.5033e+06 ps=19176 
M4668 adh6 dpc27_SBADH sb6 GND efet w=2068 l=752
+ ad=1.57369e+07 pd=40232 as=0 ps=0 
M4669 GND dpc29_0ADH17 adh6 GND efet w=2068 l=846
+ ad=0 pd=0 as=0 ps=0 
M4670 pchp0 pchp0 Vdd GND dfet w=940 l=1692
+ ad=4.23244e+06 pd=11844 as=0 ps=0 
M4671 n_835 n_919 n_1229 GND efet w=5499 l=611
+ ad=1.15928e+07 pd=32524 as=0 ps=0 
M4672 n_311 n_1010 GND GND efet w=2068 l=564
+ ad=1.02144e+07 pd=25380 as=0 ps=0 
M4673 n_835 dpc34_PCLC GND GND efet w=5217 l=611
+ ad=0 pd=0 as=0 ps=0 
M4674 n_1229 n_1229 Vdd GND dfet w=940 l=1598
+ ad=3.48138e+06 pd=10528 as=0 ps=0 
M4675 GND n_311 n_835 GND efet w=5123 l=611
+ ad=0 pd=0 as=0 ps=0 
M4676 dpc35_PCHC n_1010 GND GND efet w=5264 l=564
+ ad=0 pd=0 as=0 ps=0 
M4677 Vdd pchp1 pchp1 GND dfet w=846 l=1504
+ ad=0 pd=0 as=3.84366e+06 ps=11844 
M4678 Vdd npchp1 npchp1 GND dfet w=940 l=1504
+ ad=0 pd=0 as=9.29547e+06 ps=30644 
M4679 Vdd n_1486 n_1486 GND dfet w=846 l=1598
+ ad=0 pd=0 as=2.93355e+06 ps=8084 
M4680 n_1486 cclk n_126 GND efet w=1034 l=658
+ ad=7.72266e+06 pd=21432 as=1.46678e+06 ps=5828 
M4681 GND npchp1 pchp1 GND efet w=5734 l=564
+ ad=0 pd=0 as=0 ps=0 
M4682 pchp1 dpc33_PCHDB idb1 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M4683 n_1070 pch1 GND GND efet w=3196 l=564
+ ad=6.627e+06 pd=18612 as=0 ps=0 
M4684 GND n_126 npchp1 GND efet w=3948 l=564
+ ad=0 pd=0 as=7.50176e+06 ps=23124 
M4685 n_1486 n_200 GND GND efet w=3102 l=564
+ ad=0 pd=0 as=0 ps=0 
M4686 n_1538 n_919 n_1486 GND efet w=4042 l=564
+ ad=2.27969e+06 pd=9212 as=0 ps=0 
M4687 GND n_1070 n_1538 GND efet w=4042 l=564
+ ad=0 pd=0 as=0 ps=0 
M4688 dpc35_PCHC n_1070 GND GND efet w=5358 l=658
+ ad=0 pd=0 as=0 ps=0 
M4689 n_200 n_1070 GND GND efet w=2256 l=658
+ ad=9.96701e+06 pd=27636 as=0 ps=0 
M4690 GND n_919 n_200 GND efet w=2068 l=564
+ ad=0 pd=0 as=0 ps=0 
M4691 adh1 dpc32_PCHADH pchp1 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M4692 n_1070 n_1070 Vdd GND dfet w=940 l=1974
+ ad=1.45175e+07 pd=45120 as=0 ps=0 
M4693 n_200 n_200 Vdd GND dfet w=846 l=1316
+ ad=1.8264e+07 pd=59972 as=0 ps=0 
M4694 n_1202 n_1202 Vdd GND dfet w=940 l=1598
+ ad=1.12306e+07 pd=38352 as=0 ps=0 
M4695 GND n_1157 dpc41_DL_ADL GND efet w=9024 l=658
+ ad=0 pd=0 as=0 ps=0 
M4696 dpc42_DL_ADH n_1441 GND GND efet w=9259 l=611
+ ad=0 pd=0 as=0 ps=0 
M4697 dpc43_DL_DB n_1240 GND GND efet w=9729 l=611
+ ad=8.46489e+06 pd=22936 as=0 ps=0 
M4698 Vdd n_1566 dpc43_DL_DB GND dfet w=846 l=846
+ ad=0 pd=0 as=0 ps=0 
M4699 DBZ idb2 GND GND efet w=5076 l=564
+ ad=2.09678e+07 pd=55272 as=0 ps=0 
M4700 GND idb7 DBZ GND efet w=6392 l=564
+ ad=0 pd=0 as=0 ps=0 
M4701 DBZ idb6 GND GND efet w=4794 l=564
+ ad=0 pd=0 as=0 ps=0 
M4702 GND idb3 DBZ GND efet w=3619 l=517
+ ad=0 pd=0 as=0 ps=0 
M4703 Vdd n_206 n_206 GND dfet w=1316 l=658
+ ad=0 pd=0 as=4.98792e+07 ps=178600 
M4704 Pout0 Pout0 Vdd GND dfet w=846 l=940
+ ad=5.43414e+06 pd=20492 as=0 ps=0 
M4705 Pout1 Pout1 Vdd GND dfet w=940 l=940
+ ad=2.34154e+06 pd=8084 as=0 ps=0 
M4706 Pout0 H1x1 idb0 GND efet w=2256 l=752
+ ad=0 pd=0 as=0 ps=0 
M4707 Pout1 H1x1 idb1 GND efet w=2350 l=752
+ ad=0 pd=0 as=0 ps=0 
M4708 GND idb0 n_1224 GND efet w=6674 l=564
+ ad=0 pd=0 as=7.30737e+06 ps=20304 
M4709 n_243 idb1 GND GND efet w=6674 l=564
+ ad=6.71536e+06 pd=21056 as=0 ps=0 
M4710 n_1391 cclk pipeUNK15 GND efet w=1128 l=846
+ ad=0 pd=0 as=1.40492e+06 ps=6204 
M4711 GND pipeUNK15 H1x1 GND efet w=7849 l=517
+ ad=0 pd=0 as=1.03735e+07 ps=24064 
M4712 Vdd n_307 n_307 GND dfet w=846 l=1034
+ ad=0 pd=0 as=1.10803e+07 ps=41172 
M4713 n_90 n_90 Vdd GND dfet w=940 l=1034
+ ad=2.18779e+07 pd=79336 as=0 ps=0 
M4714 GND n_90 n_1433 GND efet w=3901 l=611
+ ad=0 pd=0 as=9.92283e+06 ps=31960 
M4715 GND n_620 n_922 GND efet w=7614 l=658
+ ad=0 pd=0 as=3.57858e+06 ps=16168 
M4716 n_922 n_270 BRtaken GND efet w=7614 l=564
+ ad=0 pd=0 as=9.43685e+06 ps=24440 
M4717 BRtaken BRtaken Vdd GND dfet w=846 l=846
+ ad=4.06633e+07 pd=148520 as=0 ps=0 
M4718 GND n_1115 BRtaken GND efet w=4841 l=705
+ ad=0 pd=0 as=0 ps=0 
M4719 n_1433 nop_branch_bit6 GND GND efet w=3854 l=658
+ ad=0 pd=0 as=0 ps=0 
M4720 n_1170 n_755 GND GND efet w=2350 l=658
+ ad=6.30007e+06 pd=16544 as=0 ps=0 
M4721 GND n_781 n_1170 GND efet w=2444 l=658
+ ad=0 pd=0 as=0 ps=0 
M4722 n_1170 n_1170 Vdd GND dfet w=940 l=1410
+ ad=6.89208e+06 pd=22184 as=0 ps=0 
M4723 n_580 nDBZ GND GND efet w=4606 l=564
+ ad=3.57858e+06 pd=12784 as=0 ps=0 
M4724 n_1224 n_1224 Vdd GND dfet w=940 l=1128
+ ad=2.57746e+07 pd=87232 as=0 ps=0 
M4725 GND n_937 dpc34_PCLC GND efet w=4559 l=611
+ ad=0 pd=0 as=0 ps=0 
M4726 n_1706 n_937 GND GND efet w=3760 l=658
+ ad=1.7672e+06 pd=8460 as=0 ps=0 
M4727 n_1500 dpc36_nIPC n_1706 GND efet w=3760 l=564
+ ad=8.09378e+06 pd=20680 as=0 ps=0 
M4728 Vdd n_1500 n_1500 GND dfet w=940 l=1504
+ ad=0 pd=0 as=2.81868e+06 ps=7708 
M4729 Vdd npclp0 npclp0 GND dfet w=940 l=1974
+ ad=0 pd=0 as=1.00024e+07 ps=32336 
M4730 n_526 cclk n_1500 GND efet w=1175 l=893
+ ad=1.47561e+06 pd=6956 as=0 ps=0 
M4731 GND n_937 n_1345 GND efet w=2303 l=611
+ ad=0 pd=0 as=1.02056e+07 ps=29892 
M4732 GND n_1345 n_1500 GND efet w=3102 l=564
+ ad=0 pd=0 as=0 ps=0 
M4733 Vdd pclp0 pclp0 GND dfet w=987 l=1457
+ ad=0 pd=0 as=3.69345e+06 ps=11656 
M4734 n_1345 dpc36_nIPC GND GND efet w=2068 l=564
+ ad=0 pd=0 as=0 ps=0 
M4735 npclp0 n_526 GND GND efet w=3290 l=658
+ ad=6.58282e+06 pd=21432 as=0 ps=0 
M4736 GND pcl0 n_937 GND efet w=3196 l=658
+ ad=0 pd=0 as=6.45028e+06 ps=17484 
M4737 pclp0 npclp0 GND GND efet w=5734 l=564
+ ad=1.44115e+07 pd=36848 as=0 ps=0 
M4738 Vdd cclk adl2 GND efet w=2068 l=564
+ ad=0 pd=0 as=0 ps=0 
M4739 Vdd n_293 n_293 GND dfet w=1034 l=1410
+ ad=0 pd=0 as=1.91564e+07 ps=65048 
M4740 n_1402 cclk npchp2 GND efet w=1034 l=752
+ ad=7.12182e+06 pd=21808 as=1.91741e+06 ps=7520 
M4741 pchp2 dpc31_PCHPCH pch2 GND efet w=1410 l=658
+ ad=1.40404e+07 pd=36660 as=5.3988e+06 ps=14852 
M4742 pch2 dpc30_ADHPCH adh2 GND efet w=1316 l=752
+ ad=0 pd=0 as=0 ps=0 
M4743 n_1592 dpc26_ACDB idb7 GND efet w=1316 l=752
+ ad=0 pd=0 as=0 ps=0 
M4744 idb7 dpc25_SBDB sb7 GND efet w=1974 l=658
+ ad=0 pd=0 as=0 ps=0 
M4745 sb7 dpc24_ACSB n_1592 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M4746 Vdd n_128 n_128 GND dfet w=940 l=1504
+ ad=0 pd=0 as=9.38383e+06 ps=26696 
M4747 adh7 dpc27_SBADH sb7 GND efet w=2068 l=752
+ ad=1.70358e+07 pd=44932 as=0 ps=0 
M4748 GND dpc29_0ADH17 adh7 GND efet w=2068 l=752
+ ad=0 pd=0 as=0 ps=0 
M4749 GND npchp2 pchp2 GND efet w=4042 l=564
+ ad=0 pd=0 as=0 ps=0 
M4750 n_1367 n_200 n_293 GND efet w=4042 l=658
+ ad=3.80832e+06 pd=11280 as=4.42684e+06 ps=13536 
M4751 GND n_1202 n_1367 GND efet w=4230 l=564
+ ad=0 pd=0 as=0 ps=0 
M4752 n_1265 pch2 GND GND efet w=4136 l=658
+ ad=4.08223e+06 pd=11844 as=0 ps=0 
M4753 Vdd n_1265 n_1265 GND dfet w=846 l=1880
+ ad=0 pd=0 as=9.71076e+06 ps=32148 
M4754 pchp2 dpc33_PCHDB idb2 GND efet w=1410 l=658
+ ad=0 pd=0 as=0 ps=0 
M4755 n_57 n_293 n_1402 GND efet w=5405 l=611
+ ad=1.09743e+07 pd=31772 as=0 ps=0 
M4756 n_1202 n_1265 GND GND efet w=2162 l=564
+ ad=1.06562e+07 pd=25568 as=0 ps=0 
M4757 Vdd n_1166 n_1166 GND dfet w=940 l=1504
+ ad=0 pd=0 as=1.20435e+07 ps=38916 
M4758 n_1345 n_1345 Vdd GND dfet w=940 l=1316
+ ad=1.74423e+07 pd=59220 as=0 ps=0 
M4759 n_937 n_937 Vdd GND dfet w=940 l=1880
+ ad=1.31921e+07 pd=40796 as=0 ps=0 
M4760 adl0 dpc38_PCLADL pclp0 GND efet w=1316 l=752
+ ad=0 pd=0 as=0 ps=0 
M4761 adl0 dpc40_ADLPCL pcl0 GND efet w=1316 l=752
+ ad=0 pd=0 as=4.20594e+06 ps=9024 
M4762 pcl0 dpc39_PCLPCL pclp0 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M4763 idb0 dpc37_PCLDB pclp0 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M4764 Vdd n_329 n_329 GND dfet w=940 l=1880
+ ad=0 pd=0 as=1.13101e+07 ps=32336 
M4765 GND pcl1 n_329 GND efet w=3901 l=611
+ ad=0 pd=0 as=3.54324e+06 ps=11468 
M4766 GND n_329 n_1166 GND efet w=2162 l=658
+ ad=0 pd=0 as=1.00465e+07 ps=25380 
M4767 n_1685 n_1166 GND GND efet w=4042 l=658
+ ad=4.0999e+06 pd=11280 as=0 ps=0 
M4768 Vdd n_1542 n_1542 GND dfet w=940 l=1222
+ ad=0 pd=0 as=1.92713e+07 ps=65236 
M4769 n_1542 n_1345 n_1685 GND efet w=4230 l=564
+ ad=5.32811e+06 pd=13724 as=0 ps=0 
M4770 npclp1 cclk n_1099 GND efet w=1034 l=752
+ ad=2.00577e+06 pd=8648 as=1.00112e+07 ps=27448 
M4771 adl1 dpc38_PCLADL pclp1 GND efet w=1316 l=658
+ ad=0 pd=0 as=1.35721e+07 ps=33088 
M4772 GND n_329 dpc34_PCLC GND efet w=5170 l=658
+ ad=0 pd=0 as=0 ps=0 
M4773 n_1568 n_1166 GND GND efet w=5264 l=658
+ ad=1.07357e+07 pd=31396 as=0 ps=0 
M4774 GND n_1345 n_1568 GND efet w=4982 l=658
+ ad=0 pd=0 as=0 ps=0 
M4775 n_1099 n_1542 n_1568 GND efet w=5452 l=564
+ ad=0 pd=0 as=0 ps=0 
M4776 pclp1 npclp1 GND GND efet w=5405 l=611
+ ad=0 pd=0 as=0 ps=0 
M4777 adl1 dpc40_ADLPCL pcl1 GND efet w=1316 l=846
+ ad=0 pd=0 as=4.08223e+06 ps=8836 
M4778 pcl1 dpc39_PCLPCL pclp1 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M4779 n_1099 n_1099 Vdd GND dfet w=940 l=1504
+ ad=3.48138e+06 pd=10528 as=0 ps=0 
M4780 idb1 dpc37_PCLDB pclp1 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M4781 adh2 dpc32_PCHADH pchp2 GND efet w=1316 l=752
+ ad=0 pd=0 as=0 ps=0 
M4782 adl3 cclk Vdd GND efet w=2162 l=658
+ ad=0 pd=0 as=0 ps=0 
M4783 pchp3 dpc31_PCHPCH pch3 GND efet w=1316 l=752
+ ad=1.46766e+07 pd=39292 as=5.26626e+06 ps=14664 
M4784 pch3 dpc30_ADHPCH adh3 GND efet w=1363 l=799
+ ad=0 pd=0 as=0 ps=0 
M4785 dpc23_SBAC cclk GND GND efet w=2444 l=658
+ ad=0 pd=0 as=0 ps=0 
M4786 dpc24_ACSB cclk GND GND efet w=2444 l=658
+ ad=0 pd=0 as=0 ps=0 
M4787 dpc26_ACDB cclk GND GND efet w=2538 l=658
+ ad=0 pd=0 as=0 ps=0 
M4788 pchp2 pchp2 Vdd GND dfet w=846 l=1786
+ ad=4.20594e+06 pd=11656 as=0 ps=0 
M4789 n_57 n_200 GND GND efet w=5123 l=611
+ ad=0 pd=0 as=0 ps=0 
M4790 n_1402 n_1402 Vdd GND dfet w=940 l=1598
+ ad=3.38419e+06 pd=10528 as=0 ps=0 
M4791 GND n_1202 n_57 GND efet w=5170 l=564
+ ad=0 pd=0 as=0 ps=0 
M4792 dpc35_PCHC n_1265 GND GND efet w=5076 l=564
+ ad=0 pd=0 as=0 ps=0 
M4793 Vdd pchp3 pchp3 GND dfet w=940 l=1504
+ ad=0 pd=0 as=3.94086e+06 ps=11656 
M4794 Vdd npchp3 npchp3 GND dfet w=940 l=1504
+ ad=0 pd=0 as=9.73727e+06 ps=30644 
M4795 Vdd n_207 n_207 GND dfet w=846 l=1504
+ ad=0 pd=0 as=2.70382e+06 ps=7896 
M4796 n_207 cclk n_1061 GND efet w=1081 l=799
+ ad=8.14679e+06 pd=22748 as=1.25471e+06 ps=6956 
M4797 GND npchp3 pchp3 GND efet w=5593 l=611
+ ad=0 pd=0 as=0 ps=0 
M4798 pchp3 dpc33_PCHDB idb3 GND efet w=1222 l=752
+ ad=0 pd=0 as=0 ps=0 
M4799 n_923 pch3 GND GND efet w=3102 l=564
+ ad=6.31774e+06 pd=18800 as=0 ps=0 
M4800 GND n_1061 npchp3 GND efet w=4230 l=658
+ ad=0 pd=0 as=7.79335e+06 ps=23500 
M4801 n_207 n_810 GND GND efet w=3102 l=564
+ ad=0 pd=0 as=0 ps=0 
M4802 n_356 n_293 n_207 GND efet w=4136 l=564
+ ad=2.72149e+06 pd=9588 as=0 ps=0 
M4803 GND n_923 n_356 GND efet w=4136 l=470
+ ad=0 pd=0 as=0 ps=0 
M4804 dpc35_PCHC n_923 GND GND efet w=5499 l=611
+ ad=0 pd=0 as=0 ps=0 
M4805 n_810 n_923 GND GND efet w=2397 l=611
+ ad=9.48986e+06 pd=29328 as=0 ps=0 
M4806 GND n_293 n_810 GND efet w=1974 l=564
+ ad=0 pd=0 as=0 ps=0 
M4807 adh3 dpc32_PCHADH pchp3 GND efet w=1316 l=752
+ ad=0 pd=0 as=0 ps=0 
M4808 pchp4 dpc31_PCHPCH pch4 GND efet w=1316 l=658
+ ad=1.40757e+07 pd=37036 as=5.53134e+06 ps=14852 
M4809 pch4 dpc30_ADHPCH adh4 GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M4810 n_923 n_923 Vdd GND dfet w=846 l=1880
+ ad=1.33335e+07 pd=44932 as=0 ps=0 
M4811 n_810 n_810 Vdd GND dfet w=940 l=1410
+ ad=7.17483e+06 pd=23688 as=0 ps=0 
M4812 n_83 n_83 Vdd GND dfet w=752 l=1504
+ ad=1.18491e+07 pd=37036 as=0 ps=0 
M4813 n_1657 cclk npchp4 GND efet w=1034 l=752
+ ad=9.91399e+06 pd=27448 as=1.69651e+06 ps=7708 
M4814 Vdd n_523 n_523 GND dfet w=940 l=1410
+ ad=0 pd=0 as=1.98898e+07 ps=64672 
M4815 GND npchp4 pchp4 GND efet w=5358 l=564
+ ad=0 pd=0 as=0 ps=0 
M4816 n_949 n_83 n_523 GND efet w=4042 l=658
+ ad=4.02038e+06 pd=10904 as=3.71112e+06 ps=12972 
M4817 GND dpc35_PCHC n_949 GND efet w=4183 l=611
+ ad=0 pd=0 as=0 ps=0 
M4818 n_1400 pch4 GND GND efet w=4042 l=658
+ ad=3.5344e+06 pd=11092 as=0 ps=0 
M4819 Vdd n_1400 n_1400 GND dfet w=846 l=1974
+ ad=0 pd=0 as=7.01578e+06 ps=20868 
M4820 pchp4 dpc33_PCHDB idb4 GND efet w=1316 l=752
+ ad=0 pd=0 as=0 ps=0 
M4821 n_1406 n_523 n_1657 GND efet w=5358 l=658
+ ad=1.05237e+07 pd=31772 as=0 ps=0 
M4822 n_83 n_1400 GND GND efet w=2068 l=564
+ ad=1.03293e+07 pd=25004 as=0 ps=0 
M4823 adh4 dpc32_PCHADH pchp4 GND efet w=1316 l=752
+ ad=0 pd=0 as=0 ps=0 
M4824 pchp5 dpc31_PCHPCH pch5 GND efet w=1316 l=658
+ ad=1.42525e+07 pd=39292 as=5.46065e+06 ps=14664 
M4825 pch5 dpc30_ADHPCH adh5 GND efet w=1222 l=658
+ ad=0 pd=0 as=0 ps=0 
M4826 pchp4 pchp4 Vdd GND dfet w=940 l=1692
+ ad=4.2943e+06 pd=11844 as=0 ps=0 
M4827 n_1406 n_83 GND GND efet w=5170 l=658
+ ad=0 pd=0 as=0 ps=0 
M4828 n_1657 n_1657 Vdd GND dfet w=940 l=1504
+ ad=3.29583e+06 pd=10340 as=0 ps=0 
M4829 GND dpc35_PCHC n_1406 GND efet w=5264 l=564
+ ad=0 pd=0 as=0 ps=0 
M4830 GND n_783 dpc34_PCLC GND efet w=5311 l=611
+ ad=0 pd=0 as=0 ps=0 
M4831 pclp1 pclp1 Vdd GND dfet w=940 l=1692
+ ad=4.3208e+06 pd=12032 as=0 ps=0 
M4832 n_1158 n_783 GND GND efet w=3666 l=564
+ ad=1.72302e+06 pd=8272 as=0 ps=0 
M4833 n_515 n_1542 n_1158 GND efet w=3666 l=658
+ ad=8.24399e+06 pd=22560 as=0 ps=0 
M4834 Vdd n_515 n_515 GND dfet w=846 l=1598
+ ad=0 pd=0 as=2.98657e+06 ps=7896 
M4835 Vdd npclp2 npclp2 GND dfet w=1034 l=1974
+ ad=0 pd=0 as=9.97584e+06 ps=32148 
M4836 GND n_783 n_1253 GND efet w=2303 l=611
+ ad=0 pd=0 as=9.78145e+06 ps=29516 
M4837 GND n_1253 n_515 GND efet w=3196 l=564
+ ad=0 pd=0 as=0 ps=0 
M4838 n_515 cclk n_1411 GND efet w=1128 l=752
+ ad=0 pd=0 as=1.41376e+06 ps=7144 
M4839 Vdd pclp2 pclp2 GND dfet w=940 l=1504
+ ad=0 pd=0 as=4.04689e+06 ps=11468 
M4840 n_1253 n_1542 GND GND efet w=2068 l=658
+ ad=0 pd=0 as=0 ps=0 
M4841 npclp2 n_1411 GND GND efet w=3102 l=658
+ ad=7.57245e+06 pd=21996 as=0 ps=0 
M4842 GND pcl2 n_783 GND efet w=3102 l=658
+ ad=0 pd=0 as=6.36192e+06 ps=16544 
M4843 pclp2 npclp2 GND GND efet w=5734 l=564
+ ad=1.48268e+07 pd=36848 as=0 ps=0 
M4844 Vdd n_163 n_163 GND dfet w=846 l=1504
+ ad=0 pd=0 as=1.25736e+07 ps=39104 
M4845 n_1253 n_1253 Vdd GND dfet w=846 l=1222
+ ad=1.67265e+07 pd=58844 as=0 ps=0 
M4846 n_783 n_783 Vdd GND dfet w=940 l=1880
+ ad=1.36958e+07 pd=44368 as=0 ps=0 
M4847 adl2 dpc38_PCLADL pclp2 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M4848 DBZ idb4 GND GND efet w=3572 l=564
+ ad=0 pd=0 as=0 ps=0 
M4849 GND idb5 DBZ GND efet w=4747 l=517
+ ad=0 pd=0 as=0 ps=0 
M4850 H1x1 H1x1 Vdd GND dfet w=1034 l=1504
+ ad=2.37247e+07 pd=68996 as=0 ps=0 
M4851 n_243 n_243 Vdd GND dfet w=940 l=1128
+ ad=1.95011e+07 pd=74636 as=0 ps=0 
M4852 DBZ idb0 GND GND efet w=4747 l=517
+ ad=0 pd=0 as=0 ps=0 
M4853 GND idb1 DBZ GND efet w=3572 l=376
+ ad=0 pd=0 as=0 ps=0 
M4854 Vdd DBZ DBZ GND dfet w=940 l=940
+ ad=0 pd=0 as=7.79335e+06 ps=23312 
M4855 n_566 n_755 n_580 GND efet w=3666 l=470
+ ad=1.18579e+07 pd=33464 as=0 ps=0 
M4856 n_661 n_1170 n_566 GND efet w=5499 l=611
+ ad=7.32504e+06 pd=17108 as=0 ps=0 
M4857 n_318 cclk pipeUNK14 GND efet w=1222 l=752
+ ad=1.41818e+07 pd=34216 as=1.3254e+06 ps=7520 
M4858 GND pipeUNK14 n_661 GND efet w=7614 l=470
+ ad=0 pd=0 as=0 ps=0 
M4859 GND p1 n_318 GND efet w=8131 l=611
+ ad=0 pd=0 as=0 ps=0 
M4860 n_1115 n_1115 Vdd GND dfet w=940 l=1128
+ ad=6.90975e+06 pd=21244 as=0 ps=0 
M4861 n_1115 n_270 GND GND efet w=3008 l=658
+ ad=5.66388e+06 pd=17108 as=0 ps=0 
M4862 GND n_201 n_1433 GND efet w=3854 l=658
+ ad=0 pd=0 as=0 ps=0 
M4863 Vdd n_1433 n_1433 GND dfet w=846 l=1034
+ ad=0 pd=0 as=1.24941e+07 ps=40796 
M4864 n_1371 n_1045 GND GND efet w=3807 l=611
+ ad=9.25129e+06 pd=32148 as=0 ps=0 
M4865 n_318 n_318 Vdd GND dfet w=846 l=1128
+ ad=2.73916e+07 pd=95692 as=0 ps=0 
M4866 Vdd n_1371 n_1371 GND dfet w=940 l=1128
+ ad=0 pd=0 as=1.17254e+07 ps=38352 
M4867 n_1115 n_620 GND GND efet w=3290 l=564
+ ad=0 pd=0 as=0 ps=0 
M4868 GND n_307 n_620 GND efet w=3760 l=564
+ ad=0 pd=0 as=1.78752e+07 ps=47564 
M4869 GND n_201 n_1371 GND efet w=3854 l=658
+ ad=0 pd=0 as=0 ps=0 
M4870 n_620 n_1433 GND GND efet w=3854 l=658
+ ad=0 pd=0 as=0 ps=0 
M4871 n_1371 n_846 GND GND efet w=3901 l=611
+ ad=0 pd=0 as=0 ps=0 
M4872 n_802 n_781 GND GND efet w=3666 l=564
+ ad=2.41223e+06 pd=8648 as=0 ps=0 
M4873 n_566 n_243 n_802 GND efet w=3666 l=470
+ ad=0 pd=0 as=0 ps=0 
M4874 Vdd n_566 n_566 GND dfet w=893 l=1269
+ ad=0 pd=0 as=3.01308e+06 ps=8648 
M4875 p1 cp1 n_566 GND efet w=1034 l=846
+ ad=1.35191e+06 pd=5452 as=0 ps=0 
M4876 GND n_1371 n_620 GND efet w=3854 l=658
+ ad=0 pd=0 as=0 ps=0 
M4877 n_620 n_620 Vdd GND dfet w=846 l=940
+ ad=1.7619e+07 pd=58656 as=0 ps=0 
M4878 GND n_1293 n_620 GND efet w=5170 l=658
+ ad=0 pd=0 as=0 ps=0 
M4879 GND n_318 n_1293 GND efet w=3854 l=658
+ ad=0 pd=0 as=1.08064e+07 ps=31584 
M4880 n_1579 cp1 notRnWprepad GND efet w=1128 l=752
+ ad=1.53746e+06 pd=7520 as=0 ps=0 
M4881 nDBE cclk GND GND efet w=11609 l=611
+ ad=1.34749e+07 pd=40796 as=0 ps=0 
M4882 GND n_251 n_1028 GND efet w=8460 l=564
+ ad=0 pd=0 as=6.93626e+06 ps=20868 
M4883 n_1028 n_1028 Vdd GND dfet w=846 l=658
+ ad=6.22054e+06 pd=21996 as=0 ps=0 
M4884 RnWstretched n_1028 Vdd GND dfet w=1974 l=470
+ ad=4.31374e+07 pd=86480 as=0 ps=0 
M4885 GND n_251 RnWstretched GND efet w=15416 l=564
+ ad=0 pd=0 as=0 ps=0 
M4886 n_251 n_221 GND GND efet w=9729 l=611
+ ad=1.46589e+07 pd=44180 as=0 ps=0 
M4887 GND nDBE n_251 GND efet w=12596 l=564
+ ad=0 pd=0 as=0 ps=0 
M4888 nDBZ DBZ GND GND efet w=5922 l=658
+ ad=8.12028e+06 pd=26508 as=0 ps=0 
M4889 RnWstretched n_251 GND GND efet w=15134 l=752
+ ad=0 pd=0 as=0 ps=0 
M4890 GND n_251 RnWstretched GND efet w=14758 l=658
+ ad=0 pd=0 as=0 ps=0 
M4891 GND n_962 nDBE GND efet w=11139 l=611
+ ad=0 pd=0 as=0 ps=0 
M4892 n_1585 cclk GND GND efet w=3290 l=658
+ ad=3.94086e+06 pd=14288 as=0 ps=0 
M4893 n_1585 n_1585 Vdd GND dfet w=846 l=1880
+ ad=7.45758e+06 pd=22748 as=0 ps=0 
M4894 GND n_1579 n_221 GND efet w=7097 l=611
+ ad=0 pd=0 as=8.04076e+06 ps=20868 
M4895 n_962 n_1585 GND GND efet w=3384 l=470
+ ad=5.65504e+06 pd=16544 as=0 ps=0 
M4896 n_1293 nop_branch_bit6 GND GND efet w=3807 l=611
+ ad=0 pd=0 as=0 ps=0 
M4897 Vdd n_1293 n_1293 GND dfet w=846 l=1034
+ ad=0 pd=0 as=1.11687e+07 ps=39856 
M4898 GND nop_branch_bit6 n_846 GND efet w=2538 l=658
+ ad=0 pd=0 as=8.5179e+06 ps=20680 
M4899 GND nop_branch_bit7 n_1293 GND efet w=3572 l=564
+ ad=0 pd=0 as=0 ps=0 
M4900 n_201 nop_branch_bit7 GND GND efet w=2538 l=564
+ ad=5.88478e+06 pd=17484 as=0 ps=0 
M4901 n_846 n_846 Vdd GND dfet w=940 l=1598
+ ad=1.63996e+07 pd=52640 as=0 ps=0 
M4902 n_201 n_201 Vdd GND dfet w=846 l=1504
+ ad=2.61899e+07 pd=90052 as=0 ps=0 
M4903 n_221 n_221 Vdd GND dfet w=940 l=1128
+ ad=1.51979e+07 pd=49068 as=0 ps=0 
M4904 nDBZ nDBZ Vdd GND dfet w=1034 l=1034
+ ad=1.47384e+07 pd=57716 as=0 ps=0 
M4905 n_719 dpc41_DL_ADL adl0 GND efet w=5922 l=658
+ ad=1.73097e+07 pd=47000 as=0 ps=0 
M4906 adl2 dpc40_ADLPCL pcl2 GND efet w=1316 l=658
+ ad=0 pd=0 as=4.32964e+06 ps=9212 
M4907 pcl2 dpc39_PCLPCL pclp2 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M4908 idb2 dpc37_PCLDB pclp2 GND efet w=1222 l=752
+ ad=0 pd=0 as=0 ps=0 
M4909 Vdd n_249 n_249 GND dfet w=940 l=1974
+ ad=0 pd=0 as=1.1204e+07 ps=31960 
M4910 GND pcl3 n_249 GND efet w=3948 l=564
+ ad=0 pd=0 as=4.35615e+06 ps=11468 
M4911 GND n_249 n_163 GND efet w=2068 l=658
+ ad=0 pd=0 as=1.04088e+07 ps=25192 
M4912 n_1498 n_163 GND GND efet w=4042 l=658
+ ad=4.10874e+06 pd=11280 as=0 ps=0 
M4913 Vdd n_1184 n_1184 GND dfet w=940 l=1316
+ ad=0 pd=0 as=1.88649e+07 ps=67680 
M4914 n_1184 n_1253 n_1498 GND efet w=4042 l=564
+ ad=4.9835e+06 pd=12972 as=0 ps=0 
M4915 npclp3 cclk n_1631 GND efet w=1128 l=658
+ ad=1.90858e+06 pd=8460 as=1.04795e+07 ps=27824 
M4916 GND n_249 dpc34_PCLC GND efet w=5170 l=658
+ ad=0 pd=0 as=0 ps=0 
M4917 n_903 n_163 GND GND efet w=5311 l=705
+ ad=1.14868e+07 pd=31960 as=0 ps=0 
M4918 GND n_1253 n_903 GND efet w=5076 l=470
+ ad=0 pd=0 as=0 ps=0 
M4919 n_1631 n_1184 n_903 GND efet w=5358 l=564
+ ad=0 pd=0 as=0 ps=0 
M4920 pclp3 npclp3 GND GND efet w=5358 l=564
+ ad=1.41818e+07 pd=34216 as=0 ps=0 
M4921 adl3 dpc38_PCLADL pclp3 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M4922 adl3 dpc40_ADLPCL pcl3 GND efet w=1316 l=752
+ ad=0 pd=0 as=4.14408e+06 ps=9024 
M4923 pcl3 dpc39_PCLPCL pclp3 GND efet w=1222 l=658
+ ad=0 pd=0 as=0 ps=0 
M4924 n_1631 n_1631 Vdd GND dfet w=940 l=1504
+ ad=3.56091e+06 pd=10340 as=0 ps=0 
M4925 idb3 dpc37_PCLDB pclp3 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M4926 pclp3 pclp3 Vdd GND dfet w=940 l=1786
+ ad=4.20594e+06 pd=12032 as=0 ps=0 
M4927 GND n_1643 dpc34_PCLC GND efet w=5358 l=564
+ ad=0 pd=0 as=0 ps=0 
M4928 n_766 n_1643 GND GND efet w=3666 l=564
+ ad=2.06762e+06 pd=8460 as=0 ps=0 
M4929 n_474 n_1184 n_766 GND efet w=3666 l=564
+ ad=8.36769e+06 pd=22560 as=0 ps=0 
M4930 Vdd n_474 n_474 GND dfet w=846 l=1410
+ ad=0 pd=0 as=2.50942e+06 ps=7520 
M4931 Vdd npclp4 npclp4 GND dfet w=846 l=1880
+ ad=0 pd=0 as=1.01526e+07 ps=31960 
M4932 GND n_1643 n_410 GND efet w=2350 l=564
+ ad=0 pd=0 as=9.98468e+06 ps=30080 
M4933 GND n_410 n_474 GND efet w=3196 l=564
+ ad=0 pd=0 as=0 ps=0 
M4934 n_474 cclk n_15 GND efet w=1128 l=752
+ ad=0 pd=0 as=1.53746e+06 ps=6956 
M4935 Vdd pclp4 pclp4 GND dfet w=846 l=1504
+ ad=0 pd=0 as=3.44604e+06 ps=10716 
M4936 n_410 n_1184 GND GND efet w=1974 l=564
+ ad=0 pd=0 as=0 ps=0 
M4937 npclp4 n_15 GND GND efet w=3102 l=564
+ ad=6.79488e+06 pd=21620 as=0 ps=0 
M4938 GND pcl4 n_1643 GND efet w=3102 l=658
+ ad=0 pd=0 as=6.57398e+06 ps=16920 
M4939 pclp4 npclp4 GND GND efet w=5687 l=611
+ ad=1.44292e+07 pd=36848 as=0 ps=0 
M4940 Vdd n_392 n_392 GND dfet w=846 l=1504
+ ad=0 pd=0 as=1.18491e+07 ps=38728 
M4941 Vdd pchp5 pchp5 GND dfet w=940 l=1410
+ ad=0 pd=0 as=3.79064e+06 ps=11468 
M4942 Vdd npchp5 npchp5 GND dfet w=940 l=1504
+ ad=0 pd=0 as=9.8433e+06 ps=31020 
M4943 Vdd n_875 n_875 GND dfet w=846 l=1598
+ ad=0 pd=0 as=2.88054e+06 ps=7896 
M4944 n_875 cclk n_469 GND efet w=1128 l=752
+ ad=8.01425e+06 pd=22372 as=1.43143e+06 ps=6580 
M4945 GND npchp5 pchp5 GND efet w=5781 l=611
+ ad=0 pd=0 as=0 ps=0 
M4946 pchp5 dpc33_PCHDB idb5 GND efet w=1128 l=752
+ ad=0 pd=0 as=0 ps=0 
M4947 n_499 pch5 GND GND efet w=3196 l=658
+ ad=6.22054e+06 pd=18800 as=0 ps=0 
M4948 GND n_469 npchp5 GND efet w=3948 l=658
+ ad=0 pd=0 as=7.17483e+06 ps=23124 
M4949 n_875 n_743 GND GND efet w=3102 l=564
+ ad=0 pd=0 as=0 ps=0 
M4950 n_1659 n_523 n_875 GND efet w=4136 l=564
+ ad=2.3327e+06 pd=9400 as=0 ps=0 
M4951 GND n_499 n_1659 GND efet w=4136 l=564
+ ad=0 pd=0 as=0 ps=0 
M4952 GND n_523 n_743 GND efet w=2068 l=564
+ ad=0 pd=0 as=9.7196e+06 ps=28012 
M4953 GND n_499 n_743 GND efet w=2726 l=564
+ ad=0 pd=0 as=0 ps=0 
M4954 adh5 dpc32_PCHADH pchp5 GND efet w=1222 l=658
+ ad=0 pd=0 as=0 ps=0 
M4955 pchp6 dpc31_PCHPCH pch6 GND efet w=1316 l=658
+ ad=1.41023e+07 pd=37788 as=5.10721e+06 ps=14664 
M4956 pch6 dpc30_ADHPCH adh6 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M4957 n_499 n_499 Vdd GND dfet w=846 l=1880
+ ad=1.48622e+07 pd=50196 as=0 ps=0 
M4958 n_410 n_410 Vdd GND dfet w=846 l=1222
+ ad=1.80696e+07 pd=59032 as=0 ps=0 
M4959 n_1643 n_1643 Vdd GND dfet w=940 l=1974
+ ad=1.36781e+07 pd=45120 as=0 ps=0 
M4960 adl4 dpc38_PCLADL pclp4 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M4961 adl4 dpc40_ADLPCL pcl4 GND efet w=1316 l=658
+ ad=0 pd=0 as=4.32964e+06 ps=9212 
M4962 pcl4 dpc39_PCLPCL pclp4 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M4963 idb4 dpc37_PCLDB pclp4 GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M4964 Vdd n_386 n_386 GND dfet w=1034 l=1974
+ ad=0 pd=0 as=1.01437e+07 ps=32148 
M4965 GND pcl5 n_386 GND efet w=3948 l=658
+ ad=0 pd=0 as=3.71112e+06 ps=11844 
M4966 GND n_386 n_392 GND efet w=2162 l=564
+ ad=0 pd=0 as=1.02056e+07 ps=25380 
M4967 n_814 n_392 GND GND efet w=4042 l=658
+ ad=3.76414e+06 pd=11092 as=0 ps=0 
M4968 Vdd n_344 n_344 GND dfet w=940 l=1222
+ ad=0 pd=0 as=1.79636e+07 ps=64860 
M4969 n_344 n_410 n_814 GND efet w=4230 l=658
+ ad=5.22208e+06 pd=13724 as=0 ps=0 
M4970 npclp5 cclk n_1073 GND efet w=1128 l=752
+ ad=1.80254e+06 pd=8272 as=1.03823e+07 ps=27636 
M4971 n_743 n_743 Vdd GND dfet w=940 l=1316
+ ad=1.83347e+07 pd=59596 as=0 ps=0 
M4972 n_1488 n_1488 Vdd GND dfet w=846 l=1504
+ ad=1.16724e+07 pd=37976 as=0 ps=0 
M4973 n_1192 cclk npchp6 GND efet w=1128 l=658
+ ad=9.64891e+06 pd=27072 as=1.70535e+06 ps=7896 
M4974 Vdd n_609 n_609 GND dfet w=846 l=1316
+ ad=0 pd=0 as=1.89179e+07 ps=64672 
M4975 GND npchp6 pchp6 GND efet w=5405 l=611
+ ad=0 pd=0 as=0 ps=0 
M4976 n_545 n_743 n_609 GND efet w=4136 l=658
+ ad=3.74646e+06 pd=11280 as=4.17059e+06 ps=13536 
M4977 GND n_1488 n_545 GND efet w=4136 l=564
+ ad=0 pd=0 as=0 ps=0 
M4978 n_278 pch6 GND GND efet w=3948 l=658
+ ad=3.60509e+06 pd=11092 as=0 ps=0 
M4979 Vdd n_278 n_278 GND dfet w=940 l=1880
+ ad=0 pd=0 as=6.90975e+06 ps=20868 
M4980 pchp6 dpc33_PCHDB idb6 GND efet w=1222 l=658
+ ad=0 pd=0 as=0 ps=0 
M4981 n_1547 n_609 n_1192 GND efet w=5311 l=611
+ ad=1.06916e+07 pd=32148 as=0 ps=0 
M4982 n_1488 n_278 GND GND efet w=2162 l=564
+ ad=9.80796e+06 pd=25380 as=0 ps=0 
M4983 GND n_386 dpc34_PCLC GND efet w=5170 l=564
+ ad=0 pd=0 as=0 ps=0 
M4984 n_557 n_392 GND GND efet w=5264 l=564
+ ad=1.07357e+07 pd=31584 as=0 ps=0 
M4985 GND n_410 n_557 GND efet w=4888 l=658
+ ad=0 pd=0 as=0 ps=0 
M4986 n_1073 n_344 n_557 GND efet w=5452 l=564
+ ad=0 pd=0 as=0 ps=0 
M4987 pclp5 npclp5 GND GND efet w=5452 l=564
+ ad=1.36958e+07 pd=33088 as=0 ps=0 
M4988 adl5 dpc38_PCLADL pclp5 GND efet w=1316 l=752
+ ad=0 pd=0 as=0 ps=0 
M4989 adl5 dpc40_ADLPCL pcl5 GND efet w=1316 l=752
+ ad=0 pd=0 as=4.08223e+06 ps=8836 
M4990 pcl5 dpc39_PCLPCL pclp5 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M4991 GND n_232 dpc34_PCLC GND efet w=5264 l=658
+ ad=0 pd=0 as=0 ps=0 
M4992 n_1073 n_1073 Vdd GND dfet w=846 l=1504
+ ad=3.48138e+06 pd=10528 as=0 ps=0 
M4993 idb5 dpc37_PCLDB pclp5 GND efet w=1316 l=564
+ ad=0 pd=0 as=0 ps=0 
M4994 pclp5 pclp5 Vdd GND dfet w=846 l=1692
+ ad=4.28546e+06 pd=12032 as=0 ps=0 
M4995 n_585 n_232 GND GND efet w=3666 l=658
+ ad=1.72302e+06 pd=8272 as=0 ps=0 
M4996 n_20 n_344 n_585 GND efet w=3666 l=564
+ ad=8.62394e+06 pd=22560 as=0 ps=0 
M4997 Vdd n_20 n_20 GND dfet w=940 l=1598
+ ad=0 pd=0 as=2.97773e+06 ps=7896 
M4998 Vdd npclp6 npclp6 GND dfet w=940 l=1880
+ ad=0 pd=0 as=9.7196e+06 ps=31584 
M4999 adh6 dpc32_PCHADH pchp6 GND efet w=1222 l=658
+ ad=0 pd=0 as=0 ps=0 
M5000 pchp7 dpc31_PCHPCH pch7 GND efet w=1316 l=752
+ ad=1.47561e+07 pd=39856 as=5.29276e+06 ps=14476 
M5001 pch7 dpc30_ADHPCH adh7 GND efet w=1222 l=658
+ ad=0 pd=0 as=0 ps=0 
M5002 pchp6 pchp6 Vdd GND dfet w=1034 l=1692
+ ad=4.01154e+06 pd=11280 as=0 ps=0 
M5003 n_1547 n_743 GND GND efet w=5217 l=611
+ ad=0 pd=0 as=0 ps=0 
M5004 n_1192 n_1192 Vdd GND dfet w=940 l=1504
+ ad=3.48138e+06 pd=10528 as=0 ps=0 
M5005 GND n_1488 n_1547 GND efet w=5123 l=611
+ ad=0 pd=0 as=0 ps=0 
M5006 Vdd pchp7 pchp7 GND dfet w=940 l=1410
+ ad=0 pd=0 as=3.77297e+06 ps=11468 
M5007 Vdd npchp7 npchp7 GND dfet w=940 l=1504
+ ad=0 pd=0 as=9.66658e+06 ps=30832 
M5008 Vdd n_1209 n_1209 GND dfet w=846 l=1598
+ ad=0 pd=0 as=2.88054e+06 ps=7896 
M5009 n_1209 cclk n_663 GND efet w=1034 l=752
+ ad=7.92589e+06 pd=21996 as=1.36958e+06 ps=7332 
M5010 GND npchp7 pchp7 GND efet w=5687 l=611
+ ad=0 pd=0 as=0 ps=0 
M5011 pchp7 dpc33_PCHDB idb7 GND efet w=1410 l=752
+ ad=0 pd=0 as=0 ps=0 
M5012 n_453 pch7 GND GND efet w=3008 l=564
+ ad=6.07917e+06 pd=18612 as=0 ps=0 
M5013 GND n_663 npchp7 GND efet w=3948 l=564
+ ad=0 pd=0 as=7.93473e+06 ps=23312 
M5014 n_1209 n_1213 GND GND efet w=3102 l=658
+ ad=0 pd=0 as=0 ps=0 
M5015 n_1264 n_609 n_1209 GND efet w=4136 l=564
+ ad=2.3327e+06 pd=9400 as=0 ps=0 
M5016 GND n_453 n_1264 GND efet w=4136 l=564
+ ad=0 pd=0 as=0 ps=0 
M5017 GND n_609 n_1213 GND efet w=2162 l=564
+ ad=0 pd=0 as=1.03293e+07 ps=29328 
M5018 n_1213 n_453 GND GND efet w=2068 l=564
+ ad=0 pd=0 as=0 ps=0 
M5019 GND n_232 n_1316 GND efet w=2256 l=658
+ ad=0 pd=0 as=1.04353e+07 ps=27448 
M5020 GND n_1316 n_20 GND efet w=3196 l=564
+ ad=0 pd=0 as=0 ps=0 
M5021 n_20 cclk n_993 GND efet w=1222 l=846
+ ad=0 pd=0 as=1.51979e+06 ps=6956 
M5022 Vdd pclp6 pclp6 GND dfet w=940 l=1504
+ ad=0 pd=0 as=3.72879e+06 ps=10904 
M5023 n_1316 n_344 GND GND efet w=1974 l=564
+ ad=0 pd=0 as=0 ps=0 
M5024 npclp6 n_993 GND GND efet w=3196 l=658
+ ad=6.96277e+06 pd=21432 as=0 ps=0 
M5025 GND pcl6 n_232 GND efet w=3102 l=658
+ ad=0 pd=0 as=6.36192e+06 ps=16544 
M5026 pclp6 npclp6 GND GND efet w=5734 l=564
+ ad=1.51361e+07 pd=37036 as=0 ps=0 
M5027 Vdd n_715 n_715 GND dfet w=940 l=1504
+ ad=0 pd=0 as=1.21672e+07 ps=38916 
M5028 n_1316 n_1316 Vdd GND dfet w=846 l=1222
+ ad=1.80166e+07 pd=59220 as=0 ps=0 
M5029 n_232 n_232 Vdd GND dfet w=940 l=1974
+ ad=1.44204e+07 pd=43804 as=0 ps=0 
M5030 adl6 dpc38_PCLADL pclp6 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M5031 nDBE nDBE Vdd GND dfet w=846 l=752
+ ad=1.34396e+07 pd=45120 as=0 ps=0 
M5032 RnWstretched n_251 GND GND efet w=16356 l=658
+ ad=0 pd=0 as=0 ps=0 
M5033 n_251 n_221 GND GND efet w=3008 l=658
+ ad=0 pd=0 as=0 ps=0 
M5034 n_962 n_962 Vdd GND dfet w=846 l=1222
+ ad=1.10185e+07 pd=35908 as=0 ps=0 
M5035 Vdd n_251 n_251 GND dfet w=1692 l=658
+ ad=0 pd=0 as=5.32899e+07 ps=172396 
M5036 Vdd n_1687 n_1687 GND dfet w=846 l=1504
+ ad=0 pd=0 as=2.84519e+06 ps=7896 
M5037 idl0 idl0 Vdd GND dfet w=940 l=1598
+ ad=2.97773e+06 pd=7896 as=0 ps=0 
M5038 n_1687 cp1 notdor0 GND efet w=1175 l=799
+ ad=7.96124e+06 pd=25380 as=1.89974e+06 ps=7896 
M5039 idl0 cp1 n_719 GND efet w=5781 l=705
+ ad=1.23085e+07 pd=31396 as=0 ps=0 
M5040 n_719 dpc42_DL_ADH adh0 GND efet w=4089 l=705
+ ad=0 pd=0 as=0 ps=0 
M5041 GND idb0 n_1687 GND efet w=4371 l=611
+ ad=0 pd=0 as=0 ps=0 
M5042 dor0 notdor0 GND GND efet w=6486 l=564
+ ad=7.54594e+06 pd=23688 as=0 ps=0 
M5043 GND notidl0 idl0 GND efet w=3572 l=564
+ ad=0 pd=0 as=0 ps=0 
M5044 Vdd n_718 n_718 GND dfet w=940 l=658
+ ad=0 pd=0 as=2.26202e+06 ps=9212 
M5045 db0 GND GND GND efet w=5076 l=658
+ ad=2.31503e+08 pd=409652 as=0 ps=0 
M5046 n_718 cclk notidl0 GND efet w=1316 l=752
+ ad=1.52244e+07 pd=35720 as=2.06762e+06 ps=7708 
M5047 GND db0 n_718 GND efet w=12596 l=564
+ ad=0 pd=0 as=0 ps=0 
M5048 n_87 dpc41_DL_ADL adl1 GND efet w=5828 l=658
+ ad=1.72479e+07 pd=47188 as=0 ps=0 
M5049 idb0 dpc43_DL_DB n_719 GND efet w=4042 l=658
+ ad=0 pd=0 as=0 ps=0 
M5050 GND notidl0 idl0 GND efet w=3149 l=517
+ ad=0 pd=0 as=0 ps=0 
M5051 db0 n_1325 Vdd GND efet w=59878 l=658
+ ad=0 pd=0 as=0 ps=0 
M5052 n_1325 RnWstretched GND GND efet w=14241 l=611
+ ad=2.07204e+07 pd=51512 as=0 ps=0 
M5053 GND RnWstretched n_1325 GND efet w=14570 l=564
+ ad=0 pd=0 as=0 ps=0 
M5054 idl0 notidl0 GND GND efet w=4653 l=611
+ ad=0 pd=0 as=0 ps=0 
M5055 GND RnWstretched n_769 GND efet w=6815 l=611
+ ad=0 pd=0 as=7.05996e+06 ps=20116 
M5056 GND n_769 n_1325 GND efet w=12972 l=564
+ ad=0 pd=0 as=0 ps=0 
M5057 Vdd cclk idb0 GND efet w=2068 l=752
+ ad=0 pd=0 as=0 ps=0 
M5058 n_1325 dor0 Vdd GND dfet w=1504 l=658
+ ad=0 pd=0 as=0 ps=0 
M5059 Vdd n_769 n_769 GND dfet w=940 l=752
+ ad=0 pd=0 as=1.29271e+07 ps=46248 
M5060 n_1072 n_769 Vdd GND dfet w=1598 l=564
+ ad=2.17101e+07 pd=51888 as=0 ps=0 
M5061 GND RnWstretched n_1072 GND efet w=8883 l=611
+ ad=0 pd=0 as=0 ps=0 
M5062 GND RnWstretched n_1072 GND efet w=18894 l=564
+ ad=0 pd=0 as=0 ps=0 
M5063 n_1072 dor0 GND GND efet w=13959 l=611
+ ad=0 pd=0 as=0 ps=0 
M5064 n_769 dor0 GND GND efet w=5546 l=564
+ ad=0 pd=0 as=0 ps=0 
M5065 db0 n_1072 GND GND efet w=10481 l=611
+ ad=0 pd=0 as=0 ps=0 
M5066 GND n_1072 db0 GND efet w=20304 l=564
+ ad=0 pd=0 as=0 ps=0 
M5067 db0 n_1072 GND GND efet w=20022 l=564
+ ad=0 pd=0 as=0 ps=0 
M5068 db0 n_1325 Vdd GND efet w=59596 l=658
+ ad=0 pd=0 as=0 ps=0 
M5069 GND n_1072 db0 GND efet w=1034 l=564
+ ad=0 pd=0 as=0 ps=0 
M5070 dor0 dor0 Vdd GND dfet w=940 l=1034
+ ad=1.88914e+07 pd=63168 as=0 ps=0 
M5071 Vdd n_1474 n_1474 GND dfet w=846 l=1504
+ ad=0 pd=0 as=2.79218e+06 ps=7708 
M5072 idl1 idl1 Vdd GND dfet w=846 l=1598
+ ad=2.80101e+06 pd=7896 as=0 ps=0 
M5073 n_1474 cp1 notdor1 GND efet w=1034 l=846
+ ad=7.57245e+06 pd=24628 as=1.90858e+06 ps=7708 
M5074 idl1 cp1 n_87 GND efet w=5922 l=658
+ ad=1.19021e+07 pd=31772 as=0 ps=0 
M5075 Vdd cclk adh3 GND efet w=2068 l=564
+ ad=0 pd=0 as=0 ps=0 
M5076 adl4 cclk Vdd GND efet w=2068 l=658
+ ad=0 pd=0 as=0 ps=0 
M5077 adl6 dpc40_ADLPCL pcl6 GND efet w=1316 l=752
+ ad=0 pd=0 as=4.25895e+06 ps=9024 
M5078 pcl6 dpc39_PCLPCL pclp6 GND efet w=1410 l=752
+ ad=0 pd=0 as=0 ps=0 
M5079 idb6 dpc37_PCLDB pclp6 GND efet w=1222 l=658
+ ad=0 pd=0 as=0 ps=0 
M5080 Vdd n_641 n_641 GND dfet w=940 l=1974
+ ad=0 pd=0 as=1.07181e+07 ps=30268 
M5081 GND pcl7 n_641 GND efet w=4042 l=564
+ ad=0 pd=0 as=4.18826e+06 ps=11280 
M5082 GND n_641 n_715 GND efet w=2162 l=658
+ ad=0 pd=0 as=1.04618e+07 ps=25944 
M5083 n_426 n_715 GND GND efet w=4136 l=658
+ ad=4.25012e+06 pd=11468 as=0 ps=0 
M5084 Vdd n_1386 n_1386 GND dfet w=940 l=1410
+ ad=0 pd=0 as=9.89632e+06 ps=30268 
M5085 n_1386 n_1316 n_426 GND efet w=4324 l=564
+ ad=4.42684e+06 pd=13536 as=0 ps=0 
M5086 npclp7 cclk n_484 GND efet w=1034 l=752
+ ad=1.91741e+06 pd=8460 as=9.4987e+06 ps=27448 
M5087 adh7 dpc32_PCHADH pchp7 GND efet w=1316 l=752
+ ad=0 pd=0 as=0 ps=0 
M5088 n_453 n_453 Vdd GND dfet w=846 l=1974
+ ad=9.86098e+06 pd=31396 as=0 ps=0 
M5089 n_1213 n_1213 Vdd GND dfet w=940 l=1316
+ ad=7.2897e+06 pd=23876 as=0 ps=0 
M5090 dpc34_PCLC dpc34_PCLC Vdd GND dfet w=1034 l=564
+ ad=8.69728e+07 pd=328812 as=0 ps=0 
M5091 GND n_641 dpc34_PCLC GND efet w=4418 l=658
+ ad=0 pd=0 as=0 ps=0 
M5092 n_914 n_715 GND GND efet w=5311 l=611
+ ad=1.05679e+07 pd=31208 as=0 ps=0 
M5093 GND n_1316 n_914 GND efet w=4935 l=611
+ ad=0 pd=0 as=0 ps=0 
M5094 n_484 n_1386 n_914 GND efet w=5405 l=611
+ ad=0 pd=0 as=0 ps=0 
M5095 pclp7 npclp7 GND GND efet w=5452 l=658
+ ad=1.36339e+07 pd=36096 as=0 ps=0 
M5096 adl7 dpc38_PCLADL pclp7 GND efet w=1316 l=752
+ ad=0 pd=0 as=0 ps=0 
M5097 adl7 dpc40_ADLPCL pcl7 GND efet w=1316 l=752
+ ad=0 pd=0 as=4.01154e+06 ps=8648 
M5098 pcl7 dpc39_PCLPCL pclp7 GND efet w=1316 l=752
+ ad=0 pd=0 as=0 ps=0 
M5099 n_484 n_484 Vdd GND dfet w=940 l=1504
+ ad=3.48138e+06 pd=10528 as=0 ps=0 
M5100 idb7 dpc37_PCLDB pclp7 GND efet w=1316 l=658
+ ad=0 pd=0 as=0 ps=0 
M5101 pclp7 pclp7 Vdd GND dfet w=940 l=1692
+ ad=4.18826e+06 pd=11844 as=0 ps=0 
M5102 GND cclk dpc30_ADHPCH GND efet w=2444 l=752
+ ad=0 pd=0 as=0 ps=0 
M5103 n_87 dpc42_DL_ADH adh1 GND efet w=4089 l=705
+ ad=0 pd=0 as=0 ps=0 
M5104 GND idb1 n_1474 GND efet w=4230 l=564
+ ad=0 pd=0 as=0 ps=0 
M5105 dor1 notdor1 GND GND efet w=6533 l=611
+ ad=7.46642e+06 pd=23500 as=0 ps=0 
M5106 GND notidl1 idl1 GND efet w=3478 l=658
+ ad=0 pd=0 as=0 ps=0 
M5107 Vdd n_213 n_213 GND dfet w=940 l=658
+ ad=0 pd=0 as=2.17366e+06 ps=9400 
M5108 db0 n_1072 GND GND efet w=19834 l=564
+ ad=0 pd=0 as=0 ps=0 
M5109 GND n_1072 db0 GND efet w=1034 l=564
+ ad=0 pd=0 as=0 ps=0 
M5110 n_213 cclk notidl1 GND efet w=1316 l=752
+ ad=1.62582e+07 pd=36660 as=2.0853e+06 ps=7332 
M5111 GND db1 n_213 GND efet w=12690 l=564
+ ad=0 pd=0 as=0 ps=0 
M5112 n_1424 dpc41_DL_ADL adl2 GND efet w=5828 l=564
+ ad=1.83082e+07 pd=47564 as=0 ps=0 
M5113 idb1 dpc43_DL_DB n_87 GND efet w=4042 l=658
+ ad=0 pd=0 as=0 ps=0 
M5114 GND notidl1 idl1 GND efet w=3149 l=611
+ ad=0 pd=0 as=0 ps=0 
M5115 n_798 RnWstretched GND GND efet w=14241 l=611
+ ad=2.02433e+07 pd=51324 as=0 ps=0 
M5116 n_798 RnWstretched GND GND efet w=14382 l=564
+ ad=0 pd=0 as=0 ps=0 
M5117 idl1 notidl1 GND GND efet w=4653 l=611
+ ad=0 pd=0 as=0 ps=0 
M5118 GND n_288 n_798 GND efet w=13066 l=564
+ ad=0 pd=0 as=0 ps=0 
M5119 GND RnWstretched n_288 GND efet w=6862 l=658
+ ad=0 pd=0 as=6.80372e+06 ps=19552 
M5120 Vdd cclk idb1 GND efet w=1974 l=846
+ ad=0 pd=0 as=0 ps=0 
M5121 n_798 dor1 Vdd GND dfet w=1598 l=658
+ ad=0 pd=0 as=0 ps=0 
M5122 Vdd n_288 n_288 GND dfet w=940 l=752
+ ad=0 pd=0 as=1.33159e+07 ps=46060 
M5123 db0 n_1072 GND GND efet w=14805 l=611
+ ad=0 pd=0 as=0 ps=0 
M5124 db0 n_1072 GND GND efet w=12220 l=658
+ ad=0 pd=0 as=0 ps=0 
M5125 GND n_794 db1 GND efet w=14758 l=658
+ ad=0 pd=0 as=2.35373e+08 ps=412284 
M5126 GND n_794 db1 GND efet w=12220 l=658
+ ad=0 pd=0 as=0 ps=0 
M5127 db1 n_798 Vdd GND efet w=60019 l=611
+ ad=0 pd=0 as=0 ps=0 
M5128 n_794 n_288 Vdd GND dfet w=1598 l=564
+ ad=2.21695e+07 pd=52452 as=0 ps=0 
M5129 GND RnWstretched n_794 GND efet w=8930 l=564
+ ad=0 pd=0 as=0 ps=0 
M5130 db1 n_794 GND GND efet w=26414 l=564
+ ad=0 pd=0 as=0 ps=0 
M5131 GND RnWstretched n_794 GND efet w=18847 l=611
+ ad=0 pd=0 as=0 ps=0 
M5132 n_794 dor1 GND GND efet w=14053 l=611
+ ad=0 pd=0 as=0 ps=0 
M5133 n_288 dor1 GND GND efet w=5452 l=564
+ ad=0 pd=0 as=0 ps=0 
M5134 GND n_794 db1 GND efet w=1128 l=564
+ ad=0 pd=0 as=0 ps=0 
M5135 dor1 dor1 Vdd GND dfet w=846 l=1128
+ ad=1.92006e+07 pd=63732 as=0 ps=0 
M5136 Vdd n_1376 n_1376 GND dfet w=940 l=1504
+ ad=0 pd=0 as=2.88054e+06 ps=7896 
M5137 idl2 idl2 Vdd GND dfet w=846 l=1504
+ ad=2.65964e+06 pd=7708 as=0 ps=0 
M5138 n_1376 cp1 notdor2 GND efet w=1034 l=752
+ ad=7.97891e+06 pd=25004 as=1.97043e+06 ps=7708 
M5139 idl2 cp1 n_1424 GND efet w=5687 l=705
+ ad=1.20876e+07 pd=31772 as=0 ps=0 
M5140 n_1424 dpc42_DL_ADH adh2 GND efet w=4136 l=752
+ ad=0 pd=0 as=0 ps=0 
M5141 GND idb2 n_1376 GND efet w=4371 l=611
+ ad=0 pd=0 as=0 ps=0 
M5142 dor2 notdor2 GND GND efet w=6580 l=564
+ ad=7.55478e+06 pd=23876 as=0 ps=0 
M5143 GND notidl2 idl2 GND efet w=3572 l=564
+ ad=0 pd=0 as=0 ps=0 
M5144 Vdd n_1199 n_1199 GND dfet w=846 l=658
+ ad=0 pd=0 as=2.21784e+06 ps=9024 
M5145 db1 n_794 GND GND efet w=21009 l=517
+ ad=0 pd=0 as=0 ps=0 
M5146 db1 n_798 Vdd GND efet w=60113 l=611
+ ad=0 pd=0 as=0 ps=0 
M5147 GND n_794 db1 GND efet w=1034 l=564
+ ad=0 pd=0 as=0 ps=0 
M5148 n_1661 dpc41_DL_ADL adl3 GND efet w=5640 l=658
+ ad=1.74246e+07 pd=47000 as=0 ps=0 
M5149 adh4 cclk Vdd GND efet w=2068 l=564
+ ad=0 pd=0 as=0 ps=0 
M5150 adl5 cclk Vdd GND efet w=2162 l=564
+ ad=0 pd=0 as=0 ps=0 
M5151 adh5 cclk Vdd GND efet w=2350 l=658
+ ad=0 pd=0 as=0 ps=0 
M5152 idb2 dpc43_DL_DB n_1424 GND efet w=4136 l=658
+ ad=0 pd=0 as=0 ps=0 
M5153 GND notidl2 idl2 GND efet w=3149 l=517
+ ad=0 pd=0 as=0 ps=0 
M5154 n_1199 cclk notidl2 GND efet w=1316 l=658
+ ad=1.52863e+07 pd=36096 as=1.93508e+06 ps=6768 
M5155 GND db2 n_1199 GND efet w=12455 l=611
+ ad=0 pd=0 as=0 ps=0 
M5156 idl2 notidl2 GND GND efet w=4606 l=658
+ ad=0 pd=0 as=0 ps=0 
M5157 n_520 RnWstretched GND GND efet w=14382 l=564
+ ad=1.96513e+07 pd=51700 as=0 ps=0 
M5158 n_520 RnWstretched GND GND efet w=14523 l=517
+ ad=0 pd=0 as=0 ps=0 
M5159 GND n_224 n_520 GND efet w=13207 l=611
+ ad=0 pd=0 as=0 ps=0 
M5160 GND RnWstretched n_224 GND efet w=7003 l=611
+ ad=0 pd=0 as=6.68002e+06 ps=19928 
M5161 Vdd cclk idb2 GND efet w=2068 l=752
+ ad=0 pd=0 as=0 ps=0 
M5162 n_520 dor2 Vdd GND dfet w=1504 l=658
+ ad=0 pd=0 as=0 ps=0 
M5163 Vdd n_224 n_224 GND dfet w=846 l=752
+ ad=0 pd=0 as=1.43408e+07 ps=46248 
M5164 n_37 n_224 Vdd GND dfet w=1598 l=658
+ ad=2.22137e+07 pd=52452 as=0 ps=0 
M5165 GND RnWstretched n_37 GND efet w=8930 l=564
+ ad=0 pd=0 as=0 ps=0 
M5166 GND RnWstretched n_37 GND efet w=18894 l=564
+ ad=0 pd=0 as=0 ps=0 
M5167 n_37 dor2 GND GND efet w=13959 l=611
+ ad=0 pd=0 as=0 ps=0 
M5168 n_224 dor2 GND GND efet w=5640 l=658
+ ad=0 pd=0 as=0 ps=0 
M5169 GND n_794 db1 GND efet w=23030 l=564
+ ad=0 pd=0 as=0 ps=0 
M5170 GND GND db1 GND efet w=5358 l=752
+ ad=0 pd=0 as=0 ps=0 
M5171 GND GND db2 GND efet w=5170 l=564
+ ad=0 pd=0 as=2.19177e+08 ps=400440 
M5172 db2 n_520 Vdd GND efet w=60066 l=658
+ ad=0 pd=0 as=0 ps=0 
M5173 dor2 dor2 Vdd GND dfet w=940 l=1128
+ ad=2.0473e+07 pd=63544 as=0 ps=0 
M5174 Vdd n_457 n_457 GND dfet w=846 l=1598
+ ad=0 pd=0 as=2.98657e+06 ps=8084 
M5175 idl3 idl3 Vdd GND dfet w=846 l=1598
+ ad=2.80101e+06 pd=7896 as=0 ps=0 
M5176 n_457 cp1 notdor3 GND efet w=1128 l=752
+ ad=8.43838e+06 pd=25756 as=1.79371e+06 ps=7520 
M5177 idl3 cp1 n_1661 GND efet w=5687 l=705
+ ad=1.16193e+07 pd=31020 as=0 ps=0 
M5178 n_1661 dpc42_DL_ADH adh3 GND efet w=4136 l=752
+ ad=0 pd=0 as=0 ps=0 
M5179 GND idb3 n_457 GND efet w=4324 l=564
+ ad=0 pd=0 as=0 ps=0 
M5180 dor3 notdor3 GND GND efet w=6439 l=611
+ ad=7.72266e+06 pd=23312 as=0 ps=0 
M5181 GND notidl3 idl3 GND efet w=3478 l=658
+ ad=0 pd=0 as=0 ps=0 
M5182 db2 n_37 db2 GND efet w=752 l=564
+ ad=0 pd=0 as=0 ps=0 
M5183 Vdd n_896 n_896 GND dfet w=940 l=658
+ ad=0 pd=0 as=2.26202e+06 ps=9212 
M5184 n_896 cclk notidl3 GND efet w=1316 l=752
+ ad=1.54983e+07 pd=36096 as=1.99694e+06 ps=6956 
M5185 db2 n_37 GND GND efet w=21197 l=611
+ ad=0 pd=0 as=0 ps=0 
M5186 GND n_37 db2 GND efet w=752 l=564
+ ad=0 pd=0 as=0 ps=0 
M5187 GND db3 n_896 GND efet w=12596 l=658
+ ad=0 pd=0 as=0 ps=0 
M5188 n_1095 dpc41_DL_ADL adl4 GND efet w=5781 l=705
+ ad=1.78929e+07 pd=47376 as=0 ps=0 
M5189 idb3 dpc43_DL_DB n_1661 GND efet w=4042 l=564
+ ad=0 pd=0 as=0 ps=0 
M5190 GND notidl3 idl3 GND efet w=3196 l=564
+ ad=0 pd=0 as=0 ps=0 
M5191 n_42 RnWstretched GND GND efet w=14288 l=564
+ ad=1.95894e+07 pd=51700 as=0 ps=0 
M5192 n_42 RnWstretched GND GND efet w=14429 l=517
+ ad=0 pd=0 as=0 ps=0 
M5193 idl3 notidl3 GND GND efet w=4559 l=611
+ ad=0 pd=0 as=0 ps=0 
M5194 GND n_1613 n_42 GND efet w=13254 l=564
+ ad=0 pd=0 as=0 ps=0 
M5195 GND RnWstretched n_1613 GND efet w=7003 l=705
+ ad=0 pd=0 as=6.627e+06 ps=19740 
M5196 Vdd cclk idb3 GND efet w=2162 l=752
+ ad=0 pd=0 as=0 ps=0 
M5197 n_42 dor3 Vdd GND dfet w=1504 l=658
+ ad=0 pd=0 as=0 ps=0 
M5198 db2 n_37 GND GND efet w=21150 l=564
+ ad=0 pd=0 as=0 ps=0 
M5199 db2 n_520 Vdd GND efet w=60019 l=611
+ ad=0 pd=0 as=0 ps=0 
M5200 GND n_37 db2 GND efet w=1034 l=564
+ ad=0 pd=0 as=0 ps=0 
M5201 Vdd n_1613 n_1613 GND dfet w=940 l=752
+ ad=0 pd=0 as=1.36251e+07 ps=46060 
M5202 n_643 n_1613 Vdd GND dfet w=1598 l=564
+ ad=2.24788e+07 pd=52264 as=0 ps=0 
M5203 GND RnWstretched n_643 GND efet w=8883 l=611
+ ad=0 pd=0 as=0 ps=0 
M5204 GND RnWstretched n_643 GND efet w=18847 l=611
+ ad=0 pd=0 as=0 ps=0 
M5205 n_643 dor3 GND GND efet w=13959 l=611
+ ad=0 pd=0 as=0 ps=0 
M5206 n_1613 dor3 GND GND efet w=5546 l=658
+ ad=0 pd=0 as=0 ps=0 
M5207 dor3 dor3 Vdd GND dfet w=940 l=1128
+ ad=2.04642e+07 pd=63356 as=0 ps=0 
M5208 Vdd n_797 n_797 GND dfet w=846 l=1598
+ ad=0 pd=0 as=3.07493e+06 ps=8084 
M5209 idl4 idl4 Vdd GND dfet w=940 l=1598
+ ad=3.03075e+06 pd=8084 as=0 ps=0 
M5210 n_797 cp1 notdor4 GND efet w=1034 l=752
+ ad=7.45758e+06 pd=25192 as=1.71418e+06 ps=7332 
M5211 idl4 cp1 n_1095 GND efet w=5875 l=705
+ ad=1.14073e+07 pd=31396 as=0 ps=0 
M5212 n_1095 dpc42_DL_ADH adh4 GND efet w=4042 l=752
+ ad=0 pd=0 as=0 ps=0 
M5213 GND idb4 n_797 GND efet w=4324 l=564
+ ad=0 pd=0 as=0 ps=0 
M5214 dor4 notdor4 GND GND efet w=6486 l=564
+ ad=7.75801e+06 pd=23500 as=0 ps=0 
M5215 GND notidl4 idl4 GND efet w=3572 l=658
+ ad=0 pd=0 as=0 ps=0 
M5216 db2 n_37 GND GND efet w=22748 l=564
+ ad=0 pd=0 as=0 ps=0 
M5217 GND n_37 db2 GND efet w=1034 l=564
+ ad=0 pd=0 as=0 ps=0 
M5218 db2 n_37 GND GND efet w=17155 l=611
+ ad=0 pd=0 as=0 ps=0 
M5219 db2 n_37 GND GND efet w=14664 l=564
+ ad=0 pd=0 as=0 ps=0 
M5220 GND n_643 db3 GND efet w=14664 l=658
+ ad=0 pd=0 as=2.27297e+08 ps=408900 
M5221 GND n_643 db3 GND efet w=22184 l=658
+ ad=0 pd=0 as=0 ps=0 
M5222 Vdd n_490 n_490 GND dfet w=940 l=752
+ ad=0 pd=0 as=2.46524e+06 ps=9400 
M5223 db3 n_42 Vdd GND efet w=59831 l=611
+ ad=0 pd=0 as=0 ps=0 
M5224 db3 n_643 GND GND efet w=19928 l=564
+ ad=0 pd=0 as=0 ps=0 
M5225 n_490 cclk notidl4 GND efet w=1222 l=752
+ ad=1.5463e+07 pd=35532 as=1.8909e+06 ps=7144 
M5226 GND db4 n_490 GND efet w=12455 l=611
+ ad=0 pd=0 as=0 ps=0 
M5227 n_1387 dpc41_DL_ADL adl5 GND efet w=5781 l=611
+ ad=1.79017e+07 pd=47564 as=0 ps=0 
M5228 adl6 cclk Vdd GND efet w=2162 l=658
+ ad=0 pd=0 as=0 ps=0 
M5229 Vdd cclk adh6 GND efet w=2350 l=658
+ ad=0 pd=0 as=0 ps=0 
M5230 Vdd cclk adl7 GND efet w=2162 l=658
+ ad=0 pd=0 as=0 ps=0 
M5231 dpc31_PCHPCH cclk GND GND efet w=2444 l=658
+ ad=0 pd=0 as=0 ps=0 
M5232 aluvout aluvout Vdd GND dfet w=940 l=658
+ ad=9.17972e+07 pd=332196 as=0 ps=0 
M5233 n_1267 n_1267 Vdd GND dfet w=846 l=940
+ ad=2.04995e+06 pd=6956 as=0 ps=0 
M5234 n_676 abh1 GND GND efet w=13818 l=658
+ ad=9.64891e+06 pd=33088 as=0 ps=0 
M5235 Vdd n_617 n_676 GND dfet w=1786 l=658
+ ad=0 pd=0 as=0 ps=0 
M5236 nABH1 cclk n_676 GND efet w=1128 l=752
+ ad=3.60509e+06 pd=11092 as=0 ps=0 
M5237 n_1298 ADH_ABH nABH1 GND efet w=1128 l=752
+ ad=636192 pd=3384 as=0 ps=0 
M5238 n_1267 cp1 n_1298 GND efet w=1128 l=658
+ ad=8.14679e+06 pd=22748 as=0 ps=0 
M5239 GND adh1 n_1267 GND efet w=7050 l=658
+ ad=0 pd=0 as=0 ps=0 
M5240 n_168 adh2 GND GND efet w=7050 l=658
+ ad=7.69616e+06 pd=22936 as=0 ps=0 
M5241 Vdd n_168 n_168 GND dfet w=940 l=846
+ ad=0 pd=0 as=1.79371e+06 ps=6768 
M5242 abh2 nABH2 GND GND efet w=6204 l=658
+ ad=4.61239e+06 pd=17860 as=0 ps=0 
M5243 Vdd abh2 abh2 GND dfet w=846 l=1410
+ ad=0 pd=0 as=1.91388e+07 ps=62228 
M5244 GND n_1034 n_1545 GND efet w=10622 l=470
+ ad=0 pd=0 as=1.70888e+07 ps=37976 
M5245 GND n_1346 n_1296 GND efet w=10622 l=470
+ ad=0 pd=0 as=1.69828e+07 ps=37976 
M5246 n_1545 abh2 Vdd GND dfet w=1598 l=564
+ ad=0 pd=0 as=0 ps=0 
M5247 Vdd n_1034 n_1034 GND dfet w=846 l=940
+ ad=0 pd=0 as=1.74423e+07 ps=63920 
M5248 GND abh2 n_1034 GND efet w=4136 l=658
+ ad=0 pd=0 as=4.16176e+06 ps=13724 
M5249 n_836 cp1 n_168 GND efet w=1128 l=752
+ ad=530160 pd=3196 as=0 ps=0 
M5250 nABH2 ADH_ABH n_836 GND efet w=1128 l=752
+ ad=3.50789e+06 pd=10716 as=0 ps=0 
M5251 nABH2 cclk n_994 GND efet w=1128 l=752
+ ad=0 pd=0 as=1.04265e+07 ps=33464 
M5252 Vdd n_1034 n_994 GND dfet w=1692 l=752
+ ad=0 pd=0 as=0 ps=0 
M5253 GND abh2 n_994 GND efet w=13912 l=658
+ ad=0 pd=0 as=0 ps=0 
M5254 GND n_676 ab9 GND efet w=3854 l=470
+ ad=0 pd=0 as=0 ps=0 
M5255 GND n_676 ab9 GND efet w=1128 l=470
+ ad=0 pd=0 as=0 ps=0 
M5256 GND n_994 ab10 GND efet w=1222 l=564
+ ad=0 pd=0 as=1.66099e+08 ps=217328 
M5257 GND n_994 ab10 GND efet w=3854 l=564
+ ad=0 pd=0 as=0 ps=0 
M5258 GND n_676 ab9 GND efet w=15322 l=658
+ ad=0 pd=0 as=0 ps=0 
M5259 ab9 n_676 GND GND efet w=15322 l=658
+ ad=0 pd=0 as=0 ps=0 
M5260 GND n_676 ab9 GND efet w=15322 l=564
+ ad=0 pd=0 as=0 ps=0 
M5261 ab9 n_676 GND GND efet w=15322 l=658
+ ad=0 pd=0 as=0 ps=0 
M5262 GND n_676 ab9 GND efet w=15322 l=658
+ ad=0 pd=0 as=0 ps=0 
M5263 ab10 n_994 GND GND efet w=15322 l=564
+ ad=0 pd=0 as=0 ps=0 
M5264 GND n_994 ab10 GND efet w=15322 l=564
+ ad=0 pd=0 as=0 ps=0 
M5265 ab10 n_994 GND GND efet w=15322 l=564
+ ad=0 pd=0 as=0 ps=0 
M5266 GND n_994 ab10 GND efet w=15322 l=658
+ ad=0 pd=0 as=0 ps=0 
M5267 ab10 n_994 GND GND efet w=15322 l=658
+ ad=0 pd=0 as=0 ps=0 
M5268 Vdd n_1545 ab10 GND efet w=39151 l=611
+ ad=0 pd=0 as=0 ps=0 
M5269 Vdd n_1545 ab10 GND efet w=29704 l=564
+ ad=0 pd=0 as=0 ps=0 
M5270 Vdd n_1545 ab10 GND efet w=14946 l=658
+ ad=0 pd=0 as=0 ps=0 
M5271 ab11 n_1296 Vdd GND efet w=14946 l=658
+ ad=1.63537e+08 pd=217328 as=0 ps=0 
M5272 Vdd n_1296 ab11 GND efet w=29892 l=564
+ ad=0 pd=0 as=0 ps=0 
M5273 Vdd n_1296 ab11 GND efet w=39292 l=658
+ ad=0 pd=0 as=0 ps=0 
M5274 Vdd abh3 n_1296 GND dfet w=1598 l=658
+ ad=0 pd=0 as=0 ps=0 
M5275 n_1346 abh3 GND GND efet w=4324 l=658
+ ad=4.09107e+06 pd=12596 as=0 ps=0 
M5276 Vdd n_1346 n_1346 GND dfet w=846 l=940
+ ad=0 pd=0 as=1.65498e+07 ps=63920 
M5277 abh3 abh3 Vdd GND dfet w=752 l=1222
+ ad=2.0367e+07 pd=62040 as=0 ps=0 
M5278 GND nABH3 abh3 GND efet w=6110 l=564
+ ad=0 pd=0 as=5.49599e+06 ps=17672 
M5279 n_883 n_883 Vdd GND dfet w=846 l=846
+ ad=1.88207e+06 pd=6768 as=0 ps=0 
M5280 n_359 abh3 GND GND efet w=14006 l=658
+ ad=9.23362e+06 pd=32524 as=0 ps=0 
M5281 Vdd n_1346 n_359 GND dfet w=1786 l=564
+ ad=0 pd=0 as=0 ps=0 
M5282 nABH3 cclk n_359 GND efet w=1034 l=658
+ ad=3.46371e+06 pd=11092 as=0 ps=0 
M5283 n_1667 ADH_ABH nABH3 GND efet w=1034 l=752
+ ad=485980 pd=3008 as=0 ps=0 
M5284 n_883 cp1 n_1667 GND efet w=1034 l=658
+ ad=8.45605e+06 pd=22560 as=0 ps=0 
M5285 GND adh3 n_883 GND efet w=7050 l=564
+ ad=0 pd=0 as=0 ps=0 
M5286 n_212 adh4 GND GND efet w=7050 l=564
+ ad=7.08647e+06 pd=22936 as=0 ps=0 
M5287 Vdd n_212 n_212 GND dfet w=846 l=940
+ ad=0 pd=0 as=2.13831e+06 ps=7144 
M5288 abh4 nABH4 GND GND efet w=6110 l=658
+ ad=4.44451e+06 pd=17296 as=0 ps=0 
M5289 Vdd abh4 abh4 GND dfet w=846 l=1316
+ ad=0 pd=0 as=1.9934e+07 ps=62040 
M5290 GND n_1677 n_475 GND efet w=10528 l=658
+ ad=0 pd=0 as=1.48533e+07 ps=36284 
M5291 GND n_1423 n_1608 GND efet w=10622 l=658
+ ad=0 pd=0 as=1.52244e+07 ps=36472 
M5292 n_475 abh4 Vdd GND dfet w=1598 l=658
+ ad=0 pd=0 as=0 ps=0 
M5293 Vdd n_1677 n_1677 GND dfet w=940 l=846
+ ad=0 pd=0 as=1.91034e+07 ps=63544 
M5294 GND abh4 n_1677 GND efet w=4277 l=611
+ ad=0 pd=0 as=4.87747e+06 ps=14476 
M5295 n_1451 cp1 n_212 GND efet w=1128 l=752
+ ad=424128 pd=3008 as=0 ps=0 
M5296 nABH4 ADH_ABH n_1451 GND efet w=1128 l=752
+ ad=3.40186e+06 pd=10528 as=0 ps=0 
M5297 nABH4 cclk n_999 GND efet w=1034 l=752
+ ad=0 pd=0 as=1.07446e+07 ps=33464 
M5298 Vdd n_1677 n_999 GND dfet w=1880 l=658
+ ad=0 pd=0 as=0 ps=0 
M5299 GND abh4 n_999 GND efet w=13865 l=611
+ ad=0 pd=0 as=0 ps=0 
M5300 GND n_359 ab11 GND efet w=3854 l=564
+ ad=0 pd=0 as=0 ps=0 
M5301 GND n_359 ab11 GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M5302 GND n_359 ab11 GND efet w=15322 l=564
+ ad=0 pd=0 as=0 ps=0 
M5303 ab11 n_359 GND GND efet w=15322 l=564
+ ad=0 pd=0 as=0 ps=0 
M5304 GND n_359 ab11 GND efet w=15322 l=564
+ ad=0 pd=0 as=0 ps=0 
M5305 ab11 n_359 GND GND efet w=15322 l=752
+ ad=0 pd=0 as=0 ps=0 
M5306 GND n_359 ab11 GND efet w=15322 l=658
+ ad=0 pd=0 as=0 ps=0 
M5307 GND n_999 ab12 GND efet w=1222 l=470
+ ad=0 pd=0 as=1.65825e+08 ps=218080 
M5308 GND n_999 ab12 GND efet w=3854 l=470
+ ad=0 pd=0 as=0 ps=0 
M5309 ab12 n_999 GND GND efet w=15416 l=658
+ ad=0 pd=0 as=0 ps=0 
M5310 GND n_999 ab12 GND efet w=15416 l=564
+ ad=0 pd=0 as=0 ps=0 
M5311 ab12 n_999 GND GND efet w=15416 l=564
+ ad=0 pd=0 as=0 ps=0 
M5312 GND n_999 ab12 GND efet w=15322 l=564
+ ad=0 pd=0 as=0 ps=0 
M5313 ab12 n_999 GND GND efet w=15322 l=564
+ ad=0 pd=0 as=0 ps=0 
M5314 Vdd n_475 ab12 GND efet w=39104 l=658
+ ad=0 pd=0 as=0 ps=0 
M5315 Vdd n_475 ab12 GND efet w=29610 l=564
+ ad=0 pd=0 as=0 ps=0 
M5316 Vdd n_475 ab12 GND efet w=15040 l=658
+ ad=0 pd=0 as=0 ps=0 
M5317 ab13 n_1608 Vdd GND efet w=15040 l=658
+ ad=1.61284e+08 pd=217140 as=0 ps=0 
M5318 Vdd n_1608 ab13 GND efet w=29704 l=564
+ ad=0 pd=0 as=0 ps=0 
M5319 Vdd n_1608 ab13 GND efet w=39104 l=658
+ ad=0 pd=0 as=0 ps=0 
M5320 Vdd abh5 n_1608 GND dfet w=1598 l=658
+ ad=0 pd=0 as=0 ps=0 
M5321 n_1423 abh5 GND GND efet w=4136 l=658
+ ad=3.91435e+06 pd=12596 as=0 ps=0 
M5322 Vdd n_1423 n_1423 GND dfet w=846 l=1034
+ ad=0 pd=0 as=1.95717e+07 ps=64108 
M5323 abh5 abh5 Vdd GND dfet w=940 l=1222
+ ad=1.89974e+07 pd=62040 as=0 ps=0 
M5324 GND nABH5 abh5 GND efet w=6204 l=658
+ ad=0 pd=0 as=5.82292e+06 ps=18048 
M5325 Vdd cclk adh7 GND efet w=2162 l=658
+ ad=0 pd=0 as=0 ps=0 
M5326 dpc39_PCLPCL cclk GND GND efet w=2538 l=846
+ ad=0 pd=0 as=0 ps=0 
M5327 dpc40_ADLPCL cclk GND GND efet w=2444 l=846
+ ad=0 pd=0 as=0 ps=0 
M5328 idb4 dpc43_DL_DB n_1095 GND efet w=4136 l=658
+ ad=0 pd=0 as=0 ps=0 
M5329 GND notidl4 idl4 GND efet w=3149 l=611
+ ad=0 pd=0 as=0 ps=0 
M5330 n_1076 RnWstretched GND GND efet w=14335 l=611
+ ad=2.05084e+07 pd=51700 as=0 ps=0 
M5331 GND RnWstretched n_1076 GND efet w=14664 l=564
+ ad=0 pd=0 as=0 ps=0 
M5332 idl4 notidl4 GND GND efet w=4512 l=658
+ ad=0 pd=0 as=0 ps=0 
M5333 GND RnWstretched n_1463 GND efet w=6909 l=611
+ ad=0 pd=0 as=6.75954e+06 ps=19552 
M5334 GND n_1463 n_1076 GND efet w=12925 l=611
+ ad=0 pd=0 as=0 ps=0 
M5335 Vdd cclk idb4 GND efet w=2068 l=752
+ ad=0 pd=0 as=0 ps=0 
M5336 n_1076 dor4 Vdd GND dfet w=1504 l=658
+ ad=0 pd=0 as=0 ps=0 
M5337 GND n_643 db3 GND efet w=1128 l=564
+ ad=0 pd=0 as=0 ps=0 
M5338 Vdd n_1463 n_1463 GND dfet w=846 l=752
+ ad=0 pd=0 as=1.37311e+07 ps=46248 
M5339 n_147 n_1463 Vdd GND dfet w=1598 l=658
+ ad=2.18338e+07 pd=51512 as=0 ps=0 
M5340 GND RnWstretched n_147 GND efet w=8977 l=611
+ ad=0 pd=0 as=0 ps=0 
M5341 GND RnWstretched n_147 GND efet w=18941 l=611
+ ad=0 pd=0 as=0 ps=0 
M5342 n_147 dor4 GND GND efet w=13865 l=611
+ ad=0 pd=0 as=0 ps=0 
M5343 n_1463 dor4 GND GND efet w=5452 l=564
+ ad=0 pd=0 as=0 ps=0 
M5344 dor4 dor4 Vdd GND dfet w=846 l=1034
+ ad=1.90504e+07 pd=63356 as=0 ps=0 
M5345 Vdd n_961 n_961 GND dfet w=940 l=1598
+ ad=0 pd=0 as=2.93355e+06 ps=7896 
M5346 idl5 idl5 Vdd GND dfet w=846 l=1598
+ ad=2.80101e+06 pd=7896 as=0 ps=0 
M5347 n_961 cp1 notdor5 GND efet w=1034 l=752
+ ad=7.62547e+06 pd=25380 as=1.89974e+06 ps=7332 
M5348 idl5 cp1 n_1387 GND efet w=5922 l=658
+ ad=1.20965e+07 pd=31584 as=0 ps=0 
M5349 n_1387 dpc42_DL_ADH adh5 GND efet w=4042 l=752
+ ad=0 pd=0 as=0 ps=0 
M5350 GND idb5 n_961 GND efet w=4324 l=564
+ ad=0 pd=0 as=0 ps=0 
M5351 dor5 notdor5 GND GND efet w=6533 l=611
+ ad=8.12912e+06 pd=23876 as=0 ps=0 
M5352 GND notidl5 idl5 GND efet w=3572 l=658
+ ad=0 pd=0 as=0 ps=0 
M5353 Vdd n_568 n_568 GND dfet w=940 l=658
+ ad=0 pd=0 as=2.31503e+06 ps=9212 
M5354 n_568 cclk notidl5 GND efet w=1316 l=752
+ ad=1.63024e+07 pd=35908 as=1.91741e+06 ps=7144 
M5355 GND db5 n_568 GND efet w=12502 l=564
+ ad=0 pd=0 as=0 ps=0 
M5356 n_1014 dpc41_DL_ADL adl6 GND efet w=6016 l=658
+ ad=1.76897e+07 pd=47564 as=0 ps=0 
M5357 idb5 dpc43_DL_DB n_1387 GND efet w=4042 l=658
+ ad=0 pd=0 as=0 ps=0 
M5358 GND notidl5 idl5 GND efet w=3149 l=611
+ ad=0 pd=0 as=0 ps=0 
M5359 db3 n_643 GND GND efet w=19928 l=564
+ ad=0 pd=0 as=0 ps=0 
M5360 GND n_643 db3 GND efet w=1034 l=564
+ ad=0 pd=0 as=0 ps=0 
M5361 db3 n_42 Vdd GND efet w=60207 l=611
+ ad=0 pd=0 as=0 ps=0 
M5362 GND n_643 db3 GND efet w=21996 l=564
+ ad=0 pd=0 as=0 ps=0 
M5363 GND GND db3 GND efet w=5123 l=705
+ ad=0 pd=0 as=0 ps=0 
M5364 GND GND db4 GND efet w=5170 l=658
+ ad=0 pd=0 as=2.43644e+08 ps=442552 
M5365 n_373 RnWstretched GND GND efet w=14335 l=611
+ ad=2.0314e+07 pd=51512 as=0 ps=0 
M5366 n_373 RnWstretched GND GND efet w=14570 l=564
+ ad=0 pd=0 as=0 ps=0 
M5367 idl5 notidl5 GND GND efet w=4559 l=705
+ ad=0 pd=0 as=0 ps=0 
M5368 GND n_1720 n_373 GND efet w=13066 l=564
+ ad=0 pd=0 as=0 ps=0 
M5369 GND RnWstretched n_1720 GND efet w=6956 l=658
+ ad=0 pd=0 as=6.59166e+06 ps=19928 
M5370 Vdd cclk idb5 GND efet w=1974 l=752
+ ad=0 pd=0 as=0 ps=0 
M5371 n_373 dor5 Vdd GND dfet w=1598 l=658
+ ad=0 pd=0 as=0 ps=0 
M5372 db4 n_1076 Vdd GND efet w=60066 l=658
+ ad=0 pd=0 as=0 ps=0 
M5373 db4 n_147 db4 GND efet w=846 l=470
+ ad=0 pd=0 as=0 ps=0 
M5374 Vdd n_1720 n_1720 GND dfet w=940 l=752
+ ad=0 pd=0 as=1.32982e+07 ps=46060 
M5375 n_612 n_1720 Vdd GND dfet w=1598 l=564
+ ad=2.07204e+07 pd=51888 as=0 ps=0 
M5376 GND RnWstretched n_612 GND efet w=8930 l=658
+ ad=0 pd=0 as=0 ps=0 
M5377 GND RnWstretched n_612 GND efet w=18894 l=658
+ ad=0 pd=0 as=0 ps=0 
M5378 n_612 dor5 GND GND efet w=13865 l=611
+ ad=0 pd=0 as=0 ps=0 
M5379 n_1720 dor5 GND GND efet w=5546 l=658
+ ad=0 pd=0 as=0 ps=0 
M5380 db4 n_147 GND GND efet w=20304 l=564
+ ad=0 pd=0 as=0 ps=0 
M5381 GND n_147 db4 GND efet w=846 l=470
+ ad=0 pd=0 as=0 ps=0 
M5382 dor5 dor5 Vdd GND dfet w=893 l=1175
+ ad=2.04642e+07 pd=63356 as=0 ps=0 
M5383 Vdd n_1684 n_1684 GND dfet w=846 l=1598
+ ad=0 pd=0 as=3.03075e+06 ps=8084 
M5384 idl6 idl6 Vdd GND dfet w=846 l=1504
+ ad=2.80101e+06 pd=7896 as=0 ps=0 
M5385 n_1684 cp1 notdor6 GND efet w=1128 l=752
+ ad=7.52827e+06 pd=25568 as=1.67884e+06 ps=7332 
M5386 idl6 cp1 n_1014 GND efet w=6110 l=658
+ ad=1.23527e+07 pd=32148 as=0 ps=0 
M5387 n_1014 dpc42_DL_ADH adh6 GND efet w=4042 l=752
+ ad=0 pd=0 as=0 ps=0 
M5388 GND idb6 n_1684 GND efet w=4371 l=611
+ ad=0 pd=0 as=0 ps=0 
M5389 dor6 notdor6 GND GND efet w=6580 l=564
+ ad=7.8552e+06 pd=23688 as=0 ps=0 
M5390 GND notidl6 idl6 GND efet w=3478 l=564
+ ad=0 pd=0 as=0 ps=0 
M5391 Vdd n_1638 n_1638 GND dfet w=752 l=658
+ ad=0 pd=0 as=2.26202e+06 ps=9212 
M5392 n_1638 cclk notidl6 GND efet w=1316 l=752
+ ad=1.63113e+07 pd=35908 as=1.93508e+06 ps=6956 
M5393 GND db6 n_1638 GND efet w=12502 l=564
+ ad=0 pd=0 as=0 ps=0 
M5394 n_1147 dpc41_DL_ADL adl7 GND efet w=5828 l=658
+ ad=1.81845e+07 pd=47940 as=0 ps=0 
M5395 idb6 dpc43_DL_DB n_1014 GND efet w=4042 l=658
+ ad=0 pd=0 as=0 ps=0 
M5396 GND notidl6 idl6 GND efet w=3196 l=564
+ ad=0 pd=0 as=0 ps=0 
M5397 n_7 RnWstretched GND GND efet w=14335 l=611
+ ad=2.01814e+07 pd=51512 as=0 ps=0 
M5398 n_7 RnWstretched GND GND efet w=14476 l=564
+ ad=0 pd=0 as=0 ps=0 
M5399 idl6 notidl6 GND GND efet w=4747 l=611
+ ad=0 pd=0 as=0 ps=0 
M5400 GND n_466 n_7 GND efet w=13019 l=611
+ ad=0 pd=0 as=0 ps=0 
M5401 GND RnWstretched n_466 GND efet w=7050 l=658
+ ad=0 pd=0 as=7.10414e+06 ps=20116 
M5402 Vdd cclk idb6 GND efet w=2068 l=658
+ ad=0 pd=0 as=0 ps=0 
M5403 n_7 dor6 Vdd GND dfet w=1598 l=658
+ ad=0 pd=0 as=0 ps=0 
M5404 Vdd n_466 n_466 GND dfet w=752 l=752
+ ad=0 pd=0 as=1.36958e+07 ps=46248 
M5405 n_471 n_466 Vdd GND dfet w=1598 l=658
+ ad=2.32917e+07 pd=51888 as=0 ps=0 
M5406 GND RnWstretched n_471 GND efet w=8977 l=611
+ ad=0 pd=0 as=0 ps=0 
M5407 db4 n_147 GND GND efet w=20116 l=564
+ ad=0 pd=0 as=0 ps=0 
M5408 db4 n_1076 Vdd GND efet w=59596 l=658
+ ad=0 pd=0 as=0 ps=0 
M5409 GND n_147 db4 GND efet w=1034 l=470
+ ad=0 pd=0 as=0 ps=0 
M5410 db4 n_147 GND GND efet w=20210 l=564
+ ad=0 pd=0 as=0 ps=0 
M5411 GND n_147 db4 GND efet w=1034 l=470
+ ad=0 pd=0 as=0 ps=0 
M5412 db4 n_147 GND GND efet w=14664 l=658
+ ad=0 pd=0 as=0 ps=0 
M5413 db4 n_147 GND GND efet w=21479 l=611
+ ad=0 pd=0 as=0 ps=0 
M5414 GND n_612 db5 GND efet w=14570 l=658
+ ad=0 pd=0 as=2.62491e+08 ps=475640 
M5415 GND n_612 db5 GND efet w=21432 l=658
+ ad=0 pd=0 as=0 ps=0 
M5416 GND RnWstretched n_471 GND efet w=18894 l=564
+ ad=0 pd=0 as=0 ps=0 
M5417 n_471 dor6 GND GND efet w=13959 l=611
+ ad=0 pd=0 as=0 ps=0 
M5418 n_466 dor6 GND GND efet w=5640 l=564
+ ad=0 pd=0 as=0 ps=0 
M5419 db5 n_373 Vdd GND efet w=59925 l=611
+ ad=0 pd=0 as=0 ps=0 
M5420 dor6 dor6 Vdd GND dfet w=940 l=1128
+ ad=1.90062e+07 pd=63732 as=0 ps=0 
M5421 db5 n_612 GND GND efet w=20022 l=564
+ ad=0 pd=0 as=0 ps=0 
M5422 Vdd n_789 n_789 GND dfet w=846 l=1598
+ ad=0 pd=0 as=3.03075e+06 ps=8084 
M5423 idl7 idl7 Vdd GND dfet w=846 l=1598
+ ad=2.95122e+06 pd=8084 as=0 ps=0 
M5424 n_789 cp1 notdor7 GND efet w=1128 l=752
+ ad=8.42071e+06 pd=25192 as=2.01461e+06 ps=8084 
M5425 idl7 cp1 n_1147 GND efet w=6110 l=658
+ ad=1.19374e+07 pd=31960 as=0 ps=0 
M5426 n_1147 dpc42_DL_ADH adh7 GND efet w=4042 l=658
+ ad=0 pd=0 as=0 ps=0 
M5427 GND idb7 n_789 GND efet w=4183 l=611
+ ad=0 pd=0 as=0 ps=0 
M5428 dor7 notdor7 GND GND efet w=6486 l=564
+ ad=7.81102e+06 pd=23500 as=0 ps=0 
M5429 GND notidl7 idl7 GND efet w=3384 l=564
+ ad=0 pd=0 as=0 ps=0 
M5430 GND n_612 db5 GND efet w=1222 l=658
+ ad=0 pd=0 as=0 ps=0 
M5431 Vdd n_588 n_588 GND dfet w=940 l=658
+ ad=0 pd=0 as=2.26202e+06 ps=9212 
M5432 idb7 dpc43_DL_DB n_1147 GND efet w=4136 l=658
+ ad=0 pd=0 as=0 ps=0 
M5433 GND notidl7 idl7 GND efet w=3290 l=564
+ ad=0 pd=0 as=0 ps=0 
M5434 n_588 cclk notidl7 GND efet w=1316 l=752
+ ad=1.55514e+07 pd=35908 as=1.8644e+06 ps=6768 
M5435 GND db7 n_588 GND efet w=12596 l=658
+ ad=0 pd=0 as=0 ps=0 
M5436 GND notidl7 idl7 GND efet w=4512 l=658
+ ad=0 pd=0 as=0 ps=0 
M5437 n_298 RnWstretched GND GND efet w=14288 l=564
+ ad=1.98368e+07 pd=51888 as=0 ps=0 
M5438 n_298 RnWstretched GND GND efet w=14758 l=564
+ ad=0 pd=0 as=0 ps=0 
M5439 GND n_23 n_298 GND efet w=13019 l=611
+ ad=0 pd=0 as=0 ps=0 
M5440 GND RnWstretched n_23 GND efet w=7003 l=611
+ ad=0 pd=0 as=6.96277e+06 ps=20116 
M5441 Vdd cclk idb7 GND efet w=2162 l=658
+ ad=0 pd=0 as=0 ps=0 
M5442 n_298 dor7 Vdd GND dfet w=1551 l=705
+ ad=0 pd=0 as=0 ps=0 
M5443 Vdd n_23 n_23 GND dfet w=846 l=752
+ ad=0 pd=0 as=1.41553e+07 ps=46624 
M5444 n_1501 n_23 Vdd GND dfet w=1598 l=658
+ ad=2.20281e+07 pd=51512 as=0 ps=0 
M5445 GND RnWstretched n_1501 GND efet w=8977 l=611
+ ad=0 pd=0 as=0 ps=0 
M5446 GND RnWstretched n_1501 GND efet w=18706 l=564
+ ad=0 pd=0 as=0 ps=0 
M5447 n_1501 dor7 GND GND efet w=13959 l=611
+ ad=0 pd=0 as=0 ps=0 
M5448 n_23 dor7 GND GND efet w=5640 l=658
+ ad=0 pd=0 as=0 ps=0 
M5449 dor7 dor7 Vdd GND dfet w=940 l=1128
+ ad=2.03935e+07 pd=63356 as=0 ps=0 
M5450 db5 n_612 GND GND efet w=19928 l=564
+ ad=0 pd=0 as=0 ps=0 
M5451 db5 n_373 Vdd GND efet w=60113 l=611
+ ad=0 pd=0 as=0 ps=0 
M5452 GND n_612 db5 GND efet w=1034 l=658
+ ad=0 pd=0 as=0 ps=0 
M5453 GND n_612 db5 GND efet w=21855 l=611
+ ad=0 pd=0 as=0 ps=0 
M5454 GND GND db5 GND efet w=5076 l=658
+ ad=0 pd=0 as=0 ps=0 
M5455 GND GND db6 GND efet w=5264 l=658
+ ad=0 pd=0 as=2.26034e+08 ps=409652 
M5456 n_254 n_254 Vdd GND dfet w=940 l=940
+ ad=1.87323e+06 pd=6768 as=0 ps=0 
M5457 n_869 abh5 GND GND efet w=13959 l=611
+ ad=1.03116e+07 pd=33276 as=0 ps=0 
M5458 Vdd n_1423 n_869 GND dfet w=1880 l=658
+ ad=0 pd=0 as=0 ps=0 
M5459 nABH5 cclk n_869 GND efet w=1128 l=752
+ ad=3.57858e+06 pd=11092 as=0 ps=0 
M5460 n_1353 ADH_ABH nABH5 GND efet w=1034 l=752
+ ad=485980 pd=3008 as=0 ps=0 
M5461 n_254 cp1 n_1353 GND efet w=1034 l=658
+ ad=8.64161e+06 pd=22560 as=0 ps=0 
M5462 GND adh5 n_254 GND efet w=7144 l=564
+ ad=0 pd=0 as=0 ps=0 
M5463 n_880 adh6 GND GND efet w=7144 l=658
+ ad=7.05996e+06 pd=23124 as=0 ps=0 
M5464 Vdd n_880 n_880 GND dfet w=846 l=846
+ ad=0 pd=0 as=1.82022e+06 ps=6580 
M5465 abh6 nABH6 GND GND efet w=6204 l=658
+ ad=5.16022e+06 pd=18048 as=0 ps=0 
M5466 Vdd abh6 abh6 GND dfet w=846 l=1316
+ ad=0 pd=0 as=1.87853e+07 ps=62228 
M5467 GND n_1523 n_963 GND efet w=10622 l=564
+ ad=0 pd=0 as=1.67884e+07 ps=37412 
M5468 n_963 abh6 Vdd GND dfet w=1598 l=658
+ ad=0 pd=0 as=0 ps=0 
M5469 Vdd n_1523 n_1523 GND dfet w=846 l=940
+ ad=0 pd=0 as=1.73097e+07 ps=62980 
M5470 GND abh6 n_1523 GND efet w=4277 l=611
+ ad=0 pd=0 as=4.49752e+06 ps=13536 
M5471 n_1514 cp1 n_880 GND efet w=1128 l=658
+ ad=530160 pd=3196 as=0 ps=0 
M5472 nABH6 ADH_ABH n_1514 GND efet w=1128 l=752
+ ad=3.55207e+06 pd=10340 as=0 ps=0 
M5473 n_635 cclk nABH6 GND efet w=1316 l=846
+ ad=1.04795e+07 pd=33652 as=0 ps=0 
M5474 Vdd n_1523 n_635 GND dfet w=1880 l=564
+ ad=0 pd=0 as=0 ps=0 
M5475 GND abh6 n_635 GND efet w=13865 l=611
+ ad=0 pd=0 as=0 ps=0 
M5476 GND n_869 ab13 GND efet w=3854 l=564
+ ad=0 pd=0 as=0 ps=0 
M5477 GND n_869 ab13 GND efet w=1222 l=564
+ ad=0 pd=0 as=0 ps=0 
M5478 GND n_869 ab13 GND efet w=15322 l=564
+ ad=0 pd=0 as=0 ps=0 
M5479 ab13 n_869 GND GND efet w=15322 l=564
+ ad=0 pd=0 as=0 ps=0 
M5480 GND n_869 ab13 GND efet w=15416 l=564
+ ad=0 pd=0 as=0 ps=0 
M5481 ab13 n_869 GND GND efet w=15416 l=752
+ ad=0 pd=0 as=0 ps=0 
M5482 GND n_869 ab13 GND efet w=15416 l=658
+ ad=0 pd=0 as=0 ps=0 
M5483 GND n_635 ab14 GND efet w=1222 l=470
+ ad=0 pd=0 as=1.648e+08 ps=218456 
M5484 GND n_635 ab14 GND efet w=3948 l=470
+ ad=0 pd=0 as=0 ps=0 
M5485 ab14 n_635 GND GND efet w=15416 l=564
+ ad=0 pd=0 as=0 ps=0 
M5486 GND n_635 ab14 GND efet w=15416 l=658
+ ad=0 pd=0 as=0 ps=0 
M5487 ab14 n_635 GND GND efet w=15416 l=564
+ ad=0 pd=0 as=0 ps=0 
M5488 GND n_635 ab14 GND efet w=15416 l=564
+ ad=0 pd=0 as=0 ps=0 
M5489 ab14 n_635 GND GND efet w=15416 l=564
+ ad=0 pd=0 as=0 ps=0 
M5490 Vdd n_963 ab14 GND efet w=39386 l=658
+ ad=0 pd=0 as=0 ps=0 
M5491 Vdd n_963 ab14 GND efet w=29798 l=564
+ ad=0 pd=0 as=0 ps=0 
M5492 Vdd n_963 ab14 GND efet w=15040 l=658
+ ad=0 pd=0 as=0 ps=0 
M5493 db6 n_7 Vdd GND efet w=13724 l=658
+ ad=0 pd=0 as=0 ps=0 
M5494 GND n_1153 n_1639 GND efet w=12314 l=564
+ ad=0 pd=0 as=1.8856e+07 ps=40420 
M5495 n_494 adh7 GND GND efet w=7144 l=658
+ ad=6.60049e+06 pd=21996 as=0 ps=0 
M5496 Vdd n_494 n_494 GND dfet w=940 l=940
+ ad=0 pd=0 as=2.04995e+06 ps=6956 
M5497 abh7 nABH7 GND GND efet w=6298 l=658
+ ad=4.60356e+06 pd=16732 as=0 ps=0 
M5498 Vdd abh7 abh7 GND dfet w=940 l=1175
+ ad=0 pd=0 as=1.77339e+07 ps=61852 
M5499 n_1639 abh7 Vdd GND dfet w=1598 l=564
+ ad=0 pd=0 as=0 ps=0 
M5500 Vdd n_1153 n_1153 GND dfet w=846 l=846
+ ad=0 pd=0 as=1.73274e+07 ps=62604 
M5501 GND abh7 n_1153 GND efet w=4418 l=564
+ ad=0 pd=0 as=4.6389e+06 ps=13536 
M5502 n_514 cp1 n_494 GND efet w=1128 l=658
+ ad=636192 pd=3384 as=0 ps=0 
M5503 nABH7 ADH_ABH n_514 GND efet w=1128 l=658
+ ad=3.42837e+06 pd=11280 as=0 ps=0 
M5504 n_659 cclk nABH7 GND efet w=1034 l=752
+ ad=1.00465e+07 pd=34592 as=0 ps=0 
M5505 Vdd n_1153 n_659 GND dfet w=1786 l=658
+ ad=0 pd=0 as=0 ps=0 
M5506 GND abh7 n_659 GND efet w=13959 l=611
+ ad=0 pd=0 as=0 ps=0 
M5507 ab15 n_659 GND GND efet w=16732 l=564
+ ad=1.7156e+08 pd=219396 as=0 ps=0 
M5508 GND n_659 ab15 GND efet w=4794 l=564
+ ad=0 pd=0 as=0 ps=0 
M5509 GND n_659 ab15 GND efet w=15228 l=564
+ ad=0 pd=0 as=0 ps=0 
M5510 ab15 n_659 GND GND efet w=15228 l=564
+ ad=0 pd=0 as=0 ps=0 
M5511 GND n_659 ab15 GND efet w=15228 l=564
+ ad=0 pd=0 as=0 ps=0 
M5512 ab15 n_659 GND GND efet w=15228 l=658
+ ad=0 pd=0 as=0 ps=0 
M5513 Vdd n_1639 ab15 GND efet w=38681 l=611
+ ad=0 pd=0 as=0 ps=0 
M5514 Vdd n_1639 ab15 GND efet w=29657 l=611
+ ad=0 pd=0 as=0 ps=0 
M5515 Vdd n_1639 ab15 GND efet w=15369 l=611
+ ad=0 pd=0 as=0 ps=0 
M5516 db6 n_471 db6 GND efet w=752 l=564
+ ad=0 pd=0 as=0 ps=0 
M5517 db6 n_7 Vdd GND efet w=44180 l=564
+ ad=0 pd=0 as=0 ps=0 
M5518 db6 n_471 GND GND efet w=20022 l=564
+ ad=0 pd=0 as=0 ps=0 
M5519 GND n_471 db6 GND efet w=846 l=564
+ ad=0 pd=0 as=0 ps=0 
M5520 db6 n_471 GND GND efet w=19834 l=564
+ ad=0 pd=0 as=0 ps=0 
M5521 db6 n_7 Vdd GND efet w=58891 l=611
+ ad=0 pd=0 as=0 ps=0 
M5522 GND n_471 db6 GND efet w=1034 l=564
+ ad=0 pd=0 as=0 ps=0 
M5523 db6 n_471 GND GND efet w=20210 l=564
+ ad=0 pd=0 as=0 ps=0 
M5524 GND n_471 db6 GND efet w=1034 l=564
+ ad=0 pd=0 as=0 ps=0 
M5525 db6 n_471 GND GND efet w=14100 l=564
+ ad=0 pd=0 as=0 ps=0 
M5526 db6 n_471 GND GND efet w=21573 l=611
+ ad=0 pd=0 as=0 ps=0 
M5527 GND GND db7 GND efet w=4371 l=705
+ ad=0 pd=0 as=2.51331e+08 ps=421684 
M5528 Vdd n_298 db7 GND efet w=27918 l=564
+ ad=0 pd=0 as=0 ps=0 
M5529 db7 n_1501 GND GND efet w=24581 l=611
+ ad=0 pd=0 as=0 ps=0 
M5530 Vdd n_298 db7 GND efet w=27589 l=611
+ ad=0 pd=0 as=0 ps=0 
M5531 Vdd n_298 db7 GND efet w=27542 l=658
+ ad=0 pd=0 as=0 ps=0 
M5532 Vdd n_298 db7 GND efet w=27354 l=658
+ ad=0 pd=0 as=0 ps=0 
M5533 GND n_1501 db7 GND efet w=24581 l=517
+ ad=0 pd=0 as=0 ps=0 
M5534 db7 n_1501 GND GND efet w=24628 l=564
+ ad=0 pd=0 as=0 ps=0 
M5535 db7 n_1501 GND GND efet w=24581 l=611
+ ad=0 pd=0 as=0 ps=0 
C0 metal_351842_6674# gnd! 3.2fF ;**FLOATING
C1 metal_349868_6674# gnd! 3.2fF ;**FLOATING
C2 metal_342630_7238# gnd! 16.7fF ;**FLOATING
C3 metal_351842_10152# gnd! 3.2fF ;**FLOATING
C4 metal_349868_9024# gnd! 3.2fF ;**FLOATING
C5 metal_23688_7896# gnd! 18.9fF ;**FLOATING
C6 testpad_8 gnd! 101.5fF ;**FLOATING
C7 metal_162902_194862# gnd! 125.6fF ;**FLOATING
C8 metal_72568_216576# gnd! 15.4fF ;**FLOATING
C9 metal_152750_223626# gnd! 100.2fF ;**FLOATING
C10 metal_74260_220712# gnd! 6.9fF ;**FLOATING
C11 metal_72568_220712# gnd! 7.6fF ;**FLOATING
C12 metal_80182_238760# gnd! 22.0fF ;**FLOATING
C13 metal_242990_287452# gnd! 120.9fF ;**FLOATING
C14 pad_nc1 gnd! 330.2fF ;**FLOATING
C15 diff_348082_6674# gnd! 4.2fF ;**FLOATING
C16 diff_346014_6674# gnd! 4.4fF ;**FLOATING
C17 n_915 gnd! 21.2fF ;**FLOATING
C18 n_749 gnd! 20.5fF ;**FLOATING
C19 diff_348082_10246# gnd! 3.2fF ;**FLOATING
C20 diff_346014_9118# gnd! 4.1fF ;**FLOATING
C21 n_1208 gnd! 22.7fF ;**FLOATING
C22 n_908 gnd! 22.7fF ;**FLOATING
C23 n_144 gnd! 76.6fF ;**FLOATING
C24 ab15 gnd! 2566.8fF
C25 n_659 gnd! 421.1fF
C26 n_514 gnd! 9.7fF
C27 n_1639 gnd! 514.2fF
C28 abh7 gnd! 171.1fF
C29 n_494 gnd! 101.5fF
C30 n_1153 gnd! 149.5fF
C31 nABH7 gnd! 77.3fF
C32 ab14 gnd! 2450.1fF
C33 n_635 gnd! 413.4fF
C34 n_1514 gnd! 8.5fF
C35 n_963 gnd! 499.2fF
C36 n_1523 gnd! 149.6fF
C37 abh6 gnd! 182.0fF
C38 n_1353 gnd! 7.9fF
C39 n_869 gnd! 432.7fF
C40 n_880 gnd! 105.0fF
C41 nABH6 gnd! 76.9fF
C42 n_1501 gnd! 734.9fF
C43 n_23 gnd! 162.4fF
C44 n_298 gnd! 753.5fF
C45 n_588 gnd! 203.9fF
C46 dor7 gnd! 225.5fF
C47 notdor7 gnd! 52.8fF
C48 n_789 gnd! 126.4fF
C49 notidl7 gnd! 83.1fF
C50 idl7 gnd! 167.0fF
C51 n_471 gnd! 734.4fF
C52 n_466 gnd! 162.4fF
C53 n_7 gnd! 785.0fF
C54 n_1147 gnd! 271.1fF
C55 n_1638 gnd! 211.6fF
C56 dor6 gnd! 215.8fF
C57 notdor6 gnd! 48.6fF
C58 n_1684 gnd! 117.9fF
C59 notidl6 gnd! 84.4fF
C60 idl6 gnd! 170.9fF
C61 n_612 gnd! 656.5fF
C62 n_1720 gnd! 154.0fF
C63 n_373 gnd! 755.2fF
C64 n_542 gnd! 600.1fF ;**FLOATING
C65 n_1014 gnd! 266.0fF
C66 n_568 gnd! 212.3fF
C67 dor5 gnd! 227.5fF
C68 notdor5 gnd! 51.8fF
C69 n_961 gnd! 117.9fF
C70 notidl5 gnd! 89.0fF
C71 idl5 gnd! 167.9fF
C72 n_147 gnd! 691.9fF
C73 n_1463 gnd! 157.7fF
C74 n_1076 gnd! 747.1fF
C75 n_254 gnd! 120.0fF
C76 ab13 gnd! 2412.3fF
C77 ab12 gnd! 2457.8fF
C78 n_999 gnd! 416.4fF
C79 n_1451 gnd! 7.2fF
C80 n_1608 gnd! 478.5fF
C81 n_475 gnd! 479.8fF
C82 abh5 gnd! 187.4fF
C83 nABH5 gnd! 78.6fF
C84 n_1423 gnd! 153.6fF
C85 n_1677 gnd! 162.1fF
C86 abh4 gnd! 177.7fF
C87 n_212 gnd! 106.6fF
C88 nABH4 gnd! 76.8fF
C89 n_1667 gnd! 7.9fF
C90 n_359 gnd! 424.0fF
C91 n_883 gnd! 118.6fF
C92 nABH3 gnd! 73.6fF
C93 ab11 gnd! 2430.4fF
C94 ab10 gnd! 2460.7fF
C95 n_994 gnd! 429.6fF
C96 n_836 gnd! 8.5fF
C97 n_1296 gnd! 498.9fF
C98 n_1545 gnd! 496.5fF
C99 abh3 gnd! 191.1fF
C100 n_1346 gnd! 140.5fF
C101 n_1034 gnd! 145.9fF
C102 abh2 gnd! 176.3fF
C103 n_1298 gnd! 9.7fF
C104 n_676 gnd! 427.5fF
C105 n_168 gnd! 110.4fF
C106 nABH2 gnd! 76.8fF
C107 n_1387 gnd! 268.4fF
C108 n_490 gnd! 203.6fF
C109 dor4 gnd! 215.3fF
C110 notdor4 gnd! 48.7fF
C111 n_797 gnd! 117.3fF
C112 notidl4 gnd! 87.1fF
C113 idl4 gnd! 162.1fF
C114 n_643 gnd! 653.1fF
C115 n_1613 gnd! 155.2fF
C116 n_42 gnd! 749.8fF
C117 n_1095 gnd! 267.7fF
C118 n_896 gnd! 203.6fF
C119 dor3 gnd! 223.0fF
C120 notdor3 gnd! 51.8fF
C121 n_457 gnd! 126.7fF
C122 notidl3 gnd! 83.9fF
C123 idl3 gnd! 162.3fF
C124 n_37 gnd! 688.3fF
C125 n_224 gnd! 160.5fF
C126 n_520 gnd! 710.7fF
C127 n_1661 gnd! 262.0fF
C128 n_1199 gnd! 201.4fF
C129 dor2 gnd! 221.4fF
C130 notdor2 gnd! 51.5fF
C131 n_1376 gnd! 120.8fF
C132 notidl2 gnd! 81.4fF
C133 idl2 gnd! 167.3fF
C134 n_794 gnd! 678.8fF
C135 n_288 gnd! 156.2fF
C136 n_798 gnd! 709.0fF
C137 n_1424 gnd! 271.6fF
C138 n_213 gnd! 211.6fF
C139 dor1 gnd! 213.7fF
C140 pclp7 gnd! 211.6fF
C141 n_914 gnd! 136.9fF
C142 n_484 gnd! 143.1fF
C143 npclp7 gnd! 59.7fF
C144 n_1386 gnd! 109.7fF
C145 n_426 gnd! 54.0fF
C146 pcl7 gnd! 121.2fF
C147 n_641 gnd! 110.4fF
C148 notdor1 gnd! 53.4fF
C149 n_1474 gnd! 116.0fF
C150 notidl1 gnd! 88.1fF
C151 idl1 gnd! 166.1fF
C152 n_769 gnd! 157.6fF
C153 n_87 gnd! 260.4fF
C154 n_1325 gnd! 705.6fF
C155 n_1072 gnd! 654.7fF
C156 n_718 gnd! 201.2fF
C157 dor0 gnd! 212.9fF
C158 notdor0 gnd! 51.6fF
C159 n_1687 gnd! 121.1fF
C160 notidl0 gnd! 83.5fF
C161 idl0 gnd! 170.9fF
C162 n_715 gnd! 209.1fF
C163 pcl6 gnd! 107.3fF
C164 n_993 gnd! 40.0fF
C165 n_1264 gnd! 32.7fF
C166 n_663 gnd! 39.4fF
C167 n_1213 gnd! 171.9fF
C168 n_453 gnd! 157.3fF
C169 n_1209 gnd! 117.5fF
C170 npchp7 gnd! 153.3fF
C171 pchp7 gnd! 227.8fF
C172 n_1316 gnd! 228.7fF
C173 pclp6 gnd! 227.5fF
C174 npclp6 gnd! 143.4fF
C175 n_585 gnd! 25.5fF
C176 n_20 gnd! 125.2fF
C177 n_232 gnd! 181.4fF
C178 pclp5 gnd! 213.3fF
C179 n_557 gnd! 138.9fF
C180 n_1547 gnd! 139.1fF
C181 n_278 gnd! 84.1fF
C182 n_545 gnd! 48.7fF
C183 n_1192 gnd! 143.7fF
C184 npchp6 gnd! 56.1fF
C185 n_609 gnd! 153.5fF
C186 n_1488 gnd! 200.5fF
C187 n_1073 gnd! 152.1fF
C188 npclp5 gnd! 56.5fF
C189 n_344 gnd! 159.3fF
C190 n_814 gnd! 48.7fF
C191 pcl5 gnd! 124.8fF
C192 n_386 gnd! 101.5fF
C193 pch7 gnd! 127.4fF
C194 pchp6 gnd! 218.4fF
C195 pch6 gnd! 144.2fF
C196 n_1659 gnd! 32.7fF
C197 n_469 gnd! 40.4fF
C198 n_743 gnd! 220.3fF
C199 n_499 gnd! 182.8fF
C200 n_875 gnd! 118.3fF
C201 npchp5 gnd! 147.0fF
C202 n_392 gnd! 210.1fF
C203 pcl4 gnd! 106.3fF
C204 n_15 gnd! 37.7fF
C205 n_410 gnd! 223.1fF
C206 pclp4 gnd! 217.5fF
C207 npclp4 gnd! 143.7fF
C208 n_766 gnd! 29.1fF
C209 n_474 gnd! 119.8fF
C210 n_1643 gnd! 178.4fF
C211 pclp3 gnd! 212.0fF
C212 n_903 gnd! 146.8fF
C213 n_1631 gnd! 154.0fF
C214 npclp3 gnd! 57.2fF
C215 n_1184 gnd! 160.3fF
C216 n_1498 gnd! 52.4fF
C217 pcl3 gnd! 124.1fF
C218 n_249 gnd! 115.9fF
C219 n_719 gnd! 265.2fF
C220 n_1585 gnd! 92.8fF
C221 RnWstretched gnd! 2566.1fF
C222 n_221 gnd! 214.6fF
C223 n_1028 gnd! 126.2fF
C224 n_251 gnd! 462.4fF
C225 n_962 gnd! 131.6fF
C226 n_1579 gnd! 52.6fF
C227 nDBE gnd! 247.3fF
C228 n_1293 gnd! 198.4fF
C229 n_802 gnd! 32.8fF
C230 n_1371 gnd! 185.1fF
C231 n_201 gnd! 236.2fF
C232 p1 gnd! 53.7fF
C233 n_661 gnd! 90.4fF
C234 n_163 gnd! 210.8fF
C235 pcl2 gnd! 108.0fF
C236 n_1411 gnd! 40.1fF
C237 n_1253 gnd! 215.7fF
C238 pclp2 gnd! 225.2fF
C239 npclp2 gnd! 151.8fF
C240 n_1158 gnd! 25.5fF
C241 n_515 gnd! 122.1fF
C242 pchp5 gnd! 219.5fF
C243 n_1406 gnd! 137.0fF
C244 n_1400 gnd! 83.4fF
C245 n_949 gnd! 51.1fF
C246 n_1657 gnd! 146.9fF
C247 npchp4 gnd! 52.9fF
C248 n_523 gnd! 153.6fF
C249 n_83 gnd! 213.3fF
C250 pch5 gnd! 129.8fF
C251 pchp4 gnd! 218.6fF
C252 n_356 gnd! 36.8fF
C253 n_1061 gnd! 40.8fF
C254 n_810 gnd! 163.5fF
C255 n_923 gnd! 176.3fF
C256 n_207 gnd! 119.2fF
C257 npchp3 gnd! 153.0fF
C258 pch4 gnd! 148.7fF
C259 pchp3 gnd! 225.4fF
C260 pch3 gnd! 125.7fF
C261 n_783 gnd! 178.1fF
C262 pclp1 gnd! 211.0fF
C263 n_1568 gnd! 138.8fF
C264 n_1099 gnd! 148.2fF
C265 npclp1 gnd! 58.7fF
C266 n_1542 gnd! 166.4fF
C267 n_1685 gnd! 52.3fF
C268 pcl1 gnd! 124.0fF
C269 n_329 gnd! 105.8fF
C270 n_57 gnd! 141.5fF
C271 n_1265 gnd! 102.3fF
C272 adh7 gnd! 496.2fF
C273 pchp2 gnd! 213.2fF
C274 n_1402 gnd! 114.9fF
C275 npchp2 gnd! 43.8fF
C276 n_1367 gnd! 49.4fF
C277 n_293 gnd! 156.3fF
C278 n_1166 gnd! 212.5fF
C279 pcl0 gnd! 112.7fF
C280 n_526 gnd! 39.8fF
C281 n_1345 gnd! 221.7fF
C282 pclp0 gnd! 219.4fF
C283 npclp0 gnd! 138.8fF
C284 n_1706 gnd! 26.1fF
C285 n_1500 gnd! 118.9fF
C286 n_937 gnd! 178.0fF
C287 n_580 gnd! 48.6fF
C288 n_566 gnd! 215.5fF
C289 pipeUNK14 gnd! 52.5fF
C290 n_1170 gnd! 116.1fF
C291 nDBZ gnd! 185.4fF
C292 n_1115 gnd! 109.3fF
C293 n_922 gnd! 52.0fF
C294 n_620 gnd! 319.6fF
C295 n_1433 gnd! 195.1fF
C296 pipeUNK15 gnd! 49.6fF
C297 n_243 gnd! 251.2fF
C298 DBZ gnd! 414.2fF
C299 dpc43_DL_DB gnd! 531.4fF
C300 n_1202 gnd! 211.3fF
C301 pch2 gnd! 157.0fF
C302 n_1538 gnd! 32.0fF
C303 n_126 gnd! 40.1fF
C304 n_200 gnd! 222.6fF
C305 n_1070 gnd! 185.5fF
C306 n_1486 gnd! 115.2fF
C307 npchp1 gnd! 147.0fF
C308 n_835 gnd! 148.5fF
C309 adh6 gnd! 563.9fF
C310 n_128 gnd! 134.2fF
C311 n_1592 gnd! 198.9fF
C312 n_569 gnd! 23.6fF
C313 n_260 gnd! 119.2fF
C314 a7 gnd! 72.8fF
C315 adh5 gnd! 596.6fF
C316 n_1356 gnd! 132.2fF
C317 n_1454 gnd! 27.0fF
C318 n_100 gnd! 35.8fF
C319 n_1205 gnd! 186.8fF
C320 n_852 gnd! 108.0fF
C321 dasb7 gnd! 96.3fF
C322 n_1018 gnd! 105.5fF
C323 n_711 gnd! 25.5fF
C324 n_1080 gnd! 23.0fF
C325 n_479 gnd! 118.9fF
C326 n_326 gnd! 210.2fF
C327 a6 gnd! 78.9fF
C328 adh4 gnd! 879.4fF
C329 n_1719 gnd! 128.4fF
C330 n_1554 gnd! 27.0fF
C331 n_739 gnd! 183.8fF
C332 n_61 gnd! 108.5fF
C333 dasb6 gnd! 94.4fF
C334 n_1056 gnd! 91.3fF
C335 n_1629 gnd! 114.1fF
C336 n_831 gnd! 211.6fF
C337 a5 gnd! 78.9fF
C338 adh3 gnd! 822.5fF
C339 n_556 gnd! 134.7fF
C340 n_1344 gnd! 206.2fF
C341 n_1203 gnd! 35.0fF
C342 n_408 gnd! 100.1fF
C343 n_1267 gnd! 116.6fF
C344 ab9 gnd! 2416.2fF
C345 diff_25568_7426# gnd! 20.7fF ;**FLOATING
C346 diff_23218_7426# gnd! 19.3fF ;**FLOATING
C347 diff_25568_10058# gnd! 17.1fF ;**FLOATING
C348 n_290 gnd! 16.0fF ;**FLOATING
C349 n_1461 gnd! 18.4fF ;**FLOATING
C350 diff_23218_11280# gnd! 17.6fF ;**FLOATING
C351 diff_25568_13912# gnd! 18.0fF ;**FLOATING
C352 diff_23218_13160# gnd! 17.4fF ;**FLOATING
C353 diff_25568_15134# gnd! 18.0fF ;**FLOATING
C354 diff_23218_15134# gnd! 17.4fF ;**FLOATING
C355 diff_25568_17766# gnd! 18.0fF ;**FLOATING
C356 n_30 gnd! 17.4fF ;**FLOATING
C357 ab8 gnd! 2393.4fF
C358 n_381 gnd! 448.0fF
C359 ab7 gnd! 2644.8fF
C360 n_705 gnd! 9.0fF
C361 n_826 gnd! 489.6fF
C362 n_1140 gnd! 492.2fF
C363 abh1 gnd! 195.2fF
C364 nABH1 gnd! 78.8fF
C365 n_617 gnd! 145.3fF
C366 n_1315 gnd! 164.8fF
C367 alu7 gnd! 160.9fF
C368 notalu7 gnd! 65.1fF
C369 n_762 gnd! 181.8fF
C370 n_1135 gnd! 205.3fF
C371 dasb5 gnd! 94.7fF
C372 n_970 gnd! 46.5fF
C373 n_149 gnd! 143.6fF
C374 n_233 gnd! 243.4fF
C375 n_761 gnd! 237.9fF
C376 n_838 gnd! 119.0fF
C377 a4 gnd! 71.5fF
C378 n_753 gnd! 178.8fF
C379 n_811 gnd! 284.8fF
C380 n_947 gnd! 132.5fF
C381 n_581 gnd! 43.1fF
C382 n_306 gnd! 110.8fF
C383 n_393 gnd! 38.0fF
C384 n_551 gnd! 139.7fF
C385 n_1279 gnd! 29.1fF
C386 n_1097 gnd! 113.4fF
C387 n_1654 gnd! 222.0fF
C388 a3 gnd! 76.0fF
C389 pchp1 gnd! 228.6fF
C390 pch1 gnd! 124.6fF
C391 n_1010 gnd! 98.2fF
C392 pchp0 gnd! 207.1fF
C393 n_1229 gnd! 125.8fF
C394 npchp0 gnd! 47.3fF
C395 n_856 gnd! 53.3fF
C396 n_919 gnd! 157.9fF
C397 pch0 gnd! 143.5fF
C398 n_311 gnd! 209.4fF
C399 adh1 gnd! 955.4fF
C400 n_419 gnd! 131.8fF
C401 n_1686 gnd! 22.4fF
C402 n_1584 gnd! 34.8fF
C403 n_1179 gnd! 174.3fF
C404 n_345 gnd! 178.2fF
C405 n_432 gnd! 153.9fF
C406 dasb3 gnd! 99.7fF
C407 n_1159 gnd! 103.2fF
C408 n_1618 gnd! 218.1fF
C409 a2 gnd! 73.0fF
C410 n_1656 gnd! 26.9fF
C411 n_1580 gnd! 116.7fF
C412 dasb2 gnd! 106.1fF
C413 n_1549 gnd! 128.7fF
C414 n_929 gnd! 210.4fF
C415 n_619 gnd! 34.7fF
C416 n_695 gnd! 120.0fF
C417 n_735 gnd! 108.0fF
C418 a1 gnd! 73.1fF
C419 n_1322 gnd! 26.3fF
C420 n_320 gnd! 103.9fF
C421 dasb1 gnd! 100.9fF
C422 n_5 gnd! 133.9fF
C423 a0 gnd! 67.9fF
C424 dpc41_DL_ADL gnd! 609.2fF
C425 dpc42_DL_ADH gnd! 582.7fF
C426 Pout1 gnd! 153.3fF
C427 Pout0 gnd! 155.8fF
C428 n_318 gnd! 393.2fF
C429 n_846 gnd! 235.3fF
C430 n_1625 gnd! 52.9fF
C431 n_307 gnd! 219.1fF
C432 pipeUNK05 gnd! 65.1fF
C433 n_1616 gnd! 60.0fF
C434 n_69 gnd! 50.6fF
C435 n_1445 gnd! 21.1fF
C436 n_1546 gnd! 24.1fF
C437 n_1470 gnd! 24.1fF
C438 pipeUNK13 gnd! 47.9fF
C439 n_793 gnd! 62.4fF
C440 n_1595 gnd! 93.0fF
C441 n_1181 gnd! 200.2fF
C442 n_1614 gnd! 239.2fF
C443 pipeUNK03 gnd! 85.3fF
C444 n_1723 gnd! 64.4fF
C445 n_1177 gnd! 61.2fF
C446 n_299 gnd! 236.0fF
C447 n_648 gnd! 34.1fF
C448 n_1644 gnd! 75.4fF
C449 n_1457 gnd! 153.6fF
C450 n_1495 gnd! 193.9fF
C451 p3 gnd! 50.1fF
C452 pipeUNK04 gnd! 65.2fF
C453 db6 gnd! 4084.6fF
C454 db2 gnd! 3674.4fF
C455 n_1492 gnd! 201.5fF
C456 db0 gnd! 4829.9fF
C457 db5 gnd! 4363.2fF
C458 pipeUNK02 gnd! 35.4fF
C459 p4 gnd! 190.2fF
C460 n_1471 gnd! 119.6fF
C461 p0 gnd! 49.7fF
C462 n_455 gnd! 44.9fF
C463 p6 gnd! 148.5fF
C464 n_1240 gnd! 101.4fF
C465 n_1441 gnd! 112.9fF
C466 n_1157 gnd! 98.3fF
C467 dpc35_PCHC gnd! 598.7fF
C468 H1x1 gnd! 363.1fF
C469 n_1416 gnd! 364.8fF
C470 n_1600 gnd! 290.2fF
C471 n_90 gnd! 346.5fF
C472 p7 gnd! 145.5fF
C473 Pout2 gnd! 148.4fF
C474 n_1566 gnd! 142.2fF
C475 dpc40_ADLPCL gnd! 631.0fF
C476 n_146 gnd! 220.7fF
C477 n_1341 gnd! 49.5fF
C478 n_876 gnd! 146.2fF
C479 n_1362 gnd! 55.3fF
C480 n_600 gnd! 325.8fF
C481 n_150 gnd! 43.2fF
C482 n_613 gnd! 271.2fF
C483 n_867 gnd! 166.1fF
C484 n_8 gnd! 260.0fF
C485 n_1682 gnd! 79.2fF
C486 n_986 gnd! 217.3fF
C487 n_1556 gnd! 28.0fF
C488 nDA_ADD2 gnd! 155.5fF
C489 nDA_ADD1 gnd! 178.3fF
C490 notalu6 gnd! 59.1fF
C491 alu6 gnd! 234.2fF
C492 C78 gnd! 138.0fF
C493 C78_phi2 gnd! 36.9fF
C494 DC78_phi2 gnd! 38.6fF
C495 notaluvout gnd! 158.1fF
C496 adh2 gnd! 1013.0fF
C497 n_637 gnd! 122.0fF
C498 n_1489 gnd! 65.2fF
C499 notalu5 gnd! 61.4fF
C500 alu5 gnd! 238.5fF
C501 notalu4 gnd! 60.2fF
C502 alu4 gnd! 198.9fF
C503 notalu3 gnd! 59.5fF
C504 alu3 gnd! 192.7fF
C505 notalu2 gnd! 58.4fF
C506 alu2 gnd! 255.9fF
C507 dpc38_PCLADL gnd! 567.3fF
C508 dpc39_PCLPCL gnd! 596.7fF
C509 dpc32_PCHADH gnd! 522.8fF
C510 dpc37_PCLDB gnd! 507.1fF
C511 n_1007 gnd! 92.8fF
C512 dpc34_PCLC gnd! 1031.4fF
C513 n_1043 gnd! 105.1fF
C514 n_1462 gnd! 99.5fF
C515 dpc33_PCHDB gnd! 492.1fF
C516 n_36 gnd! 187.0fF
C517 n_1277 gnd! 142.8fF
C518 n_291 gnd! 156.5fF
C519 n_1221 gnd! 52.4fF
C520 n_1020 gnd! 52.0fF
C521 n_1121 gnd! 50.3fF
C522 n_1045 gnd! 500.0fF
C523 n_186 gnd! 20.5fF
C524 n_367 gnd! 40.3fF
C525 n_1224 gnd! 223.7fF
C526 pipeUNK16 gnd! 69.4fF
C527 n_756 gnd! 80.5fF
C528 n_1110 gnd! 273.9fF
C529 n_626 gnd! 138.5fF
C530 pipeUNK12 gnd! 41.7fF
C531 n_1198 gnd! 68.7fF
C532 n_1249 gnd! 81.8fF
C533 pipeUNK01 gnd! 46.5fF
C534 n_755 gnd! 297.3fF
C535 n_1692 gnd! 24.8fF
C536 n_1082 gnd! 335.8fF
C537 n_279 gnd! 190.0fF
C538 n_507 gnd! 128.2fF
C539 n_1049 gnd! 46.2fF
C540 n_1194 gnd! 343.9fF
C541 n_160 gnd! 135.5fF
C542 db4 gnd! 4125.7fF
C543 n_374 gnd! 175.4fF
C544 n_111 gnd! 171.1fF
C545 n_62 gnd! 167.2fF
C546 db7 gnd! 4555.5fF
C547 db1 gnd! 4967.1fF
C548 n_1319 gnd! 173.0fF
C549 n_93 gnd! 183.3fF
C550 n_1588 gnd! 182.1fF
C551 n_1281 gnd! 171.4fF
C552 db3 gnd! 3983.1fF
C553 n_1075 gnd! 171.8fF
C554 n_587 gnd! 243.6fF
C555 n_503 gnd! 89.6fF
C556 n_340 gnd! 89.1fF
C557 pd4 gnd! 59.0fF
C558 n_1214 gnd! 108.6fF
C559 n_1401 gnd! 127.5fF
C560 n_1269 gnd! 74.6fF
C561 DBNeg gnd! 497.7fF
C562 n_1673 gnd! 40.8fF
C563 n_754 gnd! 420.5fF
C564 n_1422 gnd! 63.7fF
C565 pipeUNK06 gnd! 82.0fF
C566 n_1111 gnd! 333.8fF
C567 pipeUNK11 gnd! 51.6fF
C568 pipeUNK07 gnd! 46.2fF
C569 n_941 gnd! 59.3fF
C570 pipeUNK09 gnd! 176.6fF
C571 n_954 gnd! 343.8fF
C572 pipeUNK08 gnd! 57.0fF
C573 n_818 gnd! 153.2fF
C574 n_1518 gnd! 100.7fF
C575 n_1413 gnd! 99.5fF
C576 dpc31_PCHPCH gnd! 573.0fF
C577 n_1323 gnd! 94.6fF
C578 n_849 gnd! 99.6fF
C579 dpc30_ADHPCH gnd! 592.8fF
C580 n_AxB7__C67 gnd! 93.2fF
C581 DC78 gnd! 188.7fF
C582 n_AxBxC_7 gnd! 117.7fF
C583 n_1013 gnd! 23.0fF
C584 n_AxB_7 gnd! 75.7fF
C585 nC78 gnd! 156.8fF
C586 n_1617 gnd! 37.5fF
C587 n_1030 gnd! 202.0fF
C588 nC67 gnd! 88.5fF
C589 n_269 gnd! 119.6fF
C590 AxB7 gnd! 238.8fF
C591 A_B7 gnd! 115.7fF
C592 n_748 gnd! 153.4fF
C593 n_A_B_7 gnd! 280.7fF
C594 naluresult7 gnd! 268.1fF
C595 _AxB_6_nC56 gnd! 106.2fF
C596 n_1038 gnd! 85.0fF
C597 n_AxBxC_6 gnd! 116.5fF
C598 n_1390 gnd! 23.0fF
C599 n_112 gnd! 40.3fF
C600 C67 gnd! 234.4fF
C601 n_482 gnd! 25.5fF
C602 n_AxB_6 gnd! 250.0fF
C603 C56 gnd! 98.4fF
C604 nA_B7 gnd! 272.3fF
C605 n_1695 gnd! 44.9fF
C606 alua7 gnd! 107.7fF
C607 n_423 gnd! 129.9fF
C608 idb7 gnd! 1102.7fF
C609 alub7 gnd! 161.3fF
C610 n_A_B_6 gnd! 221.0fF
C611 naluresult6 gnd! 335.3fF
C612 A_B6 gnd! 101.4fF
C613 n_570 gnd! 257.7fF
C614 n_AxB5__C45 gnd! 98.3fF
C615 n_122 gnd! 122.7fF
C616 n_1257 gnd! 369.7fF
C617 n_AxBxC_5 gnd! 119.8fF
C618 n_547 gnd! 26.3fF
C619 n_AxB_5 gnd! 75.7fF
C620 nC56 gnd! 158.9fF
C621 n_165 gnd! 40.4fF
C622 AxB5 gnd! 205.9fF
C623 n_939 gnd! 44.1fF
C624 n_757 gnd! 225.7fF
C625 notalucout gnd! 295.3fF
C626 alucout gnd! 717.5fF
C627 A_B5 gnd! 109.5fF
C628 n_647 gnd! 235.5fF
C629 nC45 gnd! 152.2fF
C630 _AxB_4_nC34 gnd! 105.4fF
C631 DA_C45 gnd! 119.4fF
C632 n_AxBxC_4 gnd! 124.4fF
C633 n_375 gnd! 26.3fF
C634 n_1310 gnd! 35.6fF
C635 C45 gnd! 150.4fF
C636 n_1583 gnd! 24.8fF
C637 nA_B6 gnd! 311.5fF
C638 n_1483 gnd! 44.9fF
C639 alua6 gnd! 105.9fF
C640 n_351 gnd! 128.9fF
C641 idb6 gnd! 1086.2fF
C642 alub6 gnd! 159.4fF
C643 s7 gnd! 66.8fF
C644 nots7 gnd! 51.3fF
C645 n_548 gnd! 122.5fF
C646 n_721 gnd! 262.7fF
C647 n_A_B_5 gnd! 215.8fF
C648 naluresult5 gnd! 357.7fF
C649 nA_B5 gnd! 206.2fF
C650 n_1559 gnd! 39.4fF
C651 alua5 gnd! 109.8fF
C652 n_AxB_4 gnd! 177.5fF
C653 n_1218 gnd! 137.3fF
C654 C34 gnd! 244.3fF
C655 n_1565 gnd! 50.5fF
C656 n_700 gnd! 214.0fF
C657 notalu1 gnd! 61.2fF
C658 alu1 gnd! 242.7fF
C659 notalu0 gnd! 60.7fF
C660 alu0 gnd! 200.8fF
C661 n_972 gnd! 189.8fF
C662 n_1383 gnd! 128.0fF
C663 idb5 gnd! 1015.4fF
C664 alub5 gnd! 155.1fF
C665 n_A_B_4 gnd! 219.5fF
C666 naluresult4 gnd! 328.0fF
C667 A_B4 gnd! 100.7fF
C668 DC34 gnd! 209.6fF
C669 n_AxB3__C23 gnd! 99.6fF
C670 n_AxBxC_3 gnd! 116.1fF
C671 n_136 gnd! 26.3fF
C672 nC34 gnd! 177.3fF
C673 n_924 gnd! 39.2fF
C674 n_AxB_3 gnd! 77.5fF
C675 nC23 gnd! 91.8fF
C676 A_B3 gnd! 110.3fF
C677 n_988 gnd! 152.9fF
C678 nA_B4 gnd! 248.6fF
C679 n_185 gnd! 44.9fF
C680 alua4 gnd! 101.5fF
C681 n_478 gnd! 123.4fF
C682 idb4 gnd! 1004.3fF
C683 alub4 gnd! 154.4fF
C684 n_A_B_3 gnd! 225.0fF
C685 naluresult3 gnd! 364.9fF
C686 _AxB_2_nC12 gnd! 120.9fF
C687 n_1610 gnd! 176.6fF
C688 AxB3 gnd! 277.1fF
C689 DA_AB2 gnd! 195.7fF
C690 n_AxBxC_2 gnd! 129.2fF
C691 n_1572 gnd! 27.0fF
C692 n_433 gnd! 59.4fF
C693 C23 gnd! 164.7fF
C694 n_716 gnd! 25.3fF
C695 n_AxB_2 gnd! 166.0fF
C696 nA_B3 gnd! 209.5fF
C697 n_313 gnd! 44.9fF
C698 alua3 gnd! 106.8fF
C699 n_1621 gnd! 124.8fF
C700 idb3 gnd! 990.3fF
C701 alub3 gnd! 153.3fF
C702 n_A_B_2 gnd! 348.0fF
C703 naluresult2 gnd! 332.9fF
C704 C12 gnd! 82.2fF
C705 A_B2 gnd! 76.1fF
C706 n_AxB1__C01 gnd! 97.4fF
C707 DA_AxB2 gnd! 186.3fF
C708 n_388 gnd! 307.5fF
C709 n_AxBxC_1 gnd! 118.2fF
C710 n_1388 gnd! 26.3fF
C711 n_AxB_1 gnd! 75.1fF
C712 nC12 gnd! 162.0fF
C713 n_1510 gnd! 39.2fF
C714 n_1354 gnd! 34.3fF
C715 n_319 gnd! 244.0fF
C716 n_1707 gnd! 39.9fF
C717 AxB1 gnd! 209.7fF
C718 nC01 gnd! 87.2fF
C719 n_936 gnd! 236.5fF
C720 A_B1 gnd! 108.5fF
C721 _AxB_0_nC0in gnd! 123.2fF
C722 DA_C01 gnd! 170.0fF
C723 dpc26_ACDB gnd! 605.0fF
C724 n_1369 gnd! 151.5fF
C725 n_1270 gnd! 157.5fF
C726 n_1260 gnd! 144.8fF
C727 n_255 gnd! 93.7fF
C728 n_631 gnd! 150.4fF
C729 n_228 gnd! 99.7fF
C730 dpc24_ACSB gnd! 522.9fF
C731 dpc29_0ADH17 gnd! 569.2fF
C732 dpc27_SBADH gnd! 485.1fF
C733 n_800 gnd! 96.2fF
C734 n_321 gnd! 145.7fF
C735 n_1335 gnd! 91.9fF
C736 dpc23_SBAC gnd! 531.5fF
C737 dpc25_SBDB gnd! 541.5fF
C738 n_1635 gnd! 95.8fF
C739 n_265 gnd! 42.7fF
C740 n_897 gnd! 49.8fF
C741 n_611 gnd! 155.9fF
C742 n_21 gnd! 160.4fF
C743 n_525 gnd! 159.1fF
C744 n_598 gnd! 51.8fF
C745 n_878 gnd! 53.9fF
C746 n_509 gnd! 38.8fF
C747 n_398 gnd! 52.6fF
C748 n_1509 gnd! 40.8fF
C749 n_1162 gnd! 40.0fF
C750 n_266 gnd! 40.1fF
C751 n_1271 gnd! 99.0fF
C752 n_628 gnd! 146.1fF
C753 n_1047 gnd! 95.7fF
C754 n_1238 gnd! 100.5fF
C755 n_966 gnd! 148.9fF
C756 n_1596 gnd! 152.5fF
C757 n_830 gnd! 158.5fF
C758 n_1295 gnd! 153.6fF
C759 n_55 gnd! 43.2fF
C760 n_1683 gnd! 50.3fF
C761 n_1602 gnd! 48.4fF
C762 n_1505 gnd! 42.8fF
C763 n_1527 gnd! 51.7fF
C764 n_1581 gnd! 73.2fF
C765 n_1480 gnd! 361.6fF
C766 dpc36_nIPC gnd! 340.4fF
C767 n_1275 gnd! 195.4fF
C768 n_1570 gnd! 70.9fF
C769 n_1472 gnd! 85.5fF
C770 pipeBRtaken gnd! 88.0fF
C771 n_1446 gnd! 138.6fF
C772 n_465 gnd! 141.8fF
C773 pipeUNK20 gnd! 74.5fF
C774 n_850 gnd! 149.4fF
C775 short_circuit_branch_add gnd! 283.0fF
C776 n_323 gnd! 40.7fF
C777 n_1550 gnd! 40.6fF
C778 pipeUNK18 gnd! 58.3fF
C779 n_771 gnd! 348.2fF
C780 n_959 gnd! 237.1fF
C781 n_671 gnd! 42.4fF
C782 n_1573 gnd! 251.5fF
C783 n_511 gnd! 59.0fF
C784 pipeUNK17 gnd! 56.6fF
C785 n_270 gnd! 731.6fF
C786 n_1426 gnd! 72.2fF
C787 n_513 gnd! 153.4fF
C788 pd6 gnd! 80.3fF
C789 pd2 gnd! 69.0fF
C790 pd7 gnd! 65.8fF
C791 pd1 gnd! 61.1fF
C792 pd0 gnd! 68.9fF
C793 pd5 gnd! 63.4fF
C794 pd3 gnd! 63.4fF
C795 clearIR gnd! 337.7fF
C796 n_380 gnd! 41.3fF
C797 n_1662 gnd! 194.9fF
C798 n_553 gnd! 199.9fF
C799 n_845 gnd! 238.2fF
C800 p2 gnd! 54.2fF
C801 n_31 gnd! 714.2fF
C802 n_24 gnd! 77.0fF
C803 n_1528 gnd! 78.5fF
C804 n_106 gnd! 118.5fF
C805 n_231 gnd! 206.8fF
C806 PD_0xx0xx0x gnd! 276.4fF
C807 PD_n_0xx0xx0x gnd! 165.7fF
C808 n_1515 gnd! 87.0fF
C809 n_1379 gnd! 229.2fF
C810 n_1161 gnd! 78.3fF
C811 n_253 gnd! 304.3fF
C812 n_19 gnd! 103.7fF
C813 n_442 gnd! 207.2fF
C814 n_1619 gnd! 186.0fF
C815 pipeUNK21 gnd! 78.6fF
C816 n_1231 gnd! 123.9fF
C817 n_781 gnd! 613.8fF
C818 n_1154 gnd! 165.9fF
C819 n_1409 gnd! 63.8fF
C820 n_1448 gnd! 101.2fF
C821 n_1330 gnd! 74.6fF
C822 nTWOCYCLE_phi1 gnd! 86.1fF
C823 PD_xxxx10x0 gnd! 368.6fF
C824 pd2_clearIR gnd! 226.2fF
C825 pd3_clearIR gnd! 284.1fF
C826 pd5_clearIR gnd! 283.4fF
C827 PD_1xx000x0 gnd! 370.1fF
C828 n_732 gnd! 284.5fF
C829 n_1124 gnd! 111.5fF
C830 n_2 gnd! 94.7fF
C831 n_1039 gnd! 152.9fF
C832 pipeUNK39 gnd! 57.1fF
C833 n_137 gnd! 25.5fF
C834 n_1718 gnd! 137.9fF
C835 n_770 gnd! 141.4fF
C836 n_812 gnd! 124.5fF
C837 pd4_clearIR gnd! 293.7fF
C838 pd7_clearIR gnd! 230.8fF
C839 pd1_clearIR gnd! 226.6fF
C840 pd0_clearIR gnd! 219.2fF
C841 PD_xxx010x1 gnd! 287.6fF
C842 n_17 gnd! 180.3fF
C843 n_504 gnd! 161.7fF
C844 pipeUNK42 gnd! 96.4fF
C845 nTWOCYCLE gnd! 281.1fF
C846 pipeUNK40 gnd! 57.0fF
C847 n_1380 gnd! 188.2fF
C848 n_14 gnd! 335.6fF
C849 n_666 gnd! 68.1fF
C850 ONEBYTE gnd! 464.8fF
C851 pipenWR_phi2 gnd! 63.9fF
C852 pipeUNK41 gnd! 52.5fF
C853 n_1497 gnd! 137.7fF
C854 n_964 gnd! 174.4fF
C855 n_653 gnd! 53.3fF
C856 pipenT0 gnd! 113.6fF
C857 n_1180 gnd! 143.4fF
C858 n_1533 gnd! 119.0fF
C859 n_664 gnd! 101.9fF
C860 n_889 gnd! 129.0fF
C861 n_390 gnd! 131.9fF
C862 n_1120 gnd! 112.6fF
C863 n_424 gnd! 137.7fF
C864 n_109 gnd! 377.8fF
C865 n_816 gnd! 53.0fF
C866 n_774 gnd! 353.4fF
C867 n_327 gnd! 239.9fF
C868 n_591 gnd! 63.2fF
C869 nop_set_C gnd! 519.2fF
C870 n_191 gnd! 155.2fF
C871 nWR gnd! 374.0fF
C872 n_387 gnd! 81.4fF
C873 n_586 gnd! 380.5fF
C874 n_1517 gnd! 197.3fF
C875 n_853 gnd! 135.7fF
C876 n_206 gnd! 602.7fF
C877 n_559 gnd! 54.6fF
C878 n_608 gnd! 101.1fF
C879 n_1278 gnd! 58.4fF
C880 n_1642 gnd! 470.3fF
C881 n_176 gnd! 235.5fF
C882 n_1655 gnd! 80.9fF
C883 n_1697 gnd! 505.7fF
C884 n_275 gnd! 129.1fF
C885 n_1272 gnd! 71.8fF
C886 n_773 gnd! 140.0fF
C887 n_759 gnd! 51.2fF
C888 n_198 gnd! 204.8fF
C889 pipeUNK37 gnd! 69.7fF
C890 n_944 gnd! 174.5fF
C891 n_218 gnd! 128.5fF
C892 n_470 gnd! 146.8fF
C893 n_1276 gnd! 67.6fF
C894 n_AxBxC_0 gnd! 115.7fF
C895 n_406 gnd! 23.0fF
C896 n_942 gnd! 57.6fF
C897 C01 gnd! 169.0fF
C898 nA_B2 gnd! 303.9fF
C899 n_452 gnd! 39.4fF
C900 alua2 gnd! 114.0fF
C901 n_458 gnd! 127.3fF
C902 idb2 gnd! 935.9fF
C903 alub2 gnd! 157.3fF
C904 s6 gnd! 63.3fF
C905 nots6 gnd! 52.4fF
C906 x7 gnd! 48.4fF
C907 notx7 gnd! 106.8fF
C908 n_871 gnd! 175.8fF
C909 n_1187 gnd! 118.1fF
C910 n_618 gnd! 257.3fF
C911 s5 gnd! 65.6fF
C912 nots5 gnd! 51.1fF
C913 x6 gnd! 48.8fF
C914 notx6 gnd! 109.6fF
C915 sb7 gnd! 819.2fF
C916 y7 gnd! 50.0fF
C917 noty7 gnd! 106.2fF
C918 n_1251 gnd! 184.6fF
C919 abh0 gnd! 180.3fF
C920 nABH0 gnd! 88.4fF
C921 n_1668 gnd! 142.4fF
C922 adh0 gnd! 1179.1fF
C923 n_577 gnd! 11.0fF
C924 nABL7 gnd! 69.2fF
C925 n_1046 gnd! 128.2fF
C926 adl7 gnd! 824.5fF
C927 sb6 gnd! 827.5fF
C928 y6 gnd! 48.0fF
C929 noty6 gnd! 107.1fF
C930 n_1724 gnd! 185.8fF
C931 n_496 gnd! 122.7fF
C932 n_280 gnd! 262.8fF
C933 s4 gnd! 64.6fF
C934 nots4 gnd! 51.3fF
C935 x5 gnd! 51.4fF
C936 notx5 gnd! 106.2fF
C937 n_578 gnd! 187.1fF
C938 n_973 gnd! 123.8fF
C939 n_3 gnd! 262.7fF
C940 s3 gnd! 64.8fF
C941 nots3 gnd! 52.4fF
C942 x4 gnd! 48.2fF
C943 notx4 gnd! 106.7fF
C944 n_436 gnd! 176.1fF
C945 n_34 gnd! 125.4fF
C946 n_998 gnd! 266.2fF
C947 n_A_B_1 gnd! 227.3fF
C948 naluresult1 gnd! 368.3fF
C949 n_1348 gnd! 24.4fF
C950 n_AxB_0 gnd! 168.6fF
C951 A_B0 gnd! 79.0fF
C952 n_105 gnd! 94.8fF
C953 dpc21_ADDADL gnd! 475.8fF
C954 dpc20_ADDSB06 gnd! 422.0fF
C955 n_1033 gnd! 100.3fF
C956 n_75 gnd! 102.8fF
C957 dpc19_ADDSB7 gnd! 407.9fF
C958 nA_B1 gnd! 198.7fF
C959 n_189 gnd! 44.9fF
C960 alua1 gnd! 108.7fF
C961 n_583 gnd! 129.2fF
C962 idb1 gnd! 914.9fF
C963 alub1 gnd! 154.5fF
C964 n_A_B_0 gnd! 316.8fF
C965 naluresult0 gnd! 341.1fF
C966 nA_B0 gnd! 361.3fF
C967 n_316 gnd! 39.4fF
C968 alua0 gnd! 108.4fF
C969 n_624 gnd! 122.0fF
C970 idb0 gnd! 898.8fF
C971 dpc18_nDAA gnd! 506.9fF
C972 n_241 gnd! 147.8fF
C973 n_714 gnd! 89.0fF
C974 n_709 gnd! 101.0fF
C975 n_154 gnd! 138.2fF
C976 n_745 gnd! 52.6fF
C977 n_906 gnd! 182.9fF
C978 n_1499 gnd! 154.0fF
C979 dpc17_SUMS gnd! 449.6fF
C980 n_1305 gnd! 106.0fF
C981 n_1552 gnd! 103.5fF
C982 n_772 gnd! 137.3fF
C983 n_1593 gnd! 151.9fF
C984 n_512 gnd! 57.7fF
C985 n_1333 gnd! 50.5fF
C986 n_1450 gnd! 67.4fF
C987 n_1674 gnd! 64.4fF
C988 n_226 gnd! 65.0fF
C989 n_1705 gnd! 418.3fF
C990 n_930 gnd! 205.6fF
C991 n_1427 gnd! 243.4fF
C992 n_1151 gnd! 50.7fF
C993 n_467 gnd! 197.7fF
C994 n_1286 gnd! 231.9fF
C995 aluvout gnd! 658.3fF
C996 n_1245 gnd! 645.2fF
C997 n_80 gnd! 117.3fF
C998 dpc22_nDSA gnd! 409.6fF
C999 n_674 gnd! 148.1fF
C1000 dpc14_SRS gnd! 461.6fF
C1001 dpc13_ORS gnd! 478.6fF
C1002 dpc16_EORS gnd! 437.0fF
C1003 alub0 gnd! 159.4fF
C1004 s2 gnd! 67.9fF
C1005 nots2 gnd! 54.0fF
C1006 x3 gnd! 51.3fF
C1007 notx3 gnd! 108.2fF
C1008 n_242 gnd! 188.0fF
C1009 n_1190 gnd! 122.0fF
C1010 n_1389 gnd! 261.9fF
C1011 s1 gnd! 68.7fF
C1012 nots1 gnd! 51.5fF
C1013 x2 gnd! 52.6fF
C1014 notx2 gnd! 106.3fF
C1015 n_1694 gnd! 180.2fF
C1016 n_518 gnd! 178.6fF
C1017 abl7 gnd! 233.3fF
C1018 n_1026 gnd! 127.5fF
C1019 n_322 gnd! 603.5fF
C1020 ab6 gnd! 2435.5fF
C1021 n_171 gnd! 582.2fF
C1022 n_524 gnd! 11.0fF
C1023 nABL6 gnd! 70.4fF
C1024 n_1548 gnd! 122.2fF
C1025 adl6 gnd! 854.8fF
C1026 sb5 gnd! 812.5fF
C1027 y5 gnd! 50.0fF
C1028 noty5 gnd! 101.6fF
C1029 n_733 gnd! 178.3fF
C1030 sb4 gnd! 827.2fF
C1031 abl6 gnd! 232.6fF
C1032 n_1195 gnd! 127.5fF
C1033 n_1191 gnd! 528.3fF
C1034 n_1254 gnd! 655.7fF
C1035 n_463 gnd! 10.2fF
C1036 nABL5 gnd! 67.8fF
C1037 n_1094 gnd! 123.3fF
C1038 adl5 gnd! 848.4fF
C1039 y4 gnd! 50.2fF
C1040 noty4 gnd! 106.5fF
C1041 ab5 gnd! 2405.5fF
C1042 abl5 gnd! 233.2fF
C1043 n_172 gnd! 126.5fF
C1044 n_1633 gnd! 538.5fF
C1045 n_210 gnd! 637.6fF
C1046 ab4 gnd! 2383.5fF
C1047 n_738 gnd! 11.0fF
C1048 nABL4 gnd! 68.0fF
C1049 n_1519 gnd! 116.8fF
C1050 adl4 gnd! 866.2fF
C1051 n_658 gnd! 173.6fF
C1052 abl4 gnd! 223.9fF
C1053 n_1676 gnd! 136.0fF
C1054 n_634 gnd! 532.0fF
C1055 n_86 gnd! 621.4fF
C1056 sb3 gnd! 819.2fF
C1057 y3 gnd! 49.4fF
C1058 noty3 gnd! 104.6fF
C1059 n_1531 gnd! 180.2fF
C1060 sb2 gnd! 824.4fF
C1061 n_864 gnd! 11.0fF
C1062 nABL3 gnd! 70.2fF
C1063 n_1507 gnd! 136.7fF
C1064 adl3 gnd! 857.0fF
C1065 y2 gnd! 53.2fF
C1066 noty2 gnd! 106.0fF
C1067 n_1711 gnd! 122.5fF
C1068 n_694 gnd! 260.4fF
C1069 s0 gnd! 67.9fF
C1070 nots0 gnd! 58.7fF
C1071 x1 gnd! 50.8fF
C1072 notx1 gnd! 106.6fF
C1073 n_1709 gnd! 177.0fF
C1074 n_983 gnd! 119.9fF
C1075 n_332 gnd! 266.0fF
C1076 x0 gnd! 50.1fF
C1077 notx0 gnd! 102.1fF
C1078 n_1169 gnd! 181.1fF
C1079 n_1491 gnd! 185.8fF
C1080 sb1 gnd! 817.6fF
C1081 ab3 gnd! 2397.6fF
C1082 abl3 gnd! 224.0fF
C1083 n_990 gnd! 132.2fF
C1084 n_1041 gnd! 541.3fF
C1085 n_138 gnd! 616.0fF
C1086 n_1636 gnd! 12.2fF
C1087 nABL2 gnd! 69.5fF
C1088 n_935 gnd! 114.7fF
C1089 adl2 gnd! 883.8fF
C1090 y1 gnd! 50.7fF
C1091 noty1 gnd! 110.3fF
C1092 n_767 gnd! 185.4fF
C1093 sb0 gnd! 872.6fF
C1094 y0 gnd! 47.3fF
C1095 noty0 gnd! 103.8fF
C1096 abl2 gnd! 230.0fF
C1097 n_951 gnd! 133.3fF
C1098 ab2 gnd! 2427.5fF
C1099 n_1152 gnd! 503.5fF
C1100 n_642 gnd! 572.2fF
C1101 n_416 gnd! 11.3fF
C1102 nABL1 gnd! 66.7fF
C1103 n_1016 gnd! 120.7fF
C1104 adl1 gnd! 886.6fF
C1105 n_564 gnd! 181.9fF
C1106 abl1 gnd! 233.5fF
C1107 n_842 gnd! 129.7fF
C1108 ab1 gnd! 2386.0fF
C1109 n_1479 gnd! 496.4fF
C1110 n_66 gnd! 562.2fF
C1111 n_246 gnd! 12.2fF
C1112 nABL0 gnd! 70.3fF
C1113 n_123 gnd! 125.0fF
C1114 adl0 gnd! 924.1fF
C1115 n_1255 gnd! 104.0fF
C1116 n_108 gnd! 95.3fF
C1117 n_531 gnd! 152.3fF
C1118 dpc15_ANDS gnd! 468.9fF
C1119 dpc10_ADLADD gnd! 689.9fF
C1120 n_1256 gnd! 118.7fF
C1121 dpc11_SBADD gnd! 625.9fF
C1122 n_491 gnd! 95.5fF
C1123 dpc12_0ADD gnd! 544.7fF
C1124 n_1364 gnd! 147.2fF
C1125 n_708 gnd! 98.9fF
C1126 dpc9_DBADD gnd! 585.3fF
C1127 n_956 gnd! 100.5fF
C1128 dpc8_nDBADD gnd! 553.7fF
C1129 n_225 gnd! 102.3fF
C1130 dpc7_SS gnd! 625.0fF
C1131 n_763 gnd! 96.8fF
C1132 dpc6_SBS gnd! 547.7fF
C1133 dpc5_SADL gnd! 464.3fF
C1134 n_95 gnd! 66.4fF
C1135 n_91 gnd! 154.3fF
C1136 n_1541 gnd! 153.1fF
C1137 n_1230 gnd! 153.0fF
C1138 n_71 gnd! 98.2fF
C1139 dpc4_SSB gnd! 557.3fF
C1140 n_282 gnd! 95.4fF
C1141 dpc3_SBX gnd! 568.2fF
C1142 n_196 gnd! 94.4fF
C1143 dpc1_SBY gnd! 527.9fF
C1144 n_593 gnd! 92.2fF
C1145 n_476 gnd! 154.9fF
C1146 n_1223 gnd! 155.1fF
C1147 n_1534 gnd! 157.2fF
C1148 n_35 gnd! 152.7fF
C1149 n_6 gnd! 155.0fF
C1150 n_662 gnd! 95.2fF
C1151 n_543 gnd! 154.1fF
C1152 n_101 gnd! 64.6fF
C1153 n_1529 gnd! 63.7fF
C1154 n_1477 gnd! 41.3fF
C1155 n_360 gnd! 39.6fF
C1156 n_1027 gnd! 39.0fF
C1157 n_441 gnd! 96.3fF
C1158 n_355 gnd! 150.7fF
C1159 n_625 gnd! 154.8fF
C1160 n_692 gnd! 148.9fF
C1161 n_688 gnd! 35.9fF
C1162 n_805 gnd! 38.7fF
C1163 n_931 gnd! 147.8fF
C1164 n_1526 gnd! 145.2fF
C1165 n_968 gnd! 46.8fF
C1166 n_1093 gnd! 150.4fF
C1167 n_1375 gnd! 127.4fF
C1168 notalucin gnd! 320.9fF
C1169 n_415 gnd! 59.7fF
C1170 n_599 gnd! 76.1fF
C1171 dpc28_0ADH0 gnd! 399.6fF
C1172 n_182 gnd! 540.5fF
C1173 n_462 gnd! 320.0fF
C1174 n_1338 gnd! 54.6fF
C1175 n_180 gnd! 151.6fF
C1176 n_1716 gnd! 396.4fF
C1177 n_1211 gnd! 588.0fF
C1178 n_916 gnd! 289.1fF
C1179 n_1708 gnd! 286.9fF
C1180 op_rmw gnd! 78.8fF
C1181 n_1137 gnd! 205.0fF
C1182 pipeUNK36 gnd! 114.5fF
C1183 short_circuit_idx_add gnd! 232.0fF
C1184 n_347 gnd! 535.6fF
C1185 n_1065 gnd! 160.6fF
C1186 n_790 gnd! 279.0fF
C1187 n_368 gnd! 283.7fF
C1188 n_1391 gnd! 535.6fF
C1189 nop_store gnd! 170.1fF
C1190 n_510 gnd! 219.8fF
C1191 n_10 gnd! 359.1fF
C1192 n_1407 gnd! 55.1fF
C1193 n_933 gnd! 163.3fF
C1194 pipedpc28 gnd! 60.5fF
C1195 n_1141 gnd! 140.8fF
C1196 n_1089 gnd! 132.6fF
C1197 n_88 gnd! 45.6fF
C1198 n_982 gnd! 45.5fF
C1199 n_680 gnd! 83.6fF
C1200 n_572 gnd! 326.8fF
C1201 n_261 gnd! 144.1fF
C1202 pipeUNK35 gnd! 43.6fF
C1203 n_720 gnd! 271.6fF
C1204 pipeUNK34 gnd! 49.0fF
C1205 n_238 gnd! 194.9fF
C1206 n_501 gnd! 300.0fF
C1207 n_636 gnd! 117.1fF
C1208 n_726 gnd! 252.4fF
C1209 n_1280 gnd! 46.7fF
C1210 n_1262 gnd! 243.7fF
C1211 n_1679 gnd! 52.7fF
C1212 n_1574 gnd! 53.6fF
C1213 n_796 gnd! 37.6fF
C1214 op_SUMS gnd! 234.4fF
C1215 alucin gnd! 139.3fF
C1216 n_590 gnd! 49.7fF
C1217 n_1215 gnd! 787.6fF
C1218 n_223 gnd! 79.1fF
C1219 n_533 gnd! 170.2fF
C1220 pipeUNK22 gnd! 47.1fF
C1221 pipeUNK23 gnd! 52.9fF
C1222 n_819 gnd! 594.6fF
C1223 pipephi2Reset0 gnd! 48.0fF
C1224 n_29 gnd! 156.2fF
C1225 n_51 gnd! 40.0fF
C1226 n_1688 gnd! 251.6fF
C1227 n_334 gnd! 749.1fF
C1228 n_1508 gnd! 94.0fF
C1229 n_46 gnd! 162.3fF
C1230 n_272 gnd! 696.5fF
C1231 n_239 gnd! 31.8fF
C1232 n_992 gnd! 102.4fF
C1233 n_813 gnd! 156.1fF
C1234 n_25 gnd! 287.9fF
C1235 n_1053 gnd! 57.9fF
C1236 n_1440 gnd! 82.2fF
C1237 Pout3 gnd! 738.6fF
C1238 n_506 gnd! 411.6fF
C1239 n_550 gnd! 162.5fF
C1240 n_885 gnd! 553.6fF
C1241 n_1219 gnd! 85.2fF
C1242 n_1004 gnd! 48.8fF
C1243 n_979 gnd! 89.2fF
C1244 n_1347 gnd! 659.4fF
C1245 n_134 gnd! 421.2fF
C1246 n_1037 gnd! 563.0fF
C1247 n_824 gnd! 551.1fF
C1248 n_1012 gnd! 44.9fF
C1249 n_366 gnd! 140.9fF
C1250 nop_branch_done gnd! 100.4fF
C1251 n_595 gnd! 149.3fF
C1252 n_669 gnd! 105.6fF
C1253 n_1225 gnd! 977.0fF
C1254 n_1412 gnd! 95.9fF
C1255 n_1222 gnd! 127.5fF
C1256 n_384 gnd! 335.3fF
C1257 n_1681 gnd! 34.8fF
C1258 n_905 gnd! 97.0fF
C1259 n_1090 gnd! 477.7fF
C1260 n_1563 gnd! 32.9fF
C1261 n_397 gnd! 111.4fF
C1262 n_11 gnd! 573.5fF
C1263 n_1455 gnd! 664.9fF
C1264 n_928 gnd! 240.0fF
C1265 n_1378 gnd! 15.4fF
C1266 n_605 gnd! 205.3fF
C1267 n_673 gnd! 116.6fF
C1268 n_1304 gnd! 177.9fF
C1269 n_521 gnd! 39.6fF
C1270 n_339 gnd! 46.4fF
C1271 n_621 gnd! 47.0fF
C1272 n_459 gnd! 41.3fF
C1273 n_460 gnd! 41.3fF
C1274 n_795 gnd! 101.2fF
C1275 n_656 gnd! 34.9fF
C1276 n_396 gnd! 92.6fF
C1277 n_1594 gnd! 139.6fF
C1278 D1x1 gnd! 1086.5fF
C1279 n_760 gnd! 63.7fF
C1280 n_236 gnd! 773.2fF
C1281 n_405 gnd! 60.3fF
C1282 n_1343 gnd! 125.0fF
C1283 n_877 gnd! 349.4fF
C1284 n_779 gnd! 379.8fF
C1285 n_1172 gnd! 133.7fF
C1286 BRtaken gnd! 903.6fF
C1287 n_1085 gnd! 272.2fF
C1288 n_1365 gnd! 29.9fF
C1289 n_104 gnd! 956.0fF
C1290 n_1408 gnd! 135.7fF
C1291 n_1044 gnd! 575.1fF
C1292 INTG gnd! 263.2fF
C1293 n_372 gnd! 86.6fF
C1294 op_EORS gnd! 219.3fF
C1295 n_630 gnd! 624.5fF
C1296 n_256 gnd! 801.6fF
C1297 n_847 gnd! 120.1fF
C1298 n_1258 gnd! 649.6fF
C1299 n_1130 gnd! 517.2fF
C1300 n_192 gnd! 427.8fF
C1301 n_1081 gnd! 285.2fF
C1302 pipeUNK32 gnd! 66.5fF
C1303 pipeUNK33 gnd! 54.9fF
C1304 n_152 gnd! 213.1fF
C1305 abl0 gnd! 225.2fF
C1306 n_1660 gnd! 135.3fF
C1307 n_855 gnd! 495.2fF
C1308 ab0 gnd! 2177.4fF
C1309 dpc2_XSB gnd! 562.2fF
C1310 dpc0_YSB gnd! 577.1fF
C1311 n_1100 gnd! 559.6fF
C1312 n_1701 gnd! 256.3fF
C1313 diff_22278_155664# gnd! 74.5fF
C1314 testpad_6 gnd! 182.3fF
C1315 ADL_ABL gnd! 407.0fF
C1316 ADH_ABH gnd! 1259.3fF
C1317 n_602 gnd! 94.9fF
C1318 n_969 gnd! 95.6fF
C1319 n_130 gnd! 96.8fF
C1320 n_1067 gnd! 106.5fF
C1321 n_38 gnd! 116.4fF
C1322 testpad_4 gnd! 121.8fF
C1323 testpad_2 gnd! 880.6fF
C1324 n_1127 gnd! 204.3fF
C1325 testpad_5 gnd! 637.1fF
C1326 testpad_1 gnd! 382.3fF
C1327 n_1247 gnd! 1362.2fF
C1328 n_133 gnd! 150.4fF
C1329 n_1404 gnd! 39.9fF
C1330 n_161 gnd! 145.8fF
C1331 n_220 gnd! 151.7fF
C1332 n_839 gnd! 115.5fF
C1333 n_43 gnd! 1054.7fF
C1334 n_582 gnd! 157.7fF
C1335 n_1113 gnd! 44.4fF
C1336 n_190 gnd! 50.1fF
C1337 n_610 gnd! 54.1fF
C1338 n_0_ADL2 gnd! 285.6fF
C1339 n_0_ADL1 gnd! 281.5fF
C1340 pipeVectorA1 gnd! 56.9fF
C1341 n_1117 gnd! 115.3fF
C1342 n_815 gnd! 135.0fF
C1343 n_952 gnd! 581.9fF
C1344 n_50 gnd! 42.4fF
C1345 pipeUNK31 gnd! 54.3fF
C1346 n_1178 gnd! 370.8fF
C1347 pipeUNK30 gnd! 58.5fF
C1348 n_473 gnd! 268.8fF
C1349 n_1002 gnd! 477.8fF
C1350 n_629 gnd! 293.1fF
C1351 n_646 gnd! 1206.6fF
C1352 n_202 gnd! 106.5fF
C1353 op_ORS gnd! 291.7fF
C1354 n_385 gnd! 120.9fF
C1355 n_782 gnd! 306.0fF
C1356 n_1040 gnd! 123.9fF
C1357 n_1377 gnd! 104.5fF
C1358 nnT2BR gnd! 1138.1fF
C1359 n_1092 gnd! 207.0fF
C1360 n_118 gnd! 259.6fF
C1361 n_480 gnd! 196.2fF
C1362 op_ANDS gnd! 624.6fF
C1363 n_837 gnd! 252.6fF
C1364 n_1145 gnd! 154.7fF
C1365 n_980 gnd! 178.8fF
C1366 n_389 gnd! 219.9fF
C1367 n_1055 gnd! 622.5fF
C1368 n_1560 gnd! 149.2fF
C1369 n_1000 gnd! 133.4fF
C1370 n_300 gnd! 408.3fF
C1371 n_1555 gnd! 34.3fF
C1372 n_1118 gnd! 40.6fF
C1373 n_1649 gnd! 706.8fF
C1374 n_1107 gnd! 236.1fF
C1375 n_440 gnd! 837.0fF
C1376 n_638 gnd! 102.2fF
C1377 n_604 gnd! 703.6fF
C1378 pipeVectorA2 gnd! 47.9fF
C1379 n_70 gnd! 145.1fF
C1380 n_1054 gnd! 112.1fF
C1381 pipeVectorA0 gnd! 79.9fF
C1382 n_911 gnd! 404.3fF
C1383 n_0_ADL0 gnd! 384.4fF
C1384 n_696 gnd! 278.6fF
C1385 n_1361 gnd! 68.3fF ;**FLOATING
C1386 n_79 gnd! 344.2fF
C1387 diff_67022_217892# gnd! 16.2fF ;**FLOATING
C1388 diff_68244_220806# gnd! 9.5fF ;**FLOATING
C1389 diff_67022_220806# gnd! 9.5fF ;**FLOATING
C1390 n_1132 gnd! 50.8fF
C1391 pipephi2Reset0x gnd! 41.4fF
C1392 n_1087 gnd! 160.1fF
C1393 n_717 gnd! 168.2fF
C1394 n_1712 gnd! 286.7fF
C1395 n_1317 gnd! 83.5fF ;**FLOATING
C1396 n_1261 gnd! 31.9fF ;**FLOATING
C1397 n_1207 gnd! 31.9fF ;**FLOATING
C1398 n_728 gnd! 210.4fF
C1399 n_411 gnd! 10.5fF ;**FLOATING
C1400 n_1663 gnd! 98.2fF ;**FLOATING
C1401 diff_77268_238760# gnd! 35.5fF ;**FLOATING
C1402 n_497 gnd! 89.5fF ;**FLOATING
C1403 n_563 gnd! 95.5fF ;**FLOATING
C1404 op_SRS gnd! 1074.5fF
C1405 n_902 gnd! 78.4fF
C1406 n_920 gnd! 95.5fF
C1407 pipeUNK27 gnd! 39.8fF
C1408 n_1598 gnd! 59.5fF
C1409 n_1511 gnd! 98.8fF
C1410 n_785 gnd! 39.6fF
C1411 pipeUNK28 gnd! 46.3fF
C1412 n_1189 gnd! 90.1fF
C1413 n_1624 gnd! 66.3fF
C1414 n_139 gnd! 190.3fF
C1415 n_267 gnd! 630.8fF
C1416 n_383 gnd! 252.8fF
C1417 n_917 gnd! 124.3fF
C1418 n_1058 gnd! 37.8fF
C1419 n_262 gnd! 194.7fF
C1420 pipeUNK29 gnd! 110.0fF
C1421 n_169 gnd! 125.8fF
C1422 n_1175 gnd! 142.7fF
C1423 n_1447 gnd! 63.1fF
C1424 sync gnd! 2500.1fF
C1425 n_417 gnd! 524.8fF
C1426 n_1101 gnd! 770.0fF
C1427 n_132 gnd! 901.1fF
C1428 pipeUNK26 gnd! 41.2fF
C1429 n_317 gnd! 124.2fF
C1430 n_1714 gnd! 207.8fF
C1431 C1x5Reset gnd! 1074.8fF
C1432 n_1289 gnd! 169.0fF
C1433 n_1358 gnd! 452.7fF
C1434 n_632 gnd! 392.6fF
C1435 n_1109 gnd! 461.4fF
C1436 n_544 gnd! 249.5fF
C1437 n_454 gnd! 47.2fF
C1438 n_689 gnd! 218.9fF
C1439 n_1586 gnd! 408.9fF
C1440 n_946 gnd! 442.3fF
C1441 n_734 gnd! 70.5fF
C1442 n_1103 gnd! 32.2fF
C1443 n_445 gnd! 511.7fF
C1444 n_1464 gnd! 275.0fF
C1445 n_616 gnd! 561.8fF
C1446 n_844 gnd! 499.0fF
C1447 n_1351 gnd! 57.1fF
C1448 n_1244 gnd! 101.4fF
C1449 n_1106 gnd! 679.5fF
C1450 n_1604 gnd! 38.1fF
C1451 n_1397 gnd! 38.1fF
C1452 n_698 gnd! 63.6fF
C1453 VEC0 gnd! 596.0fF
C1454 n_508 gnd! 70.8fF
C1455 n_335 gnd! 1011.0fF
C1456 n_1303 gnd! 495.1fF
C1457 n_1717 gnd! 669.7fF
C1458 n_1126 gnd! 45.8fF
C1459 n_1290 gnd! 198.6fF
C1460 n_912 gnd! 51.3fF
C1461 VEC1 gnd! 245.8fF
C1462 n_1452 gnd! 61.2fF
C1463 n_861 gnd! 214.6fF
C1464 brk_done gnd! 1358.8fF
C1465 n_1291 gnd! 56.0fF
C1466 clock2 gnd! 1144.1fF
C1467 n_1312 gnd! 145.4fF
C1468 n_1609 gnd! 92.6fF
C1469 pd6_clearIR gnd! 264.8fF
C1470 n_1309 gnd! 182.8fF
C1471 n_74 gnd! 15.4fF
C1472 clock1 gnd! 1055.8fF
C1473 notir5 gnd! 1269.9fF
C1474 n_1693 gnd! 60.1fF
C1475 nNMIG gnd! 711.3fF
C1476 n_799 gnd! 61.4fF
C1477 n_1675 gnd! 95.4fF
C1478 n_1149 gnd! 63.2fF
C1479 n_1339 gnd! 103.0fF
C1480 nVEC gnd! 634.0fF
C1481 ir5 gnd! 1030.8fF
C1482 n_571 gnd! 244.6fF
C1483 n_343 gnd! 15.4fF
C1484 notir6 gnd! 1042.0fF
C1485 ir6 gnd! 1017.0fF
C1486 notir2 gnd! 1056.2fF
C1487 n_1300 gnd! 96.6fF
C1488 diff_343852_306628# gnd! 52.0fF ;**FLOATING
C1489 n_1083 gnd! 269.2fF
C1490 n_1590 gnd! 16.1fF
C1491 n_597 gnd! 47.8fF
C1492 ir2 gnd! 1023.5fF
C1493 notir3 gnd! 1028.9fF
C1494 n_1620 gnd! 99.4fF
C1495 diff_343852_309072# gnd! 47.1fF ;**FLOATING
C1496 diff_343852_311516# gnd! 44.7fF ;**FLOATING
C1497 ir3 gnd! 1026.4fF
C1498 n_1252 gnd! 68.0fF
C1499 pipenVEC gnd! 62.1fF
C1500 n_1578 gnd! 94.2fF
C1501 n_882 gnd! 160.5fF
C1502 n_562 gnd! 85.1fF
C1503 NMIL gnd! 204.5fF
C1504 n_227 gnd! 284.0fF
C1505 n_703 gnd! 16.1fF
C1506 notir4 gnd! 1056.7fF
C1507 n_927 gnd! 95.7fF
C1508 n_1368 gnd! 344.6fF
C1509 n_862 gnd! 1677.6fF
C1510 pipeT_SYNC gnd! 75.0fF
C1511 n_363 gnd! 111.5fF
C1512 n_1091 gnd! 136.8fF
C1513 n_1360 gnd! 51.3fF
C1514 ir4 gnd! 1022.9fF
C1515 diff_343946_316028# gnd! 141.9fF ;**FLOATING
C1516 diff_348176_321386# gnd! 46.3fF ;**FLOATING
C1517 diff_346014_321386# gnd! 48.8fF ;**FLOATING
C1518 n_1183 gnd! 14.8fF
C1519 n_1605 gnd! 352.0fF
C1520 notir7 gnd! 1050.7fF
C1521 n_541 gnd! 90.8fF
C1522 diff_343852_322514# gnd! 45.3fF ;**FLOATING
C1523 ir7 gnd! 1023.0fF
C1524 notir0 gnd! 996.8fF
C1525 n_409 gnd! 366.4fF
C1526 n_724 gnd! 15.4fF
C1527 n_310 gnd! 93.2fF
C1528 n_1641 gnd! 338.3fF
C1529 n_237 gnd! 14.8fF
C1530 fetch gnd! 677.6fF
C1531 irline3 gnd! 933.9fF
C1532 n_12 gnd! 72.6fF
C1533 n_1575 gnd! 178.3fF
C1534 n_644 gnd! 55.7fF
C1535 _t2 gnd! 926.2fF
C1536 pipeT2out gnd! 121.0fF
C1537 n_1558 gnd! 113.7fF
C1538 n_428 gnd! 155.0fF
C1539 _t3 gnd! 943.6fF
C1540 n_119 gnd! 100.5fF
C1541 n_1133 gnd! 185.0fF
C1542 ir1 gnd! 166.8fF
C1543 n_678 gnd! 240.1fF
C1544 notir1 gnd! 999.4fF
C1545 notRnWprepad gnd! 1134.1fF
C1546 ir0 gnd! 292.6fF
C1547 op_clv gnd! 588.5fF
C1548 op_implied gnd! 337.0fF
C1549 op_T4_mem_abs_idx gnd! 306.5fF
C1550 op_T2_mem_zp gnd! 328.1fF
C1551 nop_branch_bit7 gnd! 734.1fF
C1552 op_T5_mem_ind_idx gnd! 330.1fF
C1553 nop_branch_bit6 gnd! 709.9fF
C1554 x_op_push_pull gnd! 359.1fF
C1555 op_T__asl_rol_a gnd! 380.5fF
C1556 op_T3_mem_abs gnd! 328.0fF
C1557 op_T0_cld_sed gnd! 372.0fF
C1558 op_T__cpx_cpy_imm_zp gnd! 357.2fF
C1559 op_T__cmp gnd! 329.9fF
C1560 op_T__cpx_cpy_abs gnd! 374.5fF
C1561 op_T0_plp gnd! 385.5fF
C1562 x_op_T4_rti gnd! 396.5fF
C1563 x_op_T__adc_sbc gnd! 736.0fF
C1564 x_op_T0_bit gnd! 457.0fF
C1565 op_T0_clc_sec gnd! 427.0fF
C1566 op_T3_mem_zp_idx gnd! 295.9fF
C1567 n_1363 gnd! 195.7fF
C1568 op_T__bit gnd! 603.5fF
C1569 op_asl_rol gnd! 323.3fF
C1570 op_T0_cli_sei gnd! 365.8fF
C1571 x_op_T3_plp_pla gnd! 383.9fF
C1572 op_lsr_ror_dec_inc gnd! 258.4fF
C1573 op_T5_rti_rts gnd! 405.5fF
C1574 op_T2_jmp_abs gnd! 411.7fF
C1575 xx_op_T5_jsr gnd! 424.9fF
C1576 op_T4_jmp gnd! 508.8fF
C1577 op_T2_php gnd! 433.5fF
C1578 n_173 gnd! 188.4fF
C1579 op_T2_php_pha gnd! 410.7fF
C1580 op_store gnd! 299.5fF
C1581 op_T4_brk gnd! 472.6fF
C1582 op_push_pull gnd! 409.5fF
C1583 op_jsr gnd! 415.5fF
C1584 n_9 gnd! 29.0fF
C1585 diff_244212_338400# gnd! 16.3fF
C1586 x_op_jmp gnd! 397.2fF
C1587 op_T3_branch gnd! 382.2fF
C1588 x_op_T4_ind_y gnd! 340.4fF
C1589 op_T3_abs_idx_ind gnd! 290.5fF
C1590 op_brk_rti gnd! 371.9fF
C1591 x_op_T3_abs_idx gnd! 300.7fF
C1592 op_T0_jmp gnd! 428.5fF
C1593 op_T3 gnd! 255.7fF
C1594 op_T5_ind_x gnd! 359.2fF
C1595 op_T0_brk_rti gnd! 402.7fF
C1596 op_T5_rts gnd! 768.4fF
C1597 op_T4 gnd! 241.2fF
C1598 op_T2_ind gnd! 326.0fF
C1599 op_T2_branch gnd! 361.7fF
C1600 op_T2_abs_access gnd! 538.0fF
C1601 n_402 gnd! 58.8fF
C1602 n_400 gnd! 128.4fF
C1603 n_1059 gnd! 121.6fF
C1604 n_834 gnd! 197.6fF
C1605 rw gnd! 2521.9fF
C1606 n_633 gnd! 45.8fF
C1607 n_102 gnd! 549.1fF
C1608 n_1129 gnd! 490.8fF
C1609 n_1467 gnd! 605.6fF
C1610 n_358 gnd! 529.4fF
C1611 n_1399 gnd! 449.2fF
C1612 op_T2_zp_zp_idx gnd! 331.9fF
C1613 op_T3_jsr gnd! 446.0fF
C1614 op_sta_cmp gnd! 422.3fF
C1615 op_shift_right gnd! 321.6fF
C1616 op_T2_brk gnd! 425.7fF
C1617 op_T2_pha gnd! 439.4fF
C1618 op_T0_shift_right_a gnd! 387.3fF
C1619 op_T4_abs_idx gnd! 310.6fF
C1620 op_branch_done gnd! 547.7fF
C1621 op_T5_ind_y gnd! 332.7fF
C1622 op_T0_bit gnd! 384.5fF
C1623 op_T0_and gnd! 310.1fF
C1624 op_T0_shift_a gnd! 439.8fF
C1625 op_T0_tax gnd! 357.5fF
C1626 op_T0_acc gnd! 285.9fF
C1627 op_T0_tay gnd! 359.9fF
C1628 op_T0_pla gnd! 398.4fF
C1629 op_T0_lda gnd! 341.2fF
C1630 op_T__shift_a gnd! 374.2fF
C1631 op_T0_txa gnd! 392.6fF
C1632 op_T__ora_and_eor_adc gnd! 320.1fF
C1633 op_T__adc_sbc gnd! 343.1fF
C1634 op_T2_stack_access gnd! 410.6fF
C1635 op_T0_tya gnd! 418.0fF
C1636 op_shift gnd! 350.6fF
C1637 op_T5_jsr gnd! 541.7fF
C1638 op_rol_ror gnd! 340.1fF
C1639 op_T0_sbc gnd! 522.2fF
C1640 op_T3_jmp gnd! 414.8fF
C1641 op_T0_adc_sbc gnd! 424.7fF
C1642 op_T0_cpx_cpy_inx_iny gnd! 341.9fF
C1643 op_T0_cmp gnd! 328.0fF
C1644 op_rti_rts gnd! 523.0fF
C1645 op_T2_jsr gnd! 543.9fF
C1646 op_T4_ind_x gnd! 401.7fF
C1647 x_op_T3_ind_y gnd! 335.2fF
C1648 op_plp_pla gnd! 360.3fF
C1649 op_inc_nop gnd! 343.9fF
C1650 op_T2_ind_y gnd! 343.6fF
C1651 op_T3_abs_idx gnd! 298.9fF
C1652 op_T3_ind_x gnd! 377.7fF
C1653 op_T4_ind_y gnd! 326.6fF
C1654 op_T4_brk_jsr gnd! 416.5fF
C1655 op_T4_rti gnd! 405.8fF
C1656 op_T2_stack gnd! 505.4fF
C1657 op_T3_stack_bit_jmp gnd! 322.1fF
C1658 op_T2_ADL_ADD gnd! 324.9fF
C1659 op_T0 gnd! 250.9fF
C1660 op_T2_abs gnd! 388.7fF
C1661 op_T0_ora gnd! 391.0fF
C1662 op_T0_eor gnd! 397.5fF
C1663 op_jmp gnd! 434.4fF
C1664 op_ror gnd! 390.8fF
C1665 op_T2 gnd! 452.1fF
C1666 op_T3_plp_pla gnd! 394.6fF
C1667 n_1456 gnd! 92.3fF
C1668 op_T0_php_pha gnd! 393.0fF
C1669 op_T5_rti gnd! 646.1fF
C1670 op_T4_rts gnd! 444.4fF
C1671 op_T0_jsr gnd! 483.9fF
C1672 op_T5_brk gnd! 494.1fF
C1673 op_T0_tay_ldy_not_idx gnd! 331.8fF
C1674 op_T__iny_dey gnd! 376.5fF
C1675 op_T__inx gnd! 399.6fF
C1676 op_T0_ldy_mem gnd! 339.4fF
C1677 op_T0_tsx gnd! 426.2fF
C1678 op_T0_ldx_tax_tsx gnd! 324.4fF
C1679 op_T__dex gnd! 353.7fF
C1680 op_from_x gnd! 472.8fF
C1681 op_T0_txs gnd! 563.7fF
C1682 op_T0_dex gnd! 357.6fF
C1683 op_T2_ind_x gnd! 361.7fF
C1684 op_T0_cpx_inx gnd! 339.9fF
C1685 x_op_T0_txa gnd! 394.0fF
C1686 op_T2_idx_x_xy gnd! 394.0fF
C1687 op_T0_cpy_iny gnd! 335.1fF
C1688 op_xy gnd! 355.3fF
C1689 op_T0_iny_dey gnd! 360.0fF
C1690 x_op_T0_tya gnd! 421.3fF
C1691 op_T3_ind_y gnd! 343.7fF
C1692 op_T2_abs_y gnd! 331.7fF
C1693 n_1606 gnd! 53.1fF
C1694 _t4 gnd! 894.0fF
C1695 op_sty_cpy_mem gnd! 409.1fF
C1696 n_913 gnd! 117.0fF
C1697 n_1699 gnd! 41.1fF
C1698 n_1069 gnd! 930.5fF
C1699 n_1274 gnd! 55.2fF
C1700 n_1024 gnd! 224.4fF
C1701 n_94 gnd! 50.5fF
C1702 n_1650 gnd! 177.6fF
C1703 n_1105 gnd! 665.6fF
C1704 n_1715 gnd! 489.6fF
C1705 n_1696 gnd! 469.7fF
C1706 so gnd! 1148.8fF
C1707 n_127 gnd! 512.0fF
C1708 n_1395 gnd! 84.7fF
C1709 n_742 gnd! 30.5fF
C1710 n_975 gnd! 118.9fF
C1711 n_886 gnd! 30.5fF
C1712 n_995 gnd! 123.4fF
C1713 n_854 gnd! 188.1fF
C1714 n_312 gnd! 187.1fF
C1715 Reset0 gnd! 1529.4fF
C1716 clk2out gnd! 1570.7fF
C1717 n_603 gnd! 310.7fF
C1718 n_47 gnd! 47.9fF
C1719 n_865 gnd! 47.1fF
C1720 n_420 gnd! 130.2fF
C1721 n_1449 gnd! 769.0fF
C1722 n_958 gnd! 249.9fF
C1723 clk0 gnd! 1816.5fF
C1724 res gnd! 970.4fF
C1725 n_519 gnd! 624.5fF
C1726 n_135 gnd! 670.5fF
C1727 n_670 gnd! 579.0fF
C1728 n_747 gnd! 642.6fF
C1729 nIRQP gnd! 592.1fF
C1730 IRQP gnd! 76.0fF
C1731 n_806 gnd! 333.1fF
C1732 n_431 gnd! 73.6fF
C1733 n_330 gnd! 183.1fF
C1734 n_881 gnd! 87.6fF
C1735 n_538 gnd! 100.7fF
C1736 n_807 gnd! 147.4fF
C1737 n_1599 gnd! 195.1fF
C1738 n_346 gnd! 30.5fF
C1739 nNMIP gnd! 122.9fF
C1740 pipeT3out gnd! 110.7fF
C1741 n_1366 gnd! 123.9fF
C1742 n_188 gnd! 263.2fF
C1743 n_1357 gnd! 990.8fF
C1744 n_891 gnd! 53.7fF
C1745 n_284 gnd! 104.4fF
C1746 NMIP gnd! 177.2fF
C1747 _t5 gnd! 1020.8fF
C1748 cclk gnd! 22714.6fF
C1749 n_472 gnd! 140.6fF
C1750 cp1 gnd! 13270.9fF
C1751 n_378 gnd! 190.7fF
C1752 n_18 gnd! 62.7fF
C1753 n_395 gnd! 95.4fF
C1754 pipeT5out gnd! 72.4fF
C1755 n_468 gnd! 128.0fF
C1756 n_16 gnd! 344.0fF
C1757 pipeT4out gnd! 111.4fF
C1758 n_1703 gnd! 152.5fF
C1759 notRdy0 gnd! 2773.1fF
C1760 n_1615 gnd! 128.6fF
C1761 n_645 gnd! 372.8fF
C1762 Vdd gnd! 93485.8fF
C1763 n_1392 gnd! 189.6fF
C1764 clk1out gnd! 1867.9fF
C1765 n_1417 gnd! 750.0fF
C1766 irq gnd! 881.3fF
C1767 rdy gnd! 1015.5fF
C1768 nmi gnd! 913.2fF
