spice-netlist.txt