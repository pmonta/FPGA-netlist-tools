* SPICE3 converted from Lajos's format

M0 N0385 N0770 GND GND efet
M1 GND PC0.11 N0785 GND efet
M2 N0761 N0754 GND GND efet
M3 GND PC2.11 N0821 GND efet
M4 GND R1.0 N0903 GND efet
M5 N0920 R3.0 GND GND efet
M6 GND R5.0 N0929 GND efet
M7 N0947 R7.0 GND GND efet
M8 N0770 N0406 N0785 GND efet
M9 N0770 N0424 N0806 GND efet
M10 N0770 N0434 N0821 GND efet
M11 N0834 N0444 N0770 GND efet
M12 GND R9.0 N0956 GND efet
M13 N0966 R11.0 GND GND efet
M14 GND R13.0 N0975 GND efet
M15 N0984 R15.0 GND GND efet
M16 N0866 N0543 N0903 GND efet
M17 N0866 N0565 N0920 GND efet
M18 N0866 N0581 N0929 GND efet
M19 N0866 N0591 N0947 GND efet
M20 N0866 N0616 N0956 GND efet
M21 N0866 N0632 N0966 GND efet
M22 N0866 N0645 N0975 GND efet
M23 N0866 N0657 N0984 GND efet
M24 N0806 PC1.11 GND GND efet
M25 N0834 PC3.11 GND GND efet
M26 VDD SC(A22+M22)CLK2 N0866 GND efet
M27 VDD (~INH)(X11+X31)CLK1 N0770 GND efet
M28 N0862 WRAB1 N0866 GND efet
M29 D3 RADB1 N0386 GND efet
M30 D3 RADB2 N0385 GND efet
M31 N0770 WADB2 N0761 GND efet
M32 N0754 N0301 GND GND efet
M33 N0753 N0301 N0761 GND efet
M34 N0531 N0866 GND GND efet
M35 GND GND TEST_PAD GND efet
M36 N0497 M12+M22+CLK1~(M11+M12) D0 GND efet
M37 D0 RRAB1 N0531 GND efet
M38 VDD VDD N0531 GND efet
M39 VDD VDD N0754 GND efet
M40 VDD VDD N0385 GND efet
M41 N0385 N0381 PC0.11 GND efet
M42 N0385 N0426 PC2.11 GND efet
M43 VDD VDD N0761 GND efet
M44 PC1.11 N0410 N0385 GND efet
M45 PC3.11 N0439 N0385 GND efet
M46 N0531 N0569 R5.0 GND efet
M47 R11.0 N0619 N0531 GND efet
M48 N0862 N0497 GND GND efet
M49 D0 RRAB0 N0532 GND efet
M50 N0531 N0529 R1.0 GND efet
M51 R3.0 N0544 N0531 GND efet
M52 R7.0 N0583 N0531 GND efet
M53 N0531 N0598 R9.0 GND efet
M54 N0531 N0634 R13.0 GND efet
M55 R15.0 N0647 N0531 GND efet
M56 GND N0289 N0754 GND efet
M57 N0386 N0381 PC0.7 GND efet
M58 PC1.7 N0410 N0386 GND efet
M59 N0386 N0426 PC2.7 GND efet
M60 PC3.7 N0439 N0386 GND efet
M61 VDD VDD N0386 GND efet
M62 N0532 N0529 R0.0 GND efet
M63 R2.0 N0544 N0532 GND efet
M64 N0532 N0569 R4.0 GND efet
M65 R6.0 N0583 N0532 GND efet
M66 N0532 N0598 R8.0 GND efet
M67 N0532 N0619 R10.0 GND efet
M68 N0532 N0634 R12.0 GND efet
M69 N0532 N0647 R14.0 GND efet
M70 VDD VDD N0532 GND efet
M71 GND N0289 N0753 GND efet
M72 N0386 N0774 GND GND efet
M73 GND N0880 N0532 GND efet
M74 N0761 WADB1 N0774 GND efet
M75 N0786 N0406 N0774 GND efet
M76 GND PC0.7 N0786 GND efet
M77 GND PC1.7 N0807 GND efet
M78 N0807 N0424 N0774 GND efet
M79 N0822 N0434 N0774 GND efet
M80 GND PC2.7 N0822 GND efet
M81 GND PC3.7 N0835 GND efet
M82 N0835 N0444 N0774 GND efet
M83 N0904 N0543 N0880 GND efet
M84 GND R0.0 N0904 GND efet
M85 GND R2.0 N0921 GND efet
M86 N0921 N0565 N0880 GND efet
M87 N0930 N0581 N0880 GND efet
M88 GND R6.0 N0948 GND efet
M89 N0880 N0591 N0948 GND efet
M90 GND R8.0 N0957 GND efet
M91 N0311 N0289 GND GND efet
M92 N0880 WRAB0 N0862 GND efet
M93 GND R4.0 N0930 GND efet
M94 N0957 N0616 N0880 GND efet
M95 GND R10.0 N0967 GND efet
M96 N0967 N0632 N0880 GND efet
M97 N0976 N0645 N0880 GND efet
M98 N0976 R12.0 GND GND efet
M99 GND R14.0 N0985 GND efet
M100 N0985 N0657 N0880 GND efet
M101 VDD N0325 N0301 GND efet
M102 VDD (~INH)(X11+X31)CLK1 N0774 GND efet
M103 VDD SC(A22+M22)CLK2 N0880 GND efet
M104 VDD VDD N0862 GND efet
M105 GND GND POC_PAD GND efet
M106 GND PC0.3 N0787 GND efet
M107 GND PC2.3 N0823 GND efet
M108 D3 RADB0 N0387 GND efet
M109 N0808 PC1.3 GND GND efet
M110 N0836 PC3.3 GND GND efet
M111 N0387 N0778 GND GND efet
M112 N0778 N0406 N0787 GND efet
M113 N0778 N0424 N0808 GND efet
M114 N0778 N0434 N0823 GND efet
M115 N0778 N0444 N0836 GND efet
M116 GND R0.1 N0905 GND efet
M117 N0922 R2.1 GND GND efet
M118 GND R4.1 N0931 GND efet
M119 N0949 R6.1 GND GND efet
M120 N0968 R10.1 GND GND efet
M121 N0986 R14.1 GND GND efet
M122 N0881 N0543 N0905 GND efet
M123 N0881 N0565 N0922 GND efet
M124 N0881 N0581 N0931 GND efet
M125 N0881 N0591 N0949 GND efet
M126 N0881 N0616 N0958 GND efet
M127 GND R8.1 N0958 GND efet
M128 N0881 N0632 N0968 GND efet
M129 N0881 N0657 N0986 GND efet
M130 VDD VDD N0863 GND efet
M131 N0881 N0645 N0977 GND efet
M132 GND R12.1 N0977 GND efet
M133 VDD (~INH)(X11+X31)CLK1 N0778 GND efet
M134 VDD SC(A22+M22)CLK2 N0881 GND efet
M135 N0778 WADB0 N0761 GND efet
M136 GND N0498 N0863 GND efet
M137 N0881 WRAB0 N0863 GND efet
M138 N0533 RRAB0 D1 GND efet
M139 D3 M12+M22+CLK1~(M11+M12) N0289 GND efet
M140 N0533 N0881 GND GND efet
M141 D1 RRAB1 N0534 GND efet
M142 VDD VDD N0387 GND efet
M143 VDD VDD N0533 GND efet
M144 N0387 N0381 PC0.3 GND efet
M145 N0387 N0426 PC2.3 GND efet
M146 PC1.3 N0410 N0387 GND efet
M147 PC3.3 N0439 N0387 GND efet
M148 R14.1 N0647 N0533 GND efet
M149 N0533 N0529 R0.1 GND efet
M150 R2.1 N0544 N0533 GND efet
M151 R4.1 N0569 N0533 GND efet
M152 R6.1 N0583 N0533 GND efet
M153 N0533 N0598 R8.1 GND efet
M154 R10.1 N0619 N0533 GND efet
M155 N0533 N0634 R12.1 GND efet
M156 N0388 RADB0 D2 GND efet
M157 N0388 N0381 PC0.2 GND efet
M158 PC1.2 N0410 N0388 GND efet
M159 N0388 N0426 PC2.2 GND efet
M160 PC3.2 N0439 N0388 GND efet
M161 VDD VDD N0388 GND efet
M162 N0534 N0529 R1.1 GND efet
M163 R3.1 N0544 N0534 GND efet
M164 N0534 N0569 R5.1 GND efet
M165 R7.1 N0583 N0534 GND efet
M166 N0534 N0598 R9.1 GND efet
M167 R11.1 N0619 N0534 GND efet
M168 N0534 N0634 R13.1 GND efet
M169 N0534 N0647 R15.1 GND efet
M170 VDD VDD N0534 GND efet
M171 N0388 N0779 GND GND efet
M172 N0290 M12+M22+CLK1~(M11+M12) D2 GND efet
M173 GND N0867 N0534 GND efet
M174 D1 M12+M22+CLK1~(M11+M12) N0498 GND efet
M175 N0779 WADB0 N0762 GND efet
M176 N0788 N0406 N0779 GND efet
M177 GND PC0.2 N0788 GND efet
M178 GND PC1.2 N0809 GND efet
M179 N0809 N0424 N0779 GND efet
M180 N0824 N0434 N0779 GND efet
M181 GND PC2.2 N0824 GND efet
M182 GND PC3.2 N0837 GND efet
M183 N0837 N0444 N0779 GND efet
M184 N0906 N0543 N0867 GND efet
M185 GND R1.1 N0906 GND efet
M186 GND R3.1 N0923 GND efet
M187 N0923 N0565 N0867 GND efet
M188 N0932 N0581 N0867 GND efet
M189 GND R5.1 N0932 GND efet
M190 GND R7.1 N0950 GND efet
M191 N0950 N0591 N0867 GND efet
M192 N0959 N0616 N0867 GND efet
M193 GND R9.1 N0959 GND efet
M194 GND R11.1 N0969 GND efet
M195 N0867 N0632 N0969 GND efet
M196 N0978 N0645 N0867 GND efet
M197 GND R13.1 N0978 GND efet
M198 GND R15.1 N0987 GND efet
M199 N0863 WRAB1 N0867 GND efet
M200 N0987 N0657 N0867 GND efet
M201 N0312 N0290 N0311 GND efet
M202 N0302 N0290 N0301 GND efet
M203 VDD (~INH)(X11+X31)CLK1 N0779 GND efet
M204 N0755 N0290 GND GND efet
M205 VDD SC(A22+M22)CLK2 N0867 GND efet
M206 GND PC0.6 N0789 GND efet
M207 GND PC2.6 N0825 GND efet
M208 N0838 PC3.6 GND GND efet
M209 N0810 PC1.6 GND GND efet
M210 GND R1.2 N0907 GND efet
M211 N0389 N0775 GND GND efet
M212 N0775 N0406 N0789 GND efet
M213 N0775 N0424 N0810 GND efet
M214 N0775 N0434 N0825 GND efet
M215 N0775 N0444 N0838 GND efet
M216 N0924 R3.2 GND GND efet
M217 GND R5.2 N0933 GND efet
M218 N0951 R7.2 GND GND efet
M219 GND R9.2 N0960 GND efet
M220 N0970 R11.2 GND GND efet
M221 N0988 R15.2 GND GND efet
M222 N0868 N0543 N0907 GND efet
M223 N0868 N0565 N0924 GND efet
M224 N0868 N0581 N0933 GND efet
M225 N0868 N0591 N0951 GND efet
M226 N0868 N0616 N0960 GND efet
M227 N0868 N0632 N0970 GND efet
M228 N0868 N0645 N0979 GND efet
M229 N0868 N0657 N0988 GND efet
M230 VDD N0325 N0298 GND efet
M231 N0868 SC(A22+M22)CLK2 VDD GND efet
M232 VDD (~INH)(X11+X31)CLK1 N0775 GND efet
M233 GND R13.2 N0979 GND efet
M234 N0762 WADB1 N0775 GND efet
M235 N0864 WRAB1 N0868 GND efet
M236 N0499 M12+M22+CLK1~(M11+M12) D2 GND efet
M237 GND N0740 SYNC GND efet
M238 N0535 N0868 GND GND efet
M239 N0762 N0298 N0755 GND efet
M240 D2 RRAB1 N0535 GND efet
M241 VDD VDD N0535 GND efet
M242 VDD VDD N0389 GND efet
M243 N0756 N0290 GND GND efet
M244 D2 RADB1 N0389 GND efet
M245 PC0.6 N0381 N0389 GND efet
M246 PC1.6 N0410 N0389 GND efet
M247 N0389 N0426 PC2.6 GND efet
M248 N0390 RADB2 D2 GND efet
M249 PC3.6 N0439 N0389 GND efet
M250 N0535 N0529 R1.2 GND efet
M251 R3.2 N0544 N0535 GND efet
M252 R11.2 N0619 N0535 GND efet
M253 R15.2 N0647 N0535 GND efet
M254 N0864 N0499 GND GND efet
M255 N0536 RRAB0 D2 GND efet
M256 N0535 N0569 R5.2 GND efet
M257 R7.2 N0583 N0535 GND efet
M258 N0535 N0598 R9.2 GND efet
M259 N0535 N0634 R13.2 GND efet
M260 VDD VDD N0756 GND efet
M261 VDD VDD N0762 GND efet
M262 GND N0771 N0390 GND efet
M263 N0390 N0381 PC0.10 GND efet
M264 PC1.10 N0410 N0390 GND efet
M265 N0390 N0426 PC2.10 GND efet
M266 PC3.10 N0439 N0390 GND efet
M267 VDD VDD N0390 GND efet
M268 R0.2 N0529 N0536 GND efet
M269 R2.2 N0544 N0536 GND efet
M270 N0536 N0569 R4.2 GND efet
M271 R6.2 N0583 N0536 GND efet
M272 N0536 N0598 R8.2 GND efet
M273 R10.2 N0619 N0536 GND efet
M274 N0536 N0634 R12.2 GND efet
M275 R14.2 N0647 N0536 GND efet
M276 VDD VDD N0536 GND efet
M277 GND GND CLK2 GND efet
M278 GND N0298 N0756 GND efet
M279 GND N0882 N0536 GND efet
M280 N0790 N0406 N0771 GND efet
M281 GND PC0.10 N0790 GND efet
M282 GND PC1.10 N0811 GND efet
M283 N0811 N0424 N0771 GND efet
M284 N0771 N0434 N0826 GND efet
M285 GND PC2.10 N0826 GND efet
M286 GND PC3.10 N0839 GND efet
M287 N0839 N0444 N0771 GND efet
M288 N0771 WADB2 N0762 GND efet
M289 N0908 N0543 N0882 GND efet
M290 GND R0.2 N0908 GND efet
M291 GND R2.2 N0925 GND efet
M292 N0925 N0565 N0882 GND efet
M293 N0934 N0581 N0882 GND efet
M294 N0934 R4.2 GND GND efet
M295 GND R6.2 N0952 GND efet
M296 N0952 N0591 N0882 GND efet
M297 N0961 N0616 N0882 GND efet
M298 N0961 R8.2 GND GND efet
M299 GND R10.2 N0971 GND efet
M300 N0971 N0632 N0882 GND efet
M301 N0980 N0645 N0882 GND efet
M302 N0980 R12.2 GND GND efet
M303 GND R14.2 N0989 GND efet
M304 N0989 N0657 N0882 GND efet
M305 N0882 WRAB0 N0864 GND efet
M306 GND N0756 N0762 GND efet
M307 VDD (~INH)(X11+X31)CLK1 N0771 GND efet
M308 VDD SC(A22+M22)CLK2 N0882 GND efet
M309 VDD VDD N0864 GND efet
M310 N0391 N0772 GND GND efet
M311 GND PC0.9 N0791 GND efet
M312 GND PC2.9 N0827 GND efet
M313 N0840 PC3.9 GND GND efet
M314 N0812 PC1.9 GND GND efet
M315 GND R0.3 N0909 GND efet
M316 N0763 N0758 GND GND efet
M317 N0772 N0406 N0791 GND efet
M318 N0772 N0424 N0812 GND efet
M319 N0772 N0434 N0827 GND efet
M320 N0772 N0444 N0840 GND efet
M321 N0926 R2.3 GND GND efet
M322 GND R4.3 N0935 GND efet
M323 N0953 R6.3 GND GND efet
M324 GND R8.3 N0962 GND efet
M325 GND R10.3 N0972 GND efet
M326 N0883 N0543 N0909 GND efet
M327 N0883 N0565 N0926 GND efet
M328 N0883 N0581 N0935 GND efet
M329 N0953 N0591 N0883 GND efet
M330 N0883 N0616 N0962 GND efet
M331 N0883 N0632 N0972 GND efet
M332 N0883 N0645 N0981 GND efet
M333 GND R12.3 N0981 GND efet
M334 N0990 R14.3 GND GND efet
M335 N0883 N0657 N0990 GND efet
M336 VDD VDD N0865 GND efet
M337 VDD (~INH)(X11+X31)CLK1 N0772 GND efet
M338 VDD SC(A22+M22)CLK2 N0883 GND efet
M339 N0772 WADB2 N0763 GND efet
M340 GND N0500 N0865 GND efet
M341 N0883 WRAB0 N0865 GND efet
M342 N0758 N0293 GND GND efet
M343 D1 RADB1 N0392 GND efet
M344 D1 RADB2 N0391 GND efet
M345 N0537 RRAB0 D3 GND efet
M346 N0757 N0293 N0763 GND efet
M347 N0537 N0883 GND GND efet
M348 N0538 RRAB1 D3 GND efet
M349 VDD VDD N0758 GND efet
M350 VDD VDD N0763 GND efet
M351 VDD VDD N0391 GND efet
M352 VDD VDD N0537 GND efet
M353 N0391 N0381 PC0.9 GND efet
M354 PC1.9 N0410 N0391 GND efet
M355 N0391 N0426 PC2.9 GND efet
M356 PC3.9 N0439 N0391 GND efet
M357 N0537 N0529 R0.3 GND efet
M358 R2.3 N0544 N0537 GND efet
M359 N0537 N0569 R4.3 GND efet
M360 R6.3 N0583 N0537 GND efet
M361 R10.3 N0619 N0537 GND efet
M362 N0537 N0598 R8.3 GND efet
M363 N0537 N0634 R12.3 GND efet
M364 R14.3 N0647 N0537 GND efet
M365 GND GND CLK1 GND efet
M366 GND N0291 N0758 GND efet
M367 PC1.5 N0410 N0392 GND efet
M368 N0392 N0381 PC0.5 GND efet
M369 N0392 N0426 PC2.5 GND efet
M370 PC3.5 N0439 N0392 GND efet
M371 VDD VDD N0392 GND efet
M372 N0538 N0529 R1.3 GND efet
M373 R3.3 N0544 N0538 GND efet
M374 N0538 N0569 R5.3 GND efet
M375 R7.3 N0583 N0538 GND efet
M376 N0538 N0598 R9.3 GND efet
M377 R11.3 N0619 N0538 GND efet
M378 N0538 N0634 R13.3 GND efet
M379 R15.3 N0647 N0538 GND efet
M380 VDD VDD N0538 GND efet
M381 GND N0291 N0757 GND efet
M382 GND N0776 N0392 GND efet
M383 GND N0869 N0538 GND efet
M384 D3 M12+M22+CLK1~(M11+M12) N0500 GND efet
M385 N0763 WADB1 N0776 GND efet
M386 N0792 N0406 N0776 GND efet
M387 GND PC0.5 N0792 GND efet
M388 GND PC1.5 N0813 GND efet
M389 N0813 N0424 N0776 GND efet
M390 N0828 N0434 N0776 GND efet
M391 N0828 PC2.5 GND GND efet
M392 GND PC3.5 N0841 GND efet
M393 N0841 N0444 N0776 GND efet
M394 N0910 N0543 N0869 GND efet
M395 GND R1.3 N0910 GND efet
M396 GND R3.3 N0927 GND efet
M397 N0927 N0565 N0869 GND efet
M398 N0869 N0581 N0936 GND efet
M399 N0936 R5.3 GND GND efet
M400 GND R7.3 N0954 GND efet
M401 N0954 N0591 N0869 GND efet
M402 N0963 N0616 N0869 GND efet
M403 N0963 R9.3 GND GND efet
M404 GND R11.3 N0973 GND efet
M405 N0869 N0632 N0973 GND efet
M406 N0982 N0645 N0869 GND efet
M407 GND R13.3 N0982 GND efet
M408 GND R15.3 N0991 GND efet
M409 N0869 WRAB1 N0865 GND efet
M410 N0991 N0657 N0869 GND efet
M411 VDD N0325 N0293 GND efet
M412 VDD VDD S00531 GND efet
M413 SYNC N0738 VDD GND efet
M414 N0776 (~INH)(X11+X31)CLK1 VDD GND efet
M415 VDD SC(A22+M22)CLK2 N0869 GND efet
M416 VDD S00531 N0740 GND efet
M417 GND PC0.1 N0793 GND efet
M418 GND PC2.1 N0829 GND efet
M419 N0393 RADB0 D1 GND efet
M420 N0814 PC1.1 GND GND efet
M421 N0842 PC3.1 GND GND efet
M422 N0393 N0780 GND GND efet
M423 N0780 N0406 N0793 GND efet
M424 N0780 N0424 N0814 GND efet
M425 N0780 N0434 N0829 GND efet
M426 N0780 N0444 N0842 GND efet
M427 VDD (~INH)(X11+X31)CLK1 N0780 GND efet
M428 N0780 WADB0 N0763 GND efet
M429 D1 M12+M22+CLK1~(M11+M12) N0291 GND efet
M430 N0299 N0291 N0298 GND efet
M431 VDD S00536 N0738 GND efet
M432 N0461 N0469 GND GND efet
M433 N0313 N0291 N0312 GND efet
M434 N0303 N0291 N0302 GND efet
M435 VDD VDD N0393 GND efet
M436 GND N0461 N0469 GND efet
M437 N0393 N0381 PC0.1 GND efet
M438 PC1.1 N0410 N0393 GND efet
M439 N0393 N0426 PC2.1 GND efet
M440 PC3.1 N0439 N0393 GND efet
M441 N0543 N0902 GND GND efet
M442 N0529 N0902 GND GND efet
M443 N0544 N0919 GND GND efet
M444 N0565 N0919 GND GND efet
M445 VDD VDD N0461 GND efet
M446 N0581 N0928 GND GND efet
M447 N0569 N0928 GND GND efet
M448 N0583 N0938 GND GND efet
M449 N0591 N0938 GND GND efet
M450 N0616 N0955 GND GND efet
M451 N0598 N0955 GND GND efet
M452 N0619 N0965 GND GND efet
M453 N0632 N0965 GND GND efet
M454 N0645 N0974 GND GND efet
M455 N0634 N0974 GND GND efet
M456 N0647 N0983 GND GND efet
M457 N0657 N0983 GND GND efet
M458 VDD VDD N0469 GND efet
M459 VDD VDD S00536 GND efet
M460 N0305 N0292 N0313 GND efet
M461 N0294 N0292 N0303 GND efet
M462 N0294 N0292 N0299 GND efet
M463 N0294 N0292 N0293 GND efet
M464 N0453 N0469 GND GND efet
M465 N0394 RADB0 D0 GND efet
M466 N0394 N0381 PC0.0 GND efet
M467 PC1.0 N0410 N0394 GND efet
M468 N0394 N0426 PC2.0 GND efet
M469 PC3.0 N0439 N0394 GND efet
M470 VDD VDD N0453 GND efet
M471 VDD VDD N0394 GND efet
M472 GND N0781 N0394 GND efet
M473 GND N0461 ADDR-RFSH.1 GND efet
M474 N0292 M12+M22+CLK1~(M11+M12) D0 GND efet
M475 VDD VDD ADDR-RFSH.1 GND efet
M476 (~POC)&CLK2&SC(A32+X12) N0530 N0543 GND efet
M477 CLK2&SC(A12+M12) N0530 N0529 GND efet
M478 CLK2&SC(A12+M12) N0545 N0544 GND efet
M479 (~POC)&CLK2&SC(A32+X12) N0545 N0565 GND efet
M480 (~POC)&CLK2&SC(A32+X12) N0570 N0581 GND efet
M481 CLK2&SC(A12+M12) N0570 N0569 GND efet
M482 CLK2&SC(A12+M12) N0584 N0583 GND efet
M483 (~POC)&CLK2&SC(A32+X12) N0584 N0591 GND efet
M484 (~POC)&CLK2&SC(A32+X12) N0599 N0616 GND efet
M485 CLK2&SC(A12+M12) N0599 N0598 GND efet
M486 CLK2&SC(A12+M12) N0620 N0619 GND efet
M487 (~POC)&CLK2&SC(A32+X12) N0620 N0632 GND efet
M488 (~POC)&CLK2&SC(A32+X12) N0635 N0645 GND efet
M489 CLK2&SC(A12+M12) N0635 N0634 GND efet
M490 CLK2&SC(A12+M12) N0648 N0647 GND efet
M491 (~POC)&CLK2&SC(A32+X12) N0648 N0657 GND efet
M492 N0781 WADB0 N0764 GND efet
M493 N0794 N0406 N0781 GND efet
M494 GND PC0.0 N0794 GND efet
M495 GND PC1.0 N0815 GND efet
M496 GND PC3.0 N0843 GND efet
M497 VDD VDD N0902 GND efet
M498 N0815 N0424 N0781 GND efet
M499 N0781 N0434 N0830 GND efet
M500 N0830 PC2.0 GND GND efet
M501 N0843 N0444 N0781 GND efet
M502 N0759 N0292 GND GND efet
M503 VDD (~INH)(X11+X31)CLK1 N0781 GND efet
M504 VDD VDD N0613 GND efet
M505 N0489 N0455 ADDR-RFSH.1 GND efet
M506 N0454 N0455 N0453 GND efet
M507 N0395 N0777 GND GND efet
M508 GND PC0.4 N0795 GND efet
M509 N0816 PC1.4 GND GND efet
M510 GND PC2.4 N0831 GND efet
M511 N0844 PC3.4 GND GND efet
M512 N0777 N0406 N0795 GND efet
M513 N0777 N0424 N0816 GND efet
M514 N0777 N0434 N0831 GND efet
M515 N0777 N0444 N0844 GND efet
M516 N0305 N0325 VDD GND efet
M517 N0752 N0325 VDD GND efet
M518 VDD (~INH)(X11+X31)CLK1 N0777 GND efet
M519 N0764 WADB1 N0777 GND efet
M520 GND N0489 N0488 GND efet
M521 N0462 N0454 GND GND efet
M522 GND N0530 N0902 GND efet
M523 N0919 N0545 GND GND efet
M524 GND N0570 N0928 GND efet
M525 N0938 N0584 GND GND efet
M526 N0955 N0599 GND GND efet
M527 N0965 N0620 GND GND efet
M528 GND N0635 N0974 GND efet
M529 N0983 N0648 GND GND efet
M530 N0764 N0752 N0759 GND efet
M531 N0488 N0463 N0469 GND efet
M532 N0461 N0463 N0462 GND efet
M533 VDD VDD N0938 GND efet
M534 VDD VDD N0955 GND efet
M535 VDD VDD N0965 GND efet
M536 VDD VDD N0974 GND efet
M537 VDD VDD N0983 GND efet
M538 VDD VDD N0919 GND efet
M539 VDD VDD N0928 GND efet
M540 VDD VDD N0395 GND efet
M541 VDD S00557 RRAB1 GND efet
M542 N0760 N0292 GND GND efet
M543 N0395 N0381 PC0.4 GND efet
M544 PC1.4 N0410 N0395 GND efet
M545 D0 RADB1 N0395 GND efet
M546 N0396 RADB2 D0 GND efet
M547 N0395 N0426 PC2.4 GND efet
M548 PC3.4 N0439 N0395 GND efet
M549 VDD VDD N0760 GND efet
M550 VDD VDD N0764 GND efet
M551 GND N0773 N0396 GND efet
M552 N0396 N0381 PC0.8 GND efet
M553 PC1.8 N0410 N0396 GND efet
M554 N0396 N0426 PC2.8 GND efet
M555 PC3.8 N0439 N0396 GND efet
M556 VDD VDD N0396 GND efet
M557 VDD VDD S00557 GND efet
M558 GND N0752 N0760 GND efet
M559 VDD VDD N0540 GND efet
M560 N0539 N0540 GND GND efet
M561 N0796 N0406 N0773 GND efet
M562 GND PC0.8 N0796 GND efet
M563 GND PC1.8 N0817 GND efet
M564 N0817 N0424 N0773 GND efet
M565 N0832 N0434 N0773 GND efet
M566 N0832 PC2.8 GND GND efet
M567 GND PC3.8 N0845 GND efet
M568 N0845 N0444 N0773 GND efet
M569 N0773 WADB2 N0764 GND efet
M570 N0455 N0463 GND GND efet
M571 GND N0540 N0545 GND efet
M572 GND N0540 N0570 GND efet
M573 GND N0540 N0584 GND efet
M574 GND N0613 N0599 GND efet
M575 GND N0613 N0620 GND efet
M576 GND N0613 N0635 GND efet
M577 GND N0613 N0648 GND efet
M578 GND N0307 N0294 GND efet
M579 N0752 N0307 GND GND efet
M580 GND N0760 N0764 GND efet
M581 GND N0613 N0540 GND efet
M582 VDD (~INH)(X11+X31)CLK1 N0773 GND efet
M583 N0613 N0646 GND GND efet
M584 GND N0455 N0463 GND efet
M585 VDD VDD N0455 GND efet
M586 VDD VDD S00564 GND efet
M587 VDD VDD N0463 GND efet
M588 N0503 N0463 GND GND efet
M589 N0599 N0541 GND GND efet
M590 N0620 N0541 GND GND efet
M591 GND N0541 N0539 GND efet
M592 N0545 N0541 GND GND efet
M593 N0740 N0738 GND GND efet
M594 VDD N0325 N0306 GND efet
M595 VDD VDD N0503 GND efet
M596 GND N0455 ADDR-RFSH.0 GND efet
M597 VDD VDD ADDR-RFSH.0 GND efet
M598 RRAB0 S00564 VDD GND efet
M599 N0306 N0307 N0305 GND efet
M600 GND N0577 N0570 GND efet
M601 GND N0577 N0584 GND efet
M602 N0539 N0542 GND GND efet
M603 GND N0577 N0635 GND efet
M604 GND N0577 N0648 GND efet
M605 VDD VDD N0541 GND efet
M606 N0314 N0306 GND GND efet
M607 VDD VDD WADB2 GND efet
M608 VDD VDD WADB1 GND efet
M609 GND N0577 N0541 GND efet
M610 N0519 CLK1 ADDR-RFSH.0 GND efet
M611 N0504 CLK1 N0503 GND efet
M612 VDD VDD N0314 GND efet
M613 N0406 N0783 GND GND efet
M614 N0381 N0783 GND GND efet
M615 N0410 N0804 GND GND efet
M616 N0424 N0804 GND GND efet
M617 N0434 N0820 GND GND efet
M618 N0426 N0820 GND GND efet
M619 N0439 N0833 GND GND efet
M620 N0444 N0833 GND GND efet
M621 N0570 N0542 GND GND efet
M622 N0599 N0542 GND GND efet
M623 N0635 N0542 GND GND efet
M624 N0738 N0295 GND GND efet
M625 N0577 N0617 GND GND efet
M626 VDD VDD N0577 GND efet
M627 N0518 N0519 GND GND efet
M628 N0508 N0504 GND GND efet
M629 N0712 A32 GND GND efet
M630 N0325 VDD CLK1 GND efet
M631 WADB1 N0318 GND GND efet
M632 GND N0304 WADB2 GND efet
M633 N0314 CLK2 N0315 GND efet
M634 (~POC)CLK2(X12+X32)~INH N0382 N0406 GND efet
M635 ((~SC)(JIN+FIN))CLK1(M11+X21~INH) N0382 N0381 GND efet
M636 ((~SC)(JIN+FIN))CLK1(M11+X21~INH) N0411 N0410 GND efet
M637 (~POC)CLK2(X12+X32)~INH N0411 N0424 GND efet
M638 (~POC)CLK2(X12+X32)~INH N0427 N0434 GND efet
M639 ((~SC)(JIN+FIN))CLK1(M11+X21~INH) N0427 N0426 GND efet
M640 ((~SC)(JIN+FIN))CLK1(M11+X21~INH) N0440 N0439 GND efet
M641 (~POC)CLK2(X12+X32)~INH N0440 N0444 GND efet
M642 N0530 ~(FIN&X12) N0539 GND efet
M643 GND N0560 N0545 GND efet
M644 GND N0560 N0584 GND efet
M645 GND N0560 N0620 GND efet
M646 GND N0560 N0648 GND efet
M647 VDD VDD WADB0 GND efet
M648 N0518 (~INH)&X32&CLK2 N0463 GND efet
M649 N0455 (~INH)&X32&CLK2 N0508 GND efet
M650 VDD N0717 CMROM GND efet
M651 VDD VDD N0561 GND efet
M652 GND ~(FIN&X12) N0561 GND efet
M653 GND A22 N0712 GND efet
M654 GND N0737 CMROM GND efet
M655 GND N0300 WADB0 GND efet
M656 GND N0300 WADB1 GND efet
M657 GND N0300 WADB2 GND efet
M658 N0545 N0561 GND GND efet
M659 N0570 N0561 GND GND efet
M660 N0584 N0561 GND GND efet
M661 N0599 N0561 GND GND efet
M662 N0620 N0561 GND GND efet
M663 N0635 N0561 GND GND efet
M664 N0648 N0561 GND GND efet
M665 VDD VDD N0542 GND efet
M666 N0316 N0315 GND GND efet
M667 VDD VDD N0316 GND efet
M668 WADB0 N0326 GND GND efet
M669 GND N0560 N0542 GND efet
M670 N0711 A12 GND GND efet
M671 VDD VDD N0833 GND efet
M672 N0317 CLK1 N0316 GND efet
M673 VDD VDD N0711 GND efet
M674 GND N0427 N0820 GND efet
M675 N0560 N0582 GND GND efet
M676 GND N0382 N0783 GND efet
M677 N0804 N0411 GND GND efet
M678 N0833 N0440 GND GND efet
M679 VDD VDD N0400 GND efet
M680 VDD VDD N0560 GND efet
M681 N0712 N0732 N0711 GND efet
M682 VDD VDD N0804 GND efet
M683 VDD VDD N0820 GND efet
M684 N0464 N0475 GND GND efet
M685 VDD VDD N0783 GND efet
M686 GND N0409 N0400 GND efet
M687 VDD S00578 N0530 GND efet
M688 VDD S00579 N0545 GND efet
M689 VDD S00580 N0570 GND efet
M690 VDD S00581 N0584 GND efet
M691 VDD S00582 N0599 GND efet
M692 VDD S00583 N0620 GND efet
M693 VDD S00584 N0635 GND efet
M694 VDD S00585 N0648 GND efet
M695 GND N0464 N0475 GND efet
M696 VDD VDD N0464 GND efet
M697 N0732 N0317 GND GND efet
M698 VDD VDD N0732 GND efet
M699 VDD VDD N0475 GND efet
M700 D1 SC&M22&CLK2 N0582 GND efet
M701 RADB1 CLK2 GND GND efet
M702 GND N0384 RADB1 GND efet
M703 GND CLK2 RADB2 GND efet
M704 GND N0374 RADB2 GND efet
M705 N0457 N0475 GND GND efet
M706 GND N0416 RADB0 GND efet
M707 VDD VDD N0457 GND efet
M708 GND N0400 N0427 GND efet
M709 GND N0464 ADDR-PTR.1 GND efet
M710 VDD VDD ADDR-PTR.1 GND efet
M711 D2 SC&M22&CLK2 N0617 GND efet
M712 VDD VDD RADB2 GND efet
M713 N0646 SC&M22&CLK2 D3 GND efet
M714 N0307 N0711 GND GND efet
M715 GND N0409 N0440 GND efet
M716 N0300 CLK2 GND GND efet
M717 VDD VDD N0737 GND efet
M718 VDD VDD N0307 GND efet
M719 VDD VDD N0300 GND efet
M720 VDD VDD S00578 GND efet
M721 VDD VDD S00579 GND efet
M722 VDD VDD S00580 GND efet
M723 VDD VDD S00581 GND efet
M724 VDD VDD S00582 GND efet
M725 VDD VDD S00583 GND efet
M726 VDD VDD S00584 GND efet
M727 VDD VDD S00585 GND efet
M728 N0492 N0459 ADDR-PTR.1 GND efet
M729 N0458 N0459 N0457 GND efet
M730 VDD VDD RADB1 GND efet
M731 GND CLK1 N0307 GND efet
M732 GND N0400 N0382 GND efet
M733 GND N0409 N0411 GND efet
M734 N0491 N0492 GND GND efet
M735 N0465 N0458 GND GND efet
M736 VDD VDD RADB0 GND efet
M737 N0379 CLK2 N0384 GND efet
M738 N0365 CLK2 N0374 GND efet
M739 VDD VDD N0571 GND efet
M740 VDD VDD N0574 GND efet
M741 VDD VDD N0573 GND efet
M742 VDD VDD N0600 GND efet
M743 VDD VDD N0610 GND efet
M744 VDD VDD N0609 GND efet
M745 VDD VDD N0637 GND efet
M746 VDD VDD N0642 GND efet
M747 VDD VDD N0641 GND efet
M748 N0382 N0401 GND GND efet
M749 N0411 N0401 GND GND efet
M750 N0427 N0420 GND GND efet
M751 N0440 N0420 GND GND efet
M752 N0402 CLK2 N0416 GND efet
M753 N0737 N0717 GND GND efet
M754 VDD VDD REG-RFSH.0 GND efet
M755 VDD VDD REG-RFSH.1 GND efet
M756 VDD VDD REG-RFSH.2 GND efet
M757 GND X32 N0402 GND efet
M758 VDD VDD N0402 GND efet
M759 N0475 N0466 N0491 GND efet
M760 N0464 N0466 N0465 GND efet
M761 N0401 N0420 GND GND efet
M762 VDD VDD N0401 GND efet
M763 REG-RFSH.0 SC&A22 N0582 GND efet
M764 REG-RFSH.1 SC&A22 N0617 GND efet
M765 REG-RFSH.2 SC&A22 N0646 GND efet
M766 M12+M22+CLK1~(M11+M12) N0710 VDD GND efet
M767 GND CLK2 RADB0 GND efet
M768 N0459 N0466 GND GND efet
M769 GND N0708 M12+M22+CLK1~(M11+M12) GND efet
M770 VDD S00598 N0382 GND efet
M771 VDD S00599 N0411 GND efet
M772 VDD S00600 N0427 GND efet
M773 GND N0459 N0466 GND efet
M774 VDD S00601 N0440 GND efet
M775 N0409 X12 ADDR-RFSH.1 GND efet
M776 ADDR-PTR.1 X32 N0409 GND efet
M777 N0641 N0600 N0653 GND efet
M778 N0573 CLK1 N0586 GND efet
M779 N0625 N0571 N0609 GND efet
M780 VDD VDD N0466 GND efet
M781 VDD VDD N0459 GND efet
M782 REG-RFSH.0 CLK1 N0566 GND efet
M783 GND N0571 N0573 GND efet
M784 REG-RFSH.1 N0571 N0593 GND efet
M785 GND N0600 N0609 GND efet
M786 N0633 N0600 REG-RFSH.2 GND efet
M787 GND N0637 N0641 GND efet
M788 N0505 N0466 GND GND efet
M789 N0420 X12 ADDR-RFSH.0 GND efet
M790 ADDR-PTR.0 X32 N0420 GND efet
M791 VDD VDD N0505 GND efet
M792 GND N0574 REG-RFSH.0 GND efet
M793 GND N0574 N0571 GND efet
M794 GND N0610 REG-RFSH.1 GND efet
M795 GND N0610 N0600 GND efet
M796 GND N0642 REG-RFSH.2 GND efet
M797 GND N0642 N0637 GND efet
M798 GND N0459 ADDR-PTR.0 GND efet
M799 VDD VDD ADDR-PTR.0 GND efet
M800 N0379 A12 GND GND efet
M801 N0572 SC&A12&CLK2 N0571 GND efet
M802 N0585 SC&A12&CLK2 N0574 GND efet
M803 N0601 N0574 N0600 GND efet
M804 N0624 N0574 N0610 GND efet
M805 N0638 N0610 N0637 GND efet
M806 N0652 N0610 N0642 GND efet
M807 N0710 N0708 GND GND efet
M808 GND N0571 N0574 GND efet
M809 GND N0600 N0610 GND efet
M810 GND N0637 N0642 GND efet
M811 VDD VDD N0379 GND efet
M812 VDD VDD S00609 GND efet
M813 GND N0566 N0572 GND efet
M814 GND N0586 N0585 GND efet
M815 GND N0593 N0601 GND efet
M816 GND N0625 N0624 GND efet
M817 GND N0633 N0638 GND efet
M818 GND N0653 N0652 GND efet
M819 GND A22 N0365 GND efet
M820 VDD VDD S00598 GND efet
M821 VDD VDD S00599 GND efet
M822 VDD VDD S00600 GND efet
M823 VDD VDD S00601 GND efet
M824 VDD VDD N0450 GND efet
M825 N0521 CLK1 ADDR-PTR.0 GND efet
M826 N0506 CLK1 N0505 GND efet
M827 VDD S00609 N0710 GND efet
M828 VDD VDD N0365 GND efet
M829 N0520 N0521 GND GND efet
M830 N0509 N0506 GND GND efet
M831 N0627 N0626 GND GND efet
M832 VDD S00612 N0436 GND efet
M833 N0621 N0622 GND GND efet
M834 CLK2&SC(A12+M12) N0622 GND GND efet
M835 VDD VDD S00628 GND efet
M836 VDD VDD S00612 GND efet
M837 SC(A22+M22)CLK2 N0655 GND GND efet
M838 SC&A12&CLK2 N0649 GND GND efet
M839 (~POC)CLK2(X12+X32)~INH N0449 VDD GND efet
M840 VDD VDD N0708 GND efet
M841 VDD VDD N0437 GND efet
M842 VDD VDD N0494 GND efet
M843 WRAB1 N0578 GND GND efet
M844 (~POC)&CLK2&SC(A32+X12) N0627 GND GND efet
M845 VDD S00620 N0621 GND efet
M846 (~INH)(X11+X31)CLK1 S00628 VDD GND efet
M847 (~INH)(X11+X31)CLK1 N0517 GND GND efet
M848 N0520 CLK2(JMS&DC&M22+BBL(M22+X12+X22)) N0466 GND efet
M849 N0459 CLK2(JMS&DC&M22+BBL(M22+X12+X22)) N0509 GND efet
M850 GND DC RRAB1 GND efet
M851 (~INH)(X11+X31)CLK1 INH GND GND efet
M852 GND N0522 (~INH)(X11+X31)CLK1 GND efet
M853 GND N0592 RRAB1 GND efet
M854 GND M12 N0708 GND efet
M855 N0708 M22 GND GND efet
M856 GND CLK2 RRAB1 GND efet
M857 VDD VDD S00613 GND efet
M858 GND N0450 (~POC)CLK2(X12+X32)~INH GND efet
M859 VDD N0621 CLK2&SC(A12+M12) GND efet
M860 ((~SC)(JIN+FIN))CLK1(M11+X21~INH) N0437 GND GND efet
M861 VDD S00624 SC(A22+M22)CLK2 GND efet
M862 VDD VDD (~INH)&X32&CLK2 GND efet
M863 N0708 CLK1 N0709 GND efet
M864 VDD VDD SC&A12&CLK2 GND efet
M865 GND N0494 (~INH)&X32&CLK2 GND efet
M866 VDD VDD WRAB1 GND efet
M867 N0709 N0278 GND GND efet
M868 VDD VDD N0547 GND efet
M869 VDD VDD N0627 GND efet
M870 VDD N0436 ((~SC)(JIN+FIN))CLK1(M11+X21~INH) GND efet
M871 GND N0436 N0437 GND efet
M872 CLK2(JMS&DC&M22+BBL(M22+X12+X22)) N0467 GND GND efet
M873 VDD S00613 N0449 GND efet
M874 VDD VDD CLK2(JMS&DC&M22+BBL(M22+X12+X22)) GND efet
M875 VDD S00627 N0626 GND efet
M876 VDD VDD N0304 GND efet
M877 VDD N0626 (~POC)&CLK2&SC(A32+X12) GND efet
M878 VDD VDD S00624 GND efet
M879 N0450 N0449 GND GND efet
M880 N0436 N0443 GND GND efet
M881 VDD VDD N0451 GND efet
M882 VDD VDD S00620 GND efet
M883 VDD VDD S00627 GND efet
M884 VDD VDD N0467 GND efet
M885 VDD VDD N0279 GND efet
M886 VDD VDD N0655 GND efet
M887 VDD VDD N0318 GND efet
M888 VDD VDD N0679 GND efet
M889 VDD VDD N0443 GND efet
M890 N0441 N0435 N0436 GND efet
M891 RRAB0 DC GND GND efet
M892 RRAB0 CLK2 GND GND efet
M893 VDD VDD N0460 GND efet
M894 RRAB0 N0615 GND GND efet
M895 VDD VDD N0608 GND efet
M896 GND CLK2 N0496 GND efet
M897 VDD VDD WRAB0 GND efet
M898 VDD VDD N0649 GND efet
M899 N0449 INH GND GND efet
M900 VDD VDD N0522 GND efet
M901 N0496 X32 N0495 GND efet
M902 VDD VDD ~(FIN&X12) GND efet
M903 N0495 ~INH N0494 GND efet
M904 VDD VDD N0511 GND efet
M905 GND JUN+JMS N0309 GND efet
M906 GND JIN+FIN N0441 GND efet
M907 VDD VDD SC&M22&CLK2 GND efet
M908 N0279 CLK2 N0278 GND efet
M909 VDD VDD N0588 GND efet
M910 N0308 X22 N0304 GND efet
M911 N0309 N0310 N0308 GND efet
M912 GND M12 N0323 GND efet
M913 VDD VDD INH GND efet
M914 N0517 CLK2 N0511 GND efet
M915 VDD VDD DC GND efet
M916 GND N0451 N0449 GND efet
M917 VDD VDD SC&A22 GND efet
M918 N0615 CLK2 N0608 GND efet
M919 N0449 POC GND GND efet
M920 GND N0447 N0449 GND efet
M921 GND M12 N0279 GND efet
M922 GND N0438 N0436 GND efet
M923 VDD VDD ~INH GND efet
M924 GND N0679 SC&M22&CLK2 GND efet
M925 GND CLK2 N0451 GND efet
M926 N0656 CLK2 N0655 GND efet
M927 GND A32 N0304 GND efet
M928 N0592 CLK2 N0588 GND efet
M929 GND CLK2 N0460 GND efet
M930 GND CLK1 N0443 GND efet
M931 N0323 JUN+JMS N0324 GND efet
M932 WRAB0 N0547 GND GND efet
M933 N0680 M22 N0679 GND efet
M934 N0650 CLK2 N0649 GND efet
M935 N0279 A32 GND GND efet
M936 GND M22 N0511 GND efet
M937 VDD VDD N0622 GND efet
M938 N0602 X12 N0608 GND efet
M939 N0639 X12 ~(FIN&X12) GND efet
M940 N0654 SC N0656 GND efet
M941 N0320 SC GND GND efet
M942 N0319 JIN+FIN N0320 GND efet
M943 N0318 X22 N0319 GND efet
M944 N0324 N0310 N0318 GND efet
M945 N0321 JCN+ISZ N0323 GND efet
M946 N0318 N0322 N0321 GND efet
M947 N0522 CLK1 GND GND efet
M948 GND M22 N0654 GND efet
M949 N0681 CLK2 N0680 GND efet
M950 GND X12 N0447 GND efet
M951 DC SC GND GND efet
M952 GND N0524 INH GND efet
M953 N0614 ~OPA.0 N0602 GND efet
M954 CLK2(JMS&DC&M22+BBL(M22+X12+X22)) N0460 GND GND efet
M955 N0640 ~OPA.0 N0639 GND efet
M956 N0651 A12 N0650 GND efet
M957 GND M12 N0618 GND efet
M958 N0682 X12 N0683 GND efet
M959 GND INH ~INH GND efet
M960 GND SC N0651 GND efet
M961 N0623 CLK2 N0622 GND efet
M962 GND POC N0626 GND efet
M963 GND SC N0612 GND efet
M964 GND N0643 SC&A22 GND efet
M965 GND SC N0681 GND efet
M966 N0485 JMS GND GND efet
M967 N0484 M22 N0485 GND efet
M968 N0467 DC N0484 GND efet
M969 N0594 N0580 N0588 GND efet
M970 N0595 X12 N0594 GND efet
M971 GND INC+ISZ+ADD+SUB+XCH+LD N0595 GND efet
M972 N0626 N0630 GND GND efet
M973 GND INC+ISZ+ADD+SUB+XCH+LD N0614 GND efet
M974 GND A22 N0318 GND efet
M975 N0589 X22 GND GND efet
M976 N0588 FIN+FIM+SRC+JIN N0589 GND efet
M977 N0597 DC GND GND efet
M978 N0447 X32 GND GND efet
M979 GND X22 N0511 GND efet
M980 N0562 N0564 N0563 GND efet
M981 N0563 M12 GND GND efet
M982 GND M22 N0576 GND efet
M983 N0575 N0564 N0576 GND efet
M984 N0640 N0636 GND GND efet
M985 N0618 A12 GND GND efet
M986 N0618 SC N0623 GND efet
M987 N0683 POC GND GND efet
M988 VDD VDD N0528 GND efet
M989 GND A22 N0654 GND efet
M990 GND ~CN N0322 GND efet
M991 N0596 FIN+FIM+SRC+JIN N0597 GND efet
M992 GND DC N0526 GND efet
M993 N0602 FIN+FIM+SRC+JIN GND GND efet
M994 N0703 CLK2 N0682 GND efet
M995 N0629 X12 GND GND efet
M996 N0322 SC GND GND efet
M997 N0435 SC GND GND efet
M998 VDD VDD N0447 GND efet
M999 GND A32 N0629 GND efet
M1000 N0662 M12 GND GND efet
M1001 N0596 ~OPA.0 N0590 GND efet
M1002 N0428 CLK2 N0438 GND efet
M1003 N0611 X32 N0612 GND efet
M1004 N0562 CLK2 N0547 GND efet
M1005 GND N0590 N0564 GND efet
M1006 N0567 ~OPA.0 N0562 GND efet
M1007 N0631 SC N0629 GND efet
M1008 N0661 SC N0662 GND efet
M1009 N0429 X12 GND GND efet
M1010 GND BBL N0468 GND efet
M1011 N0467 M22 N0468 GND efet
M1012 N0467 X12 N0468 GND efet
M1013 N0428 ~INH N0429 GND efet
M1014 N0631 CLK2 N0630 GND efet
M1015 VDD VDD N0435 GND efet
M1016 GND ~CN N0528 GND efet
M1017 N0467 X22 N0468 GND efet
M1018 N0579 N0568 GND GND efet
M1019 N0525 SC GND GND efet
M1020 GND N0568 N0567 GND efet
M1021 N0575 N0580 N0579 GND efet
M1022 N0578 CLK2 N0575 GND efet
M1023 N0580 ~OPA.0 GND GND efet
M1024 VDD VDD N0578 GND efet
M1025 GND N0603 N0568 GND efet
M1026 N0660 CLK2 N0661 GND efet
M1027 VDD VDD N0428 GND efet
M1028 GND IOR N0683 GND efet
M1029 N0643 A22 N0644 GND efet
M1030 GND SC N0644 GND efet
M1031 N0524 JIN+FIN N0525 GND efet
M1032 GND A32 N0682 GND efet
M1033 GND N0703 L GND efet
M1034 GND N0703 L GND efet
M1035 VDD VDD N0660 GND efet
M1036 N0428 A32 GND GND efet
M1037 N0682 M12 GND GND efet
M1038 VDD VDD N0568 GND efet
M1039 N0333 SC N0326 GND efet
M1040 N0334 JIN+FIN N0333 GND efet
M1041 GND X32 N0334 GND efet
M1042 N0341 JUN+JMS N0326 GND efet
M1043 N0338 JCN+ISZ N0326 GND efet
M1044 N0339 N0322 N0338 GND efet
M1045 GND M22 N0339 GND efet
M1046 VDD VDD N0564 GND efet
M1047 VDD VDD N0590 GND efet
M1048 N0341 N0310 N0339 GND efet
M1049 N0603 INC+ISZ+XCH N0611 GND efet
M1050 VDD VDD N0630 GND efet
M1051 N0527 N0528 N0526 GND efet
M1052 VDD VDD N0322 GND efet
M1053 SC&M12&CLK2 N0660 GND GND efet
M1054 VDD VDD N0643 GND efet
M1055 N0326 A12 GND GND efet
M1056 VDD VDD N0603 GND efet
M1057 N0524 JCN+ISZ N0527 GND efet
M1058 N0524 JUN+JMS N0526 GND efet
M1059 VDD VDD N0580 GND efet
M1060 VDD VDD N0682 GND efet
M1061 VDD VDD SC&M12&CLK2 GND efet
M1062 VDD VDD L GND efet
M1063 VDD VDD N0524 GND efet
M1064 VDD VDD N0326 GND efet
M1065 N0310 SC GND GND efet
M1066 INC/ISZ DC GND GND efet
M1067 OPR.3 N0993 VDD GND efet
M1068 VDD VDD N0310 GND efet
M1069 N1011 SC&M12&CLK2 D0 GND efet
M1070 OPR.2 N0995 VDD GND efet
M1071 GND ~OPR.3 IO GND efet
M1072 GND ~OPR.3 OPE GND efet
M1073 GND ~OPR.3 XCH GND efet
M1074 GND ~OPR.3 BBL GND efet
M1075 GND ~OPR.3 N0628 GND efet
M1076 N0587 ~OPR.3 INC+ISZ+XCH GND efet
M1077 GND ~OPR.3 LD GND efet
M1078 GND ~OPR.3 SUB GND efet
M1079 GND ~OPR.3 ADD GND efet
M1080 GND ~OPR.3 LDM/BBL GND efet
M1081 VDD N0992 ~OPR.3 GND efet
M1082 VDD N0994 ~OPR.2 GND efet
M1083 D2 SC&M12&CLK2 N1009 GND efet
M1084 GND OPR.3 JCN+ISZ GND efet
M1085 JCN OPR.3 GND GND efet
M1086 FIN+FIM OPR.3 GND GND efet
M1087 ISZ OPR.3 GND GND efet
M1088 FIM+SRC OPR.3 GND GND efet
M1089 JIN+FIN OPR.3 GND GND efet
M1090 JUN+JMS OPR.3 GND GND efet
M1091 INC/ISZ OPR.3 GND GND efet
M1092 JMS OPR.3 GND GND efet
M1093 N0636 OPR.3 GND GND efet
M1094 N0628 OPR.3 INC+ISZ+ADD+SUB+XCH+LD GND efet
M1095 GND OPR.3 N0587 GND efet
M1096 FIN+FIM+SRC+JIN OPR.3 GND GND efet
M1097 JUN2+JMS2 OPR.3 GND GND efet
M1098 N0344 S00654 VDD GND efet
M1099 D1 SC&M12&CLK2 N1010 GND efet
M1100 SC N0344 VDD GND efet
M1101 VDD VDD S00654 GND efet
M1102 GND N1008 N0992 GND efet
M1103 N0523 ~OPR.2 GND GND efet
M1104 GND ~OPR.2 ISZ GND efet
M1105 GND ~OPR.2 IO GND efet
M1106 GND ~OPR.2 OPE GND efet
M1107 GND ~OPR.2 JUN+JMS GND efet
M1108 OPR.3 N0992 GND GND efet
M1109 VDD VDD N0361 GND efet
M1110 GND ~OPR.2 INC/ISZ GND efet
M1111 GND ~OPR.2 BBL GND efet
M1112 GND ~OPR.2 JMS GND efet
M1113 INC+ISZ+ADD+SUB+XCH+LD ~OPR.2 N0628 GND efet
M1114 GND ~OPR.2 LDM/BBL GND efet
M1115 GND ~OPR.2 JUN2+JMS2 GND efet
M1116 N0587 ~OPR.2 GND GND efet
M1117 VDD VDD N0998 GND efet
M1118 VDD VDD N0996 GND efet
M1119 D3 SC&M12&CLK2 N1008 GND efet
M1120 VDD VDD N0994 GND efet
M1121 VDD VDD N0992 GND efet
M1122 JCN+ISZ OPR.2 N0523 GND efet
M1123 N0372 JCN+ISZ N0373 GND efet
M1124 GND N0995 ~OPR.2 GND efet
M1125 GND N0993 ~OPR.3 GND efet
M1126 N0998 N1011 GND GND efet
M1127 GND N1009 N0994 GND efet
M1128 GND N1010 N0996 GND efet
M1129 OPR.2 N0994 GND GND efet
M1130 FIN+FIM OPR.2 GND GND efet
M1131 JCN OPR.2 GND GND efet
M1132 FIM+SRC OPR.2 GND GND efet
M1133 GND N0343 N0344 GND efet
M1134 JIN+FIN OPR.2 GND GND efet
M1135 XCH OPR.2 GND GND efet
M1136 N0636 OPR.2 GND GND efet
M1137 N0628 OPR.2 GND GND efet
M1138 INC+ISZ+XCH OPR.2 N0587 GND efet
M1139 FIN+FIM+SRC+JIN OPR.2 GND GND efet
M1140 LD OPR.2 GND GND efet
M1141 SUB OPR.2 GND GND efet
M1142 ADD OPR.2 GND GND efet
M1143 GND N0343 SC GND efet
M1144 N0373 FIN+FIM N0372 GND efet
M1145 GND ~OPR.1 FIN+FIM GND efet
M1146 GND ~OPR.1 ISZ GND efet
M1147 GND ~OPR.1 FIM+SRC GND efet
M1148 GND ~OPR.1 IO GND efet
M1149 GND ~OPR.1 OPE GND efet
M1150 GND ~OPR.1 JIN+FIN GND efet
M1151 GND ~OPR.1 XCH GND efet
M1152 GND ~OPR.1 INC/ISZ GND efet
M1153 INC+ISZ+ADD+SUB+XCH+LD ~OPR.1 N0628 GND efet
M1154 N0587 ~OPR.1 GND GND efet
M1155 N0587 ~OPR.1 INC+ISZ+XCH GND efet
M1156 GND ~OPR.1 FIN+FIM+SRC+JIN GND efet
M1157 GND ~OPR.1 LD GND efet
M1158 N0999 N0998 GND GND efet
M1159 N0995 N0994 GND GND efet
M1160 N0993 N0992 GND GND efet
M1161 ~OPR.1 N0996 VDD GND efet
M1162 N0997 N0996 GND GND efet
M1163 GND ~OPR.1 N0636 GND efet
M1164 N0523 ~OPR.1 GND GND efet
M1165 OPR.0 N0999 VDD GND efet
M1166 JCN OPR.1 GND GND efet
M1167 JUN+JMS OPR.1 GND GND efet
M1168 BBL OPR.1 GND GND efet
M1169 JMS OPR.1 GND GND efet
M1170 SUB OPR.1 GND GND efet
M1171 ADD OPR.1 GND GND efet
M1172 LDM/BBL OPR.1 GND GND efet
M1173 JUN2+JMS2 OPR.1 GND GND efet
M1174 JCN+ISZ OPR.1 N0523 GND efet
M1175 VDD N0998 ~OPR.0 GND efet
M1176 N0361 CLK1 N0343 GND efet
M1177 N0372 X32 GND GND efet
M1178 N0373 JUN+JMS N0372 GND efet
M1179 N0373 SC N0368 GND efet
M1180 GND N0362 N0361 GND efet
M1181 OPR.1 N0997 VDD GND efet
M1182 GND ~OPR.0 ISZ GND efet
M1183 GND ~OPR.0 JCN GND efet
M1184 GND ~OPR.0 OPE GND efet
M1185 GND ~OPR.0 JIN+FIN GND efet
M1186 GND ~OPR.0 XCH GND efet
M1187 GND ~OPR.0 JMS GND efet
M1188 N0587 ~OPR.0 INC+ISZ+XCH GND efet
M1189 GND ~OPR.0 SUB GND efet
M1190 GND ~OPR.0 JCN+ISZ GND efet
M1191 VDD VDD N0352 GND efet
M1192 VDD VDD N0999 GND efet
M1193 VDD VDD N0995 GND efet
M1194 VDD VDD N0997 GND efet
M1195 GND ~OPR.0 N0636 GND efet
M1196 VDD VDD N0368 GND efet
M1197 VDD VDD N0993 GND efet
M1198 FIN+FIM OPA.0 GND GND efet
M1199 FIM+SRC OPR.0 GND GND efet
M1200 IO OPR.0 GND GND efet
M1201 BBL OPR.0 GND GND efet
M1202 LD OPR.0 GND GND efet
M1203 ADD OPR.0 GND GND efet
M1204 N0367 N0352 GND GND efet
M1205 N0368 N0343 N0367 GND efet
M1206 N0368 CLK2 N0362 GND efet
M1207 GND N0998 OPR.0 GND efet
M1208 GND N0997 ~OPR.1 GND efet
M1209 GND X32 N0352 GND efet
M1210 GND N0996 OPR.1 GND efet
M1211 GND N0999 ~OPR.0 GND efet
M1212 VDD VDD FIN+FIM GND efet
M1213 VDD VDD ISZ GND efet
M1214 VDD VDD JCN GND efet
M1215 VDD VDD JUN2+JMS2 GND efet
M1216 VDD VDD JIN+FIN GND efet
M1217 VDD VDD JCN+ISZ GND efet
M1218 VDD VDD INC/ISZ GND efet
M1219 VDD VDD XCH GND efet
M1220 VDD VDD BBL GND efet
M1221 VDD VDD JMS GND efet
M1222 VDD VDD N0636 GND efet
M1223 VDD VDD FIM+SRC GND efet
M1224 VDD VDD IO GND efet
M1225 VDD VDD INC+ISZ+ADD+SUB+XCH+LD GND efet
M1226 VDD VDD ADD GND efet
M1227 VDD VDD LDM/BBL GND efet
M1228 VDD VDD OPE GND efet
M1229 VDD VDD LD GND efet
M1230 VDD VDD JUN+JMS GND efet
M1231 VDD VDD INC+ISZ+XCH GND efet
M1232 VDD VDD SUB GND efet
M1233 VDD VDD FIN+FIM+SRC+JIN GND efet
M1234 VDD VDD N0510 GND efet
M1235 D3 OPA-IB OPA.3 GND efet
M1236 VDD VDD N0493 GND efet
M1237 VDD VDD DCL GND efet
M1238 VDD VDD O-IB GND efet
M1239 VDD VDD KBP GND efet
M1240 VDD VDD STC GND efet
M1241 N0480 ~(X31&~CLK2) GND GND efet
M1242 VDD VDD CLC GND efet
M1243 VDD VDD CLB GND efet
M1244 VDD VDD TCC GND efet
M1245 VDD VDD IOW GND efet
M1246 VDD VDD RAR GND efet
M1247 VDD VDD RAL GND efet
M1248 VDD VDD CMA GND efet
M1249 VDD VDD IAC GND efet
M1250 VDD VDD SBM GND efet
M1251 VDD VDD CMC GND efet
M1252 VDD VDD DAC GND efet
M1253 VDD VDD N0477 GND efet
M1254 VDD VDD TCS GND efet
M1255 VDD VDD DAA GND efet
M1256 VDD VDD N0480 GND efet
M1257 N0482 N0480 N0477 GND efet
M1258 GND OPE N0510 GND efet
M1259 VDD VDD ADM GND efet
M1260 GND IO N0493 GND efet
M1261 VDD VDD IOR GND efet
M1262 VDD VDD N0479 GND efet
M1263 GND OPA.0 N0516 GND efet
M1264 GND N0479 N0482 GND efet
M1265 N0516 FIM+SRC ~SRC GND efet
M1266 ~OPE N0510 VDD GND efet
M1267 D2 OPA-IB OPA.2 GND efet
M1268 GND IO ~I/O GND efet
M1269 ~OPE OPE GND GND efet
M1270 GND IOR N0479 GND efet
M1271 ~I/O N0493 VDD GND efet
M1272 VDD VDD N0769 GND efet
M1273 VDD VDD POC GND efet
M1274 VDD VDD ~CN GND efet
M1275 GND ~I/O IOW GND efet
M1276 GND ~I/O SBM GND efet
M1277 GND ~I/O ADM GND efet
M1278 N0483 A12 N0477 GND efet
M1279 IOR ~I/O GND GND efet
M1280 N0417 SC GND GND efet
M1281 N0476 JCN GND GND efet
M1282 ~OPA.2 N1003 GND GND efet
M1283 GND IOR N0483 GND efet
M1284 ~OPA.3 N1001 GND GND efet
M1285 OPA.2 N1002 GND GND efet
M1286 OPA.3 N1000 GND GND efet
M1287 DCL ~OPE GND GND efet
M1288 O-IB ~OPE GND GND efet
M1289 KBP ~OPE GND GND efet
M1290 TCS ~OPE GND GND efet
M1291 DAA ~OPE GND GND efet
M1292 GND N0397 ~CN GND efet
M1293 N0412 N0397 GND GND efet
M1294 RAR ~OPE GND GND efet
M1295 RAL ~OPE GND GND efet
M1296 CMA ~OPE GND GND efet
M1297 TCC ~OPE GND GND efet
M1298 STC ~OPE GND GND efet
M1299 CMC ~OPE GND GND efet
M1300 DAC ~OPE GND GND efet
M1301 IAC ~OPE GND GND efet
M1302 N0769 A12 GND GND efet
M1303 N0399 X32 GND GND efet
M1304 N0418 X32 N0417 GND efet
M1305 CLC ~OPE GND GND efet
M1306 CLB ~OPE GND GND efet
M1307 GND N0327 N0769 GND efet
M1308 GND N0327 POC GND efet
M1309 N0456 ISZ GND GND efet
M1310 N0327 POC_PAD GND GND efet
M1311 N0478 N0476 GND GND efet
M1312 N0481 N0487 N0478 GND efet
M1313 N0481 ~OPA.3 N0478 GND efet
M1314 GND ~OPA.3 DCL GND efet
M1315 D1 OPA-IB OPA.1 GND efet
M1316 GND ~OPA.3 KBP GND efet
M1317 GND ~OPA.3 TCS GND efet
M1318 GND ~OPA.3 DAA GND efet
M1319 GND ~OPA.3 STC GND efet
M1320 GND CLK2 N0702 GND efet
M1321 GND ~OPA.3 DAC GND efet
M1322 GND ~OPA.3 SBM GND efet
M1323 GND ~OPA.3 ADM GND efet
M1324 GND ~OPA.3 IOR GND efet
M1325 N0413 N0399 N0412 GND efet
M1326 N0413 N0419 N0418 GND efet
M1327 N0419 N0456 N0478 GND efet
M1328 GND N0486 N0481 GND efet
M1329 GND OPA.3 N0481 GND efet
M1330 VDD VDD N0399 GND efet
M1331 VDD VDD N0456 GND efet
M1332 VDD VDD N0413 GND efet
M1333 O-IB OPA.3 GND GND efet
M1334 N0478 ADD_0 N0419 GND efet
M1335 IOW OPA.3 GND GND efet
M1336 RAR OPA.3 GND GND efet
M1337 RAL OPA.3 GND GND efet
M1338 CMA OPA.3 GND GND efet
M1339 TCC OPA.3 GND GND efet
M1340 CMC OPA.3 GND GND efet
M1341 IAC OPA.3 GND GND efet
M1342 CLC OPA.3 GND GND efet
M1343 CLB OPA.3 GND GND efet
M1344 VDD VDD N0476 GND efet
M1345 N0405 CLK2 N0413 GND efet
M1346 VDD VDD S00676 GND efet
M1347 GND N0769 N0327 GND efet
M1348 N0404 CLK1 N0397 GND efet
M1349 N0404 N0405 GND GND efet
M1350 VDD VDD N0671 GND efet
M1351 N0487 N0486 GND GND efet
M1352 VDD N1000 ~OPA.3 GND efet
M1353 VDD VDD N0419 GND efet
M1354 GND ~OPA.2 DCL GND efet
M1355 VDD N1001 OPA.3 GND efet
M1356 N0501 OPA.2 GND GND efet
M1357 GND ~OPA.2 KBP GND efet
M1358 GND ~OPA.2 RAR GND efet
M1359 GND ~OPA.2 RAL GND efet
M1360 GND ~OPA.2 CMA GND efet
M1361 GND ~OPA.2 TCC GND efet
M1362 N0486 ACC_0 N0501 GND efet
M1363 VDD N1002 ~OPA.2 GND efet
M1364 VDD N1003 OPA.2 GND efet
M1365 N0297 CLK2 GND GND efet
M1366 N0702 S00676 VDD GND efet
M1367 VDD VDD N0487 GND efet
M1368 D0 OPA-IB OPA.0 GND efet
M1369 VDD S00678 N0297 GND efet
M1370 N0432 TEST_PAD GND GND efet
M1371 VDD VDD N0327 GND efet
M1372 VDD VDD N0404 GND efet
M1373 TCS OPA.2 GND GND efet
M1374 DAA OPA.2 GND GND efet
M1375 VDD VDD N0486 GND efet
M1376 STC OPA.2 GND GND efet
M1377 CMC OPA.2 GND GND efet
M1378 DAC OPA.2 GND GND efet
M1379 IAC OPA.2 GND GND efet
M1380 CLC OPA.2 GND GND efet
M1381 CLB OPA.2 GND GND efet
M1382 SBM OPA.2 GND GND efet
M1383 ADM OPA.2 GND GND efet
M1384 N0280 CLK2 X22 GND efet
M1385 OPA.1 N1004 GND GND efet
M1386 VDD VDD N0432 GND efet
M1387 ~OPA.1 N1005 GND GND efet
M1388 ~OPA.0 N1007 GND GND efet
M1389 OPA.0 N1006 GND GND efet
M1390 N0688 N0702 N0671 GND efet
M1391 VDD VDD S00678 GND efet
M1392 GND D3 N0671 GND efet
M1393 GND ~OPA.1 DAA GND efet
M1394 VDD VDD ~SRC GND efet
M1395 GND ~OPA.1 RAR GND efet
M1396 GND ~OPA.1 TCC GND efet
M1397 GND ~OPA.1 STC GND efet
M1398 GND ~OPA.1 CMC GND efet
M1399 GND ~OPA.1 IAC GND efet
M1400 GND ~OPA.1 ADM GND efet
M1401 VDD VDD N0398 GND efet
M1402 N0507 CY_1 N0486 GND efet
M1403 N0507 OPA.1 GND GND efet
M1404 VDD VDD N0329 GND efet
M1405 VDD VDD S00685 GND efet
M1406 N0296 N0297 N0295 GND efet
M1407 DCL OPA.1 GND GND efet
M1408 KBP OPA.1 GND GND efet
M1409 TCS OPA.1 GND GND efet
M1410 RAL OPA.1 GND GND efet
M1411 CMA OPA.1 GND GND efet
M1412 GND CLK2 N0398 GND efet
M1413 DAC OPA.1 GND GND efet
M1414 CLC OPA.1 GND GND efet
M1415 CLB OPA.1 GND GND efet
M1416 SBM OPA.1 GND GND efet
M1417 VDD VDD N0784 GND efet
M1418 GND N0280 N0296 GND efet
M1419 VDD N1004 ~OPA.1 GND efet
M1420 VDD N1006 ~OPA.0 GND efet
M1421 N0415 S00685 VDD GND efet
M1422 N0512 N0432 N0486 GND efet
M1423 N0329 ~I/O GND GND efet
M1424 VDD VDD N0799 GND efet
M1425 VDD VDD N0296 GND efet
M1426 N0414 CLK2 A22 GND efet
M1427 GND ~OPA.0 DCL GND efet
M1428 GND ~OPA.0 TCS GND efet
M1429 GND ~OPA.0 DAA GND efet
M1430 GND ~OPA.0 RAL GND efet
M1431 GND ~OPA.0 TCC GND efet
M1432 GND ~OPA.0 CMC GND efet
M1433 GND ~OPA.0 CLC GND efet
M1434 N0739 CLK1 N0296 GND efet
M1435 N0512 OPA.0 GND GND efet
M1436 GND ~OPA.0 ADM GND efet
M1437 VDD VDD S00689 GND efet
M1438 VDD N1005 OPA.1 GND efet
M1439 VDD VDD S00687 GND efet
M1440 VDD N1007 OPA.0 GND efet
M1441 N0407 N0414 GND GND efet
M1442 N0689 S00689 VDD GND efet
M1443 KBP OPA.0 GND GND efet
M1444 RAR OPA.0 GND GND efet
M1445 DAC OPA.0 GND GND efet
M1446 CMA OPA.0 GND GND efet
M1447 STC OPA.0 GND GND efet
M1448 IAC OPA.0 GND GND efet
M1449 CLB OPA.0 GND GND efet
M1450 SBM OPA.0 GND GND efet
M1451 GND N0739 N0741 GND efet
M1452 N0687 S00687 VDD GND efet
M1453 GND ~SRC N0799 GND efet
M1454 N0741 S00690 VDD GND efet
M1455 GND N0782 N0784 GND efet
M1456 N0407 N0398 N0408 GND efet
M1457 GND ~OPE N0415 GND efet
M1458 VDD VDD N0407 GND efet
M1459 VDD VDD S00690 GND efet
M1460 VDD VDD N1001 GND efet
M1461 N0782 N0799 N0798 GND efet
M1462 VDD VDD N1005 GND efet
M1463 VDD VDD N1003 GND efet
M1464 VDD VDD N1007 GND efet
M1465 N0351 N0353 GND GND efet
M1466 N0351 ~(X21&~CLK2) GND GND efet
M1467 GND DCL N0353 GND efet
M1468 WRITE_ACC(1) KBP GND GND efet
M1469 GND TCS WRITE_ACC(1) GND efet
M1470 WRITE_ACC(1) DAA GND GND efet
M1471 GND XCH WRITE_ACC(1) GND efet
M1472 WRITE_ACC(1) POC GND GND efet
M1473 GND CMA WRITE_ACC(1) GND efet
M1474 WRITE_ACC(1) TCC GND GND efet
M1475 GND N0700 N0687 GND efet
M1476 GND DAC WRITE_ACC(1) GND efet
M1477 WRITE_ACC(1) IAC GND GND efet
M1478 WRITE_ACC(1) CLB GND GND efet
M1479 GND LD WRITE_ACC(1) GND efet
M1480 GND SUB WRITE_ACC(1) GND efet
M1481 GND ADD WRITE_ACC(1) GND efet
M1482 GND LDM/BBL WRITE_ACC(1) GND efet
M1483 GND IOR WRITE_ACC(1) GND efet
M1484 GND CLK2 N0375 GND efet
M1485 GND N0408 N0797 GND efet
M1486 X32 N0739 GND GND efet
M1487 GND N0797 N0782 GND efet
M1488 VDD VDD N0797 GND efet
M1489 GND N0700 N0689 GND efet
M1490 ~COM N0782 VDD GND efet
M1491 GND N0784 ~COM GND efet
M1492 N0800 N0801 N0782 GND efet
M1493 GND N0329 N0800 GND efet
M1494 N0798 N0805 GND GND efet
M1495 X32 N0741 VDD GND efet
M1496 VDD VDD N0353 GND efet
M1497 N0415 ~(X21&~CLK2) GND GND efet
M1498 GND SUB WRITE_CARRY(2) GND efet
M1499 WRITE_CARRY(2) POC GND GND efet
M1500 GND TCS WRITE_CARRY(2) GND efet
M1501 WRITE_CARRY(2) TCC GND GND efet
M1502 GND STC WRITE_CARRY(2) GND efet
M1503 WRITE_CARRY(2) CMC GND GND efet
M1504 WRITE_CARRY(2) DAC GND GND efet
M1505 WRITE_CARRY(2) IAC GND GND efet
M1506 GND CLC WRITE_CARRY(2) GND efet
M1507 WRITE_CARRY(2) CLB GND GND efet
M1508 GND SBM WRITE_CARRY(2) GND efet
M1509 GND ADM WRITE_CARRY(2) GND efet
M1510 GND ADD WRITE_CARRY(2) GND efet
M1511 N0442 INC/ISZ GND GND efet
M1512 VDD VDD N0351 GND efet
M1513 N0383 X22 GND GND efet
M1514 D0 N0659 VDD GND efet
M1515 READ_ACC(3) DAA GND GND efet
M1516 GND RAR READ_ACC(3) GND efet
M1517 READ_ACC(3) RAL GND GND efet
M1518 GND IAC READ_ACC(3) GND efet
M1519 GND SUB READ_ACC(3) GND efet
M1520 GND ADD READ_ACC(3) GND efet
M1521 N0380 CLK2 N0383 GND efet
M1522 GND DAC READ_ACC(3) GND efet
M1523 GND SBM READ_ACC(3) GND efet
M1524 GND ADM READ_ACC(3) GND efet
M1525 N1001 N1000 GND GND efet
M1526 N1005 N1004 GND GND efet
M1527 GND N1006 N1007 GND efet
M1528 GND TCS ADD_GROUP(4) GND efet
M1529 GND N1002 N1003 GND efet
M1530 N1000 N1012 GND GND efet
M1531 GND N1014 N1004 GND efet
M1532 GND N1013 N1002 GND efet
M1533 VDD S00699 N0782 GND efet
M1534 VDD VDD N0442 GND efet
M1535 N1006 N1015 GND GND efet
M1536 VDD VDD ~(X31&~CLK2) GND efet
M1537 VDD N0742 X22 GND efet
M1538 N0687 N0688 GND GND efet
M1539 N0375 N0380 GND GND efet
M1540 N0689 N0687 GND GND efet
M1541 GND N0719 X22 GND efet
M1542 GND TCC ADD_GROUP(4) GND efet
M1543 ADD_GROUP(4) ADM GND GND efet
M1544 VDD VDD N0383 GND efet
M1545 GND ADD ADD_GROUP(4) GND efet
M1546 N0448 N0446 GND GND efet
M1547 GND N0375 ~(X31&~CLK2) GND efet
M1548 INC_GROUP(5) INC/ISZ GND GND efet
M1549 D0 SC&M22&CLK2 N1015 GND efet
M1550 VDD N0659 D2 GND efet
M1551 N0448 ~(X21&~CLK2) GND GND efet
M1552 VDD VDD S00699 GND efet
M1553 VDD VDD WRITE_CARRY(2) GND efet
M1554 INC_GROUP(5) IAC GND GND efet
M1555 VDD VDD ~(X21&~CLK2) GND efet
M1556 GND STC INC_GROUP(5) GND efet
M1557 VDD S00709 SUB_GROUP(6) GND efet
M1558 N0658 JUN2+JMS2 GND GND efet
M1559 GND X22 N0288 GND efet
M1560 VDD VDD S00710 GND efet
M1561 VDD VDD N0375 GND efet
M1562 SUB_GROUP(6) SBM GND GND efet
M1563 GND N0689 D3_PAD GND efet
M1564 N0742 N0719 GND GND efet
M1565 VDD VDD N1000 GND efet
M1566 VDD VDD N1004 GND efet
M1567 VDD VDD N1002 GND efet
M1568 VDD VDD N1006 GND efet
M1569 GND CMC SUB_GROUP(6) GND efet
M1570 D3_PAD N0687 VDD GND efet
M1571 VDD VDD N0337 GND efet
M1572 SUB_GROUP(6) SUB GND GND efet
M1573 N1013 SC&M22&CLK2 D2 GND efet
M1574 VDD VDD N0369 GND efet
M1575 VDD VDD N0328 GND efet
M1576 N0742 S00710 VDD GND efet
M1577 ~(X21&~CLK2) N0337 GND GND efet
M1578 VDD VDD INC_GROUP(5) GND efet
M1579 VDD VDD READ_ACC(3) GND efet
M1580 GND LDM/BBL N0658 GND efet
M1581 N1014 SC&M22&CLK2 D1 GND efet
M1582 ACB-IB N0445 N0448 GND efet
M1583 VDD VDD N0658 GND efet
M1584 VDD VDD ADD_GROUP(4) GND efet
M1585 OPA-IB N0658 GND GND efet
M1586 VDD N0659 D1 GND efet
M1587 N0718 CLK1 N0719 GND efet
M1588 ACB-IB ~(X31&~CLK2) N0448 GND efet
M1589 N0337 N0360 GND GND efet
M1590 VDD VDD S00709 GND efet
M1591 D3 SC&M22&CLK2 N1012 GND efet
M1592 N0718 N0281 GND GND efet
M1593 GND CLK2 N0337 GND efet
M1594 N0446 IOW GND GND efet
M1595 N0502 RAL GND GND efet
M1596 VDD VDD N0718 GND efet
M1597 N0445 XCH GND GND efet
M1598 N0328 POC GND GND efet
M1599 VDD S00716 OPA-IB GND efet
M1600 X12 CLK2 N0281 GND efet
M1601 CY-IB N0446 GND GND efet
M1602 VDD N0659 D3 GND efet
M1603 ADSR ~(X31&~CLK2) GND GND efet
M1604 GND N0329 N0328 GND efet
M1605 N0490 RAR GND GND efet
M1606 GND ~(X21&~CLK2) OPA-IB GND efet
M1607 N0515 CMA GND GND efet
M1608 ADSL ~(X31&~CLK2) GND GND efet
M1609 GND N0490 ADSR GND efet
M1610 CY-IB ~(X31&~CLK2) GND GND efet
M1611 VDD VDD S00716 GND efet
M1612 VDD VDD N0659 GND efet
M1613 GND X12 N0288 GND efet
M1614 VDD VDD N0675 GND efet
M1615 N0330 X22 N0331 GND efet
M1616 GND CLK2 N0330 GND efet
M1617 N0335 CLK1 GND GND efet
M1618 N0336 N0337 N0335 GND efet
M1619 N0332 N0328 N0336 GND efet
M1620 N0331 N0329 N0332 GND efet
M1621 N0332 POC N0331 GND efet
M1622 ADSL N0502 GND GND efet
M1623 GND N0675 N0659 GND efet
M1624 ACC-ADAC N0515 GND GND efet
M1625 ACC-ADAC N0342 GND GND efet
M1626 VDD VDD N0445 GND efet
M1627 VDD N0743 X12 GND efet
M1628 N0369 X12 GND GND efet
M1629 VDD VDD CY-IB GND efet
M1630 VDD VDD N0446 GND efet
M1631 GND N0721 X12 GND efet
M1632 GND N0442 ADD-IB GND efet
M1633 VDD VDD ADSR GND efet
M1634 VDD VDD N0502 GND efet
M1635 VDD VDD WRITE_ACC(1) GND efet
M1636 N0360 CLK2 N0369 GND efet
M1637 VDD VDD N0515 GND efet
M1638 N0686 L GND GND efet
M1639 VDD VDD N0678 GND efet
M1640 VDD VDD N0701 GND efet
M1641 VDD VDD ADSL GND efet
M1642 VDD VDD N0490 GND efet
M1643 N0546 INC_GROUP(5) GND GND efet
M1644 N0701 L GND GND efet
M1645 N0342 N0332 VDD GND efet
M1646 VDD VDD N0677 GND efet
M1647 VDD VDD S00725 GND efet
M1648 N0423 CLK2 GND GND efet
M1649 N0685 CLK1 N0701 GND efet
M1650 N0675 CLK1 N0686 GND efet
M1651 GND CLK1 N0678 GND efet
M1652 VDD VDD N0546 GND efet
M1653 ADD-IB ~(X31&~CLK2) GND GND efet
M1654 N0743 N0721 GND GND efet
M1655 N0546 N0342 GND GND efet
M1656 N0743 S00725 VDD GND efet
M1657 GND N0340 N0342 GND efet
M1658 N0678 N0699 GND GND efet
M1659 VDD VDD N0423 GND efet
M1660 GND N0678 N0677 GND efet
M1661 N0699 N0702 N0701 GND efet
M1662 N0684 CLK2 N0675 GND efet
M1663 VDD VDD N0340 GND efet
M1664 GND N0332 N0340 GND efet
M1665 CY-ADAC SUB_GROUP(6) GND GND efet
M1666 CY-ADA ADD_GROUP(4) GND GND efet
M1667 N0707 CLK1 L GND efet
M1668 GND N0685 N0684 GND efet
M1669 GND N0685 N0678 GND efet
M1670 N0720 CLK1 N0721 GND efet
M1671 CY-ADAC N0342 GND GND efet
M1672 N0720 N0282 GND GND efet
M1673 ACC-ADA READ_ACC(3) GND GND efet
M1674 VDD N0677 N0676 GND efet
M1675 VDD VDD N0720 GND efet
M1676 GND N0342 CY-ADA GND efet
M1677 N0676 N0678 GND GND efet
M1678 N0705 N0707 GND GND efet
M1679 VDD S00731 N0332 GND efet
M1680 M22 CLK2 N0282 GND efet
M1681 ADD-ACC WRITE_ACC(1) GND GND efet
M1682 N0513 ADSR CY_1 GND efet
M1683 VDD VDD S00731 GND efet
M1684 ADC-CY WRITE_CARRY(2) GND GND efet
M1685 VDD VDD N0853 GND efet
M1686 ACB-IB S00724 VDD GND efet
M1687 GND N0853 N0854 GND efet
M1688 VDD VDD N0430 GND efet
M1689 GND N0342 ACC-ADA GND efet
M1690 GND N0477 ADD-ACC GND efet
M1691 N0706 L N0705 GND efet
M1692 ADD-IB S00729 VDD GND efet
M1693 GND POC N0705 GND efet
M1694 GND N0477 ADC-CY GND efet
M1695 GND M22 N0288 GND efet
M1696 CY N0415 N0860 GND efet
M1697 VDD VDD ADD-ACC GND efet
M1698 VDD N0744 M22 GND efet
M1699 VDD N0403 N0860 GND efet
M1700 VDD S00732 CY-ADAC GND efet
M1701 VDD VDD N0805 GND efet
M1702 GND N0702 N0706 GND efet
M1703 GND N0723 M22 GND efet
M1704 N0550 CY-ADA N0470 GND efet
M1705 N0470 M12 CY GND efet
M1706 VDD VDD ADC-CY GND efet
M1707 N0425 CLK2 X12 GND efet
M1708 VDD VDD N0421 GND efet
M1709 GND X12 N0853 GND efet
M1710 VDD VDD N0705 GND efet
M1711 N0704 N0705 GND GND efet
M1712 N0513 ADSL CY GND efet
M1713 N0430 N0423 N0431 GND efet
M1714 VDD VDD S00729 GND efet
M1715 VDD VDD S00724 GND efet
M1716 N0421 N0423 N0422 GND efet
M1717 VDD VDD N0470 GND efet
M1718 GND N0855 N0470 GND efet
M1719 VDD VDD S00740 GND efet
M1720 VDD S00734 CY-ADA GND efet
M1721 N0744 N0723 GND GND efet
M1722 VDD VDD N0704 GND efet
M1723 M12 CLK2 N0433 GND efet
M1724 VDD VDD S00734 GND efet
M1725 N0861 ADC-CY CY GND efet
M1726 N0700 N0705 GND GND efet
M1727 N0550 M12 GND GND efet
M1728 N0805 N0422 GND GND efet
M1729 VDD VDD S00732 GND efet
M1730 VDD S00740 N0744 GND efet
M1731 N0855 CY GND GND efet
M1732 N0550 N0546 VDD GND efet
M1733 VDD N0704 N0700 GND efet
M1734 GND SUB_GROUP(6) N0937 GND efet
M1735 CY_1 CY-IB D0 GND efet
M1736 GND N0425 N0421 GND efet
M1737 VDD VDD N0855 GND efet
M1738 GND M12 N0937 GND efet
M1739 GND N0433 N0430 GND efet
M1740 N0846 ADSR CY GND efet
M1741 GND M12 SUB_GROUP(6) GND efet
M1742 N0722 CLK1 N0723 GND efet
M1743 N0855 N0854 N0452 GND efet
M1744 N0550 CY-ADAC N0855 GND efet
M1745 N0722 N0283 GND GND efet
M1746 N0886 N0550 N0894 GND efet
M1747 N0548 N0550 N0549 GND efet
M1748 GND N0452 CY_1 GND efet
M1749 ~TMP.0 N0940 GND GND efet
M1750 VDD VDD N0801 GND efet
M1751 VDD VDD N0722 GND efet
M1752 GND N0431 N0801 GND efet
M1753 GND N0878 N0846 GND efet
M1754 N0886 N0887 N0878 GND efet
M1755 N0846 N0874 VDD GND efet
M1756 N0894 N0870 GND GND efet
M1757 N0548 N0870 GND GND efet
M1758 N0549 N0887 GND GND efet
M1759 VDD N0939 ~TMP.0 GND efet
M1760 N0283 CLK2 M12 GND efet
M1761 VDD VDD CY_1 GND efet
M1762 N0870 ACC-ADAC N0856 GND efet
M1763 N0887 N0937 ~TMP.0 GND efet
M1764 N0346 N0849 GND GND efet
M1765 N0856 N0854 N0849 GND efet
M1766 VDD VDD N0350 GND efet
M1767 VDD VDD N0911 GND efet
M1768 GND N0939 N0940 GND efet
M1769 VDD VDD N0346 GND efet
M1770 N0549 N0870 N0911 GND efet
M1771 VDD VDD N0940 GND efet
M1772 CY_1 ADSL ACC.0 GND efet
M1773 N0911 N0887 N0548 GND efet
M1774 GND N0803 N0403 GND efet
M1775 N0403 N0802 GND GND efet
M1776 VDD VDD N0856 GND efet
M1777 N0874 N0878 GND GND efet
M1778 GND M12 N0288 GND efet
M1779 N0818 N0803 GND GND efet
M1780 N0378 DAA N0818 GND efet
M1781 N0378 O-IB GND GND efet
M1782 GND M12 N0870 GND efet
M1783 GND ACC.0 N0856 GND efet
M1784 N0604 M12 VDD GND efet
M1785 GND N0346 ACC_0 GND efet
M1786 TMP.0 N0940 VDD GND efet
M1787 GND N0939 TMP.0 GND efet
M1788 GND N0870 N0898 GND efet
M1789 N0898 N0550 GND GND efet
M1790 GND N0887 N0898 GND efet
M1791 N0350 KBP GND GND efet
M1792 VDD N0745 M12 GND efet
M1793 N0803 CY_1 GND GND efet
M1794 N0802 DAA GND GND efet
M1795 VDD VDD N0471 GND efet
M1796 GND POC N0717 GND efet
M1797 GND N0725 M12 GND efet
M1798 VDD VDD N0874 GND efet
M1799 N0846 ADD-ACC ACC.0 GND efet
M1800 N0915 N0911 GND GND efet
M1801 TMP.0 SUB_GROUP(6) N0887 GND efet
M1802 N0898 N0553 N0878 GND efet
M1803 VDD VDD N0915 GND efet
M1804 D0 N0964 N0604 GND efet
M1805 N0717 S00757 VDD GND efet
M1806 VDD VDD N0802 GND efet
M1807 N0819 N0356 N0803 GND efet
M1808 N0471 M12 ACC.0 GND efet
M1809 N0471 N0856 GND GND efet
M1810 D0 ACB-IB N0346 GND efet
M1811 N0847 ADSR ACC.0 GND efet
M1812 GND N0604 N0939 GND efet
M1813 VDD VDD N0803 GND efet
M1814 GND N0846 ADD_0 GND efet
M1815 VDD VDD N0378 GND efet
M1816 N0553 N0915 GND GND efet
M1817 VDD VDD N0878 GND efet
M1818 N0717 ~COM GND GND efet
M1819 VDD VDD S00761 GND efet
M1820 VDD VDD S00757 GND efet
M1821 N0939 S00762 VDD GND efet
M1822 VDD VDD ACC_0 GND efet
M1823 N0870 ACC-ADA N0471 GND efet
M1824 N0745 N0725 GND GND efet
M1825 GND POC D2_PAD GND efet
M1826 VDD VDD N0403 GND efet
M1827 VDD N0911 N0553 GND efet
M1828 N0672 D2 GND GND efet
M1829 VDD VDD S00766 GND efet
M1830 N0846 ADD-IB D0 GND efet
M1831 VDD S00761 N0745 GND efet
M1832 GND N0348 N0819 GND efet
M1833 N0819 N0347 GND GND efet
M1834 GND N0884 N0847 GND efet
M1835 VDD S00764 ACC-ADAC GND efet
M1836 VDD VDD S00767 GND efet
M1837 VDD VDD N0672 GND efet
M1838 VDD VDD S00765 GND efet
M1839 VDD VDD S00762 GND efet
M1840 GND N0342 N0964 GND efet
M1841 N0692 S00766 VDD GND efet
M1842 N0888 N0553 N0895 GND efet
M1843 N0552 N0553 N0551 GND efet
M1844 VDD VDD S00764 GND efet
M1845 N0888 N0889 N0875 GND efet
M1846 GND N0871 N0895 GND efet
M1847 N0551 N0871 GND GND efet
M1848 N0552 N0889 GND GND efet
M1849 N0690 S00765 VDD GND efet
M1850 N0724 CLK1 N0725 GND efet
M1851 VDD VDD ADD_0 GND efet
M1852 VDD VDD N0766 GND efet
M1853 VDD VDD N0751 GND efet
M1854 VDD VDD DCL.0 GND efet
M1855 VDD VDD N0964 GND efet
M1856 VDD VDD N0354 GND efet
M1857 VDD VDD N0363 GND efet
M1858 VDD VDD N0370 GND efet
M1859 N0724 N0284 GND GND efet
M1860 VDD VDD N0345 GND efet
M1861 N0377 N0378 N0376 GND efet
M1862 ~TMP.1 N0942 GND GND efet
M1863 N0847 N0875 VDD GND efet
M1864 VDD VDD N0724 GND efet
M1865 VDD N0941 ~TMP.1 GND efet
M1866 ADD_0 N0847 GND GND efet
M1867 D1 ADD-IB N0847 GND efet
M1868 N0284 CLK2 A32 GND efet
M1869 TMP.1 N0937 N0889 GND efet
M1870 N0691 N0702 N0672 GND efet
M1871 N0912 S00767 VDD GND efet
M1872 N0871 ACC-ADAC N0472 GND efet
M1873 N0552 N0871 N0912 GND efet
M1874 GND N0700 N0690 GND efet
M1875 N0912 N0889 N0551 GND efet
M1876 VDD VDD N0942 GND efet
M1877 GND N0700 N0692 GND efet
M1878 GND N0941 N0942 GND efet
M1879 GND A32 N0288 GND efet
M1880 VDD VDD N0377 GND efet
M1881 GND N0875 N0884 GND efet
M1882 N0347 ACB-IB D1 GND efet
M1883 N0846 ADSL ACC.1 GND efet
M1884 VDD VDD N0472 GND efet
M1885 ACC.1 M12 N0472 GND efet
M1886 GND N0857 N0472 GND efet
M1887 VDD N0746 A32 GND efet
M1888 GND N0871 N0899 GND efet
M1889 N0899 N0553 GND GND efet
M1890 GND N0889 N0899 GND efet
M1891 GND N0727 A32 GND efet
M1892 N0376 N0350 GND GND efet
M1893 VDD VDD N0371 GND efet
M1894 GND N0347 ACC_0 GND efet
M1895 N0916 N0912 GND GND efet
M1896 N0605 M12 VDD GND efet
M1897 N0899 N0556 N0875 GND efet
M1898 TMP.1 N0942 VDD GND efet
M1899 GND N0941 TMP.1 GND efet
M1900 VDD VDD N0916 GND efet
M1901 VDD VDD N0884 GND efet
M1902 VDD M12 N0871 GND efet
M1903 N0751 DCL.0 GND GND efet
M1904 DCL.0 POC GND GND efet
M1905 N0857 ACC.1 GND GND efet
M1906 N0847 ADD-ACC ACC.1 GND efet
M1907 DCL.0 N0767 GND GND efet
M1908 ~TMP.1 SUB_GROUP(6) N0889 GND efet
M1909 D1 N0964 N0605 GND efet
M1910 GND N0350 N0345 GND efet
M1911 GND N0350 N0354 GND efet
M1912 N0363 N0350 GND GND efet
M1913 N0370 N0350 GND GND efet
M1914 N0556 N0916 GND GND efet
M1915 N0766 N0351 GND GND efet
M1916 VDD VDD N0875 GND efet
M1917 GND DCL.0 N0716 GND efet
M1918 VDD VDD N0857 GND efet
M1919 VDD VDD S00778 GND efet
M1920 N0848 ADSR ACC.1 GND efet
M1921 N0746 N0727 GND GND efet
M1922 N0941 N0605 GND GND efet
M1923 N0690 N0691 GND GND efet
M1924 N0767 N0766 N0751 GND efet
M1925 N0692 N0690 GND GND efet
M1926 VDD VDD N0347 GND efet
M1927 VDD N0912 N0556 GND efet
M1928 VDD VDD N0364 GND efet
M1929 N0871 ACC-ADA N0857 GND efet
M1930 N0746 S00778 VDD GND efet
M1931 GND N0850 N0347 GND efet
M1932 N0857 N0854 N0850 GND efet
M1933 N0941 S00781 VDD GND efet
M1934 GND N0371 N0370 GND efet
M1935 GND N0879 N0848 GND efet
M1936 D2 N0964 N0606 GND efet
M1937 GND N0346 N0371 GND efet
M1938 N0767 N0351 N0371 GND efet
M1939 N0896 N0556 N0890 GND efet
M1940 N0555 N0556 N0554 GND efet
M1941 N0872 ACC-ADAC N0858 GND efet
M1942 N0848 N0876 VDD GND efet
M1943 GND N0692 D2_PAD GND efet
M1944 N0348 N0851 GND GND efet
M1945 N0345 N0346 GND GND efet
M1946 N0354 N0346 GND GND efet
M1947 N0363 N0346 GND GND efet
M1948 N0376 N0346 GND GND efet
M1949 N0858 N0854 N0851 GND efet
M1950 N0890 N0891 N0879 GND efet
M1951 GND N0872 N0896 GND efet
M1952 N0554 N0872 GND GND efet
M1953 N0555 N0891 GND GND efet
M1954 VDD VDD S00781 GND efet
M1955 N0726 CLK1 N0727 GND efet
M1956 D2_PAD N0690 VDD GND efet
M1957 VDD VDD N0348 GND efet
M1958 N0726 N0285 GND GND efet
M1959 GND DCL.1 N0716 GND efet
M1960 VDD VDD N0726 GND efet
M1961 N0847 ADSL ACC.2 GND efet
M1962 VDD VDD N0858 GND efet
M1963 N0665 N0676 GND GND efet
M1964 N0285 CLK2 A22 GND efet
M1965 ~TMP.2 N0944 GND GND efet
M1966 DCL.1 N0765 GND GND efet
M1967 VDD VDD N0913 GND efet
M1968 GND N0364 N0363 GND efet
M1969 VDD N0943 ~TMP.2 GND efet
M1970 N0765 N0351 N0364 GND efet
M1971 N0555 N0872 N0913 GND efet
M1972 GND ACC.2 N0858 GND efet
M1973 GND N0348 ACC_0 GND efet
M1974 ~TMP.2 N0937 N0891 GND efet
M1975 N0606 M12 VDD GND efet
M1976 N0913 N0891 N0554 GND efet
M1977 VDD VDD N0473 GND efet
M1978 N0364 N0347 GND GND efet
M1979 GND N0879 N0876 GND efet
M1980 GND A22 N0288 GND efet
M1981 N0848 ADD-ACC ACC.2 GND efet
M1982 GND POC DCL.1 GND efet
M1983 GND M12 N0872 GND efet
M1984 VDD VDD N0665 GND efet
M1985 VDD VDD N0944 GND efet
M1986 GND N0943 N0944 GND efet
M1987 VDD N0747 A22 GND efet
M1988 N0345 N0347 GND GND efet
M1989 N0354 N0347 GND GND efet
M1990 N0370 N0347 GND GND efet
M1991 N0376 N0347 GND GND efet
M1992 VDD VDD N0355 GND efet
M1993 GND N0872 N0900 GND efet
M1994 N0900 N0556 GND GND efet
M1995 N0900 N0891 GND GND efet
M1996 N0473 M12 ACC.2 GND efet
M1997 N0473 N0858 GND GND efet
M1998 GND N0729 A22 GND efet
M1999 D2 ACB-IB N0348 GND efet
M2000 VDD VDD N0876 GND efet
M2001 N0514 ADSR ACC.2 GND efet
M2002 VDD VDD DCL.1 GND efet
M2003 GND N0913 N0917 GND efet
M2004 N0665 N0666 GND GND efet
M2005 GND N0848 ADD_0 GND efet
M2006 N0900 N0559 N0879 GND efet
M2007 VDD VDD N0917 GND efet
M2008 N0750 DCL.1 GND GND efet
M2009 TMP.2 N0944 VDD GND efet
M2010 GND N0943 TMP.2 GND efet
M2011 VDD VDD N0750 GND efet
M2012 GND N0355 N0354 GND efet
M2013 N0872 ACC-ADA N0473 GND efet
M2014 N0355 N0351 N0768 GND efet
M2015 VDD VDD N0879 GND efet
M2016 N0559 N0917 GND GND efet
M2017 N0848 ADD-IB D2 GND efet
M2018 D2 N0666 GND GND efet
M2019 N0747 N0729 GND GND efet
M2020 VDD VDD S00800 GND efet
M2021 VDD N0665 D2 GND efet
M2022 N0765 N0766 N0750 GND efet
M2023 TMP.2 SUB_GROUP(6) N0891 GND efet
M2024 N0355 N0348 GND GND efet
M2025 VDD VDD S00804 GND efet
M2026 VDD N0913 N0559 GND efet
M2027 N0943 S00801 VDD GND efet
M2028 VDD S00800 N0747 GND efet
M2029 N0345 N0348 GND GND efet
M2030 N0363 N0348 GND GND efet
M2031 N0370 N0348 GND GND efet
M2032 N0943 N0606 GND GND efet
M2033 N0376 N0348 GND GND efet
M2034 GND N0885 N0514 GND efet
M2035 ACC-ADA S00803 VDD GND efet
M2036 N0716 DCL.2 GND GND efet
M2037 VDD VDD N0349 GND efet
M2038 N0892 N0559 N0897 GND efet
M2039 N0558 N0559 N0557 GND efet
M2040 ADD_0 N0514 GND GND efet
M2041 D3 ADD-IB N0514 GND efet
M2042 VDD VDD S00803 GND efet
M2043 N0892 N0893 N0877 GND efet
M2044 VDD VDD S00801 GND efet
M2045 GND N0873 N0897 GND efet
M2046 N0557 N0873 GND GND efet
M2047 N0558 N0893 GND GND efet
M2048 N0728 CLK1 N0729 GND efet
M2049 DCL.2 N0768 GND GND efet
M2050 VDD VDD N0666 GND efet
M2051 N0728 N0286 GND GND efet
M2052 N0345 N0349 GND GND efet
M2053 N0514 N0877 VDD GND efet
M2054 N0349 N0356 GND GND efet
M2055 VDD VDD N0728 GND efet
M2056 ~TMP.3 N0946 GND GND efet
M2057 N0474 ACC-ADAC N0873 GND efet
M2058 GND D2_PAD N0666 GND efet
M2059 GND N0676 N0666 GND efet
M2060 N0286 CLK2 A12 GND efet
M2061 VDD VDD DCL.2 GND efet
M2062 N0356 ACB-IB D3 GND efet
M2063 N0354 N0356 GND GND efet
M2064 VDD S00804 N0914 GND efet
M2065 VDD N0945 ~TMP.3 GND efet
M2066 GND POC DCL.2 GND efet
M2067 N0363 N0356 GND GND efet
M2068 N0370 N0356 GND GND efet
M2069 N0376 N0356 GND GND efet
M2070 N0848 ADSL ACC.3 GND efet
M2071 VDD VDD N0474 GND efet
M2072 ACC.3 M12 N0474 GND efet
M2073 GND N0859 N0474 GND efet
M2074 ~TMP.3 SUB_GROUP(6) N0893 GND efet
M2075 N0558 N0873 N0914 GND efet
M2076 N0914 N0893 N0557 GND efet
M2077 GND N0356 ACC_0 GND efet
M2078 VDD VDD N0749 GND efet
M2079 GND N0877 N0885 GND efet
M2080 GND A12 N0288 GND efet
M2081 GND N0852 N0356 GND efet
M2082 N0749 DCL.2 GND GND efet
M2083 VDD VDD N0946 GND efet
M2084 GND N0945 N0946 GND efet
M2085 VDD N0748 A12 GND efet
M2086 N0859 ACC.3 GND GND efet
M2087 N0514 ADD-ACC ACC.3 GND efet
M2088 GND N0873 N0901 GND efet
M2089 N0901 N0559 GND GND efet
M2090 GND N0893 N0901 GND efet
M2091 GND N0731 A12 GND efet
M2092 VDD VDD N0356 GND efet
M2093 N0513 ADSL N0514 GND efet
M2094 N0918 N0914 GND GND efet
M2095 N0901 N0861 N0877 GND efet
M2096 VDD VDD N0859 GND efet
M2097 N0607 M12 VDD GND efet
M2098 VDD VDD N0918 GND efet
M2099 VDD VDD N0885 GND efet
M2100 N0768 N0766 N0749 GND efet
M2101 GND N0377 N0358 GND efet
M2102 N0513 ADSR ACC.3 GND efet
M2103 VDD M12 N0873 GND efet
M2104 TMP.3 N0946 VDD GND efet
M2105 GND N0945 TMP.3 GND efet
M2106 GND N0354 N0358 GND efet
M2107 N0358 N0363 GND GND efet
M2108 N0358 N0370 GND GND efet
M2109 GND N0403 N0358 GND efet
M2110 N0358 N0345 GND GND efet
M2111 TMP.3 N0937 N0893 GND efet
M2112 VDD VDD N0877 GND efet
M2113 N0861 N0918 GND GND efet
M2114 N0859 N0854 N0852 GND efet
M2115 D3 N0964 N0607 GND efet
M2116 VDD VDD S00817 GND efet
M2117 VDD VDD S00814 GND efet
M2118 N0873 ACC-ADA N0859 GND efet
M2119 N0748 N0731 GND GND efet
M2120 VDD VDD N0358 GND efet
M2121 GND GND D2_PAD GND efet
M2122 VDD N0914 N0861 GND efet
M2123 VDD S00814 N0748 GND efet
M2124 D3 N0415 N0358 GND efet
M2125 D2 N0415 N0366 GND efet
M2126 GND N0607 N0945 GND efet
M2127 VDD VDD S00819 GND efet
M2128 GND N0749 N0714 GND efet
M2129 N0945 S00817 VDD GND efet
M2130 VDD VDD S00818 GND efet
M2131 GND D0_PAD N0670 GND efet
M2132 N0668 D1_PAD GND GND efet
M2133 N0730 CLK1 N0731 GND efet
M2134 N0366 N0354 GND GND efet
M2135 GND N0363 N0366 GND efet
M2136 GND N0370 N0366 GND efet
M2137 GND N0377 N0366 GND efet
M2138 N0366 TCS GND GND efet
M2139 N0730 N0287 GND GND efet
M2140 N0714 ~COM GND GND efet
M2141 N0937 S00819 VDD GND efet
M2142 VDD VDD N0730 GND efet
M2143 VDD S00818 N0714 GND efet
M2144 GND GND D0_PAD GND efet
M2145 D0 N0670 GND GND efet
M2146 N0669 N0670 GND GND efet
M2147 GND GND D1_PAD GND efet
M2148 VDD VDD N0366 GND efet
M2149 N0287 CLK2 N0288 GND efet
M2150 D1 N0415 N0359 GND efet
M2151 D0 N0415 N0357 GND efet
M2152 N0669 N0676 GND GND efet
M2153 D3 N0664 GND GND efet
M2154 VDD N0663 D3 GND efet
M2155 D1 N0668 GND GND efet
M2156 N0667 N0668 GND GND efet
M2157 GND N0750 N0715 GND efet
M2158 VDD VDD N0288 GND efet
M2159 N0667 N0676 GND GND efet
M2160 N0674 D0 GND GND efet
M2161 D3_PAD POC GND GND efet
M2162 N0673 D1 GND GND efet
M2163 VDD VDD N0359 GND efet
M2164 GND N0345 N0359 GND efet
M2165 GND N0370 N0359 GND efet
M2166 GND N0377 N0359 GND efet
M2167 N0359 TCS GND GND efet
M2168 VDD VDD N0669 GND efet
M2169 VDD VDD S00825 GND efet
M2170 GND N0676 N0670 GND efet
M2171 N0668 N0676 GND GND efet
M2172 N0715 ~COM GND GND efet
M2173 VDD VDD N0674 GND efet
M2174 N0674 N0702 N0697 GND efet
M2175 VDD VDD N0673 GND efet
M2176 GND N0714 N0734 GND efet
M2177 VDD S00825 N0715 GND efet
M2178 N0673 N0702 N0694 GND efet
M2179 VDD VDD N0667 GND efet
M2180 CMRAM3 N0714 VDD GND efet
M2181 CMRAM2 N0715 VDD GND efet
M2182 VDD VDD N0734 GND efet
M2183 VDD VDD N0735 GND efet
M2184 GND N0715 N0735 GND efet
M2185 VDD N0669 D0 GND efet
M2186 VDD N0667 D1 GND efet
M2187 VDD VDD N0357 GND efet
M2188 VDD VDD N0670 GND efet
M2189 VDD VDD N0668 GND efet
M2190 GND N0345 N0357 GND efet
M2191 GND N0363 N0357 GND efet
M2192 GND N0377 N0357 GND efet
M2193 GND N0403 N0357 GND efet
M2194 GND ~COM N0716 GND efet
M2195 N0854 S00828 VDD GND efet
M2196 GND ~COM N0713 GND efet
M2197 VDD VDD S00833 GND efet
M2198 CMRAM2 N0735 GND GND efet
M2199 GND N0751 N0713 GND efet
M2200 GND N0734 CMRAM3 GND efet
M2201 VDD S00833 N0716 GND efet
M2202 VDD VDD S00828 GND efet
M2203 GND N0697 N0696 GND efet
M2204 GND N0694 N0693 GND efet
M2205 D0_PAD N0696 VDD GND efet
M2206 GND N0700 N0696 GND efet
M2207 VDD VDD S00834 GND efet
M2208 D1_PAD N0693 VDD GND efet
M2209 GND N0700 N0693 GND efet
M2210 VDD VDD N0664 GND efet
M2211 VDD VDD S00835 GND efet
M2212 VDD VDD S00836 GND efet
M2213 N0713 S00834 VDD GND efet
M2214 N0696 S00835 VDD GND efet
M2215 N0693 S00836 VDD GND efet
M2216 VDD VDD N0663 GND efet
M2217 GND N0676 N0664 GND efet
M2218 GND N0713 N0733 GND efet
M2219 CMRAM1 N0713 VDD GND efet
M2220 CMRAM0 N0716 VDD GND efet
M2221 VDD VDD N0733 GND efet
M2222 VDD VDD N0736 GND efet
M2223 GND N0716 N0736 GND efet
M2224 D0_PAD N0698 GND GND efet
M2225 D1_PAD N0695 GND GND efet
M2226 N0664 D3_PAD GND GND efet
M2227 GND N0664 N0663 GND efet
M2228 N0698 N0696 GND GND efet
M2229 GND N0700 N0698 GND efet
M2230 VDD S00839 N0698 GND efet
M2231 N0695 N0693 GND GND efet
M2232 GND N0700 N0695 GND efet
M2233 VDD S00840 N0695 GND efet
M2234 GND GND D3_PAD GND efet
M2235 GND N0676 N0663 GND efet
M2236 GND N0733 CMRAM1 GND efet
M2237 GND N0736 CMRAM0 GND efet
M2238 VDD VDD S00839 GND efet
M2239 VDD VDD S00840 GND efet
M2240 D0_PAD POC GND GND efet
M2241 D1_PAD POC GND GND efet
