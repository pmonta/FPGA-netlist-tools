* SPICE3 file created from 4002.ext - technology: nmos

.option scale=0.01u

M1000 diff_28920_288480# diff_35880_289800# GND GND efet w=7740 l=720
+ ad=2.97504e+07 pd=58560 as=-2.91681e+08 ps=7.19088e+06 
M1001 d1 GND GND GND efet w=10560 l=840
+ ad=1.79222e+08 pd=303360 as=0 ps=0 
M1002 GND diff_8760_228840# diff_28920_288480# GND efet w=21540 l=720
+ ad=0 pd=0 as=0 ps=0 
M1003 GND d1 diff_9720_284520# GND efet w=5580 l=660
+ ad=0 pd=0 as=1.31616e+07 ps=29040 
M1004 GND diff_8760_228840# diff_35880_289800# GND efet w=22320 l=660
+ ad=0 pd=0 as=3.87216e+07 ps=76080 
M1005 diff_35880_289800# diff_45720_287880# GND GND efet w=21180 l=780
+ ad=0 pd=0 as=0 ps=0 
M1006 diff_28920_288480# diff_28920_285720# diff_28920_288480# GND efet w=4020 l=1320
+ ad=0 pd=0 as=0 ps=0 
M1007 GND diff_9720_284520# diff_16560_282240# GND efet w=2220 l=780
+ ad=0 pd=0 as=1.43856e+07 ps=27360 
M1008 diff_9720_284520# diff_9720_284520# diff_9720_284520# GND efet w=240 l=480
+ ad=0 pd=0 as=0 ps=0 
M1009 diff_9720_284520# diff_9720_284520# diff_9720_284520# GND efet w=180 l=180
+ ad=0 pd=0 as=0 ps=0 
M1010 diff_16560_282240# diff_16560_282240# diff_16560_282240# GND efet w=360 l=360
+ ad=0 pd=0 as=0 ps=0 
M1011 diff_16560_282240# diff_16560_282240# diff_16560_282240# GND efet w=120 l=480
+ ad=0 pd=0 as=0 ps=0 
M1012 diff_9720_284520# Vdd Vdd GND efet w=960 l=3540
+ ad=0 pd=0 as=1.76661e+09 ps=3.49416e+06 
M1013 GND diff_13200_279960# diff_9720_284520# GND efet w=3480 l=720
+ ad=0 pd=0 as=0 ps=0 
M1014 diff_16560_282240# diff_13200_279960# GND GND efet w=3660 l=720
+ ad=0 pd=0 as=0 ps=0 
M1015 GND diff_28920_288480# d1 GND efet w=112380 l=420
+ ad=0 pd=0 as=0 ps=0 
M1016 diff_35880_289800# diff_38640_285720# diff_35880_289800# GND efet w=4260 l=1320
+ ad=0 pd=0 as=0 ps=0 
M1017 diff_28920_288480# diff_28920_285720# Vdd GND efet w=1140 l=900
+ ad=0 pd=0 as=0 ps=0 
M1018 diff_28920_285720# diff_28920_285720# diff_28920_285720# GND efet w=300 l=420
+ ad=2.2032e+06 pd=7680 as=0 ps=0 
M1019 diff_28920_285720# diff_28920_285720# diff_28920_285720# GND efet w=180 l=780
+ ad=0 pd=0 as=0 ps=0 
M1020 diff_35880_289800# diff_38640_285720# Vdd GND efet w=1140 l=900
+ ad=0 pd=0 as=0 ps=0 
M1021 diff_38640_285720# diff_38640_285720# diff_38640_285720# GND efet w=300 l=420
+ ad=2.1168e+06 pd=7200 as=0 ps=0 
M1022 diff_38640_285720# diff_38640_285720# diff_38640_285720# GND efet w=180 l=780
+ ad=0 pd=0 as=0 ps=0 
M1023 diff_28920_285720# Vdd Vdd GND efet w=960 l=720
+ ad=0 pd=0 as=0 ps=0 
M1024 Vdd Vdd Vdd GND efet w=240 l=480
+ ad=0 pd=0 as=0 ps=0 
M1025 Vdd Vdd Vdd GND efet w=120 l=120
+ ad=0 pd=0 as=0 ps=0 
M1026 Vdd Vdd diff_16560_282240# GND efet w=840 l=3780
+ ad=0 pd=0 as=0 ps=0 
M1027 diff_25200_276600# diff_16560_282240# Vdd GND efet w=3840 l=960
+ ad=1.30234e+08 pd=281280 as=0 ps=0 
M1028 GND diff_9720_284520# diff_25200_276600# GND efet w=3840 l=720
+ ad=0 pd=0 as=0 ps=0 
M1029 d0 GND GND GND efet w=10800 l=840
+ ad=1.7437e+08 pd=305040 as=0 ps=0 
M1030 GND diff_8760_228840# diff_126240_288840# GND efet w=21120 l=720
+ ad=0 pd=0 as=2.9664e+07 ps=57840 
M1031 GND d0 diff_94320_284400# GND efet w=5520 l=720
+ ad=0 pd=0 as=1.27728e+07 ps=28560 
M1032 diff_126240_288840# diff_133080_289920# GND GND efet w=7560 l=720
+ ad=0 pd=0 as=0 ps=0 
M1033 GND diff_8760_228840# diff_133080_289920# GND efet w=21780 l=780
+ ad=0 pd=0 as=3.8304e+07 ps=71760 
M1034 diff_133080_289920# diff_142920_287880# GND GND efet w=21240 l=720
+ ad=0 pd=0 as=0 ps=0 
M1035 GND diff_94320_284400# diff_100920_281280# GND efet w=2160 l=720
+ ad=0 pd=0 as=1.46016e+07 ps=28800 
M1036 diff_94320_284400# diff_94320_284400# diff_94320_284400# GND efet w=240 l=600
+ ad=0 pd=0 as=0 ps=0 
M1037 diff_100920_281280# diff_100920_281280# diff_100920_281280# GND efet w=600 l=480
+ ad=0 pd=0 as=0 ps=0 
M1038 d1 diff_35880_289800# Vdd GND efet w=60600 l=720
+ ad=0 pd=0 as=0 ps=0 
M1039 diff_45720_287880# diff_45720_287880# diff_45720_287880# GND efet w=240 l=960
+ ad=9.9648e+06 pd=22320 as=0 ps=0 
M1040 diff_38640_285720# Vdd Vdd GND efet w=840 l=840
+ ad=0 pd=0 as=0 ps=0 
M1041 diff_45720_287880# diff_45720_287880# diff_45720_287880# GND efet w=300 l=480
+ ad=0 pd=0 as=0 ps=0 
M1042 diff_100920_281280# diff_100920_281280# diff_100920_281280# GND efet w=180 l=540
+ ad=0 pd=0 as=0 ps=0 
M1043 diff_94320_284400# Vdd Vdd GND efet w=900 l=3540
+ ad=0 pd=0 as=0 ps=0 
M1044 GND diff_13200_279960# diff_94320_284400# GND efet w=3480 l=720
+ ad=0 pd=0 as=0 ps=0 
M1045 diff_100920_281280# diff_13200_279960# GND GND efet w=3480 l=720
+ ad=0 pd=0 as=0 ps=0 
M1046 diff_126240_288840# diff_126120_285720# diff_126240_288840# GND efet w=3660 l=3180
+ ad=0 pd=0 as=0 ps=0 
M1047 GND diff_126240_288840# d0 GND efet w=111540 l=420
+ ad=0 pd=0 as=0 ps=0 
M1048 diff_133080_289920# diff_135840_285600# diff_133080_289920# GND efet w=3420 l=3360
+ ad=0 pd=0 as=0 ps=0 
M1049 o0 diff_191640_286080# GND GND efet w=19800 l=720
+ ad=3.83328e+07 pd=69120 as=0 ps=0 
M1050 diff_191640_286080# diff_201720_295920# GND GND efet w=11040 l=720
+ ad=1.37088e+07 pd=28320 as=0 ps=0 
M1051 diff_192360_286440# diff_191640_286080# GND GND efet w=4800 l=720
+ ad=9.3744e+06 pd=17280 as=0 ps=0 
M1052 diff_201600_290400# diff_191640_286080# GND GND efet w=2400 l=720
+ ad=5.6736e+06 pd=13680 as=0 ps=0 
M1053 diff_201720_295920# diff_205080_288960# diff_201600_290400# GND efet w=1320 l=720
+ ad=1.47024e+07 pd=31920 as=0 ps=0 
M1054 GND diff_207720_290040# diff_201720_295920# GND efet w=2520 l=720
+ ad=0 pd=0 as=0 ps=0 
M1055 diff_192360_286440# diff_192360_286440# diff_192360_286440# GND efet w=360 l=480
+ ad=0 pd=0 as=0 ps=0 
M1056 diff_192360_286440# diff_192360_286440# diff_192360_286440# GND efet w=120 l=240
+ ad=0 pd=0 as=0 ps=0 
M1057 o0 diff_192360_286440# Vdd GND efet w=21180 l=660
+ ad=0 pd=0 as=0 ps=0 
M1058 d0 diff_133080_289920# Vdd GND efet w=60900 l=720
+ ad=0 pd=0 as=0 ps=0 
M1059 diff_126240_288840# diff_126120_285720# Vdd GND efet w=1020 l=780
+ ad=0 pd=0 as=0 ps=0 
M1060 diff_126120_285720# diff_126120_285720# diff_126120_285720# GND efet w=240 l=420
+ ad=2.1024e+06 pd=6960 as=0 ps=0 
M1061 diff_126120_285720# diff_126120_285720# diff_126120_285720# GND efet w=120 l=600
+ ad=0 pd=0 as=0 ps=0 
M1062 diff_135840_285600# diff_135840_285600# diff_135840_285600# GND efet w=240 l=420
+ ad=1.9728e+06 pd=6720 as=0 ps=0 
M1063 diff_135840_285600# diff_135840_285600# diff_135840_285600# GND efet w=180 l=540
+ ad=0 pd=0 as=0 ps=0 
M1064 Vdd Vdd Vdd GND efet w=240 l=600
+ ad=0 pd=0 as=0 ps=0 
M1065 diff_45720_287880# diff_22200_108240# diff_25200_276600# GND efet w=2940 l=720
+ ad=0 pd=0 as=0 ps=0 
M1066 Vdd Vdd diff_100920_281280# GND efet w=840 l=3720
+ ad=0 pd=0 as=0 ps=0 
M1067 diff_34920_109680# diff_100920_281280# Vdd GND efet w=3720 l=720
+ ad=1.1844e+08 pd=248160 as=0 ps=0 
M1068 GND diff_94320_284400# diff_34920_109680# GND efet w=3900 l=780
+ ad=0 pd=0 as=0 ps=0 
M1069 diff_126120_285720# Vdd Vdd GND efet w=1020 l=900
+ ad=0 pd=0 as=0 ps=0 
M1070 diff_133080_289920# diff_135840_285600# Vdd GND efet w=960 l=840
+ ad=0 pd=0 as=0 ps=0 
M1071 Vdd Vdd diff_135840_285600# GND efet w=780 l=840
+ ad=0 pd=0 as=0 ps=0 
M1072 Vdd Vdd Vdd GND efet w=120 l=120
+ ad=0 pd=0 as=0 ps=0 
M1073 diff_192360_286440# Vdd Vdd GND efet w=960 l=1920
+ ad=0 pd=0 as=0 ps=0 
M1074 diff_201600_290400# Vdd Vdd GND efet w=720 l=3000
+ ad=0 pd=0 as=0 ps=0 
M1075 GND diff_207480_277200# diff_205080_288960# GND efet w=1320 l=720
+ ad=0 pd=0 as=2.9664e+06 ps=7440 
M1076 diff_205080_288960# Vdd Vdd GND efet w=780 l=5700
+ ad=0 pd=0 as=0 ps=0 
M1077 Vdd Vdd Vdd GND efet w=480 l=840
+ ad=0 pd=0 as=0 ps=0 
M1078 Vdd Vdd Vdd GND efet w=540 l=420
+ ad=0 pd=0 as=0 ps=0 
M1079 diff_191640_286080# Vdd Vdd GND efet w=1140 l=1860
+ ad=0 pd=0 as=0 ps=0 
M1080 GND diff_241560_285240# diff_237360_275280# GND efet w=4920 l=720
+ ad=0 pd=0 as=1.15056e+07 ps=18720 
M1081 GND diff_241560_285240# o1 GND efet w=20280 l=600
+ ad=0 pd=0 as=4.12416e+07 ps=70800 
M1082 diff_201720_295920# diff_207480_277200# diff_210480_277440# GND efet w=1920 l=660
+ ad=0 pd=0 as=2.88e+06 ps=7920 
M1083 Vdd diff_6840_236160# d2 GND efet w=62340 l=660
+ ad=0 pd=0 as=1.89403e+08 ps=306960 
M1084 GND diff_6960_253440# d2 GND efet w=114420 l=420
+ ad=0 pd=0 as=0 ps=0 
M1085 diff_142920_287880# diff_22200_108240# diff_34920_109680# GND efet w=2640 l=720
+ ad=8.208e+06 pd=17040 as=0 ps=0 
M1086 diff_210480_277440# clk2 diff_34920_109680# GND efet w=1800 l=720
+ ad=0 pd=0 as=0 ps=0 
M1087 diff_237360_275280# Vdd Vdd GND efet w=1080 l=1920
+ ad=0 pd=0 as=0 ps=0 
M1088 diff_237360_275280# diff_237360_275280# diff_237360_275280# GND efet w=420 l=420
+ ad=0 pd=0 as=0 ps=0 
M1089 o1 diff_237360_275280# Vdd GND efet w=20940 l=660
+ ad=0 pd=0 as=0 ps=0 
M1090 GND diff_241560_285240# diff_245400_273720# GND efet w=2640 l=840
+ ad=0 pd=0 as=6.5952e+06 ps=14640 
M1091 diff_245400_273720# Vdd Vdd GND efet w=1080 l=2880
+ ad=0 pd=0 as=0 ps=0 
M1092 Vdd Vdd Vdd GND efet w=360 l=840
+ ad=0 pd=0 as=0 ps=0 
M1093 Vdd Vdd Vdd GND efet w=360 l=840
+ ad=0 pd=0 as=0 ps=0 
M1094 GND diff_234600_265200# diff_241560_285240# GND efet w=11160 l=540
+ ad=0 pd=0 as=1.4112e+07 ps=27600 
M1095 diff_245400_273720# diff_242400_271320# diff_234600_265200# GND efet w=1440 l=840
+ ad=0 pd=0 as=1.6344e+07 ps=32640 
M1096 diff_242400_271320# Vdd Vdd GND efet w=840 l=5760
+ ad=3.456e+06 pd=7920 as=0 ps=0 
M1097 diff_242400_271320# diff_207480_277200# GND GND efet w=1500 l=660
+ ad=0 pd=0 as=0 ps=0 
M1098 diff_234600_265200# diff_207720_290040# GND GND efet w=2520 l=660
+ ad=0 pd=0 as=0 ps=0 
M1099 Vdd Vdd Vdd GND efet w=300 l=420
+ ad=0 pd=0 as=0 ps=0 
M1100 Vdd Vdd Vdd GND efet w=240 l=720
+ ad=0 pd=0 as=0 ps=0 
M1101 diff_48720_260280# diff_32640_245760# diff_34920_109680# GND efet w=3840 l=720
+ ad=9.8928e+06 pd=22800 as=0 ps=0 
M1102 diff_48720_260280# diff_52320_146760# diff_50640_260400# GND efet w=3840 l=720
+ ad=0 pd=0 as=1.73808e+07 ps=34080 
M1103 diff_54840_260160# diff_42600_159120# diff_48720_260280# GND efet w=4620 l=780
+ ad=3.17376e+07 pd=86400 as=0 ps=0 
M1104 diff_232560_264480# clk2 diff_25200_276600# GND efet w=2040 l=720
+ ad=3.2112e+06 pd=8160 as=0 ps=0 
M1105 diff_234600_265200# diff_207480_277200# diff_232560_264480# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M1106 diff_56760_259080# Vdd Vdd GND efet w=840 l=3000
+ ad=9.1872e+06 pd=22560 as=0 ps=0 
M1107 Vdd diff_66360_261120# diff_50640_260400# GND efet w=1560 l=720
+ ad=0 pd=0 as=0 ps=0 
M1108 diff_56760_259080# diff_42360_242040# diff_54840_260160# GND efet w=3240 l=720
+ ad=0 pd=0 as=0 ps=0 
M1109 diff_48720_255480# diff_32640_245760# diff_25200_276600# GND efet w=3840 l=720
+ ad=9.8928e+06 pd=22800 as=0 ps=0 
M1110 diff_56760_255360# diff_42360_242040# diff_54840_253440# GND efet w=3180 l=780
+ ad=9.216e+06 pd=21840 as=3.20976e+07 ps=88560 
M1111 diff_50640_260400# diff_56760_259080# GND GND efet w=5520 l=840
+ ad=0 pd=0 as=0 ps=0 
M1112 diff_56760_259080# diff_66360_261120# GND GND efet w=2700 l=780
+ ad=0 pd=0 as=0 ps=0 
M1113 GND diff_56760_255360# diff_50640_253320# GND efet w=5400 l=840
+ ad=0 pd=0 as=1.7352e+07 ps=33360 
M1114 diff_81360_258480# diff_80400_261120# GND GND efet w=2280 l=720
+ ad=2.4048e+06 pd=7200 as=0 ps=0 
M1115 diff_54840_260160# diff_84360_149760# diff_80400_261120# GND efet w=960 l=720
+ ad=0 pd=0 as=2.6928e+06 ps=7440 
M1116 diff_88080_261360# diff_87240_145800# diff_54840_260160# GND efet w=960 l=720
+ ad=2.6208e+06 pd=7440 as=0 ps=0 
M1117 diff_66360_261120# diff_80760_144360# diff_81360_258480# GND efet w=2160 l=840
+ ad=6.47136e+07 pd=154080 as=0 ps=0 
M1118 diff_66480_253440# diff_80760_144360# diff_81360_254280# GND efet w=2220 l=960
+ ad=6.18336e+07 pd=154800 as=2.4192e+06 ps=7440 
M1119 diff_6840_236160# diff_8760_249240# GND GND efet w=21540 l=660
+ ad=3.94128e+07 pd=78720 as=0 ps=0 
M1120 diff_8760_249240# diff_8760_249240# diff_8760_249240# GND efet w=180 l=660
+ ad=1.1592e+07 pd=21840 as=0 ps=0 
M1121 diff_8760_249240# diff_8760_249240# diff_8760_249240# GND efet w=300 l=420
+ ad=0 pd=0 as=0 ps=0 
M1122 diff_23040_212640# diff_22200_108240# diff_8760_249240# GND efet w=2760 l=720
+ ad=1.18325e+08 pd=248400 as=0 ps=0 
M1123 diff_48720_249120# diff_32640_245760# diff_23040_212640# GND efet w=3840 l=720
+ ad=9.6048e+06 pd=22800 as=0 ps=0 
M1124 diff_48720_255480# diff_52320_146760# diff_50640_253320# GND efet w=3840 l=720
+ ad=0 pd=0 as=0 ps=0 
M1125 diff_54840_253440# diff_42600_159120# diff_48720_255480# GND efet w=4500 l=780
+ ad=0 pd=0 as=0 ps=0 
M1126 GND diff_66480_253440# diff_56760_255360# GND efet w=2640 l=720
+ ad=0 pd=0 as=0 ps=0 
M1127 GND diff_32640_245760# diff_44040_244680# GND efet w=5220 l=780
+ ad=0 pd=0 as=5.7456e+06 ps=12720 
M1128 diff_48720_249120# diff_52320_146760# diff_50640_246720# GND efet w=3720 l=720
+ ad=0 pd=0 as=1.7136e+07 ps=32400 
M1129 diff_54840_246000# diff_42600_159120# diff_48720_249120# GND efet w=4500 l=780
+ ad=3.11616e+07 pd=85920 as=0 ps=0 
M1130 Vdd diff_66480_253440# diff_50640_253320# GND efet w=1500 l=720
+ ad=0 pd=0 as=0 ps=0 
M1131 diff_81360_254280# diff_80400_252840# GND GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1132 diff_56760_255360# Vdd Vdd GND efet w=720 l=2760
+ ad=0 pd=0 as=0 ps=0 
M1133 Vdd Vdd Vdd GND efet w=600 l=360
+ ad=0 pd=0 as=0 ps=0 
M1134 Vdd Vdd Vdd GND efet w=420 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1135 diff_56760_245040# Vdd Vdd GND efet w=720 l=2760
+ ad=9.6912e+06 pd=23280 as=0 ps=0 
M1136 diff_56760_245040# diff_42360_242040# diff_54840_246000# GND efet w=3240 l=720
+ ad=0 pd=0 as=0 ps=0 
M1137 diff_44040_244680# diff_42600_159120# diff_42360_242040# GND efet w=4860 l=780
+ ad=0 pd=0 as=9.864e+06 ps=20400 
M1138 diff_6840_236160# diff_8760_228840# GND GND efet w=21540 l=780
+ ad=0 pd=0 as=0 ps=0 
M1139 Vdd diff_16200_238800# diff_6840_236160# GND efet w=1080 l=840
+ ad=0 pd=0 as=0 ps=0 
M1140 Vdd Vdd diff_42360_242040# GND efet w=1200 l=3900
+ ad=0 pd=0 as=0 ps=0 
M1141 diff_6840_236160# diff_16200_238800# diff_6840_236160# GND efet w=4860 l=1800
+ ad=0 pd=0 as=0 ps=0 
M1142 diff_16200_238800# diff_16200_238800# diff_16200_238800# GND efet w=300 l=780
+ ad=2.376e+06 pd=7680 as=0 ps=0 
M1143 Vdd Vdd diff_16200_238800# GND efet w=960 l=840
+ ad=0 pd=0 as=0 ps=0 
M1144 diff_16200_238800# diff_16200_238800# diff_16200_238800# GND efet w=180 l=360
+ ad=0 pd=0 as=0 ps=0 
M1145 Vdd Vdd Vdd GND efet w=240 l=720
+ ad=0 pd=0 as=0 ps=0 
M1146 Vdd Vdd Vdd GND efet w=180 l=360
+ ad=0 pd=0 as=0 ps=0 
M1147 Vdd diff_66360_247080# diff_50640_246720# GND efet w=1320 l=660
+ ad=0 pd=0 as=0 ps=0 
M1148 diff_50640_246720# diff_56760_245040# GND GND efet w=5220 l=780
+ ad=0 pd=0 as=0 ps=0 
M1149 diff_95160_258480# diff_94080_261120# GND GND efet w=2280 l=960
+ ad=2.376e+06 pd=7440 as=0 ps=0 
M1150 diff_90480_258120# diff_89400_145800# diff_66360_261120# GND efet w=2160 l=720
+ ad=2.6496e+06 pd=7680 as=0 ps=0 
M1151 GND diff_88080_261360# diff_90480_258120# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1152 diff_54840_260160# diff_98160_145800# diff_94080_261120# GND efet w=1020 l=720
+ ad=0 pd=0 as=2.6784e+06 ps=7440 
M1153 diff_101760_261360# diff_100920_145800# diff_54840_260160# GND efet w=960 l=720
+ ad=2.592e+06 pd=7680 as=0 ps=0 
M1154 diff_66360_261120# diff_94560_144240# diff_95160_258480# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1155 diff_90480_254760# diff_89400_145800# diff_66480_253440# GND efet w=2160 l=720
+ ad=2.6784e+06 pd=7680 as=0 ps=0 
M1156 diff_66480_253440# diff_94560_144240# diff_95040_256560# GND efet w=2160 l=900
+ ad=0 pd=0 as=2.4336e+06 ps=7920 
M1157 GND diff_88080_252840# diff_90480_254760# GND efet w=2340 l=780
+ ad=0 pd=0 as=0 ps=0 
M1158 diff_54840_253440# diff_84360_149760# diff_80400_252840# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6928e+06 ps=7680 
M1159 diff_88080_252840# diff_87240_145800# diff_54840_253440# GND efet w=840 l=720
+ ad=2.448e+06 pd=7440 as=0 ps=0 
M1160 diff_56760_245040# diff_66360_247080# GND GND efet w=2640 l=720
+ ad=0 pd=0 as=0 ps=0 
M1161 diff_56760_241080# diff_42360_242040# diff_54840_239280# GND efet w=3240 l=780
+ ad=9.6768e+06 pd=23280 as=3.15216e+07 ps=86640 
M1162 diff_81360_244320# diff_80400_246960# GND GND efet w=2280 l=720
+ ad=2.3184e+06 pd=7200 as=0 ps=0 
M1163 diff_54840_246000# diff_84360_149760# diff_80400_246960# GND efet w=840 l=720
+ ad=0 pd=0 as=2.5344e+06 ps=7440 
M1164 diff_88080_247200# diff_87240_145800# diff_54840_246000# GND efet w=840 l=720
+ ad=2.5056e+06 pd=7440 as=0 ps=0 
M1165 diff_66360_247080# diff_80760_144360# diff_81360_244320# GND efet w=2160 l=840
+ ad=6.49152e+07 pd=154320 as=0 ps=0 
M1166 diff_66480_239280# diff_80760_144360# diff_81360_240120# GND efet w=2220 l=780
+ ad=6.31296e+07 pd=155280 as=2.4336e+06 ps=7680 
M1167 GND diff_56760_241080# diff_50640_239280# GND efet w=5040 l=720
+ ad=0 pd=0 as=1.68624e+07 ps=32640 
M1168 GND diff_66480_239280# diff_56760_241080# GND efet w=2640 l=840
+ ad=0 pd=0 as=0 ps=0 
M1169 diff_6960_253440# diff_6840_236160# GND GND efet w=7920 l=600
+ ad=3.16368e+07 pd=60960 as=0 ps=0 
M1170 diff_48720_236880# diff_32640_245760# diff_23160_135720# GND efet w=3840 l=720
+ ad=9.6768e+06 pd=22800 as=1.27973e+08 ps=271680 
M1171 diff_48720_236880# diff_52320_146760# diff_50640_239280# GND efet w=3780 l=780
+ ad=0 pd=0 as=0 ps=0 
M1172 diff_54840_239280# diff_42600_159120# diff_48720_236880# GND efet w=4560 l=840
+ ad=0 pd=0 as=0 ps=0 
M1173 diff_50640_239280# diff_66480_239280# Vdd GND efet w=1380 l=780
+ ad=0 pd=0 as=0 ps=0 
M1174 diff_81360_240120# diff_80400_238680# GND GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M1175 diff_6960_253440# diff_8760_228840# GND GND efet w=21600 l=900
+ ad=0 pd=0 as=0 ps=0 
M1176 Vdd diff_16200_228600# diff_6960_253440# GND efet w=1140 l=780
+ ad=0 pd=0 as=0 ps=0 
M1177 diff_6960_253440# diff_16200_228600# diff_6960_253440# GND efet w=4020 l=1680
+ ad=0 pd=0 as=0 ps=0 
M1178 diff_16200_228600# diff_16200_228600# diff_16200_228600# GND efet w=240 l=720
+ ad=2.2464e+06 pd=7680 as=0 ps=0 
M1179 Vdd Vdd diff_16200_228600# GND efet w=840 l=840
+ ad=0 pd=0 as=0 ps=0 
M1180 diff_48720_231240# diff_32760_140400# diff_34920_109680# GND efet w=3840 l=720
+ ad=1.10448e+07 pd=25200 as=0 ps=0 
M1181 diff_48720_231240# diff_52320_146760# diff_50640_232080# GND efet w=3960 l=720
+ ad=0 pd=0 as=1.6704e+07 ps=33600 
M1182 diff_56760_241080# Vdd Vdd GND efet w=720 l=2760
+ ad=0 pd=0 as=0 ps=0 
M1183 Vdd Vdd Vdd GND efet w=360 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1184 Vdd Vdd Vdd GND efet w=600 l=360
+ ad=0 pd=0 as=0 ps=0 
M1185 diff_54840_231960# diff_42600_159120# diff_48720_231240# GND efet w=4500 l=780
+ ad=3.11328e+07 pd=86640 as=0 ps=0 
M1186 diff_56760_230880# Vdd Vdd GND efet w=720 l=2880
+ ad=8.928e+06 pd=21840 as=0 ps=0 
M1187 Vdd diff_66480_232800# diff_50640_232080# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M1188 diff_56760_230880# diff_42360_213840# diff_54840_231960# GND efet w=3240 l=720
+ ad=0 pd=0 as=0 ps=0 
M1189 diff_16200_228600# diff_16200_228600# diff_16200_228600# GND efet w=300 l=360
+ ad=0 pd=0 as=0 ps=0 
M1190 diff_48720_225840# diff_32760_140400# diff_25200_276600# GND efet w=3720 l=720
+ ad=9.5616e+06 pd=23040 as=0 ps=0 
M1191 diff_56760_227400# diff_42360_213840# diff_54840_225240# GND efet w=3180 l=780
+ ad=8.9136e+06 pd=21600 as=3.10608e+07 ps=85920 
M1192 diff_50640_232080# diff_56760_230880# GND GND efet w=5460 l=780
+ ad=0 pd=0 as=0 ps=0 
M1193 diff_95040_256560# diff_94080_252840# GND GND efet w=2340 l=780
+ ad=0 pd=0 as=0 ps=0 
M1194 diff_90480_243960# diff_89400_145800# diff_66360_247080# GND efet w=2160 l=720
+ ad=2.6352e+06 pd=7440 as=0 ps=0 
M1195 GND diff_88080_247200# diff_90480_243960# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1196 diff_95040_244320# diff_94080_247080# GND GND efet w=2340 l=780
+ ad=2.592e+06 pd=7440 as=0 ps=0 
M1197 diff_104280_258120# diff_103200_145800# diff_66360_261120# GND efet w=2160 l=720
+ ad=2.3904e+06 pd=7440 as=0 ps=0 
M1198 GND diff_101760_261360# diff_104280_258120# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1199 diff_108840_258480# diff_107880_261120# GND GND efet w=2280 l=720
+ ad=2.376e+06 pd=7200 as=0 ps=0 
M1200 diff_54840_260160# diff_111840_149760# diff_107880_261120# GND efet w=960 l=720
+ ad=0 pd=0 as=2.6928e+06 ps=7440 
M1201 diff_115560_261360# diff_114720_145800# diff_54840_260160# GND efet w=1140 l=660
+ ad=2.5776e+06 pd=7200 as=0 ps=0 
M1202 diff_66360_261120# diff_108240_144360# diff_108840_258480# GND efet w=2160 l=840
+ ad=0 pd=0 as=0 ps=0 
M1203 diff_104280_254640# diff_103200_145800# diff_66480_253440# GND efet w=2160 l=840
+ ad=2.3904e+06 pd=7440 as=0 ps=0 
M1204 diff_66480_253440# diff_108240_144360# diff_108840_254280# GND efet w=2160 l=900
+ ad=0 pd=0 as=2.376e+06 ps=7200 
M1205 diff_54840_253440# diff_98160_145800# diff_94080_252840# GND efet w=840 l=840
+ ad=0 pd=0 as=2.7216e+06 ps=7680 
M1206 diff_101760_252840# diff_100920_145800# diff_54840_253440# GND efet w=840 l=720
+ ad=2.592e+06 pd=7680 as=0 ps=0 
M1207 diff_54840_246000# diff_98160_145800# diff_94080_247080# GND efet w=840 l=840
+ ad=0 pd=0 as=2.5056e+06 ps=7680 
M1208 diff_101760_247200# diff_100920_145800# diff_54840_246000# GND efet w=840 l=720
+ ad=2.5776e+06 pd=7920 as=0 ps=0 
M1209 diff_66360_247080# diff_94560_144240# diff_95040_244320# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1210 diff_90480_240600# diff_89400_145800# diff_66480_239280# GND efet w=2160 l=720
+ ad=2.7072e+06 pd=7680 as=0 ps=0 
M1211 GND diff_88080_238680# diff_90480_240600# GND efet w=2340 l=780
+ ad=0 pd=0 as=0 ps=0 
M1212 diff_54840_239280# diff_84360_149760# diff_80400_238680# GND efet w=840 l=720
+ ad=0 pd=0 as=2.7072e+06 ps=7680 
M1213 diff_88080_238680# diff_87240_145800# diff_54840_239280# GND efet w=840 l=720
+ ad=2.5632e+06 pd=7200 as=0 ps=0 
M1214 diff_54840_231960# diff_84360_149760# diff_80400_232800# GND efet w=840 l=720
+ ad=0 pd=0 as=2.7072e+06 ps=7440 
M1215 diff_88080_233040# diff_87240_145800# diff_54840_231960# GND efet w=840 l=720
+ ad=2.592e+06 pd=7200 as=0 ps=0 
M1216 diff_56760_230880# diff_66480_232800# GND GND efet w=2700 l=780
+ ad=0 pd=0 as=0 ps=0 
M1217 diff_81360_230160# diff_80400_232800# GND GND efet w=2280 l=720
+ ad=2.3328e+06 pd=7200 as=0 ps=0 
M1218 GND diff_56760_227400# diff_50640_225120# GND efet w=5040 l=840
+ ad=0 pd=0 as=1.6488e+07 ps=32160 
M1219 diff_66480_232800# diff_80760_144360# diff_81360_230160# GND efet w=2160 l=840
+ ad=6.48e+07 pd=154320 as=0 ps=0 
M1220 diff_48720_220920# diff_32760_140400# diff_23040_212640# GND efet w=3720 l=720
+ ad=9.72e+06 pd=22800 as=0 ps=0 
M1221 diff_48720_225840# diff_52320_146760# diff_50640_225120# GND efet w=3720 l=720
+ ad=0 pd=0 as=0 ps=0 
M1222 diff_54840_225240# diff_42600_159120# diff_48720_225840# GND efet w=4680 l=720
+ ad=0 pd=0 as=0 ps=0 
M1223 GND diff_32760_140400# diff_44040_216360# GND efet w=5640 l=720
+ ad=0 pd=0 as=5.2992e+06 ps=12240 
M1224 diff_48720_220920# diff_52320_146760# diff_50640_218640# GND efet w=3840 l=720
+ ad=0 pd=0 as=1.6776e+07 ps=32880 
M1225 diff_54840_217800# diff_42600_159120# diff_48720_220920# GND efet w=4560 l=720
+ ad=3.14208e+07 pd=86640 as=0 ps=0 
M1226 GND diff_66480_225120# diff_56760_227400# GND efet w=2640 l=720
+ ad=0 pd=0 as=0 ps=0 
M1227 diff_50640_225120# diff_66480_225120# Vdd GND efet w=1380 l=720
+ ad=0 pd=0 as=0 ps=0 
M1228 diff_81360_225960# diff_80400_224520# GND GND efet w=2400 l=720
+ ad=2.4192e+06 pd=7440 as=0 ps=0 
M1229 diff_66480_225120# diff_80760_144360# diff_81360_225960# GND efet w=2160 l=840
+ ad=6.13728e+07 pd=152880 as=0 ps=0 
M1230 diff_56760_227400# Vdd Vdd GND efet w=600 l=2640
+ ad=0 pd=0 as=0 ps=0 
M1231 Vdd Vdd Vdd GND efet w=600 l=360
+ ad=0 pd=0 as=0 ps=0 
M1232 Vdd Vdd Vdd GND efet w=360 l=840
+ ad=0 pd=0 as=0 ps=0 
M1233 diff_56880_216720# Vdd Vdd GND efet w=600 l=2640
+ ad=9.6912e+06 pd=23280 as=0 ps=0 
M1234 diff_56880_216720# diff_42360_213840# diff_54840_217800# GND efet w=3360 l=840
+ ad=0 pd=0 as=0 ps=0 
M1235 diff_44040_216360# diff_42600_159120# diff_42360_213840# GND efet w=4680 l=840
+ ad=0 pd=0 as=9.6192e+06 ps=20400 
M1236 GND diff_16320_201240# diff_23040_212640# GND efet w=3840 l=720
+ ad=0 pd=0 as=0 ps=0 
M1237 d2 GND GND GND efet w=10560 l=720
+ ad=0 pd=0 as=0 ps=0 
M1238 diff_23040_212640# diff_17040_204360# Vdd GND efet w=3840 l=720
+ ad=0 pd=0 as=0 ps=0 
M1239 Vdd Vdd diff_42360_213840# GND efet w=1200 l=3840
+ ad=0 pd=0 as=0 ps=0 
M1240 Vdd Vdd Vdd GND efet w=240 l=720
+ ad=0 pd=0 as=0 ps=0 
M1241 Vdd Vdd Vdd GND efet w=180 l=360
+ ad=0 pd=0 as=0 ps=0 
M1242 Vdd diff_66480_218640# diff_50640_218640# GND efet w=1380 l=780
+ ad=0 pd=0 as=0 ps=0 
M1243 diff_50640_218640# diff_56880_216720# GND GND efet w=5280 l=840
+ ad=0 pd=0 as=0 ps=0 
M1244 diff_95040_240840# diff_94080_238680# GND GND efet w=2580 l=900
+ ad=2.5776e+06 pd=7920 as=0 ps=0 
M1245 diff_66480_239280# diff_94560_144240# diff_95040_240840# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1246 diff_90480_229800# diff_89400_145800# diff_66480_232800# GND efet w=2160 l=720
+ ad=2.6496e+06 pd=7680 as=0 ps=0 
M1247 GND diff_88080_233040# diff_90480_229800# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1248 diff_95160_230160# diff_94080_232920# GND GND efet w=2280 l=840
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1249 GND diff_101760_252840# diff_104280_254640# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1250 diff_108840_254280# diff_107760_253200# GND GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1251 diff_104280_243960# diff_103200_145800# diff_66360_247080# GND efet w=2160 l=720
+ ad=2.376e+06 pd=7200 as=0 ps=0 
M1252 GND diff_101760_247200# diff_104280_243960# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1253 diff_108840_244320# diff_107880_246960# GND GND efet w=2280 l=720
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1254 diff_117960_258120# diff_116880_145800# diff_66360_261120# GND efet w=2160 l=720
+ ad=2.6496e+06 pd=7440 as=0 ps=0 
M1255 GND diff_115560_261360# diff_117960_258120# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1256 diff_122640_258480# diff_121560_261120# GND GND efet w=2280 l=840
+ ad=2.376e+06 pd=7440 as=0 ps=0 
M1257 diff_54840_260160# diff_125640_145800# diff_121560_261120# GND efet w=960 l=780
+ ad=0 pd=0 as=2.5776e+06 ps=7680 
M1258 diff_129240_261360# diff_128400_145800# diff_54840_260160# GND efet w=960 l=720
+ ad=2.5344e+06 pd=7440 as=0 ps=0 
M1259 diff_66360_261120# diff_122040_144240# diff_122640_258480# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1260 diff_117960_254760# diff_116880_145800# diff_66480_253440# GND efet w=2160 l=720
+ ad=2.6496e+06 pd=7440 as=0 ps=0 
M1261 diff_54840_253440# diff_111840_149760# diff_107760_253200# GND efet w=840 l=720
+ ad=0 pd=0 as=2.664e+06 ps=7440 
M1262 diff_115560_252840# diff_114720_145800# diff_54840_253440# GND efet w=960 l=720
+ ad=2.5344e+06 pd=7200 as=0 ps=0 
M1263 diff_54840_246000# diff_111840_149760# diff_107880_246960# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6784e+06 ps=7440 
M1264 diff_115560_247200# diff_114720_145800# diff_54840_246000# GND efet w=900 l=720
+ ad=2.5056e+06 pd=7440 as=0 ps=0 
M1265 diff_66360_247080# diff_108240_144360# diff_108840_244320# GND efet w=2160 l=840
+ ad=0 pd=0 as=0 ps=0 
M1266 diff_104280_240480# diff_103200_145800# diff_66480_239280# GND efet w=2160 l=720
+ ad=2.4624e+06 pd=7440 as=0 ps=0 
M1267 diff_101760_238680# diff_100920_145800# diff_54840_239280# GND efet w=840 l=780
+ ad=2.592e+06 pd=7680 as=0 ps=0 
M1268 diff_54840_239280# diff_98160_145800# diff_94080_238680# GND efet w=840 l=840
+ ad=0 pd=0 as=2.664e+06 ps=7680 
M1269 diff_54840_231960# diff_98160_145800# diff_94080_232920# GND efet w=840 l=840
+ ad=0 pd=0 as=2.6208e+06 ps=7680 
M1270 diff_101760_233040# diff_100920_145800# diff_54840_231960# GND efet w=840 l=720
+ ad=2.6208e+06 pd=7680 as=0 ps=0 
M1271 diff_66480_232800# diff_94560_144240# diff_95160_230160# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1272 diff_90480_226440# diff_89400_145800# diff_66480_225120# GND efet w=2040 l=720
+ ad=2.6496e+06 pd=7440 as=0 ps=0 
M1273 diff_66480_225120# diff_94560_144240# diff_95160_225960# GND efet w=2100 l=900
+ ad=0 pd=0 as=2.4048e+06 ps=7440 
M1274 GND diff_88080_224520# diff_90480_226440# GND efet w=2340 l=780
+ ad=0 pd=0 as=0 ps=0 
M1275 diff_54840_225240# diff_84360_149760# diff_80400_224520# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6352e+06 ps=7440 
M1276 diff_88080_224520# diff_87240_145800# diff_54840_225240# GND efet w=840 l=720
+ ad=2.5776e+06 pd=7440 as=0 ps=0 
M1277 diff_54840_217800# diff_84360_149760# diff_80400_218760# GND efet w=960 l=720
+ ad=0 pd=0 as=2.6064e+06 ps=7440 
M1278 diff_88080_218880# diff_87240_145800# diff_54840_217800# GND efet w=960 l=720
+ ad=2.5632e+06 pd=7200 as=0 ps=0 
M1279 diff_95160_225960# diff_94080_224640# GND GND efet w=2400 l=900
+ ad=0 pd=0 as=0 ps=0 
M1280 diff_56880_216720# diff_66480_218640# GND GND efet w=2700 l=780
+ ad=0 pd=0 as=0 ps=0 
M1281 diff_56880_212760# diff_42360_213840# diff_54840_210960# GND efet w=3360 l=840
+ ad=9.36e+06 pd=23280 as=3.14064e+07 ps=87600 
M1282 GND diff_56880_212760# diff_50640_210960# GND efet w=5220 l=720
+ ad=0 pd=0 as=1.68624e+07 ps=32400 
M1283 diff_81360_216000# diff_80400_218760# GND GND efet w=2400 l=840
+ ad=2.6064e+06 pd=7440 as=0 ps=0 
M1284 diff_66480_218640# diff_80760_144360# diff_81360_216000# GND efet w=2100 l=780
+ ad=6.37488e+07 pd=154080 as=0 ps=0 
M1285 diff_48720_208560# diff_32760_140400# diff_23160_135720# GND efet w=3900 l=780
+ ad=9.9504e+06 pd=22800 as=0 ps=0 
M1286 diff_17040_204360# diff_16320_201240# GND GND efet w=2160 l=720
+ ad=1.50624e+07 pd=27600 as=0 ps=0 
M1287 diff_17040_204360# diff_17040_204360# diff_17040_204360# GND efet w=240 l=360
+ ad=0 pd=0 as=0 ps=0 
M1288 diff_17040_204360# diff_17040_204360# diff_17040_204360# GND efet w=240 l=840
+ ad=0 pd=0 as=0 ps=0 
M1289 Vdd Vdd diff_17040_204360# GND efet w=840 l=3720
+ ad=0 pd=0 as=0 ps=0 
M1290 diff_48720_208560# diff_52320_146760# diff_50640_210960# GND efet w=3840 l=720
+ ad=0 pd=0 as=0 ps=0 
M1291 diff_54840_210960# diff_42600_159120# diff_48720_208560# GND efet w=4500 l=780
+ ad=0 pd=0 as=0 ps=0 
M1292 GND diff_66480_210960# diff_56880_212760# GND efet w=2760 l=840
+ ad=0 pd=0 as=0 ps=0 
M1293 diff_81360_211920# diff_80400_210360# GND GND efet w=2280 l=720
+ ad=2.6064e+06 pd=7440 as=0 ps=0 
M1294 diff_66480_210960# diff_80760_144360# diff_81360_211920# GND efet w=2160 l=720
+ ad=6.44688e+07 pd=155040 as=0 ps=0 
M1295 diff_50640_210960# diff_66480_210960# Vdd GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M1296 diff_56880_212760# Vdd Vdd GND efet w=600 l=2640
+ ad=0 pd=0 as=0 ps=0 
M1297 diff_16320_201240# diff_16320_201240# diff_16320_201240# GND efet w=240 l=720
+ ad=1.19808e+07 pd=28080 as=0 ps=0 
M1298 diff_16320_201240# diff_16320_201240# diff_16320_201240# GND efet w=180 l=780
+ ad=0 pd=0 as=0 ps=0 
M1299 diff_16320_201240# d2 GND GND efet w=5640 l=840
+ ad=0 pd=0 as=0 ps=0 
M1300 diff_17040_204360# diff_13200_279960# GND GND efet w=3480 l=660
+ ad=0 pd=0 as=0 ps=0 
M1301 diff_48720_202920# diff_33120_151080# diff_34920_109680# GND efet w=3840 l=720
+ ad=1.09728e+07 pd=24720 as=0 ps=0 
M1302 diff_48720_202920# diff_52320_146760# diff_50640_203760# GND efet w=3840 l=720
+ ad=0 pd=0 as=1.68192e+07 ps=32640 
M1303 Vdd Vdd Vdd GND efet w=600 l=360
+ ad=0 pd=0 as=0 ps=0 
M1304 diff_54840_203640# diff_42600_159120# diff_48720_202920# GND efet w=4500 l=780
+ ad=3.18528e+07 pd=86400 as=0 ps=0 
M1305 Vdd Vdd Vdd GND efet w=360 l=840
+ ad=0 pd=0 as=0 ps=0 
M1306 diff_56880_202560# Vdd Vdd GND efet w=660 l=2700
+ ad=8.7552e+06 pd=21840 as=0 ps=0 
M1307 Vdd diff_66480_204480# diff_50640_203760# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M1308 diff_56880_202560# diff_42360_185400# diff_54840_203640# GND efet w=3180 l=780
+ ad=0 pd=0 as=0 ps=0 
M1309 GND diff_13200_279960# diff_16320_201240# GND efet w=3480 l=660
+ ad=0 pd=0 as=0 ps=0 
M1310 GND GND GND GND efet w=60 l=180
+ ad=0 pd=0 as=0 ps=0 
M1311 Vdd Vdd Vdd GND efet w=240 l=840
+ ad=0 pd=0 as=0 ps=0 
M1312 Vdd Vdd Vdd GND efet w=180 l=480
+ ad=0 pd=0 as=0 ps=0 
M1313 Vdd Vdd diff_16320_201240# GND efet w=840 l=3600
+ ad=0 pd=0 as=0 ps=0 
M1314 diff_48720_197520# diff_33120_151080# diff_25200_276600# GND efet w=3720 l=720
+ ad=9.7344e+06 pd=22320 as=0 ps=0 
M1315 diff_50640_203760# diff_56880_202560# GND GND efet w=5280 l=840
+ ad=0 pd=0 as=0 ps=0 
M1316 diff_56880_202560# diff_66480_204480# GND GND efet w=2820 l=780
+ ad=0 pd=0 as=0 ps=0 
M1317 diff_81360_201840# diff_80400_204480# GND GND efet w=2460 l=780
+ ad=2.6496e+06 pd=7680 as=0 ps=0 
M1318 diff_90480_215640# diff_89400_145800# diff_66480_218640# GND efet w=2280 l=780
+ ad=2.4336e+06 pd=7680 as=0 ps=0 
M1319 GND diff_88080_218880# diff_90480_215640# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1320 diff_95160_216000# diff_94080_218760# GND GND efet w=2280 l=840
+ ad=2.3472e+06 pd=7440 as=0 ps=0 
M1321 GND diff_101760_238680# diff_104280_240480# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1322 diff_108840_240120# diff_107880_238680# GND GND efet w=2340 l=780
+ ad=2.4336e+06 pd=7440 as=0 ps=0 
M1323 diff_66480_239280# diff_108240_144360# diff_108840_240120# GND efet w=2340 l=900
+ ad=0 pd=0 as=0 ps=0 
M1324 GND diff_115560_252840# diff_117960_254760# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1325 diff_122640_254280# diff_121560_252840# GND GND efet w=2280 l=840
+ ad=2.376e+06 pd=7440 as=0 ps=0 
M1326 diff_66480_253440# diff_122040_144240# diff_122640_254280# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1327 diff_117960_243960# diff_116880_145800# diff_66360_247080# GND efet w=2160 l=720
+ ad=2.6208e+06 pd=7440 as=0 ps=0 
M1328 GND diff_115560_247200# diff_117960_243960# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1329 diff_122640_244320# diff_121560_247080# GND GND efet w=2280 l=840
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1330 diff_131760_258120# diff_130680_145800# diff_66360_261120# GND efet w=2160 l=720
+ ad=2.3904e+06 pd=7440 as=0 ps=0 
M1331 GND diff_129240_261360# diff_131760_258120# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1332 diff_136320_258480# diff_135360_261120# GND GND efet w=2280 l=720
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1333 diff_54840_260160# diff_139320_149640# diff_135360_261120# GND efet w=960 l=720
+ ad=0 pd=0 as=2.6928e+06 ps=7440 
M1334 diff_143040_261360# diff_142200_145800# diff_54840_260160# GND efet w=960 l=780
+ ad=2.5776e+06 pd=7200 as=0 ps=0 
M1335 diff_66360_261120# diff_135720_144480# diff_136320_258480# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1336 diff_131760_254760# diff_130680_145800# diff_66480_253440# GND efet w=2100 l=780
+ ad=2.376e+06 pd=7440 as=0 ps=0 
M1337 diff_54840_253440# diff_125640_145800# diff_121560_252840# GND efet w=840 l=960
+ ad=0 pd=0 as=2.5056e+06 ps=7440 
M1338 diff_129240_252840# diff_128400_145800# diff_54840_253440# GND efet w=840 l=840
+ ad=2.5488e+06 pd=7680 as=0 ps=0 
M1339 diff_54840_246000# diff_125640_145800# diff_121560_247080# GND efet w=840 l=840
+ ad=0 pd=0 as=2.52e+06 ps=7440 
M1340 diff_129240_247200# diff_128400_145800# diff_54840_246000# GND efet w=840 l=720
+ ad=2.5776e+06 pd=7680 as=0 ps=0 
M1341 diff_66360_247080# diff_122040_144240# diff_122640_244320# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1342 diff_117960_240600# diff_116880_145800# diff_66480_239280# GND efet w=2100 l=720
+ ad=2.664e+06 pd=7440 as=0 ps=0 
M1343 diff_66480_239280# diff_122040_144240# diff_122640_240120# GND efet w=2160 l=960
+ ad=0 pd=0 as=2.3904e+06 ps=7440 
M1344 diff_54840_239280# diff_111840_149760# diff_107880_238680# GND efet w=840 l=720
+ ad=0 pd=0 as=2.664e+06 ps=7440 
M1345 diff_115560_238680# diff_114720_145800# diff_54840_239280# GND efet w=960 l=840
+ ad=2.5632e+06 pd=7200 as=0 ps=0 
M1346 diff_104280_229800# diff_103200_145800# diff_66480_232800# GND efet w=2160 l=720
+ ad=2.3904e+06 pd=7440 as=0 ps=0 
M1347 GND diff_101760_233040# diff_104280_229800# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1348 diff_108840_230040# diff_107880_232800# GND GND efet w=2280 l=720
+ ad=2.3904e+06 pd=7440 as=0 ps=0 
M1349 diff_54840_231960# diff_111840_149760# diff_107880_232800# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6928e+06 ps=7440 
M1350 diff_115560_233040# diff_114720_145800# diff_54840_231960# GND efet w=840 l=840
+ ad=2.592e+06 pd=7200 as=0 ps=0 
M1351 diff_66480_232800# diff_108240_144360# diff_108840_230040# GND efet w=2160 l=840
+ ad=0 pd=0 as=0 ps=0 
M1352 diff_104280_226320# diff_103200_145800# diff_66480_225120# GND efet w=2160 l=960
+ ad=2.4192e+06 pd=7440 as=0 ps=0 
M1353 diff_66480_225120# diff_108240_144360# diff_108840_225960# GND efet w=2100 l=1020
+ ad=0 pd=0 as=2.4336e+06 ps=7440 
M1354 diff_54840_225240# diff_98160_145800# diff_94080_224640# GND efet w=960 l=840
+ ad=0 pd=0 as=2.6928e+06 ps=8160 
M1355 diff_101760_224520# diff_100920_145800# diff_54840_225240# GND efet w=840 l=720
+ ad=2.736e+06 pd=7920 as=0 ps=0 
M1356 diff_54840_217800# diff_98160_145800# diff_94080_218760# GND efet w=1080 l=780
+ ad=0 pd=0 as=2.664e+06 ps=8160 
M1357 diff_101760_218880# diff_100920_145800# diff_54840_217800# GND efet w=960 l=720
+ ad=2.592e+06 pd=7680 as=0 ps=0 
M1358 diff_66480_218640# diff_94560_144240# diff_95160_216000# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1359 diff_90480_213840# diff_89400_145800# diff_66480_210960# GND efet w=2400 l=840
+ ad=2.448e+06 pd=7680 as=0 ps=0 
M1360 GND diff_88080_210480# diff_90480_213840# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1361 diff_95160_211920# diff_94080_210360# GND GND efet w=2280 l=840
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1362 diff_66480_210960# diff_94560_144240# diff_95160_211920# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1363 diff_54840_210960# diff_84360_149760# diff_80400_210360# GND efet w=960 l=780
+ ad=0 pd=0 as=2.7072e+06 ps=7440 
M1364 diff_88080_210480# diff_87240_145800# diff_54840_210960# GND efet w=840 l=720
+ ad=2.5488e+06 pd=7200 as=0 ps=0 
M1365 diff_54840_203640# diff_84360_149760# diff_80400_204480# GND efet w=900 l=900
+ ad=0 pd=0 as=2.7072e+06 ps=7680 
M1366 diff_88080_204720# diff_87240_145800# diff_54840_203640# GND efet w=900 l=780
+ ad=2.5776e+06 pd=7200 as=0 ps=0 
M1367 diff_56880_198480# diff_42360_185400# diff_54840_196800# GND efet w=3240 l=960
+ ad=8.8992e+06 pd=21600 as=3.19104e+07 ps=90720 
M1368 GND diff_56880_198480# diff_50640_196800# GND efet w=5160 l=720
+ ad=0 pd=0 as=1.63584e+07 ps=32640 
M1369 diff_66480_204480# diff_80760_144360# diff_81360_201840# GND efet w=2160 l=720
+ ad=6.43248e+07 pd=154080 as=0 ps=0 
M1370 Vdd diff_6840_159480# d3 GND efet w=61260 l=660
+ ad=0 pd=0 as=1.86926e+08 ps=302880 
M1371 GND diff_6960_191160# d3 GND efet w=114660 l=420
+ ad=0 pd=0 as=0 ps=0 
M1372 diff_48720_192480# diff_33120_151080# diff_23040_212640# GND efet w=3840 l=720
+ ad=1.00368e+07 pd=23280 as=0 ps=0 
M1373 diff_48720_197520# diff_52320_146760# diff_50640_196800# GND efet w=3720 l=720
+ ad=0 pd=0 as=0 ps=0 
M1374 diff_54840_196800# diff_42600_159120# diff_48720_197520# GND efet w=4500 l=780
+ ad=0 pd=0 as=0 ps=0 
M1375 diff_48720_192480# diff_52320_146760# diff_50640_190200# GND efet w=4080 l=720
+ ad=0 pd=0 as=1.6704e+07 ps=32880 
M1376 GND diff_66480_196680# diff_56880_198480# GND efet w=2640 l=720
+ ad=0 pd=0 as=0 ps=0 
M1377 diff_50640_196800# diff_66480_196680# Vdd GND efet w=1440 l=660
+ ad=0 pd=0 as=0 ps=0 
M1378 diff_81360_197640# diff_80400_196200# GND GND efet w=2400 l=720
+ ad=2.7072e+06 pd=7680 as=0 ps=0 
M1379 diff_66480_196680# diff_80760_144360# diff_81360_197640# GND efet w=2160 l=720
+ ad=6.17472e+07 pd=153600 as=0 ps=0 
M1380 Vdd Vdd Vdd GND efet w=600 l=360
+ ad=0 pd=0 as=0 ps=0 
M1381 GND diff_33120_151080# diff_44040_187920# GND efet w=5280 l=660
+ ad=0 pd=0 as=5.4576e+06 ps=12480 
M1382 diff_54840_189360# diff_42600_159120# diff_48720_192480# GND efet w=4620 l=780
+ ad=3.16656e+07 pd=87600 as=0 ps=0 
M1383 diff_56880_198480# Vdd Vdd GND efet w=720 l=2640
+ ad=0 pd=0 as=0 ps=0 
M1384 Vdd Vdd Vdd GND efet w=360 l=840
+ ad=0 pd=0 as=0 ps=0 
M1385 diff_56880_188280# Vdd Vdd GND efet w=780 l=2700
+ ad=9.8352e+06 pd=23280 as=0 ps=0 
M1386 diff_56880_188280# diff_42360_185400# diff_54840_189360# GND efet w=3300 l=780
+ ad=0 pd=0 as=0 ps=0 
M1387 Vdd diff_66480_190200# diff_50640_190200# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M1388 diff_44040_187920# diff_42600_159120# diff_42360_185400# GND efet w=5100 l=780
+ ad=0 pd=0 as=9.8496e+06 ps=21120 
M1389 Vdd Vdd diff_42360_185400# GND efet w=1140 l=3900
+ ad=0 pd=0 as=0 ps=0 
M1390 Vdd Vdd Vdd GND efet w=240 l=720
+ ad=0 pd=0 as=0 ps=0 
M1391 Vdd Vdd Vdd GND efet w=240 l=420
+ ad=0 pd=0 as=0 ps=0 
M1392 diff_50640_190200# diff_56880_188280# GND GND efet w=5160 l=840
+ ad=0 pd=0 as=0 ps=0 
M1393 diff_56880_188280# diff_66480_190200# GND GND efet w=2700 l=780
+ ad=0 pd=0 as=0 ps=0 
M1394 diff_81360_187680# diff_80400_190320# GND GND efet w=2280 l=720
+ ad=2.6352e+06 pd=7440 as=0 ps=0 
M1395 diff_90600_201480# diff_89400_145800# diff_66480_204480# GND efet w=2160 l=840
+ ad=2.3904e+06 pd=7440 as=0 ps=0 
M1396 GND diff_88080_204720# diff_90600_201480# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1397 diff_95160_201840# diff_94080_204480# GND GND efet w=2460 l=780
+ ad=2.376e+06 pd=7440 as=0 ps=0 
M1398 GND diff_101760_224520# diff_104280_226320# GND efet w=2460 l=900
+ ad=0 pd=0 as=0 ps=0 
M1399 diff_108840_225960# diff_107880_224520# GND GND efet w=2400 l=960
+ ad=0 pd=0 as=0 ps=0 
M1400 diff_104280_215640# diff_103200_145800# diff_66480_218640# GND efet w=2160 l=720
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1401 GND diff_101760_218880# diff_104280_215640# GND efet w=2340 l=780
+ ad=0 pd=0 as=0 ps=0 
M1402 diff_108840_216000# diff_107880_218760# GND GND efet w=2280 l=720
+ ad=2.3328e+06 pd=7200 as=0 ps=0 
M1403 GND diff_115560_238680# diff_117960_240600# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1404 diff_122640_240120# diff_121560_238680# GND GND efet w=2280 l=840
+ ad=0 pd=0 as=0 ps=0 
M1405 diff_117960_229800# diff_116880_145800# diff_66480_232800# GND efet w=2640 l=720
+ ad=2.592e+06 pd=8400 as=0 ps=0 
M1406 GND diff_115560_233040# diff_117960_229800# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1407 diff_122640_230160# diff_121560_232920# GND GND efet w=2280 l=840
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1408 GND diff_129240_252840# diff_131760_254760# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1409 diff_136320_254280# diff_135360_252840# GND GND efet w=2280 l=720
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1410 diff_66480_253440# diff_135720_144480# diff_136320_254280# GND efet w=2100 l=780
+ ad=0 pd=0 as=0 ps=0 
M1411 diff_131760_243960# diff_130680_145800# diff_66360_247080# GND efet w=2160 l=720
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1412 GND diff_129240_247200# diff_131760_243960# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1413 diff_136320_244320# diff_135360_246960# GND GND efet w=2280 l=720
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1414 diff_145440_258120# diff_144360_145800# diff_66360_261120# GND efet w=2160 l=720
+ ad=2.6352e+06 pd=7440 as=0 ps=0 
M1415 GND diff_143040_261360# diff_145440_258120# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1416 diff_150120_258480# diff_149040_261240# GND GND efet w=2280 l=840
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1417 diff_54840_260160# diff_153120_145800# diff_149040_261240# GND efet w=1020 l=840
+ ad=0 pd=0 as=2.5776e+06 ps=7680 
M1418 diff_156720_261360# diff_155880_145800# diff_54840_260160# GND efet w=900 l=780
+ ad=2.6784e+06 pd=7440 as=0 ps=0 
M1419 diff_66360_261120# diff_149520_144360# diff_150120_258480# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1420 diff_145440_254760# diff_144360_145800# diff_66480_253440# GND efet w=2100 l=780
+ ad=2.6208e+06 pd=7440 as=0 ps=0 
M1421 diff_54840_253440# diff_139320_149640# diff_135360_252840# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6208e+06 ps=7440 
M1422 diff_143040_252840# diff_142200_145800# diff_54840_253440# GND efet w=840 l=840
+ ad=2.5488e+06 pd=7440 as=0 ps=0 
M1423 diff_54840_246000# diff_139320_149640# diff_135360_246960# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6352e+06 ps=7440 
M1424 diff_143040_247200# diff_142200_145800# diff_54840_246000# GND efet w=840 l=840
+ ad=2.5488e+06 pd=7200 as=0 ps=0 
M1425 diff_66360_247080# diff_135720_144480# diff_136320_244320# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1426 diff_131760_240600# diff_130680_145800# diff_66480_239280# GND efet w=2160 l=720
+ ad=2.4336e+06 pd=7440 as=0 ps=0 
M1427 diff_54840_239280# diff_125640_145800# diff_121560_238680# GND efet w=840 l=840
+ ad=0 pd=0 as=2.5632e+06 ps=7680 
M1428 diff_129240_238680# diff_128400_145800# diff_54840_239280# GND efet w=840 l=720
+ ad=2.592e+06 pd=7680 as=0 ps=0 
M1429 diff_54840_231960# diff_125640_145800# diff_121560_232920# GND efet w=840 l=840
+ ad=0 pd=0 as=2.6064e+06 ps=7680 
M1430 diff_129240_233040# diff_128400_145800# diff_54840_231960# GND efet w=840 l=720
+ ad=2.5776e+06 pd=7680 as=0 ps=0 
M1431 diff_66480_232800# diff_122040_144240# diff_122640_230160# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1432 diff_117960_226800# diff_116880_145800# diff_66480_225120# GND efet w=2280 l=840
+ ad=2.592e+06 pd=7680 as=0 ps=0 
M1433 GND diff_115560_224520# diff_117960_226800# GND efet w=2340 l=780
+ ad=0 pd=0 as=0 ps=0 
M1434 diff_122640_225960# diff_121560_224640# GND GND efet w=2400 l=840
+ ad=2.3472e+06 pd=7440 as=0 ps=0 
M1435 diff_66480_225120# diff_122040_144240# diff_122640_225960# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M1436 diff_54840_225240# diff_111840_149760# diff_107880_224520# GND efet w=840 l=720
+ ad=0 pd=0 as=2.7072e+06 ps=7680 
M1437 diff_115560_224520# diff_114720_145800# diff_54840_225240# GND efet w=960 l=780
+ ad=2.5488e+06 pd=7200 as=0 ps=0 
M1438 diff_54840_217800# diff_111840_149760# diff_107880_218760# GND efet w=960 l=720
+ ad=0 pd=0 as=2.7504e+06 ps=7680 
M1439 diff_115560_218880# diff_114720_145800# diff_54840_217800# GND efet w=960 l=720
+ ad=2.4336e+06 pd=6960 as=0 ps=0 
M1440 diff_66480_218640# diff_108240_144360# diff_108840_216000# GND efet w=2160 l=840
+ ad=0 pd=0 as=0 ps=0 
M1441 diff_104280_212280# diff_103200_145800# diff_66480_210960# GND efet w=2160 l=720
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1442 diff_54840_210960# diff_98160_145800# diff_94080_210360# GND efet w=1020 l=720
+ ad=0 pd=0 as=2.6928e+06 ps=8160 
M1443 diff_101760_210360# diff_100920_145800# diff_54840_210960# GND efet w=840 l=720
+ ad=2.5632e+06 pd=7680 as=0 ps=0 
M1444 diff_54840_203640# diff_98160_145800# diff_94080_204480# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6784e+06 ps=7440 
M1445 diff_101760_204840# diff_100920_145800# diff_54840_203640# GND efet w=840 l=720
+ ad=2.52e+06 pd=7440 as=0 ps=0 
M1446 diff_66480_204480# diff_94560_144240# diff_95160_201840# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1447 diff_90600_197760# diff_89400_145800# diff_66480_196680# GND efet w=2220 l=900
+ ad=2.448e+06 pd=7440 as=0 ps=0 
M1448 diff_54840_196800# diff_84360_149760# diff_80400_196200# GND efet w=1260 l=1560
+ ad=0 pd=0 as=2.6352e+06 ps=7440 
M1449 diff_88080_196200# diff_87240_145800# diff_54840_196800# GND efet w=840 l=720
+ ad=2.6496e+06 pd=7440 as=0 ps=0 
M1450 diff_54840_189360# diff_84360_149760# diff_80400_190320# GND efet w=840 l=840
+ ad=0 pd=0 as=2.6496e+06 ps=7440 
M1451 diff_88080_190440# diff_87240_145800# diff_54840_189360# GND efet w=840 l=720
+ ad=2.5632e+06 pd=7200 as=0 ps=0 
M1452 diff_66480_190200# diff_80760_144360# diff_81360_187680# GND efet w=2040 l=720
+ ad=6.3432e+07 pd=152880 as=0 ps=0 
M1453 diff_56880_184320# diff_42360_185400# diff_54840_182640# GND efet w=3180 l=720
+ ad=9.6912e+06 pd=23280 as=3.12192e+07 ps=86880 
M1454 GND diff_56880_184320# diff_50640_182520# GND efet w=5160 l=840
+ ad=0 pd=0 as=1.6848e+07 ps=32400 
M1455 GND diff_66480_182520# diff_56880_184320# GND efet w=2760 l=720
+ ad=0 pd=0 as=0 ps=0 
M1456 diff_48720_180120# diff_33120_151080# diff_23160_135720# GND efet w=3900 l=780
+ ad=1.01088e+07 pd=23040 as=0 ps=0 
M1457 diff_48720_180120# diff_52320_146760# diff_50640_182520# GND efet w=3840 l=720
+ ad=0 pd=0 as=0 ps=0 
M1458 diff_54840_182640# diff_42600_159120# diff_48720_180120# GND efet w=4500 l=780
+ ad=0 pd=0 as=0 ps=0 
M1459 diff_50640_182520# diff_66480_182520# Vdd GND efet w=1380 l=780
+ ad=0 pd=0 as=0 ps=0 
M1460 diff_81360_183480# diff_80400_181920# GND GND efet w=2280 l=720
+ ad=2.6064e+06 pd=7440 as=0 ps=0 
M1461 diff_66480_182520# diff_80760_144360# diff_81360_183480# GND efet w=2160 l=720
+ ad=6.44112e+07 pd=153840 as=0 ps=0 
M1462 diff_56880_184320# Vdd Vdd GND efet w=660 l=2760
+ ad=0 pd=0 as=0 ps=0 
M1463 diff_6840_159480# diff_8880_168480# GND GND efet w=21840 l=720
+ ad=4.01904e+07 pd=79680 as=0 ps=0 
M1464 diff_48720_174000# diff_43680_161280# diff_34920_109680# GND efet w=3720 l=720
+ ad=1.15344e+07 pd=25920 as=0 ps=0 
M1465 diff_48720_174000# diff_52320_146760# diff_50640_174720# GND efet w=3960 l=720
+ ad=0 pd=0 as=1.7064e+07 ps=33600 
M1466 Vdd Vdd Vdd GND efet w=660 l=420
+ ad=0 pd=0 as=0 ps=0 
M1467 diff_54840_175200# diff_42600_159120# diff_48720_174000# GND efet w=4500 l=780
+ ad=3.15936e+07 pd=85920 as=0 ps=0 
M1468 Vdd Vdd Vdd GND efet w=360 l=840
+ ad=0 pd=0 as=0 ps=0 
M1469 diff_56880_174120# Vdd Vdd GND efet w=600 l=2640
+ ad=8.8272e+06 pd=21600 as=0 ps=0 
M1470 Vdd diff_66480_176040# diff_50640_174720# GND efet w=1380 l=720
+ ad=0 pd=0 as=0 ps=0 
M1471 diff_8880_168480# diff_8880_168480# diff_8880_168480# GND efet w=240 l=480
+ ad=1.1808e+07 pd=21600 as=0 ps=0 
M1472 diff_8880_168480# diff_8880_168480# diff_8880_168480# GND efet w=360 l=480
+ ad=0 pd=0 as=0 ps=0 
M1473 diff_23160_135720# diff_22200_108240# diff_8880_168480# GND efet w=2760 l=720
+ ad=0 pd=0 as=0 ps=0 
M1474 diff_48720_169080# diff_43680_161280# diff_25200_276600# GND efet w=3720 l=720
+ ad=9.7056e+06 pd=22800 as=0 ps=0 
M1475 diff_56880_174120# diff_42360_157080# diff_54840_175200# GND efet w=3120 l=720
+ ad=0 pd=0 as=0 ps=0 
M1476 diff_56880_170160# diff_42360_157080# diff_54840_168480# GND efet w=3180 l=780
+ ad=8.7408e+06 pd=21600 as=3.1608e+07 ps=86640 
M1477 diff_50640_174720# diff_56880_174120# GND GND efet w=5040 l=720
+ ad=0 pd=0 as=0 ps=0 
M1478 diff_56880_174120# diff_66480_176040# GND GND efet w=2640 l=720
+ ad=0 pd=0 as=0 ps=0 
M1479 GND diff_56880_170160# diff_50640_168360# GND efet w=5160 l=720
+ ad=0 pd=0 as=1.6416e+07 ps=32400 
M1480 diff_81360_173400# diff_80400_176040# GND GND efet w=2580 l=780
+ ad=2.6784e+06 pd=7920 as=0 ps=0 
M1481 GND diff_88080_196200# diff_90600_197760# GND efet w=2340 l=780
+ ad=0 pd=0 as=0 ps=0 
M1482 diff_95160_197640# diff_94080_196200# GND GND efet w=2640 l=720
+ ad=2.4336e+06 pd=7440 as=0 ps=0 
M1483 diff_66480_196680# diff_94560_144240# diff_95160_197640# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1484 diff_90600_187200# diff_89400_145800# diff_66480_190200# GND efet w=2220 l=900
+ ad=2.4768e+06 pd=7440 as=0 ps=0 
M1485 GND diff_88080_190440# diff_90600_187200# GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M1486 diff_95160_187560# diff_94080_190320# GND GND efet w=2580 l=780
+ ad=2.4048e+06 pd=7440 as=0 ps=0 
M1487 GND diff_101760_210360# diff_104280_212280# GND efet w=2280 l=780
+ ad=0 pd=0 as=0 ps=0 
M1488 diff_108840_211920# diff_107880_210360# GND GND efet w=2280 l=720
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1489 diff_66480_210960# diff_108240_144360# diff_108840_211920# GND efet w=2160 l=840
+ ad=0 pd=0 as=0 ps=0 
M1490 diff_118080_215640# diff_116880_145800# diff_66480_218640# GND efet w=2160 l=840
+ ad=2.376e+06 pd=7200 as=0 ps=0 
M1491 GND diff_115560_218880# diff_118080_215640# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1492 diff_122640_216000# diff_121560_218760# GND GND efet w=2280 l=840
+ ad=2.3472e+06 pd=7440 as=0 ps=0 
M1493 diff_66480_239280# diff_135720_144480# diff_136320_240120# GND efet w=2160 l=960
+ ad=0 pd=0 as=2.3904e+06 ps=7440 
M1494 GND diff_129240_238680# diff_131760_240600# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1495 diff_136320_240120# diff_135360_238680# GND GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1496 diff_131760_229800# diff_130680_145800# diff_66480_232800# GND efet w=2160 l=720
+ ad=2.376e+06 pd=7440 as=0 ps=0 
M1497 GND diff_129240_233040# diff_131760_229800# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1498 diff_136320_230160# diff_135360_232800# GND GND efet w=2280 l=720
+ ad=2.3328e+06 pd=7200 as=0 ps=0 
M1499 GND diff_143040_252840# diff_145440_254760# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1500 diff_150120_254280# diff_149040_252840# GND GND efet w=2280 l=840
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1501 diff_66480_253440# diff_149520_144360# diff_150120_254280# GND efet w=2100 l=780
+ ad=0 pd=0 as=0 ps=0 
M1502 diff_145440_243960# diff_144360_145800# diff_66360_247080# GND efet w=2160 l=720
+ ad=2.6064e+06 pd=7440 as=0 ps=0 
M1503 GND diff_143040_247200# diff_145440_243960# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1504 diff_150120_244320# diff_149040_247080# GND GND efet w=2280 l=840
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1505 diff_159240_258120# diff_158160_145800# diff_66360_261120# GND efet w=2160 l=720
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1506 GND diff_156720_261360# diff_159240_258120# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1507 diff_163800_258480# diff_162840_261120# GND GND efet w=2280 l=720
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1508 diff_54840_260160# diff_166800_149760# diff_162840_261120# GND efet w=900 l=780
+ ad=0 pd=0 as=2.5632e+06 ps=7680 
M1509 diff_170520_261360# diff_169680_145800# diff_54840_260160# GND efet w=900 l=780
+ ad=2.5488e+06 pd=7440 as=0 ps=0 
M1510 diff_66360_261120# diff_163320_144240# diff_163800_258480# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1511 diff_159240_254760# diff_158160_145800# diff_66480_253440# GND efet w=2100 l=780
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1512 diff_54840_253440# diff_153120_145800# diff_149040_252840# GND efet w=840 l=840
+ ad=0 pd=0 as=2.52e+06 ps=7200 
M1513 diff_156720_252840# diff_155880_145800# diff_54840_253440# GND efet w=840 l=720
+ ad=2.6496e+06 pd=7440 as=0 ps=0 
M1514 diff_54840_246000# diff_153120_145800# diff_149040_247080# GND efet w=840 l=840
+ ad=0 pd=0 as=2.4768e+06 ps=7680 
M1515 diff_156720_247200# diff_155880_145800# diff_54840_246000# GND efet w=840 l=720
+ ad=2.5344e+06 pd=7440 as=0 ps=0 
M1516 diff_66360_247080# diff_149520_144360# diff_150120_244320# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1517 diff_145440_240600# diff_144360_145800# diff_66480_239280# GND efet w=2040 l=720
+ ad=2.6064e+06 pd=7440 as=0 ps=0 
M1518 diff_54840_239280# diff_139320_149640# diff_135360_238680# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6352e+06 ps=7440 
M1519 diff_143040_238680# diff_142200_145800# diff_54840_239280# GND efet w=840 l=840
+ ad=2.5344e+06 pd=7200 as=0 ps=0 
M1520 diff_54840_231960# diff_139320_149640# diff_135360_232800# GND efet w=840 l=720
+ ad=0 pd=0 as=2.664e+06 ps=7440 
M1521 diff_143040_233040# diff_142200_145800# diff_54840_231960# GND efet w=840 l=840
+ ad=2.5488e+06 pd=7440 as=0 ps=0 
M1522 diff_66480_232800# diff_135720_144480# diff_136320_230160# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1523 diff_131760_226440# diff_130680_145800# diff_66480_225120# GND efet w=2040 l=720
+ ad=2.376e+06 pd=7440 as=0 ps=0 
M1524 diff_54840_225240# diff_125640_145800# diff_121560_224640# GND efet w=840 l=840
+ ad=0 pd=0 as=2.5488e+06 ps=7680 
M1525 diff_129240_224520# diff_128400_145800# diff_54840_225240# GND efet w=840 l=720
+ ad=2.5488e+06 pd=7680 as=0 ps=0 
M1526 diff_54840_217800# diff_125640_145800# diff_121560_218760# GND efet w=840 l=840
+ ad=0 pd=0 as=2.5776e+06 ps=7680 
M1527 diff_129240_218880# diff_128400_145800# diff_54840_217800# GND efet w=840 l=720
+ ad=2.6064e+06 pd=7680 as=0 ps=0 
M1528 diff_66480_218640# diff_122040_144240# diff_122640_216000# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1529 diff_118080_212040# diff_116880_145800# diff_66480_210960# GND efet w=2160 l=840
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1530 diff_54840_210960# diff_111840_149760# diff_107880_210360# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6496e+06 ps=7440 
M1531 diff_115560_210360# diff_114720_145800# diff_54840_210960# GND efet w=840 l=720
+ ad=2.5632e+06 pd=7200 as=0 ps=0 
M1532 diff_104280_201480# diff_103200_145800# diff_66480_204480# GND efet w=2160 l=720
+ ad=2.3904e+06 pd=7440 as=0 ps=0 
M1533 GND diff_101760_204840# diff_104280_201480# GND efet w=2280 l=840
+ ad=0 pd=0 as=0 ps=0 
M1534 diff_108840_201840# diff_107880_204480# GND GND efet w=2280 l=720
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1535 diff_54840_203640# diff_111840_149760# diff_107880_204480# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6784e+06 ps=7440 
M1536 diff_115560_204840# diff_114720_145800# diff_54840_203640# GND efet w=840 l=720
+ ad=2.5632e+06 pd=7200 as=0 ps=0 
M1537 diff_66480_204480# diff_108240_144360# diff_108840_201840# GND efet w=2160 l=840
+ ad=0 pd=0 as=0 ps=0 
M1538 diff_104280_198120# diff_103200_145800# diff_66480_196680# GND efet w=2220 l=780
+ ad=2.4336e+06 pd=7440 as=0 ps=0 
M1539 diff_66480_196680# diff_108240_144360# diff_108840_197640# GND efet w=2220 l=900
+ ad=0 pd=0 as=2.448e+06 ps=7680 
M1540 GND diff_101760_196200# diff_104280_198120# GND efet w=2340 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1541 diff_54840_196800# diff_98160_145800# diff_94080_196200# GND efet w=840 l=720
+ ad=0 pd=0 as=2.808e+06 ps=7920 
M1542 diff_101760_196200# diff_100920_145800# diff_54840_196800# GND efet w=840 l=720
+ ad=2.6208e+06 pd=7920 as=0 ps=0 
M1543 diff_54840_189360# diff_98160_145800# diff_94080_190320# GND efet w=900 l=780
+ ad=0 pd=0 as=2.7072e+06 ps=8160 
M1544 diff_101760_190560# diff_100920_145800# diff_54840_189360# GND efet w=840 l=720
+ ad=2.5488e+06 pd=7680 as=0 ps=0 
M1545 diff_66480_190200# diff_94560_144240# diff_95160_187560# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1546 diff_90600_183600# diff_89400_145800# diff_66480_182520# GND efet w=2160 l=840
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1547 diff_54840_182640# diff_84360_149760# diff_80400_181920# GND efet w=840 l=840
+ ad=0 pd=0 as=2.6928e+06 ps=7680 
M1548 diff_88080_182040# diff_87240_145800# diff_54840_182640# GND efet w=840 l=720
+ ad=2.6064e+06 pd=7440 as=0 ps=0 
M1549 GND diff_88080_182040# diff_90600_183600# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1550 diff_95160_183480# diff_94080_181920# GND GND efet w=2280 l=720
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1551 diff_66480_182520# diff_94560_144240# diff_95160_183480# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1552 diff_54840_175200# diff_84360_149760# diff_80400_176040# GND efet w=840 l=840
+ ad=0 pd=0 as=2.664e+06 ps=7440 
M1553 diff_88080_176280# diff_87240_145800# diff_54840_175200# GND efet w=840 l=720
+ ad=2.5776e+06 pd=7200 as=0 ps=0 
M1554 diff_66480_176040# diff_80760_144360# diff_81360_173400# GND efet w=2160 l=720
+ ad=6.40512e+07 pd=153840 as=0 ps=0 
M1555 diff_48720_169080# diff_52320_146760# diff_50640_168360# GND efet w=3900 l=780
+ ad=0 pd=0 as=0 ps=0 
M1556 diff_6840_159480# diff_8760_228840# GND GND efet w=21840 l=720
+ ad=0 pd=0 as=0 ps=0 
M1557 Vdd diff_16200_162120# diff_6840_159480# GND efet w=1080 l=780
+ ad=0 pd=0 as=0 ps=0 
M1558 diff_6840_159480# diff_16200_162120# diff_6840_159480# GND efet w=4980 l=1680
+ ad=0 pd=0 as=0 ps=0 
M1559 diff_16200_162120# diff_16200_162120# diff_16200_162120# GND efet w=240 l=840
+ ad=2.2896e+06 pd=8160 as=0 ps=0 
M1560 Vdd Vdd diff_16200_162120# GND efet w=840 l=720
+ ad=0 pd=0 as=0 ps=0 
M1561 diff_16200_162120# diff_16200_162120# diff_16200_162120# GND efet w=360 l=420
+ ad=0 pd=0 as=0 ps=0 
M1562 diff_6960_191160# diff_6840_159480# GND GND efet w=7920 l=600
+ ad=3.12624e+07 pd=60720 as=0 ps=0 
M1563 diff_6960_191160# diff_8760_228840# GND GND efet w=21480 l=780
+ ad=0 pd=0 as=0 ps=0 
M1564 diff_6960_191160# diff_16200_152040# diff_6960_191160# GND efet w=3900 l=1860
+ ad=0 pd=0 as=0 ps=0 
M1565 Vdd diff_16200_152040# diff_6960_191160# GND efet w=1080 l=840
+ ad=0 pd=0 as=0 ps=0 
M1566 diff_16200_152040# diff_16200_152040# diff_16200_152040# GND efet w=240 l=960
+ ad=2.1168e+06 pd=6960 as=0 ps=0 
M1567 Vdd Vdd diff_16200_152040# GND efet w=840 l=840
+ ad=0 pd=0 as=0 ps=0 
M1568 diff_16200_152040# diff_16200_152040# diff_16200_152040# GND efet w=60 l=300
+ ad=0 pd=0 as=0 ps=0 
M1569 diff_48720_164160# diff_43680_161280# diff_23040_212640# GND efet w=3720 l=720
+ ad=9.4176e+06 pd=22560 as=0 ps=0 
M1570 diff_54840_168480# diff_42600_159120# diff_48720_169080# GND efet w=4560 l=840
+ ad=0 pd=0 as=0 ps=0 
M1571 GND diff_43680_161280# diff_44040_159600# GND efet w=5280 l=660
+ ad=0 pd=0 as=5.5584e+06 ps=12480 
M1572 diff_48720_164160# diff_52320_146760# diff_50640_161880# GND efet w=3840 l=840
+ ad=0 pd=0 as=1.67328e+07 ps=32640 
M1573 diff_54840_161040# diff_42600_159120# diff_48720_164160# GND efet w=4500 l=780
+ ad=3.07728e+07 pd=86160 as=0 ps=0 
M1574 GND diff_66480_168360# diff_56880_170160# GND efet w=2820 l=780
+ ad=0 pd=0 as=0 ps=0 
M1575 diff_50640_168360# diff_66480_168360# Vdd GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M1576 diff_81360_169200# diff_80400_167760# GND GND efet w=2520 l=720
+ ad=2.664e+06 pd=7920 as=0 ps=0 
M1577 diff_66480_168360# diff_80760_144360# diff_81360_169200# GND efet w=2160 l=720
+ ad=6.16752e+07 pd=155520 as=0 ps=0 
M1578 diff_56880_170160# Vdd Vdd GND efet w=600 l=2640
+ ad=0 pd=0 as=0 ps=0 
M1579 Vdd Vdd Vdd GND efet w=600 l=360
+ ad=0 pd=0 as=0 ps=0 
M1580 Vdd Vdd Vdd GND efet w=360 l=840
+ ad=0 pd=0 as=0 ps=0 
M1581 diff_56880_159960# Vdd Vdd GND efet w=720 l=2760
+ ad=9.2736e+06 pd=22800 as=0 ps=0 
M1582 diff_56880_159960# diff_42360_157080# diff_54840_161040# GND efet w=3420 l=900
+ ad=0 pd=0 as=0 ps=0 
M1583 diff_44040_159600# diff_42600_159120# diff_42360_157080# GND efet w=4680 l=720
+ ad=0 pd=0 as=1.0008e+07 ps=20400 
M1584 Vdd Vdd diff_42360_157080# GND efet w=1200 l=3960
+ ad=0 pd=0 as=0 ps=0 
M1585 Vdd Vdd Vdd GND efet w=180 l=540
+ ad=0 pd=0 as=0 ps=0 
M1586 Vdd Vdd Vdd GND efet w=120 l=120
+ ad=0 pd=0 as=0 ps=0 
M1587 Vdd Vdd Vdd GND efet w=300 l=420
+ ad=0 pd=0 as=0 ps=0 
M1588 Vdd diff_66480_162000# diff_50640_161880# GND efet w=1380 l=780
+ ad=0 pd=0 as=0 ps=0 
M1589 diff_50640_161880# diff_56880_159960# GND GND efet w=5160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1590 diff_56880_159960# diff_66480_162000# GND GND efet w=2640 l=840
+ ad=0 pd=0 as=0 ps=0 
M1591 diff_56880_156000# diff_42360_157080# diff_54840_154320# GND efet w=3240 l=720
+ ad=9.648e+06 pd=23040 as=3.14496e+07 ps=86160 
M1592 diff_81360_159720# diff_80400_162000# GND GND efet w=2520 l=780
+ ad=2.3616e+06 pd=7680 as=0 ps=0 
M1593 GND diff_88080_176280# diff_90600_173040# GND efet w=2340 l=780
+ ad=0 pd=0 as=2.376e+06 ps=7440 
M1594 diff_95160_173400# diff_94080_176160# GND GND efet w=2580 l=780
+ ad=2.4336e+06 pd=7440 as=0 ps=0 
M1595 diff_90600_173040# diff_89400_145800# diff_66480_176040# GND efet w=2340 l=900
+ ad=0 pd=0 as=0 ps=0 
M1596 diff_108840_197640# diff_107880_196080# GND GND efet w=2280 l=840
+ ad=0 pd=0 as=0 ps=0 
M1597 GND diff_115560_210360# diff_118080_212040# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1598 diff_122640_211920# diff_121560_210360# GND GND efet w=2280 l=780
+ ad=2.3328e+06 pd=7200 as=0 ps=0 
M1599 diff_66480_210960# diff_122040_144240# diff_122640_211920# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1600 diff_118080_201480# diff_116880_145800# diff_66480_204480# GND efet w=2160 l=840
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1601 GND diff_115560_204840# diff_118080_201480# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1602 diff_122640_201840# diff_121560_204480# GND GND efet w=2580 l=780
+ ad=2.3616e+06 pd=7440 as=0 ps=0 
M1603 GND diff_129240_224520# diff_131760_226440# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1604 diff_136320_225960# diff_135360_224520# GND GND efet w=2280 l=720
+ ad=2.376e+06 pd=7200 as=0 ps=0 
M1605 diff_66480_225120# diff_135720_144480# diff_136320_225960# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M1606 GND diff_143040_238680# diff_145440_240600# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1607 diff_150000_242040# diff_149040_238680# GND GND efet w=2400 l=780
+ ad=2.3328e+06 pd=7680 as=0 ps=0 
M1608 diff_66480_239280# diff_149520_144360# diff_150000_242040# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M1609 diff_145440_229800# diff_144360_145800# diff_66480_232800# GND efet w=2160 l=720
+ ad=2.592e+06 pd=7440 as=0 ps=0 
M1610 GND diff_143040_233040# diff_145440_229800# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1611 diff_150120_230160# diff_149040_232920# GND GND efet w=2280 l=840
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1612 GND diff_156720_252840# diff_159240_254760# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1613 diff_163800_254280# diff_162840_252840# GND GND efet w=2280 l=720
+ ad=2.376e+06 pd=7440 as=0 ps=0 
M1614 diff_66480_253440# diff_163320_144240# diff_163800_254280# GND efet w=2100 l=780
+ ad=0 pd=0 as=0 ps=0 
M1615 diff_159240_243960# diff_158160_145800# diff_66360_247080# GND efet w=2160 l=720
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1616 GND diff_156720_247200# diff_159240_243960# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1617 diff_163800_244320# diff_162840_247080# GND GND efet w=2280 l=720
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1618 diff_172920_258840# diff_171960_145800# diff_66360_261120# GND efet w=2580 l=780
+ ad=2.4768e+06 pd=8400 as=0 ps=0 
M1619 GND diff_170520_261360# diff_172920_258840# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1620 diff_177600_258480# diff_176520_261240# GND GND efet w=2280 l=720
+ ad=2.376e+06 pd=7440 as=0 ps=0 
M1621 diff_54840_260160# diff_180600_149640# diff_176520_261240# GND efet w=960 l=720
+ ad=0 pd=0 as=2.664e+06 ps=7680 
M1622 diff_184200_262200# diff_183480_145800# diff_54840_260160# GND efet w=1020 l=780
+ ad=2.592e+06 pd=7920 as=0 ps=0 
M1623 diff_66360_261120# diff_177000_144360# diff_177600_258480# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1624 diff_172920_254760# diff_171960_145800# diff_66480_253440# GND efet w=2520 l=780
+ ad=2.5776e+06 pd=8400 as=0 ps=0 
M1625 diff_54840_253440# diff_166800_149760# diff_162840_252840# GND efet w=840 l=720
+ ad=0 pd=0 as=2.5056e+06 ps=7440 
M1626 diff_170520_252840# diff_169680_145800# diff_54840_253440# GND efet w=840 l=720
+ ad=2.5488e+06 pd=7680 as=0 ps=0 
M1627 diff_54840_246000# diff_166800_149760# diff_162840_247080# GND efet w=840 l=720
+ ad=0 pd=0 as=2.52e+06 ps=7680 
M1628 diff_170520_247200# diff_169680_145800# diff_54840_246000# GND efet w=840 l=720
+ ad=2.5056e+06 pd=7440 as=0 ps=0 
M1629 diff_66360_247080# diff_163320_144240# diff_163800_244320# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1630 diff_159240_240600# diff_158160_145800# diff_66480_239280# GND efet w=2040 l=780
+ ad=2.4048e+06 pd=7440 as=0 ps=0 
M1631 diff_54840_239280# diff_153120_145800# diff_149040_238680# GND efet w=840 l=780
+ ad=0 pd=0 as=2.5488e+06 ps=7200 
M1632 diff_156720_238680# diff_155880_145800# diff_54840_239280# GND efet w=840 l=720
+ ad=2.6496e+06 pd=7440 as=0 ps=0 
M1633 diff_54840_231960# diff_153120_145800# diff_149040_232920# GND efet w=840 l=840
+ ad=0 pd=0 as=2.592e+06 ps=7440 
M1634 diff_156720_233040# diff_155880_145800# diff_54840_231960# GND efet w=840 l=720
+ ad=2.6064e+06 pd=7680 as=0 ps=0 
M1635 diff_66480_232800# diff_149520_144360# diff_150120_230160# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1636 diff_145440_226440# diff_144360_145800# diff_66480_225120# GND efet w=2040 l=720
+ ad=2.6208e+06 pd=7440 as=0 ps=0 
M1637 diff_54840_225240# diff_139320_149640# diff_135360_224520# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6496e+06 ps=7680 
M1638 diff_143040_224520# diff_142200_145800# diff_54840_225240# GND efet w=840 l=840
+ ad=2.52e+06 pd=7200 as=0 ps=0 
M1639 diff_131760_215640# diff_130680_145800# diff_66480_218640# GND efet w=2160 l=720
+ ad=2.3616e+06 pd=7440 as=0 ps=0 
M1640 GND diff_129240_218880# diff_131760_215640# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1641 diff_136320_216000# diff_135360_218760# GND GND efet w=2280 l=720
+ ad=2.3328e+06 pd=7200 as=0 ps=0 
M1642 diff_54840_217800# diff_139320_149640# diff_135360_218760# GND efet w=840 l=720
+ ad=0 pd=0 as=2.592e+06 ps=7920 
M1643 diff_143040_218880# diff_142200_145800# diff_54840_217800# GND efet w=840 l=840
+ ad=2.5632e+06 pd=7200 as=0 ps=0 
M1644 diff_66480_218640# diff_135720_144480# diff_136320_216000# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1645 diff_131760_212280# diff_130680_145800# diff_66480_210960# GND efet w=2160 l=720
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1646 diff_129240_210480# diff_128400_145800# diff_54840_210960# GND efet w=1080 l=1260
+ ad=2.592e+06 pd=8400 as=0 ps=0 
M1647 diff_54840_210960# diff_125640_145800# diff_121560_210360# GND efet w=840 l=840
+ ad=0 pd=0 as=2.592e+06 ps=7680 
M1648 diff_54840_203640# diff_125640_145800# diff_121560_204480# GND efet w=840 l=720
+ ad=0 pd=0 as=2.7072e+06 ps=7920 
M1649 diff_129240_204720# diff_128400_145800# diff_54840_203640# GND efet w=840 l=720
+ ad=2.5776e+06 pd=7440 as=0 ps=0 
M1650 diff_66480_204480# diff_122040_144240# diff_122640_201840# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1651 diff_118080_198000# diff_116880_145800# diff_66480_196680# GND efet w=2160 l=960
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1652 diff_66480_196680# diff_122040_144240# diff_122640_197640# GND efet w=2100 l=900
+ ad=0 pd=0 as=2.3616e+06 ps=7440 
M1653 diff_54840_196800# diff_111840_149760# diff_107880_196080# GND efet w=840 l=720
+ ad=0 pd=0 as=2.7648e+06 ps=7680 
M1654 diff_115560_196200# diff_114720_145800# diff_54840_196800# GND efet w=840 l=720
+ ad=2.6496e+06 pd=7440 as=0 ps=0 
M1655 diff_104280_187200# diff_103200_145800# diff_66480_190200# GND efet w=2160 l=720
+ ad=2.4624e+06 pd=7440 as=0 ps=0 
M1656 GND diff_101760_190560# diff_104280_187200# GND efet w=2400 l=840
+ ad=0 pd=0 as=0 ps=0 
M1657 diff_108840_187560# diff_107880_190320# GND GND efet w=2400 l=720
+ ad=2.4624e+06 pd=7680 as=0 ps=0 
M1658 diff_54840_189360# diff_111840_149760# diff_107880_190320# GND efet w=900 l=720
+ ad=0 pd=0 as=2.6928e+06 ps=7680 
M1659 diff_115560_190440# diff_114720_145800# diff_54840_189360# GND efet w=840 l=720
+ ad=2.5632e+06 pd=7200 as=0 ps=0 
M1660 diff_66480_190200# diff_108240_144360# diff_108840_187560# GND efet w=2280 l=840
+ ad=0 pd=0 as=0 ps=0 
M1661 diff_104280_183840# diff_103200_145800# diff_66480_182520# GND efet w=2160 l=720
+ ad=2.376e+06 pd=7200 as=0 ps=0 
M1662 diff_54840_182640# diff_98160_145800# diff_94080_181920# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6928e+06 ps=8160 
M1663 diff_101760_182040# diff_100920_145800# diff_54840_182640# GND efet w=840 l=720
+ ad=2.5632e+06 pd=7920 as=0 ps=0 
M1664 diff_54840_175200# diff_98160_145800# diff_94080_176160# GND efet w=840 l=720
+ ad=0 pd=0 as=2.7072e+06 ps=7920 
M1665 diff_101760_176400# diff_100920_145800# diff_54840_175200# GND efet w=840 l=720
+ ad=2.6496e+06 pd=7440 as=0 ps=0 
M1666 diff_66480_176040# diff_94560_144240# diff_95160_173400# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1667 diff_90600_169320# diff_89400_145800# diff_66480_168360# GND efet w=2280 l=1020
+ ad=2.4192e+06 pd=7200 as=0 ps=0 
M1668 diff_54840_168480# diff_84360_149760# diff_80400_167760# GND efet w=840 l=840
+ ad=0 pd=0 as=2.6496e+06 ps=7440 
M1669 diff_88080_167760# diff_87240_145800# diff_54840_168480# GND efet w=840 l=720
+ ad=2.5488e+06 pd=7200 as=0 ps=0 
M1670 GND diff_88080_167760# diff_90600_169320# GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M1671 diff_95160_169200# diff_94080_167760# GND GND efet w=2580 l=780
+ ad=2.4336e+06 pd=7440 as=0 ps=0 
M1672 diff_66480_168360# diff_94560_144240# diff_95160_169200# GND efet w=2220 l=780
+ ad=0 pd=0 as=0 ps=0 
M1673 diff_54840_161040# diff_84360_149760# diff_80400_162000# GND efet w=840 l=840
+ ad=0 pd=0 as=2.6496e+06 ps=7440 
M1674 diff_88080_162120# diff_87240_145800# diff_54840_161040# GND efet w=840 l=720
+ ad=2.5776e+06 pd=7200 as=0 ps=0 
M1675 diff_66480_162000# diff_80760_144360# diff_81360_159720# GND efet w=2160 l=720
+ ad=6.21648e+07 pd=152880 as=0 ps=0 
M1676 GND diff_56880_156000# diff_50640_154200# GND efet w=5160 l=720
+ ad=0 pd=0 as=1.71792e+07 ps=32640 
M1677 diff_48720_152160# diff_43680_161280# diff_23160_135720# GND efet w=4020 l=900
+ ad=9.288e+06 pd=22800 as=0 ps=0 
M1678 diff_48720_152160# diff_52320_146760# diff_50640_154200# GND efet w=3720 l=840
+ ad=0 pd=0 as=0 ps=0 
M1679 diff_54840_154320# diff_42600_159120# diff_48720_152160# GND efet w=4500 l=780
+ ad=0 pd=0 as=0 ps=0 
M1680 GND diff_66480_154320# diff_56880_156000# GND efet w=2640 l=840
+ ad=0 pd=0 as=0 ps=0 
M1681 diff_50640_154200# diff_66480_154320# Vdd GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M1682 diff_81480_155160# diff_80400_153720# GND GND efet w=2280 l=840
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1683 diff_66480_154320# diff_80760_144360# diff_81480_155160# GND efet w=2160 l=720
+ ad=6.28704e+07 pd=154320 as=0 ps=0 
M1684 diff_56880_156000# Vdd Vdd GND efet w=660 l=2700
+ ad=0 pd=0 as=0 ps=0 
M1685 Vdd Vdd Vdd GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M1686 Vdd Vdd Vdd GND efet w=180 l=660
+ ad=0 pd=0 as=0 ps=0 
M1687 diff_90600_158880# diff_89400_145800# diff_66480_162000# GND efet w=2160 l=840
+ ad=2.376e+06 pd=7200 as=0 ps=0 
M1688 GND diff_88080_162120# diff_90600_158880# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1689 diff_95160_159240# diff_94080_162000# GND GND efet w=2580 l=780
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1690 GND diff_101760_182040# diff_104280_183840# GND efet w=2280 l=840
+ ad=0 pd=0 as=0 ps=0 
M1691 diff_108840_183480# diff_107880_181920# GND GND efet w=2280 l=720
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1692 diff_66480_182520# diff_108240_144360# diff_108840_183480# GND efet w=2160 l=840
+ ad=0 pd=0 as=0 ps=0 
M1693 GND diff_115560_196200# diff_118080_198000# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1694 diff_122640_197640# diff_121560_196200# GND GND efet w=2520 l=780
+ ad=0 pd=0 as=0 ps=0 
M1695 GND diff_129240_210480# diff_131760_212280# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1696 diff_136320_211920# diff_135360_210360# GND GND efet w=2280 l=720
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1697 diff_66480_210960# diff_135720_144480# diff_136320_211920# GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M1698 GND diff_143040_224520# diff_145440_226440# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1699 diff_150120_225960# diff_149040_224640# GND GND efet w=2280 l=840
+ ad=2.3328e+06 pd=7440 as=0 ps=0 
M1700 diff_66480_225120# diff_149520_144360# diff_150120_225960# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M1701 diff_145440_215640# diff_144360_145800# diff_66480_218640# GND efet w=2160 l=720
+ ad=2.6064e+06 pd=7440 as=0 ps=0 
M1702 GND diff_143040_218880# diff_145440_215640# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1703 diff_150120_216000# diff_149040_218760# GND GND efet w=2280 l=840
+ ad=2.3472e+06 pd=7440 as=0 ps=0 
M1704 GND diff_156720_238680# diff_159240_240600# GND efet w=2280 l=840
+ ad=0 pd=0 as=0 ps=0 
M1705 diff_163800_240120# diff_162840_238680# GND GND efet w=2280 l=720
+ ad=2.3616e+06 pd=7440 as=0 ps=0 
M1706 diff_66480_239280# diff_163320_144240# diff_163800_240120# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M1707 diff_159240_229800# diff_158160_145800# diff_66480_232800# GND efet w=2160 l=720
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1708 GND diff_156720_233040# diff_159240_229800# GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M1709 diff_163800_230160# diff_162840_232800# GND GND efet w=2280 l=720
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1710 GND diff_170520_252840# diff_172920_254760# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1711 diff_177600_254280# diff_176520_252960# GND GND efet w=2280 l=720
+ ad=2.376e+06 pd=7440 as=0 ps=0 
M1712 diff_66480_253440# diff_177000_144360# diff_177600_254280# GND efet w=2100 l=780
+ ad=0 pd=0 as=0 ps=0 
M1713 diff_172920_243960# diff_171960_145800# diff_66360_247080# GND efet w=2160 l=720
+ ad=2.6208e+06 pd=7440 as=0 ps=0 
M1714 GND diff_170520_247200# diff_172920_243960# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1715 diff_177600_244320# diff_176520_247080# GND GND efet w=2280 l=720
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1716 diff_186720_258120# diff_185640_145800# diff_66360_261120# GND efet w=2160 l=720
+ ad=2.6208e+06 pd=7680 as=0 ps=0 
M1717 GND diff_184200_262200# diff_186720_258120# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1718 diff_191400_258480# diff_190320_261240# GND GND efet w=2280 l=720
+ ad=2.376e+06 pd=7440 as=0 ps=0 
M1719 diff_54840_260160# diff_194400_149640# diff_190320_261240# GND efet w=780 l=780
+ ad=0 pd=0 as=2.6496e+06 ps=7440 
M1720 diff_198000_261480# diff_197280_145800# diff_54840_260160# GND efet w=840 l=720
+ ad=2.6208e+06 pd=7920 as=0 ps=0 
M1721 diff_66360_261120# diff_190800_144240# diff_191400_258480# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1722 diff_186720_254760# diff_185640_145800# diff_66480_253440# GND efet w=2040 l=720
+ ad=2.664e+06 pd=7680 as=0 ps=0 
M1723 diff_54840_253440# diff_180600_149640# diff_176520_252960# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6496e+06 ps=7440 
M1724 diff_184320_252840# diff_183480_145800# diff_54840_253440# GND efet w=840 l=840
+ ad=2.5488e+06 pd=7680 as=0 ps=0 
M1725 diff_54840_246000# diff_180600_149640# diff_176520_247080# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6496e+06 ps=7440 
M1726 diff_184200_247200# diff_183480_145800# diff_54840_246000# GND efet w=900 l=780
+ ad=2.5344e+06 pd=8400 as=0 ps=0 
M1727 diff_66360_247080# diff_177000_144360# diff_177600_244320# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1728 diff_172920_240720# diff_171960_145800# diff_66480_239280# GND efet w=2040 l=720
+ ad=2.6064e+06 pd=7680 as=0 ps=0 
M1729 diff_66480_239280# diff_177000_144360# diff_177600_240120# GND efet w=2160 l=840
+ ad=0 pd=0 as=2.3904e+06 ps=7440 
M1730 diff_54840_239280# diff_166800_149760# diff_162840_238680# GND efet w=840 l=720
+ ad=0 pd=0 as=2.5344e+06 ps=7680 
M1731 diff_170520_238680# diff_169680_145800# diff_54840_239280# GND efet w=840 l=720
+ ad=2.592e+06 pd=7680 as=0 ps=0 
M1732 diff_54840_231960# diff_166800_149760# diff_162840_232800# GND efet w=840 l=720
+ ad=0 pd=0 as=2.4048e+06 ps=7440 
M1733 diff_170520_233040# diff_169680_145800# diff_54840_231960# GND efet w=840 l=720
+ ad=2.3904e+06 pd=7200 as=0 ps=0 
M1734 diff_66480_232800# diff_163320_144240# diff_163800_230160# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1735 diff_159240_226440# diff_158160_145800# diff_66480_225120# GND efet w=2040 l=720
+ ad=2.3616e+06 pd=7440 as=0 ps=0 
M1736 diff_54840_225240# diff_153120_145800# diff_149040_224640# GND efet w=840 l=840
+ ad=0 pd=0 as=2.5056e+06 ps=7440 
M1737 diff_156720_224520# diff_155880_145800# diff_54840_225240# GND efet w=840 l=720
+ ad=2.6064e+06 pd=7440 as=0 ps=0 
M1738 diff_54840_217800# diff_153120_145800# diff_149040_218760# GND efet w=960 l=720
+ ad=0 pd=0 as=2.4912e+06 ps=7440 
M1739 diff_156720_218880# diff_155880_145800# diff_54840_217800# GND efet w=840 l=720
+ ad=2.6496e+06 pd=7440 as=0 ps=0 
M1740 diff_66480_218640# diff_149520_144360# diff_150120_216000# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1741 diff_145440_212400# diff_144360_145800# diff_66480_210960# GND efet w=2160 l=720
+ ad=2.592e+06 pd=7440 as=0 ps=0 
M1742 diff_54840_210960# diff_139320_149640# diff_135360_210360# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6352e+06 ps=7440 
M1743 diff_143040_210480# diff_142200_145800# diff_54840_210960# GND efet w=960 l=720
+ ad=2.6208e+06 pd=7440 as=0 ps=0 
M1744 diff_131760_201480# diff_130680_145800# diff_66480_204480# GND efet w=2160 l=720
+ ad=2.3904e+06 pd=7440 as=0 ps=0 
M1745 GND diff_129240_204720# diff_131760_201480# GND efet w=2700 l=780
+ ad=0 pd=0 as=0 ps=0 
M1746 diff_136320_201840# diff_135360_204480# GND GND efet w=2280 l=720
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1747 diff_54840_203640# diff_139320_149640# diff_135360_204480# GND efet w=840 l=720
+ ad=0 pd=0 as=2.664e+06 ps=7440 
M1748 diff_143040_204840# diff_142200_145800# diff_54840_203640# GND efet w=840 l=720
+ ad=2.592e+06 pd=7440 as=0 ps=0 
M1749 diff_66480_204480# diff_135720_144480# diff_136320_201840# GND efet w=2160 l=840
+ ad=0 pd=0 as=0 ps=0 
M1750 diff_131760_198120# diff_130680_145800# diff_66480_196680# GND efet w=2160 l=780
+ ad=2.3904e+06 pd=7440 as=0 ps=0 
M1751 GND diff_129240_196200# diff_131760_198120# GND efet w=2700 l=780
+ ad=0 pd=0 as=0 ps=0 
M1752 diff_54840_196800# diff_125640_145800# diff_121560_196200# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6352e+06 ps=7680 
M1753 diff_129240_196200# diff_128400_145800# diff_54840_196800# GND efet w=840 l=720
+ ad=2.6928e+06 pd=7680 as=0 ps=0 
M1754 diff_118080_187200# diff_116880_145800# diff_66480_190200# GND efet w=2160 l=840
+ ad=2.448e+06 pd=7440 as=0 ps=0 
M1755 GND diff_115560_190440# diff_118080_187200# GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M1756 diff_122640_187560# diff_121560_190320# GND GND efet w=2460 l=780
+ ad=2.4048e+06 pd=7440 as=0 ps=0 
M1757 diff_54840_189360# diff_125640_145800# diff_121560_190320# GND efet w=960 l=720
+ ad=0 pd=0 as=2.736e+06 ps=7920 
M1758 diff_129240_190440# diff_128400_145800# diff_54840_189360# GND efet w=960 l=720
+ ad=2.7504e+06 pd=7920 as=0 ps=0 
M1759 diff_66480_190200# diff_122040_144240# diff_122640_187560# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1760 diff_118080_183720# diff_116880_145800# diff_66480_182520# GND efet w=2220 l=900
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1761 diff_54840_182640# diff_111840_149760# diff_107880_181920# GND efet w=840 l=720
+ ad=0 pd=0 as=2.664e+06 ps=7440 
M1762 diff_115560_181920# diff_114720_145800# diff_54840_182640# GND efet w=840 l=720
+ ad=2.6064e+06 pd=7440 as=0 ps=0 
M1763 diff_104280_173040# diff_103200_145800# diff_66480_176040# GND efet w=2160 l=720
+ ad=2.3904e+06 pd=7440 as=0 ps=0 
M1764 GND diff_101760_176400# diff_104280_173040# GND efet w=2280 l=840
+ ad=0 pd=0 as=0 ps=0 
M1765 diff_108840_173400# diff_107880_176160# GND GND efet w=2280 l=720
+ ad=2.4048e+06 pd=7440 as=0 ps=0 
M1766 diff_54840_175200# diff_111840_149760# diff_107880_176160# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6784e+06 ps=7440 
M1767 diff_115560_176280# diff_114720_145800# diff_54840_175200# GND efet w=840 l=720
+ ad=2.5488e+06 pd=7440 as=0 ps=0 
M1768 diff_66480_176040# diff_108240_144360# diff_108840_173400# GND efet w=2280 l=840
+ ad=0 pd=0 as=0 ps=0 
M1769 diff_104280_169680# diff_103200_145800# diff_66480_168360# GND efet w=2160 l=780
+ ad=2.448e+06 pd=7440 as=0 ps=0 
M1770 diff_54840_168480# diff_98160_145800# diff_94080_167760# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6208e+06 ps=7680 
M1771 diff_101760_167760# diff_100920_145800# diff_54840_168480# GND efet w=900 l=720
+ ad=2.6352e+06 pd=7440 as=0 ps=0 
M1772 diff_54840_161040# diff_98160_145800# diff_94080_162000# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6928e+06 ps=7920 
M1773 diff_101880_162120# diff_100920_145800# diff_54840_161040# GND efet w=840 l=840
+ ad=2.5776e+06 pd=7680 as=0 ps=0 
M1774 diff_66480_162000# diff_94560_144240# diff_95160_159240# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1775 diff_90600_155160# diff_89400_145800# diff_66480_154320# GND efet w=2400 l=840
+ ad=2.448e+06 pd=7440 as=0 ps=0 
M1776 diff_54840_154320# diff_84360_149760# diff_80400_153720# GND efet w=840 l=840
+ ad=0 pd=0 as=2.6496e+06 ps=7440 
M1777 diff_88080_153600# diff_87240_145800# diff_54840_154320# GND efet w=900 l=780
+ ad=2.5632e+06 pd=7200 as=0 ps=0 
M1778 GND diff_88080_153600# diff_90600_155160# GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M1779 diff_95160_155040# diff_94080_153720# GND GND efet w=2460 l=780
+ ad=2.4192e+06 pd=7440 as=0 ps=0 
M1780 diff_66480_154320# diff_94560_144240# diff_95160_155040# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1781 GND diff_101760_167760# diff_104280_169680# GND efet w=2400 l=840
+ ad=0 pd=0 as=0 ps=0 
M1782 diff_108840_169200# diff_107880_167760# GND GND efet w=2400 l=720
+ ad=2.448e+06 pd=7440 as=0 ps=0 
M1783 diff_66480_168360# diff_108240_144360# diff_108840_169200# GND efet w=2220 l=900
+ ad=0 pd=0 as=0 ps=0 
M1784 GND diff_115560_181920# diff_118080_183720# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1785 diff_122640_183480# diff_121560_181920# GND GND efet w=2460 l=780
+ ad=2.3328e+06 pd=7200 as=0 ps=0 
M1786 diff_66480_182520# diff_122040_144240# diff_122640_183480# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1787 diff_118080_173040# diff_116880_145800# diff_66480_176040# GND efet w=2160 l=840
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1788 GND diff_115560_176280# diff_118080_173040# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1789 diff_122640_173400# diff_121560_176160# GND GND efet w=2700 l=780
+ ad=2.376e+06 pd=7440 as=0 ps=0 
M1790 diff_136320_197640# diff_135360_196200# GND GND efet w=2280 l=720
+ ad=2.4048e+06 pd=7200 as=0 ps=0 
M1791 diff_66480_196680# diff_135720_144480# diff_136320_197640# GND efet w=2160 l=840
+ ad=0 pd=0 as=0 ps=0 
M1792 GND diff_143040_210480# diff_145440_212400# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1793 diff_150120_211920# diff_149040_210360# GND GND efet w=2280 l=780
+ ad=2.3328e+06 pd=7200 as=0 ps=0 
M1794 diff_66480_210960# diff_149520_144360# diff_150120_211920# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1795 diff_145440_201480# diff_144360_145800# diff_66480_204480# GND efet w=2160 l=720
+ ad=2.6064e+06 pd=7440 as=0 ps=0 
M1796 GND diff_143040_204840# diff_145440_201480# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1797 diff_150120_201840# diff_149040_204480# GND GND efet w=2400 l=780
+ ad=2.3328e+06 pd=7200 as=0 ps=0 
M1798 GND diff_156720_224520# diff_159240_226440# GND efet w=2580 l=780
+ ad=0 pd=0 as=0 ps=0 
M1799 diff_163800_225960# diff_162840_224520# GND GND efet w=2280 l=720
+ ad=2.376e+06 pd=7440 as=0 ps=0 
M1800 diff_66480_225120# diff_163320_144240# diff_163800_225960# GND efet w=2100 l=780
+ ad=0 pd=0 as=0 ps=0 
M1801 GND diff_170520_238680# diff_172920_240720# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1802 diff_177600_240120# diff_176520_238800# GND GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1803 diff_172920_229800# diff_171960_145800# diff_66480_232800# GND efet w=2280 l=720
+ ad=2.5776e+06 pd=7680 as=0 ps=0 
M1804 GND diff_170520_233040# diff_172920_229800# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1805 diff_177600_230160# diff_176520_232920# GND GND efet w=2280 l=720
+ ad=2.376e+06 pd=7200 as=0 ps=0 
M1806 GND diff_184320_252840# diff_186720_254760# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1807 diff_191400_254280# diff_190320_252960# GND GND efet w=2280 l=720
+ ad=2.4048e+06 pd=7440 as=0 ps=0 
M1808 diff_66480_253440# diff_190800_144240# diff_191400_254280# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M1809 diff_186720_243960# diff_185640_145800# diff_66360_247080# GND efet w=2160 l=720
+ ad=2.6352e+06 pd=7680 as=0 ps=0 
M1810 GND diff_184200_247200# diff_186720_243960# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1811 diff_191400_244320# diff_190320_247080# GND GND efet w=2340 l=780
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1812 diff_200520_258120# diff_199440_146040# diff_66360_261120# GND efet w=2160 l=720
+ ad=2.6064e+06 pd=7680 as=0 ps=0 
M1813 GND diff_198000_261480# diff_200520_258120# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1814 diff_205200_258480# diff_204120_261240# GND GND efet w=2520 l=720
+ ad=2.3184e+06 pd=7200 as=0 ps=0 
M1815 diff_54840_260160# diff_208200_149640# diff_204120_261240# GND efet w=720 l=720
+ ad=0 pd=0 as=2.5776e+06 ps=7440 
M1816 diff_211800_261480# diff_211080_145800# diff_54840_260160# GND efet w=720 l=720
+ ad=2.5488e+06 pd=7680 as=0 ps=0 
M1817 diff_66360_261120# diff_204600_144480# diff_205200_258480# GND efet w=2100 l=780
+ ad=0 pd=0 as=0 ps=0 
M1818 diff_200520_254880# diff_199440_146040# diff_66480_253440# GND efet w=2040 l=720
+ ad=2.6064e+06 pd=7680 as=0 ps=0 
M1819 diff_54840_253440# diff_194400_149640# diff_190320_252960# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6064e+06 ps=7440 
M1820 diff_198000_252840# diff_197280_145800# diff_54840_253440# GND efet w=840 l=720
+ ad=2.5776e+06 pd=7680 as=0 ps=0 
M1821 diff_54840_246000# diff_194400_149640# diff_190320_247080# GND efet w=840 l=720
+ ad=0 pd=0 as=2.5776e+06 ps=7920 
M1822 diff_198000_247200# diff_197280_145800# diff_54840_246000# GND efet w=840 l=720
+ ad=2.592e+06 pd=7680 as=0 ps=0 
M1823 diff_66360_247080# diff_190800_144240# diff_191400_244320# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1824 diff_66480_239280# diff_190800_144240# diff_191400_240120# GND efet w=2160 l=840
+ ad=0 pd=0 as=2.3472e+06 ps=7440 
M1825 diff_186720_240720# diff_185640_145800# diff_66480_239280# GND efet w=2040 l=720
+ ad=2.5776e+06 pd=7680 as=0 ps=0 
M1826 GND diff_184200_238920# diff_186720_240720# GND efet w=2340 l=900
+ ad=0 pd=0 as=0 ps=0 
M1827 diff_54840_239280# diff_180600_149640# diff_176520_238800# GND efet w=840 l=720
+ ad=0 pd=0 as=2.7504e+06 ps=7680 
M1828 diff_184200_238920# diff_183480_145800# diff_54840_239280# GND efet w=1080 l=780
+ ad=2.5776e+06 pd=8160 as=0 ps=0 
M1829 diff_54840_231960# diff_180600_149640# diff_176520_232920# GND efet w=840 l=720
+ ad=0 pd=0 as=2.5488e+06 ps=7680 
M1830 diff_184200_233400# diff_183480_145800# diff_54840_231960# GND efet w=960 l=720
+ ad=2.5344e+06 pd=7680 as=0 ps=0 
M1831 diff_66480_232800# diff_177000_144360# diff_177600_230160# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1832 diff_172920_226440# diff_171960_145800# diff_66480_225120# GND efet w=2160 l=720
+ ad=2.52e+06 pd=7920 as=0 ps=0 
M1833 diff_54840_225240# diff_166800_149760# diff_162840_224520# GND efet w=840 l=720
+ ad=0 pd=0 as=2.5344e+06 ps=7680 
M1834 diff_170520_224520# diff_169680_145800# diff_54840_225240# GND efet w=840 l=720
+ ad=2.6496e+06 pd=7680 as=0 ps=0 
M1835 diff_54840_217800# diff_166800_149760# diff_162840_218760# GND efet w=840 l=720
+ ad=0 pd=0 as=2.5056e+06 ps=7440 
M1836 diff_170520_218880# diff_169680_145800# diff_54840_217800# GND efet w=840 l=720
+ ad=2.5344e+06 pd=7440 as=0 ps=0 
M1837 diff_159240_215640# diff_158160_145800# diff_66480_218640# GND efet w=2160 l=720
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1838 GND diff_156720_218880# diff_159240_215640# GND efet w=2460 l=780
+ ad=0 pd=0 as=0 ps=0 
M1839 diff_163800_216000# diff_162840_218760# GND GND efet w=2280 l=720
+ ad=2.3616e+06 pd=7440 as=0 ps=0 
M1840 diff_66480_218640# diff_163320_144240# diff_163800_216000# GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M1841 diff_159240_212280# diff_158160_145800# diff_66480_210960# GND efet w=2160 l=720
+ ad=2.376e+06 pd=7200 as=0 ps=0 
M1842 diff_66480_210960# diff_163320_144240# diff_163800_211920# GND efet w=2400 l=720
+ ad=0 pd=0 as=2.4768e+06 ps=7680 
M1843 diff_54840_210960# diff_153120_145800# diff_149040_210360# GND efet w=720 l=720
+ ad=0 pd=0 as=2.6928e+06 ps=7680 
M1844 diff_156720_210360# diff_155880_145800# diff_54840_210960# GND efet w=720 l=720
+ ad=2.664e+06 pd=7440 as=0 ps=0 
M1845 diff_54840_203640# diff_153120_145800# diff_149040_204480# GND efet w=960 l=720
+ ad=0 pd=0 as=2.6784e+06 ps=7440 
M1846 diff_156720_204720# diff_155880_145800# diff_54840_203640# GND efet w=840 l=720
+ ad=2.664e+06 pd=7440 as=0 ps=0 
M1847 diff_66480_204480# diff_149520_144360# diff_150120_201840# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1848 diff_145440_198120# diff_144360_145800# diff_66480_196680# GND efet w=2100 l=780
+ ad=2.6208e+06 pd=7440 as=0 ps=0 
M1849 diff_54840_196800# diff_139320_149640# diff_135360_196200# GND efet w=960 l=720
+ ad=0 pd=0 as=2.736e+06 ps=7920 
M1850 diff_143040_196080# diff_142200_145800# diff_54840_196800# GND efet w=840 l=720
+ ad=2.736e+06 pd=7680 as=0 ps=0 
M1851 diff_131760_187200# diff_130680_145800# diff_66480_190200# GND efet w=2160 l=720
+ ad=2.232e+06 pd=7440 as=0 ps=0 
M1852 GND diff_129240_190440# diff_131760_187200# GND efet w=2460 l=780
+ ad=0 pd=0 as=0 ps=0 
M1853 diff_136320_187560# diff_135360_190320# GND GND efet w=2400 l=720
+ ad=2.4624e+06 pd=7440 as=0 ps=0 
M1854 diff_54840_189360# diff_139320_149640# diff_135360_190320# GND efet w=960 l=720
+ ad=0 pd=0 as=2.6784e+06 ps=7440 
M1855 diff_143040_190440# diff_142200_145800# diff_54840_189360# GND efet w=960 l=720
+ ad=2.6064e+06 pd=7680 as=0 ps=0 
M1856 diff_66480_190200# diff_135720_144480# diff_136320_187560# GND efet w=2160 l=840
+ ad=0 pd=0 as=0 ps=0 
M1857 diff_131760_183840# diff_130680_145800# diff_66480_182520# GND efet w=2160 l=720
+ ad=2.376e+06 pd=7200 as=0 ps=0 
M1858 diff_54840_182640# diff_125640_145800# diff_121560_181920# GND efet w=840 l=720
+ ad=0 pd=0 as=2.664e+06 ps=7920 
M1859 diff_129240_182040# diff_128400_145800# diff_54840_182640# GND efet w=840 l=720
+ ad=2.5632e+06 pd=7440 as=0 ps=0 
M1860 diff_54840_175200# diff_125640_145800# diff_121560_176160# GND efet w=900 l=720
+ ad=0 pd=0 as=2.6064e+06 ps=7920 
M1861 diff_129240_176400# diff_128400_145800# diff_54840_175200# GND efet w=840 l=720
+ ad=2.4048e+06 pd=7440 as=0 ps=0 
M1862 diff_66480_176040# diff_122040_144240# diff_122640_173400# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1863 diff_118080_169440# diff_116880_145800# diff_66480_168360# GND efet w=2160 l=960
+ ad=2.3904e+06 pd=7200 as=0 ps=0 
M1864 GND diff_115560_167760# diff_118080_169440# GND efet w=2340 l=900
+ ad=0 pd=0 as=0 ps=0 
M1865 diff_54840_168480# diff_111840_149760# diff_107880_167760# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6496e+06 ps=7440 
M1866 diff_115560_167760# diff_114720_145800# diff_54840_168480# GND efet w=840 l=720
+ ad=2.6064e+06 pd=7440 as=0 ps=0 
M1867 diff_104280_158880# diff_103200_145800# diff_66480_162000# GND efet w=2160 l=720
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1868 GND diff_101880_162120# diff_104280_158880# GND efet w=2280 l=840
+ ad=0 pd=0 as=0 ps=0 
M1869 diff_108840_159240# diff_107880_162000# GND GND efet w=2280 l=720
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1870 diff_54840_161040# diff_111840_149760# diff_107880_162000# GND efet w=840 l=720
+ ad=0 pd=0 as=2.664e+06 ps=7440 
M1871 diff_115560_162120# diff_114720_145800# diff_54840_161040# GND efet w=840 l=720
+ ad=2.5488e+06 pd=7200 as=0 ps=0 
M1872 diff_66480_162000# diff_108240_144360# diff_108840_159240# GND efet w=2160 l=840
+ ad=0 pd=0 as=0 ps=0 
M1873 diff_104280_155520# diff_103200_145800# diff_66480_154320# GND efet w=2160 l=720
+ ad=2.4336e+06 pd=7440 as=0 ps=0 
M1874 diff_54840_154320# diff_98160_145800# diff_94080_153720# GND efet w=960 l=840
+ ad=0 pd=0 as=2.7072e+06 ps=7920 
M1875 diff_101880_152880# diff_100920_145800# diff_54840_154320# GND efet w=900 l=900
+ ad=2.5776e+06 pd=7440 as=0 ps=0 
M1876 GND diff_101880_152880# diff_104280_155520# GND efet w=2400 l=840
+ ad=0 pd=0 as=0 ps=0 
M1877 diff_108840_155040# diff_107880_153720# GND GND efet w=2400 l=720
+ ad=2.4912e+06 pd=7920 as=0 ps=0 
M1878 diff_66480_154320# diff_108240_144360# diff_108840_155040# GND efet w=2400 l=840
+ ad=0 pd=0 as=0 ps=0 
M1879 diff_122640_169200# diff_121560_167760# GND GND efet w=2400 l=960
+ ad=2.4048e+06 pd=7440 as=0 ps=0 
M1880 diff_66480_168360# diff_122040_144240# diff_122640_169200# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M1881 diff_118080_158880# diff_116880_145800# diff_66480_162000# GND efet w=2160 l=840
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1882 GND diff_115560_162120# diff_118080_158880# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1883 diff_122640_159240# diff_121560_162000# GND GND efet w=2280 l=780
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1884 GND diff_129240_182040# diff_131760_183840# GND efet w=2340 l=780
+ ad=0 pd=0 as=0 ps=0 
M1885 diff_136320_183480# diff_135360_181920# GND GND efet w=2280 l=720
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1886 diff_66480_182520# diff_135720_144480# diff_136320_183480# GND efet w=2160 l=840
+ ad=0 pd=0 as=0 ps=0 
M1887 GND diff_143040_196080# diff_145440_198120# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1888 diff_150120_197640# diff_149040_196200# GND GND efet w=2280 l=780
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1889 diff_66480_196680# diff_149520_144360# diff_150120_197640# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M1890 diff_145440_187200# diff_144360_145800# diff_66480_190200# GND efet w=2160 l=720
+ ad=2.7216e+06 pd=7680 as=0 ps=0 
M1891 GND diff_143040_190440# diff_145440_187200# GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M1892 diff_150120_187560# diff_149040_190320# GND GND efet w=2460 l=780
+ ad=2.4192e+06 pd=7440 as=0 ps=0 
M1893 GND diff_156720_210360# diff_159240_212280# GND efet w=2280 l=780
+ ad=0 pd=0 as=0 ps=0 
M1894 diff_163800_211920# diff_162840_210360# GND GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1895 GND diff_156720_204720# diff_159240_201480# GND efet w=2400 l=780
+ ad=0 pd=0 as=2.376e+06 ps=7440 
M1896 diff_159240_201480# diff_158160_145800# diff_66480_204480# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1897 diff_163800_201840# diff_162840_204480# GND GND efet w=2280 l=720
+ ad=2.6352e+06 pd=7680 as=0 ps=0 
M1898 GND diff_170520_224520# diff_172920_226440# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1899 diff_177600_225960# diff_176520_224640# GND GND efet w=2280 l=720
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1900 diff_66480_225120# diff_177000_144360# diff_177600_225960# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M1901 diff_172920_215880# diff_171960_145800# diff_66480_218640# GND efet w=2280 l=780
+ ad=2.4048e+06 pd=7680 as=0 ps=0 
M1902 GND diff_170520_218880# diff_172920_215880# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1903 diff_177600_216000# diff_176520_218880# GND GND efet w=2280 l=720
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1904 diff_191400_240120# diff_190320_238680# GND GND efet w=2400 l=840
+ ad=0 pd=0 as=0 ps=0 
M1905 diff_186720_229800# diff_185640_145800# diff_66480_232800# GND efet w=2160 l=720
+ ad=2.6352e+06 pd=7680 as=0 ps=0 
M1906 GND diff_184200_233400# diff_186720_229800# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1907 diff_191400_230160# diff_190320_232920# GND GND efet w=2400 l=720
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1908 GND diff_198000_252840# diff_200520_254880# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1909 diff_205200_254280# diff_204120_252840# GND GND efet w=2460 l=780
+ ad=2.3904e+06 pd=7440 as=0 ps=0 
M1910 diff_66480_253440# diff_204600_144480# diff_205200_254280# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M1911 diff_200520_243960# diff_199440_146040# diff_66360_247080# GND efet w=2160 l=720
+ ad=2.6064e+06 pd=7680 as=0 ps=0 
M1912 GND diff_198000_247200# diff_200520_243960# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1913 diff_205080_245640# diff_204120_247080# GND GND efet w=2520 l=780
+ ad=2.3472e+06 pd=7680 as=0 ps=0 
M1914 Vdd diff_189240_66360# diff_54840_260160# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M1915 diff_214320_258120# diff_213360_145800# diff_66360_261120# GND efet w=2160 l=720
+ ad=2.6928e+06 pd=7680 as=0 ps=0 
M1916 GND diff_211800_261480# diff_214320_258120# GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M1917 Vdd diff_222480_158400# diff_66360_261120# GND efet w=1440 l=660
+ ad=0 pd=0 as=0 ps=0 
M1918 diff_241560_285240# Vdd Vdd GND efet w=1080 l=1920
+ ad=0 pd=0 as=0 ps=0 
M1919 Vdd Vdd Vdd GND efet w=540 l=300
+ ad=0 pd=0 as=0 ps=0 
M1920 Vdd Vdd Vdd GND efet w=420 l=780
+ ad=0 pd=0 as=0 ps=0 
M1921 diff_241440_260160# Vdd Vdd GND efet w=1320 l=1860
+ ad=1.25424e+07 pd=26160 as=0 ps=0 
M1922 diff_232560_257640# clk2 diff_23040_212640# GND efet w=1920 l=720
+ ad=2.736e+06 pd=7680 as=0 ps=0 
M1923 diff_234480_257040# diff_207480_277200# diff_232560_257640# GND efet w=1920 l=720
+ ad=1.67184e+07 pd=32640 as=0 ps=0 
M1924 diff_214320_254880# diff_213360_145800# diff_66480_253440# GND efet w=2040 l=720
+ ad=2.1024e+06 pd=6480 as=0 ps=0 
M1925 GND diff_211800_252840# diff_214320_254880# GND efet w=1680 l=720
+ ad=0 pd=0 as=0 ps=0 
M1926 diff_54840_253440# diff_208200_149640# diff_204120_252840# GND efet w=840 l=840
+ ad=0 pd=0 as=2.5776e+06 ps=7440 
M1927 diff_211800_252840# diff_211080_145800# diff_54840_253440# GND efet w=840 l=720
+ ad=2.5776e+06 pd=7680 as=0 ps=0 
M1928 diff_54840_246000# diff_208200_149640# diff_204120_247080# GND efet w=780 l=900
+ ad=0 pd=0 as=2.4192e+06 ps=8640 
M1929 diff_211800_247200# diff_211080_145800# diff_54840_246000# GND efet w=840 l=840
+ ad=2.5344e+06 pd=7440 as=0 ps=0 
M1930 diff_66360_247080# diff_204600_144480# diff_205080_245640# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1931 diff_200520_240720# diff_199440_146040# diff_66480_239280# GND efet w=2100 l=780
+ ad=2.52e+06 pd=7680 as=0 ps=0 
M1932 diff_54840_239280# diff_194400_149640# diff_190320_238680# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6352e+06 ps=7440 
M1933 diff_198000_238680# diff_197280_145800# diff_54840_239280# GND efet w=840 l=720
+ ad=2.6208e+06 pd=7680 as=0 ps=0 
M1934 diff_54840_231960# diff_194400_149640# diff_190320_232920# GND efet w=900 l=780
+ ad=0 pd=0 as=2.6784e+06 ps=7440 
M1935 diff_198000_233040# diff_197280_145800# diff_54840_231960# GND efet w=840 l=720
+ ad=2.6208e+06 pd=7680 as=0 ps=0 
M1936 diff_66480_232800# diff_190800_144240# diff_191400_230160# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1937 diff_186720_226560# diff_185640_145800# diff_66480_225120# GND efet w=2040 l=720
+ ad=2.592e+06 pd=7440 as=0 ps=0 
M1938 diff_54840_225240# diff_180600_149640# diff_176520_224640# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6208e+06 ps=7680 
M1939 diff_184200_225120# diff_183480_145800# diff_54840_225240# GND efet w=1020 l=720
+ ad=2.5776e+06 pd=7920 as=0 ps=0 
M1940 diff_54840_217800# diff_180600_149640# diff_176520_218880# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6496e+06 ps=7440 
M1941 diff_184320_218880# diff_183480_145800# diff_54840_217800# GND efet w=840 l=840
+ ad=2.5632e+06 pd=7680 as=0 ps=0 
M1942 diff_66480_218640# diff_177000_144360# diff_177600_216000# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1943 diff_173040_212280# diff_171960_145800# diff_66480_210960# GND efet w=2160 l=840
+ ad=2.4336e+06 pd=7440 as=0 ps=0 
M1944 diff_54840_210960# diff_166800_149760# diff_162840_210360# GND efet w=780 l=780
+ ad=0 pd=0 as=2.5344e+06 ps=7440 
M1945 diff_170520_210360# diff_169680_145800# diff_54840_210960# GND efet w=840 l=840
+ ad=2.5488e+06 pd=7440 as=0 ps=0 
M1946 GND diff_170520_210360# diff_173040_212280# GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M1947 diff_177600_211800# diff_176520_210960# GND GND efet w=2400 l=720
+ ad=2.4048e+06 pd=7440 as=0 ps=0 
M1948 diff_66480_210960# diff_177000_144360# diff_177600_211800# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1949 diff_170520_204720# diff_169680_145800# diff_54840_203640# GND efet w=960 l=840
+ ad=2.52e+06 pd=7440 as=0 ps=0 
M1950 diff_54840_203640# diff_166800_149760# diff_162840_204480# GND efet w=840 l=720
+ ad=0 pd=0 as=2.5344e+06 ps=7440 
M1951 diff_66480_204480# diff_163320_144240# diff_163800_201840# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1952 diff_159240_198120# diff_158160_145800# diff_66480_196680# GND efet w=2040 l=720
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1953 diff_54840_196800# diff_153120_145800# diff_149040_196200# GND efet w=840 l=720
+ ad=0 pd=0 as=2.592e+06 ps=7440 
M1954 diff_156720_196200# diff_155880_145800# diff_54840_196800# GND efet w=840 l=720
+ ad=2.6064e+06 pd=7920 as=0 ps=0 
M1955 diff_54840_189360# diff_153120_145800# diff_149040_190320# GND efet w=900 l=780
+ ad=0 pd=0 as=2.6784e+06 ps=7440 
M1956 diff_156720_190440# diff_155880_145800# diff_54840_189360# GND efet w=960 l=720
+ ad=2.7072e+06 pd=7920 as=0 ps=0 
M1957 diff_66480_190200# diff_149520_144360# diff_150120_187560# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1958 diff_145440_183960# diff_144360_145800# diff_66480_182520# GND efet w=2160 l=720
+ ad=2.6208e+06 pd=7440 as=0 ps=0 
M1959 diff_54840_182640# diff_139320_149640# diff_135360_181920# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6496e+06 ps=7440 
M1960 diff_143040_181920# diff_142200_145800# diff_54840_182640# GND efet w=840 l=720
+ ad=2.6208e+06 pd=7440 as=0 ps=0 
M1961 GND diff_129240_176400# diff_131760_173040# GND efet w=2580 l=780
+ ad=0 pd=0 as=2.3904e+06 ps=7440 
M1962 diff_131760_173040# diff_130680_145800# diff_66480_176040# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1963 diff_136320_173400# diff_135360_176040# GND GND efet w=2280 l=720
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M1964 diff_54840_175200# diff_139320_149640# diff_135360_176040# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6352e+06 ps=7440 
M1965 diff_143040_176400# diff_142200_145800# diff_54840_175200# GND efet w=840 l=720
+ ad=2.5056e+06 pd=7440 as=0 ps=0 
M1966 diff_66480_176040# diff_135720_144480# diff_136320_173400# GND efet w=2160 l=840
+ ad=0 pd=0 as=0 ps=0 
M1967 diff_131760_169680# diff_130680_145800# diff_66480_168360# GND efet w=2040 l=720
+ ad=2.3904e+06 pd=7440 as=0 ps=0 
M1968 diff_54840_168480# diff_125640_145800# diff_121560_167760# GND efet w=960 l=840
+ ad=0 pd=0 as=2.592e+06 ps=7920 
M1969 diff_129240_167760# diff_128400_145800# diff_54840_168480# GND efet w=840 l=720
+ ad=2.6064e+06 pd=7680 as=0 ps=0 
M1970 diff_54840_161040# diff_125640_145800# diff_121560_162000# GND efet w=1020 l=780
+ ad=0 pd=0 as=2.592e+06 ps=8400 
M1971 diff_129240_162120# diff_128400_145800# diff_54840_161040# GND efet w=840 l=720
+ ad=2.52e+06 pd=7920 as=0 ps=0 
M1972 diff_66480_162000# diff_122040_144240# diff_122640_159240# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1973 diff_118080_155400# diff_116880_145800# diff_66480_154320# GND efet w=2160 l=840
+ ad=2.4192e+06 pd=7440 as=0 ps=0 
M1974 diff_54840_154320# diff_111840_149760# diff_107880_153720# GND efet w=900 l=780
+ ad=0 pd=0 as=2.6928e+06 ps=7440 
M1975 diff_115560_153600# diff_114720_145800# diff_54840_154320# GND efet w=960 l=720
+ ad=2.5632e+06 pd=7200 as=0 ps=0 
M1976 GND diff_115560_153600# diff_118080_155400# GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M1977 diff_122640_155040# diff_121560_153720# GND GND efet w=2580 l=780
+ ad=2.376e+06 pd=7680 as=0 ps=0 
M1978 diff_66480_154320# diff_122040_144240# diff_122640_155040# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1979 GND diff_129240_167760# diff_131760_169680# GND efet w=2340 l=780
+ ad=0 pd=0 as=0 ps=0 
M1980 diff_136320_169200# diff_135360_167760# GND GND efet w=2280 l=720
+ ad=2.376e+06 pd=7200 as=0 ps=0 
M1981 diff_66480_168360# diff_135720_144480# diff_136320_169200# GND efet w=2040 l=840
+ ad=0 pd=0 as=0 ps=0 
M1982 diff_131760_158880# diff_130680_145800# diff_66480_162000# GND efet w=2160 l=720
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M1983 GND diff_129240_162120# diff_131760_158880# GND efet w=2400 l=780
+ ad=0 pd=0 as=0 ps=0 
M1984 diff_136320_159240# diff_135360_162000# GND GND efet w=2280 l=720
+ ad=2.3328e+06 pd=7200 as=0 ps=0 
M1985 GND diff_143040_181920# diff_145440_183960# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1986 diff_150120_183480# diff_149040_181920# GND GND efet w=2520 l=780
+ ad=2.3328e+06 pd=7440 as=0 ps=0 
M1987 diff_66480_182520# diff_149520_144360# diff_150120_183480# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1988 diff_145440_173040# diff_144360_145800# diff_66480_176040# GND efet w=2280 l=720
+ ad=2.592e+06 pd=7680 as=0 ps=0 
M1989 GND diff_143040_176400# diff_145440_173040# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1990 diff_150120_173400# diff_149040_176160# GND GND efet w=2280 l=840
+ ad=2.3328e+06 pd=7200 as=0 ps=0 
M1991 GND diff_156720_196200# diff_159240_198120# GND efet w=2280 l=840
+ ad=0 pd=0 as=0 ps=0 
M1992 diff_163800_197640# diff_162840_196200# GND GND efet w=2280 l=720
+ ad=2.5632e+06 pd=7680 as=0 ps=0 
M1993 diff_66480_196680# diff_163320_144240# diff_163800_197640# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M1994 diff_159240_187200# diff_158160_145800# diff_66480_190200# GND efet w=2160 l=720
+ ad=2.4624e+06 pd=7440 as=0 ps=0 
M1995 GND diff_156720_190440# diff_159240_187200# GND efet w=2400 l=840
+ ad=0 pd=0 as=0 ps=0 
M1996 diff_163800_187560# diff_162840_190320# GND GND efet w=2400 l=720
+ ad=2.6928e+06 pd=7920 as=0 ps=0 
M1997 diff_173040_201480# diff_171960_145800# diff_66480_204480# GND efet w=2160 l=840
+ ad=2.1888e+06 pd=7200 as=0 ps=0 
M1998 GND diff_170520_204720# diff_173040_201480# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M1999 diff_177600_201840# diff_176640_204480# GND GND efet w=2280 l=720
+ ad=2.376e+06 pd=7440 as=0 ps=0 
M2000 GND diff_184200_225120# diff_186720_226560# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2001 diff_191400_225960# diff_190320_224640# GND GND efet w=2700 l=780
+ ad=2.3904e+06 pd=7200 as=0 ps=0 
M2002 diff_66480_225120# diff_190800_144240# diff_191400_225960# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M2003 diff_186720_215640# diff_185640_145800# diff_66480_218640# GND efet w=2160 l=720
+ ad=2.5776e+06 pd=7680 as=0 ps=0 
M2004 GND diff_184320_218880# diff_186720_215640# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2005 diff_191400_216000# diff_190320_218760# GND GND efet w=2520 l=720
+ ad=2.3184e+06 pd=7200 as=0 ps=0 
M2006 GND diff_198000_238680# diff_200520_240720# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2007 diff_205200_240240# diff_204120_238680# GND GND efet w=2220 l=780
+ ad=2.232e+06 pd=6960 as=0 ps=0 
M2008 diff_66480_239280# diff_204600_144480# diff_205200_240240# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M2009 diff_200520_229800# diff_199440_146040# diff_66480_232800# GND efet w=2160 l=720
+ ad=2.6208e+06 pd=7680 as=0 ps=0 
M2010 GND diff_198000_233040# diff_200520_229800# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2011 diff_205200_230160# diff_204120_232920# GND GND efet w=2700 l=780
+ ad=2.3184e+06 pd=7200 as=0 ps=0 
M2012 Vdd diff_222480_158400# diff_66480_253440# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M2013 Vdd diff_189240_66360# diff_54840_253440# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2014 GND diff_207480_277200# diff_242400_251880# GND efet w=1560 l=600
+ ad=0 pd=0 as=3.8736e+06 ps=8400 
M2015 GND diff_207720_290040# diff_234480_257040# GND efet w=2820 l=660
+ ad=0 pd=0 as=0 ps=0 
M2016 diff_242400_251880# Vdd Vdd GND efet w=840 l=5760
+ ad=0 pd=0 as=0 ps=0 
M2017 Vdd Vdd Vdd GND efet w=600 l=360
+ ad=0 pd=0 as=0 ps=0 
M2018 diff_234480_257040# diff_242400_251880# diff_245520_249480# GND efet w=1440 l=720
+ ad=0 pd=0 as=6.3792e+06 ps=13920 
M2019 diff_241440_260160# diff_234480_257040# GND GND efet w=11220 l=660
+ ad=0 pd=0 as=0 ps=0 
M2020 Vdd Vdd Vdd GND efet w=420 l=900
+ ad=0 pd=0 as=0 ps=0 
M2021 diff_245520_249480# Vdd Vdd GND efet w=1080 l=2820
+ ad=0 pd=0 as=0 ps=0 
M2022 Vdd diff_189240_66360# diff_54840_246000# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M2023 diff_214320_243960# diff_213360_145800# diff_66360_247080# GND efet w=2160 l=720
+ ad=2.6064e+06 pd=7440 as=0 ps=0 
M2024 GND diff_211800_247200# diff_214320_243960# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2025 Vdd diff_222480_158400# diff_66360_247080# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2026 o2 diff_237480_243480# Vdd GND efet w=20700 l=660
+ ad=3.91536e+07 pd=69840 as=0 ps=0 
M2027 diff_214320_240720# diff_213360_145800# diff_66480_239280# GND efet w=2160 l=720
+ ad=2.592e+06 pd=7680 as=0 ps=0 
M2028 diff_54840_239280# diff_208200_149640# diff_204120_238680# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6208e+06 ps=7440 
M2029 diff_211800_238680# diff_211080_145800# diff_54840_239280# GND efet w=840 l=720
+ ad=2.592e+06 pd=7680 as=0 ps=0 
M2030 diff_54840_231960# diff_208200_149640# diff_204120_232920# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6352e+06 ps=7440 
M2031 diff_211800_233040# diff_211080_145800# diff_54840_231960# GND efet w=840 l=720
+ ad=2.592e+06 pd=7680 as=0 ps=0 
M2032 diff_66480_232800# diff_204600_144480# diff_205200_230160# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2033 diff_200520_226560# diff_199440_146040# diff_66480_225120# GND efet w=2040 l=720
+ ad=2.6064e+06 pd=7680 as=0 ps=0 
M2034 diff_54840_225240# diff_194400_149640# diff_190320_224640# GND efet w=840 l=720
+ ad=0 pd=0 as=2.664e+06 ps=7680 
M2035 diff_198000_224520# diff_197280_145800# diff_54840_225240# GND efet w=840 l=720
+ ad=2.5776e+06 pd=7680 as=0 ps=0 
M2036 diff_54840_217800# diff_194400_149640# diff_190320_218760# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6352e+06 ps=7440 
M2037 diff_198000_219000# diff_197280_145800# diff_54840_217800# GND efet w=720 l=720
+ ad=2.6064e+06 pd=7680 as=0 ps=0 
M2038 diff_66480_218640# diff_190800_144240# diff_191400_216000# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2039 diff_186720_212400# diff_185640_145800# diff_66480_210960# GND efet w=2160 l=720
+ ad=2.6064e+06 pd=7440 as=0 ps=0 
M2040 diff_54840_210960# diff_180600_149640# diff_176520_210960# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6496e+06 ps=7920 
M2041 diff_184320_210360# diff_183480_145800# diff_54840_210960# GND efet w=900 l=840
+ ad=2.6064e+06 pd=7680 as=0 ps=0 
M2042 diff_54840_203640# diff_180600_149640# diff_176640_204480# GND efet w=960 l=720
+ ad=0 pd=0 as=2.7072e+06 ps=7680 
M2043 diff_184320_204720# diff_183480_145800# diff_54840_203640# GND efet w=960 l=720
+ ad=2.6208e+06 pd=7680 as=0 ps=0 
M2044 diff_66480_204480# diff_177000_144360# diff_177600_201840# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2045 diff_173040_198120# diff_171960_145800# diff_66480_196680# GND efet w=2100 l=900
+ ad=2.376e+06 pd=7440 as=0 ps=0 
M2046 diff_54840_196800# diff_166800_149760# diff_162840_196200# GND efet w=840 l=720
+ ad=0 pd=0 as=2.4048e+06 ps=7440 
M2047 diff_170520_196200# diff_169680_145800# diff_54840_196800# GND efet w=840 l=720
+ ad=2.3904e+06 pd=7440 as=0 ps=0 
M2048 diff_54840_189360# diff_166800_149760# diff_162840_190320# GND efet w=840 l=720
+ ad=0 pd=0 as=2.52e+06 ps=7440 
M2049 diff_170520_190440# diff_169680_145800# diff_54840_189360# GND efet w=840 l=720
+ ad=2.664e+06 pd=7920 as=0 ps=0 
M2050 diff_66480_190200# diff_163320_144240# diff_163800_187560# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2051 diff_159240_183840# diff_158160_145800# diff_66480_182520# GND efet w=2160 l=720
+ ad=2.4048e+06 pd=7440 as=0 ps=0 
M2052 diff_66480_182520# diff_163320_144240# diff_163800_183360# GND efet w=2700 l=720
+ ad=0 pd=0 as=2.5632e+06 ps=8640 
M2053 diff_54840_182640# diff_153120_145800# diff_149040_181920# GND efet w=900 l=780
+ ad=0 pd=0 as=2.664e+06 ps=7440 
M2054 diff_156720_181920# diff_155880_145800# diff_54840_182640# GND efet w=960 l=840
+ ad=2.664e+06 pd=7440 as=0 ps=0 
M2055 diff_54840_175200# diff_153120_145800# diff_149040_176160# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6208e+06 ps=7440 
M2056 diff_156720_176400# diff_155880_145800# diff_54840_175200# GND efet w=840 l=720
+ ad=2.6496e+06 pd=7440 as=0 ps=0 
M2057 diff_66480_176040# diff_149520_144360# diff_150120_173400# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2058 diff_145440_169680# diff_144360_145800# diff_66480_168360# GND efet w=2040 l=720
+ ad=2.6208e+06 pd=7440 as=0 ps=0 
M2059 diff_54840_168480# diff_139320_149640# diff_135360_167760# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6928e+06 ps=7680 
M2060 diff_143040_167760# diff_142200_145800# diff_54840_168480# GND efet w=900 l=780
+ ad=2.5344e+06 pd=7200 as=0 ps=0 
M2061 diff_54840_161040# diff_139320_149640# diff_135360_162000# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6496e+06 ps=7440 
M2062 diff_143040_162120# diff_142200_145800# diff_54840_161040# GND efet w=840 l=720
+ ad=2.5344e+06 pd=7200 as=0 ps=0 
M2063 diff_66480_162000# diff_135720_144480# diff_136320_159240# GND efet w=2160 l=840
+ ad=0 pd=0 as=0 ps=0 
M2064 diff_131760_155520# diff_130680_145800# diff_66480_154320# GND efet w=2160 l=720
+ ad=2.3616e+06 pd=7440 as=0 ps=0 
M2065 diff_54840_154320# diff_125640_145800# diff_121560_153720# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6928e+06 ps=7920 
M2066 diff_129240_153600# diff_128400_145800# diff_54840_154320# GND efet w=840 l=720
+ ad=2.5776e+06 pd=7680 as=0 ps=0 
M2067 GND diff_129240_153600# diff_131760_155520# GND efet w=2280 l=840
+ ad=0 pd=0 as=0 ps=0 
M2068 diff_136320_155160# diff_135360_153720# GND GND efet w=2280 l=720
+ ad=2.3184e+06 pd=7200 as=0 ps=0 
M2069 diff_66480_154320# diff_135720_144480# diff_136320_155160# GND efet w=2160 l=840
+ ad=0 pd=0 as=0 ps=0 
M2070 GND diff_143040_167760# diff_145440_169680# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2071 diff_150120_169200# diff_149040_167760# GND GND efet w=2280 l=840
+ ad=2.3328e+06 pd=7440 as=0 ps=0 
M2072 diff_66480_168360# diff_149520_144360# diff_150120_169200# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M2073 diff_145440_158880# diff_144360_145800# diff_66480_162000# GND efet w=2160 l=720
+ ad=2.6208e+06 pd=7440 as=0 ps=0 
M2074 GND diff_143040_162120# diff_145440_158880# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2075 diff_150120_159240# diff_149040_162000# GND GND efet w=2280 l=840
+ ad=2.3328e+06 pd=7200 as=0 ps=0 
M2076 GND diff_156720_181920# diff_159240_183840# GND efet w=2340 l=900
+ ad=0 pd=0 as=0 ps=0 
M2077 diff_163800_183360# diff_162840_181920# GND GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M2078 GND diff_170520_196200# diff_173040_198120# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2079 diff_177600_197640# diff_176640_196080# GND GND efet w=2280 l=720
+ ad=2.3616e+06 pd=7440 as=0 ps=0 
M2080 diff_66480_196680# diff_177000_144360# diff_177600_197640# GND efet w=2100 l=780
+ ad=0 pd=0 as=0 ps=0 
M2081 diff_173040_187200# diff_171960_145800# diff_66480_190200# GND efet w=2160 l=840
+ ad=2.448e+06 pd=7440 as=0 ps=0 
M2082 GND diff_170520_190440# diff_173040_187200# GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M2083 diff_177600_187560# diff_176520_190440# GND GND efet w=2400 l=720
+ ad=2.4624e+06 pd=7440 as=0 ps=0 
M2084 GND diff_184320_210360# diff_186720_212400# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2085 diff_191400_211920# diff_190320_210360# GND GND efet w=2280 l=720
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M2086 diff_66480_210960# diff_190800_144240# diff_191400_211920# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2087 diff_186720_201480# diff_185640_145800# diff_66480_204480# GND efet w=2160 l=720
+ ad=2.6208e+06 pd=7680 as=0 ps=0 
M2088 GND diff_184320_204720# diff_186720_201480# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2089 diff_191400_201840# diff_190320_204480# GND GND efet w=2280 l=720
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M2090 diff_54840_210960# diff_194400_149640# diff_190320_210360# GND efet w=720 l=720
+ ad=0 pd=0 as=2.6928e+06 ps=7680 
M2091 GND diff_198000_224520# diff_200520_226560# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2092 diff_205200_225960# diff_204120_224640# GND GND efet w=2460 l=780
+ ad=2.3184e+06 pd=7200 as=0 ps=0 
M2093 diff_66480_225120# diff_204600_144480# diff_205200_225960# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M2094 diff_200520_215760# diff_199440_146040# diff_66480_218640# GND efet w=2040 l=720
+ ad=2.5488e+06 pd=7440 as=0 ps=0 
M2095 GND diff_198000_219000# diff_200520_215760# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2096 diff_205200_216000# diff_204120_218760# GND GND efet w=2280 l=780
+ ad=2.2464e+06 pd=6960 as=0 ps=0 
M2097 GND diff_211800_238680# diff_214320_240720# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2098 diff_245520_249480# diff_241440_260160# GND GND efet w=2520 l=720
+ ad=0 pd=0 as=0 ps=0 
M2099 o2 diff_241440_260160# GND GND efet w=19680 l=600
+ ad=0 pd=0 as=0 ps=0 
M2100 Vdd diff_222480_158400# diff_66480_239280# GND efet w=1440 l=840
+ ad=0 pd=0 as=0 ps=0 
M2101 Vdd diff_189240_66360# diff_54840_239280# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2102 diff_237480_243480# diff_237480_243480# diff_237480_243480# GND efet w=180 l=360
+ ad=9.8064e+06 pd=16800 as=0 ps=0 
M2103 diff_237480_243480# diff_237480_243480# diff_237480_243480# GND efet w=240 l=240
+ ad=0 pd=0 as=0 ps=0 
M2104 diff_237480_243480# Vdd Vdd GND efet w=1080 l=1920
+ ad=0 pd=0 as=0 ps=0 
M2105 GND diff_241440_260160# diff_237480_243480# GND efet w=4980 l=660
+ ad=0 pd=0 as=0 ps=0 
M2106 Vdd diff_189240_66360# diff_54840_231960# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M2107 diff_214320_229800# diff_213360_145800# diff_66480_232800# GND efet w=2160 l=720
+ ad=2.6208e+06 pd=7680 as=0 ps=0 
M2108 GND diff_211800_233040# diff_214320_229800# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2109 Vdd diff_222480_158400# diff_66480_232800# GND efet w=1440 l=660
+ ad=0 pd=0 as=0 ps=0 
M2110 diff_214320_226560# diff_213360_145800# diff_66480_225120# GND efet w=2040 l=720
+ ad=2.52e+06 pd=7680 as=0 ps=0 
M2111 diff_54840_225240# diff_208200_149640# diff_204120_224640# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6064e+06 ps=7440 
M2112 diff_211800_224520# diff_211080_145800# diff_54840_225240# GND efet w=840 l=720
+ ad=2.5776e+06 pd=7440 as=0 ps=0 
M2113 diff_54840_217800# diff_208200_149640# diff_204120_218760# GND efet w=720 l=720
+ ad=0 pd=0 as=2.6208e+06 ps=7440 
M2114 diff_211800_219000# diff_211080_145800# diff_54840_217800# GND efet w=720 l=720
+ ad=2.5632e+06 pd=7680 as=0 ps=0 
M2115 diff_66480_218640# diff_204600_144480# diff_205200_216000# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M2116 diff_200520_212400# diff_199440_146040# diff_66480_210960# GND efet w=2160 l=720
+ ad=2.592e+06 pd=7440 as=0 ps=0 
M2117 diff_198000_210480# diff_197280_145800# diff_54840_210960# GND efet w=720 l=720
+ ad=2.6496e+06 pd=7920 as=0 ps=0 
M2118 diff_54840_203640# diff_194400_149640# diff_190320_204480# GND efet w=960 l=720
+ ad=0 pd=0 as=2.7216e+06 ps=7680 
M2119 diff_198000_204720# diff_197280_145800# diff_54840_203640# GND efet w=840 l=720
+ ad=2.5776e+06 pd=7440 as=0 ps=0 
M2120 diff_66480_204480# diff_190800_144240# diff_191400_201840# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2121 diff_186720_198240# diff_185640_145800# diff_66480_196680# GND efet w=2040 l=720
+ ad=2.6208e+06 pd=7680 as=0 ps=0 
M2122 diff_54840_196800# diff_180600_149640# diff_176640_196080# GND efet w=840 l=720
+ ad=0 pd=0 as=2.592e+06 ps=8160 
M2123 diff_184320_196200# diff_183480_145800# diff_54840_196800# GND efet w=840 l=720
+ ad=2.4768e+06 pd=7920 as=0 ps=0 
M2124 diff_54840_189360# diff_180600_149640# diff_176520_190440# GND efet w=840 l=720
+ ad=0 pd=0 as=2.5488e+06 ps=7920 
M2125 diff_184320_190560# diff_183480_145800# diff_54840_189360# GND efet w=1020 l=780
+ ad=2.5488e+06 pd=7920 as=0 ps=0 
M2126 diff_66480_190200# diff_177000_144360# diff_177600_187560# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2127 diff_173040_183840# diff_171960_145800# diff_66480_182520# GND efet w=2160 l=840
+ ad=2.4192e+06 pd=7440 as=0 ps=0 
M2128 diff_54840_182640# diff_166800_149760# diff_162840_181920# GND efet w=960 l=720
+ ad=0 pd=0 as=2.5632e+06 ps=7440 
M2129 diff_170520_181920# diff_169680_145800# diff_54840_182640# GND efet w=960 l=720
+ ad=2.592e+06 pd=7680 as=0 ps=0 
M2130 GND diff_170520_181920# diff_173040_183840# GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M2131 diff_177600_183360# diff_176520_182280# GND GND efet w=2400 l=720
+ ad=2.4192e+06 pd=7440 as=0 ps=0 
M2132 diff_66480_182520# diff_177000_144360# diff_177600_183360# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2133 diff_54840_175200# diff_166800_149760# diff_162840_176040# GND efet w=720 l=780
+ ad=0 pd=0 as=2.5344e+06 ps=7680 
M2134 diff_170520_176400# diff_169680_145800# diff_54840_175200# GND efet w=780 l=780
+ ad=2.5632e+06 pd=7680 as=0 ps=0 
M2135 diff_159240_173040# diff_158160_145800# diff_66480_176040# GND efet w=2160 l=720
+ ad=2.376e+06 pd=7440 as=0 ps=0 
M2136 GND diff_156720_176400# diff_159240_173040# GND efet w=2280 l=840
+ ad=0 pd=0 as=0 ps=0 
M2137 diff_163800_173400# diff_162840_176040# GND GND efet w=2280 l=720
+ ad=2.448e+06 pd=8160 as=0 ps=0 
M2138 diff_66480_176040# diff_163320_144240# diff_163800_173400# GND efet w=2460 l=780
+ ad=0 pd=0 as=0 ps=0 
M2139 diff_159240_169680# diff_158160_145800# diff_66480_168360# GND efet w=2040 l=720
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M2140 diff_54840_168480# diff_153120_145800# diff_149040_167760# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6352e+06 ps=7440 
M2141 diff_156720_167760# diff_155880_145800# diff_54840_168480# GND efet w=840 l=720
+ ad=2.664e+06 pd=7440 as=0 ps=0 
M2142 diff_54840_161040# diff_153120_145800# diff_149040_162000# GND efet w=840 l=840
+ ad=0 pd=0 as=2.6496e+06 ps=7920 
M2143 diff_156720_162120# diff_155880_145800# diff_54840_161040# GND efet w=840 l=720
+ ad=2.52e+06 pd=7440 as=0 ps=0 
M2144 diff_66480_162000# diff_149520_144360# diff_150120_159240# GND efet w=2100 l=840
+ ad=0 pd=0 as=0 ps=0 
M2145 diff_145440_155640# diff_144360_145800# diff_66480_154320# GND efet w=2400 l=840
+ ad=2.5488e+06 pd=7920 as=0 ps=0 
M2146 diff_54840_154320# diff_139320_149640# diff_135360_153720# GND efet w=840 l=720
+ ad=0 pd=0 as=2.664e+06 ps=7440 
M2147 diff_143040_153600# diff_142200_145800# diff_54840_154320# GND efet w=840 l=720
+ ad=2.5344e+06 pd=7200 as=0 ps=0 
M2148 GND diff_143040_153600# diff_145440_155640# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2149 diff_150120_155160# diff_149040_153720# GND GND efet w=2160 l=840
+ ad=2.3184e+06 pd=7680 as=0 ps=0 
M2150 diff_66480_154320# diff_149520_144360# diff_150120_155160# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2151 GND diff_156720_167760# diff_159240_169680# GND efet w=2280 l=840
+ ad=0 pd=0 as=0 ps=0 
M2152 diff_163800_169200# diff_162840_167760# GND GND efet w=2280 l=720
+ ad=2.3616e+06 pd=7440 as=0 ps=0 
M2153 diff_66480_168360# diff_163320_144240# diff_163800_169200# GND efet w=2040 l=840
+ ad=0 pd=0 as=0 ps=0 
M2154 diff_173040_173040# diff_171960_145800# diff_66480_176040# GND efet w=2160 l=840
+ ad=2.2032e+06 pd=7440 as=0 ps=0 
M2155 GND diff_170520_176400# diff_173040_173040# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2156 diff_177600_173400# diff_176520_176280# GND GND efet w=2280 l=720
+ ad=2.376e+06 pd=7440 as=0 ps=0 
M2157 GND diff_184320_196200# diff_186720_198240# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2158 diff_191400_197640# diff_190320_196200# GND GND efet w=2280 l=720
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M2159 diff_66480_196680# diff_190800_144240# diff_191400_197640# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M2160 diff_186720_187200# diff_185640_145800# diff_66480_190200# GND efet w=2160 l=720
+ ad=2.6928e+06 pd=7680 as=0 ps=0 
M2161 GND diff_184320_190560# diff_186720_187200# GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M2162 diff_191400_187560# diff_190320_190320# GND GND efet w=2400 l=720
+ ad=2.448e+06 pd=7440 as=0 ps=0 
M2163 GND diff_198000_210480# diff_200520_212400# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2164 diff_205200_211920# diff_204120_210360# GND GND efet w=2580 l=780
+ ad=2.3184e+06 pd=7200 as=0 ps=0 
M2165 diff_66480_210960# diff_204600_144480# diff_205200_211920# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2166 diff_200520_201480# diff_199440_146040# diff_66480_204480# GND efet w=2160 l=720
+ ad=2.6208e+06 pd=7680 as=0 ps=0 
M2167 GND diff_198000_204720# diff_200520_201480# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2168 diff_205200_201840# diff_204120_204480# GND GND efet w=2340 l=780
+ ad=2.3184e+06 pd=7200 as=0 ps=0 
M2169 GND diff_211800_224520# diff_214320_226560# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2170 Vdd diff_222480_158400# diff_66480_225120# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M2171 Vdd diff_189240_66360# diff_54840_225240# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2172 Vdd diff_189240_66360# diff_54840_217800# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M2173 GND diff_211800_219000# diff_214320_215760# GND efet w=2220 l=780
+ ad=0 pd=0 as=2.52e+06 ps=7440 
M2174 diff_214320_215760# diff_213360_145800# diff_66480_218640# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M2175 Vdd diff_222480_158400# diff_66480_218640# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M2176 diff_241680_195480# Vdd Vdd GND efet w=1080 l=1920
+ ad=1.31616e+07 pd=26160 as=0 ps=0 
M2177 diff_232560_214800# clk2 diff_23160_135720# GND efet w=1920 l=720
+ ad=2.6928e+06 pd=7680 as=0 ps=0 
M2178 diff_214320_212400# diff_213360_145800# diff_66480_210960# GND efet w=2160 l=720
+ ad=2.6064e+06 pd=7440 as=0 ps=0 
M2179 diff_54840_210960# diff_208200_149640# diff_204120_210360# GND efet w=720 l=720
+ ad=0 pd=0 as=2.592e+06 ps=7440 
M2180 diff_211800_210480# diff_211080_145800# diff_54840_210960# GND efet w=720 l=720
+ ad=2.592e+06 pd=7680 as=0 ps=0 
M2181 diff_54840_203640# diff_208200_149640# diff_204120_204480# GND efet w=840 l=840
+ ad=0 pd=0 as=2.592e+06 ps=7440 
M2182 diff_211800_204840# diff_211080_145800# diff_54840_203640# GND efet w=720 l=720
+ ad=2.6064e+06 pd=7680 as=0 ps=0 
M2183 diff_66480_204480# diff_204600_144480# diff_205200_201840# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2184 diff_200520_198240# diff_199440_146040# diff_66480_196680# GND efet w=2040 l=720
+ ad=2.592e+06 pd=7440 as=0 ps=0 
M2185 diff_54840_196800# diff_194400_149640# diff_190320_196200# GND efet w=840 l=720
+ ad=0 pd=0 as=2.5632e+06 ps=7680 
M2186 diff_198000_196200# diff_197280_145800# diff_54840_196800# GND efet w=840 l=720
+ ad=2.592e+06 pd=7680 as=0 ps=0 
M2187 diff_54840_189360# diff_194400_149640# diff_190320_190320# GND efet w=840 l=720
+ ad=0 pd=0 as=2.664e+06 ps=7680 
M2188 diff_198000_190560# diff_197280_145800# diff_54840_189360# GND efet w=840 l=720
+ ad=2.6208e+06 pd=7920 as=0 ps=0 
M2189 diff_66480_190200# diff_190800_144240# diff_191400_187560# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2190 diff_186720_183960# diff_185640_145800# diff_66480_182520# GND efet w=2160 l=720
+ ad=2.6352e+06 pd=7440 as=0 ps=0 
M2191 diff_54840_182640# diff_180600_149640# diff_176520_182280# GND efet w=960 l=720
+ ad=0 pd=0 as=2.6496e+06 ps=7920 
M2192 diff_184320_181920# diff_183480_145800# diff_54840_182640# GND efet w=1140 l=780
+ ad=2.5776e+06 pd=7680 as=0 ps=0 
M2193 diff_54840_175200# diff_180600_149640# diff_176520_176280# GND efet w=840 l=720
+ ad=0 pd=0 as=2.7072e+06 ps=7680 
M2194 diff_184320_176280# diff_183480_145800# diff_54840_175200# GND efet w=840 l=840
+ ad=2.6208e+06 pd=7680 as=0 ps=0 
M2195 diff_66480_176040# diff_177000_144360# diff_177600_173400# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2196 diff_173040_169680# diff_171960_145800# diff_66480_168360# GND efet w=2040 l=840
+ ad=2.3616e+06 pd=7440 as=0 ps=0 
M2197 diff_66480_168360# diff_177000_144360# diff_177600_169200# GND efet w=2160 l=840
+ ad=0 pd=0 as=2.376e+06 ps=7200 
M2198 diff_54840_168480# diff_166800_149760# diff_162840_167760# GND efet w=840 l=720
+ ad=0 pd=0 as=2.5344e+06 ps=7680 
M2199 diff_170520_167760# diff_169680_145800# diff_54840_168480# GND efet w=840 l=720
+ ad=2.5488e+06 pd=7440 as=0 ps=0 
M2200 diff_159240_158880# diff_158160_145800# diff_66480_162000# GND efet w=2100 l=780
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M2201 GND diff_156720_162120# diff_159240_158880# GND efet w=2280 l=840
+ ad=0 pd=0 as=0 ps=0 
M2202 diff_163800_159240# diff_162840_162000# GND GND efet w=2280 l=720
+ ad=2.3904e+06 pd=7440 as=0 ps=0 
M2203 GND diff_170520_167760# diff_173040_169680# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2204 diff_177600_169200# diff_176520_167880# GND GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2205 diff_54840_161040# diff_166800_149760# diff_162840_162000# GND efet w=840 l=720
+ ad=0 pd=0 as=2.5056e+06 ps=7440 
M2206 diff_170520_162120# diff_169680_145800# diff_54840_161040# GND efet w=840 l=720
+ ad=2.4336e+06 pd=7680 as=0 ps=0 
M2207 diff_66480_162000# diff_163320_144240# diff_163800_159240# GND efet w=2220 l=900
+ ad=0 pd=0 as=0 ps=0 
M2208 diff_159240_155520# diff_158160_145800# diff_66480_154320# GND efet w=2040 l=720
+ ad=2.3472e+06 pd=7440 as=0 ps=0 
M2209 diff_66480_154320# diff_163320_144240# diff_163800_155040# GND efet w=2100 l=780
+ ad=0 pd=0 as=2.3904e+06 ps=7680 
M2210 diff_54840_154320# diff_153120_145800# diff_149040_153720# GND efet w=960 l=720
+ ad=0 pd=0 as=2.7216e+06 ps=7920 
M2211 diff_156720_153600# diff_155880_145800# diff_54840_154320# GND efet w=960 l=720
+ ad=2.6784e+06 pd=7440 as=0 ps=0 
M2212 GND diff_156720_153600# diff_159240_155520# GND efet w=2280 l=840
+ ad=0 pd=0 as=0 ps=0 
M2213 diff_163800_155040# diff_162840_153720# GND GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2214 diff_173040_158880# diff_171960_145800# diff_66480_162000# GND efet w=2100 l=900
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M2215 GND diff_170520_162120# diff_173040_158880# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2216 diff_177600_159240# diff_176520_162120# GND GND efet w=2280 l=720
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M2217 GND diff_184320_181920# diff_186720_183960# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2218 diff_191400_183480# diff_190320_182040# GND GND efet w=2280 l=720
+ ad=2.3616e+06 pd=7200 as=0 ps=0 
M2219 diff_66480_182520# diff_190800_144240# diff_191400_183480# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2220 diff_186720_173040# diff_185640_145800# diff_66480_176040# GND efet w=2160 l=720
+ ad=2.6352e+06 pd=7680 as=0 ps=0 
M2221 GND diff_184320_176280# diff_186720_173040# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2222 diff_191400_173400# diff_190320_176160# GND GND efet w=2280 l=720
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M2223 GND diff_198000_196200# diff_200520_198240# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2224 diff_205200_197640# diff_204120_196200# GND GND efet w=2280 l=720
+ ad=2.3328e+06 pd=7440 as=0 ps=0 
M2225 diff_66480_196680# diff_204600_144480# diff_205200_197640# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M2226 diff_200520_187320# diff_199440_146040# diff_66480_190200# GND efet w=2040 l=720
+ ad=2.6208e+06 pd=7440 as=0 ps=0 
M2227 GND diff_198000_190560# diff_200520_187320# GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M2228 diff_205200_187560# diff_204120_190320# GND GND efet w=2280 l=720
+ ad=2.2464e+06 pd=6960 as=0 ps=0 
M2229 GND diff_211800_210480# diff_214320_212400# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2230 diff_234480_214080# diff_207480_277200# diff_232560_214800# GND efet w=1920 l=720
+ ad=1.69488e+07 pd=33600 as=0 ps=0 
M2231 Vdd diff_222480_158400# diff_66480_210960# GND efet w=1560 l=720
+ ad=0 pd=0 as=0 ps=0 
M2232 GND diff_207480_277200# diff_242520_208920# GND efet w=1440 l=660
+ ad=0 pd=0 as=3.4704e+06 ps=7920 
M2233 GND diff_207720_290040# diff_234480_214080# GND efet w=2760 l=600
+ ad=0 pd=0 as=0 ps=0 
M2234 Vdd diff_189240_66360# diff_54840_210960# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2235 diff_242520_208920# Vdd Vdd GND efet w=900 l=5820
+ ad=0 pd=0 as=0 ps=0 
M2236 Vdd Vdd Vdd GND efet w=600 l=360
+ ad=0 pd=0 as=0 ps=0 
M2237 Vdd diff_189240_66360# diff_54840_203640# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2238 diff_234480_214080# diff_242520_208920# diff_245520_206640# GND efet w=1440 l=600
+ ad=0 pd=0 as=6.5952e+06 ps=14640 
M2239 diff_241680_195480# diff_234480_214080# GND GND efet w=11160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2240 Vdd Vdd Vdd GND efet w=480 l=840
+ ad=0 pd=0 as=0 ps=0 
M2241 diff_245520_206640# Vdd Vdd GND efet w=960 l=3060
+ ad=0 pd=0 as=0 ps=0 
M2242 diff_214320_201480# diff_213360_145800# diff_66480_204480# GND efet w=2160 l=720
+ ad=2.6208e+06 pd=7680 as=0 ps=0 
M2243 GND diff_211800_204840# diff_214320_201480# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2244 Vdd diff_222480_158400# diff_66480_204480# GND efet w=1560 l=600
+ ad=0 pd=0 as=0 ps=0 
M2245 diff_214320_198240# diff_213360_145800# diff_66480_196680# GND efet w=2040 l=720
+ ad=2.592e+06 pd=7680 as=0 ps=0 
M2246 diff_54840_196800# diff_208200_149640# diff_204120_196200# GND efet w=840 l=720
+ ad=0 pd=0 as=2.52e+06 ps=7440 
M2247 diff_211800_196200# diff_211080_145800# diff_54840_196800# GND efet w=840 l=720
+ ad=2.52e+06 pd=7920 as=0 ps=0 
M2248 diff_54840_189360# diff_208200_149640# diff_204120_190320# GND efet w=840 l=720
+ ad=0 pd=0 as=2.5632e+06 ps=7440 
M2249 diff_211800_190560# diff_211080_145800# diff_54840_189360# GND efet w=840 l=720
+ ad=2.5344e+06 pd=7680 as=0 ps=0 
M2250 diff_66480_190200# diff_204600_144480# diff_205200_187560# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M2251 diff_200520_183960# diff_199440_146040# diff_66480_182520# GND efet w=2160 l=720
+ ad=2.6064e+06 pd=7440 as=0 ps=0 
M2252 diff_54840_182640# diff_194400_149640# diff_190320_182040# GND efet w=840 l=720
+ ad=0 pd=0 as=2.664e+06 ps=7440 
M2253 diff_198000_182040# diff_197280_145800# diff_54840_182640# GND efet w=960 l=720
+ ad=2.4768e+06 pd=7680 as=0 ps=0 
M2254 diff_54840_175200# diff_194400_149640# diff_190320_176160# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6208e+06 ps=7440 
M2255 diff_198000_176400# diff_197280_145800# diff_54840_175200# GND efet w=840 l=720
+ ad=2.5632e+06 pd=7680 as=0 ps=0 
M2256 diff_66480_176040# diff_190800_144240# diff_191400_173400# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2257 diff_186720_169800# diff_185640_145800# diff_66480_168360# GND efet w=2040 l=720
+ ad=2.6208e+06 pd=7680 as=0 ps=0 
M2258 diff_54840_168480# diff_180600_149640# diff_176520_167880# GND efet w=840 l=720
+ ad=0 pd=0 as=2.664e+06 ps=7440 
M2259 diff_184320_167760# diff_183480_145800# diff_54840_168480# GND efet w=840 l=840
+ ad=2.5632e+06 pd=7680 as=0 ps=0 
M2260 diff_54840_161040# diff_180600_149640# diff_176520_162120# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6496e+06 ps=7440 
M2261 diff_184320_162120# diff_183480_145800# diff_54840_161040# GND efet w=840 l=840
+ ad=2.4912e+06 pd=7920 as=0 ps=0 
M2262 diff_66480_162000# diff_177000_144360# diff_177600_159240# GND efet w=2100 l=780
+ ad=0 pd=0 as=0 ps=0 
M2263 diff_173040_155520# diff_171960_145800# diff_66480_154320# GND efet w=2040 l=840
+ ad=2.3616e+06 pd=7440 as=0 ps=0 
M2264 diff_66480_154320# diff_177000_144360# diff_177600_155040# GND efet w=2040 l=840
+ ad=0 pd=0 as=2.376e+06 ps=7200 
M2265 diff_54840_154320# diff_166800_149760# diff_162840_153720# GND efet w=960 l=720
+ ad=0 pd=0 as=2.5488e+06 ps=7440 
M2266 diff_170520_153600# diff_169680_145800# diff_54840_154320# GND efet w=960 l=720
+ ad=2.5488e+06 pd=7440 as=0 ps=0 
M2267 GND diff_170520_153600# diff_173040_155520# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2268 diff_177600_155040# diff_176520_153840# GND GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2269 GND diff_184320_167760# diff_186720_169800# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2270 diff_191400_169200# diff_190320_167880# GND GND efet w=2520 l=840
+ ad=2.376e+06 pd=7200 as=0 ps=0 
M2271 diff_66480_168360# diff_190800_144240# diff_191400_169200# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M2272 diff_186720_158880# diff_185640_145800# diff_66480_162000# GND efet w=2100 l=780
+ ad=2.6064e+06 pd=7440 as=0 ps=0 
M2273 GND diff_184320_162120# diff_186720_158880# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2274 diff_191400_159240# diff_190320_162000# GND GND efet w=2340 l=780
+ ad=2.3472e+06 pd=7200 as=0 ps=0 
M2275 GND diff_198000_182040# diff_200520_183960# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2276 diff_205200_183480# diff_204120_182040# GND GND efet w=2280 l=720
+ ad=2.3184e+06 pd=7200 as=0 ps=0 
M2277 diff_66480_182520# diff_204600_144480# diff_205200_183480# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2278 diff_200520_173040# diff_199440_146040# diff_66480_176040# GND efet w=2160 l=720
+ ad=2.6208e+06 pd=7680 as=0 ps=0 
M2279 GND diff_198000_176400# diff_200520_173040# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2280 diff_205200_173400# diff_204120_176160# GND GND efet w=2520 l=780
+ ad=2.3184e+06 pd=7200 as=0 ps=0 
M2281 GND diff_211800_196200# diff_214320_198240# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2282 o3 diff_237480_200400# Vdd GND efet w=20640 l=720
+ ad=4.03632e+07 pd=68400 as=0 ps=0 
M2283 diff_245520_206640# diff_241680_195480# GND GND efet w=2760 l=720
+ ad=0 pd=0 as=0 ps=0 
M2284 o3 diff_241680_195480# GND GND efet w=19380 l=660
+ ad=0 pd=0 as=0 ps=0 
M2285 Vdd diff_222480_158400# diff_66480_196680# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M2286 Vdd diff_189240_66360# diff_54840_196800# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M2287 diff_237480_200400# diff_237480_200400# diff_237480_200400# GND efet w=180 l=300
+ ad=9.8496e+06 pd=17280 as=0 ps=0 
M2288 diff_237480_200400# Vdd Vdd GND efet w=1200 l=1860
+ ad=0 pd=0 as=0 ps=0 
M2289 diff_237480_200400# diff_237480_200400# diff_237480_200400# GND efet w=240 l=240
+ ad=0 pd=0 as=0 ps=0 
M2290 diff_237480_200400# diff_241680_195480# GND GND efet w=5100 l=660
+ ad=0 pd=0 as=0 ps=0 
M2291 Vdd diff_189240_66360# diff_54840_189360# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2292 diff_214320_187320# diff_213360_145800# diff_66480_190200# GND efet w=2040 l=720
+ ad=2.592e+06 pd=7440 as=0 ps=0 
M2293 GND diff_211800_190560# diff_214320_187320# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2294 Vdd diff_222480_158400# diff_66480_190200# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M2295 diff_214320_183960# diff_213360_145800# diff_66480_182520# GND efet w=2100 l=780
+ ad=2.6064e+06 pd=7440 as=0 ps=0 
M2296 diff_54840_182640# diff_208200_149640# diff_204120_182040# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6208e+06 ps=7440 
M2297 diff_211800_182040# diff_211080_145800# diff_54840_182640# GND efet w=840 l=720
+ ad=2.6784e+06 pd=7920 as=0 ps=0 
M2298 diff_54840_175200# diff_208200_149640# diff_204120_176160# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6784e+06 ps=7680 
M2299 diff_211800_176400# diff_211080_145800# diff_54840_175200# GND efet w=840 l=720
+ ad=2.5632e+06 pd=7680 as=0 ps=0 
M2300 diff_66480_176040# diff_204600_144480# diff_205200_173400# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2301 diff_200520_169800# diff_199440_146040# diff_66480_168360# GND efet w=2040 l=720
+ ad=2.592e+06 pd=7680 as=0 ps=0 
M2302 diff_54840_168480# diff_194400_149640# diff_190320_167880# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6496e+06 ps=7440 
M2303 diff_198000_167760# diff_197280_145800# diff_54840_168480# GND efet w=840 l=720
+ ad=2.6496e+06 pd=7920 as=0 ps=0 
M2304 diff_54840_161040# diff_194400_149640# diff_190320_162000# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6208e+06 ps=7440 
M2305 diff_198000_162120# diff_197280_145800# diff_54840_161040# GND efet w=840 l=720
+ ad=2.5776e+06 pd=7680 as=0 ps=0 
M2306 diff_66480_162000# diff_190800_144240# diff_191400_159240# GND efet w=2100 l=780
+ ad=0 pd=0 as=0 ps=0 
M2307 diff_186720_155640# diff_185640_145800# diff_66480_154320# GND efet w=2040 l=720
+ ad=2.6064e+06 pd=7680 as=0 ps=0 
M2308 diff_54840_154320# diff_180600_149640# diff_176520_153840# GND efet w=960 l=720
+ ad=0 pd=0 as=2.6784e+06 ps=7440 
M2309 diff_184320_153600# diff_183480_145800# diff_54840_154320# GND efet w=1080 l=840
+ ad=2.5488e+06 pd=7200 as=0 ps=0 
M2310 GND diff_184320_153600# diff_186720_155640# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2311 diff_191400_155040# diff_190320_153720# GND GND efet w=2280 l=840
+ ad=2.3328e+06 pd=7200 as=0 ps=0 
M2312 diff_66480_154320# diff_190800_144240# diff_191400_155040# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M2313 GND diff_198000_167760# diff_200520_169800# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2314 diff_205200_169200# diff_204120_167880# GND GND efet w=2340 l=780
+ ad=2.304e+06 pd=7200 as=0 ps=0 
M2315 diff_66480_168360# diff_204600_144480# diff_205200_169200# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M2316 diff_200520_158880# diff_199440_146040# diff_66480_162000# GND efet w=2100 l=780
+ ad=2.592e+06 pd=7440 as=0 ps=0 
M2317 GND diff_198000_162120# diff_200520_158880# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2318 diff_205200_159240# diff_204120_162000# GND GND efet w=2280 l=840
+ ad=2.3184e+06 pd=7200 as=0 ps=0 
M2319 GND diff_211800_182040# diff_214320_183960# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2320 Vdd diff_222480_158400# diff_66480_182520# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2321 Vdd diff_189240_66360# diff_54840_182640# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M2322 Vdd diff_189240_66360# diff_54840_175200# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2323 diff_214320_173040# diff_213360_145800# diff_66480_176040# GND efet w=2160 l=720
+ ad=2.664e+06 pd=7680 as=0 ps=0 
M2324 GND diff_211800_176400# diff_214320_173040# GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M2325 Vdd diff_222480_158400# diff_66480_176040# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2326 GND diff_179280_17640# diff_207720_290040# GND efet w=5280 l=600
+ ad=0 pd=0 as=7.4736e+06 ps=14880 
M2327 diff_214320_169800# diff_213360_145800# diff_66480_168360# GND efet w=2160 l=720
+ ad=2.592e+06 pd=7440 as=0 ps=0 
M2328 diff_54840_168480# diff_208200_149640# diff_204120_167880# GND efet w=960 l=720
+ ad=0 pd=0 as=2.6064e+06 ps=7680 
M2329 diff_211800_167760# diff_211080_145800# diff_54840_168480# GND efet w=840 l=720
+ ad=2.6496e+06 pd=7920 as=0 ps=0 
M2330 diff_54840_161040# diff_208200_149640# diff_204120_162000# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6208e+06 ps=7680 
M2331 diff_211800_162120# diff_211080_145800# diff_54840_161040# GND efet w=840 l=720
+ ad=2.6496e+06 pd=7440 as=0 ps=0 
M2332 diff_66480_162000# diff_204600_144480# diff_205200_159240# GND efet w=2100 l=780
+ ad=0 pd=0 as=0 ps=0 
M2333 diff_200520_155640# diff_199440_146040# diff_66480_154320# GND efet w=2040 l=720
+ ad=2.4912e+06 pd=7200 as=0 ps=0 
M2334 diff_54840_154320# diff_194400_149640# diff_190320_153720# GND efet w=840 l=720
+ ad=0 pd=0 as=2.6784e+06 ps=7440 
M2335 diff_198000_153720# diff_197280_145800# diff_54840_154320# GND efet w=840 l=720
+ ad=2.6352e+06 pd=7440 as=0 ps=0 
M2336 GND diff_198000_153720# diff_200520_155640# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2337 diff_205200_155160# diff_204120_153720# GND GND efet w=2160 l=840
+ ad=2.232e+06 pd=6960 as=0 ps=0 
M2338 diff_66480_154320# diff_204600_144480# diff_205200_155160# GND efet w=2040 l=720
+ ad=0 pd=0 as=0 ps=0 
M2339 GND diff_211800_167760# diff_214320_169800# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2340 Vdd diff_222480_158400# diff_66480_168360# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M2341 Vdd diff_189240_66360# diff_54840_168480# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2342 diff_207720_290040# Vdd Vdd GND efet w=1080 l=1860
+ ad=0 pd=0 as=0 ps=0 
M2343 Vdd diff_189240_66360# diff_54840_161040# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M2344 diff_222480_158400# diff_228240_160560# diff_222480_158400# GND efet w=3060 l=3180
+ ad=1.47888e+07 pd=26400 as=0 ps=0 
M2345 diff_214320_158880# diff_213360_145800# diff_66480_162000# GND efet w=2160 l=720
+ ad=2.5632e+06 pd=7440 as=0 ps=0 
M2346 GND diff_211800_162120# diff_214320_158880# GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2347 Vdd diff_222480_158400# diff_66480_162000# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M2348 diff_228240_160560# Vdd Vdd GND efet w=840 l=720
+ ad=2.6064e+06 pd=8160 as=0 ps=0 
M2349 diff_228240_160560# diff_228240_160560# diff_228240_160560# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M2350 diff_228240_160560# diff_228240_160560# diff_228240_160560# GND efet w=240 l=720
+ ad=0 pd=0 as=0 ps=0 
M2351 GND diff_234240_153840# diff_222480_158400# GND efet w=7440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2352 diff_222480_158400# diff_228240_160560# Vdd GND efet w=1080 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2353 diff_222480_158400# diff_222480_158400# diff_222480_158400# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M2354 diff_222480_158400# diff_222480_158400# diff_222480_158400# GND efet w=420 l=420
+ ad=0 pd=0 as=0 ps=0 
M2355 diff_214320_155640# diff_213360_145800# diff_66480_154320# GND efet w=2160 l=720
+ ad=2.5632e+06 pd=7440 as=0 ps=0 
M2356 diff_54840_154320# diff_208200_149640# diff_204120_153720# GND efet w=840 l=720
+ ad=0 pd=0 as=2.4768e+06 ps=7440 
M2357 diff_211800_153720# diff_211080_145800# diff_54840_154320# GND efet w=720 l=840
+ ad=2.6064e+06 pd=7440 as=0 ps=0 
M2358 GND diff_211800_153720# diff_214320_155640# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2359 Vdd diff_222480_158400# diff_66480_154320# GND efet w=1380 l=720
+ ad=0 pd=0 as=0 ps=0 
M2360 diff_234240_153840# Vdd Vdd GND efet w=1080 l=1920
+ ad=9.5184e+06 pd=17280 as=0 ps=0 
M2361 Vdd diff_189240_66360# diff_54840_154320# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M2362 diff_234240_153840# clk1 diff_234600_150240# GND efet w=7320 l=720
+ ad=0 pd=0 as=1.29024e+07 ps=26640 
M2363 GND diff_234000_148080# diff_234600_150240# GND efet w=11400 l=720
+ ad=0 pd=0 as=0 ps=0 
M2364 GND diff_79800_142440# diff_80760_144360# GND efet w=1800 l=840
+ ad=0 pd=0 as=5.4144e+06 ps=12000 
M2365 GND diff_79800_142440# diff_84360_149760# GND efet w=1200 l=840
+ ad=0 pd=0 as=2.016e+06 ps=5760 
M2366 GND diff_86760_147600# diff_87240_145800# GND efet w=1200 l=840
+ ad=0 pd=0 as=2.016e+06 ps=5760 
M2367 GND diff_86760_147600# diff_89400_145800# GND efet w=1800 l=840
+ ad=0 pd=0 as=4.9536e+06 ps=11760 
M2368 Vdd Vdd diff_43680_161280# GND efet w=1080 l=3840
+ ad=0 pd=0 as=1.09296e+07 ps=26880 
M2369 Vdd Vdd diff_33120_151080# GND efet w=1080 l=4200
+ ad=0 pd=0 as=1.54368e+07 ps=34800 
M2370 diff_32760_140400# diff_32760_140400# diff_32760_140400# GND efet w=360 l=360
+ ad=1.32912e+07 pd=28080 as=0 ps=0 
M2371 Vdd Vdd diff_32760_140400# GND efet w=1080 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2372 diff_32760_140400# diff_32760_140400# diff_32760_140400# GND efet w=180 l=360
+ ad=0 pd=0 as=0 ps=0 
M2373 diff_42600_159120# diff_71400_87600# Vdd GND efet w=3840 l=720
+ ad=2.58912e+07 pd=43920 as=0 ps=0 
M2374 GND diff_73200_137520# diff_42600_159120# GND efet w=3840 l=720
+ ad=0 pd=0 as=0 ps=0 
M2375 diff_82080_142080# diff_81000_115920# diff_80760_144360# GND efet w=3180 l=1020
+ ad=9.1728e+07 pd=228960 as=0 ps=0 
M2376 diff_84360_149760# diff_81000_115920# diff_84480_143520# GND efet w=1260 l=780
+ ad=0 pd=0 as=8.83584e+07 ps=200640 
M2377 diff_87240_145800# diff_86760_145200# diff_84480_143520# GND efet w=1260 l=780
+ ad=0 pd=0 as=0 ps=0 
M2378 diff_89400_145800# diff_86760_145200# diff_82080_142080# GND efet w=3180 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2379 diff_32640_245760# diff_32640_245760# diff_32640_245760# GND efet w=420 l=420
+ ad=1.11312e+07 pd=28800 as=0 ps=0 
M2380 Vdd Vdd diff_32640_245760# GND efet w=1080 l=3840
+ ad=0 pd=0 as=0 ps=0 
M2381 diff_32640_245760# diff_32640_245760# diff_32640_245760# GND efet w=360 l=360
+ ad=0 pd=0 as=0 ps=0 
M2382 GND diff_16320_124440# diff_23160_135720# GND efet w=3900 l=660
+ ad=0 pd=0 as=0 ps=0 
M2383 diff_73200_137520# Vdd Vdd GND efet w=840 l=3840
+ ad=4.8816e+06 pd=10800 as=0 ps=0 
M2384 GND diff_93720_142200# diff_94560_144240# GND efet w=1800 l=840
+ ad=0 pd=0 as=5.1264e+06 ps=11760 
M2385 GND diff_93720_142200# diff_98160_145800# GND efet w=1320 l=840
+ ad=0 pd=0 as=2.2176e+06 ps=6000 
M2386 GND diff_100560_147600# diff_100920_145800# GND efet w=1320 l=840
+ ad=0 pd=0 as=2.016e+06 ps=5760 
M2387 GND diff_100560_147600# diff_103200_145800# GND efet w=1680 l=840
+ ad=0 pd=0 as=4.9104e+06 ps=11760 
M2388 diff_82080_142080# diff_94680_112080# diff_94560_144240# GND efet w=3180 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2389 diff_98160_145800# diff_94680_112080# diff_84480_143520# GND efet w=1440 l=840
+ ad=0 pd=0 as=0 ps=0 
M2390 diff_100920_145800# diff_100560_145080# diff_84480_143520# GND efet w=1260 l=780
+ ad=0 pd=0 as=0 ps=0 
M2391 diff_103200_145800# diff_100560_145080# diff_82080_142080# GND efet w=3120 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2392 GND diff_107520_138960# diff_108240_144360# GND efet w=1800 l=840
+ ad=0 pd=0 as=5.3568e+06 ps=12240 
M2393 GND diff_107520_138960# diff_111840_149760# GND efet w=1200 l=840
+ ad=0 pd=0 as=2.016e+06 ps=5760 
M2394 GND diff_114240_147600# diff_114720_145800# GND efet w=1200 l=840
+ ad=0 pd=0 as=2.016e+06 ps=5760 
M2395 GND diff_114240_147600# diff_116880_145800# GND efet w=1800 l=840
+ ad=0 pd=0 as=5.1984e+06 ps=12000 
M2396 diff_82080_142080# diff_108480_116040# diff_108240_144360# GND efet w=3420 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2397 diff_111840_149760# diff_108480_116040# diff_84480_143520# GND efet w=1260 l=780
+ ad=0 pd=0 as=0 ps=0 
M2398 diff_114720_145800# diff_114240_145080# diff_84480_143520# GND efet w=1260 l=780
+ ad=0 pd=0 as=0 ps=0 
M2399 diff_116880_145800# diff_114240_145080# diff_82080_142080# GND efet w=3180 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2400 GND diff_121200_142200# diff_122040_144240# GND efet w=1680 l=840
+ ad=0 pd=0 as=5.0544e+06 ps=11760 
M2401 GND diff_121200_142200# diff_125640_145800# GND efet w=1320 l=840
+ ad=0 pd=0 as=2.2176e+06 ps=6000 
M2402 GND diff_128040_147600# diff_128400_145800# GND efet w=1320 l=840
+ ad=0 pd=0 as=2.2176e+06 ps=6000 
M2403 GND diff_128040_147600# diff_130680_145800# GND efet w=1680 l=840
+ ad=0 pd=0 as=5.0112e+06 ps=11760 
M2404 diff_82080_142080# diff_122160_115920# diff_122040_144240# GND efet w=3060 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2405 diff_125640_145800# diff_122160_115920# diff_84480_143520# GND efet w=1380 l=780
+ ad=0 pd=0 as=0 ps=0 
M2406 diff_128400_145800# diff_128040_145080# diff_84480_143520# GND efet w=1500 l=780
+ ad=0 pd=0 as=0 ps=0 
M2407 diff_130680_145800# diff_128040_145080# diff_82080_142080# GND efet w=3120 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2408 GND diff_135000_138960# diff_135720_144480# GND efet w=1800 l=840
+ ad=0 pd=0 as=5.1984e+06 ps=12000 
M2409 GND diff_135000_138960# diff_139320_149640# GND efet w=1200 l=840
+ ad=0 pd=0 as=2.016e+06 ps=5760 
M2410 GND diff_141720_147600# diff_142200_145800# GND efet w=1200 l=840
+ ad=0 pd=0 as=2.016e+06 ps=5760 
M2411 GND diff_141720_147600# diff_144360_145800# GND efet w=1800 l=840
+ ad=0 pd=0 as=5.2272e+06 ps=12000 
M2412 diff_82080_142080# diff_135960_115920# diff_135720_144480# GND efet w=3300 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2413 diff_139320_149640# diff_135960_115920# diff_84480_143520# GND efet w=1260 l=780
+ ad=0 pd=0 as=0 ps=0 
M2414 diff_142200_145800# diff_141720_145080# diff_84480_143520# GND efet w=1260 l=780
+ ad=0 pd=0 as=0 ps=0 
M2415 diff_144360_145800# diff_141720_145080# diff_82080_142080# GND efet w=3180 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2416 GND diff_148680_142200# diff_149520_144360# GND efet w=1800 l=840
+ ad=0 pd=0 as=5.04e+06 ps=12000 
M2417 GND diff_148680_142200# diff_153120_145800# GND efet w=1320 l=780
+ ad=0 pd=0 as=2.2176e+06 ps=6000 
M2418 GND diff_155520_147600# diff_155880_145800# GND efet w=1260 l=840
+ ad=0 pd=0 as=2.2176e+06 ps=6000 
M2419 GND diff_155520_147600# diff_158160_145800# GND efet w=1800 l=840
+ ad=0 pd=0 as=4.9968e+06 ps=11760 
M2420 diff_82080_142080# diff_149760_115920# diff_149520_144360# GND efet w=3180 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2421 diff_153120_145800# diff_149760_115920# diff_84480_143520# GND efet w=1380 l=780
+ ad=0 pd=0 as=0 ps=0 
M2422 diff_155880_145800# diff_155520_145080# diff_84480_143520# GND efet w=1380 l=780
+ ad=0 pd=0 as=0 ps=0 
M2423 diff_158160_145800# diff_155520_145080# diff_82080_142080# GND efet w=3240 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2424 GND diff_162480_139680# diff_163320_144240# GND efet w=1800 l=840
+ ad=0 pd=0 as=5.0112e+06 ps=11760 
M2425 GND diff_162480_139680# diff_166800_149760# GND efet w=1260 l=780
+ ad=0 pd=0 as=2.016e+06 ps=5760 
M2426 GND diff_169200_147600# diff_169680_145800# GND efet w=1200 l=840
+ ad=0 pd=0 as=2.016e+06 ps=5760 
M2427 diff_171960_145800# diff_169200_147600# GND GND efet w=1680 l=840
+ ad=5.0256e+06 pd=11760 as=0 ps=0 
M2428 diff_82080_142080# diff_163440_116040# diff_163320_144240# GND efet w=3300 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2429 diff_166800_149760# diff_163440_116040# diff_84480_143520# GND efet w=1260 l=780
+ ad=0 pd=0 as=0 ps=0 
M2430 diff_169680_145800# diff_169200_145080# diff_84480_143520# GND efet w=1260 l=780
+ ad=0 pd=0 as=0 ps=0 
M2431 diff_171960_145800# diff_169200_145080# diff_82080_142080# GND efet w=3180 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2432 GND diff_176160_142200# diff_177000_144360# GND efet w=1800 l=840
+ ad=0 pd=0 as=5.2128e+06 ps=12000 
M2433 GND diff_176160_142200# diff_180600_149640# GND efet w=1200 l=780
+ ad=0 pd=0 as=2.016e+06 ps=5760 
M2434 GND diff_183000_147600# diff_183480_145800# GND efet w=1200 l=840
+ ad=0 pd=0 as=2.016e+06 ps=5760 
M2435 GND diff_183000_147600# diff_185640_145800# GND efet w=1920 l=840
+ ad=0 pd=0 as=5.256e+06 ps=12240 
M2436 diff_82080_142080# diff_175920_112080# diff_177000_144360# GND efet w=3300 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2437 diff_180600_149640# diff_175920_112080# diff_84480_143520# GND efet w=1260 l=780
+ ad=0 pd=0 as=0 ps=0 
M2438 diff_183480_145800# diff_182040_114360# diff_84480_143520# GND efet w=1260 l=780
+ ad=0 pd=0 as=0 ps=0 
M2439 diff_185640_145800# diff_182040_114360# diff_82080_142080# GND efet w=3300 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2440 GND diff_189960_142200# diff_190800_144240# GND efet w=1980 l=780
+ ad=0 pd=0 as=5.1264e+06 ps=12720 
M2441 GND diff_189960_142200# diff_194400_149640# GND efet w=1200 l=720
+ ad=0 pd=0 as=2.16e+06 ps=6000 
M2442 GND diff_196800_147600# diff_197280_145800# GND efet w=1320 l=720
+ ad=0 pd=0 as=2.1312e+06 ps=6240 
M2443 diff_199440_146040# diff_196800_147600# GND GND efet w=1740 l=780
+ ad=5.2992e+06 pd=12240 as=0 ps=0 
M2444 diff_82080_142080# diff_189240_116040# diff_190800_144240# GND efet w=3120 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2445 diff_194400_149640# diff_189240_116040# diff_84480_143520# GND efet w=1200 l=720
+ ad=0 pd=0 as=0 ps=0 
M2446 diff_197280_145800# diff_196560_127680# diff_84480_143520# GND efet w=1260 l=780
+ ad=0 pd=0 as=0 ps=0 
M2447 diff_199440_146040# diff_196560_127680# diff_82080_142080# GND efet w=3120 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2448 GND diff_203760_142200# diff_204600_144480# GND efet w=1980 l=720
+ ad=0 pd=0 as=5.2416e+06 ps=12480 
M2449 GND diff_203760_142200# diff_208200_149640# GND efet w=1200 l=720
+ ad=0 pd=0 as=2.16e+06 ps=6000 
M2450 GND diff_210600_147600# diff_211080_145800# GND efet w=1200 l=720
+ ad=0 pd=0 as=2.16e+06 ps=6000 
M2451 diff_213360_145800# diff_210600_147600# GND GND efet w=1680 l=720
+ ad=5.2128e+06 pd=12000 as=0 ps=0 
M2452 diff_234000_148080# Vdd Vdd GND efet w=1080 l=2760
+ ad=9.216e+06 pd=21120 as=0 ps=0 
M2453 diff_234000_148080# diff_234000_148080# diff_234000_148080# GND efet w=240 l=480
+ ad=0 pd=0 as=0 ps=0 
M2454 diff_234000_148080# diff_234000_148080# diff_234000_148080# GND efet w=240 l=840
+ ad=0 pd=0 as=0 ps=0 
M2455 diff_82080_142080# diff_201120_122760# diff_204600_144480# GND efet w=3300 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2456 diff_208200_149640# diff_201120_122760# diff_84480_143520# GND efet w=1200 l=720
+ ad=0 pd=0 as=0 ps=0 
M2457 diff_211080_145800# diff_205320_118080# diff_84480_143520# GND efet w=1200 l=720
+ ad=0 pd=0 as=0 ps=0 
M2458 diff_213360_145800# diff_205320_118080# diff_82080_142080# GND efet w=3120 l=960
+ ad=0 pd=0 as=0 ps=0 
M2459 diff_79800_142440# diff_79800_142440# diff_79800_142440# GND efet w=480 l=720
+ ad=5.3712e+06 pd=14640 as=0 ps=0 
M2460 diff_79800_142440# diff_79800_142440# diff_79800_142440# GND efet w=600 l=360
+ ad=0 pd=0 as=0 ps=0 
M2461 GND diff_81000_115920# diff_79800_142440# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2462 diff_86760_147600# diff_86760_145200# GND GND efet w=1440 l=720
+ ad=5.04e+06 pd=14160 as=0 ps=0 
M2463 diff_86760_147600# diff_86760_147600# diff_86760_147600# GND efet w=480 l=720
+ ad=0 pd=0 as=0 ps=0 
M2464 diff_86760_147600# diff_86760_147600# diff_86760_147600# GND efet w=600 l=360
+ ad=0 pd=0 as=0 ps=0 
M2465 Vdd Vdd diff_79800_142440# GND efet w=720 l=3840
+ ad=0 pd=0 as=0 ps=0 
M2466 GND diff_71400_87600# diff_73200_137520# GND efet w=1920 l=720
+ ad=0 pd=0 as=0 ps=0 
M2467 d3 GND GND GND efet w=10320 l=840
+ ad=0 pd=0 as=0 ps=0 
M2468 diff_23160_135720# diff_17040_127440# Vdd GND efet w=3840 l=720
+ ad=0 pd=0 as=0 ps=0 
M2469 diff_81000_115920# diff_81000_115920# diff_81000_115920# GND efet w=300 l=300
+ ad=1.89216e+07 pd=47040 as=0 ps=0 
M2470 diff_33120_151080# diff_51600_133800# GND GND efet w=2520 l=720
+ ad=0 pd=0 as=0 ps=0 
M2471 diff_32640_245760# diff_51600_133800# GND GND efet w=2520 l=720
+ ad=0 pd=0 as=0 ps=0 
M2472 diff_17040_127440# diff_16320_124440# GND GND efet w=2280 l=720
+ ad=1.4112e+07 pd=27600 as=0 ps=0 
M2473 diff_17040_127440# diff_17040_127440# diff_17040_127440# GND efet w=240 l=240
+ ad=0 pd=0 as=0 ps=0 
M2474 diff_17040_127440# diff_17040_127440# diff_17040_127440# GND efet w=180 l=540
+ ad=0 pd=0 as=0 ps=0 
M2475 Vdd Vdd diff_17040_127440# GND efet w=840 l=3660
+ ad=0 pd=0 as=0 ps=0 
M2476 diff_81000_115920# diff_81000_115920# diff_81000_115920# GND efet w=240 l=480
+ ad=0 pd=0 as=0 ps=0 
M2477 diff_93720_142200# diff_93720_142200# diff_93720_142200# GND efet w=480 l=600
+ ad=5.2992e+06 pd=14160 as=0 ps=0 
M2478 diff_93720_142200# diff_93720_142200# diff_93720_142200# GND efet w=540 l=300
+ ad=0 pd=0 as=0 ps=0 
M2479 GND diff_94680_112080# diff_93720_142200# GND efet w=1440 l=840
+ ad=0 pd=0 as=0 ps=0 
M2480 diff_100560_147600# diff_100560_145080# GND GND efet w=1680 l=720
+ ad=5.1552e+06 pd=14640 as=0 ps=0 
M2481 diff_100560_147600# diff_100560_147600# diff_100560_147600# GND efet w=480 l=600
+ ad=0 pd=0 as=0 ps=0 
M2482 diff_100560_147600# diff_100560_147600# diff_100560_147600# GND efet w=540 l=300
+ ad=0 pd=0 as=0 ps=0 
M2483 Vdd Vdd diff_86760_147600# GND efet w=900 l=5040
+ ad=0 pd=0 as=0 ps=0 
M2484 diff_93720_142200# Vdd Vdd GND efet w=900 l=4560
+ ad=0 pd=0 as=0 ps=0 
M2485 diff_86760_145200# diff_86760_145200# diff_86760_145200# GND efet w=240 l=360
+ ad=1.95984e+07 pd=45600 as=0 ps=0 
M2486 diff_86760_145200# diff_86760_145200# diff_86760_145200# GND efet w=360 l=420
+ ad=0 pd=0 as=0 ps=0 
M2487 diff_94680_112080# diff_94680_112080# diff_94680_112080# GND efet w=300 l=300
+ ad=1.76976e+07 pd=49440 as=0 ps=0 
M2488 diff_94680_112080# diff_94680_112080# diff_94680_112080# GND efet w=240 l=600
+ ad=0 pd=0 as=0 ps=0 
M2489 diff_107520_138960# diff_107520_138960# diff_107520_138960# GND efet w=480 l=720
+ ad=5.4e+06 pd=14640 as=0 ps=0 
M2490 diff_107520_138960# diff_107520_138960# diff_107520_138960# GND efet w=600 l=360
+ ad=0 pd=0 as=0 ps=0 
M2491 GND diff_108480_116040# diff_107520_138960# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2492 diff_114240_147600# diff_114240_145080# GND GND efet w=1440 l=720
+ ad=5.1984e+06 pd=14400 as=0 ps=0 
M2493 diff_114240_147600# diff_114240_147600# diff_114240_147600# GND efet w=480 l=720
+ ad=0 pd=0 as=0 ps=0 
M2494 diff_121200_142200# diff_121200_142200# diff_121200_142200# GND efet w=480 l=720
+ ad=5.2272e+06 pd=14160 as=0 ps=0 
M2495 diff_114240_147600# diff_114240_147600# diff_114240_147600# GND efet w=600 l=360
+ ad=0 pd=0 as=0 ps=0 
M2496 Vdd Vdd diff_100560_147600# GND efet w=900 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2497 diff_107520_138960# Vdd Vdd GND efet w=900 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2498 diff_100560_145080# diff_100560_145080# diff_100560_145080# GND efet w=240 l=300
+ ad=1.89216e+07 pd=45360 as=0 ps=0 
M2499 diff_100560_145080# diff_100560_145080# diff_100560_145080# GND efet w=420 l=420
+ ad=0 pd=0 as=0 ps=0 
M2500 diff_108480_116040# diff_108480_116040# diff_108480_116040# GND efet w=360 l=360
+ ad=1.87488e+07 pd=47040 as=0 ps=0 
M2501 diff_108480_116040# diff_108480_116040# diff_108480_116040# GND efet w=240 l=480
+ ad=0 pd=0 as=0 ps=0 
M2502 GND diff_122160_115920# diff_121200_142200# GND efet w=1560 l=720
+ ad=0 pd=0 as=0 ps=0 
M2503 diff_121200_142200# diff_121200_142200# diff_121200_142200# GND efet w=540 l=300
+ ad=0 pd=0 as=0 ps=0 
M2504 diff_128040_147600# diff_128040_145080# GND GND efet w=1440 l=720
+ ad=5.2128e+06 pd=14400 as=0 ps=0 
M2505 diff_128040_147600# diff_128040_147600# diff_128040_147600# GND efet w=480 l=720
+ ad=0 pd=0 as=0 ps=0 
M2506 diff_128040_147600# diff_128040_147600# diff_128040_147600# GND efet w=600 l=360
+ ad=0 pd=0 as=0 ps=0 
M2507 diff_114240_147600# Vdd Vdd GND efet w=1020 l=4680
+ ad=0 pd=0 as=0 ps=0 
M2508 diff_121200_142200# Vdd Vdd GND efet w=1020 l=4740
+ ad=0 pd=0 as=0 ps=0 
M2509 diff_114240_145080# diff_114240_145080# diff_114240_145080# GND efet w=240 l=360
+ ad=1.91952e+07 pd=44400 as=0 ps=0 
M2510 diff_114240_145080# diff_114240_145080# diff_114240_145080# GND efet w=420 l=420
+ ad=0 pd=0 as=0 ps=0 
M2511 diff_122160_115920# diff_122160_115920# diff_122160_115920# GND efet w=300 l=300
+ ad=1.86192e+07 pd=47280 as=0 ps=0 
M2512 diff_122160_115920# diff_122160_115920# diff_122160_115920# GND efet w=300 l=600
+ ad=0 pd=0 as=0 ps=0 
M2513 diff_135000_138960# diff_135000_138960# diff_135000_138960# GND efet w=540 l=660
+ ad=5.328e+06 pd=15120 as=0 ps=0 
M2514 GND diff_135960_115920# diff_135000_138960# GND efet w=1740 l=780
+ ad=0 pd=0 as=0 ps=0 
M2515 diff_141720_147600# diff_141720_145080# GND GND efet w=1680 l=780
+ ad=5.256e+06 pd=14160 as=0 ps=0 
M2516 diff_141720_147600# diff_141720_147600# diff_141720_147600# GND efet w=480 l=600
+ ad=0 pd=0 as=0 ps=0 
M2517 diff_135000_138960# diff_135000_138960# diff_135000_138960# GND efet w=540 l=300
+ ad=0 pd=0 as=0 ps=0 
M2518 diff_141720_147600# diff_141720_147600# diff_141720_147600# GND efet w=540 l=300
+ ad=0 pd=0 as=0 ps=0 
M2519 Vdd Vdd diff_128040_147600# GND efet w=900 l=4680
+ ad=0 pd=0 as=0 ps=0 
M2520 diff_135000_138960# Vdd Vdd GND efet w=900 l=4560
+ ad=0 pd=0 as=0 ps=0 
M2521 diff_128040_145080# diff_128040_145080# diff_128040_145080# GND efet w=240 l=300
+ ad=1.87632e+07 pd=44880 as=0 ps=0 
M2522 diff_128040_145080# diff_128040_145080# diff_128040_145080# GND efet w=420 l=420
+ ad=0 pd=0 as=0 ps=0 
M2523 diff_135960_115920# diff_135960_115920# diff_135960_115920# GND efet w=240 l=360
+ ad=1.87632e+07 pd=46560 as=0 ps=0 
M2524 diff_135960_115920# diff_135960_115920# diff_135960_115920# GND efet w=240 l=480
+ ad=0 pd=0 as=0 ps=0 
M2525 diff_148680_142200# diff_148680_142200# diff_148680_142200# GND efet w=480 l=720
+ ad=5.184e+06 pd=14400 as=0 ps=0 
M2526 GND diff_149760_115920# diff_148680_142200# GND efet w=1560 l=720
+ ad=0 pd=0 as=0 ps=0 
M2527 diff_155520_147600# diff_155520_145080# GND GND efet w=1560 l=720
+ ad=5.1984e+06 pd=14400 as=0 ps=0 
M2528 diff_148680_142200# diff_148680_142200# diff_148680_142200# GND efet w=600 l=360
+ ad=0 pd=0 as=0 ps=0 
M2529 diff_155520_147600# diff_155520_147600# diff_155520_147600# GND efet w=480 l=720
+ ad=0 pd=0 as=0 ps=0 
M2530 diff_162480_139680# diff_162480_139680# diff_162480_139680# GND efet w=480 l=720
+ ad=5.2848e+06 pd=14640 as=0 ps=0 
M2531 diff_155520_147600# diff_155520_147600# diff_155520_147600# GND efet w=540 l=300
+ ad=0 pd=0 as=0 ps=0 
M2532 diff_162480_139680# diff_162480_139680# diff_162480_139680# GND efet w=540 l=300
+ ad=0 pd=0 as=0 ps=0 
M2533 GND diff_163440_116040# diff_162480_139680# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2534 diff_169200_147600# diff_169200_145080# GND GND efet w=1440 l=720
+ ad=5.2128e+06 pd=14400 as=0 ps=0 
M2535 diff_169200_147600# diff_169200_147600# diff_169200_147600# GND efet w=480 l=720
+ ad=0 pd=0 as=0 ps=0 
M2536 diff_169200_147600# diff_169200_147600# diff_169200_147600# GND efet w=600 l=360
+ ad=0 pd=0 as=0 ps=0 
M2537 Vdd Vdd diff_141720_147600# GND efet w=840 l=4740
+ ad=0 pd=0 as=0 ps=0 
M2538 diff_148680_142200# Vdd Vdd GND efet w=900 l=4860
+ ad=0 pd=0 as=0 ps=0 
M2539 diff_141720_145080# diff_141720_145080# diff_141720_145080# GND efet w=240 l=300
+ ad=1.93248e+07 pd=44400 as=0 ps=0 
M2540 diff_141720_145080# diff_141720_145080# diff_141720_145080# GND efet w=360 l=360
+ ad=0 pd=0 as=0 ps=0 
M2541 diff_149760_115920# diff_149760_115920# diff_149760_115920# GND efet w=300 l=300
+ ad=1.71504e+07 pd=42480 as=0 ps=0 
M2542 diff_149760_115920# diff_149760_115920# diff_149760_115920# GND efet w=240 l=360
+ ad=0 pd=0 as=0 ps=0 
M2543 Vdd Vdd diff_155520_147600# GND efet w=900 l=4740
+ ad=0 pd=0 as=0 ps=0 
M2544 diff_162480_139680# Vdd Vdd GND efet w=780 l=4680
+ ad=0 pd=0 as=0 ps=0 
M2545 diff_155520_145080# diff_155520_145080# diff_155520_145080# GND efet w=240 l=300
+ ad=1.94112e+07 pd=52320 as=0 ps=0 
M2546 diff_155520_145080# diff_155520_145080# diff_155520_145080# GND efet w=360 l=480
+ ad=0 pd=0 as=0 ps=0 
M2547 diff_163440_116040# diff_163440_116040# diff_163440_116040# GND efet w=300 l=300
+ ad=1.89792e+07 pd=47760 as=0 ps=0 
M2548 diff_163440_116040# diff_163440_116040# diff_163440_116040# GND efet w=240 l=480
+ ad=0 pd=0 as=0 ps=0 
M2549 diff_176160_142200# diff_176160_142200# diff_176160_142200# GND efet w=480 l=600
+ ad=5.2848e+06 pd=14160 as=0 ps=0 
M2550 diff_176160_142200# diff_176160_142200# diff_176160_142200# GND efet w=540 l=300
+ ad=0 pd=0 as=0 ps=0 
M2551 GND diff_175920_112080# diff_176160_142200# GND efet w=1440 l=840
+ ad=0 pd=0 as=0 ps=0 
M2552 diff_183000_147600# diff_182040_114360# GND GND efet w=1620 l=780
+ ad=5.2992e+06 pd=14160 as=0 ps=0 
M2553 diff_183000_147600# diff_183000_147600# diff_183000_147600# GND efet w=480 l=600
+ ad=0 pd=0 as=0 ps=0 
M2554 diff_183000_147600# diff_183000_147600# diff_183000_147600# GND efet w=540 l=300
+ ad=0 pd=0 as=0 ps=0 
M2555 Vdd Vdd diff_169200_147600# GND efet w=900 l=4680
+ ad=0 pd=0 as=0 ps=0 
M2556 diff_176160_142200# Vdd Vdd GND efet w=840 l=4620
+ ad=0 pd=0 as=0 ps=0 
M2557 diff_169200_145080# diff_169200_145080# diff_169200_145080# GND efet w=180 l=420
+ ad=2.12688e+07 pd=53040 as=0 ps=0 
M2558 diff_169200_145080# diff_169200_145080# diff_169200_145080# GND efet w=360 l=360
+ ad=0 pd=0 as=0 ps=0 
M2559 diff_175920_112080# diff_175920_112080# diff_175920_112080# GND efet w=360 l=480
+ ad=2.21328e+07 pd=55920 as=0 ps=0 
M2560 diff_175920_112080# diff_175920_112080# diff_175920_112080# GND efet w=180 l=420
+ ad=0 pd=0 as=0 ps=0 
M2561 diff_189960_142200# diff_189960_142200# diff_189960_142200# GND efet w=480 l=720
+ ad=5.4e+06 pd=14640 as=0 ps=0 
M2562 diff_189960_142200# diff_189960_142200# diff_189960_142200# GND efet w=600 l=360
+ ad=0 pd=0 as=0 ps=0 
M2563 GND diff_189240_116040# diff_189960_142200# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2564 diff_196800_147600# diff_196560_127680# GND GND efet w=1440 l=720
+ ad=5.2272e+06 pd=14400 as=0 ps=0 
M2565 diff_196800_147600# diff_196800_147600# diff_196800_147600# GND efet w=480 l=600
+ ad=0 pd=0 as=0 ps=0 
M2566 diff_203760_142200# diff_203760_142200# diff_203760_142200# GND efet w=480 l=720
+ ad=5.2272e+06 pd=14400 as=0 ps=0 
M2567 diff_196800_147600# diff_196800_147600# diff_196800_147600# GND efet w=540 l=300
+ ad=0 pd=0 as=0 ps=0 
M2568 Vdd Vdd diff_183000_147600# GND efet w=900 l=4740
+ ad=0 pd=0 as=0 ps=0 
M2569 diff_189960_142200# Vdd Vdd GND efet w=900 l=4680
+ ad=0 pd=0 as=0 ps=0 
M2570 diff_182040_114360# diff_182040_114360# diff_182040_114360# GND efet w=180 l=240
+ ad=2.35872e+07 pd=60960 as=0 ps=0 
M2571 diff_182040_114360# diff_182040_114360# diff_182040_114360# GND efet w=360 l=360
+ ad=0 pd=0 as=0 ps=0 
M2572 diff_81000_115920# diff_82440_133920# GND GND efet w=1560 l=780
+ ad=0 pd=0 as=0 ps=0 
M2573 diff_86760_145200# diff_82440_133920# GND GND efet w=1680 l=840
+ ad=0 pd=0 as=0 ps=0 
M2574 diff_94680_112080# diff_82440_133920# GND GND efet w=1620 l=900
+ ad=0 pd=0 as=0 ps=0 
M2575 diff_100560_145080# diff_82440_133920# GND GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2576 diff_108480_116040# diff_82440_133920# GND GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2577 diff_114240_145080# diff_82440_133920# GND GND efet w=1620 l=900
+ ad=0 pd=0 as=0 ps=0 
M2578 diff_122160_115920# diff_82440_133920# GND GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2579 diff_128040_145080# diff_82440_133920# GND GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2580 diff_135960_115920# diff_130200_104880# GND GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2581 diff_141720_145080# diff_130200_104880# GND GND efet w=1620 l=900
+ ad=0 pd=0 as=0 ps=0 
M2582 diff_149760_115920# diff_130200_104880# GND GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2583 diff_155520_145080# diff_130200_104880# GND GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2584 diff_163440_116040# diff_130200_104880# GND GND efet w=1680 l=840
+ ad=0 pd=0 as=0 ps=0 
M2585 diff_169200_145080# diff_130200_104880# GND GND efet w=1560 l=720
+ ad=0 pd=0 as=0 ps=0 
M2586 diff_175920_112080# diff_130200_104880# GND GND efet w=1680 l=720
+ ad=0 pd=0 as=0 ps=0 
M2587 diff_182040_114360# diff_130200_104880# GND GND efet w=1560 l=720
+ ad=0 pd=0 as=0 ps=0 
M2588 diff_203760_142200# diff_203760_142200# diff_203760_142200# GND efet w=600 l=360
+ ad=0 pd=0 as=0 ps=0 
M2589 GND diff_201120_122760# diff_203760_142200# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2590 diff_234000_148080# diff_26880_44640# diff_234960_145080# GND efet w=6900 l=660
+ ad=0 pd=0 as=9.72e+06 ps=20160 
M2591 diff_234960_145080# diff_78360_22440# GND GND efet w=7200 l=660
+ ad=0 pd=0 as=0 ps=0 
M2592 diff_210600_147600# diff_210600_147600# diff_210600_147600# GND efet w=120 l=240
+ ad=6.048e+06 pd=19440 as=0 ps=0 
M2593 Vdd Vdd diff_196800_147600# GND efet w=780 l=4620
+ ad=0 pd=0 as=0 ps=0 
M2594 diff_203760_142200# Vdd Vdd GND efet w=900 l=4680
+ ad=0 pd=0 as=0 ps=0 
M2595 diff_210600_147600# diff_210600_147600# diff_210600_147600# GND efet w=240 l=240
+ ad=0 pd=0 as=0 ps=0 
M2596 diff_82080_142080# diff_231000_136440# Vdd GND efet w=3840 l=840
+ ad=0 pd=0 as=0 ps=0 
M2597 diff_210600_147600# diff_205320_118080# GND GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2598 Vdd Vdd diff_210600_147600# GND efet w=660 l=4500
+ ad=0 pd=0 as=0 ps=0 
M2599 GND diff_233520_124920# diff_82080_142080# GND efet w=4380 l=600
+ ad=0 pd=0 as=0 ps=0 
M2600 GND diff_233520_124920# diff_231000_136440# GND efet w=4080 l=720
+ ad=0 pd=0 as=1.5552e+07 ps=38400 
M2601 GND diff_51600_131160# diff_32760_140400# GND efet w=2520 l=720
+ ad=0 pd=0 as=0 ps=0 
M2602 GND diff_51600_131160# diff_43680_161280# GND efet w=2520 l=720
+ ad=0 pd=0 as=0 ps=0 
M2603 diff_52320_146760# diff_21960_94200# Vdd GND efet w=2940 l=720
+ ad=1.49328e+07 pd=25680 as=0 ps=0 
M2604 GND diff_73200_125280# diff_52320_146760# GND efet w=2760 l=720
+ ad=0 pd=0 as=0 ps=0 
M2605 GND diff_82200_132000# diff_81000_115920# GND efet w=1680 l=840
+ ad=0 pd=0 as=0 ps=0 
M2606 diff_86760_145200# diff_82200_132000# GND GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2607 GND diff_82200_132000# diff_94680_112080# GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2608 GND diff_82200_132000# diff_100560_145080# GND efet w=1740 l=780
+ ad=0 pd=0 as=0 ps=0 
M2609 GND diff_82200_132000# diff_135960_115920# GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2610 diff_141720_145080# diff_82200_132000# GND GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2611 GND diff_82200_132000# diff_149760_115920# GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2612 diff_155520_145080# diff_82200_132000# GND GND efet w=1620 l=780
+ ad=0 pd=0 as=0 ps=0 
M2613 diff_205320_118080# diff_207600_131160# diff_205320_118080# GND efet w=8400 l=360
+ ad=2.01888e+07 pd=57600 as=0 ps=0 
M2614 diff_108480_116040# diff_109680_129600# GND GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2615 diff_114240_145080# diff_109680_129600# GND GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2616 diff_122160_115920# diff_109680_129600# GND GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2617 diff_128040_145080# diff_109680_129600# GND GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2618 diff_163440_116040# diff_109680_129600# GND GND efet w=1620 l=780
+ ad=0 pd=0 as=0 ps=0 
M2619 diff_169200_145080# diff_109680_129600# GND GND efet w=1740 l=780
+ ad=0 pd=0 as=0 ps=0 
M2620 diff_175920_112080# diff_109680_129600# GND GND efet w=1560 l=720
+ ad=0 pd=0 as=0 ps=0 
M2621 diff_182040_114360# diff_109680_129600# GND GND efet w=1560 l=780
+ ad=0 pd=0 as=0 ps=0 
M2622 Vdd diff_207600_131160# diff_205320_118080# GND efet w=840 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2623 diff_207600_131160# diff_207600_131160# diff_207600_131160# GND efet w=120 l=360
+ ad=2.4912e+06 pd=7920 as=0 ps=0 
M2624 diff_207600_131160# diff_207600_131160# diff_207600_131160# GND efet w=240 l=420
+ ad=0 pd=0 as=0 ps=0 
M2625 Vdd Vdd diff_207600_131160# GND efet w=840 l=720
+ ad=0 pd=0 as=0 ps=0 
M2626 diff_231000_136440# diff_230520_127080# Vdd GND efet w=960 l=1920
+ ad=0 pd=0 as=0 ps=0 
M2627 diff_189240_116040# diff_190200_129480# GND GND efet w=2040 l=780
+ ad=1.83888e+07 pd=38880 as=0 ps=0 
M2628 diff_32760_140400# diff_51600_126720# GND GND efet w=2520 l=720
+ ad=0 pd=0 as=0 ps=0 
M2629 diff_32640_245760# diff_51600_126720# GND GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M2630 diff_17040_127440# diff_13200_279960# GND GND efet w=3600 l=720
+ ad=0 pd=0 as=0 ps=0 
M2631 diff_16320_124440# diff_16320_124440# diff_16320_124440# GND efet w=240 l=720
+ ad=1.20384e+07 pd=28800 as=0 ps=0 
M2632 diff_16320_124440# diff_16320_124440# diff_16320_124440# GND efet w=240 l=600
+ ad=0 pd=0 as=0 ps=0 
M2633 diff_16320_124440# d3 GND GND efet w=5520 l=720
+ ad=0 pd=0 as=0 ps=0 
M2634 diff_73200_125280# Vdd Vdd GND efet w=840 l=3900
+ ad=3.7584e+06 pd=9120 as=0 ps=0 
M2635 diff_81000_115920# diff_82200_127320# GND GND efet w=1740 l=780
+ ad=0 pd=0 as=0 ps=0 
M2636 diff_86760_145200# diff_82200_127320# GND GND efet w=1560 l=720
+ ad=0 pd=0 as=0 ps=0 
M2637 GND diff_82200_127320# diff_108480_116040# GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2638 GND diff_21960_94200# diff_73200_125280# GND efet w=1980 l=900
+ ad=0 pd=0 as=0 ps=0 
M2639 diff_114240_145080# diff_82200_127320# GND GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2640 diff_205320_118080# diff_190200_129480# GND GND efet w=1920 l=840
+ ad=0 pd=0 as=0 ps=0 
M2641 diff_231000_136440# diff_230520_127080# diff_231000_136440# GND efet w=5400 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2642 GND diff_51600_124080# diff_33120_151080# GND efet w=2520 l=720
+ ad=0 pd=0 as=0 ps=0 
M2643 GND diff_51600_124080# diff_43680_161280# GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M2644 diff_135960_115920# diff_82200_127320# GND GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2645 diff_141720_145080# diff_82200_127320# GND GND efet w=1740 l=780
+ ad=0 pd=0 as=0 ps=0 
M2646 GND diff_82200_127320# diff_163440_116040# GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2647 diff_169200_145080# diff_82200_127320# GND GND efet w=1740 l=780
+ ad=0 pd=0 as=0 ps=0 
M2648 diff_230520_127080# diff_230520_127080# diff_230520_127080# GND efet w=300 l=300
+ ad=2.4624e+06 pd=7920 as=0 ps=0 
M2649 diff_230520_127080# diff_230520_127080# diff_230520_127080# GND efet w=180 l=780
+ ad=0 pd=0 as=0 ps=0 
M2650 diff_196560_127680# diff_196080_127080# GND GND efet w=3120 l=720
+ ad=1.81008e+07 pd=48480 as=0 ps=0 
M2651 GND diff_196080_127080# diff_201120_122760# GND efet w=3240 l=720
+ ad=0 pd=0 as=2.09808e+07 ps=50160 
M2652 diff_230520_127080# Vdd Vdd GND efet w=900 l=840
+ ad=0 pd=0 as=0 ps=0 
M2653 GND diff_84000_102000# diff_94680_112080# GND efet w=1560 l=780
+ ad=0 pd=0 as=0 ps=0 
M2654 GND diff_84000_102000# diff_100560_145080# GND efet w=1680 l=840
+ ad=0 pd=0 as=0 ps=0 
M2655 diff_122160_115920# diff_84000_102000# GND GND efet w=1620 l=900
+ ad=0 pd=0 as=0 ps=0 
M2656 diff_128040_145080# diff_84000_102000# GND GND efet w=1620 l=900
+ ad=0 pd=0 as=0 ps=0 
M2657 GND diff_84000_102000# diff_149760_115920# GND efet w=1680 l=960
+ ad=0 pd=0 as=0 ps=0 
M2658 diff_155520_145080# diff_84000_102000# GND GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2659 diff_175920_112080# diff_84000_102000# GND GND efet w=1620 l=720
+ ad=0 pd=0 as=0 ps=0 
M2660 diff_182040_114360# diff_84000_102000# GND GND efet w=1560 l=720
+ ad=0 pd=0 as=0 ps=0 
M2661 GND diff_13200_279960# diff_16320_124440# GND efet w=3600 l=720
+ ad=0 pd=0 as=0 ps=0 
M2662 diff_81000_115920# diff_82200_122760# GND GND efet w=1560 l=720
+ ad=0 pd=0 as=0 ps=0 
M2663 diff_108480_116040# diff_82200_122760# GND GND efet w=1740 l=780
+ ad=0 pd=0 as=0 ps=0 
M2664 diff_94680_112080# diff_82200_122760# GND GND efet w=1560 l=720
+ ad=0 pd=0 as=0 ps=0 
M2665 GND diff_82200_122760# diff_122160_115920# GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2666 GND diff_197400_124560# diff_196560_127680# GND efet w=1920 l=840
+ ad=0 pd=0 as=0 ps=0 
M2667 GND diff_197400_124560# diff_205320_118080# GND efet w=1920 l=840
+ ad=0 pd=0 as=0 ps=0 
M2668 diff_233520_124920# Vdd Vdd GND efet w=1080 l=1920
+ ad=8.856e+06 pd=18240 as=0 ps=0 
M2669 diff_135960_115920# diff_82200_122760# GND GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M2670 diff_149760_115920# diff_82200_122760# GND GND efet w=1860 l=960
+ ad=0 pd=0 as=0 ps=0 
M2671 diff_163440_116040# diff_82200_122760# GND GND efet w=1920 l=840
+ ad=0 pd=0 as=0 ps=0 
M2672 Vdd Vdd Vdd GND efet w=120 l=660
+ ad=0 pd=0 as=0 ps=0 
M2673 Vdd Vdd Vdd GND efet w=420 l=780
+ ad=0 pd=0 as=0 ps=0 
M2674 Vdd Vdd diff_16320_124440# GND efet w=900 l=3660
+ ad=0 pd=0 as=0 ps=0 
M2675 diff_100560_145080# diff_88320_120720# GND GND efet w=1740 l=780
+ ad=0 pd=0 as=0 ps=0 
M2676 diff_114240_145080# diff_88320_120720# GND GND efet w=1800 l=720
+ ad=0 pd=0 as=0 ps=0 
M2677 GND diff_82200_122760# diff_175920_112080# GND efet w=1620 l=780
+ ad=0 pd=0 as=0 ps=0 
M2678 diff_233520_124920# clk2 diff_233880_120960# GND efet w=7200 l=720
+ ad=0 pd=0 as=1.40112e+07 ps=26160 
M2679 GND diff_230880_118560# diff_233880_120960# GND efet w=11280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2680 diff_189240_116040# diff_188880_122040# GND GND efet w=3240 l=720
+ ad=0 pd=0 as=0 ps=0 
M2681 diff_201120_122760# diff_188880_122040# GND GND efet w=3240 l=720
+ ad=0 pd=0 as=0 ps=0 
M2682 diff_155520_145080# diff_88320_120720# GND GND efet w=1680 l=720
+ ad=0 pd=0 as=0 ps=0 
M2683 GND diff_88320_120720# diff_86760_145200# GND efet w=1560 l=720
+ ad=0 pd=0 as=0 ps=0 
M2684 GND diff_88320_120720# diff_128040_145080# GND efet w=1560 l=720
+ ad=0 pd=0 as=0 ps=0 
M2685 GND diff_88320_120720# diff_141720_145080# GND efet w=1620 l=780
+ ad=0 pd=0 as=0 ps=0 
M2686 diff_169200_145080# diff_88320_120720# GND GND efet w=1620 l=780
+ ad=0 pd=0 as=0 ps=0 
M2687 diff_182040_114360# diff_88320_120720# GND GND efet w=1560 l=720
+ ad=0 pd=0 as=0 ps=0 
M2688 diff_8760_228840# diff_21960_110160# GND GND efet w=6600 l=720
+ ad=1.4256e+07 pd=17520 as=0 ps=0 
M2689 Vdd diff_24840_108840# diff_8760_228840# GND efet w=6960 l=720
+ ad=0 pd=0 as=0 ps=0 
M2690 diff_51600_131160# diff_51600_133800# GND GND efet w=1920 l=720
+ ad=8.2656e+06 pd=14400 as=0 ps=0 
M2691 Vdd Vdd diff_51600_131160# GND efet w=1140 l=4740
+ ad=0 pd=0 as=0 ps=0 
M2692 diff_51600_131160# diff_56640_92400# diff_57480_108840# GND efet w=840 l=720
+ ad=0 pd=0 as=6.6528e+06 ps=16320 
M2693 diff_81000_115920# diff_80880_111840# diff_81000_115920# GND efet w=3240 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2694 diff_21960_110160# diff_21960_110160# diff_21960_110160# GND efet w=240 l=720
+ ad=1.9872e+06 pd=6240 as=0 ps=0 
M2695 diff_21960_110160# diff_21960_110160# diff_21960_110160# GND efet w=120 l=720
+ ad=0 pd=0 as=0 ps=0 
M2696 diff_24840_108840# diff_24840_108840# diff_24840_108840# GND efet w=240 l=540
+ ad=2.088e+06 pd=6720 as=0 ps=0 
M2697 diff_24840_108840# diff_24840_108840# diff_24840_108840# GND efet w=240 l=660
+ ad=0 pd=0 as=0 ps=0 
M2698 diff_34920_109680# diff_20280_51120# Vdd GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2699 diff_51600_133800# diff_57480_108840# GND GND efet w=3240 l=720
+ ad=1.14336e+07 pd=23040 as=0 ps=0 
M2700 Vdd Vdd diff_51600_133800# GND efet w=1080 l=4680
+ ad=0 pd=0 as=0 ps=0 
M2701 diff_86760_145200# diff_87000_110280# diff_86760_145200# GND efet w=3120 l=4920
+ ad=0 pd=0 as=0 ps=0 
M2702 diff_21960_110160# diff_22200_108240# diff_22440_106560# GND efet w=1500 l=660
+ ad=0 pd=0 as=1.08288e+07 ps=21120 
M2703 diff_24840_108840# diff_22200_108240# diff_21960_99120# GND efet w=1440 l=840
+ ad=0 pd=0 as=8.1648e+06 ps=18240 
M2704 diff_57480_108840# diff_56160_105120# diff_34920_109680# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2705 diff_57480_108840# diff_57480_108840# diff_57480_108840# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M2706 diff_57480_108840# diff_57480_108840# diff_57480_108840# GND efet w=180 l=360
+ ad=0 pd=0 as=0 ps=0 
M2707 diff_80880_111840# diff_80880_111840# diff_80880_111840# GND efet w=300 l=300
+ ad=1.9296e+06 pd=6960 as=0 ps=0 
M2708 diff_80880_111840# diff_80880_111840# diff_80880_111840# GND efet w=180 l=360
+ ad=0 pd=0 as=0 ps=0 
M2709 diff_81000_115920# diff_80880_111840# Vdd GND efet w=840 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2710 diff_86760_145200# diff_87000_110280# Vdd GND efet w=840 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2711 diff_87000_110280# diff_87000_110280# diff_87000_110280# GND efet w=300 l=300
+ ad=1.9584e+06 pd=6960 as=0 ps=0 
M2712 diff_80880_111840# Vdd Vdd GND efet w=720 l=720
+ ad=0 pd=0 as=0 ps=0 
M2713 diff_22440_106560# diff_21960_99120# GND GND efet w=5040 l=720
+ ad=0 pd=0 as=0 ps=0 
M2714 diff_25200_276600# diff_20280_51120# Vdd GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2715 diff_57480_106560# diff_56160_105120# diff_25200_276600# GND efet w=1320 l=720
+ ad=6.2784e+06 pd=16320 as=0 ps=0 
M2716 diff_57480_106560# diff_57480_106560# diff_57480_106560# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M2717 diff_57480_106560# diff_57480_106560# diff_57480_106560# GND efet w=240 l=360
+ ad=0 pd=0 as=0 ps=0 
M2718 diff_87000_110280# diff_87000_110280# diff_87000_110280# GND efet w=180 l=360
+ ad=0 pd=0 as=0 ps=0 
M2719 diff_87000_110280# Vdd Vdd GND efet w=840 l=720
+ ad=0 pd=0 as=0 ps=0 
M2720 Vdd Vdd diff_84000_102000# GND efet w=1020 l=2880
+ ad=0 pd=0 as=2.2536e+07 ps=63360 
M2721 Vdd Vdd diff_22440_106560# GND efet w=1080 l=1920
+ ad=0 pd=0 as=0 ps=0 
M2722 diff_23040_212640# diff_20280_51120# Vdd GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M2723 diff_51600_126720# diff_57480_106560# GND GND efet w=3240 l=720
+ ad=1.14336e+07 pd=22560 as=0 ps=0 
M2724 Vdd Vdd diff_51600_126720# GND efet w=1080 l=4680
+ ad=0 pd=0 as=0 ps=0 
M2725 GND diff_82440_102720# diff_84000_102000# GND efet w=4980 l=780
+ ad=0 pd=0 as=0 ps=0 
M2726 diff_94680_112080# diff_94800_111720# diff_94680_112080# GND efet w=5100 l=2760
+ ad=0 pd=0 as=0 ps=0 
M2727 diff_100560_145080# diff_100800_110280# diff_100560_145080# GND efet w=3060 l=4740
+ ad=0 pd=0 as=0 ps=0 
M2728 diff_94800_111720# diff_94800_111720# diff_94800_111720# GND efet w=300 l=300
+ ad=2.0304e+06 pd=7680 as=0 ps=0 
M2729 diff_94800_111720# diff_94800_111720# diff_94800_111720# GND efet w=240 l=420
+ ad=0 pd=0 as=0 ps=0 
M2730 diff_94680_112080# diff_94800_111720# Vdd GND efet w=840 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2731 diff_100560_145080# diff_100800_110280# Vdd GND efet w=840 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2732 diff_100800_110280# diff_100800_110280# diff_100800_110280# GND efet w=300 l=300
+ ad=2.0592e+06 pd=7680 as=0 ps=0 
M2733 diff_100800_110280# diff_100800_110280# diff_100800_110280# GND efet w=240 l=420
+ ad=0 pd=0 as=0 ps=0 
M2734 diff_94800_111720# Vdd Vdd GND efet w=900 l=780
+ ad=0 pd=0 as=0 ps=0 
M2735 diff_100800_110280# Vdd Vdd GND efet w=840 l=840
+ ad=0 pd=0 as=0 ps=0 
M2736 diff_82200_127320# Vdd Vdd GND efet w=840 l=3120
+ ad=1.49472e+07 pd=41520 as=0 ps=0 
M2737 diff_108480_116040# diff_108360_111840# diff_108480_116040# GND efet w=3060 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2738 diff_114240_145080# diff_114480_110280# diff_114240_145080# GND efet w=3120 l=4680
+ ad=0 pd=0 as=0 ps=0 
M2739 diff_108360_111840# diff_108360_111840# diff_108360_111840# GND efet w=300 l=300
+ ad=1.9008e+06 pd=7200 as=0 ps=0 
M2740 diff_108360_111840# diff_108360_111840# diff_108360_111840# GND efet w=180 l=360
+ ad=0 pd=0 as=0 ps=0 
M2741 diff_108480_116040# diff_108360_111840# Vdd GND efet w=840 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2742 diff_114240_145080# diff_114480_110280# Vdd GND efet w=840 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2743 diff_114480_110280# diff_114480_110280# diff_114480_110280# GND efet w=300 l=300
+ ad=1.872e+06 pd=6960 as=0 ps=0 
M2744 diff_108360_111840# Vdd Vdd GND efet w=840 l=900
+ ad=0 pd=0 as=0 ps=0 
M2745 diff_114480_110280# diff_114480_110280# diff_114480_110280# GND efet w=180 l=360
+ ad=0 pd=0 as=0 ps=0 
M2746 diff_114480_110280# Vdd Vdd GND efet w=900 l=780
+ ad=0 pd=0 as=0 ps=0 
M2747 diff_122160_115920# diff_122160_112080# diff_122160_115920# GND efet w=3240 l=3360
+ ad=0 pd=0 as=0 ps=0 
M2748 diff_128040_145080# diff_128160_110400# diff_128040_145080# GND efet w=3180 l=2760
+ ad=0 pd=0 as=0 ps=0 
M2749 diff_135960_115920# diff_135840_111600# diff_135960_115920# GND efet w=3180 l=4680
+ ad=0 pd=0 as=0 ps=0 
M2750 diff_122160_112080# diff_122160_112080# diff_122160_112080# GND efet w=300 l=300
+ ad=1.9728e+06 pd=7200 as=0 ps=0 
M2751 diff_122160_112080# diff_122160_112080# diff_122160_112080# GND efet w=180 l=360
+ ad=0 pd=0 as=0 ps=0 
M2752 diff_122160_115920# diff_122160_112080# Vdd GND efet w=840 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2753 diff_128040_145080# diff_128160_110400# Vdd GND efet w=840 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2754 diff_128160_110400# diff_128160_110400# diff_128160_110400# GND efet w=300 l=300
+ ad=2.0304e+06 pd=7200 as=0 ps=0 
M2755 diff_128160_110400# diff_128160_110400# diff_128160_110400# GND efet w=180 l=420
+ ad=0 pd=0 as=0 ps=0 
M2756 diff_122160_112080# Vdd Vdd GND efet w=840 l=720
+ ad=0 pd=0 as=0 ps=0 
M2757 diff_128160_110400# Vdd Vdd GND efet w=840 l=780
+ ad=0 pd=0 as=0 ps=0 
M2758 diff_141720_145080# diff_141960_110280# diff_141720_145080# GND efet w=3180 l=4740
+ ad=0 pd=0 as=0 ps=0 
M2759 diff_135840_111600# diff_135840_111600# diff_135840_111600# GND efet w=240 l=360
+ ad=1.8576e+06 pd=6720 as=0 ps=0 
M2760 diff_135840_111600# diff_135840_111600# diff_135840_111600# GND efet w=180 l=360
+ ad=0 pd=0 as=0 ps=0 
M2761 diff_135960_115920# diff_135840_111600# Vdd GND efet w=840 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2762 diff_141720_145080# diff_141960_110280# Vdd GND efet w=840 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2763 GND diff_169680_101760# diff_189240_116040# GND efet w=1920 l=720
+ ad=0 pd=0 as=0 ps=0 
M2764 GND diff_169680_101760# diff_196560_127680# GND efet w=1920 l=780
+ ad=0 pd=0 as=0 ps=0 
M2765 GND diff_169680_101760# diff_201120_122760# GND efet w=2160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2766 GND diff_169680_101760# diff_205320_118080# GND efet w=1920 l=720
+ ad=0 pd=0 as=0 ps=0 
M2767 diff_149760_115920# diff_149640_111600# diff_149760_115920# GND efet w=3180 l=4680
+ ad=0 pd=0 as=0 ps=0 
M2768 diff_155520_145080# diff_155640_110400# diff_155520_145080# GND efet w=4920 l=2760
+ ad=0 pd=0 as=0 ps=0 
M2769 diff_141960_110280# diff_141960_110280# diff_141960_110280# GND efet w=300 l=300
+ ad=1.872e+06 pd=6720 as=0 ps=0 
M2770 diff_135840_111600# Vdd Vdd GND efet w=780 l=900
+ ad=0 pd=0 as=0 ps=0 
M2771 Vdd Vdd diff_21960_99120# GND efet w=1020 l=1980
+ ad=0 pd=0 as=0 ps=0 
M2772 diff_21960_99120# diff_21960_94200# GND GND efet w=5160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2773 diff_23160_135720# diff_20280_51120# Vdd GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M2774 Vdd Vdd diff_51600_124080# GND efet w=960 l=4680
+ ad=0 pd=0 as=1.02672e+07 ps=25440 
M2775 GND diff_84000_102000# diff_82200_127320# GND efet w=2640 l=840
+ ad=0 pd=0 as=0 ps=0 
M2776 diff_82440_133920# diff_112680_97560# GND GND efet w=3840 l=840
+ ad=1.57536e+07 pd=40320 as=0 ps=0 
M2777 Vdd Vdd diff_82440_133920# GND efet w=840 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2778 diff_130200_104880# Vdd Vdd GND efet w=840 l=3120
+ ad=1.49328e+07 pd=42960 as=0 ps=0 
M2779 diff_141960_110280# diff_141960_110280# diff_141960_110280# GND efet w=180 l=360
+ ad=0 pd=0 as=0 ps=0 
M2780 diff_141960_110280# Vdd Vdd GND efet w=840 l=840
+ ad=0 pd=0 as=0 ps=0 
M2781 diff_149640_111600# diff_149640_111600# diff_149640_111600# GND efet w=300 l=300
+ ad=2.0736e+06 pd=7440 as=0 ps=0 
M2782 diff_149640_111600# diff_149640_111600# diff_149640_111600# GND efet w=240 l=420
+ ad=0 pd=0 as=0 ps=0 
M2783 diff_149760_115920# diff_149640_111600# Vdd GND efet w=840 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2784 diff_155520_145080# diff_155640_110400# Vdd GND efet w=840 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2785 diff_155640_110400# diff_155640_110400# diff_155640_110400# GND efet w=180 l=420
+ ad=2.0592e+06 pd=7440 as=0 ps=0 
M2786 diff_149640_111600# Vdd Vdd GND efet w=960 l=780
+ ad=0 pd=0 as=0 ps=0 
M2787 diff_155640_110400# diff_155640_110400# diff_155640_110400# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M2788 diff_155640_110400# Vdd Vdd GND efet w=960 l=720
+ ad=0 pd=0 as=0 ps=0 
M2789 diff_130200_104880# diff_82440_133920# GND GND efet w=2520 l=720
+ ad=0 pd=0 as=0 ps=0 
M2790 diff_109680_129600# diff_140160_97560# GND GND efet w=3840 l=840
+ ad=1.59408e+07 pd=42480 as=0 ps=0 
M2791 Vdd Vdd diff_109680_129600# GND efet w=840 l=3120
+ ad=0 pd=0 as=0 ps=0 
M2792 diff_82200_132000# Vdd Vdd GND efet w=780 l=3060
+ ad=1.3896e+07 pd=40080 as=0 ps=0 
M2793 diff_163440_116040# diff_163320_111840# diff_163440_116040# GND efet w=3060 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2794 diff_169200_145080# diff_169440_110280# diff_169200_145080# GND efet w=4860 l=2460
+ ad=0 pd=0 as=0 ps=0 
M2795 diff_163320_111840# diff_163320_111840# diff_163320_111840# GND efet w=240 l=360
+ ad=1.8864e+06 pd=6720 as=0 ps=0 
M2796 diff_163320_111840# diff_163320_111840# diff_163320_111840# GND efet w=180 l=360
+ ad=0 pd=0 as=0 ps=0 
M2797 diff_163440_116040# diff_163320_111840# Vdd GND efet w=840 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2798 diff_169200_145080# diff_169440_110280# Vdd GND efet w=840 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2799 diff_169440_110280# diff_169440_110280# diff_169440_110280# GND efet w=240 l=300
+ ad=2.016e+06 pd=7440 as=0 ps=0 
M2800 diff_163320_111840# Vdd Vdd GND efet w=840 l=780
+ ad=0 pd=0 as=0 ps=0 
M2801 diff_169440_110280# diff_169440_110280# diff_169440_110280# GND efet w=300 l=360
+ ad=0 pd=0 as=0 ps=0 
M2802 diff_175920_112080# diff_176640_109320# diff_175920_112080# GND efet w=4800 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2803 diff_182040_114360# diff_181920_110280# diff_182040_114360# GND efet w=4860 l=2460
+ ad=0 pd=0 as=0 ps=0 
M2804 diff_176640_109320# diff_176640_109320# diff_176640_109320# GND efet w=240 l=360
+ ad=2.2176e+06 pd=7440 as=0 ps=0 
M2805 diff_176640_109320# diff_176640_109320# diff_176640_109320# GND efet w=240 l=360
+ ad=0 pd=0 as=0 ps=0 
M2806 diff_175920_112080# diff_176640_109320# Vdd GND efet w=840 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2807 diff_182040_114360# diff_181920_110280# Vdd GND efet w=840 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2808 diff_181920_110280# diff_181920_110280# diff_181920_110280# GND efet w=240 l=300
+ ad=2.0304e+06 pd=7440 as=0 ps=0 
M2809 diff_169440_110280# Vdd Vdd GND efet w=900 l=780
+ ad=0 pd=0 as=0 ps=0 
M2810 Vdd Vdd Vdd GND efet w=360 l=960
+ ad=0 pd=0 as=0 ps=0 
M2811 Vdd Vdd Vdd GND efet w=360 l=960
+ ad=0 pd=0 as=0 ps=0 
M2812 Vdd Vdd Vdd GND efet w=660 l=420
+ ad=0 pd=0 as=0 ps=0 
M2813 Vdd Vdd Vdd GND efet w=360 l=840
+ ad=0 pd=0 as=0 ps=0 
M2814 Vdd Vdd diff_82200_122760# GND efet w=960 l=3120
+ ad=0 pd=0 as=5.112e+06 ps=14880 
M2815 diff_82200_132000# diff_109680_129600# GND GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M2816 diff_176640_109320# Vdd Vdd GND efet w=840 l=840
+ ad=0 pd=0 as=0 ps=0 
M2817 diff_181920_110280# diff_181920_110280# diff_181920_110280# GND efet w=300 l=360
+ ad=0 pd=0 as=0 ps=0 
M2818 diff_181920_110280# Vdd Vdd GND efet w=900 l=720
+ ad=0 pd=0 as=0 ps=0 
M2819 Vdd Vdd Vdd GND efet w=180 l=660
+ ad=0 pd=0 as=0 ps=0 
M2820 Vdd Vdd Vdd GND efet w=300 l=900
+ ad=0 pd=0 as=0 ps=0 
M2821 Vdd Vdd Vdd GND efet w=180 l=540
+ ad=0 pd=0 as=0 ps=0 
M2822 Vdd Vdd Vdd GND efet w=660 l=420
+ ad=0 pd=0 as=0 ps=0 
M2823 diff_82200_122760# diff_82200_122760# diff_82200_122760# GND efet w=240 l=300
+ ad=0 pd=0 as=0 ps=0 
M2824 diff_82200_122760# diff_82200_122760# diff_82200_122760# GND efet w=300 l=420
+ ad=0 pd=0 as=0 ps=0 
M2825 Vdd Vdd diff_88320_120720# GND efet w=840 l=3000
+ ad=0 pd=0 as=4.7808e+06 ps=14160 
M2826 diff_189240_116040# diff_189000_112080# diff_189240_116040# GND efet w=3120 l=4920
+ ad=0 pd=0 as=0 ps=0 
M2827 diff_189000_112080# diff_189000_112080# diff_189000_112080# GND efet w=300 l=300
+ ad=1.9872e+06 pd=7440 as=0 ps=0 
M2828 diff_189000_112080# diff_189000_112080# diff_189000_112080# GND efet w=300 l=360
+ ad=0 pd=0 as=0 ps=0 
M2829 diff_189240_116040# diff_189000_112080# Vdd GND efet w=840 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2830 diff_189000_112080# Vdd Vdd GND efet w=840 l=840
+ ad=0 pd=0 as=0 ps=0 
M2831 diff_230880_118560# Vdd Vdd GND efet w=1080 l=2760
+ ad=5.1552e+06 pd=11280 as=0 ps=0 
M2832 GND diff_232800_116760# diff_230880_118560# GND efet w=3900 l=660
+ ad=0 pd=0 as=0 ps=0 
M2833 diff_196560_127680# diff_197040_110280# diff_196560_127680# GND efet w=5340 l=2580
+ ad=0 pd=0 as=0 ps=0 
M2834 diff_196560_127680# diff_197040_110280# Vdd GND efet w=840 l=3840
+ ad=0 pd=0 as=0 ps=0 
M2835 diff_201120_122760# diff_202080_109320# diff_201120_122760# GND efet w=5040 l=2820
+ ad=0 pd=0 as=0 ps=0 
M2836 diff_232800_116760# diff_232800_116760# diff_232800_116760# GND efet w=120 l=480
+ ad=5.7024e+06 pd=11040 as=0 ps=0 
M2837 diff_197040_110280# diff_197040_110280# diff_197040_110280# GND efet w=240 l=360
+ ad=1.8288e+06 pd=6960 as=0 ps=0 
M2838 diff_197040_110280# diff_197040_110280# diff_197040_110280# GND efet w=240 l=360
+ ad=0 pd=0 as=0 ps=0 
M2839 diff_169680_101760# Vdd Vdd GND efet w=900 l=3180
+ ad=8.568e+06 pd=20880 as=0 ps=0 
M2840 diff_88320_120720# diff_88320_120720# diff_88320_120720# GND efet w=180 l=360
+ ad=0 pd=0 as=0 ps=0 
M2841 diff_88320_120720# diff_88320_120720# diff_88320_120720# GND efet w=240 l=360
+ ad=0 pd=0 as=0 ps=0 
M2842 diff_202080_109320# diff_202080_109320# diff_202080_109320# GND efet w=240 l=360
+ ad=1.872e+06 pd=6720 as=0 ps=0 
M2843 diff_202080_109320# diff_202080_109320# diff_202080_109320# GND efet w=180 l=540
+ ad=0 pd=0 as=0 ps=0 
M2844 diff_201120_122760# diff_202080_109320# Vdd GND efet w=840 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2845 diff_197040_110280# Vdd Vdd GND efet w=720 l=780
+ ad=0 pd=0 as=0 ps=0 
M2846 diff_202080_109320# Vdd Vdd GND efet w=720 l=720
+ ad=0 pd=0 as=0 ps=0 
M2847 Vdd Vdd Vdd GND efet w=660 l=420
+ ad=0 pd=0 as=0 ps=0 
M2848 Vdd Vdd Vdd GND efet w=300 l=840
+ ad=0 pd=0 as=0 ps=0 
M2849 Vdd Vdd Vdd GND efet w=660 l=420
+ ad=0 pd=0 as=0 ps=0 
M2850 diff_197400_124560# diff_197400_124560# diff_197400_124560# GND efet w=360 l=600
+ ad=1.00368e+07 pd=19680 as=0 ps=0 
M2851 Vdd Vdd Vdd GND efet w=360 l=840
+ ad=0 pd=0 as=0 ps=0 
M2852 Vdd Vdd diff_197400_124560# GND efet w=840 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2853 diff_197400_124560# diff_188880_122040# GND GND efet w=4200 l=720
+ ad=0 pd=0 as=0 ps=0 
M2854 diff_197400_124560# diff_197400_124560# diff_197400_124560# GND efet w=240 l=240
+ ad=0 pd=0 as=0 ps=0 
M2855 diff_169680_101760# diff_169680_101760# diff_169680_101760# GND efet w=180 l=720
+ ad=0 pd=0 as=0 ps=0 
M2856 diff_169680_101760# diff_169680_101760# diff_169680_101760# GND efet w=300 l=480
+ ad=0 pd=0 as=0 ps=0 
M2857 diff_190200_129480# Vdd Vdd GND efet w=900 l=3660
+ ad=6.4944e+06 pd=14160 as=0 ps=0 
M2858 diff_190200_129480# diff_190200_129480# diff_190200_129480# GND efet w=360 l=840
+ ad=0 pd=0 as=0 ps=0 
M2859 diff_190200_129480# diff_190200_129480# diff_190200_129480# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M2860 diff_169680_101760# diff_187920_102120# GND GND efet w=4680 l=780
+ ad=0 pd=0 as=0 ps=0 
M2861 diff_57480_106560# diff_56640_92400# diff_51600_124080# GND efet w=840 l=720
+ ad=0 pd=0 as=0 ps=0 
M2862 diff_51600_124080# diff_51600_126720# GND GND efet w=1920 l=720
+ ad=0 pd=0 as=0 ps=0 
M2863 diff_82200_122760# diff_169680_101760# diff_170040_100680# GND efet w=4920 l=720
+ ad=0 pd=0 as=4.7232e+06 ps=11760 
M2864 diff_88320_120720# diff_169680_101760# diff_177840_100680# GND efet w=4920 l=720
+ ad=0 pd=0 as=6.2928e+06 ps=16080 
M2865 GND diff_196080_127080# diff_190200_129480# GND efet w=3720 l=720
+ ad=0 pd=0 as=0 ps=0 
M2866 diff_232800_116760# diff_232800_116760# diff_232800_116760# GND efet w=360 l=360
+ ad=0 pd=0 as=0 ps=0 
M2867 diff_232800_116760# Vdd Vdd GND efet w=900 l=5820
+ ad=0 pd=0 as=0 ps=0 
M2868 diff_239520_113040# diff_179280_17640# diff_232800_116760# GND efet w=2640 l=720
+ ad=8.928e+06 pd=18480 as=0 ps=0 
M2869 diff_239520_113040# diff_88080_99240# GND GND efet w=2760 l=720
+ ad=0 pd=0 as=0 ps=0 
M2870 GND diff_84840_96840# diff_239520_113040# GND efet w=3000 l=660
+ ad=0 pd=0 as=0 ps=0 
M2871 diff_26880_44640# clk1 diff_243600_101280# GND efet w=1500 l=660
+ ad=1.08576e+07 pd=23760 as=2.5488e+06 ps=6480 
M2872 diff_177360_99960# diff_177360_99960# diff_177360_99960# GND efet w=180 l=360
+ ad=8.5968e+06 pd=20160 as=0 ps=0 
M2873 diff_187920_102120# diff_187920_102120# diff_187920_102120# GND efet w=180 l=420
+ ad=8.928e+06 pd=20160 as=0 ps=0 
M2874 diff_188880_122040# diff_188880_122040# diff_188880_122040# GND efet w=180 l=420
+ ad=8.4672e+06 pd=19440 as=0 ps=0 
M2875 diff_177360_99960# diff_177360_99960# diff_177360_99960# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M2876 diff_187920_102120# diff_187920_102120# diff_187920_102120# GND efet w=240 l=240
+ ad=0 pd=0 as=0 ps=0 
M2877 diff_188880_122040# diff_188880_122040# diff_188880_122040# GND efet w=240 l=240
+ ad=0 pd=0 as=0 ps=0 
M2878 diff_88080_94680# diff_88080_99240# diff_82440_102720# GND efet w=1320 l=720
+ ad=1.56528e+07 pd=30960 as=8.2512e+06 ps=16800 
M2879 diff_112680_97560# diff_88080_99240# diff_115560_93600# GND efet w=1440 l=720
+ ad=1.0224e+07 pd=20880 as=1.4616e+07 ps=31200 
M2880 diff_170040_100680# diff_88320_120720# GND GND efet w=5100 l=780
+ ad=0 pd=0 as=0 ps=0 
M2881 diff_140160_97560# diff_88080_99240# diff_143040_93480# GND efet w=1320 l=720
+ ad=9.7056e+06 pd=20640 as=1.44288e+07 ps=30720 
M2882 diff_177840_100680# diff_177360_99960# GND GND efet w=7560 l=720
+ ad=0 pd=0 as=0 ps=0 
M2883 diff_82440_102720# diff_84840_96840# diff_76800_82320# GND efet w=1320 l=720
+ ad=0 pd=0 as=1.30032e+07 ps=33360 
M2884 diff_56160_105120# diff_56640_92400# GND GND efet w=1440 l=720
+ ad=4.32e+06 pd=10800 as=0 ps=0 
M2885 Vdd Vdd diff_56160_105120# GND efet w=840 l=5880
+ ad=0 pd=0 as=0 ps=0 
M2886 diff_112680_97560# diff_84840_96840# diff_104280_82320# GND efet w=1320 l=720
+ ad=0 pd=0 as=1.31328e+07 ps=34560 
M2887 diff_177360_99960# diff_88080_99240# diff_178440_81000# GND efet w=1440 l=720
+ ad=0 pd=0 as=1.5552e+07 ps=31920 
M2888 GND diff_243600_101280# diff_84840_96840# GND efet w=5280 l=600
+ ad=0 pd=0 as=1.7496e+07 ps=36240 
M2889 diff_196080_127080# diff_196080_127080# diff_196080_127080# GND efet w=360 l=840
+ ad=1.044e+07 pd=22080 as=0 ps=0 
M2890 diff_187920_102120# diff_88080_99240# diff_169200_62280# GND efet w=1320 l=720
+ ad=0 pd=0 as=1.26e+07 ps=29280 
M2891 diff_140160_97560# diff_84840_96840# diff_132360_82560# GND efet w=1380 l=720
+ ad=0 pd=0 as=8.856e+06 ps=25680 
M2892 diff_104280_82320# diff_104280_82320# diff_104280_82320# GND efet w=300 l=420
+ ad=0 pd=0 as=0 ps=0 
M2893 diff_104280_82320# diff_104280_82320# diff_104280_82320# GND efet w=120 l=480
+ ad=0 pd=0 as=0 ps=0 
M2894 Vdd Vdd diff_23760_86280# GND efet w=840 l=960
+ ad=0 pd=0 as=1.7568e+06 ps=6480 
M2895 diff_23760_86280# diff_23760_86280# diff_23760_86280# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M2896 diff_23760_86280# diff_23760_86280# diff_23760_86280# GND efet w=180 l=540
+ ad=0 pd=0 as=0 ps=0 
M2897 Vdd diff_23760_86280# diff_22200_108240# GND efet w=960 l=960
+ ad=0 pd=0 as=1.44432e+07 ps=25200 
M2898 diff_22200_108240# diff_23760_86280# diff_22200_108240# GND efet w=3660 l=2700
+ ad=0 pd=0 as=0 ps=0 
M2899 diff_115560_93600# diff_115560_93600# diff_115560_93600# GND efet w=240 l=480
+ ad=0 pd=0 as=0 ps=0 
M2900 diff_115560_93600# diff_115560_93600# diff_115560_93600# GND efet w=120 l=480
+ ad=0 pd=0 as=0 ps=0 
M2901 diff_177360_99960# diff_84840_96840# diff_159840_82560# GND efet w=1320 l=720
+ ad=0 pd=0 as=9.2016e+06 ps=26160 
M2902 diff_132360_82560# diff_132360_82560# diff_132360_82560# GND efet w=300 l=660
+ ad=0 pd=0 as=0 ps=0 
M2903 diff_132360_82560# diff_132360_82560# diff_132360_82560# GND efet w=120 l=360
+ ad=0 pd=0 as=0 ps=0 
M2904 diff_22200_108240# clk2 GND GND efet w=5100 l=660
+ ad=0 pd=0 as=0 ps=0 
M2905 Vdd Vdd diff_76800_82320# GND efet w=1080 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2906 diff_76440_81600# Vdd Vdd GND efet w=720 l=4560
+ ad=7.3152e+06 pd=18960 as=0 ps=0 
M2907 diff_76800_82320# diff_76440_81600# GND GND efet w=3360 l=840
+ ad=0 pd=0 as=0 ps=0 
M2908 diff_76440_81600# diff_76440_81600# diff_76440_81600# GND efet w=240 l=720
+ ad=0 pd=0 as=0 ps=0 
M2909 diff_76440_81600# diff_76440_81600# diff_76440_81600# GND efet w=180 l=420
+ ad=0 pd=0 as=0 ps=0 
M2910 Vdd Vdd diff_83880_78000# GND efet w=840 l=5760
+ ad=0 pd=0 as=6.2928e+06 ps=15120 
M2911 diff_77520_78480# Vdd Vdd GND efet w=720 l=4560
+ ad=7.5888e+06 pd=18000 as=0 ps=0 
M2912 diff_77520_78480# diff_77520_78480# diff_77520_78480# GND efet w=240 l=720
+ ad=0 pd=0 as=0 ps=0 
M2913 diff_77520_78480# diff_77520_78480# diff_77520_78480# GND efet w=240 l=480
+ ad=0 pd=0 as=0 ps=0 
M2914 GND diff_77520_78480# diff_83880_78000# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M2915 GND diff_38640_64440# diff_54360_73680# GND efet w=1440 l=720
+ ad=0 pd=0 as=8.136e+06 ps=21120 
M2916 GND diff_77520_78480# diff_76440_81600# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M2917 diff_54360_73680# diff_54360_73680# diff_54360_73680# GND efet w=660 l=420
+ ad=0 pd=0 as=0 ps=0 
M2918 diff_54360_73680# diff_54360_73680# diff_54360_73680# GND efet w=360 l=840
+ ad=0 pd=0 as=0 ps=0 
M2919 diff_76800_82320# diff_76800_82320# diff_76800_82320# GND efet w=300 l=420
+ ad=0 pd=0 as=0 ps=0 
M2920 diff_76800_82320# diff_76800_82320# diff_76800_82320# GND efet w=240 l=660
+ ad=0 pd=0 as=0 ps=0 
M2921 diff_83880_78000# diff_38640_64440# diff_76440_70800# GND efet w=1500 l=780
+ ad=0 pd=0 as=4.464e+06 ps=9120 
M2922 Vdd Vdd diff_88080_94680# GND efet w=1080 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2923 Vdd Vdd diff_99120_74280# GND efet w=840 l=5760
+ ad=0 pd=0 as=4.9248e+06 ps=14640 
M2924 Vdd Vdd diff_104280_82320# GND efet w=1140 l=2460
+ ad=0 pd=0 as=0 ps=0 
M2925 diff_88080_94680# diff_88080_94680# diff_88080_94680# GND efet w=180 l=540
+ ad=0 pd=0 as=0 ps=0 
M2926 GND diff_76440_81600# diff_77520_78480# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2927 diff_88080_94680# diff_88080_94680# diff_88080_94680# GND efet w=360 l=360
+ ad=0 pd=0 as=0 ps=0 
M2928 diff_99120_74280# diff_99120_74280# diff_99120_74280# GND efet w=180 l=660
+ ad=0 pd=0 as=0 ps=0 
M2929 diff_99120_74280# diff_99120_74280# diff_99120_74280# GND efet w=300 l=480
+ ad=0 pd=0 as=0 ps=0 
M2930 diff_76800_82320# diff_38640_64440# diff_86280_74040# GND efet w=1440 l=720
+ ad=0 pd=0 as=4.4784e+06 ps=9120 
M2931 diff_76440_81600# diff_54360_73680# diff_75480_71160# GND efet w=3060 l=780
+ ad=0 pd=0 as=6.8832e+06 ps=16800 
M2932 diff_37800_73440# clk2 sync GND efet w=840 l=720
+ ad=2.7936e+06 pd=7920 as=4.36176e+07 ps=100560 
M2933 diff_37800_73440# diff_37800_73440# diff_37800_73440# GND efet w=240 l=240
+ ad=0 pd=0 as=0 ps=0 
M2934 diff_37800_73440# diff_37800_73440# diff_37800_73440# GND efet w=180 l=480
+ ad=0 pd=0 as=0 ps=0 
M2935 diff_39600_69360# diff_37800_73440# GND GND efet w=3120 l=720
+ ad=6.2496e+06 pd=13200 as=0 ps=0 
M2936 Vdd Vdd diff_39600_69360# GND efet w=840 l=5760
+ ad=0 pd=0 as=0 ps=0 
M2937 diff_54360_73680# Vdd Vdd GND efet w=960 l=5880
+ ad=0 pd=0 as=0 ps=0 
M2938 GND diff_54480_70200# diff_54360_73680# GND efet w=1380 l=780
+ ad=0 pd=0 as=0 ps=0 
M2939 GND diff_76440_70800# diff_75480_71160# GND efet w=5100 l=780
+ ad=0 pd=0 as=0 ps=0 
M2940 diff_54480_70200# diff_54480_70200# diff_54480_70200# GND efet w=300 l=300
+ ad=4.8816e+06 pd=12960 as=0 ps=0 
M2941 diff_54480_70200# diff_54480_70200# diff_54480_70200# GND efet w=300 l=660
+ ad=0 pd=0 as=0 ps=0 
M2942 diff_37920_64080# clk1 diff_39600_69360# GND efet w=900 l=780
+ ad=3.4848e+06 pd=9120 as=0 ps=0 
M2943 diff_54480_70200# Vdd Vdd GND efet w=660 l=5460
+ ad=0 pd=0 as=0 ps=0 
M2944 diff_38640_64440# diff_37920_64080# GND GND efet w=2040 l=720
+ ad=4.3488e+06 pd=10800 as=0 ps=0 
M2945 diff_54480_70200# diff_39600_69360# GND GND efet w=1200 l=840
+ ad=0 pd=0 as=0 ps=0 
M2946 Vdd Vdd diff_38640_64440# GND efet w=840 l=4140
+ ad=0 pd=0 as=0 ps=0 
M2947 diff_38640_64440# clk2 diff_35400_61080# GND efet w=900 l=660
+ ad=0 pd=0 as=2.3184e+06 ps=6720 
M2948 GND diff_35400_61080# diff_35640_60240# GND efet w=1500 l=660
+ ad=0 pd=0 as=6.2064e+06 ps=15120 
M2949 diff_88080_94680# diff_95040_69120# diff_96600_67920# GND efet w=1320 l=840
+ ad=0 pd=0 as=1.07136e+07 ps=24720 
M2950 diff_77520_78480# diff_54360_73680# diff_90480_74640# GND efet w=2760 l=720
+ ad=0 pd=0 as=7.8912e+06 ps=18000 
M2951 diff_90480_74640# diff_86280_74040# GND GND efet w=5160 l=720
+ ad=0 pd=0 as=0 ps=0 
M2952 GND diff_99120_74280# diff_88080_94680# GND efet w=2520 l=720
+ ad=0 pd=0 as=0 ps=0 
M2953 diff_103920_81600# Vdd Vdd GND efet w=720 l=4560
+ ad=7.5744e+06 pd=19440 as=0 ps=0 
M2954 diff_104280_82320# diff_103920_81600# GND GND efet w=3360 l=840
+ ad=0 pd=0 as=0 ps=0 
M2955 diff_103920_81600# diff_103920_81600# diff_103920_81600# GND efet w=240 l=720
+ ad=0 pd=0 as=0 ps=0 
M2956 diff_103920_81600# diff_103920_81600# diff_103920_81600# GND efet w=240 l=420
+ ad=0 pd=0 as=0 ps=0 
M2957 Vdd Vdd diff_111360_78000# GND efet w=840 l=5760
+ ad=0 pd=0 as=6.048e+06 ps=15120 
M2958 diff_105000_78480# Vdd Vdd GND efet w=780 l=4500
+ ad=7.416e+06 pd=17760 as=0 ps=0 
M2959 diff_105000_78480# diff_105000_78480# diff_105000_78480# GND efet w=180 l=660
+ ad=0 pd=0 as=0 ps=0 
M2960 diff_105000_78480# diff_105000_78480# diff_105000_78480# GND efet w=240 l=480
+ ad=0 pd=0 as=0 ps=0 
M2961 GND diff_105000_78480# diff_111360_78000# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M2962 GND diff_105000_78480# diff_103920_81600# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2963 diff_104280_82320# diff_104280_82320# diff_104280_82320# GND efet w=240 l=420
+ ad=0 pd=0 as=0 ps=0 
M2964 diff_104280_82320# diff_104280_82320# diff_104280_82320# GND efet w=240 l=540
+ ad=0 pd=0 as=0 ps=0 
M2965 diff_111360_78000# diff_76440_81600# diff_103920_70800# GND efet w=1500 l=900
+ ad=0 pd=0 as=4.4064e+06 ps=9120 
M2966 diff_143040_93480# diff_143040_93480# diff_143040_93480# GND efet w=240 l=360
+ ad=0 pd=0 as=0 ps=0 
M2967 diff_159840_82560# diff_159840_82560# diff_159840_82560# GND efet w=420 l=420
+ ad=0 pd=0 as=0 ps=0 
M2968 diff_178440_81000# diff_178440_81000# diff_178440_81000# GND efet w=240 l=480
+ ad=0 pd=0 as=0 ps=0 
M2969 diff_143040_93480# diff_143040_93480# diff_143040_93480# GND efet w=120 l=480
+ ad=0 pd=0 as=0 ps=0 
M2970 diff_159840_82560# diff_159840_82560# diff_159840_82560# GND efet w=180 l=180
+ ad=0 pd=0 as=0 ps=0 
M2971 diff_188880_122040# diff_88080_99240# diff_148920_43440# GND efet w=1440 l=720
+ ad=0 pd=0 as=1.2024e+07 ps=28320 
M2972 Vdd Vdd Vdd GND efet w=180 l=360
+ ad=0 pd=0 as=0 ps=0 
M2973 diff_196080_127080# diff_196080_127080# diff_196080_127080# GND efet w=540 l=420
+ ad=0 pd=0 as=0 ps=0 
M2974 diff_187920_102120# diff_84840_96840# diff_187320_82560# GND efet w=1440 l=720
+ ad=0 pd=0 as=9.9216e+06 ps=27360 
M2975 diff_188880_122040# diff_84840_96840# diff_104280_82320# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M2976 diff_178440_81000# diff_178440_81000# diff_178440_81000# GND efet w=120 l=480
+ ad=0 pd=0 as=0 ps=0 
M2977 diff_187320_82560# diff_187320_82560# diff_187320_82560# GND efet w=420 l=420
+ ad=0 pd=0 as=0 ps=0 
M2978 diff_169200_62280# diff_169200_62280# diff_169200_62280# GND efet w=300 l=480
+ ad=0 pd=0 as=0 ps=0 
M2979 diff_187320_82560# diff_187320_82560# diff_187320_82560# GND efet w=120 l=480
+ ad=0 pd=0 as=0 ps=0 
M2980 diff_169200_62280# diff_169200_62280# diff_169200_62280# GND efet w=120 l=480
+ ad=0 pd=0 as=0 ps=0 
M2981 Vdd Vdd Vdd GND efet w=360 l=540
+ ad=0 pd=0 as=0 ps=0 
M2982 diff_84840_96840# Vdd Vdd GND efet w=1080 l=1920
+ ad=0 pd=0 as=0 ps=0 
M2983 diff_196080_127080# diff_88080_99240# diff_158520_43200# GND efet w=1320 l=720
+ ad=0 pd=0 as=1.2168e+07 ps=29040 
M2984 diff_148920_43440# diff_148920_43440# diff_148920_43440# GND efet w=240 l=420
+ ad=0 pd=0 as=0 ps=0 
M2985 diff_196080_127080# diff_84840_96840# diff_76800_82320# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M2986 diff_115560_93600# Vdd Vdd GND efet w=1020 l=3780
+ ad=0 pd=0 as=0 ps=0 
M2987 Vdd Vdd diff_126600_74280# GND efet w=840 l=5760
+ ad=0 pd=0 as=4.9248e+06 ps=14640 
M2988 Vdd Vdd diff_132360_82560# GND efet w=1080 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2989 diff_131520_76200# Vdd Vdd GND efet w=720 l=5040
+ ad=7.4592e+06 pd=19920 as=0 ps=0 
M2990 diff_115560_93600# diff_115560_93600# diff_115560_93600# GND efet w=180 l=540
+ ad=0 pd=0 as=0 ps=0 
M2991 GND diff_103920_81600# diff_105000_78480# GND efet w=1500 l=780
+ ad=0 pd=0 as=0 ps=0 
M2992 diff_115560_93600# diff_115560_93600# diff_115560_93600# GND efet w=360 l=360
+ ad=0 pd=0 as=0 ps=0 
M2993 diff_126600_74280# diff_126600_74280# diff_126600_74280# GND efet w=180 l=660
+ ad=0 pd=0 as=0 ps=0 
M2994 diff_126600_74280# diff_126600_74280# diff_126600_74280# GND efet w=300 l=360
+ ad=0 pd=0 as=0 ps=0 
M2995 diff_104280_82320# diff_76440_81600# diff_113760_74280# GND efet w=1560 l=720
+ ad=0 pd=0 as=4.4496e+06 ps=9120 
M2996 diff_103920_81600# diff_77520_78480# diff_102720_72840# GND efet w=2940 l=720
+ ad=0 pd=0 as=8.0928e+06 ps=18480 
M2997 diff_96600_67920# diff_96600_67920# diff_96600_67920# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M2998 diff_96600_67920# diff_96600_67920# diff_96600_67920# GND efet w=180 l=180
+ ad=0 pd=0 as=0 ps=0 
M2999 diff_99120_74280# diff_96600_67920# GND GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M3000 GND diff_103920_70800# diff_102720_72840# GND efet w=5820 l=780
+ ad=0 pd=0 as=0 ps=0 
M3001 diff_115560_93600# diff_95040_69120# diff_124080_67440# GND efet w=1320 l=780
+ ad=0 pd=0 as=1.11024e+07 ps=25680 
M3002 diff_105000_78480# diff_77520_78480# diff_117960_74760# GND efet w=2760 l=720
+ ad=0 pd=0 as=7.92e+06 ps=17760 
M3003 GND diff_113760_74280# diff_117960_74760# GND efet w=5100 l=780
+ ad=0 pd=0 as=0 ps=0 
M3004 GND diff_126600_74280# diff_115560_93600# GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M3005 diff_132360_82560# diff_131520_76200# GND GND efet w=2520 l=780
+ ad=0 pd=0 as=0 ps=0 
M3006 diff_131520_76200# diff_131520_76200# diff_131520_76200# GND efet w=120 l=600
+ ad=0 pd=0 as=0 ps=0 
M3007 diff_131520_76200# diff_131520_76200# diff_131520_76200# GND efet w=300 l=480
+ ad=0 pd=0 as=0 ps=0 
M3008 Vdd Vdd diff_138960_78000# GND efet w=840 l=5760
+ ad=0 pd=0 as=5.5728e+06 ps=14160 
M3009 diff_132480_78480# Vdd Vdd GND efet w=720 l=4560
+ ad=7.4016e+06 pd=18000 as=0 ps=0 
M3010 diff_132480_78480# diff_132480_78480# diff_132480_78480# GND efet w=120 l=600
+ ad=0 pd=0 as=0 ps=0 
M3011 diff_132480_78480# diff_132480_78480# diff_132480_78480# GND efet w=240 l=480
+ ad=0 pd=0 as=0 ps=0 
M3012 GND diff_132480_78480# diff_138960_78000# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M3013 GND diff_132480_78480# diff_131520_76200# GND efet w=1440 l=840
+ ad=0 pd=0 as=0 ps=0 
M3014 diff_132360_82560# diff_132360_82560# diff_132360_82560# GND efet w=240 l=420
+ ad=0 pd=0 as=0 ps=0 
M3015 diff_132360_82560# diff_132360_82560# diff_132360_82560# GND efet w=240 l=300
+ ad=0 pd=0 as=0 ps=0 
M3016 diff_148920_43440# diff_148920_43440# diff_148920_43440# GND efet w=120 l=600
+ ad=0 pd=0 as=0 ps=0 
M3017 diff_84840_96840# diff_84840_96840# diff_84840_96840# GND efet w=180 l=540
+ ad=0 pd=0 as=0 ps=0 
M3018 diff_84840_96840# diff_84840_96840# diff_84840_96840# GND efet w=360 l=360
+ ad=0 pd=0 as=0 ps=0 
M3019 diff_158520_43200# diff_158520_43200# diff_158520_43200# GND efet w=240 l=480
+ ad=0 pd=0 as=0 ps=0 
M3020 diff_84840_96840# clk2 diff_243600_92760# GND efet w=1440 l=720
+ ad=0 pd=0 as=2.5632e+06 ps=6480 
M3021 diff_158520_43200# diff_158520_43200# diff_158520_43200# GND efet w=120 l=480
+ ad=0 pd=0 as=0 ps=0 
M3022 Vdd Vdd diff_143040_93480# GND efet w=960 l=3720
+ ad=0 pd=0 as=0 ps=0 
M3023 Vdd Vdd diff_154080_74280# GND efet w=840 l=5760
+ ad=0 pd=0 as=5.904e+06 ps=15120 
M3024 Vdd Vdd diff_159840_82560# GND efet w=960 l=3720
+ ad=0 pd=0 as=0 ps=0 
M3025 diff_159000_76200# Vdd Vdd GND efet w=720 l=4560
+ ad=7.3728e+06 pd=19680 as=0 ps=0 
M3026 GND diff_243600_92760# diff_218760_63360# GND efet w=2580 l=720
+ ad=0 pd=0 as=2.96928e+07 ps=82080 
M3027 diff_143040_93480# diff_143040_93480# diff_143040_93480# GND efet w=180 l=540
+ ad=0 pd=0 as=0 ps=0 
M3028 GND diff_131520_76200# diff_132480_78480# GND efet w=1500 l=720
+ ad=0 pd=0 as=0 ps=0 
M3029 diff_143040_93480# diff_143040_93480# diff_143040_93480# GND efet w=360 l=360
+ ad=0 pd=0 as=0 ps=0 
M3030 diff_154080_74280# diff_154080_74280# diff_154080_74280# GND efet w=180 l=660
+ ad=0 pd=0 as=0 ps=0 
M3031 diff_154080_74280# diff_154080_74280# diff_154080_74280# GND efet w=300 l=360
+ ad=0 pd=0 as=0 ps=0 
M3032 diff_138960_78000# diff_103920_81600# diff_131400_70800# GND efet w=1320 l=840
+ ad=0 pd=0 as=4.3056e+06 ps=9600 
M3033 diff_132360_82560# diff_103920_81600# diff_141240_74160# GND efet w=1440 l=840
+ ad=0 pd=0 as=4.464e+06 ps=9120 
M3034 diff_124080_67440# diff_124080_67440# diff_124080_67440# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M3035 diff_131520_76200# diff_105000_78480# diff_130320_71160# GND efet w=3180 l=780
+ ad=0 pd=0 as=7.8768e+06 ps=18480 
M3036 diff_124080_67440# diff_124080_67440# diff_124080_67440# GND efet w=180 l=180
+ ad=0 pd=0 as=0 ps=0 
M3037 diff_126600_74280# diff_124080_67440# GND GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M3038 GND diff_131400_70800# diff_130320_71160# GND efet w=5880 l=720
+ ad=0 pd=0 as=0 ps=0 
M3039 diff_143040_93480# diff_95040_69120# diff_151200_67920# GND efet w=1320 l=780
+ ad=0 pd=0 as=1.0512e+07 ps=24720 
M3040 diff_132480_78480# diff_105000_78480# diff_145440_75120# GND efet w=2760 l=840
+ ad=0 pd=0 as=7.6752e+06 ps=18000 
M3041 diff_145440_75120# diff_141240_74160# GND GND efet w=5040 l=720
+ ad=0 pd=0 as=0 ps=0 
M3042 GND diff_154080_74280# diff_143040_93480# GND efet w=2400 l=720
+ ad=0 pd=0 as=0 ps=0 
M3043 GND diff_159000_76200# diff_159840_82560# GND efet w=2400 l=780
+ ad=0 pd=0 as=0 ps=0 
M3044 diff_159000_76200# diff_159000_76200# diff_159000_76200# GND efet w=120 l=600
+ ad=0 pd=0 as=0 ps=0 
M3045 diff_159000_76200# diff_159000_76200# diff_159000_76200# GND efet w=240 l=420
+ ad=0 pd=0 as=0 ps=0 
M3046 Vdd Vdd diff_166440_78000# GND efet w=840 l=5760
+ ad=0 pd=0 as=5.688e+06 ps=14400 
M3047 diff_159960_78480# Vdd Vdd GND efet w=720 l=4560
+ ad=7.2288e+06 pd=17520 as=0 ps=0 
M3048 diff_159960_78480# diff_159960_78480# diff_159960_78480# GND efet w=180 l=660
+ ad=0 pd=0 as=0 ps=0 
M3049 diff_159960_78480# diff_159960_78480# diff_159960_78480# GND efet w=240 l=420
+ ad=0 pd=0 as=0 ps=0 
M3050 GND diff_159960_78480# diff_166440_78000# GND efet w=1380 l=900
+ ad=0 pd=0 as=0 ps=0 
M3051 GND diff_159960_78480# diff_159000_76200# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M3052 diff_159840_82560# diff_159840_82560# diff_159840_82560# GND efet w=240 l=420
+ ad=0 pd=0 as=0 ps=0 
M3053 diff_159840_82560# diff_159840_82560# diff_159840_82560# GND efet w=240 l=540
+ ad=0 pd=0 as=0 ps=0 
M3054 diff_166440_78000# diff_131520_76200# diff_158880_70800# GND efet w=1380 l=780
+ ad=0 pd=0 as=4.1184e+06 ps=8880 
M3055 Vdd Vdd diff_178440_81000# GND efet w=960 l=3840
+ ad=0 pd=0 as=0 ps=0 
M3056 Vdd Vdd diff_181680_74280# GND efet w=840 l=5760
+ ad=0 pd=0 as=5.76e+06 ps=14400 
M3057 Vdd Vdd diff_187320_82560# GND efet w=1080 l=3720
+ ad=0 pd=0 as=0 ps=0 
M3058 diff_186600_76200# Vdd Vdd GND efet w=660 l=4620
+ ad=7.3152e+06 pd=20160 as=0 ps=0 
M3059 diff_178440_81000# diff_178440_81000# diff_178440_81000# GND efet w=180 l=540
+ ad=0 pd=0 as=0 ps=0 
M3060 diff_178440_81000# diff_178440_81000# diff_178440_81000# GND efet w=300 l=420
+ ad=0 pd=0 as=0 ps=0 
M3061 GND diff_159000_76200# diff_159960_78480# GND efet w=1380 l=720
+ ad=0 pd=0 as=0 ps=0 
M3062 diff_181680_74280# diff_181680_74280# diff_181680_74280# GND efet w=120 l=600
+ ad=0 pd=0 as=0 ps=0 
M3063 diff_181680_74280# diff_181680_74280# diff_181680_74280# GND efet w=240 l=480
+ ad=0 pd=0 as=0 ps=0 
M3064 GND diff_181680_74280# diff_178440_81000# GND efet w=2820 l=780
+ ad=0 pd=0 as=0 ps=0 
M3065 diff_159840_82560# diff_131520_76200# diff_168840_74040# GND efet w=1320 l=720
+ ad=0 pd=0 as=4.1184e+06 ps=8880 
M3066 diff_159000_76200# diff_132480_78480# diff_157800_71160# GND efet w=2940 l=780
+ ad=0 pd=0 as=7.848e+06 ps=17760 
M3067 diff_151200_67920# diff_151200_67920# diff_151200_67920# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M3068 diff_151200_67920# diff_151200_67920# diff_151200_67920# GND efet w=180 l=180
+ ad=0 pd=0 as=0 ps=0 
M3069 diff_96600_67920# diff_96240_67320# diff_34920_109680# GND efet w=1320 l=600
+ ad=0 pd=0 as=0 ps=0 
M3070 diff_124080_67440# diff_96240_67320# diff_25200_276600# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M3071 Vdd Vdd diff_35640_60240# GND efet w=840 l=5880
+ ad=0 pd=0 as=0 ps=0 
M3072 GND GND diff_55440_53520# GND efet w=3840 l=780
+ ad=0 pd=0 as=1.67328e+07 ps=40080 
M3073 diff_35640_60240# clk1 diff_35400_55320# GND efet w=900 l=660
+ ad=0 pd=0 as=2.4624e+06 ps=9120 
M3074 GND diff_23160_135720# diff_55440_53520# GND efet w=8520 l=720
+ ad=0 pd=0 as=0 ps=0 
M3075 diff_35400_55320# diff_35400_55320# diff_35400_55320# GND efet w=420 l=420
+ ad=0 pd=0 as=0 ps=0 
M3076 GND diff_35400_55320# diff_35640_54240# GND efet w=1440 l=660
+ ad=0 pd=0 as=6.6672e+06 ps=15840 
M3077 diff_35400_55320# diff_35400_55320# diff_35400_55320# GND efet w=300 l=480
+ ad=0 pd=0 as=0 ps=0 
M3078 diff_55440_49920# Vdd diff_55440_53520# GND efet w=4140 l=780
+ ad=2.22048e+07 pd=50160 as=0 ps=0 
M3079 Vdd Vdd diff_35640_54240# GND efet w=840 l=5760
+ ad=0 pd=0 as=0 ps=0 
M3080 GND diff_23040_212640# diff_63240_48000# GND efet w=8880 l=840
+ ad=0 pd=0 as=2.45808e+07 ps=49680 
M3081 diff_60480_40320# diff_23040_212640# GND GND efet w=4680 l=840
+ ad=9.3024e+06 pd=23280 as=0 ps=0 
M3082 diff_55440_53520# diff_55080_52800# diff_55440_49920# GND efet w=5400 l=720
+ ad=0 pd=0 as=0 ps=0 
M3083 clk1 GND GND GND efet w=10560 l=600
+ ad=3.75264e+07 pd=63840 as=0 ps=0 
M3084 GND diff_28560_45600# diff_26880_44640# GND efet w=5040 l=720
+ ad=0 pd=0 as=0 ps=0 
M3085 diff_35640_54240# clk2 diff_35280_49320# GND efet w=840 l=600
+ ad=0 pd=0 as=2.5344e+06 ps=9120 
M3086 diff_35280_49320# diff_35280_49320# diff_35280_49320# GND efet w=360 l=360
+ ad=0 pd=0 as=0 ps=0 
M3087 GND diff_35280_49320# diff_35640_48240# GND efet w=1440 l=660
+ ad=0 pd=0 as=6.0336e+06 ps=14640 
M3088 GND diff_23160_135720# diff_55080_52800# GND efet w=4080 l=840
+ ad=0 pd=0 as=4.968e+06 ps=12000 
M3089 diff_56640_92400# diff_56640_92400# diff_56640_92400# GND efet w=420 l=420
+ ad=2.85408e+07 pd=84480 as=0 ps=0 
M3090 diff_56640_92400# diff_56640_92400# diff_56640_92400# GND efet w=300 l=360
+ ad=0 pd=0 as=0 ps=0 
M3091 diff_74400_51600# diff_73320_44160# GND GND efet w=1440 l=720
+ ad=6.048e+06 pd=14400 as=0 ps=0 
M3092 diff_35280_49320# diff_35280_49320# diff_35280_49320# GND efet w=300 l=480
+ ad=0 pd=0 as=0 ps=0 
M3093 GND diff_30720_47640# diff_31080_46560# GND efet w=3480 l=600
+ ad=0 pd=0 as=7.7184e+06 ps=17040 
M3094 Vdd Vdd diff_35640_48240# GND efet w=840 l=5760
+ ad=0 pd=0 as=0 ps=0 
M3095 diff_55080_52800# Vdd Vdd GND efet w=1080 l=3840
+ ad=0 pd=0 as=0 ps=0 
M3096 GND p0 diff_63240_48000# GND efet w=4140 l=780
+ ad=0 pd=0 as=0 ps=0 
M3097 GND p0 diff_65640_39960# GND efet w=1440 l=720
+ ad=0 pd=0 as=5.4288e+06 ps=14880 
M3098 diff_72960_46200# diff_56640_92400# diff_74400_51600# GND efet w=1380 l=780
+ ad=5.7168e+06 pd=14880 as=0 ps=0 
M3099 GND diff_56640_92400# diff_77640_44520# GND efet w=1380 l=900
+ ad=0 pd=0 as=5.1984e+06 ps=13200 
M3100 diff_35640_48240# clk1 diff_30720_47640# GND efet w=1500 l=660
+ ad=0 pd=0 as=2.232e+06 ps=6000 
M3101 diff_28560_45600# diff_28560_45600# diff_28560_45600# GND efet w=240 l=720
+ ad=2.4192e+06 pd=7680 as=0 ps=0 
M3102 diff_26880_44640# Vdd Vdd GND efet w=960 l=1800
+ ad=0 pd=0 as=0 ps=0 
M3103 diff_28560_45600# diff_28560_45600# diff_28560_45600# GND efet w=360 l=360
+ ad=0 pd=0 as=0 ps=0 
M3104 diff_31080_46560# clk2 diff_28560_45600# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M3105 diff_63240_48000# diff_60480_40320# diff_55440_49920# GND efet w=5520 l=840
+ ad=0 pd=0 as=0 ps=0 
M3106 diff_31080_46560# Vdd Vdd GND efet w=1020 l=2700
+ ad=0 pd=0 as=0 ps=0 
M3107 diff_65640_39960# diff_65640_39960# diff_65640_39960# GND efet w=360 l=480
+ ad=0 pd=0 as=0 ps=0 
M3108 diff_73320_44160# diff_72960_46200# GND GND efet w=2460 l=780
+ ad=3.4704e+06 pd=8400 as=0 ps=0 
M3109 diff_65640_39960# diff_65640_39960# diff_65640_39960# GND efet w=300 l=600
+ ad=0 pd=0 as=0 ps=0 
M3110 diff_77640_44520# diff_77640_44520# diff_77640_44520# GND efet w=300 l=360
+ ad=0 pd=0 as=0 ps=0 
M3111 diff_81000_47280# diff_77640_44520# diff_55440_49920# GND efet w=1320 l=840
+ ad=4.4496e+06 pd=12000 as=0 ps=0 
M3112 diff_55440_49920# diff_65640_39960# diff_63240_48000# GND efet w=5400 l=840
+ ad=0 pd=0 as=0 ps=0 
M3113 Vdd Vdd diff_33840_28200# GND efet w=900 l=660
+ ad=0 pd=0 as=2.5632e+06 ps=8400 
M3114 diff_20280_51120# diff_33840_28200# diff_20280_51120# GND efet w=5220 l=1080
+ ad=1.5192e+07 pd=36720 as=0 ps=0 
M3115 diff_33840_28200# diff_33840_28200# diff_33840_28200# GND efet w=300 l=540
+ ad=0 pd=0 as=0 ps=0 
M3116 diff_33840_28200# diff_33840_28200# diff_33840_28200# GND efet w=120 l=480
+ ad=0 pd=0 as=0 ps=0 
M3117 diff_20280_51120# diff_33840_28200# Vdd GND efet w=1200 l=2040
+ ad=0 pd=0 as=0 ps=0 
M3118 Vdd Vdd diff_36600_23040# GND efet w=840 l=5760
+ ad=0 pd=0 as=3.9456e+06 ps=9360 
M3119 Vdd diff_47760_32880# diff_13200_279960# GND efet w=2040 l=660
+ ad=0 pd=0 as=3.72816e+07 ps=94560 
M3120 diff_13200_279960# diff_46080_27240# GND GND efet w=1920 l=720
+ ad=0 pd=0 as=0 ps=0 
M3121 diff_36600_23040# clk1 diff_41400_25920# GND efet w=2760 l=840
+ ad=0 pd=0 as=4.32e+06 ps=9600 
M3122 diff_20280_51120# diff_36600_23040# GND GND efet w=4440 l=660
+ ad=0 pd=0 as=0 ps=0 
M3123 diff_41400_25920# diff_41040_25200# GND GND efet w=2640 l=720
+ ad=0 pd=0 as=0 ps=0 
M3124 Vdd Vdd diff_46080_27240# GND efet w=840 l=5760
+ ad=0 pd=0 as=3.9456e+06 ps=9120 
M3125 diff_60480_40320# Vdd Vdd GND efet w=960 l=3120
+ ad=0 pd=0 as=0 ps=0 
M3126 Vdd Vdd diff_55440_49920# GND efet w=1080 l=3960
+ ad=0 pd=0 as=0 ps=0 
M3127 diff_65640_39960# Vdd Vdd GND efet w=840 l=5820
+ ad=0 pd=0 as=0 ps=0 
M3128 diff_77640_44520# diff_77640_44520# diff_77640_44520# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M3129 diff_154080_74280# diff_151200_67920# GND GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M3130 GND diff_158880_70800# diff_157800_71160# GND efet w=5700 l=780
+ ad=0 pd=0 as=0 ps=0 
M3131 diff_178440_81000# diff_95040_69120# diff_179040_69240# GND efet w=1440 l=780
+ ad=0 pd=0 as=1.03392e+07 ps=23280 
M3132 diff_159960_78480# diff_132480_78480# diff_173040_74640# GND efet w=2640 l=720
+ ad=0 pd=0 as=7.2144e+06 ps=17520 
M3133 diff_173040_74640# diff_168840_74040# GND GND efet w=5040 l=720
+ ad=0 pd=0 as=0 ps=0 
M3134 diff_187320_82560# diff_186600_76200# GND GND efet w=2520 l=720
+ ad=0 pd=0 as=0 ps=0 
M3135 diff_186600_76200# diff_186600_76200# diff_186600_76200# GND efet w=180 l=660
+ ad=0 pd=0 as=0 ps=0 
M3136 diff_186600_76200# diff_186600_76200# diff_186600_76200# GND efet w=300 l=360
+ ad=0 pd=0 as=0 ps=0 
M3137 Vdd Vdd diff_194040_77880# GND efet w=840 l=5760
+ ad=0 pd=0 as=5.5584e+06 ps=14160 
M3138 diff_187440_78480# Vdd Vdd GND efet w=720 l=5100
+ ad=7.6752e+06 pd=18960 as=0 ps=0 
M3139 diff_187440_78480# diff_187440_78480# diff_187440_78480# GND efet w=120 l=600
+ ad=0 pd=0 as=0 ps=0 
M3140 diff_187440_78480# diff_187440_78480# diff_187440_78480# GND efet w=300 l=360
+ ad=0 pd=0 as=0 ps=0 
M3141 GND diff_187440_78480# diff_194040_77880# GND efet w=1320 l=840
+ ad=0 pd=0 as=0 ps=0 
M3142 GND diff_187440_78480# diff_186600_76200# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M3143 diff_187320_82560# diff_187320_82560# diff_187320_82560# GND efet w=180 l=300
+ ad=0 pd=0 as=0 ps=0 
M3144 diff_187320_82560# diff_187320_82560# diff_187320_82560# GND efet w=300 l=360
+ ad=0 pd=0 as=0 ps=0 
M3145 GND diff_186600_76200# diff_187440_78480# GND efet w=1440 l=720
+ ad=0 pd=0 as=0 ps=0 
M3146 diff_194040_77880# diff_159000_76200# diff_186480_70800# GND efet w=1380 l=780
+ ad=0 pd=0 as=4.1616e+06 ps=9120 
M3147 diff_187320_82560# diff_159000_76200# diff_196320_74400# GND efet w=1440 l=720
+ ad=0 pd=0 as=4.4352e+06 ps=9120 
M3148 diff_186600_76200# diff_159960_78480# diff_185280_73440# GND efet w=2640 l=720
+ ad=0 pd=0 as=8.0496e+06 ps=18000 
M3149 diff_179040_69240# diff_179040_69240# diff_179040_69240# GND efet w=360 l=360
+ ad=0 pd=0 as=0 ps=0 
M3150 diff_179040_69240# diff_179040_69240# diff_179040_69240# GND efet w=240 l=240
+ ad=0 pd=0 as=0 ps=0 
M3151 diff_181680_74280# diff_179040_69240# GND GND efet w=2280 l=720
+ ad=0 pd=0 as=0 ps=0 
M3152 GND diff_186480_70800# diff_185280_73440# GND efet w=5760 l=720
+ ad=0 pd=0 as=0 ps=0 
M3153 diff_187440_78480# diff_159960_78480# diff_200640_74640# GND efet w=2640 l=720
+ ad=0 pd=0 as=7.2576e+06 ps=18000 
M3154 GND diff_196320_74400# diff_200640_74640# GND efet w=5280 l=720
+ ad=0 pd=0 as=0 ps=0 
M3155 diff_179040_69240# diff_96240_67320# diff_23160_135720# GND efet w=1740 l=720
+ ad=0 pd=0 as=0 ps=0 
M3156 GND diff_188760_69960# diff_189240_66360# GND efet w=6480 l=720
+ ad=0 pd=0 as=2.42784e+07 ps=58080 
M3157 diff_151200_67920# diff_96240_67320# diff_23040_212640# GND efet w=1320 l=720
+ ad=0 pd=0 as=0 ps=0 
M3158 diff_189240_66360# diff_188760_65280# diff_189240_66360# GND efet w=4320 l=2160
+ ad=0 pd=0 as=0 ps=0 
M3159 diff_164040_60000# Vdd Vdd GND efet w=1140 l=3480
+ ad=6.9696e+06 pd=14880 as=0 ps=0 
M3160 diff_189240_66360# diff_188760_65280# Vdd GND efet w=1020 l=1140
+ ad=0 pd=0 as=0 ps=0 
M3161 GND diff_73320_44160# diff_85080_45720# GND efet w=3480 l=720
+ ad=0 pd=0 as=9.5184e+06 ps=20880 
M3162 diff_108600_45960# diff_81000_47280# GND GND efet w=2400 l=720
+ ad=8.2944e+06 pd=21600 as=0 ps=0 
M3163 Vdd Vdd diff_169200_62280# GND efet w=1080 l=1920
+ ad=0 pd=0 as=0 ps=0 
M3164 diff_188760_65280# diff_188760_65280# diff_188760_65280# GND efet w=120 l=480
+ ad=2.2032e+06 pd=7440 as=0 ps=0 
M3165 diff_188760_65280# diff_188760_65280# diff_188760_65280# GND efet w=300 l=420
+ ad=0 pd=0 as=0 ps=0 
M3166 diff_173760_44760# Vdd Vdd GND efet w=1080 l=3840
+ ad=1.1232e+07 pd=29280 as=0 ps=0 
M3167 Vdd Vdd diff_179040_45000# GND efet w=1020 l=3780
+ ad=0 pd=0 as=1.44288e+07 ps=36240 
M3168 diff_158880_60960# diff_85080_45720# diff_23040_212640# GND efet w=1320 l=720
+ ad=2.0736e+06 pd=6000 as=0 ps=0 
M3169 diff_164040_60000# diff_164040_60000# diff_164040_60000# GND efet w=180 l=300
+ ad=0 pd=0 as=0 ps=0 
M3170 diff_169200_62280# diff_164040_60000# GND GND efet w=5820 l=780
+ ad=0 pd=0 as=0 ps=0 
M3171 diff_169200_62280# diff_169200_62280# diff_169200_62280# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M3172 diff_173760_44760# diff_169200_62280# GND GND efet w=3240 l=720
+ ad=0 pd=0 as=0 ps=0 
M3173 diff_169200_62280# diff_169200_62280# diff_169200_62280# GND efet w=240 l=360
+ ad=0 pd=0 as=0 ps=0 
M3174 diff_164040_60000# diff_164040_60000# diff_164040_60000# GND efet w=180 l=180
+ ad=0 pd=0 as=0 ps=0 
M3175 diff_25200_276600# diff_85080_45720# diff_142440_51840# GND efet w=1320 l=720
+ ad=0 pd=0 as=2.5344e+06 ps=6480 
M3176 diff_34920_109680# diff_85080_45720# diff_148320_51840# GND efet w=1320 l=720
+ ad=0 pd=0 as=2.5344e+06 ps=6480 
M3177 GND diff_38640_64440# diff_81000_47280# GND efet w=1500 l=780
+ ad=0 pd=0 as=0 ps=0 
M3178 diff_108600_45960# diff_108600_45960# diff_108600_45960# GND efet w=660 l=420
+ ad=0 pd=0 as=0 ps=0 
M3179 diff_108600_45960# diff_98040_40560# GND GND efet w=1440 l=840
+ ad=0 pd=0 as=0 ps=0 
M3180 GND clk2 diff_117120_48960# GND efet w=2280 l=840
+ ad=0 pd=0 as=3.0672e+06 ps=8160 
M3181 diff_108600_45960# diff_108600_45960# diff_108600_45960# GND efet w=420 l=900
+ ad=0 pd=0 as=0 ps=0 
M3182 GND diff_108600_45960# diff_111840_45720# GND efet w=1380 l=780
+ ad=0 pd=0 as=2.592e+06 ps=6960 
M3183 diff_117120_48960# diff_66120_24960# diff_117120_47280# GND efet w=3060 l=780
+ ad=0 pd=0 as=2.5344e+06 ps=7920 
M3184 diff_117120_47280# diff_111840_45720# diff_117120_45480# GND efet w=3000 l=840
+ ad=0 pd=0 as=7.1424e+06 ps=15600 
M3185 diff_73320_44160# Vdd Vdd GND efet w=840 l=5760
+ ad=0 pd=0 as=0 ps=0 
M3186 diff_74400_51600# Vdd Vdd GND efet w=840 l=5700
+ ad=0 pd=0 as=0 ps=0 
M3187 diff_77640_44520# Vdd Vdd GND efet w=840 l=5760
+ ad=0 pd=0 as=0 ps=0 
M3188 diff_55440_49920# diff_77640_44520# diff_72960_46200# GND efet w=1440 l=840
+ ad=0 pd=0 as=0 ps=0 
M3189 GND diff_87360_43320# diff_85080_45720# GND efet w=3360 l=720
+ ad=0 pd=0 as=0 ps=0 
M3190 diff_95160_41640# clk2 diff_56640_92400# GND efet w=3120 l=840
+ ad=4.1904e+06 pd=10080 as=0 ps=0 
M3191 diff_85080_45720# Vdd Vdd GND efet w=960 l=2880
+ ad=0 pd=0 as=0 ps=0 
M3192 diff_56640_92400# Vdd Vdd GND efet w=840 l=5760
+ ad=0 pd=0 as=0 ps=0 
M3193 diff_46080_27240# diff_47760_32880# GND GND efet w=1440 l=840
+ ad=0 pd=0 as=0 ps=0 
M3194 Vdd Vdd diff_47760_32880# GND efet w=840 l=5760
+ ad=0 pd=0 as=9.6768e+06 ps=19200 
M3195 diff_54960_30360# Vdd Vdd GND efet w=720 l=5520
+ ad=2.952e+06 pd=8160 as=0 ps=0 
M3196 Vdd Vdd diff_58800_24960# GND efet w=720 l=4560
+ ad=0 pd=0 as=8.8848e+06 ps=17520 
M3197 diff_62760_30240# diff_41040_25200# Vdd GND efet w=1380 l=780
+ ad=2.7792e+06 pd=7440 as=0 ps=0 
M3198 diff_62760_30240# clk1 diff_61200_23040# GND efet w=840 l=720
+ ad=0 pd=0 as=6.3072e+06 ps=14400 
M3199 GND diff_69720_28560# diff_54960_30360# GND efet w=1260 l=900
+ ad=0 pd=0 as=0 ps=0 
M3200 diff_61200_23040# diff_61200_23040# diff_61200_23040# GND efet w=420 l=420
+ ad=0 pd=0 as=0 ps=0 
M3201 diff_61200_23040# diff_61200_23040# diff_61200_23040# GND efet w=240 l=600
+ ad=0 pd=0 as=0 ps=0 
M3202 diff_58800_24960# diff_58800_24960# diff_58800_24960# GND efet w=420 l=420
+ ad=0 pd=0 as=0 ps=0 
M3203 GND diff_61200_23040# diff_58800_24960# GND efet w=4260 l=780
+ ad=0 pd=0 as=0 ps=0 
M3204 diff_58800_24960# diff_58800_24960# diff_58800_24960# GND efet w=180 l=960
+ ad=0 pd=0 as=0 ps=0 
M3205 GND diff_66120_24960# diff_61200_23040# GND efet w=1620 l=780
+ ad=0 pd=0 as=0 ps=0 
M3206 diff_97080_40800# diff_96240_30240# diff_95160_41640# GND efet w=4020 l=900
+ ad=3.9168e+06 pd=10080 as=0 ps=0 
M3207 GND diff_98040_40560# diff_97080_40800# GND efet w=4080 l=840
+ ad=0 pd=0 as=0 ps=0 
M3208 diff_108600_45960# Vdd Vdd GND efet w=840 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3209 Vdd Vdd diff_41040_25200# GND efet w=960 l=3780
+ ad=0 pd=0 as=6.0624e+06 ps=12960 
M3210 diff_104040_40440# diff_98040_40560# diff_87360_43320# GND efet w=3120 l=840
+ ad=2.9952e+06 pd=8160 as=5.0976e+06 ps=11280 
M3211 diff_105720_40560# diff_105000_25200# diff_104040_40440# GND efet w=3060 l=780
+ ad=2.7648e+06 pd=8160 as=0 ps=0 
M3212 GND clk2 diff_105720_40560# GND efet w=2340 l=900
+ ad=0 pd=0 as=0 ps=0 
M3213 diff_87360_43320# Vdd Vdd GND efet w=840 l=7440
+ ad=0 pd=0 as=0 ps=0 
M3214 GND diff_78360_22440# diff_41040_25200# GND efet w=2220 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3215 diff_47760_32880# diff_54960_30360# GND GND efet w=1560 l=720
+ ad=0 pd=0 as=0 ps=0 
M3216 GND diff_58800_24960# diff_47760_32880# GND efet w=1560 l=720
+ ad=0 pd=0 as=0 ps=0 
M3217 clk2 GND GND GND efet w=10560 l=840
+ ad=5.32224e+07 pd=91440 as=0 ps=0 
M3218 diff_111840_45720# Vdd Vdd GND efet w=840 l=5880
+ ad=0 pd=0 as=0 ps=0 
M3219 Vdd Vdd diff_117120_45480# GND efet w=840 l=7320
+ ad=0 pd=0 as=0 ps=0 
M3220 diff_96240_67320# diff_117120_45480# GND GND efet w=3480 l=840
+ ad=6.0192e+06 pd=15600 as=0 ps=0 
M3221 diff_95040_69120# diff_95040_69120# diff_95040_69120# GND efet w=180 l=540
+ ad=8.9424e+06 pd=24480 as=0 ps=0 
M3222 diff_95040_69120# diff_95040_69120# diff_95040_69120# GND efet w=360 l=360
+ ad=0 pd=0 as=0 ps=0 
M3223 diff_95040_69120# diff_96240_67320# GND GND efet w=4320 l=840
+ ad=0 pd=0 as=0 ps=0 
M3224 diff_164040_60000# diff_158880_60960# GND GND efet w=4080 l=720
+ ad=0 pd=0 as=0 ps=0 
M3225 Vdd Vdd Vdd GND efet w=240 l=360
+ ad=0 pd=0 as=0 ps=0 
M3226 Vdd Vdd Vdd GND efet w=180 l=180
+ ad=0 pd=0 as=0 ps=0 
M3227 Vdd diff_212400_75480# diff_84480_143520# GND efet w=2220 l=660
+ ad=0 pd=0 as=0 ps=0 
M3228 Vdd Vdd Vdd GND efet w=120 l=300
+ ad=0 pd=0 as=0 ps=0 
M3229 diff_218760_63360# Vdd Vdd GND efet w=1080 l=3720
+ ad=0 pd=0 as=0 ps=0 
M3230 Vdd Vdd Vdd GND efet w=300 l=480
+ ad=0 pd=0 as=0 ps=0 
M3231 Vdd Vdd diff_217080_82200# GND efet w=1080 l=2760
+ ad=0 pd=0 as=7.7184e+06 ps=18000 
M3232 diff_218760_63360# clk1 diff_241800_85320# GND efet w=1440 l=720
+ ad=0 pd=0 as=2.4768e+06 ps=6720 
M3233 GND diff_241800_85320# diff_105000_25200# GND efet w=5100 l=660
+ ad=0 pd=0 as=2.19456e+07 ps=59520 
M3234 Vdd Vdd diff_212280_78840# GND efet w=840 l=720
+ ad=0 pd=0 as=2.16e+06 ps=7680 
M3235 diff_84480_143520# diff_217080_82200# GND GND efet w=2040 l=600
+ ad=0 pd=0 as=0 ps=0 
M3236 diff_217080_82200# diff_217080_82200# diff_217080_82200# GND efet w=240 l=600
+ ad=0 pd=0 as=0 ps=0 
M3237 diff_212280_78840# diff_212280_78840# diff_212280_78840# GND efet w=240 l=600
+ ad=0 pd=0 as=0 ps=0 
M3238 diff_212280_78840# diff_212280_78840# diff_212280_78840# GND efet w=300 l=360
+ ad=0 pd=0 as=0 ps=0 
M3239 diff_219600_75600# clk2 diff_217080_82200# GND efet w=5220 l=660
+ ad=1.30032e+07 pd=25440 as=0 ps=0 
M3240 diff_217080_82200# diff_217080_82200# diff_217080_82200# GND efet w=180 l=420
+ ad=0 pd=0 as=0 ps=0 
M3241 GND diff_217080_82200# diff_212400_75480# GND efet w=2280 l=720
+ ad=0 pd=0 as=1.21104e+07 ps=33600 
M3242 Vdd diff_212280_78840# diff_212400_75480# GND efet w=960 l=2640
+ ad=0 pd=0 as=0 ps=0 
M3243 Vdd Vdd Vdd GND efet w=240 l=420
+ ad=0 pd=0 as=0 ps=0 
M3244 Vdd Vdd Vdd GND efet w=360 l=780
+ ad=0 pd=0 as=0 ps=0 
M3245 diff_105000_25200# Vdd Vdd GND efet w=1080 l=1920
+ ad=0 pd=0 as=0 ps=0 
M3246 GND diff_105000_25200# diff_219600_75600# GND efet w=7200 l=720
+ ad=0 pd=0 as=0 ps=0 
M3247 diff_105000_25200# diff_105000_25200# diff_105000_25200# GND efet w=180 l=600
+ ad=0 pd=0 as=0 ps=0 
M3248 diff_105000_25200# diff_105000_25200# diff_105000_25200# GND efet w=360 l=480
+ ad=0 pd=0 as=0 ps=0 
M3249 diff_105000_25200# clk2 diff_241440_77880# GND efet w=1440 l=660
+ ad=0 pd=0 as=2.5488e+06 ps=6480 
M3250 diff_212400_75480# diff_212280_78840# diff_212400_75480# GND efet w=5340 l=1860
+ ad=0 pd=0 as=0 ps=0 
M3251 GND diff_241440_77880# diff_78360_22440# GND efet w=5220 l=660
+ ad=0 pd=0 as=1.06992e+07 ps=23040 
M3252 Vdd Vdd Vdd GND efet w=180 l=360
+ ad=0 pd=0 as=0 ps=0 
M3253 diff_219600_75600# diff_71400_87600# GND GND efet w=4680 l=720
+ ad=0 pd=0 as=0 ps=0 
M3254 GND diff_210600_67320# diff_212160_65400# GND efet w=10200 l=720
+ ad=0 pd=0 as=1.49472e+07 ps=32400 
M3255 Vdd Vdd Vdd GND efet w=300 l=840
+ ad=0 pd=0 as=0 ps=0 
M3256 diff_78360_22440# Vdd Vdd GND efet w=1080 l=1920
+ ad=0 pd=0 as=0 ps=0 
M3257 diff_78360_22440# clk1 diff_239640_70440# GND efet w=1440 l=720
+ ad=0 pd=0 as=2.4912e+06 ps=6720 
M3258 diff_219240_64080# diff_203520_42720# GND GND efet w=8040 l=720
+ ad=1.91664e+07 pd=37440 as=0 ps=0 
M3259 Vdd Vdd Vdd GND efet w=180 l=300
+ ad=0 pd=0 as=0 ps=0 
M3260 GND diff_239640_70440# diff_88080_99240# GND efet w=5040 l=720
+ ad=0 pd=0 as=1.02672e+07 ps=22080 
M3261 Vdd Vdd Vdd GND efet w=300 l=540
+ ad=0 pd=0 as=0 ps=0 
M3262 diff_88080_99240# Vdd Vdd GND efet w=1080 l=1920
+ ad=0 pd=0 as=0 ps=0 
M3263 diff_219240_64080# diff_190320_40200# GND GND efet w=7920 l=720
+ ad=0 pd=0 as=0 ps=0 
M3264 diff_188760_69960# clk1 diff_212160_65400# GND efet w=7680 l=720
+ ad=8.8848e+06 pd=18240 as=0 ps=0 
M3265 diff_188760_65280# Vdd Vdd GND efet w=840 l=720
+ ad=0 pd=0 as=0 ps=0 
M3266 diff_179040_45000# diff_169200_62280# GND GND efet w=3060 l=780
+ ad=0 pd=0 as=0 ps=0 
M3267 Vdd Vdd Vdd GND efet w=420 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3268 Vdd Vdd Vdd GND efet w=660 l=420
+ ad=0 pd=0 as=0 ps=0 
M3269 GND diff_148920_43440# diff_179040_45000# GND efet w=3060 l=720
+ ad=0 pd=0 as=0 ps=0 
M3270 diff_173760_44760# diff_143520_44160# GND GND efet w=3180 l=780
+ ad=0 pd=0 as=0 ps=0 
M3271 diff_200760_57720# Vdd Vdd GND efet w=780 l=780
+ ad=2.448e+06 pd=7440 as=0 ps=0 
M3272 diff_200760_57720# diff_200760_57720# diff_200760_57720# GND efet w=120 l=480
+ ad=0 pd=0 as=0 ps=0 
M3273 diff_200760_57720# diff_200760_57720# diff_200760_57720# GND efet w=180 l=540
+ ad=0 pd=0 as=0 ps=0 
M3274 diff_21960_94200# diff_200760_57720# diff_21960_94200# GND efet w=6840 l=2280
+ ad=4.14144e+07 pd=108480 as=0 ps=0 
M3275 diff_188760_69960# Vdd Vdd GND efet w=960 l=1920
+ ad=0 pd=0 as=0 ps=0 
M3276 diff_219240_64080# diff_218760_63360# diff_210600_67320# GND efet w=6660 l=780
+ ad=0 pd=0 as=7.3008e+06 ps=15360 
M3277 diff_71400_87600# diff_208200_54000# diff_71400_87600# GND efet w=6660 l=3300
+ ad=3.53232e+07 pd=93120 as=0 ps=0 
M3278 diff_21960_94200# diff_200760_57720# Vdd GND efet w=960 l=1080
+ ad=0 pd=0 as=0 ps=0 
M3279 GND diff_158520_43200# diff_173760_44760# GND efet w=2400 l=960
+ ad=0 pd=0 as=0 ps=0 
M3280 GND diff_38640_64440# diff_133800_46680# GND efet w=1380 l=780
+ ad=0 pd=0 as=2.6928e+06 ps=6720 
M3281 diff_96240_67320# diff_96240_67320# diff_96240_67320# GND efet w=240 l=360
+ ad=0 pd=0 as=0 ps=0 
M3282 diff_96240_67320# diff_96240_67320# diff_96240_67320# GND efet w=180 l=540
+ ad=0 pd=0 as=0 ps=0 
M3283 GND diff_126960_46200# diff_95040_69120# GND efet w=3600 l=720
+ ad=0 pd=0 as=0 ps=0 
M3284 diff_160800_51480# diff_85080_45720# diff_23160_135720# GND efet w=1320 l=720
+ ad=2.0448e+06 pd=7440 as=0 ps=0 
M3285 diff_160800_51480# diff_160800_51480# diff_160800_51480# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M3286 diff_160800_51480# diff_160800_51480# diff_160800_51480# GND efet w=300 l=360
+ ad=0 pd=0 as=0 ps=0 
M3287 diff_133800_46680# diff_85080_45720# Vdd GND efet w=1440 l=780
+ ad=0 pd=0 as=0 ps=0 
M3288 diff_96240_67320# Vdd Vdd GND efet w=1020 l=2940
+ ad=0 pd=0 as=0 ps=0 
M3289 diff_138480_43680# diff_133800_46680# GND GND efet w=6300 l=780
+ ad=6.8688e+06 pd=16080 as=0 ps=0 
M3290 diff_95040_69120# Vdd Vdd GND efet w=1080 l=3120
+ ad=0 pd=0 as=0 ps=0 
M3291 diff_126960_46200# diff_78360_22440# GND GND efet w=3780 l=1020
+ ad=3.4704e+06 pd=8640 as=0 ps=0 
M3292 diff_143520_44160# diff_142440_51840# GND GND efet w=4920 l=720
+ ad=7.6464e+06 pd=17040 as=0 ps=0 
M3293 diff_143520_44160# diff_143520_44160# diff_143520_44160# GND efet w=360 l=360
+ ad=0 pd=0 as=0 ps=0 
M3294 diff_143520_44160# diff_143520_44160# diff_143520_44160# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M3295 diff_148920_43440# diff_143520_44160# GND GND efet w=3240 l=840
+ ad=0 pd=0 as=0 ps=0 
M3296 GND diff_151560_43560# diff_179040_45000# GND efet w=3060 l=780
+ ad=0 pd=0 as=0 ps=0 
M3297 diff_179040_45000# diff_160800_51480# GND GND efet w=5100 l=780
+ ad=0 pd=0 as=0 ps=0 
M3298 GND diff_138480_43680# diff_179040_45000# GND efet w=2460 l=780
+ ad=0 pd=0 as=0 ps=0 
M3299 Vdd Vdd diff_208200_54000# GND efet w=780 l=780
+ ad=0 pd=0 as=2.3904e+06 ps=7920 
M3300 diff_210600_67320# Vdd Vdd GND efet w=1020 l=2820
+ ad=0 pd=0 as=0 ps=0 
M3301 diff_88080_99240# clk2 diff_240120_63120# GND efet w=1440 l=600
+ ad=0 pd=0 as=2.5344e+06 ps=6480 
M3302 GND diff_240120_63120# diff_203520_42720# GND efet w=4140 l=660
+ ad=0 pd=0 as=4.12992e+07 ps=115440 
M3303 Vdd Vdd Vdd GND efet w=180 l=240
+ ad=0 pd=0 as=0 ps=0 
M3304 Vdd Vdd Vdd GND efet w=240 l=300
+ ad=0 pd=0 as=0 ps=0 
M3305 diff_203520_42720# Vdd Vdd GND efet w=1140 l=2820
+ ad=0 pd=0 as=0 ps=0 
M3306 diff_208200_54000# diff_208200_54000# diff_208200_54000# GND efet w=120 l=600
+ ad=0 pd=0 as=0 ps=0 
M3307 diff_208200_54000# diff_208200_54000# diff_208200_54000# GND efet w=240 l=360
+ ad=0 pd=0 as=0 ps=0 
M3308 Vdd Vdd Vdd GND efet w=540 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3309 Vdd Vdd Vdd GND efet w=300 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3310 diff_203520_42720# clk1 diff_237840_55440# GND efet w=1380 l=600
+ ad=0 pd=0 as=2.2608e+06 ps=6240 
M3311 Vdd Vdd diff_207480_277200# GND efet w=1020 l=1920
+ ad=0 pd=0 as=3.46176e+07 ps=83520 
M3312 Vdd diff_208200_54000# diff_71400_87600# GND efet w=960 l=1920
+ ad=0 pd=0 as=0 ps=0 
M3313 diff_21960_94200# diff_197400_51840# GND GND efet w=7560 l=720
+ ad=0 pd=0 as=0 ps=0 
M3314 diff_71400_87600# diff_197400_51840# GND GND efet w=4620 l=660
+ ad=0 pd=0 as=0 ps=0 
M3315 Vdd Vdd diff_207120_49680# GND efet w=960 l=2760
+ ad=0 pd=0 as=6.048e+06 ps=14640 
M3316 GND diff_237840_55440# diff_96240_30240# GND efet w=5340 l=660
+ ad=0 pd=0 as=2.72016e+07 ps=65520 
M3317 Vdd Vdd Vdd GND efet w=300 l=360
+ ad=0 pd=0 as=0 ps=0 
M3318 Vdd Vdd Vdd GND efet w=360 l=780
+ ad=0 pd=0 as=0 ps=0 
M3319 diff_96240_30240# Vdd Vdd GND efet w=1080 l=1920
+ ad=0 pd=0 as=0 ps=0 
M3320 diff_207480_277200# diff_197400_51840# GND GND efet w=5760 l=720
+ ad=0 pd=0 as=0 ps=0 
M3321 diff_179280_49800# diff_160800_51480# GND GND efet w=4920 l=720
+ ad=1.60704e+07 pd=38880 as=0 ps=0 
M3322 GND diff_187080_39600# diff_21960_94200# GND efet w=7200 l=720
+ ad=0 pd=0 as=0 ps=0 
M3323 GND diff_207120_49680# diff_71400_87600# GND efet w=4320 l=720
+ ad=0 pd=0 as=0 ps=0 
M3324 diff_148920_43440# diff_148920_43440# diff_148920_43440# GND efet w=240 l=600
+ ad=0 pd=0 as=0 ps=0 
M3325 GND diff_148320_51840# diff_151560_43560# GND efet w=4500 l=780
+ ad=0 pd=0 as=8.6832e+06 ps=20160 
M3326 Vdd Vdd diff_126960_46200# GND efet w=1020 l=3060
+ ad=0 pd=0 as=0 ps=0 
M3327 diff_138480_43680# Vdd Vdd GND efet w=960 l=2880
+ ad=0 pd=0 as=0 ps=0 
M3328 diff_148920_43440# diff_148920_43440# diff_148920_43440# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M3329 diff_151560_43560# diff_151560_43560# diff_151560_43560# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M3330 diff_143520_44160# Vdd Vdd GND efet w=960 l=3840
+ ad=0 pd=0 as=0 ps=0 
M3331 diff_158520_43200# diff_151560_43560# GND GND efet w=3360 l=840
+ ad=0 pd=0 as=0 ps=0 
M3332 GND diff_160800_51480# diff_162600_41640# GND efet w=4560 l=720
+ ad=0 pd=0 as=7.2e+06 ps=17280 
M3333 diff_158520_43200# diff_158520_43200# diff_158520_43200# GND efet w=180 l=540
+ ad=0 pd=0 as=0 ps=0 
M3334 diff_151560_43560# diff_151560_43560# diff_151560_43560# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M3335 diff_158520_43200# diff_158520_43200# diff_158520_43200# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M3336 diff_69720_28560# diff_162600_41640# GND GND efet w=2520 l=720
+ ad=1.13472e+07 pd=27840 as=0 ps=0 
M3337 GND diff_138480_43680# diff_69720_28560# GND efet w=3300 l=720
+ ad=0 pd=0 as=0 ps=0 
M3338 diff_69720_28560# diff_173760_44760# GND GND efet w=2520 l=840
+ ad=0 pd=0 as=0 ps=0 
M3339 GND diff_138480_43680# diff_179280_49800# GND efet w=3120 l=720
+ ad=0 pd=0 as=0 ps=0 
M3340 diff_179280_49800# diff_179040_45000# GND GND efet w=3180 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3341 diff_69720_28560# diff_69720_28560# diff_69720_28560# GND efet w=240 l=300
+ ad=0 pd=0 as=0 ps=0 
M3342 diff_162600_41640# diff_162600_41640# diff_162600_41640# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M3343 diff_69720_28560# diff_69720_28560# diff_69720_28560# GND efet w=240 l=300
+ ad=0 pd=0 as=0 ps=0 
M3344 diff_148920_43440# Vdd Vdd GND efet w=1080 l=2880
+ ad=0 pd=0 as=0 ps=0 
M3345 diff_162600_41640# diff_162600_41640# diff_162600_41640# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M3346 diff_158520_43200# Vdd Vdd GND efet w=1020 l=3120
+ ad=0 pd=0 as=0 ps=0 
M3347 Vdd Vdd diff_162600_41640# GND efet w=1080 l=3960
+ ad=0 pd=0 as=0 ps=0 
M3348 Vdd Vdd diff_151560_43560# GND efet w=960 l=3960
+ ad=0 pd=0 as=0 ps=0 
M3349 diff_69720_28560# Vdd Vdd GND efet w=960 l=3840
+ ad=0 pd=0 as=0 ps=0 
M3350 GND diff_207120_49680# diff_207480_277200# GND efet w=5400 l=720
+ ad=0 pd=0 as=0 ps=0 
M3351 diff_197400_51840# diff_179280_17640# GND GND efet w=3120 l=720
+ ad=6.336e+06 pd=15840 as=0 ps=0 
M3352 GND diff_203520_42720# diff_21960_94200# GND efet w=5940 l=1140
+ ad=0 pd=0 as=0 ps=0 
M3353 diff_71400_87600# diff_190320_40200# GND GND efet w=4440 l=720
+ ad=0 pd=0 as=0 ps=0 
M3354 GND diff_173760_44760# diff_179280_49800# GND efet w=2580 l=780
+ ad=0 pd=0 as=0 ps=0 
M3355 GND diff_179280_49800# diff_190320_40200# GND efet w=2160 l=720
+ ad=0 pd=0 as=4.7232e+06 ps=10080 
M3356 GND diff_96240_30240# diff_207120_49680# GND efet w=3840 l=720
+ ad=0 pd=0 as=0 ps=0 
M3357 diff_207480_277200# diff_195120_40920# GND GND efet w=5700 l=780
+ ad=0 pd=0 as=0 ps=0 
M3358 GND diff_179040_45000# diff_195120_40920# GND efet w=2160 l=720
+ ad=0 pd=0 as=4.0608e+06 ps=9840 
M3359 diff_179280_49800# Vdd Vdd GND efet w=960 l=3720
+ ad=0 pd=0 as=0 ps=0 
M3360 diff_187080_39600# diff_69720_28560# GND GND efet w=2040 l=840
+ ad=5.0544e+06 pd=9600 as=0 ps=0 
M3361 Vdd Vdd diff_187080_39600# GND efet w=1080 l=5040
+ ad=0 pd=0 as=0 ps=0 
M3362 Vdd Vdd diff_190320_40200# GND efet w=1080 l=4680
+ ad=0 pd=0 as=0 ps=0 
M3363 diff_195120_40920# Vdd Vdd GND efet w=1080 l=4680
+ ad=0 pd=0 as=0 ps=0 
M3364 diff_197400_51840# Vdd Vdd GND efet w=720 l=2340
+ ad=0 pd=0 as=0 ps=0 
M3365 diff_96240_30240# clk2 diff_238320_47040# GND efet w=1440 l=600
+ ad=0 pd=0 as=2.4048e+06 ps=6240 
M3366 Vdd Vdd Vdd GND efet w=180 l=240
+ ad=0 pd=0 as=0 ps=0 
M3367 diff_235920_44880# Vdd Vdd GND efet w=1140 l=5580
+ ad=7.0848e+06 pd=16320 as=0 ps=0 
M3368 GND diff_238320_47040# diff_235920_44880# GND efet w=1800 l=720
+ ad=0 pd=0 as=0 ps=0 
M3369 Vdd Vdd Vdd GND efet w=300 l=420
+ ad=0 pd=0 as=0 ps=0 
M3370 diff_237840_42120# clk1 diff_235920_44880# GND efet w=1320 l=720
+ ad=2.2176e+06 pd=6000 as=0 ps=0 
M3371 GND diff_237840_42120# diff_66120_24960# GND efet w=5100 l=660
+ ad=0 pd=0 as=8.3664e+06 ps=17520 
M3372 Vdd Vdd Vdd GND efet w=180 l=180
+ ad=0 pd=0 as=0 ps=0 
M3373 Vdd Vdd Vdd GND efet w=300 l=360
+ ad=0 pd=0 as=0 ps=0 
M3374 Vdd Vdd Vdd GND efet w=240 l=600
+ ad=0 pd=0 as=0 ps=0 
M3375 Vdd Vdd Vdd GND efet w=120 l=180
+ ad=0 pd=0 as=0 ps=0 
M3376 diff_179280_17640# Vdd Vdd GND efet w=1080 l=1920
+ ad=2.628e+07 pd=55440 as=0 ps=0 
M3377 diff_66120_24960# Vdd Vdd GND efet w=1080 l=1980
+ ad=0 pd=0 as=0 ps=0 
M3378 Vdd Vdd diff_98040_40560# GND efet w=1080 l=2760
+ ad=0 pd=0 as=7.56e+06 ps=17520 
M3379 Vdd Vdd diff_214320_16200# GND efet w=1320 l=4500
+ ad=0 pd=0 as=8.6976e+06 ps=19440 
M3380 diff_179280_17640# reset GND GND efet w=12600 l=720
+ ad=0 pd=0 as=0 ps=0 
M3381 sync GND GND GND efet w=10560 l=840
+ ad=0 pd=0 as=0 ps=0 
M3382 reset GND GND GND efet w=10800 l=840
+ ad=3.53376e+07 pd=77280 as=0 ps=0 
M3383 GND GND p0 GND efet w=10560 l=840
+ ad=0 pd=0 as=3.11328e+07 ps=74880 
M3384 diff_214320_16200# diff_214320_16200# diff_214320_16200# GND efet w=300 l=300
+ ad=0 pd=0 as=0 ps=0 
M3385 diff_214320_16200# diff_214320_16200# diff_214320_16200# GND efet w=180 l=540
+ ad=0 pd=0 as=0 ps=0 
M3386 diff_98040_40560# diff_214320_16200# GND GND efet w=3840 l=600
+ ad=0 pd=0 as=0 ps=0 
M3387 GND cm diff_214320_16200# GND efet w=5040 l=720
+ ad=0 pd=0 as=0 ps=0 
M3388 cm GND GND GND efet w=10620 l=780
+ ad=3.3768e+07 pd=77760 as=0 ps=0 
C0 metal_241200_4080# gnd! 43.2fF ;**FLOATING
C1 metal_235680_4920# gnd! 46.1fF ;**FLOATING
C2 metal_230160_5160# gnd! 48.2fF ;**FLOATING
C3 metal_224640_6240# gnd! 42.4fF ;**FLOATING
C4 metal_69600_5520# gnd! 6.8fF ;**FLOATING
C5 metal_67560_6360# gnd! 3.8fF ;**FLOATING
C6 metal_66000_7680# gnd! 10.7fF ;**FLOATING
C7 metal_67440_7680# gnd! 26.5fF ;**FLOATING
C8 metal_71760_11160# gnd! 75.9fF ;**FLOATING
C9 metal_15600_16200# gnd! 8.7fF ;**FLOATING
C10 metal_235440_295080# gnd! 54.0fF ;**FLOATING
C11 diff_214320_16200# gnd! 133.4fF
C12 cm gnd! 1276.1fF
C13 reset gnd! 960.4fF
C14 diff_237840_42120# gnd! 73.6fF
C15 diff_235920_44880# gnd! 87.0fF
C16 diff_238320_47040# gnd! 63.2fF
C17 diff_195120_40920# gnd! 186.0fF
C18 diff_162600_41640# gnd! 139.4fF
C19 diff_187080_39600# gnd! 167.8fF
C20 diff_179280_49800# gnd! 307.7fF
C21 diff_207120_49680# gnd! 140.2fF
C22 diff_197400_51840# gnd! 192.1fF
C23 diff_237840_55440# gnd! 70.5fF
C24 diff_240120_63120# gnd! 68.0fF
C25 diff_133800_46680# gnd! 103.6fF
C26 diff_126960_46200# gnd! 97.5fF
C27 diff_138480_43680# gnd! 343.5fF
C28 diff_160800_51480# gnd! 211.7fF
C29 diff_151560_43560# gnd! 281.0fF
C30 diff_208200_54000# gnd! 127.9fF
C31 diff_143520_44160# gnd! 278.3fF
C32 diff_200760_57720# gnd! 120.2fF
C33 diff_190320_40200# gnd! 324.5fF
C34 diff_239640_70440# gnd! 74.3fF
C35 diff_203520_42720# gnd! 844.3fF
C36 diff_219240_64080# gnd! 254.1fF
C37 diff_212160_65400# gnd! 181.9fF
C38 diff_210600_67320# gnd! 178.8fF
C39 diff_241440_77880# gnd! 73.0fF
C40 diff_219600_75600# gnd! 185.5fF
C41 diff_212280_78840# gnd! 122.6fF
C42 diff_217080_82200# gnd! 135.6fF
C43 diff_241800_85320# gnd! 72.3fF
C44 diff_212400_75480# gnd! 242.1fF
C45 diff_179040_45000# gnd! 371.6fF
C46 diff_148320_51840# gnd! 93.8fF
C47 diff_105720_40560# gnd! 35.8fF
C48 diff_104040_40440# gnd! 38.1fF
C49 diff_105000_25200# gnd! 1085.0fF
C50 diff_97080_40800# gnd! 49.2fF
C51 diff_95160_41640# gnd! 51.9fF
C52 diff_58800_24960# gnd! 133.8fF
C53 diff_61200_23040# gnd! 112.4fF
C54 diff_69720_28560# gnd! 683.5fF
C55 diff_62760_30240# gnd! 35.2fF
C56 diff_16320_16920# gnd! 13.7fF ;**FLOATING
C57 diff_15840_18000# gnd! 18.5fF ;**FLOATING
C58 diff_15480_18720# gnd! 100.7fF ;**FLOATING
C59 diff_54960_30360# gnd! 141.2fF
C60 diff_96240_30240# gnd! 1095.7fF
C61 diff_87360_43320# gnd! 139.5fF
C62 diff_117120_47280# gnd! 33.3fF
C63 diff_66120_24960# gnd! 840.1fF
C64 diff_111840_45720# gnd! 83.7fF
C65 diff_117120_48960# gnd! 38.8fF
C66 diff_117120_45480# gnd! 132.4fF
C67 diff_98040_40560# gnd! 826.5fF
C68 diff_142440_51840# gnd! 80.2fF
C69 diff_173760_44760# gnd! 271.8fF
C70 diff_158880_60960# gnd! 74.5fF
C71 diff_164040_60000# gnd! 122.0fF
C72 diff_108600_45960# gnd! 136.2fF
C73 diff_85080_45720# gnd! 568.3fF
C74 diff_188760_65280# gnd! 109.6fF
C75 diff_188760_69960# gnd! 228.3fF
C76 diff_200640_74640# gnd! 90.6fF
C77 diff_196320_74400# gnd! 102.7fF
C78 diff_185280_73440# gnd! 98.5fF
C79 diff_186480_70800# gnd! 104.3fF
C80 diff_194040_77880# gnd! 98.6fF
C81 diff_187440_78480# gnd! 209.8fF
C82 diff_186600_76200# gnd! 249.3fF
C83 diff_173040_74640# gnd! 89.7fF
C84 diff_179040_69240# gnd! 153.6fF
C85 diff_168840_74040# gnd! 99.6fF
C86 diff_41040_25200# gnd! 251.1fF
C87 diff_41400_25920# gnd! 52.8fF
C88 diff_36600_23040# gnd! 105.5fF
C89 diff_46080_27240# gnd! 103.9fF
C90 diff_47760_32880# gnd! 198.5fF
C91 diff_33840_28200# gnd! 118.1fF
C92 diff_81000_47280# gnd! 188.2fF
C93 diff_77640_44520# gnd! 106.3fF
C94 diff_65640_39960# gnd! 112.9fF
C95 diff_72960_46200# gnd! 131.5fF
C96 p0 gnd! 1530.0fF
C97 diff_31080_46560# gnd! 94.1fF
C98 diff_30720_47640# gnd! 72.3fF
C99 diff_35640_48240# gnd! 75.0fF
C100 diff_74400_51600# gnd! 138.1fF
C101 diff_35280_49320# gnd! 54.6fF
C102 diff_28560_45600# gnd! 68.6fF
C103 diff_55080_52800# gnd! 122.2fF
C104 diff_60480_40320# gnd! 222.7fF
C105 diff_73320_44160# gnd! 200.9fF
C106 diff_63240_48000# gnd! 325.1fF
C107 diff_35640_54240# gnd! 82.5fF
C108 diff_55440_49920# gnd! 469.2fF
C109 diff_35400_55320# gnd! 54.2fF
C110 diff_55440_53520# gnd! 207.4fF
C111 diff_35640_60240# gnd! 77.2fF
C112 diff_96240_67320# gnd! 539.1fF
C113 diff_158880_70800# gnd! 106.2fF
C114 diff_157800_71160# gnd! 96.2fF
C115 diff_181680_74280# gnd! 126.7fF
C116 diff_166440_78000# gnd! 97.9fF
C117 diff_159960_78480# gnd! 382.4fF
C118 diff_159000_76200# gnd! 379.1fF
C119 diff_151200_67920# gnd! 157.6fF
C120 diff_145440_75120# gnd! 94.6fF
C121 diff_141240_74160# gnd! 107.0fF
C122 diff_130320_71160# gnd! 97.2fF
C123 diff_131400_70800# gnd! 109.5fF
C124 diff_154080_74280# gnd! 127.9fF
C125 diff_218760_63360# gnd! 604.2fF
C126 diff_243600_92760# gnd! 64.6fF
C127 diff_138960_78000# gnd! 96.5fF
C128 diff_132480_78480# gnd! 388.1fF
C129 diff_131520_76200# gnd! 378.9fF
C130 diff_124080_67440# gnd! 164.9fF
C131 diff_117960_74760# gnd! 97.0fF
C132 diff_113760_74280# gnd! 106.7fF
C133 diff_103920_70800# gnd! 113.6fF
C134 diff_102720_72840# gnd! 99.4fF
C135 diff_126600_74280# gnd! 118.0fF
C136 diff_158520_43200# gnd! 590.1fF
C137 diff_148920_43440# gnd! 590.6fF
C138 diff_187320_82560# gnd! 295.9fF
C139 diff_169200_62280# gnd! 452.7fF
C140 diff_111360_78000# gnd! 102.6fF
C141 diff_105000_78480# gnd! 389.2fF
C142 diff_103920_81600# gnd! 384.7fF
C143 diff_96600_67920# gnd! 159.8fF
C144 diff_90480_74640# gnd! 96.9fF
C145 diff_86280_74040# gnd! 107.1fF
C146 diff_35400_61080# gnd! 59.0fF
C147 diff_37920_64080# gnd! 79.5fF
C148 diff_76440_70800# gnd! 108.3fF
C149 diff_54480_70200# gnd! 96.8fF
C150 diff_37800_73440# gnd! 62.1fF
C151 sync gnd! 1636.2fF
C152 diff_75480_71160# gnd! 85.6fF
C153 diff_95040_69120# gnd! 711.5fF
C154 diff_99120_74280# gnd! 118.0fF
C155 diff_39600_69360# gnd! 213.1fF
C156 diff_54360_73680# gnd! 294.3fF
C157 diff_83880_78000# gnd! 105.3fF
C158 diff_77520_78480# gnd! 387.2fF
C159 diff_76440_81600# gnd! 380.0fF
C160 diff_38640_64440# gnd! 832.0fF
C161 diff_159840_82560# gnd! 384.4fF
C162 diff_132360_82560# gnd! 255.6fF
C163 diff_360_80280# gnd! 1745.2fF ;**FLOATING
C164 diff_23760_86280# gnd! 107.9fF
C165 diff_178440_81000# gnd! 358.3fF
C166 diff_143040_93480# gnd! 288.6fF
C167 diff_104280_82320# gnd! 709.2fF
C168 diff_76800_82320# gnd! 746.0fF
C169 diff_115560_93600# gnd! 281.8fF
C170 diff_88080_94680# gnd! 291.8fF
C171 diff_243600_101280# gnd! 70.8fF
C172 diff_177840_100680# gnd! 79.0fF
C173 diff_170040_100680# gnd! 59.0fF
C174 diff_177360_99960# gnd! 215.2fF
C175 diff_239520_113040# gnd! 131.3fF
C176 diff_187920_102120# gnd! 209.2fF
C177 diff_84840_96840# gnd! 1058.8fF
C178 diff_202080_109320# gnd! 146.1fF
C179 diff_88080_99240# gnd! 1032.6fF
C180 diff_197040_110280# gnd! 138.2fF
C181 diff_189000_112080# gnd! 149.1fF
C182 diff_181920_110280# gnd! 132.1fF
C183 diff_176640_109320# gnd! 133.2fF
C184 diff_169440_110280# gnd! 132.4fF
C185 diff_163320_111840# gnd! 147.8fF
C186 diff_140160_97560# gnd! 167.5fF
C187 diff_155640_110400# gnd! 144.5fF
C188 diff_149640_111600# gnd! 148.7fF
C189 diff_232800_116760# gnd! 106.3fF
C190 diff_169680_101760# gnd! 339.4fF
C191 diff_141960_110280# gnd! 146.6fF
C192 diff_135840_111600# gnd! 148.3fF
C193 diff_128160_110400# gnd! 143.7fF
C194 diff_122160_112080# gnd! 146.6fF
C195 diff_112680_97560# gnd! 178.3fF
C196 diff_114480_110280# gnd! 146.5fF
C197 diff_108360_111840# gnd! 149.4fF
C198 diff_100800_110280# gnd! 145.4fF
C199 diff_94800_111720# gnd! 145.9fF
C200 diff_82440_102720# gnd! 152.7fF
C201 diff_57480_106560# gnd! 142.1fF
C202 diff_21960_99120# gnd! 184.9fF
C203 diff_22440_106560# gnd! 146.3fF
C204 diff_56160_105120# gnd! 125.5fF
C205 diff_87000_110280# gnd! 149.8fF
C206 diff_20280_51120# gnd! 653.3fF
C207 diff_80880_111840# gnd! 148.6fF
C208 diff_57480_108840# gnd! 139.9fF
C209 diff_56640_92400# gnd! 801.8fF
C210 diff_24840_108840# gnd! 67.8fF
C211 diff_21960_110160# gnd! 70.1fF
C212 diff_188880_122040# gnd! 389.5fF
C213 diff_233880_120960# gnd! 166.3fF
C214 diff_88320_120720# gnd! 589.5fF
C215 diff_82200_122760# gnd! 613.9fF
C216 diff_197400_124560# gnd! 277.6fF
C217 diff_230880_118560# gnd! 149.6fF
C218 diff_84000_102000# gnd! 796.0fF
C219 diff_51600_124080# gnd! 293.3fF
C220 diff_196080_127080# gnd! 342.1fF
C221 diff_82200_127320# gnd! 650.4fF
C222 diff_51600_126720# gnd! 326.3fF
C223 diff_190200_129480# gnd! 285.8fF
C224 diff_230520_127080# gnd! 119.9fF
C225 diff_109680_129600# gnd! 631.6fF
C226 diff_207600_131160# gnd! 142.9fF
C227 diff_82200_132000# gnd! 615.4fF
C228 diff_51600_131160# gnd! 207.3fF
C229 diff_73200_125280# gnd! 95.1fF
C230 diff_21960_94200# gnd! 1616.5fF
C231 diff_233520_124920# gnd! 194.7fF
C232 diff_231000_136440# gnd! 254.4fF
C233 diff_78360_22440# gnd! 1317.5fF
C234 diff_234960_145080# gnd! 117.4fF
C235 diff_26880_44640# gnd! 1521.3fF
C236 diff_82440_133920# gnd! 538.3fF
C237 diff_130200_104880# gnd! 469.0fF
C238 diff_51600_133800# gnd! 309.5fF
C239 diff_17040_127440# gnd! 239.3fF
C240 diff_205320_118080# gnd! 412.1fF
C241 diff_201120_122760# gnd! 413.2fF
C242 diff_210600_147600# gnd! 127.9fF
C243 diff_196560_127680# gnd! 359.4fF
C244 diff_189240_116040# gnd! 363.0fF
C245 diff_203760_142200# gnd! 128.2fF
C246 diff_196800_147600# gnd! 125.8fF
C247 diff_182040_114360# gnd! 424.5fF
C248 diff_175920_112080# gnd! 404.2fF
C249 diff_189960_142200# gnd! 133.6fF
C250 diff_183000_147600# gnd! 128.6fF
C251 diff_169200_145080# gnd! 383.5fF
C252 diff_163440_116040# gnd! 364.5fF
C253 diff_176160_142200# gnd! 132.6fF
C254 diff_169200_147600# gnd! 132.7fF
C255 diff_155520_145080# gnd! 367.4fF
C256 diff_149760_115920# gnd! 338.7fF
C257 diff_162480_139680# gnd! 130.0fF
C258 diff_155520_147600# gnd! 129.6fF
C259 diff_141720_145080# gnd! 361.8fF
C260 diff_135960_115920# gnd! 363.0fF
C261 diff_148680_142200# gnd! 133.1fF
C262 diff_141720_147600# gnd! 132.5fF
C263 diff_135000_138960# gnd! 131.0fF
C264 diff_128040_145080# gnd! 353.5fF
C265 diff_122160_115920# gnd! 360.8fF
C266 diff_128040_147600# gnd! 132.6fF
C267 diff_114240_145080# gnd! 359.3fF
C268 diff_108480_116040# gnd! 361.9fF
C269 diff_121200_142200# gnd! 133.3fF
C270 diff_114240_147600# gnd! 132.7fF
C271 diff_100560_145080# gnd! 357.2fF
C272 diff_94680_112080# gnd! 355.8fF
C273 diff_107520_138960# gnd! 133.2fF
C274 diff_100560_147600# gnd! 128.7fF
C275 diff_16320_124440# gnd! 246.9fF
C276 diff_82080_142080# gnd! 1693.1fF
C277 diff_84480_143520# gnd! 1684.2fF
C278 diff_86760_145200# gnd! 360.4fF
C279 diff_81000_115920# gnd! 361.8fF
C280 diff_73200_137520# gnd! 108.3fF
C281 diff_71400_87600# gnd! 1483.9fF
C282 diff_93720_142200# gnd! 133.1fF
C283 diff_86760_147600# gnd! 131.1fF
C284 diff_79800_142440# gnd! 137.8fF
C285 diff_234600_150240# gnd! 155.7fF
C286 diff_234000_148080# gnd! 190.5fF
C287 clk1 gnd! 2731.9fF
C288 diff_214320_155640# gnd! 33.1fF
C289 diff_234240_153840# gnd! 178.6fF
C290 diff_211800_153720# gnd! 69.6fF
C291 diff_214320_158880# gnd! 33.1fF
C292 diff_228240_160560# gnd! 115.1fF
C293 diff_205200_155160# gnd! 29.3fF
C294 diff_204120_153720# gnd! 70.1fF
C295 diff_198000_153720# gnd! 69.0fF
C296 diff_200520_155640# gnd! 32.1fF
C297 diff_211800_162120# gnd! 68.7fF
C298 diff_211800_167760# gnd! 69.5fF
C299 diff_214320_169800# gnd! 33.4fF
C300 diff_179280_17640# gnd! 1138.2fF
C301 diff_214320_173040# gnd! 34.2fF
C302 diff_205200_159240# gnd! 30.4fF
C303 diff_200520_158880# gnd! 33.4fF
C304 diff_204120_162000# gnd! 70.4fF
C305 diff_191400_155040# gnd! 30.5fF
C306 diff_190320_153720# gnd! 72.4fF
C307 diff_184320_153600# gnd! 69.7fF
C308 diff_186720_155640# gnd! 33.6fF
C309 diff_198000_162120# gnd! 68.5fF
C310 diff_205200_169200# gnd! 30.2fF
C311 diff_204120_167880# gnd! 70.1fF
C312 diff_198000_167760# gnd! 69.7fF
C313 diff_200520_169800# gnd! 33.6fF
C314 diff_211800_176400# gnd! 69.2fF
C315 diff_211800_182040# gnd! 70.3fF
C316 diff_214320_183960# gnd! 33.5fF
C317 diff_214320_187320# gnd! 33.4fF
C318 o3 gnd! 1012.9fF
C319 diff_205200_173400# gnd! 30.4fF
C320 diff_200520_173040# gnd! 33.9fF
C321 diff_204120_176160# gnd! 72.0fF
C322 diff_191400_159240# gnd! 30.7fF
C323 diff_186720_158880# gnd! 33.5fF
C324 diff_190320_162000# gnd! 70.1fF
C325 diff_177600_155040# gnd! 30.8fF
C326 diff_176520_153840# gnd! 71.5fF
C327 diff_173040_155520# gnd! 30.9fF
C328 diff_170520_153600# gnd! 69.8fF
C329 diff_184320_162120# gnd! 68.0fF
C330 diff_191400_169200# gnd! 30.8fF
C331 diff_190320_167880# gnd! 70.3fF
C332 diff_184320_167760# gnd! 68.5fF
C333 diff_186720_169800# gnd! 33.9fF
C334 diff_198000_176400# gnd! 69.7fF
C335 diff_205200_183480# gnd! 30.4fF
C336 diff_200520_183960# gnd! 33.5fF
C337 diff_204120_182040# gnd! 69.9fF
C338 diff_198000_182040# gnd! 68.5fF
C339 diff_211800_190560# gnd! 67.5fF
C340 diff_211800_196200# gnd! 68.1fF
C341 diff_214320_198240# gnd! 33.6fF
C342 diff_237480_200400# gnd! 222.4fF
C343 diff_245520_206640# gnd! 80.5fF
C344 diff_242520_208920# gnd! 70.7fF
C345 diff_214320_201480# gnd! 33.9fF
C346 diff_205200_187560# gnd! 29.4fF
C347 diff_200520_187320# gnd! 33.6fF
C348 diff_204120_190320# gnd! 68.5fF
C349 diff_191400_173400# gnd! 30.7fF
C350 diff_186720_173040# gnd! 34.0fF
C351 diff_190320_176160# gnd! 70.3fF
C352 diff_177600_159240# gnd! 30.8fF
C353 diff_173040_158880# gnd! 30.8fF
C354 diff_176520_162120# gnd! 69.3fF
C355 diff_163800_155040# gnd! 31.2fF
C356 diff_159240_155520# gnd! 30.8fF
C357 diff_162840_153720# gnd! 69.8fF
C358 diff_156720_153600# gnd! 72.7fF
C359 diff_170520_162120# gnd! 66.8fF
C360 diff_163800_159240# gnd! 31.3fF
C361 diff_159240_158880# gnd! 30.8fF
C362 diff_162840_162000# gnd! 68.1fF
C363 diff_177600_169200# gnd! 30.8fF
C364 diff_176520_167880# gnd! 69.1fF
C365 diff_170520_167760# gnd! 67.9fF
C366 diff_173040_169680# gnd! 30.9fF
C367 diff_184320_176280# gnd! 70.4fF
C368 diff_191400_183480# gnd! 30.8fF
C369 diff_184320_181920# gnd! 69.7fF
C370 diff_186720_183960# gnd! 33.8fF
C371 diff_190320_182040# gnd! 70.1fF
C372 diff_198000_190560# gnd! 69.4fF
C373 diff_205200_197640# gnd! 30.6fF
C374 diff_204120_196200# gnd! 68.3fF
C375 diff_200520_198240# gnd! 33.4fF
C376 diff_198000_196200# gnd! 68.8fF
C377 diff_211800_204840# gnd! 68.4fF
C378 diff_214320_212400# gnd! 33.5fF
C379 diff_234480_214080# gnd! 310.7fF
C380 diff_232560_214800# gnd! 34.6fF
C381 diff_211800_210480# gnd! 69.1fF
C382 diff_241680_195480# gnd! 394.4fF
C383 diff_214320_215760# gnd! 32.6fF
C384 diff_205200_201840# gnd! 30.4fF
C385 diff_200520_201480# gnd! 33.9fF
C386 diff_204120_204480# gnd! 68.9fF
C387 diff_191400_187560# gnd! 31.8fF
C388 diff_186720_187200# gnd! 34.6fF
C389 diff_190320_190320# gnd! 70.0fF
C390 diff_177600_173400# gnd! 31.2fF
C391 diff_173040_173040# gnd! 29.5fF
C392 diff_176520_176280# gnd! 71.1fF
C393 diff_150120_155160# gnd! 30.9fF
C394 diff_149040_153720# gnd! 73.6fF
C395 diff_145440_155640# gnd! 33.3fF
C396 diff_143040_153600# gnd! 69.6fF
C397 diff_156720_162120# gnd! 70.0fF
C398 diff_163800_169200# gnd! 30.9fF
C399 diff_162840_167760# gnd! 68.3fF
C400 diff_159240_169680# gnd! 30.6fF
C401 diff_156720_167760# gnd! 71.2fF
C402 diff_163800_173400# gnd! 32.6fF
C403 diff_170520_176400# gnd! 69.3fF
C404 diff_159240_173040# gnd! 31.2fF
C405 diff_162840_176040# gnd! 69.5fF
C406 diff_177600_183360# gnd! 31.5fF
C407 diff_176520_182280# gnd! 70.6fF
C408 diff_170520_181920# gnd! 69.2fF
C409 diff_173040_183840# gnd! 31.5fF
C410 diff_184320_190560# gnd! 68.8fF
C411 diff_191400_197640# gnd! 30.6fF
C412 diff_190320_196200# gnd! 68.8fF
C413 diff_184320_196200# gnd! 68.3fF
C414 diff_186720_198240# gnd! 33.9fF
C415 diff_198000_204720# gnd! 68.2fF
C416 diff_205200_211920# gnd! 30.4fF
C417 diff_200520_212400# gnd! 33.4fF
C418 diff_204120_210360# gnd! 69.9fF
C419 diff_198000_210480# gnd! 70.2fF
C420 diff_211800_219000# gnd! 67.9fF
C421 diff_211800_224520# gnd! 68.5fF
C422 diff_214320_226560# gnd! 32.9fF
C423 diff_214320_229800# gnd! 33.9fF
C424 diff_205200_216000# gnd! 29.4fF
C425 diff_200520_215760# gnd! 32.9fF
C426 diff_204120_218760# gnd! 70.1fF
C427 diff_191400_201840# gnd! 30.7fF
C428 diff_186720_201480# gnd! 33.9fF
C429 diff_190320_204480# gnd! 70.4fF
C430 diff_177600_187560# gnd! 31.9fF
C431 diff_173040_187200# gnd! 31.8fF
C432 diff_176520_190440# gnd! 68.4fF
C433 diff_150120_159240# gnd! 30.5fF
C434 diff_145440_158880# gnd! 33.6fF
C435 diff_149040_162000# gnd! 72.0fF
C436 diff_136320_155160# gnd! 30.4fF
C437 diff_135360_153720# gnd! 71.2fF
C438 diff_129240_153600# gnd! 71.8fF
C439 diff_131760_155520# gnd! 30.9fF
C440 diff_143040_162120# gnd! 69.2fF
C441 diff_150120_169200# gnd! 30.8fF
C442 diff_149040_167760# gnd! 70.7fF
C443 diff_143040_167760# gnd! 67.9fF
C444 diff_145440_169680# gnd! 33.5fF
C445 diff_156720_176400# gnd! 72.5fF
C446 diff_163800_183360# gnd! 34.2fF
C447 diff_162840_181920# gnd! 69.0fF
C448 diff_156720_181920# gnd! 71.6fF
C449 diff_159240_183840# gnd! 31.4fF
C450 diff_170520_190440# gnd! 69.4fF
C451 diff_177600_197640# gnd! 31.1fF
C452 diff_176640_196080# gnd! 69.4fF
C453 diff_170520_196200# gnd! 66.5fF
C454 diff_173040_198120# gnd! 31.2fF
C455 diff_184320_204720# gnd! 69.0fF
C456 diff_191400_211920# gnd! 30.7fF
C457 diff_190320_210360# gnd! 70.0fF
C458 diff_184320_210360# gnd! 68.9fF
C459 diff_186720_212400# gnd! 33.5fF
C460 diff_198000_219000# gnd! 68.8fF
C461 diff_205200_225960# gnd! 30.3fF
C462 diff_204120_224640# gnd! 70.3fF
C463 diff_200520_226560# gnd! 33.6fF
C464 diff_198000_224520# gnd! 69.6fF
C465 diff_211800_233040# gnd! 68.0fF
C466 diff_211800_238680# gnd! 68.1fF
C467 diff_214320_240720# gnd! 33.6fF
C468 o2 gnd! 1004.4fF
C469 diff_237480_243480# gnd! 218.7fF
C470 diff_214320_243960# gnd! 33.5fF
C471 diff_245520_249480# gnd! 77.6fF
C472 diff_242400_251880# gnd! 75.6fF
C473 diff_205200_230160# gnd! 30.4fF
C474 diff_200520_229800# gnd! 33.9fF
C475 diff_204120_232920# gnd! 69.5fF
C476 diff_191400_216000# gnd! 30.4fF
C477 diff_186720_215640# gnd! 33.5fF
C478 diff_190320_218760# gnd! 69.2fF
C479 diff_173040_201480# gnd! 29.1fF
C480 diff_177600_201840# gnd! 31.2fF
C481 diff_176640_204480# gnd! 69.8fF
C482 diff_163800_187560# gnd! 34.7fF
C483 diff_159240_187200# gnd! 31.9fF
C484 diff_162840_190320# gnd! 67.6fF
C485 diff_150120_173400# gnd! 30.5fF
C486 diff_145440_173040# gnd! 33.6fF
C487 diff_149040_176160# gnd! 71.7fF
C488 diff_136320_159240# gnd! 30.5fF
C489 diff_131760_158880# gnd! 30.8fF
C490 diff_135360_162000# gnd! 70.7fF
C491 diff_136320_169200# gnd! 30.8fF
C492 diff_135360_167760# gnd! 69.5fF
C493 diff_122640_155040# gnd! 31.4fF
C494 diff_121560_153720# gnd! 72.8fF
C495 diff_118080_155400# gnd! 31.4fF
C496 diff_115560_153600# gnd! 70.1fF
C497 diff_129240_162120# gnd! 71.2fF
C498 diff_129240_167760# gnd! 69.1fF
C499 diff_131760_169680# gnd! 31.1fF
C500 diff_143040_176400# gnd! 69.0fF
C501 diff_136320_173400# gnd! 30.7fF
C502 diff_131760_173040# gnd! 31.2fF
C503 diff_135360_176040# gnd! 70.3fF
C504 diff_150120_183480# gnd! 30.8fF
C505 diff_149040_181920# gnd! 70.9fF
C506 diff_143040_181920# gnd! 70.0fF
C507 diff_145440_183960# gnd! 33.6fF
C508 diff_156720_190440# gnd! 71.7fF
C509 diff_163800_197640# gnd! 33.3fF
C510 diff_162840_196200# gnd! 66.7fF
C511 diff_159240_198120# gnd! 30.6fF
C512 diff_156720_196200# gnd! 71.3fF
C513 diff_170520_204720# gnd! 67.8fF
C514 diff_177600_211800# gnd! 31.4fF
C515 diff_176520_210960# gnd! 69.3fF
C516 diff_170520_210360# gnd! 67.6fF
C517 diff_173040_212280# gnd! 31.7fF
C518 diff_184320_218880# gnd! 68.2fF
C519 diff_191400_225960# gnd! 30.9fF
C520 diff_190320_224640# gnd! 70.9fF
C521 diff_184200_225120# gnd! 69.9fF
C522 diff_186720_226560# gnd! 33.4fF
C523 diff_198000_233040# gnd! 68.6fF
C524 diff_205200_240240# gnd! 29.2fF
C525 diff_204120_238680# gnd! 69.8fF
C526 diff_198000_238680# gnd! 68.9fF
C527 diff_200520_240720# gnd! 32.9fF
C528 diff_211800_247200# gnd! 67.2fF
C529 diff_211800_252840# gnd! 68.3fF
C530 diff_214320_254880# gnd! 27.5fF
C531 diff_234480_257040# gnd! 307.1fF
C532 diff_232560_257640# gnd! 34.9fF
C533 diff_241440_260160# gnd! 388.5fF
C534 diff_222480_158400# gnd! 794.2fF
C535 diff_214320_258120# gnd! 34.5fF
C536 diff_205080_245640# gnd! 31.2fF
C537 diff_200520_243960# gnd! 33.7fF
C538 diff_204120_247080# gnd! 68.8fF
C539 diff_191400_230160# gnd! 30.7fF
C540 diff_186720_229800# gnd! 34.0fF
C541 diff_190320_232920# gnd! 69.5fF
C542 diff_177600_216000# gnd! 30.8fF
C543 diff_172920_215880# gnd! 31.6fF
C544 diff_176520_218880# gnd! 68.8fF
C545 diff_163800_201840# gnd! 34.0fF
C546 diff_159240_201480# gnd! 31.2fF
C547 diff_162840_204480# gnd! 68.2fF
C548 diff_150120_187560# gnd! 31.6fF
C549 diff_145440_187200# gnd! 34.9fF
C550 diff_149040_190320# gnd! 70.6fF
C551 diff_122640_159240# gnd! 30.7fF
C552 diff_118080_158880# gnd! 30.6fF
C553 diff_121560_162000# gnd! 72.4fF
C554 diff_108840_155040# gnd! 32.6fF
C555 diff_104280_155520# gnd! 31.7fF
C556 diff_107880_153720# gnd! 71.6fF
C557 diff_101880_152880# gnd! 71.9fF
C558 diff_115560_162120# gnd! 69.7fF
C559 diff_108840_159240# gnd! 30.7fF
C560 diff_104280_158880# gnd! 30.8fF
C561 diff_107880_162000# gnd! 70.9fF
C562 diff_122640_169200# gnd! 31.4fF
C563 diff_121560_167760# gnd! 70.8fF
C564 diff_115560_167760# gnd! 68.8fF
C565 diff_118080_169440# gnd! 30.9fF
C566 diff_129240_176400# gnd! 69.0fF
C567 diff_136320_183480# gnd! 30.8fF
C568 diff_135360_181920# gnd! 70.4fF
C569 diff_129240_182040# gnd! 70.7fF
C570 diff_131760_183840# gnd! 30.8fF
C571 diff_143040_190440# gnd! 69.1fF
C572 diff_136320_187560# gnd! 31.9fF
C573 diff_131760_187200# gnd! 29.8fF
C574 diff_135360_190320# gnd! 69.7fF
C575 diff_150120_197640# gnd! 30.6fF
C576 diff_149040_196200# gnd! 70.1fF
C577 diff_145440_198120# gnd! 33.6fF
C578 diff_143040_196080# gnd! 70.4fF
C579 diff_156720_204720# gnd! 70.7fF
C580 diff_163800_211920# gnd! 32.3fF
C581 diff_162840_210360# gnd! 68.4fF
C582 diff_156720_210360# gnd! 71.0fF
C583 diff_159240_212280# gnd! 30.8fF
C584 diff_159240_215640# gnd! 30.7fF
C585 diff_163800_216000# gnd! 31.1fF
C586 diff_170520_218880# gnd! 67.1fF
C587 diff_162840_218760# gnd! 67.7fF
C588 diff_177600_225960# gnd! 30.7fF
C589 diff_176520_224640# gnd! 69.5fF
C590 diff_170520_224520# gnd! 69.9fF
C591 diff_172920_226440# gnd! 33.0fF
C592 diff_184200_233400# gnd! 67.9fF
C593 diff_191400_240120# gnd! 30.9fF
C594 diff_190320_238680# gnd! 69.0fF
C595 diff_184200_238920# gnd! 68.8fF
C596 diff_186720_240720# gnd! 33.5fF
C597 diff_198000_247200# gnd! 68.3fF
C598 diff_205200_254280# gnd! 31.1fF
C599 diff_204120_252840# gnd! 69.7fF
C600 diff_198000_252840# gnd! 68.6fF
C601 diff_200520_254880# gnd! 33.7fF
C602 diff_213360_145800# gnd! 494.7fF
C603 diff_211080_145800# gnd! 457.6fF
C604 diff_208200_149640# gnd! 461.4fF
C605 diff_205200_258480# gnd! 30.4fF
C606 diff_200520_258120# gnd! 33.7fF
C607 diff_204600_144480# gnd! 494.3fF
C608 diff_211800_261480# gnd! 66.7fF
C609 diff_204120_261240# gnd! 67.4fF
C610 diff_199440_146040# gnd! 496.0fF
C611 diff_191400_244320# gnd! 30.7fF
C612 diff_186720_243960# gnd! 34.0fF
C613 diff_190320_247080# gnd! 68.7fF
C614 diff_177600_230160# gnd! 31.0fF
C615 diff_172920_229800# gnd! 33.5fF
C616 diff_176520_232920# gnd! 68.6fF
C617 diff_150120_201840# gnd! 30.5fF
C618 diff_145440_201480# gnd! 33.5fF
C619 diff_149040_204480# gnd! 71.2fF
C620 diff_118080_173040# gnd! 30.7fF
C621 diff_122640_173400# gnd! 31.2fF
C622 diff_121560_176160# gnd! 71.5fF
C623 diff_95160_155040# gnd! 31.6fF
C624 diff_90600_155160# gnd! 31.6fF
C625 diff_94080_153720# gnd! 72.0fF
C626 diff_88080_153600# gnd! 69.3fF
C627 diff_101880_162120# gnd! 71.4fF
C628 diff_108840_169200# gnd! 31.9fF
C629 diff_107880_167760# gnd! 69.3fF
C630 diff_101760_167760# gnd! 70.6fF
C631 diff_104280_169680# gnd! 31.9fF
C632 diff_115560_176280# gnd! 69.3fF
C633 diff_108840_173400# gnd! 31.4fF
C634 diff_104280_173040# gnd! 31.2fF
C635 diff_107880_176160# gnd! 70.8fF
C636 diff_122640_183480# gnd! 30.5fF
C637 diff_115560_181920# gnd! 69.6fF
C638 diff_118080_183720# gnd! 30.7fF
C639 diff_121560_181920# gnd! 71.7fF
C640 diff_129240_190440# gnd! 72.2fF
C641 diff_122640_187560# gnd! 31.5fF
C642 diff_118080_187200# gnd! 31.8fF
C643 diff_121560_190320# gnd! 71.9fF
C644 diff_136320_197640# gnd! 31.1fF
C645 diff_135360_196200# gnd! 70.8fF
C646 diff_129240_196200# gnd! 70.9fF
C647 diff_131760_198120# gnd! 31.3fF
C648 diff_143040_204840# gnd! 69.0fF
C649 diff_136320_201840# gnd! 30.7fF
C650 diff_131760_201480# gnd! 31.2fF
C651 diff_135360_204480# gnd! 69.8fF
C652 diff_150120_211920# gnd! 30.5fF
C653 diff_149040_210360# gnd! 71.5fF
C654 diff_145440_212400# gnd! 33.4fF
C655 diff_143040_210480# gnd! 69.6fF
C656 diff_156720_218880# gnd! 70.6fF
C657 diff_163800_225960# gnd! 31.2fF
C658 diff_162840_224520# gnd! 68.8fF
C659 diff_156720_224520# gnd! 70.4fF
C660 diff_159240_226440# gnd! 30.9fF
C661 diff_170520_233040# gnd! 66.2fF
C662 diff_177600_240120# gnd! 31.1fF
C663 diff_176520_238800# gnd! 70.1fF
C664 diff_170520_238680# gnd! 68.6fF
C665 diff_172920_240720# gnd! 33.7fF
C666 diff_184200_247200# gnd! 68.0fF
C667 diff_191400_254280# gnd! 31.2fF
C668 diff_190320_252960# gnd! 68.6fF
C669 diff_184320_252840# gnd! 68.2fF
C670 diff_186720_254760# gnd! 34.2fF
C671 diff_197280_145800# gnd! 461.8fF
C672 diff_191400_258480# gnd! 31.2fF
C673 diff_186720_258120# gnd! 33.9fF
C674 diff_194400_149640# gnd! 458.2fF
C675 diff_198000_261480# gnd! 68.1fF
C676 diff_190320_261240# gnd! 67.8fF
C677 diff_190800_144240# gnd! 493.2fF
C678 diff_177600_244320# gnd! 30.8fF
C679 diff_172920_243960# gnd! 33.6fF
C680 diff_176520_247080# gnd! 68.7fF
C681 diff_163800_230160# gnd! 30.8fF
C682 diff_159240_229800# gnd! 30.7fF
C683 diff_162840_232800# gnd! 67.0fF
C684 diff_145440_215640# gnd! 33.5fF
C685 diff_150120_216000# gnd! 30.9fF
C686 diff_149040_218760# gnd! 69.1fF
C687 diff_95160_159240# gnd! 30.7fF
C688 diff_90600_158880# gnd! 30.6fF
C689 diff_94080_162000# gnd! 71.9fF
C690 diff_48720_152160# gnd! 137.3fF
C691 diff_50640_154200# gnd! 245.4fF
C692 diff_66480_154320# gnd! 1396.2fF
C693 diff_81480_155160# gnd! 30.7fF
C694 diff_80400_153720# gnd! 72.6fF
C695 diff_88080_162120# gnd! 69.2fF
C696 diff_95160_169200# gnd! 31.8fF
C697 diff_94080_167760# gnd! 69.7fF
C698 diff_88080_167760# gnd! 67.7fF
C699 diff_90600_169320# gnd! 31.0fF
C700 diff_101760_176400# gnd! 72.4fF
C701 diff_108840_183480# gnd! 30.8fF
C702 diff_107880_181920# gnd! 70.0fF
C703 diff_101760_182040# gnd! 70.7fF
C704 diff_104280_183840# gnd! 30.8fF
C705 diff_115560_190440# gnd! 67.7fF
C706 diff_108840_187560# gnd! 32.2fF
C707 diff_104280_187200# gnd! 31.9fF
C708 diff_107880_190320# gnd! 69.5fF
C709 diff_122640_197640# gnd! 31.1fF
C710 diff_121560_196200# gnd! 70.9fF
C711 diff_118080_198000# gnd! 30.7fF
C712 diff_115560_196200# gnd! 69.4fF
C713 diff_129240_204720# gnd! 69.7fF
C714 diff_136320_211920# gnd! 30.7fF
C715 diff_135360_210360# gnd! 69.7fF
C716 diff_129240_210480# gnd! 69.9fF
C717 diff_131760_212280# gnd! 30.7fF
C718 diff_143040_218880# gnd! 67.8fF
C719 diff_136320_216000# gnd! 30.5fF
C720 diff_131760_215640# gnd! 30.9fF
C721 diff_135360_218760# gnd! 68.7fF
C722 diff_150120_225960# gnd! 30.8fF
C723 diff_149040_224640# gnd! 69.8fF
C724 diff_145440_226440# gnd! 33.5fF
C725 diff_143040_224520# gnd! 68.4fF
C726 diff_156720_233040# gnd! 69.1fF
C727 diff_163800_240120# gnd! 30.9fF
C728 diff_162840_238680# gnd! 68.0fF
C729 diff_156720_238680# gnd! 68.7fF
C730 diff_159240_240600# gnd! 31.2fF
C731 diff_170520_247200# gnd! 67.0fF
C732 diff_177600_254280# gnd! 31.2fF
C733 diff_176520_252960# gnd! 69.0fF
C734 diff_170520_252840# gnd! 68.0fF
C735 diff_172920_254760# gnd! 34.2fF
C736 diff_183480_145800# gnd! 500.4fF
C737 diff_180600_149640# gnd! 456.1fF
C738 diff_177000_144360# gnd! 493.2fF
C739 diff_177600_258480# gnd! 31.2fF
C740 diff_172920_258840# gnd! 32.9fF
C741 diff_185640_145800# gnd! 494.7fF
C742 diff_184200_262200# gnd! 67.0fF
C743 diff_176520_261240# gnd! 68.0fF
C744 diff_189240_66360# gnd! 1337.8fF
C745 diff_163800_244320# gnd! 30.8fF
C746 diff_159240_243960# gnd! 30.8fF
C747 diff_162840_247080# gnd! 67.4fF
C748 diff_150120_230160# gnd! 30.8fF
C749 diff_145440_229800# gnd! 33.4fF
C750 diff_149040_232920# gnd! 70.1fF
C751 diff_118080_201480# gnd! 30.6fF
C752 diff_122640_201840# gnd! 31.1fF
C753 diff_121560_204480# gnd! 71.7fF
C754 diff_95160_173400# gnd! 31.8fF
C755 diff_90600_173040# gnd! 31.0fF
C756 diff_94080_176160# gnd! 71.7fF
C757 diff_81360_159720# gnd! 31.3fF
C758 diff_54840_154320# gnd! 1101.4fF
C759 diff_56880_156000# gnd! 197.4fF
C760 diff_80400_162000# gnd! 71.9fF
C761 diff_66480_162000# gnd! 1400.7fF
C762 diff_56880_159960# gnd! 192.5fF
C763 diff_54840_161040# gnd! 1106.0fF
C764 diff_44040_159600# gnd! 67.9fF
C765 diff_50640_161880# gnd! 240.7fF
C766 diff_48720_164160# gnd! 139.7fF
C767 diff_16200_152040# gnd! 115.0fF
C768 diff_16200_162120# gnd! 113.8fF
C769 diff_50640_168360# gnd! 238.3fF
C770 diff_66480_168360# gnd! 1386.0fF
C771 diff_81360_169200# gnd! 34.4fF
C772 diff_80400_167760# gnd! 69.3fF
C773 diff_88080_176280# gnd! 69.2fF
C774 diff_95160_183480# gnd! 30.8fF
C775 diff_94080_181920# gnd! 71.2fF
C776 diff_88080_182040# gnd! 69.4fF
C777 diff_90600_183600# gnd! 30.5fF
C778 diff_101760_190560# gnd! 69.7fF
C779 diff_108840_197640# gnd! 32.2fF
C780 diff_107880_196080# gnd! 71.3fF
C781 diff_101760_196200# gnd! 71.7fF
C782 diff_104280_198120# gnd! 31.8fF
C783 diff_115560_204840# gnd! 68.1fF
C784 diff_108840_201840# gnd! 30.7fF
C785 diff_104280_201480# gnd! 31.2fF
C786 diff_107880_204480# gnd! 69.8fF
C787 diff_122640_211920# gnd! 30.5fF
C788 diff_121560_210360# gnd! 70.8fF
C789 diff_115560_210360# gnd! 68.4fF
C790 diff_118080_212040# gnd! 30.5fF
C791 diff_129240_218880# gnd! 68.9fF
C792 diff_136320_225960# gnd! 30.8fF
C793 diff_135360_224520# gnd! 70.4fF
C794 diff_131760_226440# gnd! 31.1fF
C795 diff_129240_224520# gnd! 69.6fF
C796 diff_143040_233040# gnd! 68.1fF
C797 diff_150000_242040# gnd! 31.0fF
C798 diff_149040_238680# gnd! 69.1fF
C799 diff_145440_240600# gnd! 33.4fF
C800 diff_143040_238680# gnd! 67.7fF
C801 diff_156720_247200# gnd! 67.3fF
C802 diff_163800_254280# gnd! 31.2fF
C803 diff_162840_252840# gnd! 67.4fF
C804 diff_156720_252840# gnd! 69.0fF
C805 diff_159240_254760# gnd! 30.7fF
C806 diff_171960_145800# gnd! 532.1fF
C807 diff_169680_145800# gnd! 456.4fF
C808 diff_166800_149760# gnd! 456.5fF
C809 diff_163800_258480# gnd! 30.8fF
C810 diff_159240_258120# gnd! 30.7fF
C811 diff_163320_144240# gnd! 504.8fF
C812 diff_170520_261360# gnd! 66.5fF
C813 diff_162840_261120# gnd! 67.2fF
C814 diff_158160_145800# gnd! 491.3fF
C815 diff_150120_244320# gnd! 30.7fF
C816 diff_145440_243960# gnd! 33.4fF
C817 diff_149040_247080# gnd! 68.3fF
C818 diff_136320_230160# gnd! 30.5fF
C819 diff_131760_229800# gnd! 31.2fF
C820 diff_135360_232800# gnd! 69.1fF
C821 diff_136320_240120# gnd! 31.2fF
C822 diff_135360_238680# gnd! 68.9fF
C823 diff_118080_215640# gnd! 30.6fF
C824 diff_122640_216000# gnd! 30.9fF
C825 diff_121560_218760# gnd! 70.2fF
C826 diff_95160_187560# gnd! 31.5fF
C827 diff_90600_187200# gnd! 31.8fF
C828 diff_94080_190320# gnd! 70.7fF
C829 diff_81360_173400# gnd! 34.7fF
C830 diff_80400_176040# gnd! 70.9fF
C831 diff_54840_168480# gnd! 1091.2fF
C832 diff_56880_170160# gnd! 189.2fF
C833 diff_42360_157080# gnd! 288.0fF
C834 diff_48720_169080# gnd! 156.1fF
C835 diff_66480_176040# gnd! 1424.5fF
C836 diff_56880_174120# gnd! 190.9fF
C837 diff_54840_175200# gnd! 1090.1fF
C838 diff_43680_161280# gnd! 432.9fF
C839 diff_8880_168480# gnd! 250.8fF
C840 diff_50640_174720# gnd! 247.3fF
C841 diff_48720_174000# gnd! 161.9fF
C842 diff_48720_180120# gnd! 145.6fF
C843 diff_50640_182520# gnd! 241.5fF
C844 diff_81360_183480# gnd! 33.5fF
C845 diff_80400_181920# gnd! 70.7fF
C846 diff_66480_182520# gnd! 1408.6fF
C847 diff_54840_182640# gnd! 1087.9fF
C848 diff_56880_184320# gnd! 201.3fF
C849 diff_88080_190440# gnd! 68.0fF
C850 diff_94080_196200# gnd! 71.5fF
C851 diff_95160_197640# gnd! 31.7fF
C852 diff_88080_196200# gnd! 69.0fF
C853 diff_90600_197760# gnd! 31.4fF
C854 diff_101760_204840# gnd! 69.8fF
C855 diff_108840_211920# gnd! 30.7fF
C856 diff_107880_210360# gnd! 69.6fF
C857 diff_101760_210360# gnd! 70.5fF
C858 diff_104280_212280# gnd! 30.6fF
C859 diff_115560_218880# gnd! 66.4fF
C860 diff_122640_225960# gnd! 30.8fF
C861 diff_121560_224640# gnd! 70.8fF
C862 diff_115560_224520# gnd! 69.1fF
C863 diff_117960_226800# gnd! 33.2fF
C864 diff_129240_233040# gnd! 68.5fF
C865 diff_129240_238680# gnd! 68.8fF
C866 diff_131760_240600# gnd! 31.5fF
C867 diff_143040_247200# gnd! 67.5fF
C868 diff_150120_254280# gnd! 30.7fF
C869 diff_145440_254760# gnd! 33.5fF
C870 diff_143040_252840# gnd! 68.1fF
C871 diff_149040_252840# gnd! 68.5fF
C872 diff_155880_145800# gnd! 458.0fF
C873 diff_153120_145800# gnd! 481.6fF
C874 diff_149520_144360# gnd! 491.7fF
C875 diff_150120_258480# gnd! 30.7fF
C876 diff_145440_258120# gnd! 33.8fF
C877 diff_156720_261360# gnd! 68.4fF
C878 diff_149040_261240# gnd! 68.9fF
C879 diff_136320_244320# gnd! 30.7fF
C880 diff_131760_243960# gnd! 30.8fF
C881 diff_135360_246960# gnd! 68.9fF
C882 diff_122640_230160# gnd! 30.7fF
C883 diff_117960_229800# gnd! 34.3fF
C884 diff_121560_232920# gnd! 70.2fF
C885 diff_108840_216000# gnd! 30.5fF
C886 diff_104280_215640# gnd! 30.7fF
C887 diff_107880_218760# gnd! 71.1fF
C888 diff_95160_201840# gnd! 31.2fF
C889 diff_90600_201480# gnd! 30.9fF
C890 diff_94080_204480# gnd! 69.6fF
C891 diff_81360_187680# gnd! 33.6fF
C892 diff_80400_190320# gnd! 69.1fF
C893 diff_66480_190200# gnd! 1396.0fF
C894 diff_56880_188280# gnd! 203.1fF
C895 diff_44040_187920# gnd! 67.1fF
C896 diff_54840_189360# gnd! 1135.8fF
C897 diff_50640_190200# gnd! 240.4fF
C898 diff_48720_192480# gnd! 146.6fF
C899 diff_6960_191160# gnd! 901.3fF
C900 d3 gnd! 3107.4fF
C901 diff_6840_159480# gnd! 835.6fF
C902 diff_50640_196800# gnd! 237.0fF
C903 diff_66480_196680# gnd! 1379.3fF
C904 diff_81360_197640# gnd! 34.8fF
C905 diff_80400_196200# gnd! 69.6fF
C906 diff_54840_196800# gnd! 1103.8fF
C907 diff_56880_198480# gnd! 191.0fF
C908 diff_88080_204720# gnd! 68.0fF
C909 diff_95160_211920# gnd! 30.8fF
C910 diff_94080_210360# gnd! 72.1fF
C911 diff_88080_210480# gnd! 68.4fF
C912 diff_90480_213840# gnd! 31.8fF
C913 diff_101760_218880# gnd! 70.7fF
C914 diff_108840_225960# gnd! 31.8fF
C915 diff_107880_224520# gnd! 71.3fF
C916 diff_101760_224520# gnd! 72.0fF
C917 diff_104280_226320# gnd! 31.4fF
C918 diff_115560_233040# gnd! 68.1fF
C919 diff_108840_230040# gnd! 31.2fF
C920 diff_104280_229800# gnd! 31.2fF
C921 diff_107880_232800# gnd! 69.5fF
C922 diff_122640_240120# gnd! 31.3fF
C923 diff_121560_238680# gnd! 70.0fF
C924 diff_117960_240600# gnd! 34.0fF
C925 diff_115560_238680# gnd! 67.8fF
C926 diff_129240_247200# gnd! 68.5fF
C927 diff_136320_254280# gnd! 30.7fF
C928 diff_135360_252840# gnd! 68.7fF
C929 diff_129240_252840# gnd! 68.3fF
C930 diff_131760_254760# gnd! 31.2fF
C931 diff_144360_145800# gnd! 495.8fF
C932 diff_143040_261360# gnd! 67.8fF
C933 diff_142200_145800# gnd! 483.6fF
C934 diff_136320_258480# gnd! 30.7fF
C935 diff_131760_258120# gnd! 31.2fF
C936 diff_139320_149640# gnd! 456.6fF
C937 diff_135360_261120# gnd! 68.4fF
C938 diff_135720_144480# gnd! 529.2fF
C939 diff_122640_244320# gnd! 30.7fF
C940 diff_117960_243960# gnd! 33.6fF
C941 diff_121560_247080# gnd! 68.6fF
C942 diff_95160_216000# gnd! 30.9fF
C943 diff_90480_215640# gnd! 32.0fF
C944 diff_81360_201840# gnd! 34.2fF
C945 diff_80400_204480# gnd! 70.1fF
C946 diff_48720_197520# gnd! 155.1fF
C947 diff_42360_185400# gnd! 287.2fF
C948 diff_66480_204480# gnd! 1406.8fF
C949 diff_56880_202560# gnd! 192.8fF
C950 diff_54840_203640# gnd! 1087.3fF
C951 diff_50640_203760# gnd! 241.7fF
C952 diff_33120_151080# gnd! 656.8fF
C953 diff_48720_202920# gnd! 155.7fF
C954 diff_48720_208560# gnd! 143.7fF
C955 diff_50640_210960# gnd! 241.4fF
C956 diff_66480_210960# gnd! 1442.8fF
C957 diff_81360_211920# gnd! 33.5fF
C958 diff_80400_210360# gnd! 70.3fF
C959 diff_81360_216000# gnd! 33.5fF
C960 diff_54840_210960# gnd! 1085.9fF
C961 diff_56880_212760# gnd! 194.9fF
C962 diff_94080_218760# gnd! 71.6fF
C963 diff_88080_218880# gnd! 68.0fF
C964 diff_80400_218760# gnd! 68.8fF
C965 diff_95160_225960# gnd! 31.5fF
C966 diff_94080_224640# gnd! 72.2fF
C967 diff_88080_224520# gnd! 69.0fF
C968 diff_90480_226440# gnd! 33.8fF
C969 diff_101760_233040# gnd! 68.7fF
C970 diff_101760_238680# gnd! 68.3fF
C971 diff_108840_240120# gnd! 31.8fF
C972 diff_107880_238680# gnd! 69.2fF
C973 diff_104280_240480# gnd! 31.7fF
C974 diff_115560_247200# gnd! 67.0fF
C975 diff_115560_252840# gnd! 67.2fF
C976 diff_117960_254760# gnd! 33.9fF
C977 diff_122640_254280# gnd! 31.2fF
C978 diff_121560_252840# gnd! 69.0fF
C979 diff_128400_145800# gnd! 458.1fF
C980 diff_125640_145800# gnd! 495.8fF
C981 diff_122040_144240# gnd! 491.4fF
C982 diff_117960_258120# gnd! 33.9fF
C983 diff_122640_258480# gnd! 31.2fF
C984 diff_130680_145800# gnd! 491.7fF
C985 diff_129240_261360# gnd! 66.8fF
C986 diff_121560_261120# gnd! 69.5fF
C987 diff_116880_145800# gnd! 537.9fF
C988 diff_108840_244320# gnd! 30.7fF
C989 diff_104280_243960# gnd! 30.8fF
C990 diff_107880_246960# gnd! 69.1fF
C991 diff_95160_230160# gnd! 30.8fF
C992 diff_90480_229800# gnd! 34.2fF
C993 diff_94080_232920# gnd! 70.4fF
C994 diff_66480_218640# gnd! 1420.9fF
C995 diff_17040_204360# gnd! 248.6fF
C996 diff_16320_201240# gnd! 245.7fF
C997 diff_56880_216720# gnd! 201.6fF
C998 diff_54840_217800# gnd! 1086.9fF
C999 diff_44040_216360# gnd! 65.2fF
C1000 diff_50640_218640# gnd! 241.4fF
C1001 diff_48720_220920# gnd! 143.1fF
C1002 diff_50640_225120# gnd! 237.4fF
C1003 diff_66480_225120# gnd! 1399.7fF
C1004 diff_81360_225960# gnd! 31.6fF
C1005 diff_80400_224520# gnd! 69.4fF
C1006 diff_81360_230160# gnd! 30.5fF
C1007 diff_88080_233040# gnd! 68.3fF
C1008 diff_80400_232800# gnd! 69.3fF
C1009 diff_95040_240840# gnd! 33.7fF
C1010 diff_94080_238680# gnd! 70.3fF
C1011 diff_88080_238680# gnd! 68.5fF
C1012 diff_90480_240600# gnd! 34.6fF
C1013 diff_101760_247200# gnd! 68.6fF
C1014 diff_108840_254280# gnd! 31.0fF
C1015 diff_107760_253200# gnd! 69.3fF
C1016 diff_101760_252840# gnd! 68.8fF
C1017 diff_104280_254640# gnd! 31.2fF
C1018 diff_108840_258480# gnd! 31.0fF
C1019 diff_114720_145800# gnd! 472.9fF
C1020 diff_111840_149760# gnd! 459.0fF
C1021 diff_108240_144360# gnd! 555.8fF
C1022 diff_115560_261360# gnd! 67.2fF
C1023 diff_107880_261120# gnd! 68.6fF
C1024 diff_104280_258120# gnd! 31.2fF
C1025 diff_95040_244320# gnd! 33.4fF
C1026 diff_90480_243960# gnd! 33.8fF
C1027 diff_94080_247080# gnd! 67.6fF
C1028 diff_54840_225240# gnd! 1082.8fF
C1029 diff_56760_227400# gnd! 192.8fF
C1030 diff_48720_225840# gnd! 155.4fF
C1031 diff_42360_213840# gnd! 281.6fF
C1032 diff_66480_232800# gnd! 1432.4fF
C1033 diff_56760_230880# gnd! 191.4fF
C1034 diff_54840_231960# gnd! 1080.7fF
C1035 diff_50640_232080# gnd! 240.9fF
C1036 diff_16200_228600# gnd! 114.9fF
C1037 diff_32760_140400# gnd! 738.4fF
C1038 diff_48720_231240# gnd! 158.2fF
C1039 diff_48720_236880# gnd! 141.3fF
C1040 diff_23160_135720# gnd! 3699.5fF
C1041 diff_50640_239280# gnd! 242.8fF
C1042 diff_66480_239280# gnd! 1400.2fF
C1043 diff_81360_240120# gnd! 32.0fF
C1044 diff_80400_238680# gnd! 69.8fF
C1045 diff_88080_247200# gnd! 67.7fF
C1046 diff_81360_244320# gnd! 30.4fF
C1047 diff_54840_239280# gnd! 1082.4fF
C1048 diff_56760_241080# gnd! 198.5fF
C1049 diff_80400_246960# gnd! 67.6fF
C1050 diff_95040_256560# gnd! 32.0fF
C1051 diff_94080_252840# gnd! 71.3fF
C1052 diff_90480_254760# gnd! 34.5fF
C1053 diff_88080_252840# gnd! 67.2fF
C1054 diff_100920_145800# gnd! 465.5fF
C1055 diff_98160_145800# gnd! 486.7fF
C1056 diff_94560_144240# gnd! 492.4fF
C1057 diff_95160_258480# gnd! 31.2fF
C1058 diff_90480_258120# gnd! 34.2fF
C1059 diff_103200_145800# gnd! 491.0fF
C1060 diff_101760_261360# gnd! 67.8fF
C1061 diff_94080_261120# gnd! 70.2fF
C1062 diff_89400_145800# gnd! 526.1fF
C1063 diff_16200_238800# gnd! 112.5fF
C1064 diff_66360_247080# gnd! 1448.3fF
C1065 diff_56760_245040# gnd! 198.5fF
C1066 diff_54840_246000# gnd! 1079.1fF
C1067 diff_44040_244680# gnd! 70.2fF
C1068 diff_50640_246720# gnd! 244.9fF
C1069 diff_48720_249120# gnd! 142.5fF
C1070 diff_8760_249240# gnd! 246.6fF
C1071 diff_50640_253320# gnd! 248.0fF
C1072 diff_66480_253440# gnd! 1381.8fF
C1073 diff_81360_254280# gnd! 31.5fF
C1074 diff_80400_252840# gnd! 68.9fF
C1075 diff_81360_258480# gnd! 31.1fF
C1076 diff_87240_145800# gnd! 459.6fF
C1077 diff_84360_149760# gnd! 493.2fF
C1078 diff_80760_144360# gnd! 515.3fF
C1079 diff_88080_261360# gnd! 68.0fF
C1080 diff_80400_261120# gnd! 68.4fF
C1081 diff_54840_253440# gnd! 1123.8fF
C1082 diff_56760_255360# gnd! 197.2fF
C1083 diff_48720_255480# gnd! 158.5fF
C1084 diff_23040_212640# gnd! 3323.5fF
C1085 diff_42360_242040# gnd! 281.0fF
C1086 diff_66360_261120# gnd! 1408.6fF
C1087 diff_56760_259080# gnd! 195.2fF
C1088 diff_42600_159120# gnd! 1371.5fF
C1089 diff_54840_260160# gnd! 1051.2fF
C1090 diff_50640_260400# gnd! 250.9fF
C1091 diff_48720_260280# gnd! 143.8fF
C1092 diff_52320_146760# gnd! 737.8fF
C1093 diff_32640_245760# gnd! 843.4fF
C1094 diff_232560_264480# gnd! 40.3fF
C1095 diff_242400_271320# gnd! 71.3fF
C1096 diff_234600_265200# gnd! 299.9fF
C1097 diff_245400_273720# gnd! 80.5fF
C1098 clk2 gnd! 3716.3fF
C1099 diff_210480_277440# gnd! 36.7fF
C1100 diff_6960_253440# gnd! 903.5fF
C1101 d2 gnd! 3131.8fF
C1102 diff_6840_236160# gnd! 833.1fF
C1103 o1 gnd! 1073.5fF
C1104 diff_237360_275280# gnd! 235.8fF
C1105 diff_241560_285240# gnd! 405.3fF
C1106 diff_207480_277200# gnd! 1558.0fF
C1107 diff_22200_108240# gnd! 1302.3fF
C1108 diff_34920_109680# gnd! 2998.9fF
C1109 diff_205080_288960# gnd! 66.3fF
C1110 diff_201600_290400# gnd! 70.4fF
C1111 diff_192360_286440# gnd! 218.2fF
C1112 diff_207720_290040# gnd! 780.4fF
C1113 o0 gnd! 1015.4fF
C1114 diff_135840_285600# gnd! 113.6fF
C1115 diff_126120_285720# gnd! 116.5fF
C1116 diff_100920_281280# gnd! 245.1fF
C1117 diff_94320_284400# gnd! 258.0fF
C1118 diff_142920_287880# gnd! 225.6fF
C1119 diff_126240_288840# gnd! 909.5fF
C1120 diff_133080_289920# gnd! 817.1fF
C1121 diff_25200_276600# gnd! 3238.3fF
C1122 diff_38640_285720# gnd! 116.3fF
C1123 Vdd gnd! 40389.6fF
C1124 diff_13200_279960# gnd! 1886.4fF
C1125 diff_16560_282240# gnd! 244.5fF
C1126 diff_9720_284520# gnd! 261.9fF
C1127 diff_28920_285720# gnd! 119.2fF
C1128 diff_45720_287880# gnd! 244.2fF
C1129 diff_8760_228840# gnd! 2092.1fF
C1130 diff_28920_288480# gnd! 907.9fF
C1131 diff_35880_289800# gnd! 830.3fF
C1132 diff_191640_286080# gnd! 411.9fF
C1133 d0 gnd! 2932.6fF
C1134 d1 gnd! 2915.7fF
C1135 diff_201720_295920# gnd! 288.6fF
