* SPICE3 file created from 4002.ext - technology: nmos

.option scale=0.001u

M1000 diff_306070_3053080# diff_379730_3067050# GND GND efet w=81915 l=7620
+ ad=-9.62716e+08 pd=619760 as=1.71928e+09 ps=7.61035e+07 
M1001 d1 GND GND GND efet w=111760 l=8890
+ ad=-1.40068e+09 pd=3.21056e+06 as=0 ps=0 
M1002 GND diff_92710_2421890# diff_306070_3053080# GND efet w=227965 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1003 GND d1 diff_102870_3011170# GND efet w=59055 l=6985
+ ad=0 pd=0 as=1.47419e+09 ps=307340 
M1004 GND diff_92710_2421890# diff_379730_3067050# GND efet w=236220 l=6985
+ ad=0 pd=0 as=4.21208e+07 ps=805180 
M1005 diff_379730_3067050# diff_483870_3046730# GND GND efet w=224155 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1006 diff_306070_3053080# diff_306070_3023870# diff_306070_3053080# GND efet w=42545 l=13970
+ ad=0 pd=0 as=0 ps=0 
M1007 GND diff_102870_3011170# diff_175260_2987040# GND efet w=23495 l=8255
+ ad=0 pd=0 as=1.61129e+09 ps=289560 
M1008 diff_102870_3011170# diff_102870_3011170# diff_102870_3011170# GND efet w=2540 l=5080
+ ad=0 pd=0 as=0 ps=0 
M1009 diff_102870_3011170# diff_102870_3011170# diff_102870_3011170# GND efet w=1905 l=1905
+ ad=0 pd=0 as=0 ps=0 
M1010 diff_175260_2987040# diff_175260_2987040# diff_175260_2987040# GND efet w=3810 l=3810
+ ad=0 pd=0 as=0 ps=0 
M1011 diff_175260_2987040# diff_175260_2987040# diff_175260_2987040# GND efet w=1270 l=5080
+ ad=0 pd=0 as=0 ps=0 
M1012 diff_102870_3011170# Vdd Vdd GND efet w=10160 l=37465
+ ad=0 pd=0 as=3.03689e+08 ps=3.69799e+07 
M1013 GND diff_139700_2962910# diff_102870_3011170# GND efet w=36830 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1014 diff_175260_2987040# diff_139700_2962910# GND GND efet w=38735 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1015 GND diff_306070_3053080# d1 GND efet w=1189355 l=4445
+ ad=0 pd=0 as=0 ps=0 
M1016 diff_379730_3067050# diff_408940_3023870# diff_379730_3067050# GND efet w=45085 l=13970
+ ad=0 pd=0 as=0 ps=0 
M1017 diff_306070_3053080# diff_306070_3023870# Vdd GND efet w=12065 l=9525
+ ad=0 pd=0 as=0 ps=0 
M1018 diff_306070_3023870# diff_306070_3023870# diff_306070_3023870# GND efet w=3175 l=4445
+ ad=2.46774e+08 pd=81280 as=0 ps=0 
M1019 diff_306070_3023870# diff_306070_3023870# diff_306070_3023870# GND efet w=1905 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1020 diff_379730_3067050# diff_408940_3023870# Vdd GND efet w=12065 l=9525
+ ad=0 pd=0 as=0 ps=0 
M1021 diff_408940_3023870# diff_408940_3023870# diff_408940_3023870# GND efet w=3175 l=4445
+ ad=2.37096e+08 pd=76200 as=0 ps=0 
M1022 diff_408940_3023870# diff_408940_3023870# diff_408940_3023870# GND efet w=1905 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1023 diff_306070_3023870# Vdd Vdd GND efet w=10160 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1024 Vdd Vdd Vdd GND efet w=2540 l=5080
+ ad=0 pd=0 as=0 ps=0 
M1025 Vdd Vdd Vdd GND efet w=1270 l=1270
+ ad=0 pd=0 as=0 ps=0 
M1026 Vdd Vdd diff_175260_2987040# GND efet w=8890 l=40005
+ ad=0 pd=0 as=0 ps=0 
M1027 diff_266700_2927350# diff_175260_2987040# Vdd GND efet w=40640 l=10160
+ ad=1.70217e+09 pd=2.97688e+06 as=0 ps=0 
M1028 GND diff_102870_3011170# diff_266700_2927350# GND efet w=40640 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1029 d0 GND GND GND efet w=114300 l=8890
+ ad=-1.94423e+09 pd=3.22834e+06 as=0 ps=0 
M1030 GND diff_92710_2421890# diff_1336040_3056890# GND efet w=223520 l=7620
+ ad=0 pd=0 as=-9.72393e+08 ps=612140 
M1031 GND d0 diff_998220_3009900# GND efet w=58420 l=7620
+ ad=0 pd=0 as=1.43064e+09 ps=302260 
M1032 diff_1336040_3056890# diff_1408430_3068320# GND GND efet w=80010 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1033 GND diff_92710_2421890# diff_1408430_3068320# GND efet w=230505 l=8255
+ ad=0 pd=0 as=-4.6533e+06 ps=759460 
M1034 diff_1408430_3068320# diff_1512570_3046730# GND GND efet w=224790 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1035 GND diff_998220_3009900# diff_1068070_2976880# GND efet w=22860 l=7620
+ ad=0 pd=0 as=1.63548e+09 ps=304800 
M1036 diff_998220_3009900# diff_998220_3009900# diff_998220_3009900# GND efet w=2540 l=6350
+ ad=0 pd=0 as=0 ps=0 
M1037 diff_1068070_2976880# diff_1068070_2976880# diff_1068070_2976880# GND efet w=6350 l=5080
+ ad=0 pd=0 as=0 ps=0 
M1038 d1 diff_379730_3067050# Vdd GND efet w=641350 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1039 diff_483870_3046730# diff_483870_3046730# diff_483870_3046730# GND efet w=2540 l=10160
+ ad=1.11613e+09 pd=236220 as=0 ps=0 
M1040 diff_408940_3023870# Vdd Vdd GND efet w=8890 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1041 diff_483870_3046730# diff_483870_3046730# diff_483870_3046730# GND efet w=3175 l=5080
+ ad=0 pd=0 as=0 ps=0 
M1042 diff_1068070_2976880# diff_1068070_2976880# diff_1068070_2976880# GND efet w=1905 l=5715
+ ad=0 pd=0 as=0 ps=0 
M1043 diff_998220_3009900# Vdd Vdd GND efet w=9525 l=37465
+ ad=0 pd=0 as=0 ps=0 
M1044 GND diff_139700_2962910# diff_998220_3009900# GND efet w=36830 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1045 diff_1068070_2976880# diff_139700_2962910# GND GND efet w=36830 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1046 diff_1336040_3056890# diff_1334770_3023870# diff_1336040_3056890# GND efet w=38735 l=33655
+ ad=0 pd=0 as=0 ps=0 
M1047 GND diff_1336040_3056890# d0 GND efet w=1180465 l=4445
+ ad=0 pd=0 as=0 ps=0 
M1048 diff_1408430_3068320# diff_1437640_3022600# diff_1408430_3068320# GND efet w=36195 l=35560
+ ad=0 pd=0 as=0 ps=0 
M1049 o0 diff_2028190_3027680# GND GND efet w=209550 l=7620
+ ad=-1.4275e+06 pd=731520 as=0 ps=0 
M1050 diff_2028190_3027680# diff_2134870_3131820# GND GND efet w=116840 l=7620
+ ad=1.53548e+09 pd=299720 as=0 ps=0 
M1051 diff_2035810_3031490# diff_2028190_3027680# GND GND efet w=50800 l=7620
+ ad=1.05e+09 pd=182880 as=0 ps=0 
M1052 diff_2133600_3073400# diff_2028190_3027680# GND GND efet w=25400 l=7620
+ ad=6.35483e+08 pd=144780 as=0 ps=0 
M1053 diff_2134870_3131820# diff_2170430_3058160# diff_2133600_3073400# GND efet w=13970 l=7620
+ ad=1.64677e+09 pd=337820 as=0 ps=0 
M1054 GND diff_2198370_3069590# diff_2134870_3131820# GND efet w=26670 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1055 diff_2035810_3031490# diff_2035810_3031490# diff_2035810_3031490# GND efet w=3810 l=5080
+ ad=0 pd=0 as=0 ps=0 
M1056 diff_2035810_3031490# diff_2035810_3031490# diff_2035810_3031490# GND efet w=1270 l=2540
+ ad=0 pd=0 as=0 ps=0 
M1057 o0 diff_2035810_3031490# Vdd GND efet w=224155 l=6985
+ ad=0 pd=0 as=0 ps=0 
M1058 d0 diff_1408430_3068320# Vdd GND efet w=644525 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1059 diff_1336040_3056890# diff_1334770_3023870# Vdd GND efet w=10795 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1060 diff_1334770_3023870# diff_1334770_3023870# diff_1334770_3023870# GND efet w=2540 l=4445
+ ad=2.35483e+08 pd=73660 as=0 ps=0 
M1061 diff_1334770_3023870# diff_1334770_3023870# diff_1334770_3023870# GND efet w=1270 l=6350
+ ad=0 pd=0 as=0 ps=0 
M1062 diff_1437640_3022600# diff_1437640_3022600# diff_1437640_3022600# GND efet w=2540 l=4445
+ ad=2.20967e+08 pd=71120 as=0 ps=0 
M1063 diff_1437640_3022600# diff_1437640_3022600# diff_1437640_3022600# GND efet w=1905 l=5715
+ ad=0 pd=0 as=0 ps=0 
M1064 Vdd Vdd Vdd GND efet w=2540 l=6350
+ ad=0 pd=0 as=0 ps=0 
M1065 diff_483870_3046730# diff_234950_1145540# diff_266700_2927350# GND efet w=31115 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1066 Vdd Vdd diff_1068070_2976880# GND efet w=8890 l=39370
+ ad=0 pd=0 as=0 ps=0 
M1067 diff_369570_1160780# diff_1068070_2976880# Vdd GND efet w=39370 l=7620
+ ad=3.81201e+08 pd=2.62636e+06 as=0 ps=0 
M1068 GND diff_998220_3009900# diff_369570_1160780# GND efet w=41275 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1069 diff_1334770_3023870# Vdd Vdd GND efet w=10795 l=9525
+ ad=0 pd=0 as=0 ps=0 
M1070 diff_1408430_3068320# diff_1437640_3022600# Vdd GND efet w=10160 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1071 Vdd Vdd diff_1437640_3022600# GND efet w=8255 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1072 Vdd Vdd Vdd GND efet w=1270 l=1270
+ ad=0 pd=0 as=0 ps=0 
M1073 diff_2035810_3031490# Vdd Vdd GND efet w=10160 l=20320
+ ad=0 pd=0 as=0 ps=0 
M1074 diff_2133600_3073400# Vdd Vdd GND efet w=7620 l=31750
+ ad=0 pd=0 as=0 ps=0 
M1075 GND diff_2195830_2933700# diff_2170430_3058160# GND efet w=13970 l=7620
+ ad=0 pd=0 as=3.32257e+08 ps=78740 
M1076 diff_2170430_3058160# Vdd Vdd GND efet w=8255 l=60325
+ ad=0 pd=0 as=0 ps=0 
M1077 Vdd Vdd Vdd GND efet w=5080 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1078 Vdd Vdd Vdd GND efet w=5715 l=4445
+ ad=0 pd=0 as=0 ps=0 
M1079 diff_2028190_3027680# Vdd Vdd GND efet w=12065 l=19685
+ ad=0 pd=0 as=0 ps=0 
M1080 GND diff_2556510_3018790# diff_2512060_2913380# GND efet w=52070 l=7620
+ ad=0 pd=0 as=1.28871e+09 ps=198120 
M1081 GND diff_2556510_3018790# o1 GND efet w=214630 l=6350
+ ad=0 pd=0 as=3.24378e+08 ps=749300 
M1082 diff_2134870_3131820# diff_2195830_2933700# diff_2227580_2936240# GND efet w=20320 l=6985
+ ad=0 pd=0 as=3.2258e+08 ps=83820 
M1083 Vdd diff_72390_2499360# d2 GND efet w=659765 l=6985
+ ad=0 pd=0 as=-2.60363e+08 ps=3.24866e+06 
M1084 GND diff_73660_2682240# d2 GND efet w=1210945 l=4445
+ ad=0 pd=0 as=0 ps=0 
M1085 diff_1512570_3046730# diff_234950_1145540# diff_369570_1160780# GND efet w=27940 l=7620
+ ad=9.19353e+08 pd=180340 as=0 ps=0 
M1086 diff_2227580_2936240# clk2 diff_369570_1160780# GND efet w=19050 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1087 diff_2512060_2913380# Vdd Vdd GND efet w=11430 l=20320
+ ad=0 pd=0 as=0 ps=0 
M1088 diff_2512060_2913380# diff_2512060_2913380# diff_2512060_2913380# GND efet w=4445 l=4445
+ ad=0 pd=0 as=0 ps=0 
M1089 o1 diff_2512060_2913380# Vdd GND efet w=221615 l=6985
+ ad=0 pd=0 as=0 ps=0 
M1090 GND diff_2556510_3018790# diff_2597150_2896870# GND efet w=27940 l=8890
+ ad=0 pd=0 as=7.38708e+08 ps=154940 
M1091 diff_2597150_2896870# Vdd Vdd GND efet w=11430 l=30480
+ ad=0 pd=0 as=0 ps=0 
M1092 Vdd Vdd Vdd GND efet w=3810 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1093 Vdd Vdd Vdd GND efet w=3810 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1094 GND diff_2482850_2806700# diff_2556510_3018790# GND efet w=118110 l=5715
+ ad=0 pd=0 as=1.58064e+09 ps=292100 
M1095 diff_2597150_2896870# diff_2565400_2871470# diff_2482850_2806700# GND efet w=15240 l=8890
+ ad=0 pd=0 as=1.83064e+09 ps=345440 
M1096 diff_2565400_2871470# Vdd Vdd GND efet w=8890 l=60960
+ ad=3.87096e+08 pd=83820 as=0 ps=0 
M1097 diff_2565400_2871470# diff_2195830_2933700# GND GND efet w=15875 l=6985
+ ad=0 pd=0 as=0 ps=0 
M1098 diff_2482850_2806700# diff_2198370_3069590# GND GND efet w=26670 l=6985
+ ad=0 pd=0 as=0 ps=0 
M1099 Vdd Vdd Vdd GND efet w=3175 l=4445
+ ad=0 pd=0 as=0 ps=0 
M1100 Vdd Vdd Vdd GND efet w=2540 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1101 diff_515620_2754630# diff_345440_2600960# diff_369570_1160780# GND efet w=40640 l=7620
+ ad=1.10806e+09 pd=241300 as=0 ps=0 
M1102 diff_515620_2754630# diff_553720_1553210# diff_535940_2755900# GND efet w=40640 l=7620
+ ad=0 pd=0 as=1.94677e+09 ps=360680 
M1103 diff_580390_2753360# diff_450850_1684020# diff_515620_2754630# GND efet w=48895 l=8255
+ ad=-7.40136e+08 pd=914400 as=0 ps=0 
M1104 diff_2461260_2799080# clk2 diff_266700_2927350# GND efet w=21590 l=7620
+ ad=3.59677e+08 pd=86360 as=0 ps=0 
M1105 diff_2482850_2806700# diff_2195830_2933700# diff_2461260_2799080# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1106 diff_600710_2741930# Vdd Vdd GND efet w=8890 l=31750
+ ad=1.02903e+09 pd=238760 as=0 ps=0 
M1107 Vdd diff_702310_2763520# diff_535940_2755900# GND efet w=16510 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1108 diff_600710_2741930# diff_448310_2561590# diff_580390_2753360# GND efet w=34290 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1109 diff_515620_2703830# diff_345440_2600960# diff_266700_2927350# GND efet w=40640 l=7620
+ ad=1.10806e+09 pd=241300 as=0 ps=0 
M1110 diff_600710_2702560# diff_448310_2561590# diff_580390_2682240# GND efet w=33655 l=8255
+ ad=1.03226e+09 pd=231140 as=-6.99813e+08 ps=937260 
M1111 diff_535940_2755900# diff_600710_2741930# GND GND efet w=58420 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1112 diff_600710_2741930# diff_702310_2763520# GND GND efet w=28575 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1113 GND diff_600710_2702560# diff_535940_2680970# GND efet w=57150 l=8890
+ ad=0 pd=0 as=1.94354e+09 ps=353060 
M1114 diff_861060_2735580# diff_850900_2763520# GND GND efet w=24130 l=7620
+ ad=2.69354e+08 pd=76200 as=0 ps=0 
M1115 diff_580390_2753360# diff_892810_1584960# diff_850900_2763520# GND efet w=10160 l=7620
+ ad=0 pd=0 as=3.01612e+08 ps=78740 
M1116 diff_932180_2766060# diff_923290_1543050# diff_580390_2753360# GND efet w=10160 l=7620
+ ad=2.93548e+08 pd=78740 as=0 ps=0 
M1117 diff_702310_2763520# diff_854710_1527810# diff_861060_2735580# GND efet w=22860 l=8890
+ ad=-1.34156e+09 pd=1.63068e+06 as=0 ps=0 
M1118 diff_703580_2682240# diff_854710_1527810# diff_861060_2691130# GND efet w=23495 l=10160
+ ad=-1.66414e+09 pd=1.6383e+06 as=2.70967e+08 ps=78740 
M1119 diff_72390_2499360# diff_92710_2637790# GND GND efet w=227965 l=6985
+ ad=1.1954e+08 pd=833120 as=0 ps=0 
M1120 diff_92710_2637790# diff_92710_2637790# diff_92710_2637790# GND efet w=1905 l=6985
+ ad=1.29838e+09 pd=231140 as=0 ps=0 
M1121 diff_92710_2637790# diff_92710_2637790# diff_92710_2637790# GND efet w=3175 l=4445
+ ad=0 pd=0 as=0 ps=0 
M1122 diff_243840_2250440# diff_234950_1145540# diff_92710_2637790# GND efet w=29210 l=7620
+ ad=3.68297e+08 pd=2.6289e+06 as=0 ps=0 
M1123 diff_515620_2636520# diff_345440_2600960# diff_243840_2250440# GND efet w=40640 l=7620
+ ad=1.0758e+09 pd=241300 as=0 ps=0 
M1124 diff_515620_2703830# diff_553720_1553210# diff_535940_2680970# GND efet w=40640 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1125 diff_580390_2682240# diff_450850_1684020# diff_515620_2703830# GND efet w=47625 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1126 GND diff_703580_2682240# diff_600710_2702560# GND efet w=27940 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1127 GND diff_345440_2600960# diff_466090_2589530# GND efet w=55245 l=8255
+ ad=0 pd=0 as=6.43547e+08 ps=134620 
M1128 diff_515620_2636520# diff_553720_1553210# diff_535940_2611120# GND efet w=39370 l=7620
+ ad=0 pd=0 as=1.91935e+09 ps=342900 
M1129 diff_580390_2603500# diff_450850_1684020# diff_515620_2636520# GND efet w=47625 l=8255
+ ad=-8.04652e+08 pd=909320 as=0 ps=0 
M1130 Vdd diff_703580_2682240# diff_535940_2680970# GND efet w=15875 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1131 diff_861060_2691130# diff_850900_2675890# GND GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1132 diff_600710_2702560# Vdd Vdd GND efet w=7620 l=29210
+ ad=0 pd=0 as=0 ps=0 
M1133 Vdd Vdd Vdd GND efet w=6350 l=3810
+ ad=0 pd=0 as=0 ps=0 
M1134 Vdd Vdd Vdd GND efet w=4445 l=12065
+ ad=0 pd=0 as=0 ps=0 
M1135 diff_600710_2593340# Vdd Vdd GND efet w=7620 l=29210
+ ad=1.08548e+09 pd=246380 as=0 ps=0 
M1136 diff_600710_2593340# diff_448310_2561590# diff_580390_2603500# GND efet w=34290 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1137 diff_466090_2589530# diff_450850_1684020# diff_448310_2561590# GND efet w=51435 l=8255
+ ad=0 pd=0 as=1.10484e+09 ps=215900 
M1138 diff_72390_2499360# diff_92710_2421890# GND GND efet w=227965 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1139 Vdd diff_171450_2527300# diff_72390_2499360# GND efet w=11430 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1140 Vdd Vdd diff_448310_2561590# GND efet w=12700 l=41275
+ ad=0 pd=0 as=0 ps=0 
M1141 diff_72390_2499360# diff_171450_2527300# diff_72390_2499360# GND efet w=51435 l=19050
+ ad=0 pd=0 as=0 ps=0 
M1142 diff_171450_2527300# diff_171450_2527300# diff_171450_2527300# GND efet w=3175 l=8255
+ ad=2.66128e+08 pd=81280 as=0 ps=0 
M1143 Vdd Vdd diff_171450_2527300# GND efet w=10160 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1144 diff_171450_2527300# diff_171450_2527300# diff_171450_2527300# GND efet w=1905 l=3810
+ ad=0 pd=0 as=0 ps=0 
M1145 Vdd Vdd Vdd GND efet w=2540 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1146 Vdd Vdd Vdd GND efet w=1905 l=3810
+ ad=0 pd=0 as=0 ps=0 
M1147 Vdd diff_702310_2614930# diff_535940_2611120# GND efet w=13970 l=6985
+ ad=0 pd=0 as=0 ps=0 
M1148 diff_535940_2611120# diff_600710_2593340# GND GND efet w=55245 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1149 diff_1007110_2735580# diff_995680_2763520# GND GND efet w=24130 l=10160
+ ad=2.66128e+08 pd=78740 as=0 ps=0 
M1150 diff_957580_2731770# diff_946150_1543050# diff_702310_2763520# GND efet w=22860 l=7620
+ ad=2.96774e+08 pd=81280 as=0 ps=0 
M1151 GND diff_932180_2766060# diff_957580_2731770# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1152 diff_580390_2753360# diff_1038860_1543050# diff_995680_2763520# GND efet w=10795 l=7620
+ ad=0 pd=0 as=2.99999e+08 ps=78740 
M1153 diff_1076960_2766060# diff_1068070_1543050# diff_580390_2753360# GND efet w=10160 l=7620
+ ad=2.90322e+08 pd=81280 as=0 ps=0 
M1154 diff_702310_2763520# diff_1000760_1526540# diff_1007110_2735580# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1155 diff_957580_2696210# diff_946150_1543050# diff_703580_2682240# GND efet w=22860 l=7620
+ ad=2.99999e+08 pd=81280 as=0 ps=0 
M1156 diff_703580_2682240# diff_1000760_1526540# diff_1005840_2715260# GND efet w=22860 l=9525
+ ad=0 pd=0 as=2.7258e+08 ps=83820 
M1157 GND diff_932180_2675890# diff_957580_2696210# GND efet w=24765 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1158 diff_580390_2682240# diff_892810_1584960# diff_850900_2675890# GND efet w=8890 l=7620
+ ad=0 pd=0 as=3.01612e+08 ps=81280 
M1159 diff_932180_2675890# diff_923290_1543050# diff_580390_2682240# GND efet w=8890 l=7620
+ ad=2.74193e+08 pd=78740 as=0 ps=0 
M1160 diff_600710_2593340# diff_702310_2614930# GND GND efet w=27940 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1161 diff_600710_2551430# diff_448310_2561590# diff_580390_2532380# GND efet w=34290 l=8255
+ ad=1.08387e+09 pd=246380 as=-7.64329e+08 ps=916940 
M1162 diff_861060_2585720# diff_850900_2613660# GND GND efet w=24130 l=7620
+ ad=2.59677e+08 pd=76200 as=0 ps=0 
M1163 diff_580390_2603500# diff_892810_1584960# diff_850900_2613660# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.8387e+08 ps=78740 
M1164 diff_932180_2616200# diff_923290_1543050# diff_580390_2603500# GND efet w=8890 l=7620
+ ad=2.80645e+08 pd=78740 as=0 ps=0 
M1165 diff_702310_2614930# diff_854710_1527810# diff_861060_2585720# GND efet w=22860 l=8890
+ ad=-1.31898e+09 pd=1.63322e+06 as=0 ps=0 
M1166 diff_703580_2532380# diff_854710_1527810# diff_861060_2541270# GND efet w=23495 l=8255
+ ad=-1.51898e+09 pd=1.64338e+06 as=2.7258e+08 ps=81280 
M1167 GND diff_600710_2551430# diff_535940_2532380# GND efet w=53340 l=7620
+ ad=0 pd=0 as=1.88871e+09 ps=345440 
M1168 GND diff_703580_2532380# diff_600710_2551430# GND efet w=27940 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1169 diff_73660_2682240# diff_72390_2499360# GND GND efet w=83820 l=6350
+ ad=-7.51426e+08 pd=645160 as=0 ps=0 
M1170 diff_515620_2506980# diff_345440_2600960# diff_245110_1436370# GND efet w=40640 l=7620
+ ad=1.08387e+09 pd=241300 as=1.44894e+09 ps=2.87528e+06 
M1171 diff_515620_2506980# diff_553720_1553210# diff_535940_2532380# GND efet w=40005 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1172 diff_580390_2532380# diff_450850_1684020# diff_515620_2506980# GND efet w=48260 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1173 diff_535940_2532380# diff_703580_2532380# Vdd GND efet w=14605 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1174 diff_861060_2541270# diff_850900_2526030# GND GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1175 diff_73660_2682240# diff_92710_2421890# GND GND efet w=228600 l=9525
+ ad=0 pd=0 as=0 ps=0 
M1176 Vdd diff_171450_2419350# diff_73660_2682240# GND efet w=12065 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1177 diff_73660_2682240# diff_171450_2419350# diff_73660_2682240# GND efet w=42545 l=17780
+ ad=0 pd=0 as=0 ps=0 
M1178 diff_171450_2419350# diff_171450_2419350# diff_171450_2419350# GND efet w=2540 l=7620
+ ad=2.51612e+08 pd=81280 as=0 ps=0 
M1179 Vdd Vdd diff_171450_2419350# GND efet w=8890 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1180 diff_515620_2447290# diff_346710_1485900# diff_369570_1160780# GND efet w=40640 l=7620
+ ad=1.23709e+09 pd=266700 as=0 ps=0 
M1181 diff_515620_2447290# diff_553720_1553210# diff_535940_2456180# GND efet w=41910 l=7620
+ ad=0 pd=0 as=1.87096e+09 ps=355600 
M1182 diff_600710_2551430# Vdd Vdd GND efet w=7620 l=29210
+ ad=0 pd=0 as=0 ps=0 
M1183 Vdd Vdd Vdd GND efet w=3810 l=11430
+ ad=0 pd=0 as=0 ps=0 
M1184 Vdd Vdd Vdd GND efet w=6350 l=3810
+ ad=0 pd=0 as=0 ps=0 
M1185 diff_580390_2454910# diff_450850_1684020# diff_515620_2447290# GND efet w=47625 l=8255
+ ad=-8.07878e+08 pd=916940 as=0 ps=0 
M1186 diff_600710_2443480# Vdd Vdd GND efet w=7620 l=30480
+ ad=9.99998e+08 pd=231140 as=0 ps=0 
M1187 Vdd diff_703580_2463800# diff_535940_2456180# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1188 diff_600710_2443480# diff_448310_2263140# diff_580390_2454910# GND efet w=34290 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1189 diff_171450_2419350# diff_171450_2419350# diff_171450_2419350# GND efet w=3175 l=3810
+ ad=0 pd=0 as=0 ps=0 
M1190 diff_515620_2390140# diff_346710_1485900# diff_266700_2927350# GND efet w=39370 l=7620
+ ad=1.07097e+09 pd=243840 as=0 ps=0 
M1191 diff_600710_2406650# diff_448310_2263140# diff_580390_2383790# GND efet w=33655 l=8255
+ ad=9.98385e+08 pd=228600 as=-8.15942e+08 ps=909320 
M1192 diff_535940_2456180# diff_600710_2443480# GND GND efet w=57785 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1193 diff_1005840_2715260# diff_995680_2675890# GND GND efet w=24765 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1194 diff_957580_2581910# diff_946150_1543050# diff_702310_2614930# GND efet w=22860 l=7620
+ ad=2.95161e+08 pd=78740 as=0 ps=0 
M1195 GND diff_932180_2616200# diff_957580_2581910# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1196 diff_1005840_2585720# diff_995680_2614930# GND GND efet w=24765 l=8255
+ ad=2.90322e+08 pd=78740 as=0 ps=0 
M1197 diff_1103630_2731770# diff_1092200_1543050# diff_702310_2763520# GND efet w=22860 l=7620
+ ad=2.67741e+08 pd=78740 as=0 ps=0 
M1198 GND diff_1076960_2766060# diff_1103630_2731770# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1199 diff_1151890_2735580# diff_1141730_2763520# GND GND efet w=24130 l=7620
+ ad=2.66128e+08 pd=76200 as=0 ps=0 
M1200 diff_580390_2753360# diff_1183640_1584960# diff_1141730_2763520# GND efet w=10160 l=7620
+ ad=0 pd=0 as=3.01612e+08 ps=78740 
M1201 diff_1223010_2766060# diff_1214120_1543050# diff_580390_2753360# GND efet w=12065 l=6985
+ ad=2.88709e+08 pd=76200 as=0 ps=0 
M1202 diff_702310_2763520# diff_1145540_1527810# diff_1151890_2735580# GND efet w=22860 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1203 diff_1103630_2694940# diff_1092200_1543050# diff_703580_2682240# GND efet w=22860 l=8890
+ ad=2.67741e+08 pd=78740 as=0 ps=0 
M1204 diff_703580_2682240# diff_1145540_1527810# diff_1151890_2691130# GND efet w=22860 l=9525
+ ad=0 pd=0 as=2.66128e+08 ps=76200 
M1205 diff_580390_2682240# diff_1038860_1543050# diff_995680_2675890# GND efet w=8890 l=8890
+ ad=0 pd=0 as=3.04838e+08 ps=81280 
M1206 diff_1076960_2675890# diff_1068070_1543050# diff_580390_2682240# GND efet w=8890 l=7620
+ ad=2.90322e+08 pd=81280 as=0 ps=0 
M1207 diff_580390_2603500# diff_1038860_1543050# diff_995680_2614930# GND efet w=8890 l=8890
+ ad=0 pd=0 as=2.80645e+08 ps=81280 
M1208 diff_1076960_2616200# diff_1068070_1543050# diff_580390_2603500# GND efet w=8890 l=7620
+ ad=2.88709e+08 pd=83820 as=0 ps=0 
M1209 diff_702310_2614930# diff_1000760_1526540# diff_1005840_2585720# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1210 diff_957580_2546350# diff_946150_1543050# diff_703580_2532380# GND efet w=22860 l=7620
+ ad=3.03225e+08 pd=81280 as=0 ps=0 
M1211 GND diff_932180_2526030# diff_957580_2546350# GND efet w=24765 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1212 diff_580390_2532380# diff_892810_1584960# diff_850900_2526030# GND efet w=8890 l=7620
+ ad=0 pd=0 as=3.03225e+08 ps=81280 
M1213 diff_932180_2526030# diff_923290_1543050# diff_580390_2532380# GND efet w=8890 l=7620
+ ad=2.87096e+08 pd=76200 as=0 ps=0 
M1214 diff_580390_2454910# diff_892810_1584960# diff_850900_2463800# GND efet w=8890 l=7620
+ ad=0 pd=0 as=3.03225e+08 ps=78740 
M1215 diff_932180_2466340# diff_923290_1543050# diff_580390_2454910# GND efet w=8890 l=7620
+ ad=2.90322e+08 pd=76200 as=0 ps=0 
M1216 diff_600710_2443480# diff_703580_2463800# GND GND efet w=28575 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1217 diff_861060_2435860# diff_850900_2463800# GND GND efet w=24130 l=7620
+ ad=2.6129e+08 pd=76200 as=0 ps=0 
M1218 GND diff_600710_2406650# diff_535940_2382520# GND efet w=53340 l=8890
+ ad=0 pd=0 as=1.84677e+09 ps=340360 
M1219 diff_703580_2463800# diff_854710_1527810# diff_861060_2435860# GND efet w=22860 l=8890
+ ad=-1.33188e+09 pd=1.63322e+06 as=0 ps=0 
M1220 diff_515620_2338070# diff_346710_1485900# diff_243840_2250440# GND efet w=39370 l=7620
+ ad=1.08871e+09 pd=241300 as=0 ps=0 
M1221 diff_515620_2390140# diff_553720_1553210# diff_535940_2382520# GND efet w=39370 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1222 diff_580390_2383790# diff_450850_1684020# diff_515620_2390140# GND efet w=49530 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1223 GND diff_346710_1485900# diff_466090_2289810# GND efet w=59690 l=7620
+ ad=0 pd=0 as=5.93547e+08 ps=129540 
M1224 diff_515620_2338070# diff_553720_1553210# diff_535940_2313940# GND efet w=40640 l=7620
+ ad=0 pd=0 as=1.87903e+09 ps=347980 
M1225 diff_580390_2305050# diff_450850_1684020# diff_515620_2338070# GND efet w=48260 l=7620
+ ad=-7.7562e+08 pd=916940 as=0 ps=0 
M1226 GND diff_703580_2382520# diff_600710_2406650# GND efet w=27940 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1227 diff_535940_2382520# diff_703580_2382520# Vdd GND efet w=14605 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1228 diff_861060_2391410# diff_850900_2376170# GND GND efet w=25400 l=7620
+ ad=2.70967e+08 pd=78740 as=0 ps=0 
M1229 diff_703580_2382520# diff_854710_1527810# diff_861060_2391410# GND efet w=22860 l=8890
+ ad=-1.71575e+09 pd=1.61798e+06 as=0 ps=0 
M1230 diff_600710_2406650# Vdd Vdd GND efet w=6350 l=27940
+ ad=0 pd=0 as=0 ps=0 
M1231 Vdd Vdd Vdd GND efet w=6350 l=3810
+ ad=0 pd=0 as=0 ps=0 
M1232 Vdd Vdd Vdd GND efet w=3810 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1233 diff_601980_2293620# Vdd Vdd GND efet w=6350 l=27940
+ ad=1.08548e+09 pd=246380 as=0 ps=0 
M1234 diff_601980_2293620# diff_448310_2263140# diff_580390_2305050# GND efet w=35560 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1235 diff_466090_2289810# diff_450850_1684020# diff_448310_2263140# GND efet w=49530 l=8890
+ ad=0 pd=0 as=1.07742e+09 ps=215900 
M1236 GND diff_172720_2129790# diff_243840_2250440# GND efet w=40640 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1237 d2 GND GND GND efet w=111760 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1238 diff_243840_2250440# diff_180340_2162810# Vdd GND efet w=40640 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1239 Vdd Vdd diff_448310_2263140# GND efet w=12700 l=40640
+ ad=0 pd=0 as=0 ps=0 
M1240 Vdd Vdd Vdd GND efet w=2540 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1241 Vdd Vdd Vdd GND efet w=1905 l=3810
+ ad=0 pd=0 as=0 ps=0 
M1242 Vdd diff_703580_2313940# diff_535940_2313940# GND efet w=14605 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1243 diff_535940_2313940# diff_601980_2293620# GND GND efet w=55880 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1244 diff_1005840_2548890# diff_995680_2526030# GND GND efet w=27305 l=9525
+ ad=2.88709e+08 pd=83820 as=0 ps=0 
M1245 diff_703580_2532380# diff_1000760_1526540# diff_1005840_2548890# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1246 diff_957580_2432050# diff_946150_1543050# diff_703580_2463800# GND efet w=22860 l=7620
+ ad=2.96774e+08 pd=81280 as=0 ps=0 
M1247 GND diff_932180_2466340# diff_957580_2432050# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1248 diff_1007110_2435860# diff_995680_2465070# GND GND efet w=24130 l=8890
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1249 GND diff_1076960_2675890# diff_1103630_2694940# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1250 diff_1151890_2691130# diff_1140460_2679700# GND GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1251 diff_1103630_2581910# diff_1092200_1543050# diff_702310_2614930# GND efet w=22860 l=7620
+ ad=2.66128e+08 pd=76200 as=0 ps=0 
M1252 GND diff_1076960_2616200# diff_1103630_2581910# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1253 diff_1151890_2585720# diff_1141730_2613660# GND GND efet w=24130 l=7620
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1254 diff_1248410_2731770# diff_1236980_1543050# diff_702310_2763520# GND efet w=22860 l=7620
+ ad=2.96774e+08 pd=78740 as=0 ps=0 
M1255 GND diff_1223010_2766060# diff_1248410_2731770# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1256 diff_1297940_2735580# diff_1286510_2763520# GND GND efet w=24130 l=8890
+ ad=2.66128e+08 pd=78740 as=0 ps=0 
M1257 diff_580390_2753360# diff_1329690_1543050# diff_1286510_2763520# GND efet w=10160 l=8255
+ ad=0 pd=0 as=2.88709e+08 ps=81280 
M1258 diff_1367790_2766060# diff_1358900_1543050# diff_580390_2753360# GND efet w=10160 l=7620
+ ad=2.8387e+08 pd=78740 as=0 ps=0 
M1259 diff_702310_2763520# diff_1291590_1526540# diff_1297940_2735580# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1260 diff_1248410_2696210# diff_1236980_1543050# diff_703580_2682240# GND efet w=22860 l=7620
+ ad=2.96774e+08 pd=78740 as=0 ps=0 
M1261 diff_580390_2682240# diff_1183640_1584960# diff_1140460_2679700# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.98386e+08 ps=78740 
M1262 diff_1223010_2675890# diff_1214120_1543050# diff_580390_2682240# GND efet w=10160 l=7620
+ ad=2.8387e+08 pd=76200 as=0 ps=0 
M1263 diff_580390_2603500# diff_1183640_1584960# diff_1141730_2613660# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.99999e+08 ps=78740 
M1264 diff_1223010_2616200# diff_1214120_1543050# diff_580390_2603500# GND efet w=9525 l=7620
+ ad=2.80645e+08 pd=78740 as=0 ps=0 
M1265 diff_702310_2614930# diff_1145540_1527810# diff_1151890_2585720# GND efet w=22860 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1266 diff_1103630_2545080# diff_1092200_1543050# diff_703580_2532380# GND efet w=22860 l=7620
+ ad=2.75806e+08 pd=78740 as=0 ps=0 
M1267 diff_1076960_2526030# diff_1068070_1543050# diff_580390_2532380# GND efet w=8890 l=8255
+ ad=2.90322e+08 pd=81280 as=0 ps=0 
M1268 diff_580390_2532380# diff_1038860_1543050# diff_995680_2526030# GND efet w=8890 l=8890
+ ad=0 pd=0 as=2.98386e+08 ps=81280 
M1269 diff_580390_2454910# diff_1038860_1543050# diff_995680_2465070# GND efet w=8890 l=8890
+ ad=0 pd=0 as=2.93548e+08 ps=81280 
M1270 diff_1076960_2466340# diff_1068070_1543050# diff_580390_2454910# GND efet w=8890 l=7620
+ ad=2.93548e+08 pd=81280 as=0 ps=0 
M1271 diff_703580_2463800# diff_1000760_1526540# diff_1007110_2435860# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1272 diff_957580_2396490# diff_946150_1543050# diff_703580_2382520# GND efet w=21590 l=7620
+ ad=2.96774e+08 pd=78740 as=0 ps=0 
M1273 diff_703580_2382520# diff_1000760_1526540# diff_1007110_2391410# GND efet w=22225 l=9525
+ ad=0 pd=0 as=2.69354e+08 ps=78740 
M1274 GND diff_932180_2376170# diff_957580_2396490# GND efet w=24765 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1275 diff_580390_2383790# diff_892810_1584960# diff_850900_2376170# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.95161e+08 ps=78740 
M1276 diff_932180_2376170# diff_923290_1543050# diff_580390_2383790# GND efet w=8890 l=7620
+ ad=2.88709e+08 pd=78740 as=0 ps=0 
M1277 diff_580390_2305050# diff_892810_1584960# diff_850900_2315210# GND efet w=10160 l=7620
+ ad=0 pd=0 as=2.91935e+08 ps=78740 
M1278 diff_932180_2316480# diff_923290_1543050# diff_580390_2305050# GND efet w=10160 l=7620
+ ad=2.87096e+08 pd=76200 as=0 ps=0 
M1279 diff_1007110_2391410# diff_995680_2377440# GND GND efet w=25400 l=9525
+ ad=0 pd=0 as=0 ps=0 
M1280 diff_601980_2293620# diff_703580_2313940# GND GND efet w=28575 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1281 diff_601980_2251710# diff_448310_2263140# diff_580390_2232660# GND efet w=35560 l=8890
+ ad=1.04839e+09 pd=246380 as=-7.77232e+08 ps=927100 
M1282 GND diff_601980_2251710# diff_535940_2232660# GND efet w=55245 l=7620
+ ad=0 pd=0 as=1.88871e+09 ps=342900 
M1283 diff_861060_2286000# diff_850900_2315210# GND GND efet w=25400 l=8890
+ ad=2.91935e+08 pd=78740 as=0 ps=0 
M1284 diff_703580_2313940# diff_854710_1527810# diff_861060_2286000# GND efet w=22225 l=8255
+ ad=-1.44963e+09 pd=1.63068e+06 as=0 ps=0 
M1285 diff_515620_2207260# diff_346710_1485900# diff_245110_1436370# GND efet w=41275 l=8255
+ ad=1.11451e+09 pd=241300 as=0 ps=0 
M1286 diff_180340_2162810# diff_172720_2129790# GND GND efet w=22860 l=7620
+ ad=1.68709e+09 pd=292100 as=0 ps=0 
M1287 diff_180340_2162810# diff_180340_2162810# diff_180340_2162810# GND efet w=2540 l=3810
+ ad=0 pd=0 as=0 ps=0 
M1288 diff_180340_2162810# diff_180340_2162810# diff_180340_2162810# GND efet w=2540 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1289 Vdd Vdd diff_180340_2162810# GND efet w=8890 l=39370
+ ad=0 pd=0 as=0 ps=0 
M1290 diff_515620_2207260# diff_553720_1553210# diff_535940_2232660# GND efet w=40640 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1291 diff_580390_2232660# diff_450850_1684020# diff_515620_2207260# GND efet w=47625 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1292 GND diff_703580_2232660# diff_601980_2251710# GND efet w=29210 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1293 diff_861060_2242820# diff_850900_2226310# GND GND efet w=24130 l=7620
+ ad=2.91935e+08 pd=78740 as=0 ps=0 
M1294 diff_703580_2232660# diff_854710_1527810# diff_861060_2242820# GND efet w=22860 l=7620
+ ad=-1.36898e+09 pd=1.64084e+06 as=0 ps=0 
M1295 diff_535940_2232660# diff_703580_2232660# Vdd GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1296 diff_601980_2251710# Vdd Vdd GND efet w=6350 l=27940
+ ad=0 pd=0 as=0 ps=0 
M1297 diff_172720_2129790# diff_172720_2129790# diff_172720_2129790# GND efet w=2540 l=7620
+ ad=1.34193e+09 pd=297180 as=0 ps=0 
M1298 diff_172720_2129790# diff_172720_2129790# diff_172720_2129790# GND efet w=1905 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1299 diff_172720_2129790# d2 GND GND efet w=59690 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1300 diff_180340_2162810# diff_139700_2962910# GND GND efet w=36830 l=6985
+ ad=0 pd=0 as=0 ps=0 
M1301 diff_515620_2147570# diff_350520_1598930# diff_369570_1160780# GND efet w=40640 l=7620
+ ad=1.22903e+09 pd=261620 as=0 ps=0 
M1302 diff_515620_2147570# diff_553720_1553210# diff_535940_2156460# GND efet w=40640 l=7620
+ ad=0 pd=0 as=1.88387e+09 ps=345440 
M1303 Vdd Vdd Vdd GND efet w=6350 l=3810
+ ad=0 pd=0 as=0 ps=0 
M1304 diff_580390_2155190# diff_450850_1684020# diff_515620_2147570# GND efet w=47625 l=8255
+ ad=-7.27233e+08 pd=914400 as=0 ps=0 
M1305 Vdd Vdd Vdd GND efet w=3810 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1306 diff_601980_2143760# Vdd Vdd GND efet w=6985 l=28575
+ ad=9.80643e+08 pd=231140 as=0 ps=0 
M1307 Vdd diff_703580_2164080# diff_535940_2156460# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1308 diff_601980_2143760# diff_448310_1962150# diff_580390_2155190# GND efet w=33655 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1309 GND diff_139700_2962910# diff_172720_2129790# GND efet w=36830 l=6985
+ ad=0 pd=0 as=0 ps=0 
M1310 GND GND GND GND efet w=635 l=1905
+ ad=0 pd=0 as=0 ps=0 
M1311 Vdd Vdd Vdd GND efet w=2540 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1312 Vdd Vdd Vdd GND efet w=1905 l=5080
+ ad=0 pd=0 as=0 ps=0 
M1313 Vdd Vdd diff_172720_2129790# GND efet w=8890 l=38100
+ ad=0 pd=0 as=0 ps=0 
M1314 diff_515620_2090420# diff_350520_1598930# diff_266700_2927350# GND efet w=39370 l=7620
+ ad=1.09032e+09 pd=236220 as=0 ps=0 
M1315 diff_535940_2156460# diff_601980_2143760# GND GND efet w=55880 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1316 diff_601980_2143760# diff_703580_2164080# GND GND efet w=29845 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1317 diff_861060_2136140# diff_850900_2164080# GND GND efet w=26035 l=8255
+ ad=2.96774e+08 pd=81280 as=0 ps=0 
M1318 diff_957580_2282190# diff_946150_1543050# diff_703580_2313940# GND efet w=24130 l=8255
+ ad=2.7258e+08 pd=81280 as=0 ps=0 
M1319 GND diff_932180_2316480# diff_957580_2282190# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1320 diff_1007110_2286000# diff_995680_2315210# GND GND efet w=24130 l=8890
+ ad=2.62903e+08 pd=78740 as=0 ps=0 
M1321 GND diff_1076960_2526030# diff_1103630_2545080# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1322 diff_1151890_2541270# diff_1141730_2526030# GND GND efet w=24765 l=8255
+ ad=2.7258e+08 pd=78740 as=0 ps=0 
M1323 diff_703580_2532380# diff_1145540_1527810# diff_1151890_2541270# GND efet w=24765 l=9525
+ ad=0 pd=0 as=0 ps=0 
M1324 GND diff_1223010_2675890# diff_1248410_2696210# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1325 diff_1297940_2691130# diff_1286510_2675890# GND GND efet w=24130 l=8890
+ ad=2.66128e+08 pd=78740 as=0 ps=0 
M1326 diff_703580_2682240# diff_1291590_1526540# diff_1297940_2691130# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1327 diff_1248410_2581910# diff_1236980_1543050# diff_702310_2614930# GND efet w=22860 l=7620
+ ad=2.93548e+08 pd=78740 as=0 ps=0 
M1328 GND diff_1223010_2616200# diff_1248410_2581910# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1329 diff_1297940_2585720# diff_1286510_2614930# GND GND efet w=24130 l=8890
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1330 diff_1394460_2731770# diff_1383030_1543050# diff_702310_2763520# GND efet w=22860 l=7620
+ ad=2.67741e+08 pd=78740 as=0 ps=0 
M1331 GND diff_1367790_2766060# diff_1394460_2731770# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1332 diff_1442720_2735580# diff_1432560_2763520# GND GND efet w=24130 l=7620
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1333 diff_580390_2753360# diff_1474470_1583690# diff_1432560_2763520# GND efet w=10160 l=7620
+ ad=0 pd=0 as=3.01612e+08 ps=78740 
M1334 diff_1513840_2766060# diff_1504950_1543050# diff_580390_2753360# GND efet w=10160 l=8255
+ ad=2.88709e+08 pd=76200 as=0 ps=0 
M1335 diff_702310_2763520# diff_1436370_1529080# diff_1442720_2735580# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1336 diff_1394460_2696210# diff_1383030_1543050# diff_703580_2682240# GND efet w=22225 l=8255
+ ad=2.66128e+08 pd=78740 as=0 ps=0 
M1337 diff_580390_2682240# diff_1329690_1543050# diff_1286510_2675890# GND efet w=8890 l=10160
+ ad=0 pd=0 as=2.80645e+08 ps=78740 
M1338 diff_1367790_2675890# diff_1358900_1543050# diff_580390_2682240# GND efet w=8890 l=8890
+ ad=2.85483e+08 pd=81280 as=0 ps=0 
M1339 diff_580390_2603500# diff_1329690_1543050# diff_1286510_2614930# GND efet w=8890 l=8890
+ ad=0 pd=0 as=2.82258e+08 ps=78740 
M1340 diff_1367790_2616200# diff_1358900_1543050# diff_580390_2603500# GND efet w=8890 l=7620
+ ad=2.88709e+08 pd=81280 as=0 ps=0 
M1341 diff_702310_2614930# diff_1291590_1526540# diff_1297940_2585720# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1342 diff_1248410_2546350# diff_1236980_1543050# diff_703580_2532380# GND efet w=22225 l=7620
+ ad=2.98386e+08 pd=78740 as=0 ps=0 
M1343 diff_703580_2532380# diff_1291590_1526540# diff_1297940_2541270# GND efet w=22860 l=10160
+ ad=0 pd=0 as=2.67741e+08 ps=78740 
M1344 diff_580390_2532380# diff_1183640_1584960# diff_1141730_2526030# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.98386e+08 ps=78740 
M1345 diff_1223010_2526030# diff_1214120_1543050# diff_580390_2532380# GND efet w=10160 l=8890
+ ad=2.87096e+08 pd=76200 as=0 ps=0 
M1346 diff_1103630_2432050# diff_1092200_1543050# diff_703580_2463800# GND efet w=22860 l=7620
+ ad=2.67741e+08 pd=78740 as=0 ps=0 
M1347 GND diff_1076960_2466340# diff_1103630_2432050# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1348 diff_1151890_2434590# diff_1141730_2463800# GND GND efet w=24130 l=7620
+ ad=2.67741e+08 pd=78740 as=0 ps=0 
M1349 diff_580390_2454910# diff_1183640_1584960# diff_1141730_2463800# GND efet w=8890 l=7620
+ ad=0 pd=0 as=3.01612e+08 ps=78740 
M1350 diff_1223010_2466340# diff_1214120_1543050# diff_580390_2454910# GND efet w=8890 l=8890
+ ad=2.90322e+08 pd=76200 as=0 ps=0 
M1351 diff_703580_2463800# diff_1145540_1527810# diff_1151890_2434590# GND efet w=22860 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1352 diff_1103630_2395220# diff_1092200_1543050# diff_703580_2382520# GND efet w=22860 l=10160
+ ad=2.70967e+08 pd=78740 as=0 ps=0 
M1353 diff_703580_2382520# diff_1145540_1527810# diff_1151890_2391410# GND efet w=22225 l=10795
+ ad=0 pd=0 as=2.7258e+08 ps=78740 
M1354 diff_580390_2383790# diff_1038860_1543050# diff_995680_2377440# GND efet w=10160 l=8890
+ ad=0 pd=0 as=3.01612e+08 ps=86360 
M1355 diff_1076960_2376170# diff_1068070_1543050# diff_580390_2383790# GND efet w=8890 l=7620
+ ad=3.06451e+08 pd=83820 as=0 ps=0 
M1356 diff_580390_2305050# diff_1038860_1543050# diff_995680_2315210# GND efet w=11430 l=8255
+ ad=0 pd=0 as=2.98386e+08 ps=86360 
M1357 diff_1076960_2316480# diff_1068070_1543050# diff_580390_2305050# GND efet w=10160 l=7620
+ ad=2.90322e+08 pd=81280 as=0 ps=0 
M1358 diff_703580_2313940# diff_1000760_1526540# diff_1007110_2286000# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1359 diff_957580_2263140# diff_946150_1543050# diff_703580_2232660# GND efet w=25400 l=8890
+ ad=2.74193e+08 pd=81280 as=0 ps=0 
M1360 GND diff_932180_2227580# diff_957580_2263140# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1361 diff_1007110_2242820# diff_995680_2226310# GND GND efet w=24130 l=8890
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1362 diff_703580_2232660# diff_1000760_1526540# diff_1007110_2242820# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1363 diff_580390_2232660# diff_892810_1584960# diff_850900_2226310# GND efet w=10160 l=8255
+ ad=0 pd=0 as=3.03225e+08 ps=78740 
M1364 diff_932180_2227580# diff_923290_1543050# diff_580390_2232660# GND efet w=8890 l=7620
+ ad=2.85483e+08 pd=76200 as=0 ps=0 
M1365 diff_580390_2155190# diff_892810_1584960# diff_850900_2164080# GND efet w=9525 l=9525
+ ad=0 pd=0 as=3.03225e+08 ps=81280 
M1366 diff_932180_2166620# diff_923290_1543050# diff_580390_2155190# GND efet w=9525 l=8255
+ ad=2.88709e+08 pd=76200 as=0 ps=0 
M1367 diff_601980_2100580# diff_448310_1962150# diff_580390_2082800# GND efet w=34290 l=10160
+ ad=9.96772e+08 pd=228600 as=-7.20781e+08 ps=960120 
M1368 GND diff_601980_2100580# diff_535940_2082800# GND efet w=54610 l=7620
+ ad=0 pd=0 as=1.83225e+09 ps=345440 
M1369 diff_703580_2164080# diff_854710_1527810# diff_861060_2136140# GND efet w=22860 l=7620
+ ad=-1.38511e+09 pd=1.63068e+06 as=0 ps=0 
M1370 Vdd diff_72390_1687830# d3 GND efet w=648335 l=6985
+ ad=0 pd=0 as=-5.37782e+08 ps=3.20548e+06 
M1371 GND diff_73660_2023110# d3 GND efet w=1213485 l=4445
+ ad=0 pd=0 as=0 ps=0 
M1372 diff_515620_2037080# diff_350520_1598930# diff_243840_2250440# GND efet w=40640 l=7620
+ ad=1.12419e+09 pd=246380 as=0 ps=0 
M1373 diff_515620_2090420# diff_553720_1553210# diff_535940_2082800# GND efet w=39370 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1374 diff_580390_2082800# diff_450850_1684020# diff_515620_2090420# GND efet w=47625 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1375 diff_515620_2037080# diff_553720_1553210# diff_535940_2012950# GND efet w=43180 l=7620
+ ad=0 pd=0 as=1.87096e+09 ps=347980 
M1376 GND diff_703580_2081530# diff_601980_2100580# GND efet w=27940 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1377 diff_535940_2082800# diff_703580_2081530# Vdd GND efet w=15240 l=6985
+ ad=0 pd=0 as=0 ps=0 
M1378 diff_861060_2091690# diff_850900_2076450# GND GND efet w=25400 l=7620
+ ad=3.03225e+08 pd=81280 as=0 ps=0 
M1379 diff_703580_2081530# diff_854710_1527810# diff_861060_2091690# GND efet w=22860 l=7620
+ ad=-1.67382e+09 pd=1.6256e+06 as=0 ps=0 
M1380 Vdd Vdd Vdd GND efet w=6350 l=3810
+ ad=0 pd=0 as=0 ps=0 
M1381 GND diff_350520_1598930# diff_466090_1988820# GND efet w=55880 l=6985
+ ad=0 pd=0 as=6.11289e+08 ps=132080 
M1382 diff_580390_2004060# diff_450850_1684020# diff_515620_2037080# GND efet w=48895 l=8255
+ ad=-7.482e+08 pd=927100 as=0 ps=0 
M1383 diff_601980_2100580# Vdd Vdd GND efet w=7620 l=27940
+ ad=0 pd=0 as=0 ps=0 
M1384 Vdd Vdd Vdd GND efet w=3810 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1385 diff_601980_1992630# Vdd Vdd GND efet w=8255 l=28575
+ ad=1.10161e+09 pd=246380 as=0 ps=0 
M1386 diff_601980_1992630# diff_448310_1962150# diff_580390_2004060# GND efet w=34925 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1387 Vdd diff_703580_2012950# diff_535940_2012950# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1388 diff_466090_1988820# diff_450850_1684020# diff_448310_1962150# GND efet w=53975 l=8255
+ ad=0 pd=0 as=1.10322e+09 ps=223520 
M1389 Vdd Vdd diff_448310_1962150# GND efet w=12065 l=41275
+ ad=0 pd=0 as=0 ps=0 
M1390 Vdd Vdd Vdd GND efet w=2540 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1391 Vdd Vdd Vdd GND efet w=2540 l=4445
+ ad=0 pd=0 as=0 ps=0 
M1392 diff_535940_2012950# diff_601980_1992630# GND GND efet w=54610 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1393 diff_601980_1992630# diff_703580_2012950# GND GND efet w=28575 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1394 diff_861060_1986280# diff_850900_2014220# GND GND efet w=24130 l=7620
+ ad=2.95161e+08 pd=78740 as=0 ps=0 
M1395 diff_958850_2132330# diff_946150_1543050# diff_703580_2164080# GND efet w=22860 l=8890
+ ad=2.67741e+08 pd=78740 as=0 ps=0 
M1396 GND diff_932180_2166620# diff_958850_2132330# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1397 diff_1007110_2136140# diff_995680_2164080# GND GND efet w=26035 l=8255
+ ad=2.66128e+08 pd=78740 as=0 ps=0 
M1398 GND diff_1076960_2376170# diff_1103630_2395220# GND efet w=26035 l=9525
+ ad=0 pd=0 as=0 ps=0 
M1399 diff_1151890_2391410# diff_1141730_2376170# GND GND efet w=25400 l=10160
+ ad=0 pd=0 as=0 ps=0 
M1400 diff_1103630_2282190# diff_1092200_1543050# diff_703580_2313940# GND efet w=22860 l=7620
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1401 GND diff_1076960_2316480# diff_1103630_2282190# GND efet w=24765 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1402 diff_1151890_2286000# diff_1141730_2315210# GND GND efet w=24130 l=7620
+ ad=2.6129e+08 pd=76200 as=0 ps=0 
M1403 GND diff_1223010_2526030# diff_1248410_2546350# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1404 diff_1297940_2541270# diff_1286510_2526030# GND GND efet w=24130 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1405 diff_1248410_2432050# diff_1236980_1543050# diff_703580_2463800# GND efet w=27940 l=7620
+ ad=2.90322e+08 pd=88900 as=0 ps=0 
M1406 GND diff_1223010_2466340# diff_1248410_2432050# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1407 diff_1297940_2435860# diff_1286510_2465070# GND GND efet w=24130 l=8890
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1408 GND diff_1367790_2675890# diff_1394460_2696210# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1409 diff_1442720_2691130# diff_1432560_2675890# GND GND efet w=24130 l=7620
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1410 diff_703580_2682240# diff_1436370_1529080# diff_1442720_2691130# GND efet w=22225 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1411 diff_1394460_2581910# diff_1383030_1543050# diff_702310_2614930# GND efet w=22860 l=7620
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1412 GND diff_1367790_2616200# diff_1394460_2581910# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1413 diff_1442720_2585720# diff_1432560_2613660# GND GND efet w=24130 l=7620
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1414 diff_1539240_2731770# diff_1527810_1543050# diff_702310_2763520# GND efet w=22860 l=7620
+ ad=2.95161e+08 pd=78740 as=0 ps=0 
M1415 GND diff_1513840_2766060# diff_1539240_2731770# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1416 diff_1588770_2735580# diff_1577340_2764790# GND GND efet w=24130 l=8890
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1417 diff_580390_2753360# diff_1620520_1543050# diff_1577340_2764790# GND efet w=10795 l=8890
+ ad=0 pd=0 as=2.88709e+08 ps=81280 
M1418 diff_1658620_2766060# diff_1649730_1543050# diff_580390_2753360# GND efet w=9525 l=8255
+ ad=2.99999e+08 pd=78740 as=0 ps=0 
M1419 diff_702310_2763520# diff_1582420_1527810# diff_1588770_2735580# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1420 diff_1539240_2696210# diff_1527810_1543050# diff_703580_2682240# GND efet w=22225 l=8255
+ ad=2.93548e+08 pd=78740 as=0 ps=0 
M1421 diff_580390_2682240# diff_1474470_1583690# diff_1432560_2675890# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.93548e+08 ps=78740 
M1422 diff_1513840_2675890# diff_1504950_1543050# diff_580390_2682240# GND efet w=8890 l=8890
+ ad=2.85483e+08 pd=78740 as=0 ps=0 
M1423 diff_580390_2603500# diff_1474470_1583690# diff_1432560_2613660# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.95161e+08 ps=78740 
M1424 diff_1513840_2616200# diff_1504950_1543050# diff_580390_2603500# GND efet w=8890 l=8890
+ ad=2.85483e+08 pd=76200 as=0 ps=0 
M1425 diff_702310_2614930# diff_1436370_1529080# diff_1442720_2585720# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1426 diff_1394460_2546350# diff_1383030_1543050# diff_703580_2532380# GND efet w=22860 l=7620
+ ad=2.7258e+08 pd=78740 as=0 ps=0 
M1427 diff_580390_2532380# diff_1329690_1543050# diff_1286510_2526030# GND efet w=8890 l=8890
+ ad=0 pd=0 as=2.87096e+08 ps=81280 
M1428 diff_1367790_2526030# diff_1358900_1543050# diff_580390_2532380# GND efet w=8890 l=7620
+ ad=2.90322e+08 pd=81280 as=0 ps=0 
M1429 diff_580390_2454910# diff_1329690_1543050# diff_1286510_2465070# GND efet w=8890 l=8890
+ ad=0 pd=0 as=2.91935e+08 ps=81280 
M1430 diff_1367790_2466340# diff_1358900_1543050# diff_580390_2454910# GND efet w=8890 l=7620
+ ad=2.88709e+08 pd=81280 as=0 ps=0 
M1431 diff_703580_2463800# diff_1291590_1526540# diff_1297940_2435860# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1432 diff_1248410_2400300# diff_1236980_1543050# diff_703580_2382520# GND efet w=24130 l=8890
+ ad=2.90322e+08 pd=81280 as=0 ps=0 
M1433 GND diff_1223010_2376170# diff_1248410_2400300# GND efet w=24765 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1434 diff_1297940_2391410# diff_1286510_2377440# GND GND efet w=25400 l=8890
+ ad=2.62903e+08 pd=78740 as=0 ps=0 
M1435 diff_703580_2382520# diff_1291590_1526540# diff_1297940_2391410# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1436 diff_580390_2383790# diff_1183640_1584960# diff_1141730_2376170# GND efet w=8890 l=7620
+ ad=0 pd=0 as=3.03225e+08 ps=81280 
M1437 diff_1223010_2376170# diff_1214120_1543050# diff_580390_2383790# GND efet w=10160 l=8255
+ ad=2.85483e+08 pd=76200 as=0 ps=0 
M1438 diff_580390_2305050# diff_1183640_1584960# diff_1141730_2315210# GND efet w=10160 l=7620
+ ad=0 pd=0 as=3.08064e+08 ps=81280 
M1439 diff_1223010_2316480# diff_1214120_1543050# diff_580390_2305050# GND efet w=10160 l=7620
+ ad=2.7258e+08 pd=73660 as=0 ps=0 
M1440 diff_703580_2313940# diff_1145540_1527810# diff_1151890_2286000# GND efet w=22860 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1441 diff_1103630_2246630# diff_1092200_1543050# diff_703580_2232660# GND efet w=22860 l=7620
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1442 diff_580390_2232660# diff_1038860_1543050# diff_995680_2226310# GND efet w=10795 l=7620
+ ad=0 pd=0 as=3.01612e+08 ps=86360 
M1443 diff_1076960_2226310# diff_1068070_1543050# diff_580390_2232660# GND efet w=8890 l=7620
+ ad=2.87096e+08 pd=81280 as=0 ps=0 
M1444 diff_580390_2155190# diff_1038860_1543050# diff_995680_2164080# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.99999e+08 ps=78740 
M1445 diff_1076960_2167890# diff_1068070_1543050# diff_580390_2155190# GND efet w=8890 l=7620
+ ad=2.82258e+08 pd=78740 as=0 ps=0 
M1446 diff_703580_2164080# diff_1000760_1526540# diff_1007110_2136140# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1447 diff_958850_2092960# diff_946150_1543050# diff_703580_2081530# GND efet w=23495 l=9525
+ ad=2.74193e+08 pd=78740 as=0 ps=0 
M1448 diff_580390_2082800# diff_892810_1584960# diff_850900_2076450# GND efet w=13335 l=16510
+ ad=0 pd=0 as=2.95161e+08 ps=78740 
M1449 diff_932180_2076450# diff_923290_1543050# diff_580390_2082800# GND efet w=8890 l=7620
+ ad=2.96774e+08 pd=78740 as=0 ps=0 
M1450 diff_580390_2004060# diff_892810_1584960# diff_850900_2014220# GND efet w=8890 l=8890
+ ad=0 pd=0 as=2.96774e+08 ps=78740 
M1451 diff_932180_2015490# diff_923290_1543050# diff_580390_2004060# GND efet w=8890 l=7620
+ ad=2.87096e+08 pd=76200 as=0 ps=0 
M1452 diff_703580_2012950# diff_854710_1527810# diff_861060_1986280# GND efet w=21590 l=7620
+ ad=-1.48511e+09 pd=1.61798e+06 as=0 ps=0 
M1453 diff_601980_1950720# diff_448310_1962150# diff_580390_1932940# GND efet w=33655 l=7620
+ ad=1.08548e+09 pd=246380 as=-7.982e+08 ps=919480 
M1454 GND diff_601980_1950720# diff_535940_1931670# GND efet w=54610 l=8890
+ ad=0 pd=0 as=1.88709e+09 ps=342900 
M1455 GND diff_703580_1931670# diff_601980_1950720# GND efet w=29210 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1456 diff_515620_1906270# diff_350520_1598930# diff_245110_1436370# GND efet w=41275 l=8255
+ ad=1.13226e+09 pd=243840 as=0 ps=0 
M1457 diff_515620_1906270# diff_553720_1553210# diff_535940_1931670# GND efet w=40640 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1458 diff_580390_1932940# diff_450850_1684020# diff_515620_1906270# GND efet w=47625 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1459 diff_535940_1931670# diff_703580_1931670# Vdd GND efet w=14605 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1460 diff_861060_1941830# diff_850900_1925320# GND GND efet w=24130 l=7620
+ ad=2.91935e+08 pd=78740 as=0 ps=0 
M1461 diff_703580_1931670# diff_854710_1527810# diff_861060_1941830# GND efet w=22860 l=7620
+ ad=-1.37543e+09 pd=1.62814e+06 as=0 ps=0 
M1462 diff_601980_1950720# Vdd Vdd GND efet w=6985 l=29210
+ ad=0 pd=0 as=0 ps=0 
M1463 diff_72390_1687830# diff_93980_1783080# GND GND efet w=231140 l=7620
+ ad=2.06637e+08 pd=843280 as=0 ps=0 
M1464 diff_515620_1841500# diff_462280_1706880# diff_369570_1160780# GND efet w=39370 l=7620
+ ad=1.29193e+09 pd=274320 as=0 ps=0 
M1465 diff_515620_1841500# diff_553720_1553210# diff_535940_1849120# GND efet w=41910 l=7620
+ ad=0 pd=0 as=1.91129e+09 ps=355600 
M1466 Vdd Vdd Vdd GND efet w=6985 l=4445
+ ad=0 pd=0 as=0 ps=0 
M1467 diff_580390_1854200# diff_450850_1684020# diff_515620_1841500# GND efet w=47625 l=8255
+ ad=-7.56265e+08 pd=909320 as=0 ps=0 
M1468 Vdd Vdd Vdd GND efet w=3810 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1469 diff_601980_1842770# Vdd Vdd GND efet w=6350 l=27940
+ ad=9.88708e+08 pd=228600 as=0 ps=0 
M1470 Vdd diff_703580_1863090# diff_535940_1849120# GND efet w=14605 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1471 diff_93980_1783080# diff_93980_1783080# diff_93980_1783080# GND efet w=2540 l=5080
+ ad=1.32258e+09 pd=228600 as=0 ps=0 
M1472 diff_93980_1783080# diff_93980_1783080# diff_93980_1783080# GND efet w=3810 l=5080
+ ad=0 pd=0 as=0 ps=0 
M1473 diff_245110_1436370# diff_234950_1145540# diff_93980_1783080# GND efet w=29210 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1474 diff_515620_1789430# diff_462280_1706880# diff_266700_2927350# GND efet w=39370 l=7620
+ ad=1.08709e+09 pd=241300 as=0 ps=0 
M1475 diff_601980_1842770# diff_448310_1662430# diff_580390_1854200# GND efet w=33020 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1476 diff_601980_1800860# diff_448310_1662430# diff_580390_1783080# GND efet w=33655 l=8255
+ ad=9.7903e+08 pd=228600 as=-7.54652e+08 ps=916940 
M1477 diff_535940_1849120# diff_601980_1842770# GND GND efet w=53340 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1478 diff_601980_1842770# diff_703580_1863090# GND GND efet w=27940 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1479 GND diff_601980_1800860# diff_535940_1781810# GND efet w=54610 l=7620
+ ad=0 pd=0 as=1.83871e+09 ps=342900 
M1480 diff_861060_1835150# diff_850900_1863090# GND GND efet w=27305 l=8255
+ ad=2.99999e+08 pd=83820 as=0 ps=0 
M1481 GND diff_932180_2076450# diff_958850_2092960# GND efet w=24765 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1482 diff_1007110_2091690# diff_995680_2076450# GND GND efet w=27940 l=7620
+ ad=2.7258e+08 pd=78740 as=0 ps=0 
M1483 diff_703580_2081530# diff_1000760_1526540# diff_1007110_2091690# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1484 diff_958850_1981200# diff_946150_1543050# diff_703580_2012950# GND efet w=23495 l=9525
+ ad=2.77419e+08 pd=78740 as=0 ps=0 
M1485 GND diff_932180_2015490# diff_958850_1981200# GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1486 diff_1007110_1985010# diff_995680_2014220# GND GND efet w=27305 l=8255
+ ad=2.69354e+08 pd=78740 as=0 ps=0 
M1487 GND diff_1076960_2226310# diff_1103630_2246630# GND efet w=24130 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1488 diff_1151890_2242820# diff_1141730_2226310# GND GND efet w=24130 l=7620
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1489 diff_703580_2232660# diff_1145540_1527810# diff_1151890_2242820# GND efet w=22860 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1490 diff_1249680_2282190# diff_1236980_1543050# diff_703580_2313940# GND efet w=22860 l=8890
+ ad=2.66128e+08 pd=76200 as=0 ps=0 
M1491 GND diff_1223010_2316480# diff_1249680_2282190# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1492 diff_1297940_2286000# diff_1286510_2315210# GND GND efet w=24130 l=8890
+ ad=2.62903e+08 pd=78740 as=0 ps=0 
M1493 diff_703580_2532380# diff_1436370_1529080# diff_1442720_2541270# GND efet w=22860 l=10160
+ ad=0 pd=0 as=2.67741e+08 ps=78740 
M1494 GND diff_1367790_2526030# diff_1394460_2546350# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1495 diff_1442720_2541270# diff_1432560_2526030# GND GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1496 diff_1394460_2432050# diff_1383030_1543050# diff_703580_2463800# GND efet w=22860 l=7620
+ ad=2.66128e+08 pd=78740 as=0 ps=0 
M1497 GND diff_1367790_2466340# diff_1394460_2432050# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1498 diff_1442720_2435860# diff_1432560_2463800# GND GND efet w=24130 l=7620
+ ad=2.6129e+08 pd=76200 as=0 ps=0 
M1499 GND diff_1513840_2675890# diff_1539240_2696210# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1500 diff_1588770_2691130# diff_1577340_2675890# GND GND efet w=24130 l=8890
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1501 diff_703580_2682240# diff_1582420_1527810# diff_1588770_2691130# GND efet w=22225 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1502 diff_1539240_2581910# diff_1527810_1543050# diff_702310_2614930# GND efet w=22860 l=7620
+ ad=2.91935e+08 pd=78740 as=0 ps=0 
M1503 GND diff_1513840_2616200# diff_1539240_2581910# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1504 diff_1588770_2585720# diff_1577340_2614930# GND GND efet w=24130 l=8890
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1505 diff_1685290_2731770# diff_1673860_1543050# diff_702310_2763520# GND efet w=22860 l=7620
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1506 GND diff_1658620_2766060# diff_1685290_2731770# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1507 diff_1733550_2735580# diff_1723390_2763520# GND GND efet w=24130 l=7620
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1508 diff_580390_2753360# diff_1765300_1584960# diff_1723390_2763520# GND efet w=9525 l=8255
+ ad=0 pd=0 as=2.87096e+08 ps=81280 
M1509 diff_1804670_2766060# diff_1795780_1543050# diff_580390_2753360# GND efet w=9525 l=8255
+ ad=2.85483e+08 pd=78740 as=0 ps=0 
M1510 diff_702310_2763520# diff_1728470_1526540# diff_1733550_2735580# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1511 diff_1685290_2696210# diff_1673860_1543050# diff_703580_2682240# GND efet w=22225 l=8255
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1512 diff_580390_2682240# diff_1620520_1543050# diff_1577340_2675890# GND efet w=8890 l=8890
+ ad=0 pd=0 as=2.82258e+08 ps=76200 
M1513 diff_1658620_2675890# diff_1649730_1543050# diff_580390_2682240# GND efet w=8890 l=7620
+ ad=2.96774e+08 pd=78740 as=0 ps=0 
M1514 diff_580390_2603500# diff_1620520_1543050# diff_1577340_2614930# GND efet w=8890 l=8890
+ ad=0 pd=0 as=2.77419e+08 ps=81280 
M1515 diff_1658620_2616200# diff_1649730_1543050# diff_580390_2603500# GND efet w=8890 l=7620
+ ad=2.8387e+08 pd=78740 as=0 ps=0 
M1516 diff_702310_2614930# diff_1582420_1527810# diff_1588770_2585720# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1517 diff_1539240_2546350# diff_1527810_1543050# diff_703580_2532380# GND efet w=21590 l=7620
+ ad=2.91935e+08 pd=78740 as=0 ps=0 
M1518 diff_580390_2532380# diff_1474470_1583690# diff_1432560_2526030# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.95161e+08 ps=78740 
M1519 diff_1513840_2526030# diff_1504950_1543050# diff_580390_2532380# GND efet w=8890 l=8890
+ ad=2.8387e+08 pd=76200 as=0 ps=0 
M1520 diff_580390_2454910# diff_1474470_1583690# diff_1432560_2463800# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.98386e+08 ps=78740 
M1521 diff_1513840_2466340# diff_1504950_1543050# diff_580390_2454910# GND efet w=8890 l=8890
+ ad=2.85483e+08 pd=78740 as=0 ps=0 
M1522 diff_703580_2463800# diff_1436370_1529080# diff_1442720_2435860# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1523 diff_1394460_2396490# diff_1383030_1543050# diff_703580_2382520# GND efet w=21590 l=7620
+ ad=2.66128e+08 pd=78740 as=0 ps=0 
M1524 diff_580390_2383790# diff_1329690_1543050# diff_1286510_2377440# GND efet w=8890 l=8890
+ ad=0 pd=0 as=2.85483e+08 ps=81280 
M1525 diff_1367790_2376170# diff_1358900_1543050# diff_580390_2383790# GND efet w=8890 l=7620
+ ad=2.85483e+08 pd=81280 as=0 ps=0 
M1526 diff_580390_2305050# diff_1329690_1543050# diff_1286510_2315210# GND efet w=8890 l=8890
+ ad=0 pd=0 as=2.88709e+08 ps=81280 
M1527 diff_1367790_2316480# diff_1358900_1543050# diff_580390_2305050# GND efet w=8890 l=7620
+ ad=2.91935e+08 pd=81280 as=0 ps=0 
M1528 diff_703580_2313940# diff_1291590_1526540# diff_1297940_2286000# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1529 diff_1249680_2244090# diff_1236980_1543050# diff_703580_2232660# GND efet w=22860 l=8890
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1530 diff_580390_2232660# diff_1183640_1584960# diff_1141730_2226310# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.96774e+08 ps=78740 
M1531 diff_1223010_2226310# diff_1214120_1543050# diff_580390_2232660# GND efet w=8890 l=7620
+ ad=2.87096e+08 pd=76200 as=0 ps=0 
M1532 diff_1103630_2132330# diff_1092200_1543050# diff_703580_2164080# GND efet w=22860 l=7620
+ ad=2.67741e+08 pd=78740 as=0 ps=0 
M1533 GND diff_1076960_2167890# diff_1103630_2132330# GND efet w=24130 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1534 diff_1151890_2136140# diff_1141730_2164080# GND GND efet w=24130 l=7620
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1535 diff_580390_2155190# diff_1183640_1584960# diff_1141730_2164080# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.99999e+08 ps=78740 
M1536 diff_1223010_2167890# diff_1214120_1543050# diff_580390_2155190# GND efet w=8890 l=7620
+ ad=2.87096e+08 pd=76200 as=0 ps=0 
M1537 diff_703580_2164080# diff_1145540_1527810# diff_1151890_2136140# GND efet w=22860 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1538 diff_1103630_2096770# diff_1092200_1543050# diff_703580_2081530# GND efet w=23495 l=8255
+ ad=2.7258e+08 pd=78740 as=0 ps=0 
M1539 diff_703580_2081530# diff_1145540_1527810# diff_1151890_2091690# GND efet w=23495 l=9525
+ ad=0 pd=0 as=2.74193e+08 ps=81280 
M1540 GND diff_1076960_2076450# diff_1103630_2096770# GND efet w=24765 l=10795
+ ad=0 pd=0 as=0 ps=0 
M1541 diff_580390_2082800# diff_1038860_1543050# diff_995680_2076450# GND efet w=8890 l=7620
+ ad=0 pd=0 as=3.14515e+08 ps=83820 
M1542 diff_1076960_2076450# diff_1068070_1543050# diff_580390_2082800# GND efet w=8890 l=7620
+ ad=2.93548e+08 pd=83820 as=0 ps=0 
M1543 diff_580390_2004060# diff_1038860_1543050# diff_995680_2014220# GND efet w=9525 l=8255
+ ad=0 pd=0 as=3.03225e+08 ps=86360 
M1544 diff_1076960_2016760# diff_1068070_1543050# diff_580390_2004060# GND efet w=8890 l=7620
+ ad=2.85483e+08 pd=81280 as=0 ps=0 
M1545 diff_703580_2012950# diff_1000760_1526540# diff_1007110_1985010# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1546 diff_958850_1943100# diff_946150_1543050# diff_703580_1931670# GND efet w=22860 l=8890
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1547 diff_580390_1932940# diff_892810_1584960# diff_850900_1925320# GND efet w=8890 l=8890
+ ad=0 pd=0 as=3.01612e+08 ps=81280 
M1548 diff_932180_1926590# diff_923290_1543050# diff_580390_1932940# GND efet w=8890 l=7620
+ ad=2.91935e+08 pd=78740 as=0 ps=0 
M1549 GND diff_932180_1926590# diff_958850_1943100# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1550 diff_1007110_1941830# diff_995680_1925320# GND GND efet w=24130 l=7620
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1551 diff_703580_1931670# diff_1000760_1526540# diff_1007110_1941830# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1552 diff_580390_1854200# diff_892810_1584960# diff_850900_1863090# GND efet w=8890 l=8890
+ ad=0 pd=0 as=2.98386e+08 ps=78740 
M1553 diff_932180_1865630# diff_923290_1543050# diff_580390_1854200# GND efet w=8890 l=7620
+ ad=2.88709e+08 pd=76200 as=0 ps=0 
M1554 diff_703580_1863090# diff_854710_1527810# diff_861060_1835150# GND efet w=22860 l=7620
+ ad=-1.41576e+09 pd=1.62814e+06 as=0 ps=0 
M1555 diff_515620_1789430# diff_553720_1553210# diff_535940_1781810# GND efet w=41275 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1556 diff_72390_1687830# diff_92710_2421890# GND GND efet w=231140 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1557 Vdd diff_171450_1715770# diff_72390_1687830# GND efet w=11430 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1558 diff_72390_1687830# diff_171450_1715770# diff_72390_1687830# GND efet w=52705 l=17780
+ ad=0 pd=0 as=0 ps=0 
M1559 diff_171450_1715770# diff_171450_1715770# diff_171450_1715770# GND efet w=2540 l=8890
+ ad=2.56451e+08 pd=86360 as=0 ps=0 
M1560 Vdd Vdd diff_171450_1715770# GND efet w=8890 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1561 diff_171450_1715770# diff_171450_1715770# diff_171450_1715770# GND efet w=3810 l=4445
+ ad=0 pd=0 as=0 ps=0 
M1562 diff_73660_2023110# diff_72390_1687830# GND GND efet w=83820 l=6350
+ ad=-7.93361e+08 pd=642620 as=0 ps=0 
M1563 diff_73660_2023110# diff_92710_2421890# GND GND efet w=227330 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1564 diff_73660_2023110# diff_171450_1609090# diff_73660_2023110# GND efet w=41275 l=19685
+ ad=0 pd=0 as=0 ps=0 
M1565 Vdd diff_171450_1609090# diff_73660_2023110# GND efet w=11430 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1566 diff_171450_1609090# diff_171450_1609090# diff_171450_1609090# GND efet w=2540 l=10160
+ ad=2.37096e+08 pd=73660 as=0 ps=0 
M1567 Vdd Vdd diff_171450_1609090# GND efet w=8890 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1568 diff_171450_1609090# diff_171450_1609090# diff_171450_1609090# GND efet w=635 l=3175
+ ad=0 pd=0 as=0 ps=0 
M1569 diff_515620_1737360# diff_462280_1706880# diff_243840_2250440# GND efet w=39370 l=7620
+ ad=1.05484e+09 pd=238760 as=0 ps=0 
M1570 diff_580390_1783080# diff_450850_1684020# diff_515620_1789430# GND efet w=48260 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1571 GND diff_462280_1706880# diff_466090_1689100# GND efet w=55880 l=6985
+ ad=0 pd=0 as=6.22579e+08 ps=132080 
M1572 diff_515620_1737360# diff_553720_1553210# diff_535940_1713230# GND efet w=40640 l=8890
+ ad=0 pd=0 as=1.87419e+09 ps=345440 
M1573 diff_580390_1704340# diff_450850_1684020# diff_515620_1737360# GND efet w=47625 l=8255
+ ad=-8.482e+08 pd=911860 as=0 ps=0 
M1574 GND diff_703580_1781810# diff_601980_1800860# GND efet w=29845 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1575 diff_535940_1781810# diff_703580_1781810# Vdd GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1576 diff_861060_1790700# diff_850900_1775460# GND GND efet w=26670 l=7620
+ ad=2.98386e+08 pd=83820 as=0 ps=0 
M1577 diff_703580_1781810# diff_854710_1527810# diff_861060_1790700# GND efet w=22860 l=7620
+ ad=-1.68188e+09 pd=1.64592e+06 as=0 ps=0 
M1578 diff_601980_1800860# Vdd Vdd GND efet w=6350 l=27940
+ ad=0 pd=0 as=0 ps=0 
M1579 Vdd Vdd Vdd GND efet w=6350 l=3810
+ ad=0 pd=0 as=0 ps=0 
M1580 Vdd Vdd Vdd GND efet w=3810 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1581 diff_601980_1692910# Vdd Vdd GND efet w=7620 l=29210
+ ad=1.03871e+09 pd=241300 as=0 ps=0 
M1582 diff_601980_1692910# diff_448310_1662430# diff_580390_1704340# GND efet w=36195 l=9525
+ ad=0 pd=0 as=0 ps=0 
M1583 diff_466090_1689100# diff_450850_1684020# diff_448310_1662430# GND efet w=49530 l=7620
+ ad=0 pd=0 as=1.12097e+09 ps=215900 
M1584 Vdd Vdd diff_448310_1662430# GND efet w=12700 l=41910
+ ad=0 pd=0 as=0 ps=0 
M1585 Vdd Vdd Vdd GND efet w=1905 l=5715
+ ad=0 pd=0 as=0 ps=0 
M1586 Vdd Vdd Vdd GND efet w=1270 l=1270
+ ad=0 pd=0 as=0 ps=0 
M1587 Vdd Vdd Vdd GND efet w=3175 l=4445
+ ad=0 pd=0 as=0 ps=0 
M1588 Vdd diff_703580_1714500# diff_535940_1713230# GND efet w=14605 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1589 diff_535940_1713230# diff_601980_1692910# GND GND efet w=54610 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1590 diff_601980_1692910# diff_703580_1714500# GND GND efet w=27940 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1591 diff_601980_1651000# diff_448310_1662430# diff_580390_1633220# GND efet w=34290 l=7620
+ ad=1.08064e+09 pd=243840 as=-7.72394e+08 ps=911860 
M1592 diff_861060_1690370# diff_850900_1714500# GND GND efet w=26670 l=8255
+ ad=2.64516e+08 pd=81280 as=0 ps=0 
M1593 GND diff_932180_1865630# diff_958850_1831340# GND efet w=24765 l=8255
+ ad=0 pd=0 as=2.66128e+08 ps=78740 
M1594 diff_1007110_1835150# diff_995680_1864360# GND GND efet w=27305 l=8255
+ ad=2.7258e+08 pd=78740 as=0 ps=0 
M1595 diff_958850_1831340# diff_946150_1543050# diff_703580_1863090# GND efet w=24765 l=9525
+ ad=0 pd=0 as=0 ps=0 
M1596 diff_1151890_2091690# diff_1141730_2075180# GND GND efet w=24130 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1597 GND diff_1223010_2226310# diff_1249680_2244090# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1598 diff_1297940_2242820# diff_1286510_2226310# GND GND efet w=24130 l=8255
+ ad=2.6129e+08 pd=76200 as=0 ps=0 
M1599 diff_703580_2232660# diff_1291590_1526540# diff_1297940_2242820# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1600 diff_1249680_2132330# diff_1236980_1543050# diff_703580_2164080# GND efet w=22860 l=8890
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1601 GND diff_1223010_2167890# diff_1249680_2132330# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1602 diff_1297940_2136140# diff_1286510_2164080# GND GND efet w=27305 l=8255
+ ad=2.64516e+08 pd=78740 as=0 ps=0 
M1603 GND diff_1367790_2376170# diff_1394460_2396490# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1604 diff_1442720_2391410# diff_1432560_2376170# GND GND efet w=24130 l=7620
+ ad=2.66128e+08 pd=76200 as=0 ps=0 
M1605 diff_703580_2382520# diff_1436370_1529080# diff_1442720_2391410# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1606 GND diff_1513840_2526030# diff_1539240_2546350# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1607 diff_1587500_2561590# diff_1577340_2526030# GND GND efet w=25400 l=8255
+ ad=2.6129e+08 pd=81280 as=0 ps=0 
M1608 diff_703580_2532380# diff_1582420_1527810# diff_1587500_2561590# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1609 diff_1539240_2432050# diff_1527810_1543050# diff_703580_2463800# GND efet w=22860 l=7620
+ ad=2.90322e+08 pd=78740 as=0 ps=0 
M1610 GND diff_1513840_2466340# diff_1539240_2432050# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1611 diff_1588770_2435860# diff_1577340_2465070# GND GND efet w=24130 l=8890
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1612 GND diff_1658620_2675890# diff_1685290_2696210# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1613 diff_1733550_2691130# diff_1723390_2675890# GND GND efet w=24130 l=7620
+ ad=2.66128e+08 pd=78740 as=0 ps=0 
M1614 diff_703580_2682240# diff_1728470_1526540# diff_1733550_2691130# GND efet w=22225 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1615 diff_1685290_2581910# diff_1673860_1543050# diff_702310_2614930# GND efet w=22860 l=7620
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1616 GND diff_1658620_2616200# diff_1685290_2581910# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1617 diff_1733550_2585720# diff_1723390_2614930# GND GND efet w=24130 l=7620
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1618 diff_1830070_2739390# diff_1819910_1543050# diff_702310_2763520# GND efet w=27305 l=8255
+ ad=2.77419e+08 pd=88900 as=0 ps=0 
M1619 GND diff_1804670_2766060# diff_1830070_2739390# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1620 diff_1879600_2735580# diff_1868170_2764790# GND GND efet w=24130 l=7620
+ ad=2.66128e+08 pd=78740 as=0 ps=0 
M1621 diff_580390_2753360# diff_1911350_1583690# diff_1868170_2764790# GND efet w=10160 l=7620
+ ad=0 pd=0 as=2.98386e+08 ps=81280 
M1622 diff_1949450_2774950# diff_1941830_1543050# diff_580390_2753360# GND efet w=10795 l=8255
+ ad=2.90322e+08 pd=83820 as=0 ps=0 
M1623 diff_702310_2763520# diff_1873250_1527810# diff_1879600_2735580# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1624 diff_1830070_2696210# diff_1819910_1543050# diff_703580_2682240# GND efet w=26670 l=8255
+ ad=2.88709e+08 pd=88900 as=0 ps=0 
M1625 diff_580390_2682240# diff_1765300_1584960# diff_1723390_2675890# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.80645e+08 ps=78740 
M1626 diff_1804670_2675890# diff_1795780_1543050# diff_580390_2682240# GND efet w=8890 l=7620
+ ad=2.85483e+08 pd=81280 as=0 ps=0 
M1627 diff_580390_2603500# diff_1765300_1584960# diff_1723390_2614930# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.82258e+08 ps=81280 
M1628 diff_1804670_2616200# diff_1795780_1543050# diff_580390_2603500# GND efet w=8890 l=7620
+ ad=2.80645e+08 pd=78740 as=0 ps=0 
M1629 diff_702310_2614930# diff_1728470_1526540# diff_1733550_2585720# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1630 diff_1685290_2546350# diff_1673860_1543050# diff_703580_2532380# GND efet w=21590 l=8255
+ ad=2.69354e+08 pd=78740 as=0 ps=0 
M1631 diff_580390_2532380# diff_1620520_1543050# diff_1577340_2526030# GND efet w=8890 l=8255
+ ad=0 pd=0 as=2.85483e+08 ps=76200 
M1632 diff_1658620_2526030# diff_1649730_1543050# diff_580390_2532380# GND efet w=8890 l=7620
+ ad=2.96774e+08 pd=78740 as=0 ps=0 
M1633 diff_580390_2454910# diff_1620520_1543050# diff_1577340_2465070# GND efet w=8890 l=8890
+ ad=0 pd=0 as=2.90322e+08 ps=78740 
M1634 diff_1658620_2466340# diff_1649730_1543050# diff_580390_2454910# GND efet w=8890 l=7620
+ ad=2.91935e+08 pd=81280 as=0 ps=0 
M1635 diff_703580_2463800# diff_1582420_1527810# diff_1588770_2435860# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1636 diff_1539240_2396490# diff_1527810_1543050# diff_703580_2382520# GND efet w=21590 l=7620
+ ad=2.93548e+08 pd=78740 as=0 ps=0 
M1637 diff_580390_2383790# diff_1474470_1583690# diff_1432560_2376170# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.96774e+08 ps=81280 
M1638 diff_1513840_2376170# diff_1504950_1543050# diff_580390_2383790# GND efet w=8890 l=8890
+ ad=2.82258e+08 pd=76200 as=0 ps=0 
M1639 diff_1394460_2282190# diff_1383030_1543050# diff_703580_2313940# GND efet w=22860 l=7620
+ ad=2.64516e+08 pd=78740 as=0 ps=0 
M1640 GND diff_1367790_2316480# diff_1394460_2282190# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1641 diff_1442720_2286000# diff_1432560_2315210# GND GND efet w=24130 l=7620
+ ad=2.6129e+08 pd=76200 as=0 ps=0 
M1642 diff_580390_2305050# diff_1474470_1583690# diff_1432560_2315210# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.90322e+08 ps=83820 
M1643 diff_1513840_2316480# diff_1504950_1543050# diff_580390_2305050# GND efet w=8890 l=8890
+ ad=2.87096e+08 pd=76200 as=0 ps=0 
M1644 diff_703580_2313940# diff_1436370_1529080# diff_1442720_2286000# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1645 diff_1394460_2246630# diff_1383030_1543050# diff_703580_2232660# GND efet w=22860 l=7620
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1646 diff_1367790_2227580# diff_1358900_1543050# diff_580390_2232660# GND efet w=11430 l=13335
+ ad=2.90322e+08 pd=88900 as=0 ps=0 
M1647 diff_580390_2232660# diff_1329690_1543050# diff_1286510_2226310# GND efet w=8890 l=8890
+ ad=0 pd=0 as=2.90322e+08 ps=81280 
M1648 diff_580390_2155190# diff_1329690_1543050# diff_1286510_2164080# GND efet w=8890 l=7620
+ ad=0 pd=0 as=3.03225e+08 ps=83820 
M1649 diff_1367790_2166620# diff_1358900_1543050# diff_580390_2155190# GND efet w=8890 l=7620
+ ad=2.88709e+08 pd=78740 as=0 ps=0 
M1650 diff_703580_2164080# diff_1291590_1526540# diff_1297940_2136140# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1651 diff_1249680_2095500# diff_1236980_1543050# diff_703580_2081530# GND efet w=22860 l=10160
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1652 diff_703580_2081530# diff_1291590_1526540# diff_1297940_2091690# GND efet w=22225 l=9525
+ ad=0 pd=0 as=2.64516e+08 ps=78740 
M1653 diff_580390_2082800# diff_1183640_1584960# diff_1141730_2075180# GND efet w=8890 l=7620
+ ad=0 pd=0 as=3.09677e+08 ps=81280 
M1654 diff_1223010_2076450# diff_1214120_1543050# diff_580390_2082800# GND efet w=8890 l=7620
+ ad=2.96774e+08 pd=78740 as=0 ps=0 
M1655 diff_1103630_1981200# diff_1092200_1543050# diff_703580_2012950# GND efet w=22860 l=7620
+ ad=2.75806e+08 pd=78740 as=0 ps=0 
M1656 GND diff_1076960_2016760# diff_1103630_1981200# GND efet w=25400 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1657 diff_1151890_1985010# diff_1141730_2014220# GND GND efet w=25400 l=7620
+ ad=2.75806e+08 pd=81280 as=0 ps=0 
M1658 diff_580390_2004060# diff_1183640_1584960# diff_1141730_2014220# GND efet w=9525 l=7620
+ ad=0 pd=0 as=3.01612e+08 ps=81280 
M1659 diff_1223010_2015490# diff_1214120_1543050# diff_580390_2004060# GND efet w=8890 l=7620
+ ad=2.87096e+08 pd=76200 as=0 ps=0 
M1660 diff_703580_2012950# diff_1145540_1527810# diff_1151890_1985010# GND efet w=24130 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1661 diff_1103630_1945640# diff_1092200_1543050# diff_703580_1931670# GND efet w=22860 l=7620
+ ad=2.66128e+08 pd=76200 as=0 ps=0 
M1662 diff_580390_1932940# diff_1038860_1543050# diff_995680_1925320# GND efet w=8890 l=7620
+ ad=0 pd=0 as=3.01612e+08 ps=86360 
M1663 diff_1076960_1926590# diff_1068070_1543050# diff_580390_1932940# GND efet w=8890 l=7620
+ ad=2.87096e+08 pd=83820 as=0 ps=0 
M1664 diff_580390_1854200# diff_1038860_1543050# diff_995680_1864360# GND efet w=8890 l=7620
+ ad=0 pd=0 as=3.03225e+08 ps=83820 
M1665 diff_1076960_1866900# diff_1068070_1543050# diff_580390_1854200# GND efet w=8890 l=7620
+ ad=2.96774e+08 pd=78740 as=0 ps=0 
M1666 diff_703580_1863090# diff_1000760_1526540# diff_1007110_1835150# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1667 diff_958850_1791970# diff_946150_1543050# diff_703580_1781810# GND efet w=24130 l=10795
+ ad=2.70967e+08 pd=76200 as=0 ps=0 
M1668 diff_580390_1783080# diff_892810_1584960# diff_850900_1775460# GND efet w=8890 l=8890
+ ad=0 pd=0 as=2.96774e+08 ps=78740 
M1669 diff_932180_1775460# diff_923290_1543050# diff_580390_1783080# GND efet w=8890 l=7620
+ ad=2.85483e+08 pd=76200 as=0 ps=0 
M1670 GND diff_932180_1775460# diff_958850_1791970# GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1671 diff_1007110_1790700# diff_995680_1775460# GND GND efet w=27305 l=8255
+ ad=2.7258e+08 pd=78740 as=0 ps=0 
M1672 diff_703580_1781810# diff_1000760_1526540# diff_1007110_1790700# GND efet w=23495 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1673 diff_580390_1704340# diff_892810_1584960# diff_850900_1714500# GND efet w=8890 l=8890
+ ad=0 pd=0 as=2.96774e+08 ps=78740 
M1674 diff_932180_1715770# diff_923290_1543050# diff_580390_1704340# GND efet w=8890 l=7620
+ ad=2.88709e+08 pd=76200 as=0 ps=0 
M1675 diff_703580_1714500# diff_854710_1527810# diff_861060_1690370# GND efet w=22860 l=7620
+ ad=-1.62705e+09 pd=1.61798e+06 as=0 ps=0 
M1676 GND diff_601980_1651000# diff_535940_1631950# GND efet w=54610 l=7620
+ ad=0 pd=0 as=1.92419e+09 ps=345440 
M1677 diff_515620_1610360# diff_462280_1706880# diff_245110_1436370# GND efet w=42545 l=9525
+ ad=1.04032e+09 pd=241300 as=0 ps=0 
M1678 diff_515620_1610360# diff_553720_1553210# diff_535940_1631950# GND efet w=39370 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1679 diff_580390_1633220# diff_450850_1684020# diff_515620_1610360# GND efet w=47625 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1680 GND diff_703580_1633220# diff_601980_1651000# GND efet w=27940 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1681 diff_535940_1631950# diff_703580_1633220# Vdd GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1682 diff_862330_1642110# diff_850900_1626870# GND GND efet w=24130 l=8890
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1683 diff_703580_1633220# diff_854710_1527810# diff_862330_1642110# GND efet w=22860 l=7620
+ ad=-1.54801e+09 pd=1.63322e+06 as=0 ps=0 
M1684 diff_601980_1651000# Vdd Vdd GND efet w=6985 l=28575
+ ad=0 pd=0 as=0 ps=0 
M1685 Vdd Vdd Vdd GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M1686 Vdd Vdd Vdd GND efet w=1905 l=6985
+ ad=0 pd=0 as=0 ps=0 
M1687 diff_958850_1681480# diff_946150_1543050# diff_703580_1714500# GND efet w=22860 l=8890
+ ad=2.66128e+08 pd=76200 as=0 ps=0 
M1688 GND diff_932180_1715770# diff_958850_1681480# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1689 diff_1007110_1685290# diff_995680_1714500# GND GND efet w=27305 l=8255
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1690 GND diff_1076960_1926590# diff_1103630_1945640# GND efet w=24130 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1691 diff_1151890_1941830# diff_1141730_1925320# GND GND efet w=24130 l=7620
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1692 diff_703580_1931670# diff_1145540_1527810# diff_1151890_1941830# GND efet w=22860 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1693 GND diff_1223010_2076450# diff_1249680_2095500# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1694 diff_1297940_2091690# diff_1286510_2076450# GND GND efet w=26670 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1695 GND diff_1367790_2227580# diff_1394460_2246630# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1696 diff_1442720_2242820# diff_1432560_2226310# GND GND efet w=24130 l=7620
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1697 diff_703580_2232660# diff_1436370_1529080# diff_1442720_2242820# GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1698 GND diff_1513840_2376170# diff_1539240_2396490# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1699 diff_1588770_2391410# diff_1577340_2377440# GND GND efet w=24130 l=8890
+ ad=2.6129e+08 pd=78740 as=0 ps=0 
M1700 diff_703580_2382520# diff_1582420_1527810# diff_1588770_2391410# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1701 diff_1539240_2282190# diff_1527810_1543050# diff_703580_2313940# GND efet w=22860 l=7620
+ ad=2.91935e+08 pd=78740 as=0 ps=0 
M1702 GND diff_1513840_2316480# diff_1539240_2282190# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1703 diff_1588770_2286000# diff_1577340_2315210# GND GND efet w=24130 l=8890
+ ad=2.62903e+08 pd=78740 as=0 ps=0 
M1704 GND diff_1658620_2526030# diff_1685290_2546350# GND efet w=24130 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1705 diff_1733550_2541270# diff_1723390_2526030# GND GND efet w=24130 l=7620
+ ad=2.64516e+08 pd=78740 as=0 ps=0 
M1706 diff_703580_2532380# diff_1728470_1526540# diff_1733550_2541270# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1707 diff_1685290_2432050# diff_1673860_1543050# diff_703580_2463800# GND efet w=22860 l=7620
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1708 GND diff_1658620_2466340# diff_1685290_2432050# GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1709 diff_1733550_2435860# diff_1723390_2463800# GND GND efet w=24130 l=7620
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1710 GND diff_1804670_2675890# diff_1830070_2696210# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1711 diff_1879600_2691130# diff_1868170_2677160# GND GND efet w=24130 l=7620
+ ad=2.66128e+08 pd=78740 as=0 ps=0 
M1712 diff_703580_2682240# diff_1873250_1527810# diff_1879600_2691130# GND efet w=22225 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1713 diff_1830070_2581910# diff_1819910_1543050# diff_702310_2614930# GND efet w=22860 l=7620
+ ad=2.93548e+08 pd=78740 as=0 ps=0 
M1714 GND diff_1804670_2616200# diff_1830070_2581910# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1715 diff_1879600_2585720# diff_1868170_2614930# GND GND efet w=24130 l=7620
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1716 diff_1976120_2731770# diff_1964690_1543050# diff_702310_2763520# GND efet w=22860 l=7620
+ ad=2.93548e+08 pd=81280 as=0 ps=0 
M1717 GND diff_1949450_2774950# diff_1976120_2731770# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1718 diff_2025650_2735580# diff_2014220_2764790# GND GND efet w=24130 l=7620
+ ad=2.66128e+08 pd=78740 as=0 ps=0 
M1719 diff_580390_2753360# diff_2057400_1583690# diff_2014220_2764790# GND efet w=8255 l=8255
+ ad=0 pd=0 as=2.96774e+08 ps=78740 
M1720 diff_2095500_2767330# diff_2087880_1543050# diff_580390_2753360# GND efet w=8890 l=7620
+ ad=2.93548e+08 pd=83820 as=0 ps=0 
M1721 diff_702310_2763520# diff_2019300_1526540# diff_2025650_2735580# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1722 diff_1976120_2696210# diff_1964690_1543050# diff_703580_2682240# GND efet w=21590 l=7620
+ ad=2.98386e+08 pd=81280 as=0 ps=0 
M1723 diff_580390_2682240# diff_1911350_1583690# diff_1868170_2677160# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.96774e+08 ps=78740 
M1724 diff_1950720_2675890# diff_1941830_1543050# diff_580390_2682240# GND efet w=8890 l=8890
+ ad=2.85483e+08 pd=81280 as=0 ps=0 
M1725 diff_580390_2603500# diff_1911350_1583690# diff_1868170_2614930# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.96774e+08 ps=78740 
M1726 diff_1949450_2616200# diff_1941830_1543050# diff_580390_2603500# GND efet w=9525 l=8255
+ ad=2.8387e+08 pd=88900 as=0 ps=0 
M1727 diff_702310_2614930# diff_1873250_1527810# diff_1879600_2585720# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1728 diff_1830070_2547620# diff_1819910_1543050# diff_703580_2532380# GND efet w=21590 l=7620
+ ad=2.91935e+08 pd=81280 as=0 ps=0 
M1729 diff_703580_2532380# diff_1873250_1527810# diff_1879600_2541270# GND efet w=22860 l=8890
+ ad=0 pd=0 as=2.67741e+08 ps=78740 
M1730 diff_580390_2532380# diff_1765300_1584960# diff_1723390_2526030# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.8387e+08 ps=81280 
M1731 diff_1804670_2526030# diff_1795780_1543050# diff_580390_2532380# GND efet w=8890 l=7620
+ ad=2.90322e+08 pd=81280 as=0 ps=0 
M1732 diff_580390_2454910# diff_1765300_1584960# diff_1723390_2463800# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.69354e+08 ps=78740 
M1733 diff_1804670_2466340# diff_1795780_1543050# diff_580390_2454910# GND efet w=8890 l=7620
+ ad=2.67741e+08 pd=76200 as=0 ps=0 
M1734 diff_703580_2463800# diff_1728470_1526540# diff_1733550_2435860# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1735 diff_1685290_2396490# diff_1673860_1543050# diff_703580_2382520# GND efet w=21590 l=7620
+ ad=2.64516e+08 pd=78740 as=0 ps=0 
M1736 diff_580390_2383790# diff_1620520_1543050# diff_1577340_2377440# GND efet w=8890 l=8890
+ ad=0 pd=0 as=2.80645e+08 ps=78740 
M1737 diff_1658620_2376170# diff_1649730_1543050# diff_580390_2383790# GND efet w=8890 l=7620
+ ad=2.91935e+08 pd=78740 as=0 ps=0 
M1738 diff_580390_2305050# diff_1620520_1543050# diff_1577340_2315210# GND efet w=10160 l=7620
+ ad=0 pd=0 as=2.79032e+08 ps=78740 
M1739 diff_1658620_2316480# diff_1649730_1543050# diff_580390_2305050# GND efet w=8890 l=7620
+ ad=2.96774e+08 pd=78740 as=0 ps=0 
M1740 diff_703580_2313940# diff_1582420_1527810# diff_1588770_2286000# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1741 diff_1539240_2247900# diff_1527810_1543050# diff_703580_2232660# GND efet w=22860 l=7620
+ ad=2.90322e+08 pd=78740 as=0 ps=0 
M1742 diff_580390_2232660# diff_1474470_1583690# diff_1432560_2226310# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.95161e+08 ps=78740 
M1743 diff_1513840_2227580# diff_1504950_1543050# diff_580390_2232660# GND efet w=10160 l=7620
+ ad=2.93548e+08 pd=78740 as=0 ps=0 
M1744 diff_1394460_2132330# diff_1383030_1543050# diff_703580_2164080# GND efet w=22860 l=7620
+ ad=2.67741e+08 pd=78740 as=0 ps=0 
M1745 GND diff_1367790_2166620# diff_1394460_2132330# GND efet w=28575 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1746 diff_1442720_2136140# diff_1432560_2164080# GND GND efet w=24130 l=7620
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1747 diff_580390_2155190# diff_1474470_1583690# diff_1432560_2164080# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.98386e+08 ps=78740 
M1748 diff_1513840_2167890# diff_1504950_1543050# diff_580390_2155190# GND efet w=8890 l=7620
+ ad=2.90322e+08 pd=78740 as=0 ps=0 
M1749 diff_703580_2164080# diff_1436370_1529080# diff_1442720_2136140# GND efet w=22860 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1750 diff_1394460_2096770# diff_1383030_1543050# diff_703580_2081530# GND efet w=22860 l=8255
+ ad=2.67741e+08 pd=78740 as=0 ps=0 
M1751 GND diff_1367790_2076450# diff_1394460_2096770# GND efet w=28575 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1752 diff_580390_2082800# diff_1329690_1543050# diff_1286510_2076450# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.95161e+08 ps=81280 
M1753 diff_1367790_2076450# diff_1358900_1543050# diff_580390_2082800# GND efet w=8890 l=7620
+ ad=3.01612e+08 pd=81280 as=0 ps=0 
M1754 diff_1249680_1981200# diff_1236980_1543050# diff_703580_2012950# GND efet w=22860 l=8890
+ ad=2.74193e+08 pd=78740 as=0 ps=0 
M1755 GND diff_1223010_2015490# diff_1249680_1981200# GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1756 diff_1297940_1985010# diff_1286510_2014220# GND GND efet w=26035 l=8255
+ ad=2.69354e+08 pd=78740 as=0 ps=0 
M1757 diff_580390_2004060# diff_1329690_1543050# diff_1286510_2014220# GND efet w=10160 l=7620
+ ad=0 pd=0 as=3.06451e+08 ps=83820 
M1758 diff_1367790_2015490# diff_1358900_1543050# diff_580390_2004060# GND efet w=10160 l=7620
+ ad=3.08064e+08 pd=83820 as=0 ps=0 
M1759 diff_703580_2012950# diff_1291590_1526540# diff_1297940_1985010# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1760 diff_1249680_1944370# diff_1236980_1543050# diff_703580_1931670# GND efet w=23495 l=9525
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1761 diff_580390_1932940# diff_1183640_1584960# diff_1141730_1925320# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.98386e+08 ps=78740 
M1762 diff_1223010_1925320# diff_1214120_1543050# diff_580390_1932940# GND efet w=8890 l=7620
+ ad=2.91935e+08 pd=78740 as=0 ps=0 
M1763 diff_1103630_1831340# diff_1092200_1543050# diff_703580_1863090# GND efet w=22860 l=7620
+ ad=2.67741e+08 pd=78740 as=0 ps=0 
M1764 GND diff_1076960_1866900# diff_1103630_1831340# GND efet w=24130 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1765 diff_1151890_1835150# diff_1141730_1864360# GND GND efet w=24130 l=7620
+ ad=2.69354e+08 pd=78740 as=0 ps=0 
M1766 diff_580390_1854200# diff_1183640_1584960# diff_1141730_1864360# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.99999e+08 ps=78740 
M1767 diff_1223010_1865630# diff_1214120_1543050# diff_580390_1854200# GND efet w=8890 l=7620
+ ad=2.85483e+08 pd=78740 as=0 ps=0 
M1768 diff_703580_1863090# diff_1145540_1527810# diff_1151890_1835150# GND efet w=24130 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1769 diff_1103630_1795780# diff_1092200_1543050# diff_703580_1781810# GND efet w=22860 l=8255
+ ad=2.74193e+08 pd=78740 as=0 ps=0 
M1770 diff_580390_1783080# diff_1038860_1543050# diff_995680_1775460# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.93548e+08 ps=81280 
M1771 diff_1076960_1775460# diff_1068070_1543050# diff_580390_1783080# GND efet w=9525 l=7620
+ ad=2.95161e+08 pd=78740 as=0 ps=0 
M1772 diff_580390_1704340# diff_1038860_1543050# diff_995680_1714500# GND efet w=8890 l=7620
+ ad=0 pd=0 as=3.01612e+08 ps=83820 
M1773 diff_1078230_1715770# diff_1068070_1543050# diff_580390_1704340# GND efet w=8890 l=8890
+ ad=2.88709e+08 pd=81280 as=0 ps=0 
M1774 diff_703580_1714500# diff_1000760_1526540# diff_1007110_1685290# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1775 diff_958850_1642110# diff_946150_1543050# diff_703580_1633220# GND efet w=25400 l=8890
+ ad=2.74193e+08 pd=78740 as=0 ps=0 
M1776 diff_580390_1633220# diff_892810_1584960# diff_850900_1626870# GND efet w=8890 l=8890
+ ad=0 pd=0 as=2.96774e+08 ps=78740 
M1777 diff_932180_1625600# diff_923290_1543050# diff_580390_1633220# GND efet w=9525 l=8255
+ ad=2.87096e+08 pd=76200 as=0 ps=0 
M1778 GND diff_932180_1625600# diff_958850_1642110# GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1779 diff_1007110_1640840# diff_995680_1626870# GND GND efet w=26035 l=8255
+ ad=2.70967e+08 pd=78740 as=0 ps=0 
M1780 diff_703580_1633220# diff_1000760_1526540# diff_1007110_1640840# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1781 GND diff_1076960_1775460# diff_1103630_1795780# GND efet w=25400 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1782 diff_1151890_1790700# diff_1141730_1775460# GND GND efet w=25400 l=7620
+ ad=2.74193e+08 pd=78740 as=0 ps=0 
M1783 diff_703580_1781810# diff_1145540_1527810# diff_1151890_1790700# GND efet w=23495 l=9525
+ ad=0 pd=0 as=0 ps=0 
M1784 GND diff_1223010_1925320# diff_1249680_1944370# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1785 diff_1297940_1941830# diff_1286510_1925320# GND GND efet w=26035 l=8255
+ ad=2.6129e+08 pd=76200 as=0 ps=0 
M1786 diff_703580_1931670# diff_1291590_1526540# diff_1297940_1941830# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1787 diff_1249680_1831340# diff_1236980_1543050# diff_703580_1863090# GND efet w=22860 l=8890
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1788 GND diff_1223010_1865630# diff_1249680_1831340# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1789 diff_1297940_1835150# diff_1286510_1864360# GND GND efet w=28575 l=8255
+ ad=2.66128e+08 pd=78740 as=0 ps=0 
M1790 diff_1442720_2091690# diff_1432560_2076450# GND GND efet w=24130 l=7620
+ ad=2.69354e+08 pd=76200 as=0 ps=0 
M1791 diff_703580_2081530# diff_1436370_1529080# diff_1442720_2091690# GND efet w=22860 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1792 GND diff_1513840_2227580# diff_1539240_2247900# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1793 diff_1588770_2242820# diff_1577340_2226310# GND GND efet w=24130 l=8255
+ ad=2.6129e+08 pd=76200 as=0 ps=0 
M1794 diff_703580_2232660# diff_1582420_1527810# diff_1588770_2242820# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1795 diff_1539240_2132330# diff_1527810_1543050# diff_703580_2164080# GND efet w=22860 l=7620
+ ad=2.91935e+08 pd=78740 as=0 ps=0 
M1796 GND diff_1513840_2167890# diff_1539240_2132330# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1797 diff_1588770_2136140# diff_1577340_2164080# GND GND efet w=25400 l=8255
+ ad=2.6129e+08 pd=76200 as=0 ps=0 
M1798 GND diff_1658620_2376170# diff_1685290_2396490# GND efet w=27305 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1799 diff_1733550_2391410# diff_1723390_2376170# GND GND efet w=24130 l=7620
+ ad=2.66128e+08 pd=78740 as=0 ps=0 
M1800 diff_703580_2382520# diff_1728470_1526540# diff_1733550_2391410# GND efet w=22225 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1801 GND diff_1804670_2526030# diff_1830070_2547620# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1802 diff_1879600_2541270# diff_1868170_2527300# GND GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1803 diff_1830070_2432050# diff_1819910_1543050# diff_703580_2463800# GND efet w=24130 l=7620
+ ad=2.88709e+08 pd=81280 as=0 ps=0 
M1804 GND diff_1804670_2466340# diff_1830070_2432050# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1805 diff_1879600_2435860# diff_1868170_2465070# GND GND efet w=24130 l=7620
+ ad=2.66128e+08 pd=76200 as=0 ps=0 
M1806 GND diff_1950720_2675890# diff_1976120_2696210# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1807 diff_2025650_2691130# diff_2014220_2677160# GND GND efet w=24130 l=7620
+ ad=2.69354e+08 pd=78740 as=0 ps=0 
M1808 diff_703580_2682240# diff_2019300_1526540# diff_2025650_2691130# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1809 diff_1976120_2581910# diff_1964690_1543050# diff_702310_2614930# GND efet w=22860 l=7620
+ ad=2.95161e+08 pd=81280 as=0 ps=0 
M1810 GND diff_1949450_2616200# diff_1976120_2581910# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1811 diff_2025650_2585720# diff_2014220_2614930# GND GND efet w=24765 l=8255
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1812 diff_2122170_2731770# diff_2110740_1545590# diff_702310_2763520# GND efet w=22860 l=7620
+ ad=2.91935e+08 pd=81280 as=0 ps=0 
M1813 GND diff_2095500_2767330# diff_2122170_2731770# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1814 diff_2171700_2735580# diff_2160270_2764790# GND GND efet w=26670 l=7620
+ ad=2.59677e+08 pd=76200 as=0 ps=0 
M1815 diff_580390_2753360# diff_2203450_1583690# diff_2160270_2764790# GND efet w=7620 l=7620
+ ad=0 pd=0 as=2.88709e+08 ps=78740 
M1816 diff_2241550_2767330# diff_2233930_1543050# diff_580390_2753360# GND efet w=7620 l=7620
+ ad=2.85483e+08 pd=81280 as=0 ps=0 
M1817 diff_702310_2763520# diff_2165350_1529080# diff_2171700_2735580# GND efet w=22225 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1818 diff_2122170_2697480# diff_2110740_1545590# diff_703580_2682240# GND efet w=21590 l=7620
+ ad=2.91935e+08 pd=81280 as=0 ps=0 
M1819 diff_580390_2682240# diff_2057400_1583690# diff_2014220_2677160# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.91935e+08 ps=78740 
M1820 diff_2095500_2675890# diff_2087880_1543050# diff_580390_2682240# GND efet w=8890 l=7620
+ ad=2.88709e+08 pd=81280 as=0 ps=0 
M1821 diff_580390_2603500# diff_2057400_1583690# diff_2014220_2614930# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.88709e+08 ps=83820 
M1822 diff_2095500_2616200# diff_2087880_1543050# diff_580390_2603500# GND efet w=8890 l=7620
+ ad=2.90322e+08 pd=81280 as=0 ps=0 
M1823 diff_702310_2614930# diff_2019300_1526540# diff_2025650_2585720# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1824 diff_703580_2532380# diff_2019300_1526540# diff_2025650_2541270# GND efet w=22860 l=8890
+ ad=0 pd=0 as=2.62903e+08 ps=78740 
M1825 diff_1976120_2547620# diff_1964690_1543050# diff_703580_2532380# GND efet w=21590 l=7620
+ ad=2.88709e+08 pd=81280 as=0 ps=0 
M1826 GND diff_1949450_2528570# diff_1976120_2547620# GND efet w=24765 l=9525
+ ad=0 pd=0 as=0 ps=0 
M1827 diff_580390_2532380# diff_1911350_1583690# diff_1868170_2527300# GND efet w=8890 l=7620
+ ad=0 pd=0 as=3.08064e+08 ps=81280 
M1828 diff_1949450_2528570# diff_1941830_1543050# diff_580390_2532380# GND efet w=11430 l=8255
+ ad=2.88709e+08 pd=86360 as=0 ps=0 
M1829 diff_580390_2454910# diff_1911350_1583690# diff_1868170_2465070# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.85483e+08 ps=81280 
M1830 diff_1949450_2470150# diff_1941830_1543050# diff_580390_2454910# GND efet w=10160 l=7620
+ ad=2.8387e+08 pd=81280 as=0 ps=0 
M1831 diff_703580_2463800# diff_1873250_1527810# diff_1879600_2435860# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1832 diff_1830070_2396490# diff_1819910_1543050# diff_703580_2382520# GND efet w=22860 l=7620
+ ad=2.82258e+08 pd=83820 as=0 ps=0 
M1833 diff_580390_2383790# diff_1765300_1584960# diff_1723390_2376170# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.8387e+08 ps=81280 
M1834 diff_1804670_2376170# diff_1795780_1543050# diff_580390_2383790# GND efet w=8890 l=7620
+ ad=2.96774e+08 pd=81280 as=0 ps=0 
M1835 diff_580390_2305050# diff_1765300_1584960# diff_1723390_2315210# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.80645e+08 ps=78740 
M1836 diff_1804670_2316480# diff_1795780_1543050# diff_580390_2305050# GND efet w=8890 l=7620
+ ad=2.8387e+08 pd=78740 as=0 ps=0 
M1837 diff_1685290_2282190# diff_1673860_1543050# diff_703580_2313940# GND efet w=22860 l=7620
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1838 GND diff_1658620_2316480# diff_1685290_2282190# GND efet w=26035 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1839 diff_1733550_2286000# diff_1723390_2315210# GND GND efet w=24130 l=7620
+ ad=2.64516e+08 pd=78740 as=0 ps=0 
M1840 diff_703580_2313940# diff_1728470_1526540# diff_1733550_2286000# GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1841 diff_1685290_2246630# diff_1673860_1543050# diff_703580_2232660# GND efet w=22860 l=7620
+ ad=2.66128e+08 pd=76200 as=0 ps=0 
M1842 diff_703580_2232660# diff_1728470_1526540# diff_1733550_2242820# GND efet w=25400 l=7620
+ ad=0 pd=0 as=2.77419e+08 ps=81280 
M1843 diff_580390_2232660# diff_1620520_1543050# diff_1577340_2226310# GND efet w=7620 l=7620
+ ad=0 pd=0 as=3.01612e+08 ps=81280 
M1844 diff_1658620_2226310# diff_1649730_1543050# diff_580390_2232660# GND efet w=7620 l=7620
+ ad=2.98386e+08 pd=78740 as=0 ps=0 
M1845 diff_580390_2155190# diff_1620520_1543050# diff_1577340_2164080# GND efet w=10160 l=7620
+ ad=0 pd=0 as=2.99999e+08 ps=78740 
M1846 diff_1658620_2166620# diff_1649730_1543050# diff_580390_2155190# GND efet w=8890 l=7620
+ ad=2.98386e+08 pd=78740 as=0 ps=0 
M1847 diff_703580_2164080# diff_1582420_1527810# diff_1588770_2136140# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1848 diff_1539240_2096770# diff_1527810_1543050# diff_703580_2081530# GND efet w=22225 l=8255
+ ad=2.93548e+08 pd=78740 as=0 ps=0 
M1849 diff_580390_2082800# diff_1474470_1583690# diff_1432560_2076450# GND efet w=10160 l=7620
+ ad=0 pd=0 as=3.06451e+08 ps=83820 
M1850 diff_1513840_2075180# diff_1504950_1543050# diff_580390_2082800# GND efet w=8890 l=7620
+ ad=3.06451e+08 pd=81280 as=0 ps=0 
M1851 diff_1394460_1981200# diff_1383030_1543050# diff_703580_2012950# GND efet w=22860 l=7620
+ ad=2.5e+08 pd=78740 as=0 ps=0 
M1852 GND diff_1367790_2015490# diff_1394460_1981200# GND efet w=26035 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1853 diff_1442720_1985010# diff_1432560_2014220# GND GND efet w=25400 l=7620
+ ad=2.75806e+08 pd=78740 as=0 ps=0 
M1854 diff_580390_2004060# diff_1474470_1583690# diff_1432560_2014220# GND efet w=10160 l=7620
+ ad=0 pd=0 as=2.99999e+08 ps=78740 
M1855 diff_1513840_2015490# diff_1504950_1543050# diff_580390_2004060# GND efet w=10160 l=7620
+ ad=2.91935e+08 pd=81280 as=0 ps=0 
M1856 diff_703580_2012950# diff_1436370_1529080# diff_1442720_1985010# GND efet w=22860 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1857 diff_1394460_1945640# diff_1383030_1543050# diff_703580_1931670# GND efet w=22860 l=7620
+ ad=2.66128e+08 pd=76200 as=0 ps=0 
M1858 diff_580390_1932940# diff_1329690_1543050# diff_1286510_1925320# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.98386e+08 ps=83820 
M1859 diff_1367790_1926590# diff_1358900_1543050# diff_580390_1932940# GND efet w=8890 l=7620
+ ad=2.87096e+08 pd=78740 as=0 ps=0 
M1860 diff_580390_1854200# diff_1329690_1543050# diff_1286510_1864360# GND efet w=9525 l=7620
+ ad=0 pd=0 as=2.91935e+08 ps=83820 
M1861 diff_1367790_1866900# diff_1358900_1543050# diff_580390_1854200# GND efet w=8890 l=7620
+ ad=2.69354e+08 pd=78740 as=0 ps=0 
M1862 diff_703580_1863090# diff_1291590_1526540# diff_1297940_1835150# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1863 diff_1249680_1793240# diff_1236980_1543050# diff_703580_1781810# GND efet w=22860 l=10160
+ ad=2.67741e+08 pd=76200 as=0 ps=0 
M1864 GND diff_1223010_1775460# diff_1249680_1793240# GND efet w=24765 l=9525
+ ad=0 pd=0 as=0 ps=0 
M1865 diff_580390_1783080# diff_1183640_1584960# diff_1141730_1775460# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.96774e+08 ps=78740 
M1866 diff_1223010_1775460# diff_1214120_1543050# diff_580390_1783080# GND efet w=8890 l=7620
+ ad=2.91935e+08 pd=78740 as=0 ps=0 
M1867 diff_1103630_1681480# diff_1092200_1543050# diff_703580_1714500# GND efet w=22860 l=7620
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1868 GND diff_1078230_1715770# diff_1103630_1681480# GND efet w=24130 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1869 diff_1151890_1685290# diff_1141730_1714500# GND GND efet w=24130 l=7620
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1870 diff_580390_1704340# diff_1183640_1584960# diff_1141730_1714500# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.98386e+08 ps=78740 
M1871 diff_1223010_1715770# diff_1214120_1543050# diff_580390_1704340# GND efet w=8890 l=7620
+ ad=2.85483e+08 pd=76200 as=0 ps=0 
M1872 diff_703580_1714500# diff_1145540_1527810# diff_1151890_1685290# GND efet w=22860 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1873 diff_1103630_1645920# diff_1092200_1543050# diff_703580_1633220# GND efet w=22860 l=7620
+ ad=2.7258e+08 pd=78740 as=0 ps=0 
M1874 diff_580390_1633220# diff_1038860_1543050# diff_995680_1626870# GND efet w=10160 l=8890
+ ad=0 pd=0 as=3.03225e+08 ps=83820 
M1875 diff_1078230_1617980# diff_1068070_1543050# diff_580390_1633220# GND efet w=9525 l=9525
+ ad=2.88709e+08 pd=78740 as=0 ps=0 
M1876 GND diff_1078230_1617980# diff_1103630_1645920# GND efet w=25400 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1877 diff_1151890_1640840# diff_1141730_1626870# GND GND efet w=25400 l=7620
+ ad=2.79032e+08 pd=83820 as=0 ps=0 
M1878 diff_703580_1633220# diff_1145540_1527810# diff_1151890_1640840# GND efet w=25400 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1879 diff_1297940_1790700# diff_1286510_1775460# GND GND efet w=25400 l=10160
+ ad=2.69354e+08 pd=78740 as=0 ps=0 
M1880 diff_703580_1781810# diff_1291590_1526540# diff_1297940_1790700# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1881 diff_1249680_1681480# diff_1236980_1543050# diff_703580_1714500# GND efet w=22860 l=8890
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1882 GND diff_1223010_1715770# diff_1249680_1681480# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1883 diff_1297940_1685290# diff_1286510_1714500# GND GND efet w=24130 l=8255
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1884 GND diff_1367790_1926590# diff_1394460_1945640# GND efet w=24765 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1885 diff_1442720_1941830# diff_1432560_1925320# GND GND efet w=24130 l=7620
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1886 diff_703580_1931670# diff_1436370_1529080# diff_1442720_1941830# GND efet w=22860 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1887 GND diff_1513840_2075180# diff_1539240_2096770# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1888 diff_1588770_2091690# diff_1577340_2076450# GND GND efet w=24130 l=8255
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1889 diff_703580_2081530# diff_1582420_1527810# diff_1588770_2091690# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1890 diff_1539240_1981200# diff_1527810_1543050# diff_703580_2012950# GND efet w=22860 l=7620
+ ad=3.04838e+08 pd=81280 as=0 ps=0 
M1891 GND diff_1513840_2015490# diff_1539240_1981200# GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1892 diff_1588770_1985010# diff_1577340_2014220# GND GND efet w=26035 l=8255
+ ad=2.70967e+08 pd=78740 as=0 ps=0 
M1893 GND diff_1658620_2226310# diff_1685290_2246630# GND efet w=24130 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1894 diff_1733550_2242820# diff_1723390_2226310# GND GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1895 GND diff_1658620_2166620# diff_1685290_2132330# GND efet w=25400 l=8255
+ ad=0 pd=0 as=2.66128e+08 ps=78740 
M1896 diff_1685290_2132330# diff_1673860_1543050# diff_703580_2164080# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1897 diff_1733550_2136140# diff_1723390_2164080# GND GND efet w=24130 l=7620
+ ad=2.95161e+08 pd=81280 as=0 ps=0 
M1898 GND diff_1804670_2376170# diff_1830070_2396490# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1899 diff_1879600_2391410# diff_1868170_2377440# GND GND efet w=24130 l=7620
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1900 diff_703580_2382520# diff_1873250_1527810# diff_1879600_2391410# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1901 diff_1830070_2284730# diff_1819910_1543050# diff_703580_2313940# GND efet w=24130 l=8255
+ ad=2.69354e+08 pd=81280 as=0 ps=0 
M1902 GND diff_1804670_2316480# diff_1830070_2284730# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1903 diff_1879600_2286000# diff_1868170_2316480# GND GND efet w=24130 l=7620
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1904 diff_2025650_2541270# diff_2014220_2526030# GND GND efet w=25400 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1905 diff_1976120_2432050# diff_1964690_1543050# diff_703580_2463800# GND efet w=22860 l=7620
+ ad=2.95161e+08 pd=81280 as=0 ps=0 
M1906 GND diff_1949450_2470150# diff_1976120_2432050# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1907 diff_2025650_2435860# diff_2014220_2465070# GND GND efet w=25400 l=7620
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1908 GND diff_2095500_2675890# diff_2122170_2697480# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1909 diff_2171700_2691130# diff_2160270_2675890# GND GND efet w=26035 l=8255
+ ad=2.67741e+08 pd=78740 as=0 ps=0 
M1910 diff_703580_2682240# diff_2165350_1529080# diff_2171700_2691130# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1911 diff_2122170_2581910# diff_2110740_1545590# diff_702310_2614930# GND efet w=22860 l=7620
+ ad=2.91935e+08 pd=81280 as=0 ps=0 
M1912 GND diff_2095500_2616200# diff_2122170_2581910# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1913 diff_2170430_2599690# diff_2160270_2614930# GND GND efet w=26670 l=8255
+ ad=2.62903e+08 pd=81280 as=0 ps=0 
M1914 Vdd diff_2002790_702310# diff_580390_2753360# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1915 diff_2268220_2731770# diff_2258060_1543050# diff_702310_2763520# GND efet w=22860 l=7620
+ ad=3.01612e+08 pd=81280 as=0 ps=0 
M1916 GND diff_2241550_2767330# diff_2268220_2731770# GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1917 Vdd diff_2354580_1676400# diff_702310_2763520# GND efet w=15240 l=6985
+ ad=0 pd=0 as=0 ps=0 
M1918 diff_2556510_3018790# Vdd Vdd GND efet w=11430 l=20320
+ ad=0 pd=0 as=0 ps=0 
M1919 Vdd Vdd Vdd GND efet w=5715 l=3175
+ ad=0 pd=0 as=0 ps=0 
M1920 Vdd Vdd Vdd GND efet w=4445 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1921 diff_2555240_2753360# Vdd Vdd GND efet w=13970 l=19685
+ ad=1.40484e+09 pd=276860 as=0 ps=0 
M1922 diff_2461260_2726690# clk2 diff_243840_2250440# GND efet w=20320 l=7620
+ ad=3.06451e+08 pd=81280 as=0 ps=0 
M1923 diff_2481580_2720340# diff_2195830_2933700# diff_2461260_2726690# GND efet w=20320 l=7620
+ ad=1.87258e+09 pd=345440 as=0 ps=0 
M1924 diff_2268220_2697480# diff_2258060_1543050# diff_703580_2682240# GND efet w=21590 l=7620
+ ad=2.35483e+08 pd=68580 as=0 ps=0 
M1925 GND diff_2241550_2675890# diff_2268220_2697480# GND efet w=17780 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1926 diff_580390_2682240# diff_2203450_1583690# diff_2160270_2675890# GND efet w=8890 l=8890
+ ad=0 pd=0 as=2.88709e+08 ps=78740 
M1927 diff_2241550_2675890# diff_2233930_1543050# diff_580390_2682240# GND efet w=8890 l=7620
+ ad=2.88709e+08 pd=81280 as=0 ps=0 
M1928 diff_580390_2603500# diff_2203450_1583690# diff_2160270_2614930# GND efet w=8255 l=9525
+ ad=0 pd=0 as=2.70967e+08 ps=91440 
M1929 diff_2241550_2616200# diff_2233930_1543050# diff_580390_2603500# GND efet w=8890 l=8890
+ ad=2.8387e+08 pd=78740 as=0 ps=0 
M1930 diff_702310_2614930# diff_2165350_1529080# diff_2170430_2599690# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1931 diff_2122170_2547620# diff_2110740_1545590# diff_703580_2532380# GND efet w=22225 l=8255
+ ad=2.82258e+08 pd=81280 as=0 ps=0 
M1932 diff_580390_2532380# diff_2057400_1583690# diff_2014220_2526030# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.95161e+08 ps=78740 
M1933 diff_2095500_2526030# diff_2087880_1543050# diff_580390_2532380# GND efet w=8890 l=7620
+ ad=2.93548e+08 pd=81280 as=0 ps=0 
M1934 diff_580390_2454910# diff_2057400_1583690# diff_2014220_2465070# GND efet w=9525 l=8255
+ ad=0 pd=0 as=2.99999e+08 ps=78740 
M1935 diff_2095500_2466340# diff_2087880_1543050# diff_580390_2454910# GND efet w=8890 l=7620
+ ad=2.93548e+08 pd=81280 as=0 ps=0 
M1936 diff_703580_2463800# diff_2019300_1526540# diff_2025650_2435860# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1937 diff_1976120_2397760# diff_1964690_1543050# diff_703580_2382520# GND efet w=21590 l=7620
+ ad=2.90322e+08 pd=78740 as=0 ps=0 
M1938 diff_580390_2383790# diff_1911350_1583690# diff_1868170_2377440# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.93548e+08 ps=81280 
M1939 diff_1949450_2382520# diff_1941830_1543050# diff_580390_2383790# GND efet w=10795 l=7620
+ ad=2.88709e+08 pd=83820 as=0 ps=0 
M1940 diff_580390_2305050# diff_1911350_1583690# diff_1868170_2316480# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.96774e+08 ps=78740 
M1941 diff_1950720_2316480# diff_1941830_1543050# diff_580390_2305050# GND efet w=8890 l=8890
+ ad=2.87096e+08 pd=81280 as=0 ps=0 
M1942 diff_703580_2313940# diff_1873250_1527810# diff_1879600_2286000# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1943 diff_1831340_2246630# diff_1819910_1543050# diff_703580_2232660# GND efet w=22860 l=8890
+ ad=2.7258e+08 pd=78740 as=0 ps=0 
M1944 diff_580390_2232660# diff_1765300_1584960# diff_1723390_2226310# GND efet w=8255 l=8255
+ ad=0 pd=0 as=2.8387e+08 ps=78740 
M1945 diff_1804670_2226310# diff_1795780_1543050# diff_580390_2232660# GND efet w=8890 l=8890
+ ad=2.85483e+08 pd=78740 as=0 ps=0 
M1946 GND diff_1804670_2226310# diff_1831340_2246630# GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1947 diff_1879600_2241550# diff_1868170_2232660# GND GND efet w=25400 l=7620
+ ad=2.69354e+08 pd=78740 as=0 ps=0 
M1948 diff_703580_2232660# diff_1873250_1527810# diff_1879600_2241550# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1949 diff_1804670_2166620# diff_1795780_1543050# diff_580390_2155190# GND efet w=10160 l=8890
+ ad=2.82258e+08 pd=78740 as=0 ps=0 
M1950 diff_580390_2155190# diff_1765300_1584960# diff_1723390_2164080# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.8387e+08 ps=78740 
M1951 diff_703580_2164080# diff_1728470_1526540# diff_1733550_2136140# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1952 diff_1685290_2096770# diff_1673860_1543050# diff_703580_2081530# GND efet w=21590 l=7620
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1953 diff_580390_2082800# diff_1620520_1543050# diff_1577340_2076450# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.90322e+08 ps=78740 
M1954 diff_1658620_2076450# diff_1649730_1543050# diff_580390_2082800# GND efet w=8890 l=7620
+ ad=2.91935e+08 pd=83820 as=0 ps=0 
M1955 diff_580390_2004060# diff_1620520_1543050# diff_1577340_2014220# GND efet w=9525 l=8255
+ ad=0 pd=0 as=2.99999e+08 ps=78740 
M1956 diff_1658620_2015490# diff_1649730_1543050# diff_580390_2004060# GND efet w=10160 l=7620
+ ad=3.03225e+08 pd=83820 as=0 ps=0 
M1957 diff_703580_2012950# diff_1582420_1527810# diff_1588770_1985010# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1958 diff_1539240_1946910# diff_1527810_1543050# diff_703580_1931670# GND efet w=22860 l=7620
+ ad=2.93548e+08 pd=78740 as=0 ps=0 
M1959 diff_580390_1932940# diff_1474470_1583690# diff_1432560_1925320# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.96774e+08 ps=78740 
M1960 diff_1513840_1925320# diff_1504950_1543050# diff_580390_1932940# GND efet w=8890 l=7620
+ ad=2.93548e+08 pd=78740 as=0 ps=0 
M1961 GND diff_1367790_1866900# diff_1394460_1831340# GND efet w=27305 l=8255
+ ad=0 pd=0 as=2.67741e+08 ps=78740 
M1962 diff_1394460_1831340# diff_1383030_1543050# diff_703580_1863090# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1963 diff_1442720_1835150# diff_1432560_1863090# GND GND efet w=24130 l=7620
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M1964 diff_580390_1854200# diff_1474470_1583690# diff_1432560_1863090# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.95161e+08 ps=78740 
M1965 diff_1513840_1866900# diff_1504950_1543050# diff_580390_1854200# GND efet w=8890 l=7620
+ ad=2.80645e+08 pd=78740 as=0 ps=0 
M1966 diff_703580_1863090# diff_1436370_1529080# diff_1442720_1835150# GND efet w=22860 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1967 diff_1394460_1795780# diff_1383030_1543050# diff_703580_1781810# GND efet w=21590 l=7620
+ ad=2.67741e+08 pd=78740 as=0 ps=0 
M1968 diff_580390_1783080# diff_1329690_1543050# diff_1286510_1775460# GND efet w=10160 l=8890
+ ad=0 pd=0 as=2.90322e+08 ps=83820 
M1969 diff_1367790_1775460# diff_1358900_1543050# diff_580390_1783080# GND efet w=8890 l=7620
+ ad=2.91935e+08 pd=81280 as=0 ps=0 
M1970 diff_580390_1704340# diff_1329690_1543050# diff_1286510_1714500# GND efet w=10795 l=8255
+ ad=0 pd=0 as=2.90322e+08 ps=88900 
M1971 diff_1367790_1715770# diff_1358900_1543050# diff_580390_1704340# GND efet w=8890 l=7620
+ ad=2.82258e+08 pd=83820 as=0 ps=0 
M1972 diff_703580_1714500# diff_1291590_1526540# diff_1297940_1685290# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1973 diff_1249680_1644650# diff_1236980_1543050# diff_703580_1633220# GND efet w=22860 l=8890
+ ad=2.70967e+08 pd=78740 as=0 ps=0 
M1974 diff_580390_1633220# diff_1183640_1584960# diff_1141730_1626870# GND efet w=9525 l=8255
+ ad=0 pd=0 as=3.01612e+08 ps=78740 
M1975 diff_1223010_1625600# diff_1214120_1543050# diff_580390_1633220# GND efet w=10160 l=7620
+ ad=2.87096e+08 pd=76200 as=0 ps=0 
M1976 GND diff_1223010_1625600# diff_1249680_1644650# GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1977 diff_1297940_1640840# diff_1286510_1626870# GND GND efet w=27305 l=8255
+ ad=2.66128e+08 pd=81280 as=0 ps=0 
M1978 diff_703580_1633220# diff_1291590_1526540# diff_1297940_1640840# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1979 GND diff_1367790_1775460# diff_1394460_1795780# GND efet w=24765 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1980 diff_1442720_1790700# diff_1432560_1775460# GND GND efet w=24130 l=7620
+ ad=2.66128e+08 pd=76200 as=0 ps=0 
M1981 diff_703580_1781810# diff_1436370_1529080# diff_1442720_1790700# GND efet w=21590 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1982 diff_1394460_1681480# diff_1383030_1543050# diff_703580_1714500# GND efet w=22860 l=7620
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M1983 GND diff_1367790_1715770# diff_1394460_1681480# GND efet w=25400 l=8255
+ ad=0 pd=0 as=0 ps=0 
M1984 diff_1442720_1685290# diff_1432560_1714500# GND GND efet w=24130 l=7620
+ ad=2.6129e+08 pd=76200 as=0 ps=0 
M1985 GND diff_1513840_1925320# diff_1539240_1946910# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1986 diff_1588770_1941830# diff_1577340_1925320# GND GND efet w=26670 l=8255
+ ad=2.6129e+08 pd=78740 as=0 ps=0 
M1987 diff_703580_1931670# diff_1582420_1527810# diff_1588770_1941830# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1988 diff_1539240_1831340# diff_1527810_1543050# diff_703580_1863090# GND efet w=24130 l=7620
+ ad=2.90322e+08 pd=81280 as=0 ps=0 
M1989 GND diff_1513840_1866900# diff_1539240_1831340# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1990 diff_1588770_1835150# diff_1577340_1864360# GND GND efet w=24130 l=8890
+ ad=2.6129e+08 pd=76200 as=0 ps=0 
M1991 GND diff_1658620_2076450# diff_1685290_2096770# GND efet w=24130 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1992 diff_1733550_2091690# diff_1723390_2076450# GND GND efet w=24130 l=7620
+ ad=2.87096e+08 pd=81280 as=0 ps=0 
M1993 diff_703580_2081530# diff_1728470_1526540# diff_1733550_2091690# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1994 diff_1685290_1981200# diff_1673860_1543050# diff_703580_2012950# GND efet w=22860 l=7620
+ ad=2.75806e+08 pd=78740 as=0 ps=0 
M1995 GND diff_1658620_2015490# diff_1685290_1981200# GND efet w=25400 l=8890
+ ad=0 pd=0 as=0 ps=0 
M1996 diff_1733550_1985010# diff_1723390_2014220# GND GND efet w=25400 l=7620
+ ad=3.01612e+08 pd=83820 as=0 ps=0 
M1997 diff_1831340_2132330# diff_1819910_1543050# diff_703580_2164080# GND efet w=22860 l=8890
+ ad=2.45161e+08 pd=76200 as=0 ps=0 
M1998 GND diff_1804670_2166620# diff_1831340_2132330# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M1999 diff_1879600_2136140# diff_1869440_2164080# GND GND efet w=24130 l=7620
+ ad=2.66128e+08 pd=78740 as=0 ps=0 
M2000 GND diff_1949450_2382520# diff_1976120_2397760# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2001 diff_2025650_2391410# diff_2014220_2377440# GND GND efet w=28575 l=8255
+ ad=2.67741e+08 pd=76200 as=0 ps=0 
M2002 diff_703580_2382520# diff_2019300_1526540# diff_2025650_2391410# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2003 diff_1976120_2282190# diff_1964690_1543050# diff_703580_2313940# GND efet w=22860 l=7620
+ ad=2.88709e+08 pd=81280 as=0 ps=0 
M2004 GND diff_1950720_2316480# diff_1976120_2282190# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2005 diff_2025650_2286000# diff_2014220_2315210# GND GND efet w=26670 l=7620
+ ad=2.59677e+08 pd=76200 as=0 ps=0 
M2006 GND diff_2095500_2526030# diff_2122170_2547620# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2007 diff_2171700_2542540# diff_2160270_2526030# GND GND efet w=23495 l=8255
+ ad=2.5e+08 pd=73660 as=0 ps=0 
M2008 diff_703580_2532380# diff_2165350_1529080# diff_2171700_2542540# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2009 diff_2122170_2432050# diff_2110740_1545590# diff_703580_2463800# GND efet w=22860 l=7620
+ ad=2.93548e+08 pd=81280 as=0 ps=0 
M2010 GND diff_2095500_2466340# diff_2122170_2432050# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2011 diff_2171700_2435860# diff_2160270_2465070# GND GND efet w=28575 l=8255
+ ad=2.59677e+08 pd=76200 as=0 ps=0 
M2012 Vdd diff_2354580_1676400# diff_703580_2682240# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2013 Vdd diff_2002790_702310# diff_580390_2682240# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2014 GND diff_2195830_2933700# diff_2565400_2665730# GND efet w=16510 l=6350
+ ad=0 pd=0 as=4.3387e+08 ps=88900 
M2015 GND diff_2198370_3069590# diff_2481580_2720340# GND efet w=29845 l=6985
+ ad=0 pd=0 as=0 ps=0 
M2016 diff_2565400_2665730# Vdd Vdd GND efet w=8890 l=60960
+ ad=0 pd=0 as=0 ps=0 
M2017 Vdd Vdd Vdd GND efet w=6350 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2018 diff_2481580_2720340# diff_2565400_2665730# diff_2598420_2640330# GND efet w=15240 l=7620
+ ad=0 pd=0 as=7.14515e+08 ps=147320 
M2019 diff_2555240_2753360# diff_2481580_2720340# GND GND efet w=118745 l=6985
+ ad=0 pd=0 as=0 ps=0 
M2020 Vdd Vdd Vdd GND efet w=4445 l=9525
+ ad=0 pd=0 as=0 ps=0 
M2021 diff_2598420_2640330# Vdd Vdd GND efet w=11430 l=29845
+ ad=0 pd=0 as=0 ps=0 
M2022 Vdd diff_2002790_702310# diff_580390_2603500# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2023 diff_2268220_2581910# diff_2258060_1543050# diff_702310_2614930# GND efet w=22860 l=7620
+ ad=2.91935e+08 pd=78740 as=0 ps=0 
M2024 GND diff_2241550_2616200# diff_2268220_2581910# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2025 Vdd diff_2354580_1676400# diff_702310_2614930# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2026 o2 diff_2513330_2576830# Vdd GND efet w=219075 l=6985
+ ad=9.05078e+07 pd=739140 as=0 ps=0 
M2027 diff_2268220_2547620# diff_2258060_1543050# diff_703580_2532380# GND efet w=22860 l=7620
+ ad=2.90322e+08 pd=81280 as=0 ps=0 
M2028 diff_580390_2532380# diff_2203450_1583690# diff_2160270_2526030# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.93548e+08 ps=78740 
M2029 diff_2241550_2526030# diff_2233930_1543050# diff_580390_2532380# GND efet w=8890 l=7620
+ ad=2.90322e+08 pd=81280 as=0 ps=0 
M2030 diff_580390_2454910# diff_2203450_1583690# diff_2160270_2465070# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.95161e+08 ps=78740 
M2031 diff_2241550_2466340# diff_2233930_1543050# diff_580390_2454910# GND efet w=8890 l=7620
+ ad=2.90322e+08 pd=81280 as=0 ps=0 
M2032 diff_703580_2463800# diff_2165350_1529080# diff_2171700_2435860# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2033 diff_2122170_2397760# diff_2110740_1545590# diff_703580_2382520# GND efet w=21590 l=7620
+ ad=2.91935e+08 pd=81280 as=0 ps=0 
M2034 diff_580390_2383790# diff_2057400_1583690# diff_2014220_2377440# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.98386e+08 ps=81280 
M2035 diff_2095500_2376170# diff_2087880_1543050# diff_580390_2383790# GND efet w=8890 l=7620
+ ad=2.88709e+08 pd=81280 as=0 ps=0 
M2036 diff_580390_2305050# diff_2057400_1583690# diff_2014220_2315210# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.95161e+08 ps=78740 
M2037 diff_2095500_2317750# diff_2087880_1543050# diff_580390_2305050# GND efet w=7620 l=7620
+ ad=2.91935e+08 pd=81280 as=0 ps=0 
M2038 diff_703580_2313940# diff_2019300_1526540# diff_2025650_2286000# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2039 diff_1976120_2247900# diff_1964690_1543050# diff_703580_2232660# GND efet w=22860 l=7620
+ ad=2.91935e+08 pd=78740 as=0 ps=0 
M2040 diff_580390_2232660# diff_1911350_1583690# diff_1868170_2232660# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.96774e+08 ps=83820 
M2041 diff_1950720_2226310# diff_1941830_1543050# diff_580390_2232660# GND efet w=9525 l=8890
+ ad=2.91935e+08 pd=81280 as=0 ps=0 
M2042 diff_580390_2155190# diff_1911350_1583690# diff_1869440_2164080# GND efet w=10160 l=7620
+ ad=0 pd=0 as=3.03225e+08 ps=81280 
M2043 diff_1950720_2166620# diff_1941830_1543050# diff_580390_2155190# GND efet w=10160 l=7620
+ ad=2.93548e+08 pd=81280 as=0 ps=0 
M2044 diff_703580_2164080# diff_1873250_1527810# diff_1879600_2136140# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2045 diff_1831340_2096770# diff_1819910_1543050# diff_703580_2081530# GND efet w=22225 l=9525
+ ad=2.66128e+08 pd=78740 as=0 ps=0 
M2046 diff_580390_2082800# diff_1765300_1584960# diff_1723390_2076450# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.69354e+08 ps=78740 
M2047 diff_1804670_2076450# diff_1795780_1543050# diff_580390_2082800# GND efet w=8890 l=7620
+ ad=2.67741e+08 pd=78740 as=0 ps=0 
M2048 diff_580390_2004060# diff_1765300_1584960# diff_1723390_2014220# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.82258e+08 ps=78740 
M2049 diff_1804670_2015490# diff_1795780_1543050# diff_580390_2004060# GND efet w=8890 l=7620
+ ad=2.98386e+08 pd=83820 as=0 ps=0 
M2050 diff_703580_2012950# diff_1728470_1526540# diff_1733550_1985010# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2051 diff_1685290_1945640# diff_1673860_1543050# diff_703580_1931670# GND efet w=22860 l=7620
+ ad=2.69354e+08 pd=78740 as=0 ps=0 
M2052 diff_703580_1931670# diff_1728470_1526540# diff_1733550_1940560# GND efet w=28575 l=7620
+ ad=0 pd=0 as=2.87096e+08 ps=91440 
M2053 diff_580390_1932940# diff_1620520_1543050# diff_1577340_1925320# GND efet w=9525 l=8255
+ ad=0 pd=0 as=2.98386e+08 ps=78740 
M2054 diff_1658620_1925320# diff_1649730_1543050# diff_580390_1932940# GND efet w=10160 l=8890
+ ad=2.98386e+08 pd=78740 as=0 ps=0 
M2055 diff_580390_1854200# diff_1620520_1543050# diff_1577340_1864360# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.93548e+08 ps=78740 
M2056 diff_1658620_1866900# diff_1649730_1543050# diff_580390_1854200# GND efet w=8890 l=7620
+ ad=2.96774e+08 pd=78740 as=0 ps=0 
M2057 diff_703580_1863090# diff_1582420_1527810# diff_1588770_1835150# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2058 diff_1539240_1795780# diff_1527810_1543050# diff_703580_1781810# GND efet w=21590 l=7620
+ ad=2.93548e+08 pd=78740 as=0 ps=0 
M2059 diff_580390_1783080# diff_1474470_1583690# diff_1432560_1775460# GND efet w=8890 l=7620
+ ad=0 pd=0 as=3.01612e+08 ps=81280 
M2060 diff_1513840_1775460# diff_1504950_1543050# diff_580390_1783080# GND efet w=9525 l=8255
+ ad=2.8387e+08 pd=76200 as=0 ps=0 
M2061 diff_580390_1704340# diff_1474470_1583690# diff_1432560_1714500# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.96774e+08 ps=78740 
M2062 diff_1513840_1715770# diff_1504950_1543050# diff_580390_1704340# GND efet w=8890 l=7620
+ ad=2.8387e+08 pd=76200 as=0 ps=0 
M2063 diff_703580_1714500# diff_1436370_1529080# diff_1442720_1685290# GND efet w=22860 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2064 diff_1394460_1645920# diff_1383030_1543050# diff_703580_1633220# GND efet w=22860 l=7620
+ ad=2.64516e+08 pd=78740 as=0 ps=0 
M2065 diff_580390_1633220# diff_1329690_1543050# diff_1286510_1626870# GND efet w=8890 l=7620
+ ad=0 pd=0 as=3.01612e+08 ps=83820 
M2066 diff_1367790_1625600# diff_1358900_1543050# diff_580390_1633220# GND efet w=8890 l=7620
+ ad=2.88709e+08 pd=81280 as=0 ps=0 
M2067 GND diff_1367790_1625600# diff_1394460_1645920# GND efet w=24130 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2068 diff_1442720_1642110# diff_1432560_1626870# GND GND efet w=24130 l=7620
+ ad=2.59677e+08 pd=76200 as=0 ps=0 
M2069 diff_703580_1633220# diff_1436370_1529080# diff_1442720_1642110# GND efet w=22860 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2070 GND diff_1513840_1775460# diff_1539240_1795780# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2071 diff_1588770_1790700# diff_1577340_1775460# GND GND efet w=24130 l=8890
+ ad=2.6129e+08 pd=78740 as=0 ps=0 
M2072 diff_703580_1781810# diff_1582420_1527810# diff_1588770_1790700# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2073 diff_1539240_1681480# diff_1527810_1543050# diff_703580_1714500# GND efet w=22860 l=7620
+ ad=2.93548e+08 pd=78740 as=0 ps=0 
M2074 GND diff_1513840_1715770# diff_1539240_1681480# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2075 diff_1588770_1685290# diff_1577340_1714500# GND GND efet w=24130 l=8890
+ ad=2.6129e+08 pd=76200 as=0 ps=0 
M2076 GND diff_1658620_1925320# diff_1685290_1945640# GND efet w=24765 l=9525
+ ad=0 pd=0 as=0 ps=0 
M2077 diff_1733550_1940560# diff_1723390_1925320# GND GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2078 GND diff_1804670_2076450# diff_1831340_2096770# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2079 diff_1879600_2091690# diff_1869440_2075180# GND GND efet w=24130 l=7620
+ ad=2.64516e+08 pd=78740 as=0 ps=0 
M2080 diff_703580_2081530# diff_1873250_1527810# diff_1879600_2091690# GND efet w=22225 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2081 diff_1831340_1981200# diff_1819910_1543050# diff_703580_2012950# GND efet w=22860 l=8890
+ ad=2.74193e+08 pd=78740 as=0 ps=0 
M2082 GND diff_1804670_2015490# diff_1831340_1981200# GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2083 diff_1879600_1985010# diff_1868170_2015490# GND GND efet w=25400 l=7620
+ ad=2.75806e+08 pd=78740 as=0 ps=0 
M2084 GND diff_1950720_2226310# diff_1976120_2247900# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2085 diff_2025650_2242820# diff_2014220_2226310# GND GND efet w=24130 l=7620
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M2086 diff_703580_2232660# diff_2019300_1526540# diff_2025650_2242820# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2087 diff_1976120_2132330# diff_1964690_1543050# diff_703580_2164080# GND efet w=22860 l=7620
+ ad=2.93548e+08 pd=81280 as=0 ps=0 
M2088 GND diff_1950720_2166620# diff_1976120_2132330# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2089 diff_2025650_2136140# diff_2014220_2164080# GND GND efet w=24130 l=7620
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M2090 diff_580390_2232660# diff_2057400_1583690# diff_2014220_2226310# GND efet w=7620 l=7620
+ ad=0 pd=0 as=3.01612e+08 ps=81280 
M2091 GND diff_2095500_2376170# diff_2122170_2397760# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2092 diff_2171700_2391410# diff_2160270_2377440# GND GND efet w=26035 l=8255
+ ad=2.59677e+08 pd=76200 as=0 ps=0 
M2093 diff_703580_2382520# diff_2165350_1529080# diff_2171700_2391410# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2094 diff_2122170_2283460# diff_2110740_1545590# diff_703580_2313940# GND efet w=21590 l=7620
+ ad=2.85483e+08 pd=78740 as=0 ps=0 
M2095 GND diff_2095500_2317750# diff_2122170_2283460# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2096 diff_2171700_2286000# diff_2160270_2315210# GND GND efet w=24130 l=8255
+ ad=2.51612e+08 pd=73660 as=0 ps=0 
M2097 GND diff_2241550_2526030# diff_2268220_2547620# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2098 diff_2598420_2640330# diff_2555240_2753360# GND GND efet w=26670 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2099 o2 diff_2555240_2753360# GND GND efet w=208280 l=6350
+ ad=0 pd=0 as=0 ps=0 
M2100 Vdd diff_2354580_1676400# diff_703580_2532380# GND efet w=15240 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2101 Vdd diff_2002790_702310# diff_580390_2532380# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2102 diff_2513330_2576830# diff_2513330_2576830# diff_2513330_2576830# GND efet w=1905 l=3810
+ ad=1.09838e+09 pd=177800 as=0 ps=0 
M2103 diff_2513330_2576830# diff_2513330_2576830# diff_2513330_2576830# GND efet w=2540 l=2540
+ ad=0 pd=0 as=0 ps=0 
M2104 diff_2513330_2576830# Vdd Vdd GND efet w=11430 l=20320
+ ad=0 pd=0 as=0 ps=0 
M2105 GND diff_2555240_2753360# diff_2513330_2576830# GND efet w=52705 l=6985
+ ad=0 pd=0 as=0 ps=0 
M2106 Vdd diff_2002790_702310# diff_580390_2454910# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2107 diff_2268220_2432050# diff_2258060_1543050# diff_703580_2463800# GND efet w=22860 l=7620
+ ad=2.93548e+08 pd=81280 as=0 ps=0 
M2108 GND diff_2241550_2466340# diff_2268220_2432050# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2109 Vdd diff_2354580_1676400# diff_703580_2463800# GND efet w=15240 l=6985
+ ad=0 pd=0 as=0 ps=0 
M2110 diff_2268220_2397760# diff_2258060_1543050# diff_703580_2382520# GND efet w=21590 l=7620
+ ad=2.82258e+08 pd=81280 as=0 ps=0 
M2111 diff_580390_2383790# diff_2203450_1583690# diff_2160270_2377440# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.91935e+08 ps=78740 
M2112 diff_2241550_2376170# diff_2233930_1543050# diff_580390_2383790# GND efet w=8890 l=7620
+ ad=2.88709e+08 pd=78740 as=0 ps=0 
M2113 diff_580390_2305050# diff_2203450_1583690# diff_2160270_2315210# GND efet w=7620 l=7620
+ ad=0 pd=0 as=2.93548e+08 ps=78740 
M2114 diff_2241550_2317750# diff_2233930_1543050# diff_580390_2305050# GND efet w=7620 l=7620
+ ad=2.87096e+08 pd=81280 as=0 ps=0 
M2115 diff_703580_2313940# diff_2165350_1529080# diff_2171700_2286000# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2116 diff_2122170_2247900# diff_2110740_1545590# diff_703580_2232660# GND efet w=22860 l=7620
+ ad=2.90322e+08 pd=78740 as=0 ps=0 
M2117 diff_2095500_2227580# diff_2087880_1543050# diff_580390_2232660# GND efet w=7620 l=7620
+ ad=2.96774e+08 pd=83820 as=0 ps=0 
M2118 diff_580390_2155190# diff_2057400_1583690# diff_2014220_2164080# GND efet w=10160 l=7620
+ ad=0 pd=0 as=3.04838e+08 ps=81280 
M2119 diff_2095500_2166620# diff_2087880_1543050# diff_580390_2155190# GND efet w=8890 l=7620
+ ad=2.88709e+08 pd=78740 as=0 ps=0 
M2120 diff_703580_2164080# diff_2019300_1526540# diff_2025650_2136140# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2121 diff_1976120_2098040# diff_1964690_1543050# diff_703580_2081530# GND efet w=21590 l=7620
+ ad=2.93548e+08 pd=81280 as=0 ps=0 
M2122 diff_580390_2082800# diff_1911350_1583690# diff_1869440_2075180# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.90322e+08 ps=86360 
M2123 diff_1950720_2076450# diff_1941830_1543050# diff_580390_2082800# GND efet w=8890 l=7620
+ ad=2.77419e+08 pd=83820 as=0 ps=0 
M2124 diff_580390_2004060# diff_1911350_1583690# diff_1868170_2015490# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.85483e+08 ps=83820 
M2125 diff_1950720_2016760# diff_1941830_1543050# diff_580390_2004060# GND efet w=10795 l=8255
+ ad=2.85483e+08 pd=83820 as=0 ps=0 
M2126 diff_703580_2012950# diff_1873250_1527810# diff_1879600_1985010# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2127 diff_1831340_1945640# diff_1819910_1543050# diff_703580_1931670# GND efet w=22860 l=8890
+ ad=2.70967e+08 pd=78740 as=0 ps=0 
M2128 diff_580390_1932940# diff_1765300_1584960# diff_1723390_1925320# GND efet w=10160 l=7620
+ ad=0 pd=0 as=2.87096e+08 ps=78740 
M2129 diff_1804670_1925320# diff_1795780_1543050# diff_580390_1932940# GND efet w=10160 l=7620
+ ad=2.90322e+08 pd=81280 as=0 ps=0 
M2130 GND diff_1804670_1925320# diff_1831340_1945640# GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2131 diff_1879600_1940560# diff_1868170_1929130# GND GND efet w=25400 l=7620
+ ad=2.70967e+08 pd=78740 as=0 ps=0 
M2132 diff_703580_1931670# diff_1873250_1527810# diff_1879600_1940560# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2133 diff_580390_1854200# diff_1765300_1584960# diff_1723390_1863090# GND efet w=7620 l=8255
+ ad=0 pd=0 as=2.8387e+08 ps=81280 
M2134 diff_1804670_1866900# diff_1795780_1543050# diff_580390_1854200# GND efet w=8255 l=8255
+ ad=2.87096e+08 pd=81280 as=0 ps=0 
M2135 diff_1685290_1831340# diff_1673860_1543050# diff_703580_1863090# GND efet w=22860 l=7620
+ ad=2.66128e+08 pd=78740 as=0 ps=0 
M2136 GND diff_1658620_1866900# diff_1685290_1831340# GND efet w=24130 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2137 diff_1733550_1835150# diff_1723390_1863090# GND GND efet w=24130 l=7620
+ ad=2.74193e+08 pd=86360 as=0 ps=0 
M2138 diff_703580_1863090# diff_1728470_1526540# diff_1733550_1835150# GND efet w=26035 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2139 diff_1685290_1795780# diff_1673860_1543050# diff_703580_1781810# GND efet w=21590 l=7620
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M2140 diff_580390_1783080# diff_1620520_1543050# diff_1577340_1775460# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.95161e+08 ps=78740 
M2141 diff_1658620_1775460# diff_1649730_1543050# diff_580390_1783080# GND efet w=8890 l=7620
+ ad=2.98386e+08 pd=78740 as=0 ps=0 
M2142 diff_580390_1704340# diff_1620520_1543050# diff_1577340_1714500# GND efet w=8890 l=8890
+ ad=0 pd=0 as=2.96774e+08 ps=83820 
M2143 diff_1658620_1715770# diff_1649730_1543050# diff_580390_1704340# GND efet w=8890 l=7620
+ ad=2.82258e+08 pd=78740 as=0 ps=0 
M2144 diff_703580_1714500# diff_1582420_1527810# diff_1588770_1685290# GND efet w=22225 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2145 diff_1539240_1647190# diff_1527810_1543050# diff_703580_1633220# GND efet w=25400 l=8890
+ ad=2.85483e+08 pd=83820 as=0 ps=0 
M2146 diff_580390_1633220# diff_1474470_1583690# diff_1432560_1626870# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.98386e+08 ps=78740 
M2147 diff_1513840_1625600# diff_1504950_1543050# diff_580390_1633220# GND efet w=8890 l=7620
+ ad=2.8387e+08 pd=76200 as=0 ps=0 
M2148 GND diff_1513840_1625600# diff_1539240_1647190# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2149 diff_1588770_1642110# diff_1577340_1626870# GND GND efet w=22860 l=8890
+ ad=2.59677e+08 pd=81280 as=0 ps=0 
M2150 diff_703580_1633220# diff_1582420_1527810# diff_1588770_1642110# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2151 GND diff_1658620_1775460# diff_1685290_1795780# GND efet w=24130 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2152 diff_1733550_1790700# diff_1723390_1775460# GND GND efet w=24130 l=7620
+ ad=2.64516e+08 pd=78740 as=0 ps=0 
M2153 diff_703580_1781810# diff_1728470_1526540# diff_1733550_1790700# GND efet w=21590 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2154 diff_1831340_1831340# diff_1819910_1543050# diff_703580_1863090# GND efet w=22860 l=8890
+ ad=2.46774e+08 pd=78740 as=0 ps=0 
M2155 GND diff_1804670_1866900# diff_1831340_1831340# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2156 diff_1879600_1835150# diff_1868170_1865630# GND GND efet w=24130 l=7620
+ ad=2.66128e+08 pd=78740 as=0 ps=0 
M2157 GND diff_1950720_2076450# diff_1976120_2098040# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2158 diff_2025650_2091690# diff_2014220_2076450# GND GND efet w=24130 l=7620
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M2159 diff_703580_2081530# diff_2019300_1526540# diff_2025650_2091690# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2160 diff_1976120_1981200# diff_1964690_1543050# diff_703580_2012950# GND efet w=22860 l=7620
+ ad=3.01612e+08 pd=81280 as=0 ps=0 
M2161 GND diff_1950720_2016760# diff_1976120_1981200# GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2162 diff_2025650_1985010# diff_2014220_2014220# GND GND efet w=25400 l=7620
+ ad=2.74193e+08 pd=78740 as=0 ps=0 
M2163 GND diff_2095500_2227580# diff_2122170_2247900# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2164 diff_2171700_2242820# diff_2160270_2226310# GND GND efet w=27305 l=8255
+ ad=2.59677e+08 pd=76200 as=0 ps=0 
M2165 diff_703580_2232660# diff_2165350_1529080# diff_2171700_2242820# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2166 diff_2122170_2132330# diff_2110740_1545590# diff_703580_2164080# GND efet w=22860 l=7620
+ ad=2.93548e+08 pd=81280 as=0 ps=0 
M2167 GND diff_2095500_2166620# diff_2122170_2132330# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2168 diff_2171700_2136140# diff_2160270_2164080# GND GND efet w=24765 l=8255
+ ad=2.59677e+08 pd=76200 as=0 ps=0 
M2169 GND diff_2241550_2376170# diff_2268220_2397760# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2170 Vdd diff_2354580_1676400# diff_703580_2382520# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2171 Vdd diff_2002790_702310# diff_580390_2383790# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2172 Vdd diff_2002790_702310# diff_580390_2305050# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2173 GND diff_2241550_2317750# diff_2268220_2283460# GND efet w=23495 l=8255
+ ad=0 pd=0 as=2.82258e+08 ps=78740 
M2174 diff_2268220_2283460# diff_2258060_1543050# diff_703580_2313940# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2175 Vdd diff_2354580_1676400# diff_703580_2313940# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2176 diff_2557780_2068830# Vdd Vdd GND efet w=11430 l=20320
+ ad=1.47419e+09 pd=276860 as=0 ps=0 
M2177 diff_2461260_2273300# clk2 diff_245110_1436370# GND efet w=20320 l=7620
+ ad=3.01612e+08 pd=81280 as=0 ps=0 
M2178 diff_2268220_2247900# diff_2258060_1543050# diff_703580_2232660# GND efet w=22860 l=7620
+ ad=2.91935e+08 pd=78740 as=0 ps=0 
M2179 diff_580390_2232660# diff_2203450_1583690# diff_2160270_2226310# GND efet w=7620 l=7620
+ ad=0 pd=0 as=2.90322e+08 ps=78740 
M2180 diff_2241550_2227580# diff_2233930_1543050# diff_580390_2232660# GND efet w=7620 l=7620
+ ad=2.90322e+08 pd=81280 as=0 ps=0 
M2181 diff_580390_2155190# diff_2203450_1583690# diff_2160270_2164080# GND efet w=8890 l=8890
+ ad=0 pd=0 as=2.90322e+08 ps=78740 
M2182 diff_2241550_2167890# diff_2233930_1543050# diff_580390_2155190# GND efet w=7620 l=7620
+ ad=2.91935e+08 pd=81280 as=0 ps=0 
M2183 diff_703580_2164080# diff_2165350_1529080# diff_2171700_2136140# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2184 diff_2122170_2098040# diff_2110740_1545590# diff_703580_2081530# GND efet w=21590 l=7620
+ ad=2.90322e+08 pd=78740 as=0 ps=0 
M2185 diff_580390_2082800# diff_2057400_1583690# diff_2014220_2076450# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.87096e+08 ps=81280 
M2186 diff_2095500_2076450# diff_2087880_1543050# diff_580390_2082800# GND efet w=8890 l=7620
+ ad=2.90322e+08 pd=81280 as=0 ps=0 
M2187 diff_580390_2004060# diff_2057400_1583690# diff_2014220_2014220# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.98386e+08 ps=81280 
M2188 diff_2095500_2016760# diff_2087880_1543050# diff_580390_2004060# GND efet w=8890 l=7620
+ ad=2.93548e+08 pd=83820 as=0 ps=0 
M2189 diff_703580_2012950# diff_2019300_1526540# diff_2025650_1985010# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2190 diff_1976120_1946910# diff_1964690_1543050# diff_703580_1931670# GND efet w=22860 l=7620
+ ad=2.95161e+08 pd=78740 as=0 ps=0 
M2191 diff_580390_1932940# diff_1911350_1583690# diff_1868170_1929130# GND efet w=10160 l=7620
+ ad=0 pd=0 as=2.96774e+08 ps=83820 
M2192 diff_1950720_1925320# diff_1941830_1543050# diff_580390_1932940# GND efet w=12065 l=8255
+ ad=2.88709e+08 pd=81280 as=0 ps=0 
M2193 diff_580390_1854200# diff_1911350_1583690# diff_1868170_1865630# GND efet w=8890 l=7620
+ ad=0 pd=0 as=3.03225e+08 ps=81280 
M2194 diff_1950720_1865630# diff_1941830_1543050# diff_580390_1854200# GND efet w=8890 l=8890
+ ad=2.93548e+08 pd=81280 as=0 ps=0 
M2195 diff_703580_1863090# diff_1873250_1527810# diff_1879600_1835150# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2196 diff_1831340_1795780# diff_1819910_1543050# diff_703580_1781810# GND efet w=21590 l=8890
+ ad=2.64516e+08 pd=78740 as=0 ps=0 
M2197 diff_703580_1781810# diff_1873250_1527810# diff_1879600_1790700# GND efet w=22860 l=8890
+ ad=0 pd=0 as=2.66128e+08 ps=76200 
M2198 diff_580390_1783080# diff_1765300_1584960# diff_1723390_1775460# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.8387e+08 ps=81280 
M2199 diff_1804670_1775460# diff_1795780_1543050# diff_580390_1783080# GND efet w=8890 l=7620
+ ad=2.85483e+08 pd=78740 as=0 ps=0 
M2200 diff_1685290_1681480# diff_1673860_1543050# diff_703580_1714500# GND efet w=22225 l=8255
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M2201 GND diff_1658620_1715770# diff_1685290_1681480# GND efet w=24130 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2202 diff_1733550_1685290# diff_1723390_1714500# GND GND efet w=24130 l=7620
+ ad=2.67741e+08 pd=78740 as=0 ps=0 
M2203 GND diff_1804670_1775460# diff_1831340_1795780# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2204 diff_1879600_1790700# diff_1868170_1776730# GND GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2205 diff_580390_1704340# diff_1765300_1584960# diff_1723390_1714500# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.80645e+08 ps=78740 
M2206 diff_1804670_1715770# diff_1795780_1543050# diff_580390_1704340# GND efet w=8890 l=7620
+ ad=2.7258e+08 pd=81280 as=0 ps=0 
M2207 diff_703580_1714500# diff_1728470_1526540# diff_1733550_1685290# GND efet w=23495 l=9525
+ ad=0 pd=0 as=0 ps=0 
M2208 diff_1685290_1645920# diff_1673860_1543050# diff_703580_1633220# GND efet w=21590 l=7620
+ ad=2.62903e+08 pd=78740 as=0 ps=0 
M2209 diff_703580_1633220# diff_1728470_1526540# diff_1733550_1640840# GND efet w=22225 l=8255
+ ad=0 pd=0 as=2.67741e+08 ps=81280 
M2210 diff_580390_1633220# diff_1620520_1543050# diff_1577340_1626870# GND efet w=10160 l=7620
+ ad=0 pd=0 as=3.04838e+08 ps=83820 
M2211 diff_1658620_1625600# diff_1649730_1543050# diff_580390_1633220# GND efet w=10160 l=7620
+ ad=2.99999e+08 pd=78740 as=0 ps=0 
M2212 GND diff_1658620_1625600# diff_1685290_1645920# GND efet w=24130 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2213 diff_1733550_1640840# diff_1723390_1626870# GND GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2214 diff_1831340_1681480# diff_1819910_1543050# diff_703580_1714500# GND efet w=22225 l=9525
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M2215 GND diff_1804670_1715770# diff_1831340_1681480# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2216 diff_1879600_1685290# diff_1868170_1715770# GND GND efet w=24130 l=7620
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M2217 GND diff_1950720_1925320# diff_1976120_1946910# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2218 diff_2025650_1941830# diff_2014220_1926590# GND GND efet w=24130 l=7620
+ ad=2.64516e+08 pd=76200 as=0 ps=0 
M2219 diff_703580_1931670# diff_2019300_1526540# diff_2025650_1941830# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2220 diff_1976120_1831340# diff_1964690_1543050# diff_703580_1863090# GND efet w=22860 l=7620
+ ad=2.95161e+08 pd=81280 as=0 ps=0 
M2221 GND diff_1950720_1865630# diff_1976120_1831340# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2222 diff_2025650_1835150# diff_2014220_1864360# GND GND efet w=24130 l=7620
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M2223 GND diff_2095500_2076450# diff_2122170_2098040# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2224 diff_2171700_2091690# diff_2160270_2076450# GND GND efet w=24130 l=7620
+ ad=2.6129e+08 pd=78740 as=0 ps=0 
M2225 diff_703580_2081530# diff_2165350_1529080# diff_2171700_2091690# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2226 diff_2122170_1982470# diff_2110740_1545590# diff_703580_2012950# GND efet w=21590 l=7620
+ ad=2.93548e+08 pd=78740 as=0 ps=0 
M2227 GND diff_2095500_2016760# diff_2122170_1982470# GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2228 diff_2171700_1985010# diff_2160270_2014220# GND GND efet w=24130 l=7620
+ ad=2.51612e+08 pd=73660 as=0 ps=0 
M2229 GND diff_2241550_2227580# diff_2268220_2247900# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2230 diff_2481580_2265680# diff_2195830_2933700# diff_2461260_2273300# GND efet w=20320 l=7620
+ ad=1.89838e+09 pd=355600 as=0 ps=0 
M2231 Vdd diff_2354580_1676400# diff_703580_2232660# GND efet w=16510 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2232 GND diff_2195830_2933700# diff_2566670_2211070# GND efet w=15240 l=6985
+ ad=0 pd=0 as=3.88709e+08 ps=83820 
M2233 GND diff_2198370_3069590# diff_2481580_2265680# GND efet w=29210 l=6350
+ ad=0 pd=0 as=0 ps=0 
M2234 Vdd diff_2002790_702310# diff_580390_2232660# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2235 diff_2566670_2211070# Vdd Vdd GND efet w=9525 l=61595
+ ad=0 pd=0 as=0 ps=0 
M2236 Vdd Vdd Vdd GND efet w=6350 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2237 Vdd diff_2002790_702310# diff_580390_2155190# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2238 diff_2481580_2265680# diff_2566670_2211070# diff_2598420_2186940# GND efet w=15240 l=6350
+ ad=0 pd=0 as=7.38708e+08 ps=154940 
M2239 diff_2557780_2068830# diff_2481580_2265680# GND GND efet w=118110 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2240 Vdd Vdd Vdd GND efet w=5080 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2241 diff_2598420_2186940# Vdd Vdd GND efet w=10160 l=32385
+ ad=0 pd=0 as=0 ps=0 
M2242 diff_2268220_2132330# diff_2258060_1543050# diff_703580_2164080# GND efet w=22860 l=7620
+ ad=2.93548e+08 pd=81280 as=0 ps=0 
M2243 GND diff_2241550_2167890# diff_2268220_2132330# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2244 Vdd diff_2354580_1676400# diff_703580_2164080# GND efet w=16510 l=6350
+ ad=0 pd=0 as=0 ps=0 
M2245 diff_2268220_2098040# diff_2258060_1543050# diff_703580_2081530# GND efet w=21590 l=7620
+ ad=2.90322e+08 pd=81280 as=0 ps=0 
M2246 diff_580390_2082800# diff_2203450_1583690# diff_2160270_2076450# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.82258e+08 ps=78740 
M2247 diff_2241550_2076450# diff_2233930_1543050# diff_580390_2082800# GND efet w=8890 l=7620
+ ad=2.82258e+08 pd=83820 as=0 ps=0 
M2248 diff_580390_2004060# diff_2203450_1583690# diff_2160270_2014220# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.87096e+08 ps=78740 
M2249 diff_2241550_2016760# diff_2233930_1543050# diff_580390_2004060# GND efet w=8890 l=7620
+ ad=2.8387e+08 pd=81280 as=0 ps=0 
M2250 diff_703580_2012950# diff_2165350_1529080# diff_2171700_1985010# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2251 diff_2122170_1946910# diff_2110740_1545590# diff_703580_1931670# GND efet w=22860 l=7620
+ ad=2.91935e+08 pd=78740 as=0 ps=0 
M2252 diff_580390_1932940# diff_2057400_1583690# diff_2014220_1926590# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.98386e+08 ps=78740 
M2253 diff_2095500_1926590# diff_2087880_1543050# diff_580390_1932940# GND efet w=10160 l=7620
+ ad=2.77419e+08 pd=81280 as=0 ps=0 
M2254 diff_580390_1854200# diff_2057400_1583690# diff_2014220_1864360# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.93548e+08 ps=78740 
M2255 diff_2095500_1866900# diff_2087880_1543050# diff_580390_1854200# GND efet w=8890 l=7620
+ ad=2.87096e+08 pd=81280 as=0 ps=0 
M2256 diff_703580_1863090# diff_2019300_1526540# diff_2025650_1835150# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2257 diff_1976120_1797050# diff_1964690_1543050# diff_703580_1781810# GND efet w=21590 l=7620
+ ad=2.93548e+08 pd=81280 as=0 ps=0 
M2258 diff_580390_1783080# diff_1911350_1583690# diff_1868170_1776730# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.98386e+08 ps=78740 
M2259 diff_1950720_1775460# diff_1941830_1543050# diff_580390_1783080# GND efet w=8890 l=8890
+ ad=2.87096e+08 pd=81280 as=0 ps=0 
M2260 diff_580390_1704340# diff_1911350_1583690# diff_1868170_1715770# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.96774e+08 ps=78740 
M2261 diff_1950720_1715770# diff_1941830_1543050# diff_580390_1704340# GND efet w=8890 l=8890
+ ad=2.79032e+08 pd=83820 as=0 ps=0 
M2262 diff_703580_1714500# diff_1873250_1527810# diff_1879600_1685290# GND efet w=22225 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2263 diff_1831340_1645920# diff_1819910_1543050# diff_703580_1633220# GND efet w=21590 l=8890
+ ad=2.64516e+08 pd=78740 as=0 ps=0 
M2264 diff_703580_1633220# diff_1873250_1527810# diff_1879600_1640840# GND efet w=21590 l=8890
+ ad=0 pd=0 as=2.66128e+08 ps=76200 
M2265 diff_580390_1633220# diff_1765300_1584960# diff_1723390_1626870# GND efet w=10160 l=7620
+ ad=0 pd=0 as=2.85483e+08 ps=78740 
M2266 diff_1804670_1625600# diff_1795780_1543050# diff_580390_1633220# GND efet w=10160 l=7620
+ ad=2.85483e+08 pd=78740 as=0 ps=0 
M2267 GND diff_1804670_1625600# diff_1831340_1645920# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2268 diff_1879600_1640840# diff_1868170_1628140# GND GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2269 GND diff_1950720_1775460# diff_1976120_1797050# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2270 diff_2025650_1790700# diff_2014220_1776730# GND GND efet w=26670 l=8890
+ ad=2.66128e+08 pd=76200 as=0 ps=0 
M2271 diff_703580_1781810# diff_2019300_1526540# diff_2025650_1790700# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2272 diff_1976120_1681480# diff_1964690_1543050# diff_703580_1714500# GND efet w=22225 l=8255
+ ad=2.91935e+08 pd=78740 as=0 ps=0 
M2273 GND diff_1950720_1715770# diff_1976120_1681480# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2274 diff_2025650_1685290# diff_2014220_1714500# GND GND efet w=24765 l=8255
+ ad=2.62903e+08 pd=76200 as=0 ps=0 
M2275 GND diff_2095500_1926590# diff_2122170_1946910# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2276 diff_2171700_1941830# diff_2160270_1926590# GND GND efet w=24130 l=7620
+ ad=2.59677e+08 pd=76200 as=0 ps=0 
M2277 diff_703580_1931670# diff_2165350_1529080# diff_2171700_1941830# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2278 diff_2122170_1831340# diff_2110740_1545590# diff_703580_1863090# GND efet w=22860 l=7620
+ ad=2.93548e+08 pd=81280 as=0 ps=0 
M2279 GND diff_2095500_1866900# diff_2122170_1831340# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2280 diff_2171700_1835150# diff_2160270_1864360# GND GND efet w=26670 l=8255
+ ad=2.59677e+08 pd=76200 as=0 ps=0 
M2281 GND diff_2241550_2076450# diff_2268220_2098040# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2282 o3 diff_2513330_2120900# Vdd GND efet w=218440 l=7620
+ ad=2.25991e+08 pd=723900 as=0 ps=0 
M2283 diff_2598420_2186940# diff_2557780_2068830# GND GND efet w=29210 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2284 o3 diff_2557780_2068830# GND GND efet w=205105 l=6985
+ ad=0 pd=0 as=0 ps=0 
M2285 Vdd diff_2354580_1676400# diff_703580_2081530# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2286 Vdd diff_2002790_702310# diff_580390_2082800# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2287 diff_2513330_2120900# diff_2513330_2120900# diff_2513330_2120900# GND efet w=1905 l=3175
+ ad=1.10322e+09 pd=182880 as=0 ps=0 
M2288 diff_2513330_2120900# Vdd Vdd GND efet w=12700 l=19685
+ ad=0 pd=0 as=0 ps=0 
M2289 diff_2513330_2120900# diff_2513330_2120900# diff_2513330_2120900# GND efet w=2540 l=2540
+ ad=0 pd=0 as=0 ps=0 
M2290 diff_2513330_2120900# diff_2557780_2068830# GND GND efet w=53975 l=6985
+ ad=0 pd=0 as=0 ps=0 
M2291 Vdd diff_2002790_702310# diff_580390_2004060# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2292 diff_2268220_1982470# diff_2258060_1543050# diff_703580_2012950# GND efet w=21590 l=7620
+ ad=2.90322e+08 pd=78740 as=0 ps=0 
M2293 GND diff_2241550_2016760# diff_2268220_1982470# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2294 Vdd diff_2354580_1676400# diff_703580_2012950# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2295 diff_2268220_1946910# diff_2258060_1543050# diff_703580_1931670# GND efet w=22225 l=8255
+ ad=2.91935e+08 pd=78740 as=0 ps=0 
M2296 diff_580390_1932940# diff_2203450_1583690# diff_2160270_1926590# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.93548e+08 ps=78740 
M2297 diff_2241550_1926590# diff_2233930_1543050# diff_580390_1932940# GND efet w=8890 l=7620
+ ad=2.99999e+08 pd=83820 as=0 ps=0 
M2298 diff_580390_1854200# diff_2203450_1583690# diff_2160270_1864360# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.99999e+08 ps=81280 
M2299 diff_2241550_1866900# diff_2233930_1543050# diff_580390_1854200# GND efet w=8890 l=7620
+ ad=2.87096e+08 pd=81280 as=0 ps=0 
M2300 diff_703580_1863090# diff_2165350_1529080# diff_2171700_1835150# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2301 diff_2122170_1797050# diff_2110740_1545590# diff_703580_1781810# GND efet w=21590 l=7620
+ ad=2.90322e+08 pd=81280 as=0 ps=0 
M2302 diff_580390_1783080# diff_2057400_1583690# diff_2014220_1776730# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.96774e+08 ps=78740 
M2303 diff_2095500_1775460# diff_2087880_1543050# diff_580390_1783080# GND efet w=8890 l=7620
+ ad=2.96774e+08 pd=83820 as=0 ps=0 
M2304 diff_580390_1704340# diff_2057400_1583690# diff_2014220_1714500# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.93548e+08 ps=78740 
M2305 diff_2095500_1715770# diff_2087880_1543050# diff_580390_1704340# GND efet w=8890 l=7620
+ ad=2.88709e+08 pd=81280 as=0 ps=0 
M2306 diff_703580_1714500# diff_2019300_1526540# diff_2025650_1685290# GND efet w=22225 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2307 diff_1976120_1647190# diff_1964690_1543050# diff_703580_1633220# GND efet w=21590 l=7620
+ ad=2.91935e+08 pd=81280 as=0 ps=0 
M2308 diff_580390_1633220# diff_1911350_1583690# diff_1868170_1628140# GND efet w=10160 l=7620
+ ad=0 pd=0 as=2.99999e+08 ps=78740 
M2309 diff_1950720_1625600# diff_1941830_1543050# diff_580390_1633220# GND efet w=11430 l=8890
+ ad=2.85483e+08 pd=76200 as=0 ps=0 
M2310 GND diff_1950720_1625600# diff_1976120_1647190# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2311 diff_2025650_1640840# diff_2014220_1626870# GND GND efet w=24130 l=8890
+ ad=2.6129e+08 pd=76200 as=0 ps=0 
M2312 diff_703580_1633220# diff_2019300_1526540# diff_2025650_1640840# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2313 GND diff_2095500_1775460# diff_2122170_1797050# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2314 diff_2171700_1790700# diff_2160270_1776730# GND GND efet w=24765 l=8255
+ ad=2.58064e+08 pd=76200 as=0 ps=0 
M2315 diff_703580_1781810# diff_2165350_1529080# diff_2171700_1790700# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2316 diff_2122170_1681480# diff_2110740_1545590# diff_703580_1714500# GND efet w=22225 l=8255
+ ad=2.90322e+08 pd=78740 as=0 ps=0 
M2317 GND diff_2095500_1715770# diff_2122170_1681480# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2318 diff_2171700_1685290# diff_2160270_1714500# GND GND efet w=24130 l=8890
+ ad=2.59677e+08 pd=76200 as=0 ps=0 
M2319 GND diff_2241550_1926590# diff_2268220_1946910# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2320 Vdd diff_2354580_1676400# diff_703580_1931670# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2321 Vdd diff_2002790_702310# diff_580390_1932940# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2322 Vdd diff_2002790_702310# diff_580390_1854200# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2323 diff_2268220_1831340# diff_2258060_1543050# diff_703580_1863090# GND efet w=22860 l=7620
+ ad=2.98386e+08 pd=81280 as=0 ps=0 
M2324 GND diff_2241550_1866900# diff_2268220_1831340# GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2325 Vdd diff_2354580_1676400# diff_703580_1863090# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2326 GND diff_1897380_186690# diff_2198370_3069590# GND efet w=55880 l=6350
+ ad=0 pd=0 as=8.37095e+08 ps=157480 
M2327 diff_2268220_1797050# diff_2258060_1543050# diff_703580_1781810# GND efet w=22860 l=7620
+ ad=2.90322e+08 pd=78740 as=0 ps=0 
M2328 diff_580390_1783080# diff_2203450_1583690# diff_2160270_1776730# GND efet w=10160 l=7620
+ ad=0 pd=0 as=2.91935e+08 ps=81280 
M2329 diff_2241550_1775460# diff_2233930_1543050# diff_580390_1783080# GND efet w=8890 l=7620
+ ad=2.96774e+08 pd=83820 as=0 ps=0 
M2330 diff_580390_1704340# diff_2203450_1583690# diff_2160270_1714500# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.93548e+08 ps=81280 
M2331 diff_2241550_1715770# diff_2233930_1543050# diff_580390_1704340# GND efet w=8890 l=7620
+ ad=2.96774e+08 pd=78740 as=0 ps=0 
M2332 diff_703580_1714500# diff_2165350_1529080# diff_2171700_1685290# GND efet w=22225 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2333 diff_2122170_1647190# diff_2110740_1545590# diff_703580_1633220# GND efet w=21590 l=7620
+ ad=2.79032e+08 pd=76200 as=0 ps=0 
M2334 diff_580390_1633220# diff_2057400_1583690# diff_2014220_1626870# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.99999e+08 ps=78740 
M2335 diff_2095500_1626870# diff_2087880_1543050# diff_580390_1633220# GND efet w=8890 l=7620
+ ad=2.95161e+08 pd=78740 as=0 ps=0 
M2336 GND diff_2095500_1626870# diff_2122170_1647190# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2337 diff_2171700_1642110# diff_2160270_1626870# GND GND efet w=22860 l=8890
+ ad=2.5e+08 pd=73660 as=0 ps=0 
M2338 diff_703580_1633220# diff_2165350_1529080# diff_2171700_1642110# GND efet w=21590 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2339 GND diff_2241550_1775460# diff_2268220_1797050# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2340 Vdd diff_2354580_1676400# diff_703580_1781810# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2341 Vdd diff_2002790_702310# diff_580390_1783080# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2342 diff_2198370_3069590# Vdd Vdd GND efet w=11430 l=19685
+ ad=0 pd=0 as=0 ps=0 
M2343 Vdd diff_2002790_702310# diff_580390_1704340# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2344 diff_2354580_1676400# diff_2415540_1699260# diff_2354580_1676400# GND efet w=32385 l=33655
+ ad=1.65645e+09 pd=279400 as=0 ps=0 
M2345 diff_2268220_1681480# diff_2258060_1543050# diff_703580_1714500# GND efet w=22860 l=7620
+ ad=2.87096e+08 pd=78740 as=0 ps=0 
M2346 GND diff_2241550_1715770# diff_2268220_1681480# GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2347 Vdd diff_2354580_1676400# diff_703580_1714500# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2348 diff_2415540_1699260# Vdd Vdd GND efet w=8890 l=7620
+ ad=2.91935e+08 pd=86360 as=0 ps=0 
M2349 diff_2415540_1699260# diff_2415540_1699260# diff_2415540_1699260# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M2350 diff_2415540_1699260# diff_2415540_1699260# diff_2415540_1699260# GND efet w=2540 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2351 GND diff_2479040_1628140# diff_2354580_1676400# GND efet w=78740 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2352 diff_2354580_1676400# diff_2415540_1699260# Vdd GND efet w=11430 l=12700
+ ad=0 pd=0 as=0 ps=0 
M2353 diff_2354580_1676400# diff_2354580_1676400# diff_2354580_1676400# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M2354 diff_2354580_1676400# diff_2354580_1676400# diff_2354580_1676400# GND efet w=4445 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2355 diff_2268220_1647190# diff_2258060_1543050# diff_703580_1633220# GND efet w=22860 l=7620
+ ad=2.87096e+08 pd=78740 as=0 ps=0 
M2356 diff_580390_1633220# diff_2203450_1583690# diff_2160270_1626870# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.77419e+08 ps=78740 
M2357 diff_2241550_1626870# diff_2233930_1543050# diff_580390_1633220# GND efet w=7620 l=8890
+ ad=2.91935e+08 pd=78740 as=0 ps=0 
M2358 GND diff_2241550_1626870# diff_2268220_1647190# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2359 Vdd diff_2354580_1676400# diff_703580_1633220# GND efet w=14605 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2360 diff_2479040_1628140# Vdd Vdd GND efet w=11430 l=20320
+ ad=1.06613e+09 pd=182880 as=0 ps=0 
M2361 Vdd diff_2002790_702310# diff_580390_1633220# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2362 diff_2479040_1628140# clk1 diff_2482850_1590040# GND efet w=77470 l=7620
+ ad=0 pd=0 as=1.44516e+09 ps=281940 
M2363 GND diff_2476500_1567180# diff_2482850_1590040# GND efet w=120650 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2364 GND diff_844550_1507490# diff_854710_1527810# GND efet w=19050 l=8890
+ ad=0 pd=0 as=6.0645e+08 ps=127000 
M2365 GND diff_844550_1507490# diff_892810_1584960# GND efet w=12700 l=8890
+ ad=0 pd=0 as=2.25806e+08 ps=60960 
M2366 GND diff_918210_1562100# diff_923290_1543050# GND efet w=12700 l=8890
+ ad=0 pd=0 as=2.25806e+08 ps=60960 
M2367 GND diff_918210_1562100# diff_946150_1543050# GND efet w=19050 l=8890
+ ad=0 pd=0 as=5.54838e+08 ps=124460 
M2368 Vdd Vdd diff_462280_1706880# GND efet w=11430 l=40640
+ ad=0 pd=0 as=1.22419e+09 ps=284480 
M2369 Vdd Vdd diff_350520_1598930# GND efet w=11430 l=44450
+ ad=0 pd=0 as=1.72903e+09 ps=368300 
M2370 diff_346710_1485900# diff_346710_1485900# diff_346710_1485900# GND efet w=3810 l=3810
+ ad=1.48871e+09 pd=297180 as=0 ps=0 
M2371 Vdd Vdd diff_346710_1485900# GND efet w=11430 l=39370
+ ad=0 pd=0 as=0 ps=0 
M2372 diff_346710_1485900# diff_346710_1485900# diff_346710_1485900# GND efet w=1905 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2373 diff_450850_1684020# diff_755650_927100# Vdd GND efet w=40640 l=7620
+ ad=-1.39497e+09 pd=464820 as=0 ps=0 
M2374 GND diff_774700_1455420# diff_450850_1684020# GND efet w=40640 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2375 diff_868680_1503680# diff_857250_1226820# diff_854710_1527810# GND efet w=33655 l=10795
+ ad=1.68424e+09 pd=2.42316e+06 as=0 ps=0 
M2376 diff_892810_1584960# diff_857250_1226820# diff_894080_1518920# GND efet w=13335 l=8255
+ ad=0 pd=0 as=1.30682e+09 ps=2.12344e+06 
M2377 diff_923290_1543050# diff_918210_1536700# diff_894080_1518920# GND efet w=13335 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2378 diff_946150_1543050# diff_918210_1536700# diff_868680_1503680# GND efet w=33655 l=10795
+ ad=0 pd=0 as=0 ps=0 
M2379 diff_345440_2600960# diff_345440_2600960# diff_345440_2600960# GND efet w=4445 l=4445
+ ad=1.24677e+09 pd=304800 as=0 ps=0 
M2380 Vdd Vdd diff_345440_2600960# GND efet w=11430 l=40640
+ ad=0 pd=0 as=0 ps=0 
M2381 diff_345440_2600960# diff_345440_2600960# diff_345440_2600960# GND efet w=3810 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2382 GND diff_172720_1316990# diff_245110_1436370# GND efet w=41275 l=6985
+ ad=0 pd=0 as=0 ps=0 
M2383 diff_774700_1455420# Vdd Vdd GND efet w=8890 l=40640
+ ad=5.46773e+08 pd=114300 as=0 ps=0 
M2384 GND diff_991870_1504950# diff_1000760_1526540# GND efet w=19050 l=8890
+ ad=0 pd=0 as=5.74192e+08 ps=124460 
M2385 GND diff_991870_1504950# diff_1038860_1543050# GND efet w=13970 l=8890
+ ad=0 pd=0 as=2.48387e+08 ps=63500 
M2386 GND diff_1064260_1562100# diff_1068070_1543050# GND efet w=13970 l=8890
+ ad=0 pd=0 as=2.25806e+08 ps=60960 
M2387 GND diff_1064260_1562100# diff_1092200_1543050# GND efet w=17780 l=8890
+ ad=0 pd=0 as=5.49999e+08 ps=124460 
M2388 diff_868680_1503680# diff_1002030_1186180# diff_1000760_1526540# GND efet w=33655 l=10795
+ ad=0 pd=0 as=0 ps=0 
M2389 diff_1038860_1543050# diff_1002030_1186180# diff_894080_1518920# GND efet w=15240 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2390 diff_1068070_1543050# diff_1064260_1535430# diff_894080_1518920# GND efet w=13335 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2391 diff_1092200_1543050# diff_1064260_1535430# diff_868680_1503680# GND efet w=33020 l=11430
+ ad=0 pd=0 as=0 ps=0 
M2392 GND diff_1137920_1470660# diff_1145540_1527810# GND efet w=19050 l=8890
+ ad=0 pd=0 as=5.99999e+08 ps=129540 
M2393 GND diff_1137920_1470660# diff_1183640_1584960# GND efet w=12700 l=8890
+ ad=0 pd=0 as=2.25806e+08 ps=60960 
M2394 GND diff_1209040_1562100# diff_1214120_1543050# GND efet w=12700 l=8890
+ ad=0 pd=0 as=2.25806e+08 ps=60960 
M2395 GND diff_1209040_1562100# diff_1236980_1543050# GND efet w=19050 l=8890
+ ad=0 pd=0 as=5.82257e+08 ps=127000 
M2396 diff_868680_1503680# diff_1148080_1228090# diff_1145540_1527810# GND efet w=36195 l=10795
+ ad=0 pd=0 as=0 ps=0 
M2397 diff_1183640_1584960# diff_1148080_1228090# diff_894080_1518920# GND efet w=13335 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2398 diff_1214120_1543050# diff_1209040_1535430# diff_894080_1518920# GND efet w=13335 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2399 diff_1236980_1543050# diff_1209040_1535430# diff_868680_1503680# GND efet w=33655 l=10795
+ ad=0 pd=0 as=0 ps=0 
M2400 GND diff_1282700_1504950# diff_1291590_1526540# GND efet w=17780 l=8890
+ ad=0 pd=0 as=5.66128e+08 ps=124460 
M2401 GND diff_1282700_1504950# diff_1329690_1543050# GND efet w=13970 l=8890
+ ad=0 pd=0 as=2.48387e+08 ps=63500 
M2402 GND diff_1355090_1562100# diff_1358900_1543050# GND efet w=13970 l=8890
+ ad=0 pd=0 as=2.48387e+08 ps=63500 
M2403 GND diff_1355090_1562100# diff_1383030_1543050# GND efet w=17780 l=8890
+ ad=0 pd=0 as=5.61289e+08 ps=124460 
M2404 diff_868680_1503680# diff_1292860_1226820# diff_1291590_1526540# GND efet w=32385 l=10795
+ ad=0 pd=0 as=0 ps=0 
M2405 diff_1329690_1543050# diff_1292860_1226820# diff_894080_1518920# GND efet w=14605 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2406 diff_1358900_1543050# diff_1355090_1535430# diff_894080_1518920# GND efet w=15875 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2407 diff_1383030_1543050# diff_1355090_1535430# diff_868680_1503680# GND efet w=33020 l=11430
+ ad=0 pd=0 as=0 ps=0 
M2408 GND diff_1428750_1470660# diff_1436370_1529080# GND efet w=19050 l=8890
+ ad=0 pd=0 as=5.82257e+08 ps=127000 
M2409 GND diff_1428750_1470660# diff_1474470_1583690# GND efet w=12700 l=8890
+ ad=0 pd=0 as=2.25806e+08 ps=60960 
M2410 GND diff_1499870_1562100# diff_1504950_1543050# GND efet w=12700 l=8890
+ ad=0 pd=0 as=2.25806e+08 ps=60960 
M2411 GND diff_1499870_1562100# diff_1527810_1543050# GND efet w=19050 l=8890
+ ad=0 pd=0 as=5.85483e+08 ps=127000 
M2412 diff_868680_1503680# diff_1438910_1226820# diff_1436370_1529080# GND efet w=34925 l=10795
+ ad=0 pd=0 as=0 ps=0 
M2413 diff_1474470_1583690# diff_1438910_1226820# diff_894080_1518920# GND efet w=13335 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2414 diff_1504950_1543050# diff_1499870_1535430# diff_894080_1518920# GND efet w=13335 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2415 diff_1527810_1543050# diff_1499870_1535430# diff_868680_1503680# GND efet w=33655 l=10795
+ ad=0 pd=0 as=0 ps=0 
M2416 GND diff_1573530_1504950# diff_1582420_1527810# GND efet w=19050 l=8890
+ ad=0 pd=0 as=5.64515e+08 ps=127000 
M2417 GND diff_1573530_1504950# diff_1620520_1543050# GND efet w=13970 l=8255
+ ad=0 pd=0 as=2.48387e+08 ps=63500 
M2418 GND diff_1645920_1562100# diff_1649730_1543050# GND efet w=13335 l=8890
+ ad=0 pd=0 as=2.48387e+08 ps=63500 
M2419 GND diff_1645920_1562100# diff_1673860_1543050# GND efet w=19050 l=8890
+ ad=0 pd=0 as=5.59676e+08 ps=124460 
M2420 diff_868680_1503680# diff_1584960_1226820# diff_1582420_1527810# GND efet w=33655 l=10795
+ ad=0 pd=0 as=0 ps=0 
M2421 diff_1620520_1543050# diff_1584960_1226820# diff_894080_1518920# GND efet w=14605 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2422 diff_1649730_1543050# diff_1645920_1535430# diff_894080_1518920# GND efet w=14605 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2423 diff_1673860_1543050# diff_1645920_1535430# diff_868680_1503680# GND efet w=34290 l=11430
+ ad=0 pd=0 as=0 ps=0 
M2424 GND diff_1719580_1478280# diff_1728470_1526540# GND efet w=19050 l=8890
+ ad=0 pd=0 as=5.61289e+08 ps=124460 
M2425 GND diff_1719580_1478280# diff_1765300_1584960# GND efet w=13335 l=8255
+ ad=0 pd=0 as=2.25806e+08 ps=60960 
M2426 GND diff_1790700_1562100# diff_1795780_1543050# GND efet w=12700 l=8890
+ ad=0 pd=0 as=2.25806e+08 ps=60960 
M2427 diff_1819910_1543050# diff_1790700_1562100# GND GND efet w=17780 l=8890
+ ad=5.62902e+08 pd=124460 as=0 ps=0 
M2428 diff_868680_1503680# diff_1729740_1228090# diff_1728470_1526540# GND efet w=34925 l=10795
+ ad=0 pd=0 as=0 ps=0 
M2429 diff_1765300_1584960# diff_1729740_1228090# diff_894080_1518920# GND efet w=13335 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2430 diff_1795780_1543050# diff_1790700_1535430# diff_894080_1518920# GND efet w=13335 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2431 diff_1819910_1543050# diff_1790700_1535430# diff_868680_1503680# GND efet w=33655 l=10795
+ ad=0 pd=0 as=0 ps=0 
M2432 GND diff_1864360_1504950# diff_1873250_1527810# GND efet w=19050 l=8890
+ ad=0 pd=0 as=5.8387e+08 ps=127000 
M2433 GND diff_1864360_1504950# diff_1911350_1583690# GND efet w=12700 l=8255
+ ad=0 pd=0 as=2.25806e+08 ps=60960 
M2434 GND diff_1936750_1562100# diff_1941830_1543050# GND efet w=12700 l=8890
+ ad=0 pd=0 as=2.25806e+08 ps=60960 
M2435 GND diff_1936750_1562100# diff_1964690_1543050# GND efet w=20320 l=8890
+ ad=0 pd=0 as=5.88708e+08 ps=129540 
M2436 diff_868680_1503680# diff_1861820_1186180# diff_1873250_1527810# GND efet w=34925 l=10795
+ ad=0 pd=0 as=0 ps=0 
M2437 diff_1911350_1583690# diff_1861820_1186180# diff_894080_1518920# GND efet w=13335 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2438 diff_1941830_1543050# diff_1926590_1210310# diff_894080_1518920# GND efet w=13335 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2439 diff_1964690_1543050# diff_1926590_1210310# diff_868680_1503680# GND efet w=34925 l=10795
+ ad=0 pd=0 as=0 ps=0 
M2440 GND diff_2010410_1504950# diff_2019300_1526540# GND efet w=20955 l=8255
+ ad=0 pd=0 as=5.74192e+08 ps=134620 
M2441 GND diff_2010410_1504950# diff_2057400_1583690# GND efet w=12700 l=7620
+ ad=0 pd=0 as=2.41935e+08 ps=63500 
M2442 GND diff_2082800_1562100# diff_2087880_1543050# GND efet w=13970 l=7620
+ ad=0 pd=0 as=2.38709e+08 ps=66040 
M2443 diff_2110740_1545590# diff_2082800_1562100# GND GND efet w=18415 l=8255
+ ad=5.93547e+08 pd=129540 as=0 ps=0 
M2444 diff_868680_1503680# diff_2002790_1228090# diff_2019300_1526540# GND efet w=33020 l=11430
+ ad=0 pd=0 as=0 ps=0 
M2445 diff_2057400_1583690# diff_2002790_1228090# diff_894080_1518920# GND efet w=12700 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2446 diff_2087880_1543050# diff_2080260_1351280# diff_894080_1518920# GND efet w=13335 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2447 diff_2110740_1545590# diff_2080260_1351280# diff_868680_1503680# GND efet w=33020 l=10795
+ ad=0 pd=0 as=0 ps=0 
M2448 GND diff_2156460_1504950# diff_2165350_1529080# GND efet w=20955 l=7620
+ ad=0 pd=0 as=5.87096e+08 ps=132080 
M2449 GND diff_2156460_1504950# diff_2203450_1583690# GND efet w=12700 l=7620
+ ad=0 pd=0 as=2.41935e+08 ps=63500 
M2450 GND diff_2228850_1562100# diff_2233930_1543050# GND efet w=12700 l=7620
+ ad=0 pd=0 as=2.41935e+08 ps=63500 
M2451 diff_2258060_1543050# diff_2228850_1562100# GND GND efet w=17780 l=7620
+ ad=5.8387e+08 pd=127000 as=0 ps=0 
M2452 diff_2476500_1567180# Vdd Vdd GND efet w=11430 l=29210
+ ad=1.03226e+09 pd=223520 as=0 ps=0 
M2453 diff_2476500_1567180# diff_2476500_1567180# diff_2476500_1567180# GND efet w=2540 l=5080
+ ad=0 pd=0 as=0 ps=0 
M2454 diff_2476500_1567180# diff_2476500_1567180# diff_2476500_1567180# GND efet w=2540 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2455 diff_868680_1503680# diff_2128520_1299210# diff_2165350_1529080# GND efet w=34925 l=10795
+ ad=0 pd=0 as=0 ps=0 
M2456 diff_2203450_1583690# diff_2128520_1299210# diff_894080_1518920# GND efet w=12700 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2457 diff_2233930_1543050# diff_2172970_1249680# diff_894080_1518920# GND efet w=12700 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2458 diff_2258060_1543050# diff_2172970_1249680# diff_868680_1503680# GND efet w=33020 l=10160
+ ad=0 pd=0 as=0 ps=0 
M2459 diff_844550_1507490# diff_844550_1507490# diff_844550_1507490# GND efet w=5080 l=7620
+ ad=6.01612e+08 pd=154940 as=0 ps=0 
M2460 diff_844550_1507490# diff_844550_1507490# diff_844550_1507490# GND efet w=6350 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2461 GND diff_857250_1226820# diff_844550_1507490# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2462 diff_918210_1562100# diff_918210_1536700# GND GND efet w=15240 l=7620
+ ad=5.64515e+08 pd=149860 as=0 ps=0 
M2463 diff_918210_1562100# diff_918210_1562100# diff_918210_1562100# GND efet w=5080 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2464 diff_918210_1562100# diff_918210_1562100# diff_918210_1562100# GND efet w=6350 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2465 Vdd Vdd diff_844550_1507490# GND efet w=7620 l=40640
+ ad=0 pd=0 as=0 ps=0 
M2466 GND diff_755650_927100# diff_774700_1455420# GND efet w=20320 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2467 d3 GND GND GND efet w=109220 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2468 diff_245110_1436370# diff_180340_1348740# Vdd GND efet w=40640 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2469 diff_857250_1226820# diff_857250_1226820# diff_857250_1226820# GND efet w=3175 l=3175
+ ad=2.11935e+09 pd=497840 as=0 ps=0 
M2470 diff_350520_1598930# diff_546100_1416050# GND GND efet w=26670 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2471 diff_345440_2600960# diff_546100_1416050# GND GND efet w=26670 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2472 diff_180340_1348740# diff_172720_1316990# GND GND efet w=24130 l=7620
+ ad=1.58064e+09 pd=292100 as=0 ps=0 
M2473 diff_180340_1348740# diff_180340_1348740# diff_180340_1348740# GND efet w=2540 l=2540
+ ad=0 pd=0 as=0 ps=0 
M2474 diff_180340_1348740# diff_180340_1348740# diff_180340_1348740# GND efet w=1905 l=5715
+ ad=0 pd=0 as=0 ps=0 
M2475 Vdd Vdd diff_180340_1348740# GND efet w=8890 l=38735
+ ad=0 pd=0 as=0 ps=0 
M2476 diff_857250_1226820# diff_857250_1226820# diff_857250_1226820# GND efet w=2540 l=5080
+ ad=0 pd=0 as=0 ps=0 
M2477 diff_991870_1504950# diff_991870_1504950# diff_991870_1504950# GND efet w=5080 l=6350
+ ad=5.93547e+08 pd=149860 as=0 ps=0 
M2478 diff_991870_1504950# diff_991870_1504950# diff_991870_1504950# GND efet w=5715 l=3175
+ ad=0 pd=0 as=0 ps=0 
M2479 GND diff_1002030_1186180# diff_991870_1504950# GND efet w=15240 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2480 diff_1064260_1562100# diff_1064260_1535430# GND GND efet w=17780 l=7620
+ ad=5.77418e+08 pd=154940 as=0 ps=0 
M2481 diff_1064260_1562100# diff_1064260_1562100# diff_1064260_1562100# GND efet w=5080 l=6350
+ ad=0 pd=0 as=0 ps=0 
M2482 diff_1064260_1562100# diff_1064260_1562100# diff_1064260_1562100# GND efet w=5715 l=3175
+ ad=0 pd=0 as=0 ps=0 
M2483 Vdd Vdd diff_918210_1562100# GND efet w=9525 l=53340
+ ad=0 pd=0 as=0 ps=0 
M2484 diff_991870_1504950# Vdd Vdd GND efet w=9525 l=48260
+ ad=0 pd=0 as=0 ps=0 
M2485 diff_918210_1536700# diff_918210_1536700# diff_918210_1536700# GND efet w=2540 l=3810
+ ad=-2.09981e+09 pd=482600 as=0 ps=0 
M2486 diff_918210_1536700# diff_918210_1536700# diff_918210_1536700# GND efet w=3810 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2487 diff_1002030_1186180# diff_1002030_1186180# diff_1002030_1186180# GND efet w=3175 l=3175
+ ad=1.98225e+09 pd=523240 as=0 ps=0 
M2488 diff_1002030_1186180# diff_1002030_1186180# diff_1002030_1186180# GND efet w=2540 l=6350
+ ad=0 pd=0 as=0 ps=0 
M2489 diff_1137920_1470660# diff_1137920_1470660# diff_1137920_1470660# GND efet w=5080 l=7620
+ ad=6.04838e+08 pd=154940 as=0 ps=0 
M2490 diff_1137920_1470660# diff_1137920_1470660# diff_1137920_1470660# GND efet w=6350 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2491 GND diff_1148080_1228090# diff_1137920_1470660# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2492 diff_1209040_1562100# diff_1209040_1535430# GND GND efet w=15240 l=7620
+ ad=5.82257e+08 pd=152400 as=0 ps=0 
M2493 diff_1209040_1562100# diff_1209040_1562100# diff_1209040_1562100# GND efet w=5080 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2494 diff_1282700_1504950# diff_1282700_1504950# diff_1282700_1504950# GND efet w=5080 l=7620
+ ad=5.85483e+08 pd=149860 as=0 ps=0 
M2495 diff_1209040_1562100# diff_1209040_1562100# diff_1209040_1562100# GND efet w=6350 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2496 Vdd Vdd diff_1064260_1562100# GND efet w=9525 l=50800
+ ad=0 pd=0 as=0 ps=0 
M2497 diff_1137920_1470660# Vdd Vdd GND efet w=9525 l=50800
+ ad=0 pd=0 as=0 ps=0 
M2498 diff_1064260_1535430# diff_1064260_1535430# diff_1064260_1535430# GND efet w=2540 l=3175
+ ad=2.11935e+09 pd=480060 as=0 ps=0 
M2499 diff_1064260_1535430# diff_1064260_1535430# diff_1064260_1535430# GND efet w=4445 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2500 diff_1148080_1228090# diff_1148080_1228090# diff_1148080_1228090# GND efet w=3810 l=3810
+ ad=2.1e+09 pd=497840 as=0 ps=0 
M2501 diff_1148080_1228090# diff_1148080_1228090# diff_1148080_1228090# GND efet w=2540 l=5080
+ ad=0 pd=0 as=0 ps=0 
M2502 GND diff_1292860_1226820# diff_1282700_1504950# GND efet w=16510 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2503 diff_1282700_1504950# diff_1282700_1504950# diff_1282700_1504950# GND efet w=5715 l=3175
+ ad=0 pd=0 as=0 ps=0 
M2504 diff_1355090_1562100# diff_1355090_1535430# GND GND efet w=15240 l=7620
+ ad=5.8387e+08 pd=152400 as=0 ps=0 
M2505 diff_1355090_1562100# diff_1355090_1562100# diff_1355090_1562100# GND efet w=5080 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2506 diff_1355090_1562100# diff_1355090_1562100# diff_1355090_1562100# GND efet w=6350 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2507 diff_1209040_1562100# Vdd Vdd GND efet w=10795 l=49530
+ ad=0 pd=0 as=0 ps=0 
M2508 diff_1282700_1504950# Vdd Vdd GND efet w=10795 l=50165
+ ad=0 pd=0 as=0 ps=0 
M2509 diff_1209040_1535430# diff_1209040_1535430# diff_1209040_1535430# GND efet w=2540 l=3810
+ ad=-2.14497e+09 pd=469900 as=0 ps=0 
M2510 diff_1209040_1535430# diff_1209040_1535430# diff_1209040_1535430# GND efet w=4445 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2511 diff_1292860_1226820# diff_1292860_1226820# diff_1292860_1226820# GND efet w=3175 l=3175
+ ad=2.08548e+09 pd=500380 as=0 ps=0 
M2512 diff_1292860_1226820# diff_1292860_1226820# diff_1292860_1226820# GND efet w=3175 l=6350
+ ad=0 pd=0 as=0 ps=0 
M2513 diff_1428750_1470660# diff_1428750_1470660# diff_1428750_1470660# GND efet w=5715 l=6985
+ ad=5.96773e+08 pd=160020 as=0 ps=0 
M2514 GND diff_1438910_1226820# diff_1428750_1470660# GND efet w=18415 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2515 diff_1499870_1562100# diff_1499870_1535430# GND GND efet w=17780 l=8255
+ ad=5.88708e+08 pd=149860 as=0 ps=0 
M2516 diff_1499870_1562100# diff_1499870_1562100# diff_1499870_1562100# GND efet w=5080 l=6350
+ ad=0 pd=0 as=0 ps=0 
M2517 diff_1428750_1470660# diff_1428750_1470660# diff_1428750_1470660# GND efet w=5715 l=3175
+ ad=0 pd=0 as=0 ps=0 
M2518 diff_1499870_1562100# diff_1499870_1562100# diff_1499870_1562100# GND efet w=5715 l=3175
+ ad=0 pd=0 as=0 ps=0 
M2519 Vdd Vdd diff_1355090_1562100# GND efet w=9525 l=49530
+ ad=0 pd=0 as=0 ps=0 
M2520 diff_1428750_1470660# Vdd Vdd GND efet w=9525 l=48260
+ ad=0 pd=0 as=0 ps=0 
M2521 diff_1355090_1535430# diff_1355090_1535430# diff_1355090_1535430# GND efet w=2540 l=3175
+ ad=2.10161e+09 pd=474980 as=0 ps=0 
M2522 diff_1355090_1535430# diff_1355090_1535430# diff_1355090_1535430# GND efet w=4445 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2523 diff_1438910_1226820# diff_1438910_1226820# diff_1438910_1226820# GND efet w=2540 l=3810
+ ad=2.10161e+09 pd=492760 as=0 ps=0 
M2524 diff_1438910_1226820# diff_1438910_1226820# diff_1438910_1226820# GND efet w=2540 l=5080
+ ad=0 pd=0 as=0 ps=0 
M2525 diff_1573530_1504950# diff_1573530_1504950# diff_1573530_1504950# GND efet w=5080 l=7620
+ ad=5.80644e+08 pd=152400 as=0 ps=0 
M2526 GND diff_1584960_1226820# diff_1573530_1504950# GND efet w=16510 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2527 diff_1645920_1562100# diff_1645920_1535430# GND GND efet w=16510 l=7620
+ ad=5.82257e+08 pd=152400 as=0 ps=0 
M2528 diff_1573530_1504950# diff_1573530_1504950# diff_1573530_1504950# GND efet w=6350 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2529 diff_1645920_1562100# diff_1645920_1562100# diff_1645920_1562100# GND efet w=5080 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2530 diff_1719580_1478280# diff_1719580_1478280# diff_1719580_1478280# GND efet w=5080 l=7620
+ ad=5.91934e+08 pd=154940 as=0 ps=0 
M2531 diff_1645920_1562100# diff_1645920_1562100# diff_1645920_1562100# GND efet w=5715 l=3175
+ ad=0 pd=0 as=0 ps=0 
M2532 diff_1719580_1478280# diff_1719580_1478280# diff_1719580_1478280# GND efet w=5715 l=3175
+ ad=0 pd=0 as=0 ps=0 
M2533 GND diff_1729740_1228090# diff_1719580_1478280# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2534 diff_1790700_1562100# diff_1790700_1535430# GND GND efet w=15240 l=7620
+ ad=5.8387e+08 pd=152400 as=0 ps=0 
M2535 diff_1790700_1562100# diff_1790700_1562100# diff_1790700_1562100# GND efet w=5080 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2536 diff_1790700_1562100# diff_1790700_1562100# diff_1790700_1562100# GND efet w=6350 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2537 Vdd Vdd diff_1499870_1562100# GND efet w=8890 l=50165
+ ad=0 pd=0 as=0 ps=0 
M2538 diff_1573530_1504950# Vdd Vdd GND efet w=9525 l=51435
+ ad=0 pd=0 as=0 ps=0 
M2539 diff_1499870_1535430# diff_1499870_1535430# diff_1499870_1535430# GND efet w=2540 l=3175
+ ad=-2.13046e+09 pd=469900 as=0 ps=0 
M2540 diff_1499870_1535430# diff_1499870_1535430# diff_1499870_1535430# GND efet w=3810 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2541 diff_1584960_1226820# diff_1584960_1226820# diff_1584960_1226820# GND efet w=3175 l=3175
+ ad=1.92096e+09 pd=449580 as=0 ps=0 
M2542 diff_1584960_1226820# diff_1584960_1226820# diff_1584960_1226820# GND efet w=2540 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2543 Vdd Vdd diff_1645920_1562100# GND efet w=9525 l=50165
+ ad=0 pd=0 as=0 ps=0 
M2544 diff_1719580_1478280# Vdd Vdd GND efet w=8255 l=49530
+ ad=0 pd=0 as=0 ps=0 
M2545 diff_1645920_1535430# diff_1645920_1535430# diff_1645920_1535430# GND efet w=2540 l=3175
+ ad=-2.12078e+09 pd=553720 as=0 ps=0 
M2546 diff_1645920_1535430# diff_1645920_1535430# diff_1645920_1535430# GND efet w=3810 l=5080
+ ad=0 pd=0 as=0 ps=0 
M2547 diff_1729740_1228090# diff_1729740_1228090# diff_1729740_1228090# GND efet w=3175 l=3175
+ ad=2.1258e+09 pd=505460 as=0 ps=0 
M2548 diff_1729740_1228090# diff_1729740_1228090# diff_1729740_1228090# GND efet w=2540 l=5080
+ ad=0 pd=0 as=0 ps=0 
M2549 diff_1864360_1504950# diff_1864360_1504950# diff_1864360_1504950# GND efet w=5080 l=6350
+ ad=5.91934e+08 pd=149860 as=0 ps=0 
M2550 diff_1864360_1504950# diff_1864360_1504950# diff_1864360_1504950# GND efet w=5715 l=3175
+ ad=0 pd=0 as=0 ps=0 
M2551 GND diff_1861820_1186180# diff_1864360_1504950# GND efet w=15240 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2552 diff_1936750_1562100# diff_1926590_1210310# GND GND efet w=17145 l=8255
+ ad=5.93547e+08 pd=149860 as=0 ps=0 
M2553 diff_1936750_1562100# diff_1936750_1562100# diff_1936750_1562100# GND efet w=5080 l=6350
+ ad=0 pd=0 as=0 ps=0 
M2554 diff_1936750_1562100# diff_1936750_1562100# diff_1936750_1562100# GND efet w=5715 l=3175
+ ad=0 pd=0 as=0 ps=0 
M2555 Vdd Vdd diff_1790700_1562100# GND efet w=9525 l=49530
+ ad=0 pd=0 as=0 ps=0 
M2556 diff_1864360_1504950# Vdd Vdd GND efet w=8890 l=48895
+ ad=0 pd=0 as=0 ps=0 
M2557 diff_1790700_1535430# diff_1790700_1535430# diff_1790700_1535430# GND efet w=1905 l=4445
+ ad=-1.91271e+09 pd=561340 as=0 ps=0 
M2558 diff_1790700_1535430# diff_1790700_1535430# diff_1790700_1535430# GND efet w=3810 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2559 diff_1861820_1186180# diff_1861820_1186180# diff_1861820_1186180# GND efet w=3810 l=5080
+ ad=-1.81594e+09 pd=591820 as=0 ps=0 
M2560 diff_1861820_1186180# diff_1861820_1186180# diff_1861820_1186180# GND efet w=1905 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2561 diff_2010410_1504950# diff_2010410_1504950# diff_2010410_1504950# GND efet w=5080 l=7620
+ ad=6.04838e+08 pd=154940 as=0 ps=0 
M2562 diff_2010410_1504950# diff_2010410_1504950# diff_2010410_1504950# GND efet w=6350 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2563 GND diff_2002790_1228090# diff_2010410_1504950# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2564 diff_2082800_1562100# diff_2080260_1351280# GND GND efet w=15240 l=7620
+ ad=5.85483e+08 pd=152400 as=0 ps=0 
M2565 diff_2082800_1562100# diff_2082800_1562100# diff_2082800_1562100# GND efet w=5080 l=6350
+ ad=0 pd=0 as=0 ps=0 
M2566 diff_2156460_1504950# diff_2156460_1504950# diff_2156460_1504950# GND efet w=5080 l=7620
+ ad=5.85483e+08 pd=152400 as=0 ps=0 
M2567 diff_2082800_1562100# diff_2082800_1562100# diff_2082800_1562100# GND efet w=5715 l=3175
+ ad=0 pd=0 as=0 ps=0 
M2568 Vdd Vdd diff_1936750_1562100# GND efet w=9525 l=50165
+ ad=0 pd=0 as=0 ps=0 
M2569 diff_2010410_1504950# Vdd Vdd GND efet w=9525 l=49530
+ ad=0 pd=0 as=0 ps=0 
M2570 diff_1926590_1210310# diff_1926590_1210310# diff_1926590_1210310# GND efet w=1905 l=2540
+ ad=-1.65304e+09 pd=645160 as=0 ps=0 
M2571 diff_1926590_1210310# diff_1926590_1210310# diff_1926590_1210310# GND efet w=3810 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2572 diff_857250_1226820# diff_872490_1417320# GND GND efet w=16510 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2573 diff_918210_1536700# diff_872490_1417320# GND GND efet w=17780 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2574 diff_1002030_1186180# diff_872490_1417320# GND GND efet w=17145 l=9525
+ ad=0 pd=0 as=0 ps=0 
M2575 diff_1064260_1535430# diff_872490_1417320# GND GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2576 diff_1148080_1228090# diff_872490_1417320# GND GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2577 diff_1209040_1535430# diff_872490_1417320# GND GND efet w=17145 l=9525
+ ad=0 pd=0 as=0 ps=0 
M2578 diff_1292860_1226820# diff_872490_1417320# GND GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2579 diff_1355090_1535430# diff_872490_1417320# GND GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2580 diff_1438910_1226820# diff_1377950_1109980# GND GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2581 diff_1499870_1535430# diff_1377950_1109980# GND GND efet w=17145 l=9525
+ ad=0 pd=0 as=0 ps=0 
M2582 diff_1584960_1226820# diff_1377950_1109980# GND GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2583 diff_1645920_1535430# diff_1377950_1109980# GND GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2584 diff_1729740_1228090# diff_1377950_1109980# GND GND efet w=17780 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2585 diff_1790700_1535430# diff_1377950_1109980# GND GND efet w=16510 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2586 diff_1861820_1186180# diff_1377950_1109980# GND GND efet w=17780 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2587 diff_1926590_1210310# diff_1377950_1109980# GND GND efet w=16510 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2588 diff_2156460_1504950# diff_2156460_1504950# diff_2156460_1504950# GND efet w=6350 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2589 GND diff_2128520_1299210# diff_2156460_1504950# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2590 diff_2476500_1567180# diff_284480_472440# diff_2486660_1535430# GND efet w=73025 l=6985
+ ad=0 pd=0 as=1.08871e+09 ps=213360 
M2591 diff_2486660_1535430# diff_829310_237490# GND GND efet w=76200 l=6985
+ ad=0 pd=0 as=0 ps=0 
M2592 diff_2228850_1562100# diff_2228850_1562100# diff_2228850_1562100# GND efet w=1270 l=2540
+ ad=6.77418e+08 pd=205740 as=0 ps=0 
M2593 Vdd Vdd diff_2082800_1562100# GND efet w=8255 l=48895
+ ad=0 pd=0 as=0 ps=0 
M2594 diff_2156460_1504950# Vdd Vdd GND efet w=9525 l=49530
+ ad=0 pd=0 as=0 ps=0 
M2595 diff_2228850_1562100# diff_2228850_1562100# diff_2228850_1562100# GND efet w=2540 l=2540
+ ad=0 pd=0 as=0 ps=0 
M2596 diff_868680_1503680# diff_2444750_1443990# Vdd GND efet w=40640 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2597 diff_2228850_1562100# diff_2172970_1249680# GND GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2598 Vdd Vdd diff_2228850_1562100# GND efet w=6985 l=47625
+ ad=0 pd=0 as=0 ps=0 
M2599 GND diff_2471420_1322070# diff_868680_1503680# GND efet w=46355 l=6350
+ ad=0 pd=0 as=0 ps=0 
M2600 GND diff_2471420_1322070# diff_2444750_1443990# GND efet w=43180 l=7620
+ ad=0 pd=0 as=1.74193e+09 ps=406400 
M2601 GND diff_546100_1388110# diff_346710_1485900# GND efet w=26670 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2602 GND diff_546100_1388110# diff_462280_1706880# GND efet w=26670 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2603 diff_553720_1553210# diff_232410_996950# Vdd GND efet w=31115 l=7620
+ ad=1.67258e+09 pd=271780 as=0 ps=0 
M2604 GND diff_774700_1325880# diff_553720_1553210# GND efet w=29210 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2605 GND diff_869950_1397000# diff_857250_1226820# GND efet w=17780 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2606 diff_918210_1536700# diff_869950_1397000# GND GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2607 GND diff_869950_1397000# diff_1002030_1186180# GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2608 GND diff_869950_1397000# diff_1064260_1535430# GND efet w=18415 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2609 GND diff_869950_1397000# diff_1438910_1226820# GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2610 diff_1499870_1535430# diff_869950_1397000# GND GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2611 GND diff_869950_1397000# diff_1584960_1226820# GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2612 diff_1645920_1535430# diff_869950_1397000# GND GND efet w=17145 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2613 diff_2172970_1249680# diff_2197100_1388110# diff_2172970_1249680# GND efet w=88900 l=3810
+ ad=-2.03368e+09 pd=609600 as=0 ps=0 
M2614 diff_1148080_1228090# diff_1160780_1371600# GND GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2615 diff_1209040_1535430# diff_1160780_1371600# GND GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2616 diff_1292860_1226820# diff_1160780_1371600# GND GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2617 diff_1355090_1535430# diff_1160780_1371600# GND GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2618 diff_1729740_1228090# diff_1160780_1371600# GND GND efet w=17145 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2619 diff_1790700_1535430# diff_1160780_1371600# GND GND efet w=18415 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2620 diff_1861820_1186180# diff_1160780_1371600# GND GND efet w=16510 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2621 diff_1926590_1210310# diff_1160780_1371600# GND GND efet w=16510 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2622 Vdd diff_2197100_1388110# diff_2172970_1249680# GND efet w=8890 l=38100
+ ad=0 pd=0 as=0 ps=0 
M2623 diff_2197100_1388110# diff_2197100_1388110# diff_2197100_1388110# GND efet w=1270 l=3810
+ ad=2.79032e+08 pd=83820 as=0 ps=0 
M2624 diff_2197100_1388110# diff_2197100_1388110# diff_2197100_1388110# GND efet w=2540 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2625 Vdd Vdd diff_2197100_1388110# GND efet w=8890 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2626 diff_2444750_1443990# diff_2439670_1344930# Vdd GND efet w=10160 l=20320
+ ad=0 pd=0 as=0 ps=0 
M2627 diff_2002790_1228090# diff_2012950_1370330# GND GND efet w=21590 l=8255
+ ad=2.05967e+09 pd=411480 as=0 ps=0 
M2628 diff_346710_1485900# diff_546100_1341120# GND GND efet w=26670 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2629 diff_345440_2600960# diff_546100_1341120# GND GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2630 diff_180340_1348740# diff_139700_2962910# GND GND efet w=38100 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2631 diff_172720_1316990# diff_172720_1316990# diff_172720_1316990# GND efet w=2540 l=7620
+ ad=1.34838e+09 pd=304800 as=0 ps=0 
M2632 diff_172720_1316990# diff_172720_1316990# diff_172720_1316990# GND efet w=2540 l=6350
+ ad=0 pd=0 as=0 ps=0 
M2633 diff_172720_1316990# d3 GND GND efet w=58420 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2634 diff_774700_1325880# Vdd Vdd GND efet w=8890 l=41275
+ ad=4.20967e+08 pd=96520 as=0 ps=0 
M2635 diff_857250_1226820# diff_869950_1347470# GND GND efet w=18415 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2636 diff_918210_1536700# diff_869950_1347470# GND GND efet w=16510 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2637 GND diff_869950_1347470# diff_1148080_1228090# GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2638 GND diff_232410_996950# diff_774700_1325880# GND efet w=20955 l=9525
+ ad=0 pd=0 as=0 ps=0 
M2639 diff_1209040_1535430# diff_869950_1347470# GND GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2640 diff_2172970_1249680# diff_2012950_1370330# GND GND efet w=20320 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2641 diff_2444750_1443990# diff_2439670_1344930# diff_2444750_1443990# GND efet w=57150 l=11430
+ ad=0 pd=0 as=0 ps=0 
M2642 GND diff_546100_1313180# diff_350520_1598930# GND efet w=26670 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2643 GND diff_546100_1313180# diff_462280_1706880# GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2644 diff_1438910_1226820# diff_869950_1347470# GND GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2645 diff_1499870_1535430# diff_869950_1347470# GND GND efet w=18415 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2646 GND diff_869950_1347470# diff_1729740_1228090# GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2647 diff_1790700_1535430# diff_869950_1347470# GND GND efet w=18415 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2648 diff_2439670_1344930# diff_2439670_1344930# diff_2439670_1344930# GND efet w=3175 l=3175
+ ad=2.75806e+08 pd=83820 as=0 ps=0 
M2649 diff_2439670_1344930# diff_2439670_1344930# diff_2439670_1344930# GND efet w=1905 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2650 diff_2080260_1351280# diff_2075180_1344930# GND GND efet w=33020 l=7620
+ ad=2.02742e+09 pd=513080 as=0 ps=0 
M2651 GND diff_2075180_1344930# diff_2128520_1299210# GND efet w=34290 l=7620
+ ad=0 pd=0 as=-1.94497e+09 ps=530860 
M2652 diff_2439670_1344930# Vdd Vdd GND efet w=9525 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2653 GND diff_889000_1079500# diff_1002030_1186180# GND efet w=16510 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2654 GND diff_889000_1079500# diff_1064260_1535430# GND efet w=17780 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2655 diff_1292860_1226820# diff_889000_1079500# GND GND efet w=17145 l=9525
+ ad=0 pd=0 as=0 ps=0 
M2656 diff_1355090_1535430# diff_889000_1079500# GND GND efet w=17145 l=9525
+ ad=0 pd=0 as=0 ps=0 
M2657 GND diff_889000_1079500# diff_1584960_1226820# GND efet w=17780 l=10160
+ ad=0 pd=0 as=0 ps=0 
M2658 diff_1645920_1535430# diff_889000_1079500# GND GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2659 diff_1861820_1186180# diff_889000_1079500# GND GND efet w=17145 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2660 diff_1926590_1210310# diff_889000_1079500# GND GND efet w=16510 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2661 GND diff_139700_2962910# diff_172720_1316990# GND efet w=38100 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2662 diff_857250_1226820# diff_869950_1299210# GND GND efet w=16510 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2663 diff_1148080_1228090# diff_869950_1299210# GND GND efet w=18415 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2664 diff_1002030_1186180# diff_869950_1299210# GND GND efet w=16510 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2665 GND diff_869950_1299210# diff_1292860_1226820# GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2666 GND diff_2089150_1318260# diff_2080260_1351280# GND efet w=20320 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2667 GND diff_2089150_1318260# diff_2172970_1249680# GND efet w=20320 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2668 diff_2471420_1322070# Vdd Vdd GND efet w=11430 l=20320
+ ad=9.91934e+08 pd=193040 as=0 ps=0 
M2669 diff_1438910_1226820# diff_869950_1299210# GND GND efet w=16510 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2670 diff_1584960_1226820# diff_869950_1299210# GND GND efet w=19685 l=10160
+ ad=0 pd=0 as=0 ps=0 
M2671 diff_1729740_1228090# diff_869950_1299210# GND GND efet w=20320 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2672 Vdd Vdd Vdd GND efet w=1270 l=6985
+ ad=0 pd=0 as=0 ps=0 
M2673 Vdd Vdd Vdd GND efet w=4445 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2674 Vdd Vdd diff_172720_1316990# GND efet w=9525 l=38735
+ ad=0 pd=0 as=0 ps=0 
M2675 diff_1064260_1535430# diff_934720_1277620# GND GND efet w=18415 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2676 diff_1209040_1535430# diff_934720_1277620# GND GND efet w=19050 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2677 GND diff_869950_1299210# diff_1861820_1186180# GND efet w=17145 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2678 diff_2471420_1322070# clk2 diff_2475230_1280160# GND efet w=76200 l=7620
+ ad=0 pd=0 as=1.56935e+09 ps=276860 
M2679 GND diff_2443480_1254760# diff_2475230_1280160# GND efet w=119380 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2680 diff_2002790_1228090# diff_1998980_1291590# GND GND efet w=34290 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2681 diff_2128520_1299210# diff_1998980_1291590# GND GND efet w=34290 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2682 diff_1645920_1535430# diff_934720_1277620# GND GND efet w=17780 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2683 GND diff_934720_1277620# diff_918210_1536700# GND efet w=16510 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2684 GND diff_934720_1277620# diff_1355090_1535430# GND efet w=16510 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2685 GND diff_934720_1277620# diff_1499870_1535430# GND efet w=17145 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2686 diff_1790700_1535430# diff_934720_1277620# GND GND efet w=17145 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2687 diff_1926590_1210310# diff_934720_1277620# GND GND efet w=16510 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2688 diff_92710_2421890# diff_232410_1165860# GND GND efet w=69850 l=7620
+ ad=1.59677e+09 pd=185420 as=0 ps=0 
M2689 Vdd diff_262890_1151890# diff_92710_2421890# GND efet w=73660 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2690 diff_546100_1388110# diff_546100_1416050# GND GND efet w=20320 l=7620
+ ad=9.25805e+08 pd=152400 as=0 ps=0 
M2691 Vdd Vdd diff_546100_1388110# GND efet w=12065 l=50165
+ ad=0 pd=0 as=0 ps=0 
M2692 diff_546100_1388110# diff_599440_977900# diff_608330_1151890# GND efet w=8890 l=7620
+ ad=0 pd=0 as=7.4516e+08 ps=172720 
M2693 diff_857250_1226820# diff_855980_1183640# diff_857250_1226820# GND efet w=34290 l=50800
+ ad=0 pd=0 as=0 ps=0 
M2694 diff_232410_1165860# diff_232410_1165860# diff_232410_1165860# GND efet w=2540 l=7620
+ ad=2.2258e+08 pd=66040 as=0 ps=0 
M2695 diff_232410_1165860# diff_232410_1165860# diff_232410_1165860# GND efet w=1270 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2696 diff_262890_1151890# diff_262890_1151890# diff_262890_1151890# GND efet w=2540 l=5715
+ ad=2.3387e+08 pd=71120 as=0 ps=0 
M2697 diff_262890_1151890# diff_262890_1151890# diff_262890_1151890# GND efet w=2540 l=6985
+ ad=0 pd=0 as=0 ps=0 
M2698 diff_369570_1160780# diff_214630_541020# Vdd GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2699 diff_546100_1416050# diff_608330_1151890# GND GND efet w=34290 l=7620
+ ad=1.28064e+09 pd=243840 as=0 ps=0 
M2700 Vdd Vdd diff_546100_1416050# GND efet w=11430 l=49530
+ ad=0 pd=0 as=0 ps=0 
M2701 diff_918210_1536700# diff_920750_1167130# diff_918210_1536700# GND efet w=33020 l=52070
+ ad=0 pd=0 as=0 ps=0 
M2702 diff_232410_1165860# diff_234950_1145540# diff_237490_1127760# GND efet w=15875 l=6985
+ ad=0 pd=0 as=1.2129e+09 ps=223520 
M2703 diff_262890_1151890# diff_234950_1145540# diff_232410_1049020# GND efet w=15240 l=8890
+ ad=0 pd=0 as=9.14514e+08 ps=193040 
M2704 diff_608330_1151890# diff_594360_1112520# diff_369570_1160780# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2705 diff_608330_1151890# diff_608330_1151890# diff_608330_1151890# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M2706 diff_608330_1151890# diff_608330_1151890# diff_608330_1151890# GND efet w=1905 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2707 diff_855980_1183640# diff_855980_1183640# diff_855980_1183640# GND efet w=3175 l=3175
+ ad=2.16129e+08 pd=73660 as=0 ps=0 
M2708 diff_855980_1183640# diff_855980_1183640# diff_855980_1183640# GND efet w=1905 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2709 diff_857250_1226820# diff_855980_1183640# Vdd GND efet w=8890 l=39370
+ ad=0 pd=0 as=0 ps=0 
M2710 diff_918210_1536700# diff_920750_1167130# Vdd GND efet w=8890 l=39370
+ ad=0 pd=0 as=0 ps=0 
M2711 diff_920750_1167130# diff_920750_1167130# diff_920750_1167130# GND efet w=3175 l=3175
+ ad=2.19354e+08 pd=73660 as=0 ps=0 
M2712 diff_855980_1183640# Vdd Vdd GND efet w=7620 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2713 diff_237490_1127760# diff_232410_1049020# GND GND efet w=53340 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2714 diff_266700_2927350# diff_214630_541020# Vdd GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2715 diff_608330_1127760# diff_594360_1112520# diff_266700_2927350# GND efet w=13970 l=7620
+ ad=7.03224e+08 pd=172720 as=0 ps=0 
M2716 diff_608330_1127760# diff_608330_1127760# diff_608330_1127760# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M2717 diff_608330_1127760# diff_608330_1127760# diff_608330_1127760# GND efet w=2540 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2718 diff_920750_1167130# diff_920750_1167130# diff_920750_1167130# GND efet w=1905 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2719 diff_920750_1167130# Vdd Vdd GND efet w=8890 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2720 Vdd Vdd diff_889000_1079500# GND efet w=10795 l=30480
+ ad=0 pd=0 as=-1.77078e+09 ps=670560 
M2721 Vdd Vdd diff_237490_1127760# GND efet w=11430 l=20320
+ ad=0 pd=0 as=0 ps=0 
M2722 diff_243840_2250440# diff_214630_541020# Vdd GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2723 diff_546100_1341120# diff_608330_1127760# GND GND efet w=34290 l=7620
+ ad=1.28064e+09 pd=238760 as=0 ps=0 
M2724 Vdd Vdd diff_546100_1341120# GND efet w=11430 l=49530
+ ad=0 pd=0 as=0 ps=0 
M2725 GND diff_872490_1087120# diff_889000_1079500# GND efet w=52705 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2726 diff_1002030_1186180# diff_1003300_1182370# diff_1002030_1186180# GND efet w=53975 l=29210
+ ad=0 pd=0 as=0 ps=0 
M2727 diff_1064260_1535430# diff_1066800_1167130# diff_1064260_1535430# GND efet w=32385 l=50165
+ ad=0 pd=0 as=0 ps=0 
M2728 diff_1003300_1182370# diff_1003300_1182370# diff_1003300_1182370# GND efet w=3175 l=3175
+ ad=2.27419e+08 pd=81280 as=0 ps=0 
M2729 diff_1003300_1182370# diff_1003300_1182370# diff_1003300_1182370# GND efet w=2540 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2730 diff_1002030_1186180# diff_1003300_1182370# Vdd GND efet w=8890 l=39370
+ ad=0 pd=0 as=0 ps=0 
M2731 diff_1064260_1535430# diff_1066800_1167130# Vdd GND efet w=8890 l=39370
+ ad=0 pd=0 as=0 ps=0 
M2732 diff_1066800_1167130# diff_1066800_1167130# diff_1066800_1167130# GND efet w=3175 l=3175
+ ad=2.30645e+08 pd=81280 as=0 ps=0 
M2733 diff_1066800_1167130# diff_1066800_1167130# diff_1066800_1167130# GND efet w=2540 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2734 diff_1003300_1182370# Vdd Vdd GND efet w=9525 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2735 diff_1066800_1167130# Vdd Vdd GND efet w=8890 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2736 diff_869950_1347470# Vdd Vdd GND efet w=8890 l=33020
+ ad=1.67419e+09 pd=439420 as=0 ps=0 
M2737 diff_1148080_1228090# diff_1146810_1183640# diff_1148080_1228090# GND efet w=32385 l=50800
+ ad=0 pd=0 as=0 ps=0 
M2738 diff_1209040_1535430# diff_1211580_1167130# diff_1209040_1535430# GND efet w=33020 l=49530
+ ad=0 pd=0 as=0 ps=0 
M2739 diff_1146810_1183640# diff_1146810_1183640# diff_1146810_1183640# GND efet w=3175 l=3175
+ ad=2.12903e+08 pd=76200 as=0 ps=0 
M2740 diff_1146810_1183640# diff_1146810_1183640# diff_1146810_1183640# GND efet w=1905 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2741 diff_1148080_1228090# diff_1146810_1183640# Vdd GND efet w=8890 l=39370
+ ad=0 pd=0 as=0 ps=0 
M2742 diff_1209040_1535430# diff_1211580_1167130# Vdd GND efet w=8890 l=39370
+ ad=0 pd=0 as=0 ps=0 
M2743 diff_1211580_1167130# diff_1211580_1167130# diff_1211580_1167130# GND efet w=3175 l=3175
+ ad=2.09677e+08 pd=73660 as=0 ps=0 
M2744 diff_1146810_1183640# Vdd Vdd GND efet w=8890 l=9525
+ ad=0 pd=0 as=0 ps=0 
M2745 diff_1211580_1167130# diff_1211580_1167130# diff_1211580_1167130# GND efet w=1905 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2746 diff_1211580_1167130# Vdd Vdd GND efet w=9525 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2747 diff_1292860_1226820# diff_1292860_1186180# diff_1292860_1226820# GND efet w=34290 l=35560
+ ad=0 pd=0 as=0 ps=0 
M2748 diff_1355090_1535430# diff_1356360_1168400# diff_1355090_1535430# GND efet w=33655 l=29210
+ ad=0 pd=0 as=0 ps=0 
M2749 diff_1438910_1226820# diff_1437640_1181100# diff_1438910_1226820# GND efet w=33655 l=49530
+ ad=0 pd=0 as=0 ps=0 
M2750 diff_1292860_1186180# diff_1292860_1186180# diff_1292860_1186180# GND efet w=3175 l=3175
+ ad=2.20967e+08 pd=76200 as=0 ps=0 
M2751 diff_1292860_1186180# diff_1292860_1186180# diff_1292860_1186180# GND efet w=1905 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2752 diff_1292860_1226820# diff_1292860_1186180# Vdd GND efet w=8890 l=39370
+ ad=0 pd=0 as=0 ps=0 
M2753 diff_1355090_1535430# diff_1356360_1168400# Vdd GND efet w=8890 l=39370
+ ad=0 pd=0 as=0 ps=0 
M2754 diff_1356360_1168400# diff_1356360_1168400# diff_1356360_1168400# GND efet w=3175 l=3175
+ ad=2.27419e+08 pd=76200 as=0 ps=0 
M2755 diff_1356360_1168400# diff_1356360_1168400# diff_1356360_1168400# GND efet w=1905 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2756 diff_1292860_1186180# Vdd Vdd GND efet w=8890 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2757 diff_1356360_1168400# Vdd Vdd GND efet w=8890 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2758 diff_1499870_1535430# diff_1502410_1167130# diff_1499870_1535430# GND efet w=33655 l=50165
+ ad=0 pd=0 as=0 ps=0 
M2759 diff_1437640_1181100# diff_1437640_1181100# diff_1437640_1181100# GND efet w=2540 l=3810
+ ad=2.08064e+08 pd=71120 as=0 ps=0 
M2760 diff_1437640_1181100# diff_1437640_1181100# diff_1437640_1181100# GND efet w=1905 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2761 diff_1438910_1226820# diff_1437640_1181100# Vdd GND efet w=8890 l=39370
+ ad=0 pd=0 as=0 ps=0 
M2762 diff_1499870_1535430# diff_1502410_1167130# Vdd GND efet w=8890 l=39370
+ ad=0 pd=0 as=0 ps=0 
M2763 GND diff_1795780_1076960# diff_2002790_1228090# GND efet w=20320 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2764 GND diff_1795780_1076960# diff_2080260_1351280# GND efet w=20320 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2765 GND diff_1795780_1076960# diff_2128520_1299210# GND efet w=22860 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2766 GND diff_1795780_1076960# diff_2172970_1249680# GND efet w=20320 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2767 diff_1584960_1226820# diff_1583690_1181100# diff_1584960_1226820# GND efet w=33655 l=49530
+ ad=0 pd=0 as=0 ps=0 
M2768 diff_1645920_1535430# diff_1647190_1168400# diff_1645920_1535430# GND efet w=52070 l=29210
+ ad=0 pd=0 as=0 ps=0 
M2769 diff_1502410_1167130# diff_1502410_1167130# diff_1502410_1167130# GND efet w=3175 l=3175
+ ad=2.09677e+08 pd=71120 as=0 ps=0 
M2770 diff_1437640_1181100# Vdd Vdd GND efet w=8255 l=9525
+ ad=0 pd=0 as=0 ps=0 
M2771 Vdd Vdd diff_232410_1049020# GND efet w=10795 l=20955
+ ad=0 pd=0 as=0 ps=0 
M2772 diff_232410_1049020# diff_232410_996950# GND GND efet w=54610 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2773 diff_245110_1436370# diff_214630_541020# Vdd GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2774 Vdd Vdd diff_546100_1313180# GND efet w=10160 l=49530
+ ad=0 pd=0 as=1.15e+09 ps=269240 
M2775 GND diff_889000_1079500# diff_869950_1347470# GND efet w=27940 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2776 diff_872490_1417320# diff_1192530_1032510# GND GND efet w=40640 l=8890
+ ad=1.76451e+09 pd=426720 as=0 ps=0 
M2777 Vdd Vdd diff_872490_1417320# GND efet w=8890 l=31750
+ ad=0 pd=0 as=0 ps=0 
M2778 diff_1377950_1109980# Vdd Vdd GND efet w=8890 l=33020
+ ad=1.67258e+09 pd=454660 as=0 ps=0 
M2779 diff_1502410_1167130# diff_1502410_1167130# diff_1502410_1167130# GND efet w=1905 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2780 diff_1502410_1167130# Vdd Vdd GND efet w=8890 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2781 diff_1583690_1181100# diff_1583690_1181100# diff_1583690_1181100# GND efet w=3175 l=3175
+ ad=2.32258e+08 pd=78740 as=0 ps=0 
M2782 diff_1583690_1181100# diff_1583690_1181100# diff_1583690_1181100# GND efet w=2540 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2783 diff_1584960_1226820# diff_1583690_1181100# Vdd GND efet w=8890 l=39370
+ ad=0 pd=0 as=0 ps=0 
M2784 diff_1645920_1535430# diff_1647190_1168400# Vdd GND efet w=8890 l=39370
+ ad=0 pd=0 as=0 ps=0 
M2785 diff_1647190_1168400# diff_1647190_1168400# diff_1647190_1168400# GND efet w=1905 l=4445
+ ad=2.30645e+08 pd=78740 as=0 ps=0 
M2786 diff_1583690_1181100# Vdd Vdd GND efet w=10160 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2787 diff_1647190_1168400# diff_1647190_1168400# diff_1647190_1168400# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M2788 diff_1647190_1168400# Vdd Vdd GND efet w=10160 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2789 diff_1377950_1109980# diff_872490_1417320# GND GND efet w=26670 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2790 diff_1160780_1371600# diff_1483360_1032510# GND GND efet w=40640 l=8890
+ ad=1.78548e+09 pd=449580 as=0 ps=0 
M2791 Vdd Vdd diff_1160780_1371600# GND efet w=8890 l=33020
+ ad=0 pd=0 as=0 ps=0 
M2792 diff_869950_1397000# Vdd Vdd GND efet w=8255 l=32385
+ ad=1.55645e+09 pd=424180 as=0 ps=0 
M2793 diff_1729740_1228090# diff_1728470_1183640# diff_1729740_1228090# GND efet w=32385 l=50800
+ ad=0 pd=0 as=0 ps=0 
M2794 diff_1790700_1535430# diff_1793240_1167130# diff_1790700_1535430# GND efet w=51435 l=26035
+ ad=0 pd=0 as=0 ps=0 
M2795 diff_1728470_1183640# diff_1728470_1183640# diff_1728470_1183640# GND efet w=2540 l=3810
+ ad=2.1129e+08 pd=71120 as=0 ps=0 
M2796 diff_1728470_1183640# diff_1728470_1183640# diff_1728470_1183640# GND efet w=1905 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2797 diff_1729740_1228090# diff_1728470_1183640# Vdd GND efet w=8890 l=39370
+ ad=0 pd=0 as=0 ps=0 
M2798 diff_1790700_1535430# diff_1793240_1167130# Vdd GND efet w=8890 l=39370
+ ad=0 pd=0 as=0 ps=0 
M2799 diff_1793240_1167130# diff_1793240_1167130# diff_1793240_1167130# GND efet w=2540 l=3175
+ ad=2.25806e+08 pd=78740 as=0 ps=0 
M2800 diff_1728470_1183640# Vdd Vdd GND efet w=8890 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2801 diff_1793240_1167130# diff_1793240_1167130# diff_1793240_1167130# GND efet w=3175 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2802 diff_1861820_1186180# diff_1869440_1156970# diff_1861820_1186180# GND efet w=50800 l=25400
+ ad=0 pd=0 as=0 ps=0 
M2803 diff_1926590_1210310# diff_1925320_1167130# diff_1926590_1210310# GND efet w=51435 l=26035
+ ad=0 pd=0 as=0 ps=0 
M2804 diff_1869440_1156970# diff_1869440_1156970# diff_1869440_1156970# GND efet w=2540 l=3810
+ ad=2.48387e+08 pd=78740 as=0 ps=0 
M2805 diff_1869440_1156970# diff_1869440_1156970# diff_1869440_1156970# GND efet w=2540 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2806 diff_1861820_1186180# diff_1869440_1156970# Vdd GND efet w=8890 l=39370
+ ad=0 pd=0 as=0 ps=0 
M2807 diff_1926590_1210310# diff_1925320_1167130# Vdd GND efet w=8890 l=39370
+ ad=0 pd=0 as=0 ps=0 
M2808 diff_1925320_1167130# diff_1925320_1167130# diff_1925320_1167130# GND efet w=2540 l=3175
+ ad=2.27419e+08 pd=78740 as=0 ps=0 
M2809 diff_1793240_1167130# Vdd Vdd GND efet w=9525 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2810 Vdd Vdd Vdd GND efet w=3810 l=10160
+ ad=0 pd=0 as=0 ps=0 
M2811 Vdd Vdd Vdd GND efet w=3810 l=10160
+ ad=0 pd=0 as=0 ps=0 
M2812 Vdd Vdd Vdd GND efet w=6985 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2813 Vdd Vdd Vdd GND efet w=3810 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2814 Vdd Vdd diff_869950_1299210# GND efet w=10160 l=33020
+ ad=0 pd=0 as=5.7258e+08 ps=157480 
M2815 diff_869950_1397000# diff_1160780_1371600# GND GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2816 diff_1869440_1156970# Vdd Vdd GND efet w=8890 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2817 diff_1925320_1167130# diff_1925320_1167130# diff_1925320_1167130# GND efet w=3175 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2818 diff_1925320_1167130# Vdd Vdd GND efet w=9525 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2819 Vdd Vdd Vdd GND efet w=1905 l=6985
+ ad=0 pd=0 as=0 ps=0 
M2820 Vdd Vdd Vdd GND efet w=3175 l=9525
+ ad=0 pd=0 as=0 ps=0 
M2821 Vdd Vdd Vdd GND efet w=1905 l=5715
+ ad=0 pd=0 as=0 ps=0 
M2822 Vdd Vdd Vdd GND efet w=6985 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2823 diff_869950_1299210# diff_869950_1299210# diff_869950_1299210# GND efet w=2540 l=3175
+ ad=0 pd=0 as=0 ps=0 
M2824 diff_869950_1299210# diff_869950_1299210# diff_869950_1299210# GND efet w=3175 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2825 Vdd Vdd diff_934720_1277620# GND efet w=8890 l=31750
+ ad=0 pd=0 as=5.35483e+08 ps=149860 
M2826 diff_2002790_1228090# diff_2000250_1186180# diff_2002790_1228090# GND efet w=33020 l=52070
+ ad=0 pd=0 as=0 ps=0 
M2827 diff_2000250_1186180# diff_2000250_1186180# diff_2000250_1186180# GND efet w=3175 l=3175
+ ad=2.2258e+08 pd=78740 as=0 ps=0 
M2828 diff_2000250_1186180# diff_2000250_1186180# diff_2000250_1186180# GND efet w=3175 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2829 diff_2002790_1228090# diff_2000250_1186180# Vdd GND efet w=8890 l=39370
+ ad=0 pd=0 as=0 ps=0 
M2830 diff_2000250_1186180# Vdd Vdd GND efet w=8890 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2831 diff_2443480_1254760# Vdd Vdd GND efet w=11430 l=29210
+ ad=5.77418e+08 pd=119380 as=0 ps=0 
M2832 GND diff_2463800_1235710# diff_2443480_1254760# GND efet w=41275 l=6985
+ ad=0 pd=0 as=0 ps=0 
M2833 diff_2080260_1351280# diff_2085340_1167130# diff_2080260_1351280# GND efet w=56515 l=27305
+ ad=0 pd=0 as=0 ps=0 
M2834 diff_2080260_1351280# diff_2085340_1167130# Vdd GND efet w=8890 l=40640
+ ad=0 pd=0 as=0 ps=0 
M2835 diff_2128520_1299210# diff_2138680_1156970# diff_2128520_1299210# GND efet w=53340 l=29845
+ ad=0 pd=0 as=0 ps=0 
M2836 diff_2463800_1235710# diff_2463800_1235710# diff_2463800_1235710# GND efet w=1270 l=5080
+ ad=6.38708e+08 pd=116840 as=0 ps=0 
M2837 diff_2085340_1167130# diff_2085340_1167130# diff_2085340_1167130# GND efet w=2540 l=3810
+ ad=2.04838e+08 pd=73660 as=0 ps=0 
M2838 diff_2085340_1167130# diff_2085340_1167130# diff_2085340_1167130# GND efet w=2540 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2839 diff_1795780_1076960# Vdd Vdd GND efet w=9525 l=33655
+ ad=9.59676e+08 pd=220980 as=0 ps=0 
M2840 diff_934720_1277620# diff_934720_1277620# diff_934720_1277620# GND efet w=1905 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2841 diff_934720_1277620# diff_934720_1277620# diff_934720_1277620# GND efet w=2540 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2842 diff_2138680_1156970# diff_2138680_1156970# diff_2138680_1156970# GND efet w=2540 l=3810
+ ad=2.09677e+08 pd=71120 as=0 ps=0 
M2843 diff_2138680_1156970# diff_2138680_1156970# diff_2138680_1156970# GND efet w=1905 l=5715
+ ad=0 pd=0 as=0 ps=0 
M2844 diff_2128520_1299210# diff_2138680_1156970# Vdd GND efet w=8890 l=39370
+ ad=0 pd=0 as=0 ps=0 
M2845 diff_2085340_1167130# Vdd Vdd GND efet w=7620 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2846 diff_2138680_1156970# Vdd Vdd GND efet w=7620 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2847 Vdd Vdd Vdd GND efet w=6985 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2848 Vdd Vdd Vdd GND efet w=3175 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2849 Vdd Vdd Vdd GND efet w=6985 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2850 diff_2089150_1318260# diff_2089150_1318260# diff_2089150_1318260# GND efet w=3810 l=6350
+ ad=1.12419e+09 pd=208280 as=0 ps=0 
M2851 Vdd Vdd Vdd GND efet w=3810 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2852 Vdd Vdd diff_2089150_1318260# GND efet w=8890 l=38100
+ ad=0 pd=0 as=0 ps=0 
M2853 diff_2089150_1318260# diff_1998980_1291590# GND GND efet w=44450 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2854 diff_2089150_1318260# diff_2089150_1318260# diff_2089150_1318260# GND efet w=2540 l=2540
+ ad=0 pd=0 as=0 ps=0 
M2855 diff_1795780_1076960# diff_1795780_1076960# diff_1795780_1076960# GND efet w=1905 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2856 diff_1795780_1076960# diff_1795780_1076960# diff_1795780_1076960# GND efet w=3175 l=5080
+ ad=0 pd=0 as=0 ps=0 
M2857 diff_2012950_1370330# Vdd Vdd GND efet w=9525 l=38735
+ ad=7.27418e+08 pd=149860 as=0 ps=0 
M2858 diff_2012950_1370330# diff_2012950_1370330# diff_2012950_1370330# GND efet w=3810 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2859 diff_2012950_1370330# diff_2012950_1370330# diff_2012950_1370330# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M2860 diff_1795780_1076960# diff_1988820_1080770# GND GND efet w=49530 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2861 diff_608330_1127760# diff_599440_977900# diff_546100_1313180# GND efet w=8890 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2862 diff_546100_1313180# diff_546100_1341120# GND GND efet w=20320 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2863 diff_869950_1299210# diff_1795780_1076960# diff_1799590_1065530# GND efet w=52070 l=7620
+ ad=0 pd=0 as=5.29031e+08 ps=124460 
M2864 diff_934720_1277620# diff_1795780_1076960# diff_1882140_1065530# GND efet w=52070 l=7620
+ ad=0 pd=0 as=7.04837e+08 ps=170180 
M2865 GND diff_2075180_1344930# diff_2012950_1370330# GND efet w=39370 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2866 diff_2463800_1235710# diff_2463800_1235710# diff_2463800_1235710# GND efet w=3810 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2867 diff_2463800_1235710# Vdd Vdd GND efet w=9525 l=61595
+ ad=0 pd=0 as=0 ps=0 
M2868 diff_2534920_1196340# diff_1897380_186690# diff_2463800_1235710# GND efet w=27940 l=7620
+ ad=9.99998e+08 pd=195580 as=0 ps=0 
M2869 diff_2534920_1196340# diff_932180_1050290# GND GND efet w=29210 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2870 GND diff_897890_1024890# diff_2534920_1196340# GND efet w=31750 l=6985
+ ad=0 pd=0 as=0 ps=0 
M2871 diff_284480_472440# clk1 diff_2578100_1071880# GND efet w=15875 l=6985
+ ad=1.21613e+09 pd=251460 as=2.85483e+08 ps=68580 
M2872 diff_1877060_1057910# diff_1877060_1057910# diff_1877060_1057910# GND efet w=1905 l=3810
+ ad=9.62901e+08 pd=213360 as=0 ps=0 
M2873 diff_1988820_1080770# diff_1988820_1080770# diff_1988820_1080770# GND efet w=1905 l=4445
+ ad=9.99998e+08 pd=213360 as=0 ps=0 
M2874 diff_1998980_1291590# diff_1998980_1291590# diff_1998980_1291590# GND efet w=1905 l=4445
+ ad=9.48385e+08 pd=205740 as=0 ps=0 
M2875 diff_1877060_1057910# diff_1877060_1057910# diff_1877060_1057910# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M2876 diff_1988820_1080770# diff_1988820_1080770# diff_1988820_1080770# GND efet w=2540 l=2540
+ ad=0 pd=0 as=0 ps=0 
M2877 diff_1998980_1291590# diff_1998980_1291590# diff_1998980_1291590# GND efet w=2540 l=2540
+ ad=0 pd=0 as=0 ps=0 
M2878 diff_932180_1002030# diff_932180_1050290# diff_872490_1087120# GND efet w=13970 l=7620
+ ad=1.75322e+09 pd=327660 as=9.24192e+08 ps=177800 
M2879 diff_1192530_1032510# diff_932180_1050290# diff_1223010_990600# GND efet w=15240 l=7620
+ ad=1.14516e+09 pd=220980 as=1.63709e+09 ps=330200 
M2880 diff_1799590_1065530# diff_934720_1277620# GND GND efet w=53975 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2881 diff_1483360_1032510# diff_932180_1050290# diff_1513840_989330# GND efet w=13970 l=7620
+ ad=1.08709e+09 pd=218440 as=1.61613e+09 ps=325120 
M2882 diff_1882140_1065530# diff_1877060_1057910# GND GND efet w=80010 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2883 diff_872490_1087120# diff_897890_1024890# diff_812800_871220# GND efet w=13970 l=7620
+ ad=0 pd=0 as=1.45645e+09 ps=353060 
M2884 diff_594360_1112520# diff_599440_977900# GND GND efet w=15240 l=7620
+ ad=4.8387e+08 pd=114300 as=0 ps=0 
M2885 Vdd Vdd diff_594360_1112520# GND efet w=8890 l=62230
+ ad=0 pd=0 as=0 ps=0 
M2886 diff_1192530_1032510# diff_897890_1024890# diff_1103630_871220# GND efet w=13970 l=7620
+ ad=0 pd=0 as=1.47096e+09 ps=365760 
M2887 diff_1877060_1057910# diff_932180_1050290# diff_1888490_857250# GND efet w=15240 l=7620
+ ad=0 pd=0 as=1.74193e+09 ps=337820 
M2888 GND diff_2578100_1071880# diff_897890_1024890# GND efet w=55880 l=6350
+ ad=0 pd=0 as=1.95967e+09 ps=383540 
M2889 diff_2075180_1344930# diff_2075180_1344930# diff_2075180_1344930# GND efet w=3810 l=8890
+ ad=1.16935e+09 pd=233680 as=0 ps=0 
M2890 diff_1988820_1080770# diff_932180_1050290# diff_1790700_659130# GND efet w=13970 l=7620
+ ad=0 pd=0 as=1.41129e+09 ps=309880 
M2891 diff_1483360_1032510# diff_897890_1024890# diff_1400810_873760# GND efet w=14605 l=7620
+ ad=0 pd=0 as=9.91934e+08 ps=271780 
M2892 diff_1103630_871220# diff_1103630_871220# diff_1103630_871220# GND efet w=3175 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2893 diff_1103630_871220# diff_1103630_871220# diff_1103630_871220# GND efet w=1270 l=5080
+ ad=0 pd=0 as=0 ps=0 
M2894 Vdd Vdd diff_251460_913130# GND efet w=8890 l=10160
+ ad=0 pd=0 as=1.96774e+08 ps=68580 
M2895 diff_251460_913130# diff_251460_913130# diff_251460_913130# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M2896 diff_251460_913130# diff_251460_913130# diff_251460_913130# GND efet w=1905 l=5715
+ ad=0 pd=0 as=0 ps=0 
M2897 Vdd diff_251460_913130# diff_234950_1145540# GND efet w=10160 l=10160
+ ad=0 pd=0 as=1.61774e+09 ps=266700 
M2898 diff_234950_1145540# diff_251460_913130# diff_234950_1145540# GND efet w=38735 l=28575
+ ad=0 pd=0 as=0 ps=0 
M2899 diff_1223010_990600# diff_1223010_990600# diff_1223010_990600# GND efet w=2540 l=5080
+ ad=0 pd=0 as=0 ps=0 
M2900 diff_1223010_990600# diff_1223010_990600# diff_1223010_990600# GND efet w=1270 l=5080
+ ad=0 pd=0 as=0 ps=0 
M2901 diff_1877060_1057910# diff_897890_1024890# diff_1691640_873760# GND efet w=13970 l=7620
+ ad=0 pd=0 as=1.03064e+09 ps=276860 
M2902 diff_1400810_873760# diff_1400810_873760# diff_1400810_873760# GND efet w=3175 l=6985
+ ad=0 pd=0 as=0 ps=0 
M2903 diff_1400810_873760# diff_1400810_873760# diff_1400810_873760# GND efet w=1270 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2904 diff_234950_1145540# clk2 GND GND efet w=53975 l=6985
+ ad=0 pd=0 as=0 ps=0 
M2905 Vdd Vdd diff_812800_871220# GND efet w=11430 l=25400
+ ad=0 pd=0 as=0 ps=0 
M2906 diff_808990_863600# Vdd Vdd GND efet w=7620 l=48260
+ ad=8.19353e+08 pd=200660 as=0 ps=0 
M2907 diff_812800_871220# diff_808990_863600# GND GND efet w=35560 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2908 diff_808990_863600# diff_808990_863600# diff_808990_863600# GND efet w=2540 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2909 diff_808990_863600# diff_808990_863600# diff_808990_863600# GND efet w=1905 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2910 Vdd Vdd diff_887730_825500# GND efet w=8890 l=60960
+ ad=0 pd=0 as=7.04837e+08 ps=160020 
M2911 diff_820420_830580# Vdd Vdd GND efet w=7620 l=48260
+ ad=8.49998e+08 pd=190500 as=0 ps=0 
M2912 diff_820420_830580# diff_820420_830580# diff_820420_830580# GND efet w=2540 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2913 diff_820420_830580# diff_820420_830580# diff_820420_830580# GND efet w=2540 l=5080
+ ad=0 pd=0 as=0 ps=0 
M2914 GND diff_820420_830580# diff_887730_825500# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2915 GND diff_408940_681990# diff_575310_779780# GND efet w=15240 l=7620
+ ad=0 pd=0 as=9.11289e+08 ps=223520 
M2916 GND diff_820420_830580# diff_808990_863600# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2917 diff_575310_779780# diff_575310_779780# diff_575310_779780# GND efet w=6985 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2918 diff_575310_779780# diff_575310_779780# diff_575310_779780# GND efet w=3810 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2919 diff_812800_871220# diff_812800_871220# diff_812800_871220# GND efet w=3175 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2920 diff_812800_871220# diff_812800_871220# diff_812800_871220# GND efet w=2540 l=6985
+ ad=0 pd=0 as=0 ps=0 
M2921 diff_887730_825500# diff_408940_681990# diff_808990_749300# GND efet w=15875 l=8255
+ ad=0 pd=0 as=4.99999e+08 ps=96520 
M2922 Vdd Vdd diff_932180_1002030# GND efet w=11430 l=39370
+ ad=0 pd=0 as=0 ps=0 
M2923 Vdd Vdd diff_1049020_786130# GND efet w=8890 l=60960
+ ad=0 pd=0 as=5.51612e+08 ps=154940 
M2924 Vdd Vdd diff_1103630_871220# GND efet w=12065 l=26035
+ ad=0 pd=0 as=0 ps=0 
M2925 diff_932180_1002030# diff_932180_1002030# diff_932180_1002030# GND efet w=1905 l=5715
+ ad=0 pd=0 as=0 ps=0 
M2926 GND diff_808990_863600# diff_820420_830580# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2927 diff_932180_1002030# diff_932180_1002030# diff_932180_1002030# GND efet w=3810 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2928 diff_1049020_786130# diff_1049020_786130# diff_1049020_786130# GND efet w=1905 l=6985
+ ad=0 pd=0 as=0 ps=0 
M2929 diff_1049020_786130# diff_1049020_786130# diff_1049020_786130# GND efet w=3175 l=5080
+ ad=0 pd=0 as=0 ps=0 
M2930 diff_812800_871220# diff_408940_681990# diff_913130_783590# GND efet w=15240 l=7620
+ ad=0 pd=0 as=5.01612e+08 ps=96520 
M2931 diff_808990_863600# diff_575310_779780# diff_798830_753110# GND efet w=32385 l=8255
+ ad=0 pd=0 as=7.70966e+08 ps=177800 
M2932 diff_400050_777240# clk2 sync GND efet w=8890 l=7620
+ ad=3.12903e+08 pd=83820 as=5.90507e+08 ps=1.06426e+06 
M2933 diff_400050_777240# diff_400050_777240# diff_400050_777240# GND efet w=2540 l=2540
+ ad=0 pd=0 as=0 ps=0 
M2934 diff_400050_777240# diff_400050_777240# diff_400050_777240# GND efet w=1905 l=5080
+ ad=0 pd=0 as=0 ps=0 
M2935 diff_419100_734060# diff_400050_777240# GND GND efet w=33020 l=7620
+ ad=6.99999e+08 pd=139700 as=0 ps=0 
M2936 Vdd Vdd diff_419100_734060# GND efet w=8890 l=60960
+ ad=0 pd=0 as=0 ps=0 
M2937 diff_575310_779780# Vdd Vdd GND efet w=10160 l=62230
+ ad=0 pd=0 as=0 ps=0 
M2938 GND diff_576580_742950# diff_575310_779780# GND efet w=14605 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2939 GND diff_808990_749300# diff_798830_753110# GND efet w=53975 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2940 diff_576580_742950# diff_576580_742950# diff_576580_742950# GND efet w=3175 l=3175
+ ad=5.46773e+08 pd=137160 as=0 ps=0 
M2941 diff_576580_742950# diff_576580_742950# diff_576580_742950# GND efet w=3175 l=6985
+ ad=0 pd=0 as=0 ps=0 
M2942 diff_401320_678180# clk1 diff_419100_734060# GND efet w=9525 l=8255
+ ad=3.90322e+08 pd=96520 as=0 ps=0 
M2943 diff_576580_742950# Vdd Vdd GND efet w=6985 l=57785
+ ad=0 pd=0 as=0 ps=0 
M2944 diff_408940_681990# diff_401320_678180# GND GND efet w=21590 l=7620
+ ad=4.87096e+08 pd=114300 as=0 ps=0 
M2945 diff_576580_742950# diff_419100_734060# GND GND efet w=12700 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2946 Vdd Vdd diff_408940_681990# GND efet w=8890 l=43815
+ ad=0 pd=0 as=0 ps=0 
M2947 diff_408940_681990# clk2 diff_374650_646430# GND efet w=9525 l=6985
+ ad=0 pd=0 as=2.59677e+08 ps=71120 
M2948 GND diff_374650_646430# diff_377190_637540# GND efet w=15875 l=6985
+ ad=0 pd=0 as=6.9516e+08 ps=160020 
M2949 diff_932180_1002030# diff_1005840_731520# diff_1022350_718820# GND efet w=13970 l=8890
+ ad=0 pd=0 as=1.2e+09 ps=261620 
M2950 diff_820420_830580# diff_575310_779780# diff_957580_789940# GND efet w=29210 l=7620
+ ad=0 pd=0 as=8.83869e+08 ps=190500 
M2951 diff_957580_789940# diff_913130_783590# GND GND efet w=54610 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2952 GND diff_1049020_786130# diff_932180_1002030# GND efet w=26670 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2953 diff_1099820_863600# Vdd Vdd GND efet w=7620 l=48260
+ ad=8.48385e+08 pd=205740 as=0 ps=0 
M2954 diff_1103630_871220# diff_1099820_863600# GND GND efet w=35560 l=8890
+ ad=0 pd=0 as=0 ps=0 
M2955 diff_1099820_863600# diff_1099820_863600# diff_1099820_863600# GND efet w=2540 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2956 diff_1099820_863600# diff_1099820_863600# diff_1099820_863600# GND efet w=2540 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2957 Vdd Vdd diff_1178560_825500# GND efet w=8890 l=60960
+ ad=0 pd=0 as=6.77418e+08 ps=160020 
M2958 diff_1111250_830580# Vdd Vdd GND efet w=8255 l=47625
+ ad=8.30644e+08 pd=187960 as=0 ps=0 
M2959 diff_1111250_830580# diff_1111250_830580# diff_1111250_830580# GND efet w=1905 l=6985
+ ad=0 pd=0 as=0 ps=0 
M2960 diff_1111250_830580# diff_1111250_830580# diff_1111250_830580# GND efet w=2540 l=5080
+ ad=0 pd=0 as=0 ps=0 
M2961 GND diff_1111250_830580# diff_1178560_825500# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2962 GND diff_1111250_830580# diff_1099820_863600# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2963 diff_1103630_871220# diff_1103630_871220# diff_1103630_871220# GND efet w=2540 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2964 diff_1103630_871220# diff_1103630_871220# diff_1103630_871220# GND efet w=2540 l=5715
+ ad=0 pd=0 as=0 ps=0 
M2965 diff_1178560_825500# diff_808990_863600# diff_1099820_749300# GND efet w=15875 l=9525
+ ad=0 pd=0 as=4.93547e+08 ps=96520 
M2966 diff_1513840_989330# diff_1513840_989330# diff_1513840_989330# GND efet w=2540 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2967 diff_1691640_873760# diff_1691640_873760# diff_1691640_873760# GND efet w=4445 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2968 diff_1888490_857250# diff_1888490_857250# diff_1888490_857250# GND efet w=2540 l=5080
+ ad=0 pd=0 as=0 ps=0 
M2969 diff_1513840_989330# diff_1513840_989330# diff_1513840_989330# GND efet w=1270 l=5080
+ ad=0 pd=0 as=0 ps=0 
M2970 diff_1691640_873760# diff_1691640_873760# diff_1691640_873760# GND efet w=1905 l=1905
+ ad=0 pd=0 as=0 ps=0 
M2971 diff_1998980_1291590# diff_932180_1050290# diff_1576070_459740# GND efet w=15240 l=7620
+ ad=0 pd=0 as=1.34677e+09 ps=299720 
M2972 Vdd Vdd Vdd GND efet w=1905 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2973 diff_2075180_1344930# diff_2075180_1344930# diff_2075180_1344930# GND efet w=5715 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2974 diff_1988820_1080770# diff_897890_1024890# diff_1982470_873760# GND efet w=15240 l=7620
+ ad=0 pd=0 as=1.11129e+09 ps=289560 
M2975 diff_1998980_1291590# diff_897890_1024890# diff_1103630_871220# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2976 diff_1888490_857250# diff_1888490_857250# diff_1888490_857250# GND efet w=1270 l=5080
+ ad=0 pd=0 as=0 ps=0 
M2977 diff_1982470_873760# diff_1982470_873760# diff_1982470_873760# GND efet w=4445 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2978 diff_1790700_659130# diff_1790700_659130# diff_1790700_659130# GND efet w=3175 l=5080
+ ad=0 pd=0 as=0 ps=0 
M2979 diff_1982470_873760# diff_1982470_873760# diff_1982470_873760# GND efet w=1270 l=5080
+ ad=0 pd=0 as=0 ps=0 
M2980 diff_1790700_659130# diff_1790700_659130# diff_1790700_659130# GND efet w=1270 l=5080
+ ad=0 pd=0 as=0 ps=0 
M2981 Vdd Vdd Vdd GND efet w=3810 l=5715
+ ad=0 pd=0 as=0 ps=0 
M2982 diff_897890_1024890# Vdd Vdd GND efet w=11430 l=20320
+ ad=0 pd=0 as=0 ps=0 
M2983 diff_2075180_1344930# diff_932180_1050290# diff_1677670_457200# GND efet w=13970 l=7620
+ ad=0 pd=0 as=1.3629e+09 ps=307340 
M2984 diff_1576070_459740# diff_1576070_459740# diff_1576070_459740# GND efet w=2540 l=4445
+ ad=0 pd=0 as=0 ps=0 
M2985 diff_2075180_1344930# diff_897890_1024890# diff_812800_871220# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M2986 diff_1223010_990600# Vdd Vdd GND efet w=10795 l=40005
+ ad=0 pd=0 as=0 ps=0 
M2987 Vdd Vdd diff_1339850_786130# GND efet w=8890 l=60960
+ ad=0 pd=0 as=5.51612e+08 ps=154940 
M2988 Vdd Vdd diff_1400810_873760# GND efet w=11430 l=39370
+ ad=0 pd=0 as=0 ps=0 
M2989 diff_1391920_806450# Vdd Vdd GND efet w=7620 l=53340
+ ad=8.35482e+08 pd=210820 as=0 ps=0 
M2990 diff_1223010_990600# diff_1223010_990600# diff_1223010_990600# GND efet w=1905 l=5715
+ ad=0 pd=0 as=0 ps=0 
M2991 GND diff_1099820_863600# diff_1111250_830580# GND efet w=15875 l=8255
+ ad=0 pd=0 as=0 ps=0 
M2992 diff_1223010_990600# diff_1223010_990600# diff_1223010_990600# GND efet w=3810 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2993 diff_1339850_786130# diff_1339850_786130# diff_1339850_786130# GND efet w=1905 l=6985
+ ad=0 pd=0 as=0 ps=0 
M2994 diff_1339850_786130# diff_1339850_786130# diff_1339850_786130# GND efet w=3175 l=3810
+ ad=0 pd=0 as=0 ps=0 
M2995 diff_1103630_871220# diff_808990_863600# diff_1203960_786130# GND efet w=16510 l=7620
+ ad=0 pd=0 as=4.98386e+08 ps=96520 
M2996 diff_1099820_863600# diff_820420_830580# diff_1087120_770890# GND efet w=31115 l=7620
+ ad=0 pd=0 as=9.0645e+08 ps=195580 
M2997 diff_1022350_718820# diff_1022350_718820# diff_1022350_718820# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M2998 diff_1022350_718820# diff_1022350_718820# diff_1022350_718820# GND efet w=1905 l=1905
+ ad=0 pd=0 as=0 ps=0 
M2999 diff_1049020_786130# diff_1022350_718820# GND GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3000 GND diff_1099820_749300# diff_1087120_770890# GND efet w=61595 l=8255
+ ad=0 pd=0 as=0 ps=0 
M3001 diff_1223010_990600# diff_1005840_731520# diff_1313180_713740# GND efet w=13970 l=8255
+ ad=0 pd=0 as=1.24355e+09 ps=271780 
M3002 diff_1111250_830580# diff_820420_830580# diff_1248410_791210# GND efet w=29210 l=7620
+ ad=0 pd=0 as=8.87095e+08 ps=187960 
M3003 GND diff_1203960_786130# diff_1248410_791210# GND efet w=53975 l=8255
+ ad=0 pd=0 as=0 ps=0 
M3004 GND diff_1339850_786130# diff_1223010_990600# GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3005 diff_1400810_873760# diff_1391920_806450# GND GND efet w=26670 l=8255
+ ad=0 pd=0 as=0 ps=0 
M3006 diff_1391920_806450# diff_1391920_806450# diff_1391920_806450# GND efet w=1270 l=6350
+ ad=0 pd=0 as=0 ps=0 
M3007 diff_1391920_806450# diff_1391920_806450# diff_1391920_806450# GND efet w=3175 l=5080
+ ad=0 pd=0 as=0 ps=0 
M3008 Vdd Vdd diff_1470660_825500# GND efet w=8890 l=60960
+ ad=0 pd=0 as=6.24192e+08 ps=149860 
M3009 diff_1402080_830580# Vdd Vdd GND efet w=7620 l=48260
+ ad=8.29031e+08 pd=190500 as=0 ps=0 
M3010 diff_1402080_830580# diff_1402080_830580# diff_1402080_830580# GND efet w=1270 l=6350
+ ad=0 pd=0 as=0 ps=0 
M3011 diff_1402080_830580# diff_1402080_830580# diff_1402080_830580# GND efet w=2540 l=5080
+ ad=0 pd=0 as=0 ps=0 
M3012 GND diff_1402080_830580# diff_1470660_825500# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3013 GND diff_1402080_830580# diff_1391920_806450# GND efet w=15240 l=8890
+ ad=0 pd=0 as=0 ps=0 
M3014 diff_1400810_873760# diff_1400810_873760# diff_1400810_873760# GND efet w=2540 l=4445
+ ad=0 pd=0 as=0 ps=0 
M3015 diff_1400810_873760# diff_1400810_873760# diff_1400810_873760# GND efet w=2540 l=3175
+ ad=0 pd=0 as=0 ps=0 
M3016 diff_1576070_459740# diff_1576070_459740# diff_1576070_459740# GND efet w=1270 l=6350
+ ad=0 pd=0 as=0 ps=0 
M3017 diff_897890_1024890# diff_897890_1024890# diff_897890_1024890# GND efet w=1905 l=5715
+ ad=0 pd=0 as=0 ps=0 
M3018 diff_897890_1024890# diff_897890_1024890# diff_897890_1024890# GND efet w=3810 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3019 diff_1677670_457200# diff_1677670_457200# diff_1677670_457200# GND efet w=2540 l=5080
+ ad=0 pd=0 as=0 ps=0 
M3020 diff_897890_1024890# clk2 diff_2578100_981710# GND efet w=15240 l=7620
+ ad=0 pd=0 as=2.87096e+08 ps=68580 
M3021 diff_1677670_457200# diff_1677670_457200# diff_1677670_457200# GND efet w=1270 l=5080
+ ad=0 pd=0 as=0 ps=0 
M3022 Vdd Vdd diff_1513840_989330# GND efet w=10160 l=39370
+ ad=0 pd=0 as=0 ps=0 
M3023 Vdd Vdd diff_1630680_786130# GND efet w=8890 l=60960
+ ad=0 pd=0 as=6.61289e+08 ps=160020 
M3024 Vdd Vdd diff_1691640_873760# GND efet w=10160 l=39370
+ ad=0 pd=0 as=0 ps=0 
M3025 diff_1682750_806450# Vdd Vdd GND efet w=7620 l=48260
+ ad=8.25805e+08 pd=208280 as=0 ps=0 
M3026 GND diff_2578100_981710# diff_2315210_670560# GND efet w=27305 l=7620
+ ad=0 pd=0 as=-9.69167e+08 ps=868680 
M3027 diff_1513840_989330# diff_1513840_989330# diff_1513840_989330# GND efet w=1905 l=5715
+ ad=0 pd=0 as=0 ps=0 
M3028 GND diff_1391920_806450# diff_1402080_830580# GND efet w=15875 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3029 diff_1513840_989330# diff_1513840_989330# diff_1513840_989330# GND efet w=3810 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3030 diff_1630680_786130# diff_1630680_786130# diff_1630680_786130# GND efet w=1905 l=6985
+ ad=0 pd=0 as=0 ps=0 
M3031 diff_1630680_786130# diff_1630680_786130# diff_1630680_786130# GND efet w=3175 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3032 diff_1470660_825500# diff_1099820_863600# diff_1390650_749300# GND efet w=13970 l=8890
+ ad=0 pd=0 as=4.82257e+08 ps=101600 
M3033 diff_1400810_873760# diff_1099820_863600# diff_1494790_784860# GND efet w=15240 l=8890
+ ad=0 pd=0 as=4.99999e+08 ps=96520 
M3034 diff_1313180_713740# diff_1313180_713740# diff_1313180_713740# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M3035 diff_1391920_806450# diff_1111250_830580# diff_1379220_753110# GND efet w=33655 l=8255
+ ad=0 pd=0 as=8.82256e+08 ps=195580 
M3036 diff_1313180_713740# diff_1313180_713740# diff_1313180_713740# GND efet w=1905 l=1905
+ ad=0 pd=0 as=0 ps=0 
M3037 diff_1339850_786130# diff_1313180_713740# GND GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3038 GND diff_1390650_749300# diff_1379220_753110# GND efet w=62230 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3039 diff_1513840_989330# diff_1005840_731520# diff_1600200_718820# GND efet w=13970 l=8255
+ ad=0 pd=0 as=1.17742e+09 ps=261620 
M3040 diff_1402080_830580# diff_1111250_830580# diff_1539240_795020# GND efet w=29210 l=8890
+ ad=0 pd=0 as=8.59676e+08 ps=190500 
M3041 diff_1539240_795020# diff_1494790_784860# GND GND efet w=53340 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3042 GND diff_1630680_786130# diff_1513840_989330# GND efet w=25400 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3043 GND diff_1682750_806450# diff_1691640_873760# GND efet w=25400 l=8255
+ ad=0 pd=0 as=0 ps=0 
M3044 diff_1682750_806450# diff_1682750_806450# diff_1682750_806450# GND efet w=1270 l=6350
+ ad=0 pd=0 as=0 ps=0 
M3045 diff_1682750_806450# diff_1682750_806450# diff_1682750_806450# GND efet w=2540 l=4445
+ ad=0 pd=0 as=0 ps=0 
M3046 Vdd Vdd diff_1761490_825500# GND efet w=8890 l=60960
+ ad=0 pd=0 as=6.37095e+08 ps=152400 
M3047 diff_1692910_830580# Vdd Vdd GND efet w=7620 l=48260
+ ad=8.09676e+08 pd=185420 as=0 ps=0 
M3048 diff_1692910_830580# diff_1692910_830580# diff_1692910_830580# GND efet w=1905 l=6985
+ ad=0 pd=0 as=0 ps=0 
M3049 diff_1692910_830580# diff_1692910_830580# diff_1692910_830580# GND efet w=2540 l=4445
+ ad=0 pd=0 as=0 ps=0 
M3050 GND diff_1692910_830580# diff_1761490_825500# GND efet w=14605 l=9525
+ ad=0 pd=0 as=0 ps=0 
M3051 GND diff_1692910_830580# diff_1682750_806450# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3052 diff_1691640_873760# diff_1691640_873760# diff_1691640_873760# GND efet w=2540 l=4445
+ ad=0 pd=0 as=0 ps=0 
M3053 diff_1691640_873760# diff_1691640_873760# diff_1691640_873760# GND efet w=2540 l=5715
+ ad=0 pd=0 as=0 ps=0 
M3054 diff_1761490_825500# diff_1391920_806450# diff_1681480_749300# GND efet w=14605 l=8255
+ ad=0 pd=0 as=4.61289e+08 ps=93980 
M3055 Vdd Vdd diff_1888490_857250# GND efet w=10160 l=40640
+ ad=0 pd=0 as=0 ps=0 
M3056 Vdd Vdd diff_1922780_786130# GND efet w=8890 l=60960
+ ad=0 pd=0 as=6.4516e+08 ps=152400 
M3057 Vdd Vdd diff_1982470_873760# GND efet w=11430 l=39370
+ ad=0 pd=0 as=0 ps=0 
M3058 diff_1974850_806450# Vdd Vdd GND efet w=6985 l=48895
+ ad=8.19353e+08 pd=213360 as=0 ps=0 
M3059 diff_1888490_857250# diff_1888490_857250# diff_1888490_857250# GND efet w=1905 l=5715
+ ad=0 pd=0 as=0 ps=0 
M3060 diff_1888490_857250# diff_1888490_857250# diff_1888490_857250# GND efet w=3175 l=4445
+ ad=0 pd=0 as=0 ps=0 
M3061 GND diff_1682750_806450# diff_1692910_830580# GND efet w=14605 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3062 diff_1922780_786130# diff_1922780_786130# diff_1922780_786130# GND efet w=1270 l=6350
+ ad=0 pd=0 as=0 ps=0 
M3063 diff_1922780_786130# diff_1922780_786130# diff_1922780_786130# GND efet w=2540 l=5080
+ ad=0 pd=0 as=0 ps=0 
M3064 GND diff_1922780_786130# diff_1888490_857250# GND efet w=29845 l=8255
+ ad=0 pd=0 as=0 ps=0 
M3065 diff_1691640_873760# diff_1391920_806450# diff_1786890_783590# GND efet w=13970 l=7620
+ ad=0 pd=0 as=4.61289e+08 ps=93980 
M3066 diff_1682750_806450# diff_1402080_830580# diff_1670050_753110# GND efet w=31115 l=8255
+ ad=0 pd=0 as=8.79031e+08 ps=187960 
M3067 diff_1600200_718820# diff_1600200_718820# diff_1600200_718820# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M3068 diff_1600200_718820# diff_1600200_718820# diff_1600200_718820# GND efet w=1905 l=1905
+ ad=0 pd=0 as=0 ps=0 
M3069 diff_1022350_718820# diff_1018540_712470# diff_369570_1160780# GND efet w=13970 l=6350
+ ad=0 pd=0 as=0 ps=0 
M3070 diff_1313180_713740# diff_1018540_712470# diff_266700_2927350# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3071 Vdd Vdd diff_377190_637540# GND efet w=8890 l=62230
+ ad=0 pd=0 as=0 ps=0 
M3072 GND GND diff_586740_566420# GND efet w=40640 l=8255
+ ad=0 pd=0 as=1.87419e+09 ps=424180 
M3073 diff_377190_637540# clk1 diff_374650_585470# GND efet w=9525 l=6985
+ ad=0 pd=0 as=2.75806e+08 ps=96520 
M3074 GND diff_245110_1436370# diff_586740_566420# GND efet w=90170 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3075 diff_374650_585470# diff_374650_585470# diff_374650_585470# GND efet w=4445 l=4445
+ ad=0 pd=0 as=0 ps=0 
M3076 GND diff_374650_585470# diff_377190_574040# GND efet w=15240 l=6985
+ ad=0 pd=0 as=7.46773e+08 ps=167640 
M3077 diff_374650_585470# diff_374650_585470# diff_374650_585470# GND efet w=3175 l=5080
+ ad=0 pd=0 as=0 ps=0 
M3078 diff_586740_528320# Vdd diff_586740_566420# GND efet w=43815 l=8255
+ ad=-1.80788e+09 pd=530860 as=0 ps=0 
M3079 Vdd Vdd diff_377190_574040# GND efet w=8890 l=60960
+ ad=0 pd=0 as=0 ps=0 
M3080 GND diff_243840_2250440# diff_669290_508000# GND efet w=93980 l=8890
+ ad=0 pd=0 as=-1.54175e+09 ps=525780 
M3081 diff_640080_426720# diff_243840_2250440# GND GND efet w=49530 l=8890
+ ad=1.04193e+09 pd=246380 as=0 ps=0 
M3082 diff_586740_566420# diff_582930_558800# diff_586740_528320# GND efet w=57150 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3083 clk1 GND GND GND efet w=111760 l=6350
+ ad=-9.17499e+07 pd=675640 as=0 ps=0 
M3084 GND diff_302260_482600# diff_284480_472440# GND efet w=53340 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3085 diff_377190_574040# clk2 diff_373380_521970# GND efet w=8890 l=6350
+ ad=0 pd=0 as=2.8387e+08 ps=96520 
M3086 diff_373380_521970# diff_373380_521970# diff_373380_521970# GND efet w=3810 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3087 GND diff_373380_521970# diff_377190_510540# GND efet w=15240 l=6985
+ ad=0 pd=0 as=6.75805e+08 ps=154940 
M3088 GND diff_245110_1436370# diff_582930_558800# GND efet w=43180 l=8890
+ ad=0 pd=0 as=5.5645e+08 ps=127000 
M3089 diff_599440_977900# diff_599440_977900# diff_599440_977900# GND efet w=4445 l=4445
+ ad=-1.0982e+09 pd=894080 as=0 ps=0 
M3090 diff_599440_977900# diff_599440_977900# diff_599440_977900# GND efet w=3175 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3091 diff_787400_546100# diff_775970_467360# GND GND efet w=15240 l=7620
+ ad=6.77418e+08 pd=152400 as=0 ps=0 
M3092 diff_373380_521970# diff_373380_521970# diff_373380_521970# GND efet w=3175 l=5080
+ ad=0 pd=0 as=0 ps=0 
M3093 GND diff_325120_504190# diff_328930_492760# GND efet w=36830 l=6350
+ ad=0 pd=0 as=8.64514e+08 ps=180340 
M3094 Vdd Vdd diff_377190_510540# GND efet w=8890 l=60960
+ ad=0 pd=0 as=0 ps=0 
M3095 diff_582930_558800# Vdd Vdd GND efet w=11430 l=40640
+ ad=0 pd=0 as=0 ps=0 
M3096 GND p0 diff_669290_508000# GND efet w=43815 l=8255
+ ad=0 pd=0 as=0 ps=0 
M3097 GND p0 diff_694690_422910# GND efet w=15240 l=7620
+ ad=0 pd=0 as=6.08063e+08 ps=157480 
M3098 diff_772160_488950# diff_599440_977900# diff_787400_546100# GND efet w=14605 l=8255
+ ad=6.40321e+08 pd=157480 as=0 ps=0 
M3099 GND diff_599440_977900# diff_821690_471170# GND efet w=14605 l=9525
+ ad=0 pd=0 as=5.82257e+08 ps=139700 
M3100 diff_377190_510540# clk1 diff_325120_504190# GND efet w=15875 l=6985
+ ad=0 pd=0 as=2.5e+08 ps=63500 
M3101 diff_302260_482600# diff_302260_482600# diff_302260_482600# GND efet w=2540 l=7620
+ ad=2.70967e+08 pd=81280 as=0 ps=0 
M3102 diff_284480_472440# Vdd Vdd GND efet w=10160 l=19050
+ ad=0 pd=0 as=0 ps=0 
M3103 diff_302260_482600# diff_302260_482600# diff_302260_482600# GND efet w=3810 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3104 diff_328930_492760# clk2 diff_302260_482600# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3105 diff_669290_508000# diff_640080_426720# diff_586740_528320# GND efet w=58420 l=8890
+ ad=0 pd=0 as=0 ps=0 
M3106 diff_328930_492760# Vdd Vdd GND efet w=10795 l=28575
+ ad=0 pd=0 as=0 ps=0 
M3107 diff_694690_422910# diff_694690_422910# diff_694690_422910# GND efet w=3810 l=5080
+ ad=0 pd=0 as=0 ps=0 
M3108 diff_775970_467360# diff_772160_488950# GND GND efet w=26035 l=8255
+ ad=3.88709e+08 pd=88900 as=0 ps=0 
M3109 diff_694690_422910# diff_694690_422910# diff_694690_422910# GND efet w=3175 l=6350
+ ad=0 pd=0 as=0 ps=0 
M3110 diff_821690_471170# diff_821690_471170# diff_821690_471170# GND efet w=3175 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3111 diff_857250_500380# diff_821690_471170# diff_586740_528320# GND efet w=13970 l=8890
+ ad=4.98386e+08 pd=127000 as=0 ps=0 
M3112 diff_586740_528320# diff_694690_422910# diff_669290_508000# GND efet w=57150 l=8890
+ ad=0 pd=0 as=0 ps=0 
M3113 Vdd Vdd diff_358140_298450# GND efet w=9525 l=6985
+ ad=0 pd=0 as=2.87096e+08 ps=88900 
M3114 diff_214630_541020# diff_358140_298450# diff_214630_541020# GND efet w=55245 l=11430
+ ad=1.70161e+09 pd=388620 as=0 ps=0 
M3115 diff_358140_298450# diff_358140_298450# diff_358140_298450# GND efet w=3175 l=5715
+ ad=0 pd=0 as=0 ps=0 
M3116 diff_358140_298450# diff_358140_298450# diff_358140_298450# GND efet w=1270 l=5080
+ ad=0 pd=0 as=0 ps=0 
M3117 diff_214630_541020# diff_358140_298450# Vdd GND efet w=12700 l=21590
+ ad=0 pd=0 as=0 ps=0 
M3118 Vdd Vdd diff_387350_243840# GND efet w=8890 l=60960
+ ad=0 pd=0 as=4.41935e+08 ps=99060 
M3119 Vdd diff_505460_347980# diff_139700_2962910# GND efet w=21590 l=6985
+ ad=0 pd=0 as=-1.19169e+08 ps=1.00076e+06 
M3120 diff_139700_2962910# diff_487680_288290# GND GND efet w=20320 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3121 diff_387350_243840# clk1 diff_438150_274320# GND efet w=29210 l=8890
+ ad=0 pd=0 as=4.8387e+08 ps=101600 
M3122 diff_214630_541020# diff_387350_243840# GND GND efet w=46990 l=6985
+ ad=0 pd=0 as=0 ps=0 
M3123 diff_438150_274320# diff_434340_266700# GND GND efet w=27940 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3124 Vdd Vdd diff_487680_288290# GND efet w=8890 l=60960
+ ad=0 pd=0 as=4.41935e+08 ps=96520 
M3125 diff_640080_426720# Vdd Vdd GND efet w=10160 l=33020
+ ad=0 pd=0 as=0 ps=0 
M3126 Vdd Vdd diff_586740_528320# GND efet w=11430 l=41910
+ ad=0 pd=0 as=0 ps=0 
M3127 diff_694690_422910# Vdd Vdd GND efet w=8890 l=61595
+ ad=0 pd=0 as=0 ps=0 
M3128 diff_821690_471170# diff_821690_471170# diff_821690_471170# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M3129 diff_1630680_786130# diff_1600200_718820# GND GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3130 GND diff_1681480_749300# diff_1670050_753110# GND efet w=60325 l=8255
+ ad=0 pd=0 as=0 ps=0 
M3131 diff_1888490_857250# diff_1005840_731520# diff_1894840_732790# GND efet w=15240 l=8255
+ ad=0 pd=0 as=1.15806e+09 ps=246380 
M3132 diff_1692910_830580# diff_1402080_830580# diff_1831340_789940# GND efet w=27940 l=7620
+ ad=0 pd=0 as=8.08063e+08 ps=185420 
M3133 diff_1831340_789940# diff_1786890_783590# GND GND efet w=53340 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3134 diff_1982470_873760# diff_1974850_806450# GND GND efet w=26670 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3135 diff_1974850_806450# diff_1974850_806450# diff_1974850_806450# GND efet w=1905 l=6985
+ ad=0 pd=0 as=0 ps=0 
M3136 diff_1974850_806450# diff_1974850_806450# diff_1974850_806450# GND efet w=3175 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3137 Vdd Vdd diff_2053590_824230# GND efet w=8890 l=60960
+ ad=0 pd=0 as=6.22579e+08 ps=149860 
M3138 diff_1983740_830580# Vdd Vdd GND efet w=7620 l=53975
+ ad=8.59676e+08 pd=200660 as=0 ps=0 
M3139 diff_1983740_830580# diff_1983740_830580# diff_1983740_830580# GND efet w=1270 l=6350
+ ad=0 pd=0 as=0 ps=0 
M3140 diff_1983740_830580# diff_1983740_830580# diff_1983740_830580# GND efet w=3175 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3141 GND diff_1983740_830580# diff_2053590_824230# GND efet w=13970 l=8890
+ ad=0 pd=0 as=0 ps=0 
M3142 GND diff_1983740_830580# diff_1974850_806450# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3143 diff_1982470_873760# diff_1982470_873760# diff_1982470_873760# GND efet w=1905 l=3175
+ ad=0 pd=0 as=0 ps=0 
M3144 diff_1982470_873760# diff_1982470_873760# diff_1982470_873760# GND efet w=3175 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3145 GND diff_1974850_806450# diff_1983740_830580# GND efet w=15240 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3146 diff_2053590_824230# diff_1682750_806450# diff_1973580_749300# GND efet w=14605 l=8255
+ ad=0 pd=0 as=4.66128e+08 ps=96520 
M3147 diff_1982470_873760# diff_1682750_806450# diff_2077720_787400# GND efet w=15240 l=7620
+ ad=0 pd=0 as=4.96773e+08 ps=96520 
M3148 diff_1974850_806450# diff_1692910_830580# diff_1960880_777240# GND efet w=27940 l=7620
+ ad=0 pd=0 as=9.01611e+08 ps=190500 
M3149 diff_1894840_732790# diff_1894840_732790# diff_1894840_732790# GND efet w=3810 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3150 diff_1894840_732790# diff_1894840_732790# diff_1894840_732790# GND efet w=2540 l=2540
+ ad=0 pd=0 as=0 ps=0 
M3151 diff_1922780_786130# diff_1894840_732790# GND GND efet w=24130 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3152 GND diff_1973580_749300# diff_1960880_777240# GND efet w=60960 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3153 diff_1983740_830580# diff_1692910_830580# diff_2123440_789940# GND efet w=27940 l=7620
+ ad=0 pd=0 as=8.12902e+08 ps=190500 
M3154 GND diff_2077720_787400# diff_2123440_789940# GND efet w=55880 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3155 diff_1894840_732790# diff_1018540_712470# diff_245110_1436370# GND efet w=18415 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3156 GND diff_1997710_740410# diff_2002790_702310# GND efet w=68580 l=7620
+ ad=0 pd=0 as=-1.57562e+09 ps=614680 
M3157 diff_1600200_718820# diff_1018540_712470# diff_243840_2250440# GND efet w=13970 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3158 diff_2002790_702310# diff_1997710_690880# diff_2002790_702310# GND efet w=45720 l=22860
+ ad=0 pd=0 as=0 ps=0 
M3159 diff_1736090_635000# Vdd Vdd GND efet w=12065 l=36830
+ ad=7.80644e+08 pd=157480 as=0 ps=0 
M3160 diff_2002790_702310# diff_1997710_690880# Vdd GND efet w=10795 l=12065
+ ad=0 pd=0 as=0 ps=0 
M3161 GND diff_775970_467360# diff_900430_483870# GND efet w=36830 l=7620
+ ad=0 pd=0 as=1.06613e+09 ps=220980 
M3162 diff_1149350_486410# diff_857250_500380# GND GND efet w=25400 l=7620
+ ad=9.2903e+08 pd=228600 as=0 ps=0 
M3163 Vdd Vdd diff_1790700_659130# GND efet w=11430 l=20320
+ ad=0 pd=0 as=0 ps=0 
M3164 diff_1997710_690880# diff_1997710_690880# diff_1997710_690880# GND efet w=1270 l=5080
+ ad=2.46774e+08 pd=78740 as=0 ps=0 
M3165 diff_1997710_690880# diff_1997710_690880# diff_1997710_690880# GND efet w=3175 l=4445
+ ad=0 pd=0 as=0 ps=0 
M3166 diff_1838960_473710# Vdd Vdd GND efet w=11430 l=40640
+ ad=1.25806e+09 pd=309880 as=0 ps=0 
M3167 Vdd Vdd diff_1894840_476250# GND efet w=10795 l=40005
+ ad=0 pd=0 as=1.61613e+09 ps=383540 
M3168 diff_1681480_645160# diff_900430_483870# diff_243840_2250440# GND efet w=13970 l=7620
+ ad=2.32258e+08 pd=63500 as=0 ps=0 
M3169 diff_1736090_635000# diff_1736090_635000# diff_1736090_635000# GND efet w=1905 l=3175
+ ad=0 pd=0 as=0 ps=0 
M3170 diff_1790700_659130# diff_1736090_635000# GND GND efet w=61595 l=8255
+ ad=0 pd=0 as=0 ps=0 
M3171 diff_1790700_659130# diff_1790700_659130# diff_1790700_659130# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M3172 diff_1838960_473710# diff_1790700_659130# GND GND efet w=34290 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3173 diff_1790700_659130# diff_1790700_659130# diff_1790700_659130# GND efet w=2540 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3174 diff_1736090_635000# diff_1736090_635000# diff_1736090_635000# GND efet w=1905 l=1905
+ ad=0 pd=0 as=0 ps=0 
M3175 diff_266700_2927350# diff_900430_483870# diff_1507490_548640# GND efet w=13970 l=7620
+ ad=0 pd=0 as=2.8387e+08 ps=68580 
M3176 diff_369570_1160780# diff_900430_483870# diff_1569720_548640# GND efet w=13970 l=7620
+ ad=0 pd=0 as=2.8387e+08 ps=68580 
M3177 GND diff_408940_681990# diff_857250_500380# GND efet w=15875 l=8255
+ ad=0 pd=0 as=0 ps=0 
M3178 diff_1149350_486410# diff_1149350_486410# diff_1149350_486410# GND efet w=6985 l=4445
+ ad=0 pd=0 as=0 ps=0 
M3179 diff_1149350_486410# diff_1037590_429260# GND GND efet w=15240 l=8890
+ ad=0 pd=0 as=0 ps=0 
M3180 GND clk2 diff_1239520_518160# GND efet w=24130 l=8890
+ ad=0 pd=0 as=3.43548e+08 ps=86360 
M3181 diff_1149350_486410# diff_1149350_486410# diff_1149350_486410# GND efet w=4445 l=9525
+ ad=0 pd=0 as=0 ps=0 
M3182 GND diff_1149350_486410# diff_1183640_483870# GND efet w=14605 l=8255
+ ad=0 pd=0 as=2.90322e+08 ps=73660 
M3183 diff_1239520_518160# diff_699770_264160# diff_1239520_500380# GND efet w=32385 l=8255
+ ad=0 pd=0 as=2.8387e+08 ps=83820 
M3184 diff_1239520_500380# diff_1183640_483870# diff_1239520_481330# GND efet w=31750 l=8890
+ ad=0 pd=0 as=7.99998e+08 ps=165100 
M3185 diff_775970_467360# Vdd Vdd GND efet w=8890 l=60960
+ ad=0 pd=0 as=0 ps=0 
M3186 diff_787400_546100# Vdd Vdd GND efet w=8890 l=60325
+ ad=0 pd=0 as=0 ps=0 
M3187 diff_821690_471170# Vdd Vdd GND efet w=8890 l=60960
+ ad=0 pd=0 as=0 ps=0 
M3188 diff_586740_528320# diff_821690_471170# diff_772160_488950# GND efet w=15240 l=8890
+ ad=0 pd=0 as=0 ps=0 
M3189 GND diff_924560_458470# diff_900430_483870# GND efet w=35560 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3190 diff_1007110_440690# clk2 diff_599440_977900# GND efet w=33020 l=8890
+ ad=4.69354e+08 pd=106680 as=0 ps=0 
M3191 diff_900430_483870# Vdd Vdd GND efet w=10160 l=30480
+ ad=0 pd=0 as=0 ps=0 
M3192 diff_599440_977900# Vdd Vdd GND efet w=8890 l=60960
+ ad=0 pd=0 as=0 ps=0 
M3193 diff_487680_288290# diff_505460_347980# GND GND efet w=15240 l=8890
+ ad=0 pd=0 as=0 ps=0 
M3194 Vdd Vdd diff_505460_347980# GND efet w=8890 l=60960
+ ad=0 pd=0 as=1.08387e+09 ps=203200 
M3195 diff_581660_321310# Vdd Vdd GND efet w=7620 l=58420
+ ad=3.30645e+08 pd=86360 as=0 ps=0 
M3196 Vdd Vdd diff_622300_264160# GND efet w=7620 l=48260
+ ad=0 pd=0 as=9.95159e+08 ps=185420 
M3197 diff_664210_320040# diff_434340_266700# Vdd GND efet w=14605 l=8255
+ ad=3.1129e+08 pd=78740 as=0 ps=0 
M3198 diff_664210_320040# clk1 diff_647700_243840# GND efet w=8890 l=7620
+ ad=0 pd=0 as=7.0645e+08 ps=152400 
M3199 GND diff_737870_302260# diff_581660_321310# GND efet w=13335 l=9525
+ ad=0 pd=0 as=0 ps=0 
M3200 diff_647700_243840# diff_647700_243840# diff_647700_243840# GND efet w=4445 l=4445
+ ad=0 pd=0 as=0 ps=0 
M3201 diff_647700_243840# diff_647700_243840# diff_647700_243840# GND efet w=2540 l=6350
+ ad=0 pd=0 as=0 ps=0 
M3202 diff_622300_264160# diff_622300_264160# diff_622300_264160# GND efet w=4445 l=4445
+ ad=0 pd=0 as=0 ps=0 
M3203 GND diff_647700_243840# diff_622300_264160# GND efet w=45085 l=8255
+ ad=0 pd=0 as=0 ps=0 
M3204 diff_622300_264160# diff_622300_264160# diff_622300_264160# GND efet w=1905 l=10160
+ ad=0 pd=0 as=0 ps=0 
M3205 GND diff_699770_264160# diff_647700_243840# GND efet w=17145 l=8255
+ ad=0 pd=0 as=0 ps=0 
M3206 diff_1027430_431800# diff_1018540_320040# diff_1007110_440690# GND efet w=42545 l=9525
+ ad=4.38709e+08 pd=106680 as=0 ps=0 
M3207 GND diff_1037590_429260# diff_1027430_431800# GND efet w=43180 l=8890
+ ad=0 pd=0 as=0 ps=0 
M3208 diff_1149350_486410# Vdd Vdd GND efet w=8890 l=63500
+ ad=0 pd=0 as=0 ps=0 
M3209 Vdd Vdd diff_434340_266700# GND efet w=10160 l=40005
+ ad=0 pd=0 as=6.79031e+08 ps=137160 
M3210 diff_1101090_427990# diff_1037590_429260# diff_924560_458470# GND efet w=33020 l=8890
+ ad=3.35483e+08 pd=86360 as=5.70967e+08 ps=119380 
M3211 diff_1118870_429260# diff_1111250_266700# diff_1101090_427990# GND efet w=32385 l=8255
+ ad=3.09677e+08 pd=86360 as=0 ps=0 
M3212 GND clk2 diff_1118870_429260# GND efet w=24765 l=9525
+ ad=0 pd=0 as=0 ps=0 
M3213 diff_924560_458470# Vdd Vdd GND efet w=8890 l=78740
+ ad=0 pd=0 as=0 ps=0 
M3214 GND diff_829310_237490# diff_434340_266700# GND efet w=23495 l=10795
+ ad=0 pd=0 as=0 ps=0 
M3215 diff_505460_347980# diff_581660_321310# GND GND efet w=16510 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3216 GND diff_622300_264160# diff_505460_347980# GND efet w=16510 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3217 clk2 GND GND GND efet w=111760 l=8890
+ ad=1.66631e+09 pd=967740 as=0 ps=0 
M3218 diff_1183640_483870# Vdd Vdd GND efet w=8890 l=62230
+ ad=0 pd=0 as=0 ps=0 
M3219 Vdd Vdd diff_1239520_481330# GND efet w=8890 l=77470
+ ad=0 pd=0 as=0 ps=0 
M3220 diff_1018540_712470# diff_1239520_481330# GND GND efet w=36830 l=8890
+ ad=6.74192e+08 pd=165100 as=0 ps=0 
M3221 diff_1005840_731520# diff_1005840_731520# diff_1005840_731520# GND efet w=1905 l=5715
+ ad=1.00161e+09 pd=259080 as=0 ps=0 
M3222 diff_1005840_731520# diff_1005840_731520# diff_1005840_731520# GND efet w=3810 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3223 diff_1005840_731520# diff_1018540_712470# GND GND efet w=45720 l=8890
+ ad=0 pd=0 as=0 ps=0 
M3224 diff_1736090_635000# diff_1681480_645160# GND GND efet w=43180 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3225 Vdd Vdd Vdd GND efet w=2540 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3226 Vdd Vdd Vdd GND efet w=1905 l=1905
+ ad=0 pd=0 as=0 ps=0 
M3227 Vdd diff_2247900_798830# diff_894080_1518920# GND efet w=23495 l=6985
+ ad=0 pd=0 as=0 ps=0 
M3228 Vdd Vdd Vdd GND efet w=1270 l=3175
+ ad=0 pd=0 as=0 ps=0 
M3229 diff_2315210_670560# Vdd Vdd GND efet w=11430 l=39370
+ ad=0 pd=0 as=0 ps=0 
M3230 Vdd Vdd Vdd GND efet w=3175 l=5080
+ ad=0 pd=0 as=0 ps=0 
M3231 Vdd Vdd diff_2297430_869950# GND efet w=11430 l=29210
+ ad=0 pd=0 as=8.64514e+08 ps=190500 
M3232 diff_2315210_670560# clk1 diff_2559050_902970# GND efet w=15240 l=7620
+ ad=0 pd=0 as=2.77419e+08 ps=71120 
M3233 GND diff_2559050_902970# diff_1111250_266700# GND efet w=53975 l=6985
+ ad=0 pd=0 as=-1.83691e+09 ps=629920 
M3234 Vdd Vdd diff_2246630_834390# GND efet w=8890 l=7620
+ ad=0 pd=0 as=2.41935e+08 ps=81280 
M3235 diff_894080_1518920# diff_2297430_869950# GND GND efet w=21590 l=6350
+ ad=0 pd=0 as=0 ps=0 
M3236 diff_2297430_869950# diff_2297430_869950# diff_2297430_869950# GND efet w=2540 l=6350
+ ad=0 pd=0 as=0 ps=0 
M3237 diff_2246630_834390# diff_2246630_834390# diff_2246630_834390# GND efet w=2540 l=6350
+ ad=0 pd=0 as=0 ps=0 
M3238 diff_2246630_834390# diff_2246630_834390# diff_2246630_834390# GND efet w=3175 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3239 diff_2324100_800100# clk2 diff_2297430_869950# GND efet w=55245 l=6985
+ ad=1.45645e+09 pd=269240 as=0 ps=0 
M3240 diff_2297430_869950# diff_2297430_869950# diff_2297430_869950# GND efet w=1905 l=4445
+ ad=0 pd=0 as=0 ps=0 
M3241 GND diff_2297430_869950# diff_2247900_798830# GND efet w=24130 l=7620
+ ad=0 pd=0 as=1.35645e+09 ps=355600 
M3242 Vdd diff_2246630_834390# diff_2247900_798830# GND efet w=10160 l=27940
+ ad=0 pd=0 as=0 ps=0 
M3243 Vdd Vdd Vdd GND efet w=2540 l=4445
+ ad=0 pd=0 as=0 ps=0 
M3244 Vdd Vdd Vdd GND efet w=3810 l=8255
+ ad=0 pd=0 as=0 ps=0 
M3245 diff_1111250_266700# Vdd Vdd GND efet w=11430 l=20320
+ ad=0 pd=0 as=0 ps=0 
M3246 GND diff_1111250_266700# diff_2324100_800100# GND efet w=76200 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3247 diff_1111250_266700# diff_1111250_266700# diff_1111250_266700# GND efet w=1905 l=6350
+ ad=0 pd=0 as=0 ps=0 
M3248 diff_1111250_266700# diff_1111250_266700# diff_1111250_266700# GND efet w=3810 l=5080
+ ad=0 pd=0 as=0 ps=0 
M3249 diff_1111250_266700# clk2 diff_2555240_824230# GND efet w=15240 l=6985
+ ad=0 pd=0 as=2.85483e+08 ps=68580 
M3250 diff_2247900_798830# diff_2246630_834390# diff_2247900_798830# GND efet w=56515 l=19685
+ ad=0 pd=0 as=0 ps=0 
M3251 GND diff_2555240_824230# diff_829310_237490# GND efet w=55245 l=6985
+ ad=0 pd=0 as=1.19838e+09 ps=243840 
M3252 Vdd Vdd Vdd GND efet w=1905 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3253 diff_2324100_800100# diff_755650_927100# GND GND efet w=49530 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3254 GND diff_2228850_712470# diff_2245360_692150# GND efet w=107950 l=7620
+ ad=0 pd=0 as=1.67419e+09 ps=342900 
M3255 Vdd Vdd Vdd GND efet w=3175 l=8890
+ ad=0 pd=0 as=0 ps=0 
M3256 diff_829310_237490# Vdd Vdd GND efet w=11430 l=20320
+ ad=0 pd=0 as=0 ps=0 
M3257 diff_829310_237490# clk1 diff_2536190_745490# GND efet w=15240 l=7620
+ ad=0 pd=0 as=2.79032e+08 ps=71120 
M3258 diff_2320290_678180# diff_2153920_452120# GND GND efet w=85090 l=7620
+ ad=2.14677e+09 pd=396240 as=0 ps=0 
M3259 Vdd Vdd Vdd GND efet w=1905 l=3175
+ ad=0 pd=0 as=0 ps=0 
M3260 GND diff_2536190_745490# diff_932180_1050290# GND efet w=53340 l=7620
+ ad=0 pd=0 as=1.15e+09 ps=233680 
M3261 Vdd Vdd Vdd GND efet w=3175 l=5715
+ ad=0 pd=0 as=0 ps=0 
M3262 diff_932180_1050290# Vdd Vdd GND efet w=11430 l=20320
+ ad=0 pd=0 as=0 ps=0 
M3263 diff_2320290_678180# diff_2014220_425450# GND GND efet w=83820 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3264 diff_1997710_740410# clk1 diff_2245360_692150# GND efet w=81280 l=7620
+ ad=9.95159e+08 pd=193040 as=0 ps=0 
M3265 diff_1997710_690880# Vdd Vdd GND efet w=8890 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3266 diff_1894840_476250# diff_1790700_659130# GND GND efet w=32385 l=8255
+ ad=0 pd=0 as=0 ps=0 
M3267 Vdd Vdd Vdd GND efet w=4445 l=10795
+ ad=0 pd=0 as=0 ps=0 
M3268 Vdd Vdd Vdd GND efet w=6985 l=4445
+ ad=0 pd=0 as=0 ps=0 
M3269 GND diff_1576070_459740# diff_1894840_476250# GND efet w=32385 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3270 diff_1838960_473710# diff_1518920_467360# GND GND efet w=33655 l=8255
+ ad=0 pd=0 as=0 ps=0 
M3271 diff_2124710_610870# Vdd Vdd GND efet w=8255 l=8255
+ ad=2.74193e+08 pd=78740 as=0 ps=0 
M3272 diff_2124710_610870# diff_2124710_610870# diff_2124710_610870# GND efet w=1270 l=5080
+ ad=0 pd=0 as=0 ps=0 
M3273 diff_2124710_610870# diff_2124710_610870# diff_2124710_610870# GND efet w=1905 l=5715
+ ad=0 pd=0 as=0 ps=0 
M3274 diff_232410_996950# diff_2124710_610870# diff_232410_996950# GND efet w=72390 l=24130
+ ad=3.43733e+08 pd=1.14808e+06 as=0 ps=0 
M3275 diff_1997710_740410# Vdd Vdd GND efet w=10160 l=20320
+ ad=0 pd=0 as=0 ps=0 
M3276 diff_2320290_678180# diff_2315210_670560# diff_2228850_712470# GND efet w=70485 l=8255
+ ad=0 pd=0 as=8.1774e+08 ps=162560 
M3277 diff_755650_927100# diff_2203450_571500# diff_755650_927100# GND efet w=70485 l=34925
+ ad=-3.38524e+08 pd=985520 as=0 ps=0 
M3278 diff_232410_996950# diff_2124710_610870# Vdd GND efet w=10160 l=11430
+ ad=0 pd=0 as=0 ps=0 
M3279 GND diff_1677670_457200# diff_1838960_473710# GND efet w=25400 l=10160
+ ad=0 pd=0 as=0 ps=0 
M3280 GND diff_408940_681990# diff_1416050_494030# GND efet w=14605 l=8255
+ ad=0 pd=0 as=3.01612e+08 ps=71120 
M3281 diff_1018540_712470# diff_1018540_712470# diff_1018540_712470# GND efet w=2540 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3282 diff_1018540_712470# diff_1018540_712470# diff_1018540_712470# GND efet w=1905 l=5715
+ ad=0 pd=0 as=0 ps=0 
M3283 GND diff_1343660_488950# diff_1005840_731520# GND efet w=38100 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3284 diff_1701800_544830# diff_900430_483870# diff_245110_1436370# GND efet w=13970 l=7620
+ ad=2.29032e+08 pd=78740 as=0 ps=0 
M3285 diff_1701800_544830# diff_1701800_544830# diff_1701800_544830# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M3286 diff_1701800_544830# diff_1701800_544830# diff_1701800_544830# GND efet w=3175 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3287 diff_1416050_494030# diff_900430_483870# Vdd GND efet w=15240 l=8255
+ ad=0 pd=0 as=0 ps=0 
M3288 diff_1018540_712470# Vdd Vdd GND efet w=10795 l=31115
+ ad=0 pd=0 as=0 ps=0 
M3289 diff_1465580_462280# diff_1416050_494030# GND GND efet w=66675 l=8255
+ ad=7.69353e+08 pd=170180 as=0 ps=0 
M3290 diff_1005840_731520# Vdd Vdd GND efet w=11430 l=33020
+ ad=0 pd=0 as=0 ps=0 
M3291 diff_1343660_488950# diff_829310_237490# GND GND efet w=40005 l=10795
+ ad=3.88709e+08 pd=91440 as=0 ps=0 
M3292 diff_1518920_467360# diff_1507490_548640# GND GND efet w=52070 l=7620
+ ad=8.5645e+08 pd=180340 as=0 ps=0 
M3293 diff_1518920_467360# diff_1518920_467360# diff_1518920_467360# GND efet w=3810 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3294 diff_1518920_467360# diff_1518920_467360# diff_1518920_467360# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M3295 diff_1576070_459740# diff_1518920_467360# GND GND efet w=34290 l=8890
+ ad=0 pd=0 as=0 ps=0 
M3296 GND diff_1604010_461010# diff_1894840_476250# GND efet w=32385 l=8255
+ ad=0 pd=0 as=0 ps=0 
M3297 diff_1894840_476250# diff_1701800_544830# GND GND efet w=53975 l=8255
+ ad=0 pd=0 as=0 ps=0 
M3298 GND diff_1465580_462280# diff_1894840_476250# GND efet w=26035 l=8255
+ ad=0 pd=0 as=0 ps=0 
M3299 Vdd Vdd diff_2203450_571500# GND efet w=8255 l=8255
+ ad=0 pd=0 as=2.67741e+08 ps=83820 
M3300 diff_2228850_712470# Vdd Vdd GND efet w=10795 l=29845
+ ad=0 pd=0 as=0 ps=0 
M3301 diff_932180_1050290# clk2 diff_2541270_668020# GND efet w=15240 l=6350
+ ad=0 pd=0 as=2.8387e+08 ps=68580 
M3302 GND diff_2541270_668020# diff_2153920_452120# GND efet w=43815 l=6985
+ ad=0 pd=0 as=3.3083e+08 ps=1.22174e+06 
M3303 Vdd Vdd Vdd GND efet w=1905 l=2540
+ ad=0 pd=0 as=0 ps=0 
M3304 Vdd Vdd Vdd GND efet w=2540 l=3175
+ ad=0 pd=0 as=0 ps=0 
M3305 diff_2153920_452120# Vdd Vdd GND efet w=12065 l=29845
+ ad=0 pd=0 as=0 ps=0 
M3306 diff_2203450_571500# diff_2203450_571500# diff_2203450_571500# GND efet w=1270 l=6350
+ ad=0 pd=0 as=0 ps=0 
M3307 diff_2203450_571500# diff_2203450_571500# diff_2203450_571500# GND efet w=2540 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3308 Vdd Vdd Vdd GND efet w=5715 l=10795
+ ad=0 pd=0 as=0 ps=0 
M3309 Vdd Vdd Vdd GND efet w=3175 l=10795
+ ad=0 pd=0 as=0 ps=0 
M3310 diff_2153920_452120# clk1 diff_2517140_586740# GND efet w=14605 l=6350
+ ad=0 pd=0 as=2.53225e+08 ps=66040 
M3311 Vdd Vdd diff_2195830_2933700# GND efet w=10795 l=20320
+ ad=0 pd=0 as=-4.17556e+08 ps=883920 
M3312 Vdd diff_2203450_571500# diff_755650_927100# GND efet w=10160 l=20320
+ ad=0 pd=0 as=0 ps=0 
M3313 diff_232410_996950# diff_2089150_548640# GND GND efet w=80010 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3314 diff_755650_927100# diff_2089150_548640# GND GND efet w=48895 l=6985
+ ad=0 pd=0 as=0 ps=0 
M3315 Vdd Vdd diff_2192020_525780# GND efet w=10160 l=29210
+ ad=0 pd=0 as=6.77418e+08 ps=154940 
M3316 GND diff_2517140_586740# diff_1018540_320040# GND efet w=56515 l=6985
+ ad=0 pd=0 as=-1.2482e+09 ps=693420 
M3317 Vdd Vdd Vdd GND efet w=3175 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3318 Vdd Vdd Vdd GND efet w=3810 l=8255
+ ad=0 pd=0 as=0 ps=0 
M3319 diff_1018540_320040# Vdd Vdd GND efet w=11430 l=20320
+ ad=0 pd=0 as=0 ps=0 
M3320 diff_2195830_2933700# diff_2089150_548640# GND GND efet w=60960 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3321 diff_1897380_527050# diff_1701800_544830# GND GND efet w=52070 l=7620
+ ad=1.8e+09 pd=411480 as=0 ps=0 
M3322 GND diff_1979930_419100# diff_232410_996950# GND efet w=76200 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3323 GND diff_2192020_525780# diff_755650_927100# GND efet w=45720 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3324 diff_1576070_459740# diff_1576070_459740# diff_1576070_459740# GND efet w=2540 l=6350
+ ad=0 pd=0 as=0 ps=0 
M3325 GND diff_1569720_548640# diff_1604010_461010# GND efet w=47625 l=8255
+ ad=0 pd=0 as=9.72579e+08 ps=213360 
M3326 Vdd Vdd diff_1343660_488950# GND efet w=10795 l=32385
+ ad=0 pd=0 as=0 ps=0 
M3327 diff_1465580_462280# Vdd Vdd GND efet w=10160 l=30480
+ ad=0 pd=0 as=0 ps=0 
M3328 diff_1576070_459740# diff_1576070_459740# diff_1576070_459740# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M3329 diff_1604010_461010# diff_1604010_461010# diff_1604010_461010# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M3330 diff_1518920_467360# Vdd Vdd GND efet w=10160 l=40640
+ ad=0 pd=0 as=0 ps=0 
M3331 diff_1677670_457200# diff_1604010_461010# GND GND efet w=35560 l=8890
+ ad=0 pd=0 as=0 ps=0 
M3332 GND diff_1701800_544830# diff_1720850_440690# GND efet w=48260 l=7620
+ ad=0 pd=0 as=8.0645e+08 ps=182880 
M3333 diff_1677670_457200# diff_1677670_457200# diff_1677670_457200# GND efet w=1905 l=5715
+ ad=0 pd=0 as=0 ps=0 
M3334 diff_1604010_461010# diff_1604010_461010# diff_1604010_461010# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M3335 diff_1677670_457200# diff_1677670_457200# diff_1677670_457200# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M3336 diff_737870_302260# diff_1720850_440690# GND GND efet w=26670 l=7620
+ ad=1.27097e+09 pd=294640 as=0 ps=0 
M3337 GND diff_1465580_462280# diff_737870_302260# GND efet w=34925 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3338 diff_737870_302260# diff_1838960_473710# GND GND efet w=26670 l=8890
+ ad=0 pd=0 as=0 ps=0 
M3339 GND diff_1465580_462280# diff_1897380_527050# GND efet w=33020 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3340 diff_1897380_527050# diff_1894840_476250# GND GND efet w=33655 l=10795
+ ad=0 pd=0 as=0 ps=0 
M3341 diff_737870_302260# diff_737870_302260# diff_737870_302260# GND efet w=2540 l=3175
+ ad=0 pd=0 as=0 ps=0 
M3342 diff_1720850_440690# diff_1720850_440690# diff_1720850_440690# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M3343 diff_737870_302260# diff_737870_302260# diff_737870_302260# GND efet w=2540 l=3175
+ ad=0 pd=0 as=0 ps=0 
M3344 diff_1576070_459740# Vdd Vdd GND efet w=11430 l=30480
+ ad=0 pd=0 as=0 ps=0 
M3345 diff_1720850_440690# diff_1720850_440690# diff_1720850_440690# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M3346 diff_1677670_457200# Vdd Vdd GND efet w=10795 l=33020
+ ad=0 pd=0 as=0 ps=0 
M3347 Vdd Vdd diff_1720850_440690# GND efet w=11430 l=41910
+ ad=0 pd=0 as=0 ps=0 
M3348 Vdd Vdd diff_1604010_461010# GND efet w=10160 l=41910
+ ad=0 pd=0 as=0 ps=0 
M3349 diff_737870_302260# Vdd Vdd GND efet w=10160 l=40640
+ ad=0 pd=0 as=0 ps=0 
M3350 GND diff_2192020_525780# diff_2195830_2933700# GND efet w=57150 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3351 diff_2089150_548640# diff_1897380_186690# GND GND efet w=33020 l=7620
+ ad=7.09676e+08 pd=167640 as=0 ps=0 
M3352 GND diff_2153920_452120# diff_232410_996950# GND efet w=62865 l=12065
+ ad=0 pd=0 as=0 ps=0 
M3353 diff_755650_927100# diff_2014220_425450# GND GND efet w=46990 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3354 GND diff_1838960_473710# diff_1897380_527050# GND efet w=27305 l=8255
+ ad=0 pd=0 as=0 ps=0 
M3355 GND diff_1897380_527050# diff_2014220_425450# GND efet w=22860 l=7620
+ ad=0 pd=0 as=5.29031e+08 ps=106680 
M3356 GND diff_1018540_320040# diff_2192020_525780# GND efet w=40640 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3357 diff_2195830_2933700# diff_2065020_433070# GND GND efet w=60325 l=8255
+ ad=0 pd=0 as=0 ps=0 
M3358 GND diff_1894840_476250# diff_2065020_433070# GND efet w=22860 l=7620
+ ad=0 pd=0 as=4.54838e+08 ps=104140 
M3359 diff_1897380_527050# Vdd Vdd GND efet w=10160 l=39370
+ ad=0 pd=0 as=0 ps=0 
M3360 diff_1979930_419100# diff_737870_302260# GND GND efet w=21590 l=8890
+ ad=5.66128e+08 pd=101600 as=0 ps=0 
M3361 Vdd Vdd diff_1979930_419100# GND efet w=11430 l=53340
+ ad=0 pd=0 as=0 ps=0 
M3362 Vdd Vdd diff_2014220_425450# GND efet w=11430 l=49530
+ ad=0 pd=0 as=0 ps=0 
M3363 diff_2065020_433070# Vdd Vdd GND efet w=11430 l=49530
+ ad=0 pd=0 as=0 ps=0 
M3364 diff_2089150_548640# Vdd Vdd GND efet w=7620 l=24765
+ ad=0 pd=0 as=0 ps=0 
M3365 diff_1018540_320040# clk2 diff_2522220_497840# GND efet w=15240 l=6350
+ ad=0 pd=0 as=2.69354e+08 ps=66040 
M3366 Vdd Vdd Vdd GND efet w=1905 l=2540
+ ad=0 pd=0 as=0 ps=0 
M3367 diff_2496820_474980# Vdd Vdd GND efet w=12065 l=59055
+ ad=7.93547e+08 pd=172720 as=0 ps=0 
M3368 GND diff_2522220_497840# diff_2496820_474980# GND efet w=19050 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3369 Vdd Vdd Vdd GND efet w=3175 l=4445
+ ad=0 pd=0 as=0 ps=0 
M3370 diff_2517140_445770# clk1 diff_2496820_474980# GND efet w=13970 l=7620
+ ad=2.48387e+08 pd=63500 as=0 ps=0 
M3371 GND diff_2517140_445770# diff_699770_264160# GND efet w=53975 l=6985
+ ad=0 pd=0 as=9.37095e+08 ps=185420 
M3372 Vdd Vdd Vdd GND efet w=1905 l=1905
+ ad=0 pd=0 as=0 ps=0 
M3373 Vdd Vdd Vdd GND efet w=3175 l=3810
+ ad=0 pd=0 as=0 ps=0 
M3374 Vdd Vdd Vdd GND efet w=2540 l=6350
+ ad=0 pd=0 as=0 ps=0 
M3375 Vdd Vdd Vdd GND efet w=1270 l=1905
+ ad=0 pd=0 as=0 ps=0 
M3376 diff_1897380_186690# Vdd Vdd GND efet w=11430 l=20320
+ ad=-1.35142e+09 pd=586740 as=0 ps=0 
M3377 diff_699770_264160# Vdd Vdd GND efet w=11430 l=20955
+ ad=0 pd=0 as=0 ps=0 
M3378 Vdd Vdd diff_1037590_429260# GND efet w=11430 l=29210
+ ad=0 pd=0 as=8.46772e+08 ps=185420 
M3379 Vdd Vdd diff_2268220_171450# GND efet w=13970 l=47625
+ ad=0 pd=0 as=9.74192e+08 ps=205740 
M3380 diff_1897380_186690# reset GND GND efet w=133350 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3381 sync GND GND GND efet w=111760 l=8890
+ ad=0 pd=0 as=0 ps=0 
M3382 reset GND GND GND efet w=114300 l=8890
+ ad=-3.36911e+08 pd=817880 as=0 ps=0 
M3383 GND GND p0 GND efet w=111760 l=8890
+ ad=0 pd=0 as=-8.07878e+08 ps=792480 
M3384 diff_2268220_171450# diff_2268220_171450# diff_2268220_171450# GND efet w=3175 l=3175
+ ad=0 pd=0 as=0 ps=0 
M3385 diff_2268220_171450# diff_2268220_171450# diff_2268220_171450# GND efet w=1905 l=5715
+ ad=0 pd=0 as=0 ps=0 
M3386 diff_1037590_429260# diff_2268220_171450# GND GND efet w=40640 l=6350
+ ad=0 pd=0 as=0 ps=0 
M3387 GND cm diff_2268220_171450# GND efet w=53340 l=7620
+ ad=0 pd=0 as=0 ps=0 
M3388 cm GND GND GND efet w=112395 l=8255
+ ad=-5.12717e+08 pd=822960 as=0 ps=0 
C0 metal_2552700_43180# gnd! 48.4fF ;**FLOATING
C1 metal_2494280_52070# gnd! 51.6fF ;**FLOATING
C2 metal_2435860_54610# gnd! 54.0fF ;**FLOATING
C3 metal_2377440_66040# gnd! 47.5fF ;**FLOATING
C4 metal_736600_58420# gnd! 7.6fF ;**FLOATING
C5 metal_715010_67310# gnd! 4.3fF ;**FLOATING
C6 metal_698500_81280# gnd! 12.0fF ;**FLOATING
C7 metal_713740_81280# gnd! 29.7fF ;**FLOATING
C8 metal_759460_118110# gnd! 85.0fF ;**FLOATING
C9 metal_165100_171450# gnd! 9.8fF ;**FLOATING
C10 metal_2491740_3122930# gnd! 60.4fF ;**FLOATING
C11 diff_2268220_171450# gnd! 148.2fF
C12 cm gnd! 651.4fF
C13 reset gnd! 684.4fF
C14 diff_2517140_445770# gnd! 82.0fF
C15 diff_2496820_474980# gnd! 96.5fF
C16 diff_2522220_497840# gnd! 70.4fF
C17 diff_2065020_433070# gnd! 207.7fF
C18 diff_1720850_440690# gnd! 155.2fF
C19 diff_1979930_419100# gnd! 187.4fF
C20 diff_1897380_527050# gnd! 342.3fF
C21 diff_2192020_525780# gnd! 156.1fF
C22 diff_2089150_548640# gnd! 214.2fF
C23 diff_2517140_586740# gnd! 78.6fF
C24 diff_2541270_668020# gnd! 75.8fF
C25 diff_1416050_494030# gnd! 115.6fF
C26 diff_1343660_488950# gnd! 108.7fF
C27 diff_1465580_462280# gnd! 383.8fF
C28 diff_1701800_544830# gnd! 236.7fF
C29 diff_1604010_461010# gnd! 313.6fF
C30 diff_2203450_571500# gnd! 142.8fF
C31 diff_1518920_467360# gnd! 310.8fF
C32 diff_2124710_610870# gnd! 134.2fF
C33 diff_2014220_425450# gnd! 362.8fF
C34 diff_2536190_745490# gnd! 82.9fF
C35 diff_2153920_452120# gnd! 938.5fF
C36 diff_2320290_678180# gnd! 282.3fF
C37 diff_2245360_692150# gnd! 201.7fF
C38 diff_2228850_712470# gnd! 199.4fF
C39 diff_2555240_824230# gnd! 81.3fF
C40 diff_2324100_800100# gnd! 206.2fF
C41 diff_2246630_834390# gnd! 136.9fF
C42 diff_2297430_869950# gnd! 150.8fF
C43 diff_2559050_902970# gnd! 80.5fF
C44 diff_2247900_798830# gnd! 269.1fF
C45 diff_1894840_476250# gnd! 413.9fF
C46 diff_1569720_548640# gnd! 104.6fF
C47 diff_1118870_429260# gnd! 39.6fF
C48 diff_1101090_427990# gnd! 42.2fF
C49 diff_1111250_266700# gnd! 567.4fF
C50 diff_1027430_431800# gnd! 54.5fF
C51 diff_1007110_440690# gnd! 57.5fF
C52 diff_622300_264160# gnd! 148.8fF
C53 diff_647700_243840# gnd! 125.1fF
C54 diff_737870_302260# gnd! 635.0fF
C55 diff_664210_320040# gnd! 39.0fF
C56 diff_172720_179070# gnd! 15.2fF ;**FLOATING
C57 diff_167640_190500# gnd! 20.7fF ;**FLOATING
C58 diff_163830_198120# gnd! 112.6fF ;**FLOATING
C59 diff_581660_321310# gnd! 157.6fF
C60 diff_1018540_320040# gnd! 965.5fF
C61 diff_924560_458470# gnd! 155.6fF
C62 diff_1239520_500380# gnd! 36.8fF
C63 diff_699770_264160# gnd! 553.4fF
C64 diff_1183640_483870# gnd! 93.3fF
C65 diff_1239520_518160# gnd! 43.0fF
C66 diff_1239520_481330# gnd! 147.4fF
C67 diff_1037590_429260# gnd! 666.9fF
C68 diff_1507490_548640# gnd! 89.5fF
C69 diff_1838960_473710# gnd! 302.6fF
C70 diff_1681480_645160# gnd! 83.1fF
C71 diff_1736090_635000# gnd! 135.8fF
C72 diff_1149350_486410# gnd! 151.3fF
C73 diff_900430_483870# gnd! 635.2fF
C74 diff_1997710_690880# gnd! 122.3fF
C75 diff_1997710_740410# gnd! 254.6fF
C76 diff_2123440_789940# gnd! 100.3fF
C77 diff_2077720_787400# gnd! 114.4fF
C78 diff_1960880_777240# gnd! 109.2fF
C79 diff_1973580_749300# gnd! 116.2fF
C80 diff_2053590_824230# gnd! 109.6fF
C81 diff_1983740_830580# gnd! 233.8fF
C82 diff_1974850_806450# gnd! 278.0fF
C83 diff_1831340_789940# gnd! 99.3fF
C84 diff_1894840_732790# gnd! 170.7fF
C85 diff_1786890_783590# gnd! 111.0fF
C86 diff_434340_266700# gnd! 280.5fF
C87 diff_438150_274320# gnd! 58.5fF
C88 diff_387350_243840# gnd! 117.6fF
C89 diff_487680_288290# gnd! 115.8fF
C90 diff_505460_347980# gnd! 221.1fF
C91 diff_358140_298450# gnd! 131.9fF
C92 diff_857250_500380# gnd! 210.0fF
C93 diff_821690_471170# gnd! 118.3fF
C94 diff_694690_422910# gnd! 125.6fF
C95 diff_772160_488950# gnd! 146.4fF
C96 p0 gnd! 1236.7fF
C97 diff_328930_492760# gnd! 104.4fF
C98 diff_325120_504190# gnd! 80.7fF
C99 diff_377190_510540# gnd! 83.1fF
C100 diff_787400_546100# gnd! 153.8fF
C101 diff_373380_521970# gnd! 60.6fF
C102 diff_302260_482600# gnd! 76.4fF
C103 diff_582930_558800# gnd! 136.1fF
C104 diff_640080_426720# gnd! 248.0fF
C105 diff_775970_467360# gnd! 224.5fF
C106 diff_669290_508000# gnd! 361.1fF
C107 diff_377190_574040# gnd! 91.4fF
C108 diff_586740_528320# gnd! 522.5fF
C109 diff_374650_585470# gnd! 60.2fF
C110 diff_586740_566420# gnd! 229.8fF
C111 diff_377190_637540# gnd! 85.5fF
C112 diff_1018540_712470# gnd! 602.9fF
C113 diff_1681480_749300# gnd! 118.4fF
C114 diff_1670050_753110# gnd! 106.7fF
C115 diff_1922780_786130# gnd! 141.0fF
C116 diff_1761490_825500# gnd! 108.8fF
C117 diff_1692910_830580# gnd! 427.3fF
C118 diff_1682750_806450# gnd! 423.4fF
C119 diff_1600200_718820# gnd! 175.0fF
C120 diff_1539240_795020# gnd! 104.9fF
C121 diff_1494790_784860# gnd! 119.3fF
C122 diff_1379220_753110# gnd! 107.8fF
C123 diff_1390650_749300# gnd! 122.0fF
C124 diff_1630680_786130# gnd! 142.4fF
C125 diff_2315210_670560# gnd! 542.8fF
C126 diff_2578100_981710# gnd! 72.0fF
C127 diff_1470660_825500# gnd! 107.3fF
C128 diff_1402080_830580# gnd! 433.6fF
C129 diff_1391920_806450# gnd! 423.2fF
C130 diff_1313180_713740# gnd! 183.1fF
C131 diff_1248410_791210# gnd! 107.5fF
C132 diff_1203960_786130# gnd! 118.9fF
C133 diff_1099820_749300# gnd! 126.7fF
C134 diff_1087120_770890# gnd! 110.2fF
C135 diff_1339850_786130# gnd! 131.3fF
C136 diff_1677670_457200# gnd! 444.6fF
C137 diff_1576070_459740# gnd! 659.9fF
C138 diff_1982470_873760# gnd! 329.8fF
C139 diff_1790700_659130# gnd! 290.6fF
C140 diff_1178560_825500# gnd! 113.9fF
C141 diff_1111250_830580# gnd! 434.9fF
C142 diff_1099820_863600# gnd! 429.8fF
C143 diff_1022350_718820# gnd! 177.5fF
C144 diff_957580_789940# gnd! 107.4fF
C145 diff_913130_783590# gnd! 119.4fF
C146 diff_374650_646430# gnd! 65.7fF
C147 diff_401320_678180# gnd! 88.5fF
C148 diff_808990_749300# gnd! 120.8fF
C149 diff_576580_742950# gnd! 107.7fF
C150 diff_400050_777240# gnd! 69.1fF
C151 sync gnd! 1439.9fF
C152 diff_798830_753110# gnd! 94.9fF
C153 diff_1005840_731520# gnd! 795.5fF
C154 diff_1049020_786130# gnd! 131.3fF
C155 diff_419100_734060# gnd! 237.9fF
C156 diff_575310_779780# gnd! 328.3fF
C157 diff_887730_825500# gnd! 117.0fF
C158 diff_820420_830580# gnd! 432.7fF
C159 diff_808990_863600# gnd! 424.5fF
C160 diff_408940_681990# gnd! 802.4fF
C161 diff_1691640_873760# gnd! 429.0fF
C162 diff_1400810_873760# gnd! 284.7fF
C163 diff_3810_849630# gnd! 1393.1fF ;**FLOATING
C164 diff_251460_913130# gnd! 120.4fF
C165 diff_1888490_857250# gnd! 399.4fF
C166 diff_1513840_989330# gnd! 321.4fF
C167 diff_1103630_871220# gnd! 663.5fF
C168 diff_812800_871220# gnd! 447.0fF
C169 diff_1223010_990600# gnd! 313.9fF
C170 diff_932180_1002030# gnd! 324.9fF
C171 diff_2578100_1071880# gnd! 78.9fF
C172 diff_1882140_1065530# gnd! 87.5fF
C173 diff_1799590_1065530# gnd! 65.3fF
C174 diff_1877060_1057910# gnd! 239.8fF
C175 diff_2534920_1196340# gnd! 145.9fF
C176 diff_1988820_1080770# gnd! 233.1fF
C177 diff_897890_1024890# gnd! 1183.8fF
C178 diff_2138680_1156970# gnd! 163.2fF
C179 diff_932180_1050290# gnd! 1026.4fF
C180 diff_2085340_1167130# gnd! 154.4fF
C181 diff_2000250_1186180# gnd! 166.6fF
C182 diff_1925320_1167130# gnd! 147.5fF
C183 diff_1869440_1156970# gnd! 148.7fF
C184 diff_1793240_1167130# gnd! 147.9fF
C185 diff_1728470_1183640# gnd! 165.1fF
C186 diff_1483360_1032510# gnd! 186.4fF
C187 diff_1647190_1168400# gnd! 161.4fF
C188 diff_1583690_1181100# gnd! 166.2fF
C189 diff_2463800_1235710# gnd! 118.4fF
C190 diff_1795780_1076960# gnd! 378.9fF
C191 diff_1502410_1167130# gnd! 163.8fF
C192 diff_1437640_1181100# gnd! 165.7fF
C193 diff_1356360_1168400# gnd! 160.5fF
C194 diff_1292860_1186180# gnd! 163.8fF
C195 diff_1192530_1032510# gnd! 198.4fF
C196 diff_1211580_1167130# gnd! 163.7fF
C197 diff_1146810_1183640# gnd! 166.9fF
C198 diff_1066800_1167130# gnd! 162.4fF
C199 diff_1003300_1182370# gnd! 163.0fF
C200 diff_872490_1087120# gnd! 170.0fF
C201 diff_608330_1127760# gnd! 158.2fF
C202 diff_232410_1049020# gnd! 205.9fF
C203 diff_237490_1127760# gnd! 162.6fF
C204 diff_594360_1112520# gnd! 139.9fF
C205 diff_920750_1167130# gnd! 167.4fF
C206 diff_214630_541020# gnd! 600.7fF
C207 diff_855980_1183640# gnd! 166.1fF
C208 diff_608330_1151890# gnd! 155.7fF
C209 diff_599440_977900# gnd! 892.9fF
C210 diff_262890_1151890# gnd! 75.6fF
C211 diff_232410_1165860# gnd! 78.1fF
C212 diff_1998980_1291590# gnd! 435.1fF
C213 diff_2475230_1280160# gnd! 184.6fF
C214 diff_934720_1277620# gnd! 659.4fF
C215 diff_869950_1299210# gnd! 686.7fF
C216 diff_2089150_1318260# gnd! 309.8fF
C217 diff_2443480_1254760# gnd! 166.9fF
C218 diff_889000_1079500# gnd! 887.6fF
C219 diff_546100_1313180# gnd! 198.1fF
C220 diff_2075180_1344930# gnd! 381.9fF
C221 diff_869950_1347470# gnd! 725.9fF
C222 diff_546100_1341120# gnd! 235.3fF
C223 diff_2012950_1370330# gnd! 319.3fF
C224 diff_2439670_1344930# gnd! 133.9fF
C225 diff_1160780_1371600# gnd! 704.8fF
C226 diff_2197100_1388110# gnd! 159.6fF
C227 diff_869950_1397000# gnd! 686.8fF
C228 diff_546100_1388110# gnd! 231.4fF
C229 diff_774700_1325880# gnd! 105.9fF
C230 diff_232410_996950# gnd! 1546.2fF
C231 diff_2471420_1322070# gnd! 217.0fF
C232 diff_2444750_1443990# gnd! 282.6fF
C233 diff_829310_237490# gnd! 1087.7fF
C234 diff_2486660_1535430# gnd! 130.2fF
C235 diff_284480_472440# gnd! 1058.2fF
C236 diff_872490_1417320# gnd! 600.4fF
C237 diff_1377950_1109980# gnd! 522.7fF
C238 diff_546100_1416050# gnd! 216.4fF
C239 diff_180340_1348740# gnd! 266.4fF
C240 diff_2172970_1249680# gnd! 458.0fF
C241 diff_2128520_1299210# gnd! 459.7fF
C242 diff_2228850_1562100# gnd! 142.1fF
C243 diff_2080260_1351280# gnd! 399.6fF
C244 diff_2002790_1228090# gnd! 404.1fF
C245 diff_2156460_1504950# gnd! 142.7fF
C246 diff_2082800_1562100# gnd! 140.0fF
C247 diff_1926590_1210310# gnd! 471.8fF
C248 diff_1861820_1186180# gnd! 449.3fF
C249 diff_2010410_1504950# gnd! 148.7fF
C250 diff_1936750_1562100# gnd! 143.1fF
C251 diff_1790700_1535430# gnd! 426.3fF
C252 diff_1729740_1228090# gnd! 405.4fF
C253 diff_1864360_1504950# gnd! 147.6fF
C254 diff_1790700_1562100# gnd! 147.7fF
C255 diff_1645920_1535430# gnd! 408.4fF
C256 diff_1584960_1226820# gnd! 376.7fF
C257 diff_1719580_1478280# gnd! 144.7fF
C258 diff_1645920_1562100# gnd! 144.3fF
C259 diff_1499870_1535430# gnd! 402.5fF
C260 diff_1438910_1226820# gnd! 403.8fF
C261 diff_1573530_1504950# gnd! 148.2fF
C262 diff_1499870_1562100# gnd! 147.5fF
C263 diff_1428750_1470660# gnd! 145.8fF
C264 diff_1355090_1535430# gnd! 393.2fF
C265 diff_1292860_1226820# gnd! 401.2fF
C266 diff_1355090_1562100# gnd! 147.6fF
C267 diff_1209040_1535430# gnd! 399.7fF
C268 diff_1148080_1228090# gnd! 402.5fF
C269 diff_1282700_1504950# gnd! 148.5fF
C270 diff_1209040_1562100# gnd! 147.8fF
C271 diff_1064260_1535430# gnd! 397.3fF
C272 diff_1002030_1186180# gnd! 395.6fF
C273 diff_1137920_1470660# gnd! 148.3fF
C274 diff_1064260_1562100# gnd! 143.3fF
C275 diff_172720_1316990# gnd! 274.8fF
C276 diff_868680_1503680# gnd! 1882.4fF
C277 diff_894080_1518920# gnd! 1487.7fF
C278 diff_918210_1536700# gnd! 400.9fF
C279 diff_857250_1226820# gnd! 402.4fF
C280 diff_774700_1455420# gnd! 120.6fF
C281 diff_755650_927100# gnd! 1527.5fF
C282 diff_991870_1504950# gnd! 148.2fF
C283 diff_918210_1562100# gnd! 146.0fF
C284 diff_844550_1507490# gnd! 153.4fF
C285 diff_2482850_1590040# gnd! 172.7fF
C286 diff_2476500_1567180# gnd! 212.1fF
C287 clk1 gnd! 2154.0fF
C288 diff_2268220_1647190# gnd! 36.6fF
C289 diff_2479040_1628140# gnd! 199.0fF
C290 diff_2241550_1626870# gnd! 77.5fF
C291 diff_2268220_1681480# gnd! 36.6fF
C292 diff_2415540_1699260# gnd! 128.4fF
C293 diff_2171700_1642110# gnd! 32.4fF
C294 diff_2160270_1626870# gnd! 78.1fF
C295 diff_2095500_1626870# gnd! 76.8fF
C296 diff_2122170_1647190# gnd! 35.5fF
C297 diff_2241550_1715770# gnd! 76.5fF
C298 diff_2241550_1775460# gnd! 77.4fF
C299 diff_2268220_1797050# gnd! 36.9fF
C300 diff_1897380_186690# gnd! 884.9fF
C301 diff_2268220_1831340# gnd! 37.8fF
C302 diff_2171700_1685290# gnd! 33.6fF
C303 diff_2122170_1681480# gnd! 36.9fF
C304 diff_2160270_1714500# gnd! 78.4fF
C305 diff_2025650_1640840# gnd! 33.7fF
C306 diff_2014220_1626870# gnd! 80.7fF
C307 diff_1950720_1625600# gnd! 77.6fF
C308 diff_1976120_1647190# gnd! 37.2fF
C309 diff_2095500_1715770# gnd! 76.3fF
C310 diff_2171700_1790700# gnd! 33.4fF
C311 diff_2160270_1776730# gnd! 78.0fF
C312 diff_2095500_1775460# gnd! 77.6fF
C313 diff_2122170_1797050# gnd! 37.2fF
C314 diff_2241550_1866900# gnd! 77.0fF
C315 diff_2241550_1926590# gnd! 78.3fF
C316 diff_2268220_1946910# gnd! 37.1fF
C317 diff_2268220_1982470# gnd! 36.9fF
C318 o3 gnd! 614.9fF
C319 diff_2171700_1835150# gnd! 33.6fF
C320 diff_2122170_1831340# gnd! 37.5fF
C321 diff_2160270_1864360# gnd! 80.1fF
C322 diff_2025650_1685290# gnd! 33.9fF
C323 diff_1976120_1681480# gnd! 37.1fF
C324 diff_2014220_1714500# gnd! 78.1fF
C325 diff_1879600_1640840# gnd! 34.1fF
C326 diff_1868170_1628140# gnd! 79.6fF
C327 diff_1831340_1645920# gnd! 34.2fF
C328 diff_1804670_1625600# gnd! 77.7fF
C329 diff_1950720_1715770# gnd! 75.7fF
C330 diff_2025650_1790700# gnd! 34.1fF
C331 diff_2014220_1776730# gnd! 78.3fF
C332 diff_1950720_1775460# gnd! 76.3fF
C333 diff_1976120_1797050# gnd! 37.5fF
C334 diff_2095500_1866900# gnd! 77.6fF
C335 diff_2171700_1941830# gnd! 33.6fF
C336 diff_2122170_1946910# gnd! 37.1fF
C337 diff_2160270_1926590# gnd! 77.8fF
C338 diff_2095500_1926590# gnd! 76.3fF
C339 diff_2241550_2016760# gnd! 75.2fF
C340 diff_2241550_2076450# gnd! 75.8fF
C341 diff_2268220_2098040# gnd! 37.2fF
C342 diff_2513330_2120900# gnd! 248.0fF
C343 diff_2598420_2186940# gnd! 89.2fF
C344 diff_2566670_2211070# gnd! 78.7fF
C345 diff_2268220_2132330# gnd! 37.5fF
C346 diff_2171700_1985010# gnd! 32.5fF
C347 diff_2122170_1982470# gnd! 37.2fF
C348 diff_2160270_2014220# gnd! 76.3fF
C349 diff_2025650_1835150# gnd! 33.9fF
C350 diff_1976120_1831340# gnd! 37.6fF
C351 diff_2014220_1864360# gnd! 78.3fF
C352 diff_1879600_1685290# gnd! 34.1fF
C353 diff_1831340_1681480# gnd! 34.1fF
C354 diff_1868170_1715770# gnd! 77.1fF
C355 diff_1733550_1640840# gnd! 34.5fF
C356 diff_1685290_1645920# gnd! 34.0fF
C357 diff_1723390_1626870# gnd! 77.7fF
C358 diff_1658620_1625600# gnd! 81.0fF
C359 diff_1804670_1715770# gnd! 74.4fF
C360 diff_1733550_1685290# gnd! 34.6fF
C361 diff_1685290_1681480# gnd! 34.1fF
C362 diff_1723390_1714500# gnd! 75.8fF
C363 diff_1879600_1790700# gnd! 34.1fF
C364 diff_1868170_1776730# gnd! 77.0fF
C365 diff_1804670_1775460# gnd! 75.6fF
C366 diff_1831340_1795780# gnd! 34.2fF
C367 diff_1950720_1865630# gnd! 78.4fF
C368 diff_2025650_1941830# gnd! 34.1fF
C369 diff_1950720_1925320# gnd! 77.6fF
C370 diff_1976120_1946910# gnd! 37.4fF
C371 diff_2014220_1926590# gnd! 78.0fF
C372 diff_2095500_2016760# gnd! 77.2fF
C373 diff_2171700_2091690# gnd! 33.9fF
C374 diff_2160270_2076450# gnd! 76.0fF
C375 diff_2122170_2098040# gnd! 36.9fF
C376 diff_2095500_2076450# gnd! 76.6fF
C377 diff_2241550_2167890# gnd! 76.1fF
C378 diff_2268220_2247900# gnd! 37.1fF
C379 diff_2481580_2265680# gnd! 346.0fF
C380 diff_2461260_2273300# gnd! 38.3fF
C381 diff_2241550_2227580# gnd! 76.9fF
C382 diff_2557780_2068830# gnd! 440.2fF
C383 diff_2268220_2283460# gnd! 36.1fF
C384 diff_2171700_2136140# gnd! 33.6fF
C385 diff_2122170_2132330# gnd! 37.5fF
C386 diff_2160270_2164080# gnd! 76.7fF
C387 diff_2025650_1985010# gnd! 35.2fF
C388 diff_1976120_1981200# gnd! 38.3fF
C389 diff_2014220_2014220# gnd! 78.0fF
C390 diff_1879600_1835150# gnd! 34.5fF
C391 diff_1831340_1831340# gnd! 32.6fF
C392 diff_1868170_1865630# gnd! 79.1fF
C393 diff_1588770_1642110# gnd! 34.1fF
C394 diff_1577340_1626870# gnd! 81.9fF
C395 diff_1539240_1647190# gnd! 36.8fF
C396 diff_1513840_1625600# gnd! 77.5fF
C397 diff_1658620_1715770# gnd! 77.9fF
C398 diff_1733550_1790700# gnd! 34.2fF
C399 diff_1723390_1775460# gnd! 76.0fF
C400 diff_1685290_1795780# gnd! 33.8fF
C401 diff_1658620_1775460# gnd! 79.3fF
C402 diff_1733550_1835150# gnd! 36.1fF
C403 diff_1804670_1866900# gnd! 77.1fF
C404 diff_1685290_1831340# gnd! 34.5fF
C405 diff_1723390_1863090# gnd! 77.3fF
C406 diff_1879600_1940560# gnd! 34.8fF
C407 diff_1868170_1929130# gnd! 78.6fF
C408 diff_1804670_1925320# gnd! 77.0fF
C409 diff_1831340_1945640# gnd! 34.8fF
C410 diff_1950720_2016760# gnd! 76.6fF
C411 diff_2025650_2091690# gnd! 33.8fF
C412 diff_2014220_2076450# gnd! 76.6fF
C413 diff_1950720_2076450# gnd! 76.0fF
C414 diff_1976120_2098040# gnd! 37.5fF
C415 diff_2095500_2166620# gnd! 75.9fF
C416 diff_2171700_2242820# gnd! 33.6fF
C417 diff_2122170_2247900# gnd! 36.9fF
C418 diff_2160270_2226310# gnd! 77.8fF
C419 diff_2095500_2227580# gnd! 78.1fF
C420 diff_2241550_2317750# gnd! 75.6fF
C421 diff_2241550_2376170# gnd! 76.3fF
C422 diff_2268220_2397760# gnd! 36.4fF
C423 diff_2268220_2432050# gnd! 37.5fF
C424 diff_2171700_2286000# gnd! 32.5fF
C425 diff_2122170_2283460# gnd! 36.4fF
C426 diff_2160270_2315210# gnd! 78.0fF
C427 diff_2025650_2136140# gnd! 33.9fF
C428 diff_1976120_2132330# gnd! 37.5fF
C429 diff_2014220_2164080# gnd! 78.4fF
C430 diff_1879600_1985010# gnd! 35.3fF
C431 diff_1831340_1981200# gnd! 35.2fF
C432 diff_1868170_2015490# gnd! 76.1fF
C433 diff_1588770_1685290# gnd! 33.7fF
C434 diff_1539240_1681480# gnd! 37.2fF
C435 diff_1577340_1714500# gnd! 80.2fF
C436 diff_1442720_1642110# gnd! 33.6fF
C437 diff_1432560_1626870# gnd! 79.3fF
C438 diff_1367790_1625600# gnd! 80.0fF
C439 diff_1394460_1645920# gnd! 34.2fF
C440 diff_1513840_1715770# gnd! 77.0fF
C441 diff_1588770_1790700# gnd! 34.0fF
C442 diff_1577340_1775460# gnd! 78.7fF
C443 diff_1513840_1775460# gnd! 75.6fF
C444 diff_1539240_1795780# gnd! 37.1fF
C445 diff_1658620_1866900# gnd! 80.8fF
C446 diff_1733550_1940560# gnd! 37.7fF
C447 diff_1723390_1925320# gnd! 76.8fF
C448 diff_1658620_1925320# gnd! 79.7fF
C449 diff_1685290_1945640# gnd! 34.7fF
C450 diff_1804670_2015490# gnd! 77.3fF
C451 diff_1879600_2091690# gnd! 34.3fF
C452 diff_1869440_2075180# gnd! 77.3fF
C453 diff_1804670_2076450# gnd! 74.0fF
C454 diff_1831340_2096770# gnd! 34.5fF
C455 diff_1950720_2166620# gnd! 76.8fF
C456 diff_2025650_2242820# gnd! 33.9fF
C457 diff_2014220_2226310# gnd! 77.9fF
C458 diff_1950720_2226310# gnd! 76.7fF
C459 diff_1976120_2247900# gnd! 37.1fF
C460 diff_2095500_2317750# gnd! 76.5fF
C461 diff_2171700_2391410# gnd! 33.5fF
C462 diff_2160270_2377440# gnd! 78.3fF
C463 diff_2122170_2397760# gnd! 37.2fF
C464 diff_2095500_2376170# gnd! 77.5fF
C465 diff_2241550_2466340# gnd! 75.7fF
C466 diff_2241550_2526030# gnd! 75.8fF
C467 diff_2268220_2547620# gnd! 37.2fF
C468 o2 gnd! 734.1fF
C469 diff_2513330_2576830# gnd! 244.0fF
C470 diff_2268220_2581910# gnd! 37.1fF
C471 diff_2598420_2640330# gnd! 86.1fF
C472 diff_2565400_2665730# gnd! 84.1fF
C473 diff_2171700_2435860# gnd! 33.6fF
C474 diff_2122170_2432050# gnd! 37.5fF
C475 diff_2160270_2465070# gnd! 77.4fF
C476 diff_2025650_2286000# gnd! 33.6fF
C477 diff_1976120_2282190# gnd! 37.0fF
C478 diff_2014220_2315210# gnd! 77.1fF
C479 diff_1831340_2132330# gnd! 32.1fF
C480 diff_1879600_2136140# gnd! 34.5fF
C481 diff_1869440_2164080# gnd! 77.7fF
C482 diff_1733550_1985010# gnd! 38.4fF
C483 diff_1685290_1981200# gnd! 35.3fF
C484 diff_1723390_2014220# gnd! 75.3fF
C485 diff_1588770_1835150# gnd! 33.7fF
C486 diff_1539240_1831340# gnd! 37.2fF
C487 diff_1577340_1864360# gnd! 79.9fF
C488 diff_1442720_1685290# gnd! 33.7fF
C489 diff_1394460_1681480# gnd! 34.1fF
C490 diff_1432560_1714500# gnd! 78.7fF
C491 diff_1442720_1790700# gnd! 34.1fF
C492 diff_1432560_1775460# gnd! 77.4fF
C493 diff_1297940_1640840# gnd! 34.7fF
C494 diff_1286510_1626870# gnd! 81.1fF
C495 diff_1249680_1644650# gnd! 34.7fF
C496 diff_1223010_1625600# gnd! 78.0fF
C497 diff_1367790_1715770# gnd! 79.3fF
C498 diff_1367790_1775460# gnd! 76.9fF
C499 diff_1394460_1795780# gnd! 34.4fF
C500 diff_1513840_1866900# gnd! 76.8fF
C501 diff_1442720_1835150# gnd! 33.9fF
C502 diff_1394460_1831340# gnd! 34.5fF
C503 diff_1432560_1863090# gnd! 78.3fF
C504 diff_1588770_1941830# gnd! 34.0fF
C505 diff_1577340_1925320# gnd! 79.0fF
C506 diff_1513840_1925320# gnd! 77.9fF
C507 diff_1539240_1946910# gnd! 37.2fF
C508 diff_1658620_2015490# gnd! 79.8fF
C509 diff_1733550_2091690# gnd! 36.8fF
C510 diff_1723390_2076450# gnd! 74.3fF
C511 diff_1685290_2096770# gnd! 33.8fF
C512 diff_1658620_2076450# gnd! 79.3fF
C513 diff_1804670_2166620# gnd! 75.5fF
C514 diff_1879600_2241550# gnd! 34.7fF
C515 diff_1868170_2232660# gnd! 77.1fF
C516 diff_1804670_2226310# gnd! 75.2fF
C517 diff_1831340_2246630# gnd! 35.0fF
C518 diff_1950720_2316480# gnd! 75.9fF
C519 diff_2025650_2391410# gnd! 34.1fF
C520 diff_2014220_2377440# gnd! 79.0fF
C521 diff_1949450_2382520# gnd! 77.8fF
C522 diff_1976120_2397760# gnd! 36.9fF
C523 diff_2095500_2466340# gnd! 76.4fF
C524 diff_2171700_2542540# gnd! 32.2fF
C525 diff_2160270_2526030# gnd! 77.7fF
C526 diff_2095500_2526030# gnd! 76.7fF
C527 diff_2122170_2547620# gnd! 36.4fF
C528 diff_2241550_2616200# gnd! 74.8fF
C529 diff_2241550_2675890# gnd! 76.0fF
C530 diff_2268220_2697480# gnd! 30.4fF
C531 diff_2481580_2720340# gnd! 342.0fF
C532 diff_2461260_2726690# gnd! 38.6fF
C533 diff_2555240_2753360# gnd! 433.6fF
C534 diff_2354580_1676400# gnd! 888.0fF
C535 diff_2268220_2731770# gnd! 38.2fF
C536 diff_2170430_2599690# gnd! 34.4fF
C537 diff_2122170_2581910# gnd! 37.3fF
C538 diff_2160270_2614930# gnd! 76.5fF
C539 diff_2025650_2435860# gnd! 33.9fF
C540 diff_1976120_2432050# gnd! 37.6fF
C541 diff_2014220_2465070# gnd! 77.3fF
C542 diff_1879600_2286000# gnd! 34.1fF
C543 diff_1830070_2284730# gnd! 34.9fF
C544 diff_1868170_2316480# gnd! 76.6fF
C545 diff_1733550_2136140# gnd! 37.6fF
C546 diff_1685290_2132330# gnd! 34.5fF
C547 diff_1723390_2164080# gnd! 75.9fF
C548 diff_1588770_1985010# gnd! 35.0fF
C549 diff_1539240_1981200# gnd! 38.6fF
C550 diff_1577340_2014220# gnd! 78.6fF
C551 diff_1297940_1685290# gnd! 33.9fF
C552 diff_1249680_1681480# gnd! 33.8fF
C553 diff_1286510_1714500# gnd! 80.6fF
C554 diff_1151890_1640840# gnd! 36.0fF
C555 diff_1103630_1645920# gnd! 35.0fF
C556 diff_1141730_1626870# gnd! 79.8fF
C557 diff_1078230_1617980# gnd! 80.1fF
C558 diff_1223010_1715770# gnd! 77.6fF
C559 diff_1151890_1685290# gnd! 33.9fF
C560 diff_1103630_1681480# gnd! 34.1fF
C561 diff_1141730_1714500# gnd! 78.9fF
C562 diff_1297940_1790700# gnd! 34.7fF
C563 diff_1286510_1775460# gnd! 78.8fF
C564 diff_1223010_1775460# gnd! 76.6fF
C565 diff_1249680_1793240# gnd! 34.1fF
C566 diff_1367790_1866900# gnd! 76.8fF
C567 diff_1442720_1941830# gnd! 34.1fF
C568 diff_1432560_1925320# gnd! 78.4fF
C569 diff_1367790_1926590# gnd! 78.7fF
C570 diff_1394460_1945640# gnd! 34.1fF
C571 diff_1513840_2015490# gnd! 76.9fF
C572 diff_1442720_1985010# gnd! 35.3fF
C573 diff_1394460_1981200# gnd! 32.9fF
C574 diff_1432560_2014220# gnd! 77.6fF
C575 diff_1588770_2091690# gnd! 33.8fF
C576 diff_1577340_2076450# gnd! 78.1fF
C577 diff_1539240_2096770# gnd! 37.2fF
C578 diff_1513840_2075180# gnd! 78.4fF
C579 diff_1658620_2166620# gnd! 78.7fF
C580 diff_1733550_2242820# gnd! 35.7fF
C581 diff_1723390_2226310# gnd! 76.2fF
C582 diff_1658620_2226310# gnd! 79.0fF
C583 diff_1685290_2246630# gnd! 34.1fF
C584 diff_1685290_2282190# gnd! 33.9fF
C585 diff_1733550_2286000# gnd! 34.3fF
C586 diff_1804670_2316480# gnd! 74.7fF
C587 diff_1723390_2315210# gnd! 75.4fF
C588 diff_1879600_2391410# gnd! 33.9fF
C589 diff_1868170_2377440# gnd! 77.4fF
C590 diff_1804670_2376170# gnd! 77.8fF
C591 diff_1830070_2396490# gnd! 36.5fF
C592 diff_1949450_2470150# gnd! 75.5fF
C593 diff_2025650_2541270# gnd! 34.2fF
C594 diff_2014220_2526030# gnd! 76.9fF
C595 diff_1949450_2528570# gnd! 76.5fF
C596 diff_1976120_2547620# gnd! 37.0fF
C597 diff_2095500_2616200# gnd! 76.0fF
C598 diff_2171700_2691130# gnd! 34.4fF
C599 diff_2160270_2675890# gnd! 77.6fF
C600 diff_2095500_2675890# gnd! 76.3fF
C601 diff_2122170_2697480# gnd! 37.3fF
C602 diff_2258060_1543050# gnd! 553.3fF
C603 diff_2233930_1543050# gnd! 512.1fF
C604 diff_2203450_1583690# gnd! 516.4fF
C605 diff_2171700_2735580# gnd! 33.6fF
C606 diff_2122170_2731770# gnd! 37.3fF
C607 diff_2165350_1529080# gnd! 552.9fF
C608 diff_2241550_2767330# gnd! 74.2fF
C609 diff_2160270_2764790# gnd! 75.1fF
C610 diff_2110740_1545590# gnd! 554.8fF
C611 diff_2025650_2585720# gnd! 33.9fF
C612 diff_1976120_2581910# gnd! 37.6fF
C613 diff_2014220_2614930# gnd! 76.5fF
C614 diff_1879600_2435860# gnd! 34.2fF
C615 diff_1830070_2432050# gnd! 37.0fF
C616 diff_1868170_2465070# gnd! 76.4fF
C617 diff_1588770_2136140# gnd! 33.7fF
C618 diff_1539240_2132330# gnd! 37.1fF
C619 diff_1577340_2164080# gnd! 79.2fF
C620 diff_1249680_1831340# gnd! 33.9fF
C621 diff_1297940_1835150# gnd! 34.5fF
C622 diff_1286510_1864360# gnd! 79.6fF
C623 diff_1007110_1640840# gnd! 35.0fF
C624 diff_958850_1642110# gnd! 34.9fF
C625 diff_995680_1626870# gnd! 80.2fF
C626 diff_932180_1625600# gnd! 77.2fF
C627 diff_1078230_1715770# gnd! 79.5fF
C628 diff_1151890_1790700# gnd! 35.3fF
C629 diff_1141730_1775460# gnd! 77.1fF
C630 diff_1076960_1775460# gnd! 78.6fF
C631 diff_1103630_1795780# gnd! 35.3fF
C632 diff_1223010_1865630# gnd! 77.2fF
C633 diff_1151890_1835150# gnd! 34.7fF
C634 diff_1103630_1831340# gnd! 34.5fF
C635 diff_1141730_1864360# gnd! 78.9fF
C636 diff_1297940_1941830# gnd! 33.7fF
C637 diff_1223010_1925320# gnd! 77.5fF
C638 diff_1249680_1944370# gnd! 33.9fF
C639 diff_1286510_1925320# gnd! 79.8fF
C640 diff_1367790_2015490# gnd! 80.4fF
C641 diff_1297940_1985010# gnd! 34.8fF
C642 diff_1249680_1981200# gnd! 35.2fF
C643 diff_1286510_2014220# gnd! 80.1fF
C644 diff_1442720_2091690# gnd! 34.4fF
C645 diff_1432560_2076450# gnd! 78.8fF
C646 diff_1367790_2076450# gnd! 79.0fF
C647 diff_1394460_2096770# gnd! 34.6fF
C648 diff_1513840_2167890# gnd! 76.9fF
C649 diff_1442720_2136140# gnd! 33.9fF
C650 diff_1394460_2132330# gnd! 34.5fF
C651 diff_1432560_2164080# gnd! 77.8fF
C652 diff_1588770_2242820# gnd! 33.7fF
C653 diff_1577340_2226310# gnd! 79.6fF
C654 diff_1539240_2247900# gnd! 36.9fF
C655 diff_1513840_2227580# gnd! 77.6fF
C656 diff_1658620_2316480# gnd! 78.6fF
C657 diff_1733550_2391410# gnd! 34.5fF
C658 diff_1723390_2376170# gnd! 76.6fF
C659 diff_1658620_2376170# gnd! 78.4fF
C660 diff_1685290_2396490# gnd! 34.2fF
C661 diff_1804670_2466340# gnd! 73.7fF
C662 diff_1879600_2541270# gnd! 34.4fF
C663 diff_1868170_2527300# gnd! 78.0fF
C664 diff_1804670_2526030# gnd! 76.4fF
C665 diff_1830070_2547620# gnd! 37.3fF
C666 diff_1949450_2616200# gnd! 75.6fF
C667 diff_2025650_2691130# gnd! 34.6fF
C668 diff_2014220_2677160# gnd! 76.4fF
C669 diff_1950720_2675890# gnd! 76.0fF
C670 diff_1976120_2696210# gnd! 37.8fF
C671 diff_2087880_1543050# gnd! 516.9fF
C672 diff_2025650_2735580# gnd! 34.5fF
C673 diff_1976120_2731770# gnd! 37.5fF
C674 diff_2057400_1583690# gnd! 512.8fF
C675 diff_2095500_2767330# gnd! 75.8fF
C676 diff_2014220_2764790# gnd! 75.5fF
C677 diff_2019300_1526540# gnd! 551.7fF
C678 diff_1879600_2585720# gnd! 34.1fF
C679 diff_1830070_2581910# gnd! 37.2fF
C680 diff_1868170_2614930# gnd! 76.5fF
C681 diff_1733550_2435860# gnd! 34.1fF
C682 diff_1685290_2432050# gnd! 33.9fF
C683 diff_1723390_2463800# gnd! 74.6fF
C684 diff_1539240_2282190# gnd! 37.1fF
C685 diff_1588770_2286000# gnd! 34.2fF
C686 diff_1577340_2315210# gnd! 77.0fF
C687 diff_1007110_1685290# gnd! 33.9fF
C688 diff_958850_1681480# gnd! 33.9fF
C689 diff_995680_1714500# gnd! 80.0fF
C690 diff_515620_1610360# gnd! 152.4fF
C691 diff_535940_1631950# gnd! 272.8fF
C692 diff_703580_1633220# gnd! 1554.3fF
C693 diff_862330_1642110# gnd! 33.9fF
C694 diff_850900_1626870# gnd! 80.8fF
C695 diff_932180_1715770# gnd! 77.1fF
C696 diff_1007110_1790700# gnd! 35.1fF
C697 diff_995680_1775460# gnd! 77.6fF
C698 diff_932180_1775460# gnd! 75.4fF
C699 diff_958850_1791970# gnd! 34.3fF
C700 diff_1076960_1866900# gnd! 80.7fF
C701 diff_1151890_1941830# gnd! 34.1fF
C702 diff_1141730_1925320# gnd! 77.9fF
C703 diff_1076960_1926590# gnd! 78.7fF
C704 diff_1103630_1945640# gnd! 34.1fF
C705 diff_1223010_2015490# gnd! 75.4fF
C706 diff_1151890_1985010# gnd! 35.6fF
C707 diff_1103630_1981200# gnd! 35.3fF
C708 diff_1141730_2014220# gnd! 77.4fF
C709 diff_1297940_2091690# gnd! 34.3fF
C710 diff_1286510_2076450# gnd! 79.0fF
C711 diff_1249680_2095500# gnd! 33.9fF
C712 diff_1223010_2076450# gnd! 77.2fF
C713 diff_1367790_2166620# gnd! 77.7fF
C714 diff_1442720_2242820# gnd! 33.9fF
C715 diff_1432560_2226310# gnd! 77.6fF
C716 diff_1367790_2227580# gnd! 77.8fF
C717 diff_1394460_2246630# gnd! 33.9fF
C718 diff_1513840_2316480# gnd! 75.5fF
C719 diff_1442720_2286000# gnd! 33.7fF
C720 diff_1394460_2282190# gnd! 34.2fF
C721 diff_1432560_2315210# gnd! 76.5fF
C722 diff_1588770_2391410# gnd! 34.0fF
C723 diff_1577340_2377440# gnd! 77.7fF
C724 diff_1539240_2396490# gnd! 37.1fF
C725 diff_1513840_2376170# gnd! 76.2fF
C726 diff_1658620_2466340# gnd! 76.9fF
C727 diff_1733550_2541270# gnd! 34.2fF
C728 diff_1723390_2526030# gnd! 75.7fF
C729 diff_1658620_2526030# gnd! 76.5fF
C730 diff_1685290_2546350# gnd! 34.6fF
C731 diff_1804670_2616200# gnd! 74.6fF
C732 diff_1879600_2691130# gnd! 34.5fF
C733 diff_1868170_2677160# gnd! 76.8fF
C734 diff_1804670_2675890# gnd! 75.7fF
C735 diff_1830070_2696210# gnd! 37.8fF
C736 diff_1941830_1543050# gnd! 560.1fF
C737 diff_1911350_1583690# gnd! 510.5fF
C738 diff_1873250_1527810# gnd! 551.7fF
C739 diff_1879600_2735580# gnd! 34.5fF
C740 diff_1830070_2739390# gnd! 36.4fF
C741 diff_1964690_1543050# gnd! 553.3fF
C742 diff_1949450_2774950# gnd! 74.6fF
C743 diff_1868170_2764790# gnd! 75.7fF
C744 diff_2002790_702310# gnd! 1366.0fF
C745 diff_1733550_2585720# gnd! 34.1fF
C746 diff_1685290_2581910# gnd! 34.1fF
C747 diff_1723390_2614930# gnd! 75.0fF
C748 diff_1588770_2435860# gnd! 34.1fF
C749 diff_1539240_2432050# gnd! 36.9fF
C750 diff_1577340_2465070# gnd! 78.1fF
C751 diff_1249680_2132330# gnd! 33.8fF
C752 diff_1297940_2136140# gnd! 34.3fF
C753 diff_1286510_2164080# gnd! 79.8fF
C754 diff_1007110_1835150# gnd! 35.1fF
C755 diff_958850_1831340# gnd! 34.2fF
C756 diff_995680_1864360# gnd! 79.8fF
C757 diff_861060_1690370# gnd! 34.6fF
C758 diff_580390_1633220# gnd! 841.9fF
C759 diff_601980_1651000# gnd! 219.7fF
C760 diff_850900_1714500# gnd! 80.1fF
C761 diff_703580_1714500# gnd! 1559.5fF
C762 diff_601980_1692910# gnd! 214.2fF
C763 diff_580390_1704340# gnd! 975.8fF
C764 diff_466090_1689100# gnd! 75.3fF
C765 diff_535940_1713230# gnd! 267.5fF
C766 diff_515620_1737360# gnd! 155.1fF
C767 diff_171450_1609090# gnd! 128.4fF
C768 diff_171450_1715770# gnd! 127.0fF
C769 diff_535940_1781810# gnd! 265.0fF
C770 diff_703580_1781810# gnd! 1414.0fF
C771 diff_861060_1790700# gnd! 38.1fF
C772 diff_850900_1775460# gnd! 77.2fF
C773 diff_932180_1865630# gnd! 77.1fF
C774 diff_1007110_1941830# gnd! 34.1fF
C775 diff_995680_1925320# gnd! 79.3fF
C776 diff_932180_1926590# gnd! 77.2fF
C777 diff_958850_1943100# gnd! 33.7fF
C778 diff_1076960_2016760# gnd! 77.6fF
C779 diff_1151890_2091690# gnd! 35.5fF
C780 diff_1141730_2075180# gnd! 79.4fF
C781 diff_1076960_2076450# gnd! 79.8fF
C782 diff_1103630_2096770# gnd! 35.1fF
C783 diff_1223010_2167890# gnd! 75.8fF
C784 diff_1151890_2136140# gnd! 33.9fF
C785 diff_1103630_2132330# gnd! 34.5fF
C786 diff_1141730_2164080# gnd! 77.7fF
C787 diff_1297940_2242820# gnd! 33.7fF
C788 diff_1286510_2226310# gnd! 78.8fF
C789 diff_1223010_2226310# gnd! 76.1fF
C790 diff_1249680_2244090# gnd! 33.7fF
C791 diff_1367790_2316480# gnd! 76.7fF
C792 diff_1442720_2391410# gnd! 34.1fF
C793 diff_1432560_2376170# gnd! 78.4fF
C794 diff_1394460_2396490# gnd! 34.4fF
C795 diff_1367790_2376170# gnd! 77.5fF
C796 diff_1513840_2466340# gnd! 75.8fF
C797 diff_1587500_2561590# gnd! 34.3fF
C798 diff_1577340_2526030# gnd! 76.9fF
C799 diff_1539240_2546350# gnd! 36.9fF
C800 diff_1513840_2526030# gnd! 75.3fF
C801 diff_1658620_2616200# gnd! 74.9fF
C802 diff_1733550_2691130# gnd! 34.5fF
C803 diff_1723390_2675890# gnd! 75.0fF
C804 diff_1658620_2675890# gnd! 76.8fF
C805 diff_1685290_2696210# gnd! 33.9fF
C806 diff_1819910_1543050# gnd! 595.3fF
C807 diff_1795780_1543050# gnd! 510.8fF
C808 diff_1765300_1584960# gnd! 511.0fF
C809 diff_1733550_2735580# gnd! 34.1fF
C810 diff_1685290_2731770# gnd! 33.9fF
C811 diff_1728470_1526540# gnd! 564.7fF
C812 diff_1804670_2766060# gnd! 74.0fF
C813 diff_1723390_2763520# gnd! 74.8fF
C814 diff_1673860_1543050# gnd! 549.5fF
C815 diff_1588770_2585720# gnd! 33.9fF
C816 diff_1539240_2581910# gnd! 36.9fF
C817 diff_1577340_2614930# gnd! 76.0fF
C818 diff_1442720_2435860# gnd! 33.7fF
C819 diff_1394460_2432050# gnd! 34.5fF
C820 diff_1432560_2463800# gnd! 76.9fF
C821 diff_1442720_2541270# gnd! 34.5fF
C822 diff_1432560_2526030# gnd! 76.7fF
C823 diff_1249680_2282190# gnd! 33.9fF
C824 diff_1297940_2286000# gnd! 34.2fF
C825 diff_1286510_2315210# gnd! 78.2fF
C826 diff_1007110_1985010# gnd! 34.8fF
C827 diff_958850_1981200# gnd! 35.2fF
C828 diff_995680_2014220# gnd! 78.7fF
C829 diff_861060_1835150# gnd! 38.4fF
C830 diff_850900_1863090# gnd! 78.9fF
C831 diff_580390_1783080# gnd! 959.1fF
C832 diff_601980_1800860# gnd! 210.6fF
C833 diff_448310_1662430# gnd! 321.4fF
C834 diff_515620_1789430# gnd! 173.4fF
C835 diff_703580_1863090# gnd! 1586.1fF
C836 diff_601980_1842770# gnd! 212.5fF
C837 diff_580390_1854200# gnd! 958.0fF
C838 diff_462280_1706880# gnd! 483.2fF
C839 diff_93980_1783080# gnd! 279.6fF
C840 diff_535940_1849120# gnd! 274.9fF
C841 diff_515620_1841500# gnd! 179.7fF
C842 diff_515620_1906270# gnd! 161.6fF
C843 diff_535940_1931670# gnd! 268.5fF
C844 diff_861060_1941830# gnd! 37.1fF
C845 diff_850900_1925320# gnd! 78.7fF
C846 diff_703580_1931670# gnd! 1568.2fF
C847 diff_580390_1932940# gnd! 1213.2fF
C848 diff_601980_1950720# gnd! 224.1fF
C849 diff_932180_2015490# gnd! 75.8fF
C850 diff_995680_2076450# gnd! 79.6fF
C851 diff_1007110_2091690# gnd! 35.0fF
C852 diff_932180_2076450# gnd! 76.9fF
C853 diff_958850_2092960# gnd! 34.8fF
C854 diff_1076960_2167890# gnd! 77.7fF
C855 diff_1151890_2242820# gnd! 33.9fF
C856 diff_1141730_2226310# gnd! 77.6fF
C857 diff_1076960_2226310# gnd! 78.5fF
C858 diff_1103630_2246630# gnd! 33.8fF
C859 diff_1223010_2316480# gnd! 73.9fF
C860 diff_1297940_2391410# gnd! 34.0fF
C861 diff_1286510_2377440# gnd! 78.9fF
C862 diff_1223010_2376170# gnd! 77.0fF
C863 diff_1248410_2400300# gnd! 36.8fF
C864 diff_1367790_2466340# gnd! 76.3fF
C865 diff_1367790_2526030# gnd! 76.5fF
C866 diff_1394460_2546350# gnd! 34.9fF
C867 diff_1513840_2616200# gnd! 75.2fF
C868 diff_1588770_2691130# gnd! 33.9fF
C869 diff_1539240_2696210# gnd! 37.1fF
C870 diff_1513840_2675890# gnd! 75.8fF
C871 diff_1577340_2675890# gnd! 76.3fF
C872 diff_1649730_1543050# gnd! 512.7fF
C873 diff_1620520_1543050# gnd! 539.0fF
C874 diff_1582420_1527810# gnd! 550.0fF
C875 diff_1588770_2735580# gnd! 33.9fF
C876 diff_1539240_2731770# gnd! 37.4fF
C877 diff_1658620_2766060# gnd! 76.2fF
C878 diff_1577340_2764790# gnd! 76.7fF
C879 diff_1442720_2585720# gnd! 33.9fF
C880 diff_1394460_2581910# gnd! 34.1fF
C881 diff_1432560_2613660# gnd! 76.7fF
C882 diff_1297940_2435860# gnd! 33.9fF
C883 diff_1248410_2432050# gnd! 37.9fF
C884 diff_1286510_2465070# gnd! 78.2fF
C885 diff_1151890_2286000# gnd! 33.7fF
C886 diff_1103630_2282190# gnd! 33.9fF
C887 diff_1141730_2315210# gnd! 79.1fF
C888 diff_1007110_2136140# gnd! 34.5fF
C889 diff_958850_2132330# gnd! 34.1fF
C890 diff_995680_2164080# gnd! 77.5fF
C891 diff_861060_1986280# gnd! 37.1fF
C892 diff_850900_2014220# gnd! 76.9fF
C893 diff_703580_2012950# gnd! 1425.3fF
C894 diff_601980_1992630# gnd! 226.1fF
C895 diff_466090_1988820# gnd! 74.3fF
C896 diff_580390_2004060# gnd! 1009.0fF
C897 diff_535940_2012950# gnd! 267.2fF
C898 diff_515620_2037080# gnd! 162.8fF
C899 diff_73660_2023110# gnd! 1005.8fF
C900 d3 gnd! 2946.4fF
C901 diff_72390_1687830# gnd! 931.0fF
C902 diff_535940_2082800# gnd! 263.4fF
C903 diff_703580_2081530# gnd! 1535.4fF
C904 diff_861060_2091690# gnd! 38.5fF
C905 diff_850900_2076450# gnd! 77.5fF
C906 diff_580390_2082800# gnd! 1101.9fF
C907 diff_601980_2100580# gnd! 212.6fF
C908 diff_932180_2166620# gnd! 75.8fF
C909 diff_1007110_2242820# gnd! 34.1fF
C910 diff_995680_2226310# gnd! 80.2fF
C911 diff_932180_2227580# gnd! 76.2fF
C912 diff_957580_2263140# gnd! 35.2fF
C913 diff_1076960_2316480# gnd! 78.7fF
C914 diff_1151890_2391410# gnd! 35.1fF
C915 diff_1141730_2376170# gnd! 79.4fF
C916 diff_1076960_2376170# gnd! 80.2fF
C917 diff_1103630_2395220# gnd! 34.7fF
C918 diff_1223010_2466340# gnd! 75.8fF
C919 diff_1151890_2434590# gnd! 34.5fF
C920 diff_1103630_2432050# gnd! 34.5fF
C921 diff_1141730_2463800# gnd! 77.4fF
C922 diff_1297940_2541270# gnd! 34.6fF
C923 diff_1286510_2526030# gnd! 77.9fF
C924 diff_1248410_2546350# gnd! 37.6fF
C925 diff_1223010_2526030# gnd! 75.5fF
C926 diff_1367790_2616200# gnd! 76.3fF
C927 diff_1442720_2691130# gnd! 33.9fF
C928 diff_1432560_2675890# gnd! 76.5fF
C929 diff_1367790_2675890# gnd! 76.0fF
C930 diff_1394460_2696210# gnd! 34.5fF
C931 diff_1527810_1543050# gnd! 554.5fF
C932 diff_1513840_2766060# gnd! 75.5fF
C933 diff_1504950_1543050# gnd! 541.3fF
C934 diff_1442720_2735580# gnd! 33.9fF
C935 diff_1394460_2731770# gnd! 34.5fF
C936 diff_1474470_1583690# gnd! 511.0fF
C937 diff_1432560_2763520# gnd! 76.2fF
C938 diff_1436370_1529080# gnd! 592.0fF
C939 diff_1297940_2585720# gnd! 33.9fF
C940 diff_1248410_2581910# gnd! 37.2fF
C941 diff_1286510_2614930# gnd! 76.4fF
C942 diff_1007110_2286000# gnd! 34.2fF
C943 diff_957580_2282190# gnd! 35.4fF
C944 diff_861060_2136140# gnd! 37.8fF
C945 diff_850900_2164080# gnd! 78.0fF
C946 diff_515620_2090420# gnd! 172.4fF
C947 diff_448310_1962150# gnd! 320.4fF
C948 diff_703580_2164080# gnd! 1566.2fF
C949 diff_601980_2143760# gnd! 214.7fF
C950 diff_580390_2155190# gnd! 1083.7fF
C951 diff_535940_2156460# gnd! 268.7fF
C952 diff_350520_1598930# gnd! 733.5fF
C953 diff_515620_2147570# gnd! 172.8fF
C954 diff_515620_2207260# gnd! 159.6fF
C955 diff_535940_2232660# gnd! 268.4fF
C956 diff_703580_2232660# gnd! 1606.5fF
C957 diff_861060_2242820# gnd! 37.1fF
C958 diff_850900_2226310# gnd! 78.3fF
C959 diff_861060_2286000# gnd! 37.1fF
C960 diff_580390_2232660# gnd! 953.2fF
C961 diff_601980_2251710# gnd! 216.9fF
C962 diff_995680_2315210# gnd! 79.7fF
C963 diff_932180_2316480# gnd! 75.7fF
C964 diff_850900_2315210# gnd! 76.6fF
C965 diff_1007110_2391410# gnd! 34.8fF
C966 diff_995680_2377440# gnd! 80.3fF
C967 diff_932180_2376170# gnd! 76.9fF
C968 diff_957580_2396490# gnd! 37.4fF
C969 diff_1076960_2466340# gnd! 76.5fF
C970 diff_1076960_2526030# gnd! 76.0fF
C971 diff_1151890_2541270# gnd! 35.1fF
C972 diff_1141730_2526030# gnd! 77.1fF
C973 diff_1103630_2545080# gnd! 35.1fF
C974 diff_1223010_2616200# gnd! 74.6fF
C975 diff_1223010_2675890# gnd! 74.8fF
C976 diff_1248410_2696210# gnd! 37.6fF
C977 diff_1297940_2691130# gnd! 34.5fF
C978 diff_1286510_2675890# gnd! 76.8fF
C979 diff_1358900_1543050# gnd! 512.7fF
C980 diff_1329690_1543050# gnd! 554.9fF
C981 diff_1291590_1526540# gnd! 549.7fF
C982 diff_1248410_2731770# gnd! 37.6fF
C983 diff_1297940_2735580# gnd! 34.5fF
C984 diff_1383030_1543050# gnd! 550.0fF
C985 diff_1367790_2766060# gnd! 74.4fF
C986 diff_1286510_2763520# gnd! 77.4fF
C987 diff_1236980_1543050# gnd! 601.8fF
C988 diff_1151890_2585720# gnd! 33.9fF
C989 diff_1103630_2581910# gnd! 34.1fF
C990 diff_1141730_2613660# gnd! 76.9fF
C991 diff_1007110_2435860# gnd! 34.1fF
C992 diff_957580_2432050# gnd! 37.8fF
C993 diff_995680_2465070# gnd! 78.4fF
C994 diff_703580_2313940# gnd! 1582.0fF
C995 diff_180340_2162810# gnd! 276.8fF
C996 diff_172720_2129790# gnd! 273.5fF
C997 diff_601980_2293620# gnd! 224.4fF
C998 diff_580390_2305050# gnd! 825.5fF
C999 diff_466090_2289810# gnd! 72.3fF
C1000 diff_535940_2313940# gnd! 268.3fF
C1001 diff_515620_2338070# gnd! 158.9fF
C1002 diff_535940_2382520# gnd! 263.9fF
C1003 diff_703580_2382520# gnd! 1429.4fF
C1004 diff_861060_2391410# gnd! 35.0fF
C1005 diff_850900_2376170# gnd! 77.3fF
C1006 diff_861060_2435860# gnd! 33.7fF
C1007 diff_932180_2466340# gnd! 76.0fF
C1008 diff_850900_2463800# gnd! 77.1fF
C1009 diff_1005840_2548890# gnd! 37.3fF
C1010 diff_995680_2526030# gnd! 78.3fF
C1011 diff_932180_2526030# gnd! 76.3fF
C1012 diff_957580_2546350# gnd! 38.3fF
C1013 diff_1076960_2616200# gnd! 76.4fF
C1014 diff_1151890_2691130# gnd! 34.2fF
C1015 diff_1140460_2679700# gnd! 77.2fF
C1016 diff_1076960_2675890# gnd! 76.6fF
C1017 diff_1103630_2694940# gnd! 34.5fF
C1018 diff_1151890_2735580# gnd! 34.2fF
C1019 diff_1214120_1543050# gnd! 529.3fF
C1020 diff_1183640_1584960# gnd! 513.8fF
C1021 diff_1145540_1527810# gnd! 621.8fF
C1022 diff_1223010_2766060# gnd! 74.9fF
C1023 diff_1141730_2763520# gnd! 76.4fF
C1024 diff_1103630_2731770# gnd! 34.5fF
C1025 diff_1005840_2585720# gnd! 36.9fF
C1026 diff_957580_2581910# gnd! 37.4fF
C1027 diff_995680_2614930# gnd! 75.3fF
C1028 diff_580390_2383790# gnd! 1078.6fF
C1029 diff_600710_2406650# gnd! 214.6fF
C1030 diff_515620_2390140# gnd! 172.6fF
C1031 diff_448310_2263140# gnd! 314.1fF
C1032 diff_703580_2463800# gnd! 1466.0fF
C1033 diff_600710_2443480# gnd! 213.0fF
C1034 diff_580390_2454910# gnd! 947.4fF
C1035 diff_535940_2456180# gnd! 267.8fF
C1036 diff_171450_2419350# gnd! 128.3fF
C1037 diff_346710_1485900# gnd! 567.7fF
C1038 diff_515620_2447290# gnd! 175.6fF
C1039 diff_515620_2506980# gnd! 156.8fF
C1040 diff_245110_1436370# gnd! 2580.7fF
C1041 diff_535940_2532380# gnd! 270.0fF
C1042 diff_703580_2532380# gnd! 1429.9fF
C1043 diff_861060_2541270# gnd! 35.4fF
C1044 diff_850900_2526030# gnd! 77.7fF
C1045 diff_932180_2616200# gnd! 75.4fF
C1046 diff_861060_2585720# gnd! 33.6fF
C1047 diff_580390_2532380# gnd! 949.3fF
C1048 diff_600710_2551430# gnd! 220.9fF
C1049 diff_850900_2613660# gnd! 75.3fF
C1050 diff_1005840_2715260# gnd! 35.4fF
C1051 diff_995680_2675890# gnd! 79.4fF
C1052 diff_957580_2696210# gnd! 38.1fF
C1053 diff_932180_2675890# gnd! 74.8fF
C1054 diff_1068070_1543050# gnd! 521.0fF
C1055 diff_1038860_1543050# gnd! 544.7fF
C1056 diff_1000760_1526540# gnd! 550.8fF
C1057 diff_1007110_2735580# gnd! 34.5fF
C1058 diff_957580_2731770# gnd! 37.8fF
C1059 diff_1092200_1543050# gnd! 549.2fF
C1060 diff_1076960_2766060# gnd! 75.5fF
C1061 diff_995680_2763520# gnd! 78.2fF
C1062 diff_946150_1543050# gnd! 588.6fF
C1063 diff_171450_2527300# gnd! 125.6fF
C1064 diff_702310_2614930# gnd! 1483.8fF
C1065 diff_600710_2593340# gnd! 220.9fF
C1066 diff_580390_2603500# gnd! 945.7fF
C1067 diff_466090_2589530# gnd! 77.8fF
C1068 diff_535940_2611120# gnd! 272.3fF
C1069 diff_515620_2636520# gnd! 158.2fF
C1070 diff_92710_2637790# gnd! 274.9fF
C1071 diff_535940_2680970# gnd! 275.7fF
C1072 diff_703580_2682240# gnd! 1409.3fF
C1073 diff_861060_2691130# gnd! 34.8fF
C1074 diff_850900_2675890# gnd! 76.7fF
C1075 diff_861060_2735580# gnd! 34.4fF
C1076 diff_923290_1543050# gnd! 514.4fF
C1077 diff_892810_1584960# gnd! 552.1fF
C1078 diff_854710_1527810# gnd! 576.4fF
C1079 diff_932180_2766060# gnd! 75.7fF
C1080 diff_850900_2763520# gnd! 76.2fF
C1081 diff_580390_2682240# gnd! 995.6fF
C1082 diff_600710_2702560# gnd! 219.5fF
C1083 diff_515620_2703830# gnd! 176.1fF
C1084 diff_243840_2250440# gnd! 2418.7fF
C1085 diff_448310_2561590# gnd! 313.5fF
C1086 diff_702310_2763520# gnd! 1568.2fF
C1087 diff_600710_2741930# gnd! 217.3fF
C1088 diff_450850_1684020# gnd! 1146.9fF
C1089 diff_580390_2753360# gnd! 914.4fF
C1090 diff_535940_2755900# gnd! 278.9fF
C1091 diff_515620_2754630# gnd! 159.7fF
C1092 diff_553720_1553210# gnd! 824.8fF
C1093 diff_345440_2600960# gnd! 556.4fF
C1094 diff_2461260_2799080# gnd! 44.6fF
C1095 diff_2565400_2871470# gnd! 79.4fF
C1096 diff_2482850_2806700# gnd! 333.9fF
C1097 diff_2597150_2896870# gnd! 89.2fF
C1098 clk2 gnd! 2997.2fF
C1099 diff_2227580_2936240# gnd! 40.6fF
C1100 diff_73660_2682240# gnd! 1008.3fF
C1101 d2 gnd! 3102.4fF
C1102 diff_72390_2499360# gnd! 928.3fF
C1103 o1 gnd! 811.5fF
C1104 diff_2512060_2913380# gnd! 263.0fF
C1105 diff_2556510_3018790# gnd! 452.3fF
C1106 diff_2195830_2933700# gnd! 1224.5fF
C1107 diff_234950_1145540# gnd! 684.0fF
C1108 diff_369570_1160780# gnd! 2441.7fF
C1109 diff_2170430_3058160# gnd! 73.8fF
C1110 diff_2133600_3073400# gnd! 78.0fF
C1111 diff_2035810_3031490# gnd! 243.3fF
C1112 diff_2198370_3069590# gnd! 615.5fF
C1113 o0 gnd! 617.7fF
C1114 diff_1437640_3022600# gnd! 126.9fF
C1115 diff_1334770_3023870# gnd! 130.1fF
C1116 diff_1068070_2976880# gnd! 272.8fF
C1117 diff_998220_3009900# gnd! 287.3fF
C1118 diff_1512570_3046730# gnd! 251.7fF
C1119 diff_1336040_3056890# gnd! 1015.2fF
C1120 diff_1408430_3068320# gnd! 910.8fF
C1121 diff_266700_2927350# gnd! 2579.0fF
C1122 diff_408940_3023870# gnd! 129.9fF
C1123 Vdd gnd! 41631.7fF
C1124 diff_139700_2962910# gnd! 1205.1fF
C1125 diff_175260_2987040# gnd! 272.2fF
C1126 diff_102870_3011170# gnd! 291.6fF
C1127 diff_306070_3023870# gnd! 133.0fF
C1128 diff_483870_3046730# gnd! 272.2fF
C1129 diff_92710_2421890# gnd! 1698.0fF
C1130 diff_306070_3053080# gnd! 1013.3fF
C1131 diff_379730_3067050# gnd! 925.3fF
C1132 diff_2028190_3027680# gnd! 459.6fF
C1133 d0 gnd! 3008.2fF
C1134 d1 gnd! 2989.3fF
C1135 diff_2134870_3131820# gnd! 321.3fF
