* SPICE3 file created from 4001.ext - technology: nmos

.option scale=0.001u

M1000 clk2 GND GND GND efet w=97200 l=7200
+ ad=-1.68369e+09 pd=1.548e+06 as=-1.10908e+09 ps=3.9312e+07 
M1001 clk1 GND GND GND efet w=97200 l=7200
+ ad=4.19593e+08 pd=1.1832e+06 as=0 ps=0 
M1002 d2 GND d2 GND efet w=177000 l=112200
+ ad=2.07814e+09 pd=2.9952e+06 as=0 ps=0 
M1003 d3 GND d3 GND efet w=178800 l=115200
+ ad=1.99373e+09 pd=4.0992e+06 as=0 ps=0 
M1004 sync GND GND GND efet w=91200 l=7200
+ ad=1.84431e+09 pd=2.6184e+06 as=0 ps=0 
M1005 GND diff_338400_1662000# d3 GND efet w=933600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M1006 GND diff_494400_1662000# d2 GND efet w=932400 l=3600
+ ad=0 pd=0 as=0 ps=0 
M1007 Vdd diff_355200_1366800# d3 GND efet w=431400 l=10200
+ ad=8.29643e+08 pd=1.52592e+07 as=0 ps=0 
M1008 GND diff_649200_1662000# d1 GND efet w=932400 l=3600
+ ad=0 pd=0 as=1.99318e+09 ps=3.036e+06 
M1009 GND diff_804000_1662000# d0 GND efet w=932400 l=3600
+ ad=0 pd=0 as=1.8535e+09 ps=3.0168e+06 
M1010 GND diff_2433600_1742400# diff_2437200_1698000# GND efet w=356400 l=6000
+ ad=0 pd=0 as=7.02385e+08 ps=1.476e+06 
M1011 GND clk1 diff_2613600_1719600# GND efet w=25200 l=7200
+ ad=0 pd=0 as=4.4784e+08 ps=91200 
M1012 GND sync diff_2433600_1742400# GND efet w=76800 l=7200
+ ad=0 pd=0 as=-1.35449e+09 ps=607200 
M1013 diff_2802000_1732800# diff_2751600_1686000# GND GND efet w=27600 l=6000
+ ad=5.2992e+08 pd=182400 as=0 ps=0 
M1014 diff_2649600_1428000# diff_2802000_1732800# GND GND efet w=40800 l=6000
+ ad=7.632e+08 pd=204000 as=0 ps=0 
M1015 GND diff_2433600_1742400# diff_2743200_1714800# GND efet w=40800 l=6000
+ ad=0 pd=0 as=3.9168e+08 ps=100800 
M1016 diff_2613600_1719600# Vdd Vdd GND efet w=7200 l=9600
+ ad=0 pd=0 as=0 ps=0 
M1017 diff_2433600_1742400# diff_2664000_1686000# GND GND efet w=46800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1018 GND diff_1003200_1702800# diff_1008000_1686000# GND efet w=619200 l=7200
+ ad=0 pd=0 as=-2.06364e+09 ps=2.7792e+06 
M1019 Vdd diff_1657200_1702800# diff_1008000_1686000# GND efet w=643200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1020 diff_1008000_1686000# diff_1004400_1680000# diff_1008000_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1021 diff_1008000_1686000# diff_1004400_1680000# diff_1028400_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1022 diff_1008000_1686000# diff_1004400_1680000# diff_1048800_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1023 diff_1008000_1686000# diff_1004400_1680000# diff_1069200_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1024 diff_1008000_1686000# diff_1004400_1680000# diff_1089600_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1025 diff_1008000_1686000# diff_1004400_1680000# diff_1110000_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1026 diff_1008000_1686000# diff_1004400_1680000# diff_1130400_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1027 diff_1008000_1686000# diff_1004400_1680000# diff_1150800_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1028 diff_1008000_1686000# diff_1004400_1680000# diff_1171200_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1029 diff_1008000_1686000# diff_1004400_1680000# diff_1191600_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1030 diff_1008000_1686000# diff_1004400_1680000# diff_1212000_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1031 diff_1008000_1686000# diff_1004400_1680000# diff_1232400_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1032 diff_1008000_1686000# diff_1004400_1680000# diff_1252800_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1033 diff_1008000_1686000# diff_1004400_1680000# diff_1273200_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1034 diff_1008000_1686000# diff_1004400_1680000# diff_1293600_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1035 diff_1008000_1686000# diff_1004400_1680000# diff_1314000_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1036 diff_1008000_1686000# diff_1004400_1680000# diff_1334400_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1037 diff_1008000_1686000# diff_1004400_1680000# diff_1354800_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1038 diff_1008000_1686000# diff_1004400_1680000# diff_1375200_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1039 diff_1008000_1686000# diff_1004400_1680000# diff_1395600_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1040 diff_1008000_1686000# diff_1004400_1680000# diff_1416000_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1041 diff_1008000_1686000# diff_1004400_1680000# diff_1436400_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1042 diff_1008000_1686000# diff_1004400_1680000# diff_1456800_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1043 diff_1008000_1686000# diff_1004400_1680000# diff_1477200_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1044 diff_1008000_1686000# diff_1004400_1680000# diff_1497600_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1045 diff_1008000_1686000# diff_1004400_1680000# diff_1518000_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1046 diff_1008000_1686000# diff_1004400_1680000# diff_1538400_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1047 diff_1008000_1686000# diff_1004400_1680000# diff_1558800_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1048 diff_1008000_1686000# diff_1004400_1680000# diff_1579200_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1049 diff_1008000_1686000# diff_1004400_1680000# diff_1599600_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1050 diff_1008000_1686000# diff_1004400_1680000# diff_1620000_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1051 diff_1008000_1686000# diff_1004400_1680000# diff_1640400_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1052 diff_1008000_1686000# diff_1004400_1680000# diff_1660800_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1053 diff_1008000_1686000# diff_1004400_1680000# diff_1681200_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1054 diff_1008000_1686000# diff_1004400_1680000# diff_1701600_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1055 diff_1008000_1686000# diff_1004400_1680000# diff_1722000_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1056 diff_1008000_1686000# diff_1004400_1680000# diff_1742400_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1057 diff_1008000_1686000# diff_1004400_1680000# diff_1762800_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1058 diff_1008000_1686000# diff_1004400_1680000# diff_1783200_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1059 diff_1008000_1686000# diff_1004400_1680000# diff_1803600_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1060 diff_1008000_1686000# diff_1004400_1680000# diff_1824000_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1061 diff_1008000_1686000# diff_1004400_1680000# diff_1844400_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1062 diff_1008000_1686000# diff_1004400_1680000# diff_1864800_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1063 diff_1008000_1686000# diff_1004400_1680000# diff_1885200_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1064 diff_1008000_1686000# diff_1004400_1680000# diff_1905600_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1065 diff_1008000_1686000# diff_1004400_1680000# diff_1926000_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1066 diff_1008000_1686000# diff_1004400_1680000# diff_1946400_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1067 diff_1008000_1686000# diff_1004400_1680000# diff_1966800_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1068 diff_1008000_1686000# diff_1004400_1680000# diff_1987200_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1069 diff_1008000_1686000# diff_1004400_1680000# diff_2007600_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1070 diff_1008000_1686000# diff_1004400_1680000# diff_2028000_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1071 diff_1008000_1686000# diff_1004400_1680000# diff_2048400_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1072 diff_1008000_1686000# diff_1004400_1680000# diff_2068800_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1073 diff_1008000_1686000# diff_1004400_1680000# diff_2089200_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1074 diff_1008000_1686000# diff_1004400_1680000# diff_2109600_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1075 diff_1008000_1686000# diff_1004400_1680000# diff_2130000_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1076 diff_1008000_1686000# diff_1004400_1680000# diff_2150400_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1077 diff_1008000_1686000# diff_1004400_1680000# diff_2170800_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1078 diff_1008000_1686000# diff_1004400_1680000# diff_2191200_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1079 diff_1008000_1686000# diff_1004400_1680000# diff_2211600_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1080 diff_1008000_1686000# diff_1004400_1680000# diff_2232000_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1081 diff_1008000_1686000# diff_1004400_1680000# diff_2252400_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1082 diff_1008000_1686000# diff_1004400_1680000# diff_2272800_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1083 diff_1008000_1686000# diff_1004400_1680000# diff_2293200_1663200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1084 diff_2367600_1674000# diff_2361600_427200# diff_1004400_1680000# GND efet w=89400 l=7200
+ ad=-6.74807e+08 pd=688800 as=9.5616e+08 ps=230400 
M1085 Vdd Vdd diff_366000_1504800# GND efet w=9600 l=9600
+ ad=0 pd=0 as=2.4912e+08 ps=72000 
M1086 Vdd Vdd diff_428400_1507200# GND efet w=8400 l=10800
+ ad=0 pd=0 as=1.9872e+08 ps=67200 
M1087 diff_366000_1504800# diff_366000_1504800# diff_366000_1504800# GND efet w=1800 l=3600
+ ad=0 pd=0 as=0 ps=0 
M1088 Vdd diff_366000_1504800# diff_355200_1366800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=-1.26953e+09 ps=650400 
M1089 Vdd diff_428400_1507200# diff_338400_1662000# GND efet w=8400 l=7200
+ ad=0 pd=0 as=-5.99927e+08 ps=768000 
M1090 diff_428400_1507200# diff_428400_1507200# diff_428400_1507200# GND efet w=1800 l=4800
+ ad=0 pd=0 as=0 ps=0 
M1091 Vdd diff_510000_1366800# d2 GND efet w=429600 l=10800
+ ad=0 pd=0 as=0 ps=0 
M1092 diff_366000_1504800# diff_366000_1504800# diff_366000_1504800# GND efet w=1200 l=3600
+ ad=0 pd=0 as=0 ps=0 
M1093 diff_355200_1366800# diff_366000_1504800# diff_355200_1366800# GND efet w=42600 l=13800
+ ad=0 pd=0 as=0 ps=0 
M1094 diff_428400_1507200# diff_428400_1507200# diff_428400_1507200# GND efet w=1200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M1095 Vdd Vdd diff_520800_1503600# GND efet w=7200 l=9600
+ ad=0 pd=0 as=2.1312e+08 ps=74400 
M1096 Vdd Vdd diff_583200_1506000# GND efet w=9600 l=10800
+ ad=0 pd=0 as=2.2032e+08 ps=79200 
M1097 diff_520800_1503600# diff_520800_1503600# diff_520800_1503600# GND efet w=2400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M1098 Vdd diff_520800_1503600# diff_510000_1366800# GND efet w=8400 l=7200
+ ad=0 pd=0 as=-1.26809e+09 ps=650400 
M1099 Vdd diff_583200_1506000# diff_494400_1662000# GND efet w=8400 l=7200
+ ad=0 pd=0 as=-5.38007e+08 ps=770400 
M1100 diff_583200_1506000# diff_583200_1506000# diff_583200_1506000# GND efet w=3600 l=4200
+ ad=0 pd=0 as=0 ps=0 
M1101 diff_520800_1503600# diff_520800_1503600# diff_520800_1503600# GND efet w=1200 l=4800
+ ad=0 pd=0 as=0 ps=0 
M1102 diff_338400_1662000# diff_428400_1507200# diff_338400_1662000# GND efet w=57000 l=6600
+ ad=0 pd=0 as=0 ps=0 
M1103 diff_510000_1366800# diff_520800_1503600# diff_510000_1366800# GND efet w=43800 l=13800
+ ad=0 pd=0 as=0 ps=0 
M1104 diff_583200_1506000# diff_583200_1506000# diff_583200_1506000# GND efet w=1200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1105 Vdd diff_664800_1365600# d1 GND efet w=430800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1106 Vdd Vdd diff_673200_1506000# GND efet w=8400 l=10800
+ ad=0 pd=0 as=1.7712e+08 ps=64800 
M1107 Vdd Vdd diff_738000_1506000# GND efet w=8400 l=10800
+ ad=0 pd=0 as=1.9152e+08 ps=62400 
M1108 Vdd diff_820800_1365600# d0 GND efet w=428400 l=10200
+ ad=0 pd=0 as=0 ps=0 
M1109 Vdd diff_673200_1506000# diff_664800_1365600# GND efet w=7200 l=7200
+ ad=0 pd=0 as=-1.23929e+09 ps=696000 
M1110 diff_673200_1506000# diff_673200_1506000# diff_673200_1506000# GND efet w=2400 l=4800
+ ad=0 pd=0 as=0 ps=0 
M1111 diff_494400_1662000# diff_583200_1506000# diff_494400_1662000# GND efet w=57000 l=6600
+ ad=0 pd=0 as=0 ps=0 
M1112 Vdd diff_738000_1506000# diff_649200_1662000# GND efet w=7800 l=7800
+ ad=0 pd=0 as=-6.38807e+08 ps=765600 
M1113 diff_738000_1506000# diff_738000_1506000# diff_738000_1506000# GND efet w=1200 l=1800
+ ad=0 pd=0 as=0 ps=0 
M1114 diff_673200_1506000# diff_673200_1506000# diff_673200_1506000# GND efet w=1200 l=4800
+ ad=0 pd=0 as=0 ps=0 
M1115 diff_738000_1506000# diff_738000_1506000# diff_738000_1506000# GND efet w=600 l=1800
+ ad=0 pd=0 as=0 ps=0 
M1116 Vdd Vdd diff_831600_1504800# GND efet w=8400 l=9600
+ ad=0 pd=0 as=2.1744e+08 ps=67200 
M1117 Vdd Vdd diff_886800_1546800# GND efet w=8400 l=9600
+ ad=0 pd=0 as=1.7856e+08 ps=60000 
M1118 diff_831600_1504800# diff_831600_1504800# diff_831600_1504800# GND efet w=600 l=1800
+ ad=0 pd=0 as=0 ps=0 
M1119 Vdd diff_831600_1504800# diff_820800_1365600# GND efet w=7200 l=7200
+ ad=0 pd=0 as=-1.24937e+09 ps=648000 
M1120 Vdd diff_886800_1546800# diff_804000_1662000# GND efet w=7200 l=7200
+ ad=0 pd=0 as=-5.75447e+08 ps=748800 
M1121 diff_886800_1546800# diff_886800_1546800# diff_886800_1546800# GND efet w=1200 l=1800
+ ad=0 pd=0 as=0 ps=0 
M1122 diff_1008000_1663200# diff_1004400_1657200# diff_1008000_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1123 diff_1028400_1663200# diff_1004400_1657200# diff_1028400_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1124 diff_1048800_1663200# diff_1004400_1657200# diff_1048800_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1125 diff_1069200_1663200# diff_1004400_1657200# diff_1069200_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1126 diff_1089600_1663200# diff_1004400_1657200# diff_1089600_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1127 diff_1110000_1663200# diff_1004400_1657200# diff_1110000_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1128 diff_1130400_1663200# diff_1004400_1657200# diff_1130400_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1129 diff_1150800_1663200# diff_1004400_1657200# diff_1150800_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1130 diff_1171200_1663200# diff_1004400_1657200# diff_1171200_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1131 diff_1191600_1663200# diff_1004400_1657200# diff_1191600_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1132 diff_1212000_1663200# diff_1004400_1657200# diff_1212000_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1133 diff_1232400_1663200# diff_1004400_1657200# diff_1232400_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1134 diff_1252800_1663200# diff_1004400_1657200# diff_1252800_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1135 diff_1273200_1663200# diff_1004400_1657200# diff_1273200_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1136 diff_1293600_1663200# diff_1004400_1657200# diff_1293600_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1137 diff_1314000_1663200# diff_1004400_1657200# diff_1314000_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1138 diff_1334400_1663200# diff_1004400_1657200# diff_1334400_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1139 diff_1354800_1663200# diff_1004400_1657200# diff_1354800_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1140 diff_1375200_1663200# diff_1004400_1657200# diff_1375200_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1141 diff_1395600_1663200# diff_1004400_1657200# diff_1395600_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1142 diff_1416000_1663200# diff_1004400_1657200# diff_1416000_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1143 diff_1436400_1663200# diff_1004400_1657200# diff_1436400_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1144 diff_1456800_1663200# diff_1004400_1657200# diff_1456800_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1145 diff_1477200_1663200# diff_1004400_1657200# diff_1477200_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1146 diff_1497600_1663200# diff_1004400_1657200# diff_1497600_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1147 diff_1518000_1663200# diff_1004400_1657200# diff_1518000_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1148 diff_1538400_1663200# diff_1004400_1657200# diff_1538400_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1149 diff_1558800_1663200# diff_1004400_1657200# diff_1558800_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1150 diff_1579200_1663200# diff_1004400_1657200# diff_1579200_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1151 diff_1599600_1663200# diff_1004400_1657200# diff_1599600_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1152 diff_1620000_1663200# diff_1004400_1657200# diff_1620000_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1153 diff_1640400_1663200# diff_1004400_1657200# diff_1640400_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1154 diff_1660800_1663200# diff_1004400_1657200# diff_1660800_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1155 diff_1681200_1663200# diff_1004400_1657200# diff_1681200_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1156 diff_1701600_1663200# diff_1004400_1657200# diff_1701600_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1157 diff_1722000_1663200# diff_1004400_1657200# diff_1722000_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1158 diff_1742400_1663200# diff_1004400_1657200# diff_1742400_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1159 diff_1762800_1663200# diff_1004400_1657200# diff_1762800_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1160 diff_1783200_1663200# diff_1004400_1657200# diff_1783200_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1161 diff_1803600_1663200# diff_1004400_1657200# diff_1803600_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1162 diff_1824000_1663200# diff_1004400_1657200# diff_1824000_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1163 diff_1844400_1663200# diff_1004400_1657200# diff_1844400_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1164 diff_1864800_1663200# diff_1004400_1657200# diff_1864800_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1165 diff_1885200_1663200# diff_1004400_1657200# diff_1885200_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1166 diff_1905600_1663200# diff_1004400_1657200# diff_1905600_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1167 diff_1926000_1663200# diff_1004400_1657200# diff_1926000_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1168 diff_1946400_1663200# diff_1004400_1657200# diff_1946400_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1169 diff_1966800_1663200# diff_1004400_1657200# diff_1966800_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1170 diff_1987200_1663200# diff_1004400_1657200# diff_1987200_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1171 diff_2007600_1663200# diff_1004400_1657200# diff_2007600_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1172 diff_2028000_1663200# diff_1004400_1657200# diff_2028000_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1173 diff_2048400_1663200# diff_1004400_1657200# diff_2048400_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1174 diff_2068800_1663200# diff_1004400_1657200# diff_2068800_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1175 diff_2089200_1663200# diff_1004400_1657200# diff_2089200_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1176 diff_2109600_1663200# diff_1004400_1657200# diff_2109600_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1177 diff_2130000_1663200# diff_1004400_1657200# diff_2130000_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1178 diff_2150400_1663200# diff_1004400_1657200# diff_2150400_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1179 diff_2170800_1663200# diff_1004400_1657200# diff_2170800_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1180 diff_2191200_1663200# diff_1004400_1657200# diff_2191200_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1181 diff_2211600_1663200# diff_1004400_1657200# diff_2211600_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1182 diff_2232000_1663200# diff_1004400_1657200# diff_2232000_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1183 diff_2252400_1663200# diff_1004400_1657200# diff_2252400_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1184 diff_2272800_1663200# diff_1004400_1657200# diff_2272800_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1185 diff_2293200_1663200# diff_1004400_1657200# diff_2293200_1641600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1186 diff_1004400_1680000# Vdd Vdd GND efet w=6000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1187 diff_1008000_1641600# diff_1004400_1635600# diff_1008000_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1188 diff_1028400_1641600# diff_1004400_1635600# diff_1028400_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1189 diff_1048800_1641600# diff_1004400_1635600# diff_1048800_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1190 diff_1069200_1641600# diff_1004400_1635600# diff_1069200_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1191 diff_1089600_1641600# diff_1004400_1635600# diff_1089600_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1192 diff_1110000_1641600# diff_1004400_1635600# diff_1110000_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1193 diff_1130400_1641600# diff_1004400_1635600# diff_1130400_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1194 diff_1150800_1641600# diff_1004400_1635600# diff_1150800_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1195 diff_1171200_1641600# diff_1004400_1635600# diff_1171200_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1196 diff_1191600_1641600# diff_1004400_1635600# diff_1191600_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1197 diff_1212000_1641600# diff_1004400_1635600# diff_1212000_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1198 diff_1232400_1641600# diff_1004400_1635600# diff_1232400_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1199 diff_1252800_1641600# diff_1004400_1635600# diff_1252800_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1200 diff_1273200_1641600# diff_1004400_1635600# diff_1273200_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1201 diff_1293600_1641600# diff_1004400_1635600# diff_1293600_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1202 diff_1314000_1641600# diff_1004400_1635600# diff_1314000_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1203 diff_1334400_1641600# diff_1004400_1635600# diff_1334400_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1204 diff_1354800_1641600# diff_1004400_1635600# diff_1354800_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1205 diff_1375200_1641600# diff_1004400_1635600# diff_1375200_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1206 diff_1395600_1641600# diff_1004400_1635600# diff_1395600_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1207 diff_1416000_1641600# diff_1004400_1635600# diff_1416000_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1208 diff_1436400_1641600# diff_1004400_1635600# diff_1436400_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1209 diff_1456800_1641600# diff_1004400_1635600# diff_1456800_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1210 diff_1477200_1641600# diff_1004400_1635600# diff_1477200_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1211 diff_1497600_1641600# diff_1004400_1635600# diff_1497600_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1212 diff_1518000_1641600# diff_1004400_1635600# diff_1518000_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1213 diff_1538400_1641600# diff_1004400_1635600# diff_1538400_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1214 diff_1558800_1641600# diff_1004400_1635600# diff_1558800_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1215 diff_1579200_1641600# diff_1004400_1635600# diff_1579200_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1216 diff_1599600_1641600# diff_1004400_1635600# diff_1599600_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1217 diff_1620000_1641600# diff_1004400_1635600# diff_1620000_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1218 diff_1640400_1641600# diff_1004400_1635600# diff_1640400_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1219 diff_1660800_1641600# diff_1004400_1635600# diff_1660800_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1220 diff_1681200_1641600# diff_1004400_1635600# diff_1681200_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1221 diff_1701600_1641600# diff_1004400_1635600# diff_1701600_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1222 diff_1722000_1641600# diff_1004400_1635600# diff_1722000_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1223 diff_1742400_1641600# diff_1004400_1635600# diff_1742400_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1224 diff_1762800_1641600# diff_1004400_1635600# diff_1762800_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1225 diff_1783200_1641600# diff_1004400_1635600# diff_1783200_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1226 diff_1803600_1641600# diff_1004400_1635600# diff_1803600_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1227 diff_1824000_1641600# diff_1004400_1635600# diff_1824000_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1228 diff_1844400_1641600# diff_1004400_1635600# diff_1844400_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1229 diff_1864800_1641600# diff_1004400_1635600# diff_1864800_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1230 diff_1885200_1641600# diff_1004400_1635600# diff_1885200_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1231 diff_1905600_1641600# diff_1004400_1635600# diff_1905600_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1232 diff_1926000_1641600# diff_1004400_1635600# diff_1926000_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1233 diff_1946400_1641600# diff_1004400_1635600# diff_1946400_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1234 diff_1966800_1641600# diff_1004400_1635600# diff_1966800_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1235 diff_1987200_1641600# diff_1004400_1635600# diff_1987200_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1236 diff_2007600_1641600# diff_1004400_1635600# diff_2007600_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1237 diff_2028000_1641600# diff_1004400_1635600# diff_2028000_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1238 diff_2048400_1641600# diff_1004400_1635600# diff_2048400_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1239 diff_2068800_1641600# diff_1004400_1635600# diff_2068800_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1240 diff_2089200_1641600# diff_1004400_1635600# diff_2089200_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1241 diff_2109600_1641600# diff_1004400_1635600# diff_2109600_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1242 diff_2130000_1641600# diff_1004400_1635600# diff_2130000_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1243 diff_2150400_1641600# diff_1004400_1635600# diff_2150400_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1244 diff_2170800_1641600# diff_1004400_1635600# diff_2170800_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1245 diff_2191200_1641600# diff_1004400_1635600# diff_2191200_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1246 diff_2211600_1641600# diff_1004400_1635600# diff_2211600_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1247 diff_2232000_1641600# diff_1004400_1635600# diff_2232000_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1248 diff_2252400_1641600# diff_1004400_1635600# diff_2252400_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1249 diff_2272800_1641600# diff_1004400_1635600# diff_2272800_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1250 diff_2293200_1641600# diff_1004400_1635600# diff_2293200_1618800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1251 Vdd Vdd diff_1004400_1612800# GND efet w=6000 l=12000
+ ad=0 pd=0 as=8.5104e+08 ps=259200 
M1252 diff_1008000_1618800# diff_1004400_1612800# diff_1008000_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1253 diff_1028400_1618800# diff_1004400_1612800# diff_1028400_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1254 diff_1048800_1618800# diff_1004400_1612800# diff_1048800_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1255 diff_1069200_1618800# diff_1004400_1612800# diff_1069200_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1256 diff_1089600_1618800# diff_1004400_1612800# diff_1089600_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1257 diff_1110000_1618800# diff_1004400_1612800# diff_1110000_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1258 diff_1130400_1618800# diff_1004400_1612800# diff_1130400_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1259 diff_1150800_1618800# diff_1004400_1612800# diff_1150800_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1260 diff_1171200_1618800# diff_1004400_1612800# diff_1171200_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1261 diff_1191600_1618800# diff_1004400_1612800# diff_1191600_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1262 diff_1212000_1618800# diff_1004400_1612800# diff_1212000_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1263 diff_1232400_1618800# diff_1004400_1612800# diff_1232400_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1264 diff_1252800_1618800# diff_1004400_1612800# diff_1252800_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1265 diff_1273200_1618800# diff_1004400_1612800# diff_1273200_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1266 diff_1293600_1618800# diff_1004400_1612800# diff_1293600_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1267 diff_1314000_1618800# diff_1004400_1612800# diff_1314000_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1268 diff_1334400_1618800# diff_1004400_1612800# diff_1334400_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1269 diff_1354800_1618800# diff_1004400_1612800# diff_1354800_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1270 diff_1375200_1618800# diff_1004400_1612800# diff_1375200_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1271 diff_1395600_1618800# diff_1004400_1612800# diff_1395600_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1272 diff_1416000_1618800# diff_1004400_1612800# diff_1416000_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1273 diff_1436400_1618800# diff_1004400_1612800# diff_1436400_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1274 diff_1456800_1618800# diff_1004400_1612800# diff_1456800_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1275 diff_1477200_1618800# diff_1004400_1612800# diff_1477200_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1276 diff_1497600_1618800# diff_1004400_1612800# diff_1497600_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1277 diff_1518000_1618800# diff_1004400_1612800# diff_1518000_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1278 diff_1538400_1618800# diff_1004400_1612800# diff_1538400_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1279 diff_1558800_1618800# diff_1004400_1612800# diff_1558800_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1280 diff_1579200_1618800# diff_1004400_1612800# diff_1579200_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1281 diff_1599600_1618800# diff_1004400_1612800# diff_1599600_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1282 diff_1620000_1618800# diff_1004400_1612800# diff_1620000_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1283 diff_1640400_1618800# diff_1004400_1612800# diff_1640400_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1284 diff_1660800_1618800# diff_1004400_1612800# diff_1660800_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1285 diff_1681200_1618800# diff_1004400_1612800# diff_1681200_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1286 diff_1701600_1618800# diff_1004400_1612800# diff_1701600_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1287 diff_1722000_1618800# diff_1004400_1612800# diff_1722000_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1288 diff_1742400_1618800# diff_1004400_1612800# diff_1742400_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1289 diff_1762800_1618800# diff_1004400_1612800# diff_1762800_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1290 diff_1783200_1618800# diff_1004400_1612800# diff_1783200_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1291 diff_1803600_1618800# diff_1004400_1612800# diff_1803600_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1292 diff_1824000_1618800# diff_1004400_1612800# diff_1824000_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1293 diff_1844400_1618800# diff_1004400_1612800# diff_1844400_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1294 diff_1864800_1618800# diff_1004400_1612800# diff_1864800_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1295 diff_1885200_1618800# diff_1004400_1612800# diff_1885200_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1296 diff_1905600_1618800# diff_1004400_1612800# diff_1905600_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1297 diff_1926000_1618800# diff_1004400_1612800# diff_1926000_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1298 diff_1946400_1618800# diff_1004400_1612800# diff_1946400_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1299 diff_1966800_1618800# diff_1004400_1612800# diff_1966800_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1300 diff_1987200_1618800# diff_1004400_1612800# diff_1987200_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1301 diff_2007600_1618800# diff_1004400_1612800# diff_2007600_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1302 diff_2028000_1618800# diff_1004400_1612800# diff_2028000_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1303 diff_2048400_1618800# diff_1004400_1612800# diff_2048400_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1304 diff_2068800_1618800# diff_1004400_1612800# diff_2068800_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1305 diff_2089200_1618800# diff_1004400_1612800# diff_2089200_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1306 diff_2109600_1618800# diff_1004400_1612800# diff_2109600_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1307 diff_2130000_1618800# diff_1004400_1612800# diff_2130000_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1308 diff_2150400_1618800# diff_1004400_1612800# diff_2150400_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1309 diff_2170800_1618800# diff_1004400_1612800# diff_2170800_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1310 diff_2191200_1618800# diff_1004400_1612800# diff_2191200_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1311 diff_2211600_1618800# diff_1004400_1612800# diff_2211600_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1312 diff_2232000_1618800# diff_1004400_1612800# diff_2232000_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1313 diff_2252400_1618800# diff_1004400_1612800# diff_2252400_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1314 diff_2272800_1618800# diff_1004400_1612800# diff_2272800_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1315 diff_2293200_1618800# diff_1004400_1612800# diff_2293200_1597200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1316 diff_1004400_1612800# diff_2384400_427200# diff_2367600_1674000# GND efet w=74400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M1317 diff_2367600_1674000# diff_2413200_996000# diff_1004400_1657200# GND efet w=82800 l=7200
+ ad=0 pd=0 as=1.08e+09 ps=223200 
M1318 diff_1004400_1657200# Vdd Vdd GND efet w=7200 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1319 Vdd Vdd diff_1004400_1635600# GND efet w=7200 l=12000
+ ad=0 pd=0 as=9.4176e+08 ps=247200 
M1320 diff_1008000_1597200# diff_1004400_1591200# diff_1008000_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1321 diff_1028400_1597200# diff_1004400_1591200# diff_1028400_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1322 diff_1048800_1597200# diff_1004400_1591200# diff_1048800_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1323 diff_1069200_1597200# diff_1004400_1591200# diff_1069200_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1324 diff_1089600_1597200# diff_1004400_1591200# diff_1089600_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1325 diff_1110000_1597200# diff_1004400_1591200# diff_1110000_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1326 diff_1130400_1597200# diff_1004400_1591200# diff_1130400_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1327 diff_1150800_1597200# diff_1004400_1591200# diff_1150800_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1328 diff_1171200_1597200# diff_1004400_1591200# diff_1171200_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1329 diff_1191600_1597200# diff_1004400_1591200# diff_1191600_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1330 diff_1212000_1597200# diff_1004400_1591200# diff_1212000_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1331 diff_1232400_1597200# diff_1004400_1591200# diff_1232400_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1332 diff_1252800_1597200# diff_1004400_1591200# diff_1252800_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1333 diff_1273200_1597200# diff_1004400_1591200# diff_1273200_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1334 diff_1293600_1597200# diff_1004400_1591200# diff_1293600_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1335 diff_1314000_1597200# diff_1004400_1591200# diff_1314000_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1336 diff_1334400_1597200# diff_1004400_1591200# diff_1334400_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1337 diff_1354800_1597200# diff_1004400_1591200# diff_1354800_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1338 diff_1375200_1597200# diff_1004400_1591200# diff_1375200_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1339 diff_1395600_1597200# diff_1004400_1591200# diff_1395600_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1340 diff_1416000_1597200# diff_1004400_1591200# diff_1416000_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1341 diff_1436400_1597200# diff_1004400_1591200# diff_1436400_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1342 diff_1456800_1597200# diff_1004400_1591200# diff_1456800_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1343 diff_1477200_1597200# diff_1004400_1591200# diff_1477200_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1344 diff_1497600_1597200# diff_1004400_1591200# diff_1497600_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1345 diff_1518000_1597200# diff_1004400_1591200# diff_1518000_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1346 diff_1538400_1597200# diff_1004400_1591200# diff_1538400_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1347 diff_1558800_1597200# diff_1004400_1591200# diff_1558800_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1348 diff_1579200_1597200# diff_1004400_1591200# diff_1579200_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1349 diff_1599600_1597200# diff_1004400_1591200# diff_1599600_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1350 diff_1620000_1597200# diff_1004400_1591200# diff_1620000_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1351 diff_1640400_1597200# diff_1004400_1591200# diff_1640400_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1352 diff_1660800_1597200# diff_1004400_1591200# diff_1660800_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1353 diff_1681200_1597200# diff_1004400_1591200# diff_1681200_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1354 diff_1701600_1597200# diff_1004400_1591200# diff_1701600_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1355 diff_1722000_1597200# diff_1004400_1591200# diff_1722000_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1356 diff_1742400_1597200# diff_1004400_1591200# diff_1742400_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1357 diff_1762800_1597200# diff_1004400_1591200# diff_1762800_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1358 diff_1783200_1597200# diff_1004400_1591200# diff_1783200_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1359 diff_1803600_1597200# diff_1004400_1591200# diff_1803600_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1360 diff_1824000_1597200# diff_1004400_1591200# diff_1824000_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1361 diff_1844400_1597200# diff_1004400_1591200# diff_1844400_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1362 diff_1864800_1597200# diff_1004400_1591200# diff_1864800_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1363 diff_1885200_1597200# diff_1004400_1591200# diff_1885200_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1364 diff_1905600_1597200# diff_1004400_1591200# diff_1905600_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1365 diff_1926000_1597200# diff_1004400_1591200# diff_1926000_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1366 diff_1946400_1597200# diff_1004400_1591200# diff_1946400_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1367 diff_1966800_1597200# diff_1004400_1591200# diff_1966800_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1368 diff_1987200_1597200# diff_1004400_1591200# diff_1987200_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1369 diff_2007600_1597200# diff_1004400_1591200# diff_2007600_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1370 diff_2028000_1597200# diff_1004400_1591200# diff_2028000_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1371 diff_2048400_1597200# diff_1004400_1591200# diff_2048400_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1372 diff_2068800_1597200# diff_1004400_1591200# diff_2068800_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1373 diff_2089200_1597200# diff_1004400_1591200# diff_2089200_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1374 diff_2109600_1597200# diff_1004400_1591200# diff_2109600_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1375 diff_2130000_1597200# diff_1004400_1591200# diff_2130000_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1376 diff_2150400_1597200# diff_1004400_1591200# diff_2150400_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1377 diff_2170800_1597200# diff_1004400_1591200# diff_2170800_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1378 diff_2191200_1597200# diff_1004400_1591200# diff_2191200_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1379 diff_2211600_1597200# diff_1004400_1591200# diff_2211600_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1380 diff_2232000_1597200# diff_1004400_1591200# diff_2232000_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1381 diff_2252400_1597200# diff_1004400_1591200# diff_2252400_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1382 diff_2272800_1597200# diff_1004400_1591200# diff_2272800_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1383 diff_2293200_1597200# diff_1004400_1591200# diff_2293200_1574400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1384 diff_2367600_1585200# diff_2361600_427200# diff_1004400_1591200# GND efet w=87600 l=6600
+ ad=-4.71767e+08 pd=732000 as=8.8992e+08 ps=225600 
M1385 diff_1004400_1635600# diff_2431200_979200# diff_2367600_1674000# GND efet w=79200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M1386 diff_1008000_1574400# diff_1004400_1568400# diff_1008000_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1387 diff_1028400_1574400# diff_1004400_1568400# diff_1028400_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1388 diff_1048800_1574400# diff_1004400_1568400# diff_1048800_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1389 diff_1069200_1574400# diff_1004400_1568400# diff_1069200_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1390 diff_1089600_1574400# diff_1004400_1568400# diff_1089600_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1391 diff_1110000_1574400# diff_1004400_1568400# diff_1110000_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1392 diff_1130400_1574400# diff_1004400_1568400# diff_1130400_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1393 diff_1150800_1574400# diff_1004400_1568400# diff_1150800_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1394 diff_1171200_1574400# diff_1004400_1568400# diff_1171200_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1395 diff_1191600_1574400# diff_1004400_1568400# diff_1191600_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1396 diff_1212000_1574400# diff_1004400_1568400# diff_1212000_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1397 diff_1232400_1574400# diff_1004400_1568400# diff_1232400_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1398 diff_1252800_1574400# diff_1004400_1568400# diff_1252800_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1399 diff_1273200_1574400# diff_1004400_1568400# diff_1273200_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1400 diff_1293600_1574400# diff_1004400_1568400# diff_1293600_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1401 diff_1314000_1574400# diff_1004400_1568400# diff_1314000_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1402 diff_1334400_1574400# diff_1004400_1568400# diff_1334400_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1403 diff_1354800_1574400# diff_1004400_1568400# diff_1354800_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1404 diff_1375200_1574400# diff_1004400_1568400# diff_1375200_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1405 diff_1395600_1574400# diff_1004400_1568400# diff_1395600_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1406 diff_1416000_1574400# diff_1004400_1568400# diff_1416000_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1407 diff_1436400_1574400# diff_1004400_1568400# diff_1436400_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1408 diff_1456800_1574400# diff_1004400_1568400# diff_1456800_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1409 diff_1477200_1574400# diff_1004400_1568400# diff_1477200_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1410 diff_1497600_1574400# diff_1004400_1568400# diff_1497600_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1411 diff_1518000_1574400# diff_1004400_1568400# diff_1518000_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1412 diff_1538400_1574400# diff_1004400_1568400# diff_1538400_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1413 diff_1558800_1574400# diff_1004400_1568400# diff_1558800_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1414 diff_1579200_1574400# diff_1004400_1568400# diff_1579200_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1415 diff_1599600_1574400# diff_1004400_1568400# diff_1599600_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1416 diff_1620000_1574400# diff_1004400_1568400# diff_1620000_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1417 diff_1640400_1574400# diff_1004400_1568400# diff_1640400_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1418 diff_1660800_1574400# diff_1004400_1568400# diff_1660800_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1419 diff_1681200_1574400# diff_1004400_1568400# diff_1681200_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1420 diff_1701600_1574400# diff_1004400_1568400# diff_1701600_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1421 diff_1722000_1574400# diff_1004400_1568400# diff_1722000_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1422 diff_1742400_1574400# diff_1004400_1568400# diff_1742400_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1423 diff_1762800_1574400# diff_1004400_1568400# diff_1762800_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1424 diff_1783200_1574400# diff_1004400_1568400# diff_1783200_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1425 diff_1803600_1574400# diff_1004400_1568400# diff_1803600_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1426 diff_1824000_1574400# diff_1004400_1568400# diff_1824000_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1427 diff_1844400_1574400# diff_1004400_1568400# diff_1844400_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1428 diff_1864800_1574400# diff_1004400_1568400# diff_1864800_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1429 diff_1885200_1574400# diff_1004400_1568400# diff_1885200_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1430 diff_1905600_1574400# diff_1004400_1568400# diff_1905600_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1431 diff_1926000_1574400# diff_1004400_1568400# diff_1926000_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1432 diff_1946400_1574400# diff_1004400_1568400# diff_1946400_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1433 diff_1966800_1574400# diff_1004400_1568400# diff_1966800_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1434 diff_1987200_1574400# diff_1004400_1568400# diff_1987200_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1435 diff_2007600_1574400# diff_1004400_1568400# diff_2007600_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1436 diff_2028000_1574400# diff_1004400_1568400# diff_2028000_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1437 diff_2048400_1574400# diff_1004400_1568400# diff_2048400_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1438 diff_2068800_1574400# diff_1004400_1568400# diff_2068800_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1439 diff_2089200_1574400# diff_1004400_1568400# diff_2089200_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1440 diff_2109600_1574400# diff_1004400_1568400# diff_2109600_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1441 diff_2130000_1574400# diff_1004400_1568400# diff_2130000_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1442 diff_2150400_1574400# diff_1004400_1568400# diff_2150400_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1443 diff_2170800_1574400# diff_1004400_1568400# diff_2170800_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1444 diff_2191200_1574400# diff_1004400_1568400# diff_2191200_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1445 diff_2211600_1574400# diff_1004400_1568400# diff_2211600_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1446 diff_2232000_1574400# diff_1004400_1568400# diff_2232000_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1447 diff_2252400_1574400# diff_1004400_1568400# diff_2252400_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1448 diff_2272800_1574400# diff_1004400_1568400# diff_2272800_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1449 diff_2293200_1574400# diff_1004400_1568400# diff_2293200_1552800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1450 diff_831600_1504800# diff_831600_1504800# diff_831600_1504800# GND efet w=600 l=1800
+ ad=0 pd=0 as=0 ps=0 
M1451 diff_355200_1366800# diff_338400_1662000# GND GND efet w=97200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1452 diff_338400_1662000# diff_408000_1448400# GND GND efet w=187200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1453 diff_664800_1365600# diff_673200_1506000# diff_664800_1365600# GND efet w=61200 l=3600
+ ad=0 pd=0 as=0 ps=0 
M1454 diff_649200_1662000# diff_738000_1506000# diff_649200_1662000# GND efet w=57000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M1455 GND diff_189600_804000# diff_355200_1366800# GND efet w=189600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1456 diff_510000_1366800# diff_494400_1662000# GND GND efet w=97200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1457 diff_494400_1662000# diff_562800_1448400# GND GND efet w=188400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1458 diff_820800_1365600# diff_831600_1504800# diff_820800_1365600# GND efet w=42600 l=13800
+ ad=0 pd=0 as=0 ps=0 
M1459 diff_886800_1546800# diff_886800_1546800# diff_886800_1546800# GND efet w=600 l=1800
+ ad=0 pd=0 as=0 ps=0 
M1460 diff_1004400_1591200# Vdd Vdd GND efet w=6000 l=13200
+ ad=0 pd=0 as=0 ps=0 
M1461 diff_1008000_1552800# diff_1004400_1546800# diff_1008000_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1462 diff_1028400_1552800# diff_1004400_1546800# diff_1028400_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1463 diff_1048800_1552800# diff_1004400_1546800# diff_1048800_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1464 diff_1069200_1552800# diff_1004400_1546800# diff_1069200_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1465 diff_1089600_1552800# diff_1004400_1546800# diff_1089600_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1466 diff_1110000_1552800# diff_1004400_1546800# diff_1110000_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1467 diff_1130400_1552800# diff_1004400_1546800# diff_1130400_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1468 diff_1150800_1552800# diff_1004400_1546800# diff_1150800_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1469 diff_1171200_1552800# diff_1004400_1546800# diff_1171200_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1470 diff_1191600_1552800# diff_1004400_1546800# diff_1191600_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1471 diff_1212000_1552800# diff_1004400_1546800# diff_1212000_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1472 diff_1232400_1552800# diff_1004400_1546800# diff_1232400_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1473 diff_1252800_1552800# diff_1004400_1546800# diff_1252800_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1474 diff_1273200_1552800# diff_1004400_1546800# diff_1273200_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1475 diff_1293600_1552800# diff_1004400_1546800# diff_1293600_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1476 diff_1314000_1552800# diff_1004400_1546800# diff_1314000_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1477 diff_1334400_1552800# diff_1004400_1546800# diff_1334400_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1478 diff_1354800_1552800# diff_1004400_1546800# diff_1354800_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1479 diff_1375200_1552800# diff_1004400_1546800# diff_1375200_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1480 diff_1395600_1552800# diff_1004400_1546800# diff_1395600_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1481 diff_1416000_1552800# diff_1004400_1546800# diff_1416000_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1482 diff_1436400_1552800# diff_1004400_1546800# diff_1436400_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1483 diff_1456800_1552800# diff_1004400_1546800# diff_1456800_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1484 diff_1477200_1552800# diff_1004400_1546800# diff_1477200_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1485 diff_1497600_1552800# diff_1004400_1546800# diff_1497600_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1486 diff_1518000_1552800# diff_1004400_1546800# diff_1518000_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1487 diff_1538400_1552800# diff_1004400_1546800# diff_1538400_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1488 diff_1558800_1552800# diff_1004400_1546800# diff_1558800_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1489 diff_1579200_1552800# diff_1004400_1546800# diff_1579200_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1490 diff_1599600_1552800# diff_1004400_1546800# diff_1599600_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1491 diff_1620000_1552800# diff_1004400_1546800# diff_1620000_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1492 diff_1640400_1552800# diff_1004400_1546800# diff_1640400_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1493 diff_1660800_1552800# diff_1004400_1546800# diff_1660800_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1494 diff_1681200_1552800# diff_1004400_1546800# diff_1681200_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1495 diff_1701600_1552800# diff_1004400_1546800# diff_1701600_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1496 diff_1722000_1552800# diff_1004400_1546800# diff_1722000_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1497 diff_1742400_1552800# diff_1004400_1546800# diff_1742400_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1498 diff_1762800_1552800# diff_1004400_1546800# diff_1762800_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1499 diff_1783200_1552800# diff_1004400_1546800# diff_1783200_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1500 diff_1803600_1552800# diff_1004400_1546800# diff_1803600_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1501 diff_1824000_1552800# diff_1004400_1546800# diff_1824000_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1502 diff_1844400_1552800# diff_1004400_1546800# diff_1844400_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1503 diff_1864800_1552800# diff_1004400_1546800# diff_1864800_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1504 diff_1885200_1552800# diff_1004400_1546800# diff_1885200_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1505 diff_1905600_1552800# diff_1004400_1546800# diff_1905600_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1506 diff_1926000_1552800# diff_1004400_1546800# diff_1926000_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1507 diff_1946400_1552800# diff_1004400_1546800# diff_1946400_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1508 diff_1966800_1552800# diff_1004400_1546800# diff_1966800_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1509 diff_1987200_1552800# diff_1004400_1546800# diff_1987200_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1510 diff_2007600_1552800# diff_1004400_1546800# diff_2007600_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1511 diff_2028000_1552800# diff_1004400_1546800# diff_2028000_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1512 diff_2048400_1552800# diff_1004400_1546800# diff_2048400_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1513 diff_2068800_1552800# diff_1004400_1546800# diff_2068800_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1514 diff_2089200_1552800# diff_1004400_1546800# diff_2089200_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1515 diff_2109600_1552800# diff_1004400_1546800# diff_2109600_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1516 diff_2130000_1552800# diff_1004400_1546800# diff_2130000_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1517 diff_2150400_1552800# diff_1004400_1546800# diff_2150400_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1518 diff_2170800_1552800# diff_1004400_1546800# diff_2170800_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1519 diff_2191200_1552800# diff_1004400_1546800# diff_2191200_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1520 diff_2211600_1552800# diff_1004400_1546800# diff_2211600_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1521 diff_2232000_1552800# diff_1004400_1546800# diff_2232000_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1522 diff_2252400_1552800# diff_1004400_1546800# diff_2252400_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1523 diff_2272800_1552800# diff_1004400_1546800# diff_2272800_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1524 diff_2293200_1552800# diff_1004400_1546800# diff_2293200_1530000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1525 diff_804000_1662000# diff_886800_1546800# diff_804000_1662000# GND efet w=50400 l=10200
+ ad=0 pd=0 as=0 ps=0 
M1526 Vdd Vdd diff_1004400_1524000# GND efet w=6000 l=13200
+ ad=0 pd=0 as=8.5104e+08 ps=259200 
M1527 diff_1008000_1530000# diff_1004400_1524000# diff_1008000_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1528 diff_1028400_1530000# diff_1004400_1524000# diff_1028400_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1529 diff_1048800_1530000# diff_1004400_1524000# diff_1048800_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1530 diff_1069200_1530000# diff_1004400_1524000# diff_1069200_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1531 diff_1089600_1530000# diff_1004400_1524000# diff_1089600_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1532 diff_1110000_1530000# diff_1004400_1524000# diff_1110000_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1533 diff_1130400_1530000# diff_1004400_1524000# diff_1130400_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1534 diff_1150800_1530000# diff_1004400_1524000# diff_1150800_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1535 diff_1171200_1530000# diff_1004400_1524000# diff_1171200_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1536 diff_1191600_1530000# diff_1004400_1524000# diff_1191600_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1537 diff_1212000_1530000# diff_1004400_1524000# diff_1212000_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1538 diff_1232400_1530000# diff_1004400_1524000# diff_1232400_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1539 diff_1252800_1530000# diff_1004400_1524000# diff_1252800_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1540 diff_1273200_1530000# diff_1004400_1524000# diff_1273200_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1541 diff_1293600_1530000# diff_1004400_1524000# diff_1293600_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1542 diff_1314000_1530000# diff_1004400_1524000# diff_1314000_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1543 diff_1334400_1530000# diff_1004400_1524000# diff_1334400_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1544 diff_1354800_1530000# diff_1004400_1524000# diff_1354800_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1545 diff_1375200_1530000# diff_1004400_1524000# diff_1375200_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1546 diff_1395600_1530000# diff_1004400_1524000# diff_1395600_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1547 diff_1416000_1530000# diff_1004400_1524000# diff_1416000_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1548 diff_1436400_1530000# diff_1004400_1524000# diff_1436400_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1549 diff_1456800_1530000# diff_1004400_1524000# diff_1456800_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1550 diff_1477200_1530000# diff_1004400_1524000# diff_1477200_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1551 diff_1497600_1530000# diff_1004400_1524000# diff_1497600_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1552 diff_1518000_1530000# diff_1004400_1524000# diff_1518000_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1553 diff_1538400_1530000# diff_1004400_1524000# diff_1538400_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1554 diff_1558800_1530000# diff_1004400_1524000# diff_1558800_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1555 diff_1579200_1530000# diff_1004400_1524000# diff_1579200_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1556 diff_1599600_1530000# diff_1004400_1524000# diff_1599600_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1557 diff_1620000_1530000# diff_1004400_1524000# diff_1620000_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1558 diff_1640400_1530000# diff_1004400_1524000# diff_1640400_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1559 diff_1660800_1530000# diff_1004400_1524000# diff_1660800_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1560 diff_1681200_1530000# diff_1004400_1524000# diff_1681200_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1561 diff_1701600_1530000# diff_1004400_1524000# diff_1701600_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1562 diff_1722000_1530000# diff_1004400_1524000# diff_1722000_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1563 diff_1742400_1530000# diff_1004400_1524000# diff_1742400_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1564 diff_1762800_1530000# diff_1004400_1524000# diff_1762800_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1565 diff_1783200_1530000# diff_1004400_1524000# diff_1783200_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1566 diff_1803600_1530000# diff_1004400_1524000# diff_1803600_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1567 diff_1824000_1530000# diff_1004400_1524000# diff_1824000_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1568 diff_1844400_1530000# diff_1004400_1524000# diff_1844400_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1569 diff_1864800_1530000# diff_1004400_1524000# diff_1864800_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1570 diff_1885200_1530000# diff_1004400_1524000# diff_1885200_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1571 diff_1905600_1530000# diff_1004400_1524000# diff_1905600_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1572 diff_1926000_1530000# diff_1004400_1524000# diff_1926000_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1573 diff_1946400_1530000# diff_1004400_1524000# diff_1946400_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1574 diff_1966800_1530000# diff_1004400_1524000# diff_1966800_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1575 diff_1987200_1530000# diff_1004400_1524000# diff_1987200_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1576 diff_2007600_1530000# diff_1004400_1524000# diff_2007600_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1577 diff_2028000_1530000# diff_1004400_1524000# diff_2028000_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1578 diff_2048400_1530000# diff_1004400_1524000# diff_2048400_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1579 diff_2068800_1530000# diff_1004400_1524000# diff_2068800_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1580 diff_2089200_1530000# diff_1004400_1524000# diff_2089200_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1581 diff_2109600_1530000# diff_1004400_1524000# diff_2109600_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1582 diff_2130000_1530000# diff_1004400_1524000# diff_2130000_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1583 diff_2150400_1530000# diff_1004400_1524000# diff_2150400_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1584 diff_2170800_1530000# diff_1004400_1524000# diff_2170800_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1585 diff_2191200_1530000# diff_1004400_1524000# diff_2191200_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1586 diff_2211600_1530000# diff_1004400_1524000# diff_2211600_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1587 diff_2232000_1530000# diff_1004400_1524000# diff_2232000_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1588 diff_2252400_1530000# diff_1004400_1524000# diff_2252400_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1589 diff_2272800_1530000# diff_1004400_1524000# diff_2272800_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1590 diff_2293200_1530000# diff_1004400_1524000# diff_2293200_1508400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1591 diff_1004400_1524000# diff_2384400_427200# diff_2367600_1585200# GND efet w=74400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M1592 diff_2367600_1585200# diff_2413200_996000# diff_1004400_1568400# GND efet w=84600 l=6600
+ ad=0 pd=0 as=1.1232e+09 ps=223200 
M1593 diff_1004400_1568400# Vdd Vdd GND efet w=7200 l=14400
+ ad=0 pd=0 as=0 ps=0 
M1594 Vdd Vdd diff_1004400_1546800# GND efet w=7200 l=13200
+ ad=0 pd=0 as=9.4176e+08 ps=247200 
M1595 diff_1008000_1508400# diff_1004400_1502400# diff_1008000_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1596 diff_1028400_1508400# diff_1004400_1502400# diff_1028400_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1597 diff_1048800_1508400# diff_1004400_1502400# diff_1048800_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1598 diff_1069200_1508400# diff_1004400_1502400# diff_1069200_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1599 diff_1089600_1508400# diff_1004400_1502400# diff_1089600_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1600 diff_1110000_1508400# diff_1004400_1502400# diff_1110000_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1601 diff_1130400_1508400# diff_1004400_1502400# diff_1130400_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1602 diff_1150800_1508400# diff_1004400_1502400# diff_1150800_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1603 diff_1171200_1508400# diff_1004400_1502400# diff_1171200_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1604 diff_1191600_1508400# diff_1004400_1502400# diff_1191600_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1605 diff_1212000_1508400# diff_1004400_1502400# diff_1212000_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1606 diff_1232400_1508400# diff_1004400_1502400# diff_1232400_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1607 diff_1252800_1508400# diff_1004400_1502400# diff_1252800_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1608 diff_1273200_1508400# diff_1004400_1502400# diff_1273200_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1609 diff_1293600_1508400# diff_1004400_1502400# diff_1293600_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1610 diff_1314000_1508400# diff_1004400_1502400# diff_1314000_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1611 diff_1334400_1508400# diff_1004400_1502400# diff_1334400_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1612 diff_1354800_1508400# diff_1004400_1502400# diff_1354800_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1613 diff_1375200_1508400# diff_1004400_1502400# diff_1375200_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1614 diff_1395600_1508400# diff_1004400_1502400# diff_1395600_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1615 diff_1416000_1508400# diff_1004400_1502400# diff_1416000_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1616 diff_1436400_1508400# diff_1004400_1502400# diff_1436400_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1617 diff_1456800_1508400# diff_1004400_1502400# diff_1456800_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1618 diff_1477200_1508400# diff_1004400_1502400# diff_1477200_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1619 diff_1497600_1508400# diff_1004400_1502400# diff_1497600_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1620 diff_1518000_1508400# diff_1004400_1502400# diff_1518000_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1621 diff_1538400_1508400# diff_1004400_1502400# diff_1538400_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1622 diff_1558800_1508400# diff_1004400_1502400# diff_1558800_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1623 diff_1579200_1508400# diff_1004400_1502400# diff_1579200_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1624 diff_1599600_1508400# diff_1004400_1502400# diff_1599600_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1625 diff_1620000_1508400# diff_1004400_1502400# diff_1620000_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1626 diff_1640400_1508400# diff_1004400_1502400# diff_1640400_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1627 diff_1660800_1508400# diff_1004400_1502400# diff_1660800_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1628 diff_1681200_1508400# diff_1004400_1502400# diff_1681200_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1629 diff_1701600_1508400# diff_1004400_1502400# diff_1701600_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1630 diff_1722000_1508400# diff_1004400_1502400# diff_1722000_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1631 diff_1742400_1508400# diff_1004400_1502400# diff_1742400_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1632 diff_1762800_1508400# diff_1004400_1502400# diff_1762800_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1633 diff_1783200_1508400# diff_1004400_1502400# diff_1783200_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1634 diff_1803600_1508400# diff_1004400_1502400# diff_1803600_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1635 diff_1824000_1508400# diff_1004400_1502400# diff_1824000_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1636 diff_1844400_1508400# diff_1004400_1502400# diff_1844400_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1637 diff_1864800_1508400# diff_1004400_1502400# diff_1864800_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1638 diff_1885200_1508400# diff_1004400_1502400# diff_1885200_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1639 diff_1905600_1508400# diff_1004400_1502400# diff_1905600_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1640 diff_1926000_1508400# diff_1004400_1502400# diff_1926000_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1641 diff_1946400_1508400# diff_1004400_1502400# diff_1946400_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1642 diff_1966800_1508400# diff_1004400_1502400# diff_1966800_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1643 diff_1987200_1508400# diff_1004400_1502400# diff_1987200_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1644 diff_2007600_1508400# diff_1004400_1502400# diff_2007600_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1645 diff_2028000_1508400# diff_1004400_1502400# diff_2028000_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1646 diff_2048400_1508400# diff_1004400_1502400# diff_2048400_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1647 diff_2068800_1508400# diff_1004400_1502400# diff_2068800_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1648 diff_2089200_1508400# diff_1004400_1502400# diff_2089200_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1649 diff_2109600_1508400# diff_1004400_1502400# diff_2109600_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1650 diff_2130000_1508400# diff_1004400_1502400# diff_2130000_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1651 diff_2150400_1508400# diff_1004400_1502400# diff_2150400_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1652 diff_2170800_1508400# diff_1004400_1502400# diff_2170800_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1653 diff_2191200_1508400# diff_1004400_1502400# diff_2191200_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1654 diff_2211600_1508400# diff_1004400_1502400# diff_2211600_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1655 diff_2232000_1508400# diff_1004400_1502400# diff_2232000_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1656 diff_2252400_1508400# diff_1004400_1502400# diff_2252400_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1657 diff_2272800_1508400# diff_1004400_1502400# diff_2272800_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1658 diff_2293200_1508400# diff_1004400_1502400# diff_2293200_1485600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1659 diff_338400_1662000# diff_189600_804000# GND GND efet w=190800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1660 GND diff_189600_804000# diff_510000_1366800# GND efet w=189600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1661 diff_664800_1365600# diff_649200_1662000# GND GND efet w=97200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1662 diff_649200_1662000# diff_718800_1448400# GND GND efet w=188400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1663 diff_494400_1662000# diff_189600_804000# GND GND efet w=190800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1664 GND diff_189600_804000# diff_664800_1365600# GND efet w=190800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1665 diff_820800_1365600# diff_804000_1662000# GND GND efet w=97200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1666 diff_804000_1662000# diff_873600_1448400# GND GND efet w=188400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1667 diff_2367600_1494000# diff_2361600_427200# diff_1004400_1502400# GND efet w=88200 l=7200
+ ad=-4.32887e+08 pd=717600 as=9.4176e+08 ps=230400 
M1668 diff_1004400_1546800# diff_2431200_979200# diff_2367600_1585200# GND efet w=79200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M1669 diff_2437200_1698000# diff_2488800_853200# diff_2367600_1585200# GND efet w=154800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1670 diff_2367600_1674000# diff_2505600_919200# diff_2437200_1698000# GND efet w=160800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1671 diff_2433600_1742400# Vdd Vdd GND efet w=7200 l=14400
+ ad=0 pd=0 as=0 ps=0 
M1672 diff_2751600_1686000# diff_2751600_1686000# diff_2751600_1686000# GND efet w=1200 l=1800
+ ad=8.5968e+08 pd=232800 as=0 ps=0 
M1673 diff_2743200_1714800# diff_2664000_1422000# diff_2743200_1702800# GND efet w=40800 l=6000
+ ad=0 pd=0 as=4.3776e+08 ps=120000 
M1674 diff_2751600_1686000# diff_2751600_1686000# diff_2751600_1686000# GND efet w=600 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1675 GND diff_2682000_1690800# diff_2664000_1686000# GND efet w=22800 l=6000
+ ad=0 pd=0 as=7.4304e+08 ps=216000 
M1676 diff_2743200_1702800# diff_2649600_1519200# diff_2751600_1686000# GND efet w=42000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M1677 diff_2664000_1686000# diff_2664000_1686000# diff_2664000_1686000# GND efet w=1200 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1678 GND d3 diff_2828400_1086000# GND efet w=162000 l=6000
+ ad=0 pd=0 as=1.82592e+09 ps=355200 
M1679 diff_2664000_1686000# Vdd Vdd GND efet w=6600 l=38400
+ ad=0 pd=0 as=0 ps=0 
M1680 diff_2682000_1690800# diff_2682000_1690800# diff_2682000_1690800# GND efet w=1800 l=4200
+ ad=1.44e+08 pd=50400 as=0 ps=0 
M1681 Vdd Vdd Vdd GND efet w=600 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1682 Vdd Vdd Vdd GND efet w=1200 l=2400
+ ad=0 pd=0 as=0 ps=0 
M1683 diff_2682000_1690800# diff_2682000_1690800# diff_2682000_1690800# GND efet w=1200 l=3000
+ ad=0 pd=0 as=0 ps=0 
M1684 Vdd Vdd diff_2751600_1686000# GND efet w=7200 l=32400
+ ad=0 pd=0 as=0 ps=0 
M1685 diff_2802000_1732800# Vdd Vdd GND efet w=6000 l=21600
+ ad=0 pd=0 as=0 ps=0 
M1686 diff_2649600_1428000# Vdd Vdd GND efet w=7200 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1687 diff_2828400_1086000# Vdd Vdd GND efet w=9600 l=15600
+ ad=0 pd=0 as=0 ps=0 
M1688 diff_2682000_1690800# diff_2613600_1719600# diff_2710800_1356000# GND efet w=12000 l=7200
+ ad=0 pd=0 as=1.58256e+09 ps=362400 
M1689 diff_2828400_1273200# Vdd Vdd GND efet w=9600 l=15600
+ ad=1.20096e+09 pd=196800 as=0 ps=0 
M1690 GND diff_2828400_1086000# diff_2828400_1273200# GND efet w=45600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M1691 diff_2664000_1686000# diff_2649600_1519200# GND GND efet w=15600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M1692 sync clk2 diff_2767200_1582800# GND efet w=12000 l=6000
+ ad=0 pd=0 as=1.5264e+08 ps=52800 
M1693 diff_2767200_1582800# diff_2767200_1582800# diff_2767200_1582800# GND efet w=1200 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1694 diff_2767200_1582800# diff_2767200_1582800# diff_2767200_1582800# GND efet w=600 l=1800
+ ad=0 pd=0 as=0 ps=0 
M1695 GND diff_2649600_1519200# diff_1657200_1702800# GND efet w=294000 l=6000
+ ad=0 pd=0 as=9.33673e+08 ps=1.0632e+06 
M1696 diff_1657200_1702800# diff_2592000_1532400# diff_1657200_1702800# GND efet w=55200 l=16800
+ ad=0 pd=0 as=0 ps=0 
M1697 diff_1657200_1702800# diff_2592000_1532400# Vdd GND efet w=15600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M1698 diff_649200_1662000# diff_189600_804000# GND GND efet w=189600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1699 GND diff_189600_804000# diff_820800_1365600# GND efet w=189600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1700 diff_1008000_1485600# diff_1004400_1479600# diff_1008000_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1701 diff_1028400_1485600# diff_1004400_1479600# diff_1028400_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1702 diff_1048800_1485600# diff_1004400_1479600# diff_1048800_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1703 diff_1069200_1485600# diff_1004400_1479600# diff_1069200_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1704 diff_1089600_1485600# diff_1004400_1479600# diff_1089600_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1705 diff_1110000_1485600# diff_1004400_1479600# diff_1110000_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1706 diff_1130400_1485600# diff_1004400_1479600# diff_1130400_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1707 diff_1150800_1485600# diff_1004400_1479600# diff_1150800_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1708 diff_1171200_1485600# diff_1004400_1479600# diff_1171200_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1709 diff_1191600_1485600# diff_1004400_1479600# diff_1191600_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1710 diff_1212000_1485600# diff_1004400_1479600# diff_1212000_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1711 diff_1232400_1485600# diff_1004400_1479600# diff_1232400_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1712 diff_1252800_1485600# diff_1004400_1479600# diff_1252800_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1713 diff_1273200_1485600# diff_1004400_1479600# diff_1273200_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1714 diff_1293600_1485600# diff_1004400_1479600# diff_1293600_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1715 diff_1314000_1485600# diff_1004400_1479600# diff_1314000_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1716 diff_1334400_1485600# diff_1004400_1479600# diff_1334400_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1717 diff_1354800_1485600# diff_1004400_1479600# diff_1354800_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1718 diff_1375200_1485600# diff_1004400_1479600# diff_1375200_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1719 diff_1395600_1485600# diff_1004400_1479600# diff_1395600_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1720 diff_1416000_1485600# diff_1004400_1479600# diff_1416000_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1721 diff_1436400_1485600# diff_1004400_1479600# diff_1436400_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1722 diff_1456800_1485600# diff_1004400_1479600# diff_1456800_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1723 diff_1477200_1485600# diff_1004400_1479600# diff_1477200_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1724 diff_1497600_1485600# diff_1004400_1479600# diff_1497600_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1725 diff_1518000_1485600# diff_1004400_1479600# diff_1518000_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1726 diff_1538400_1485600# diff_1004400_1479600# diff_1538400_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1727 diff_1558800_1485600# diff_1004400_1479600# diff_1558800_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1728 diff_1579200_1485600# diff_1004400_1479600# diff_1579200_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1729 diff_1599600_1485600# diff_1004400_1479600# diff_1599600_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1730 diff_1620000_1485600# diff_1004400_1479600# diff_1620000_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1731 diff_1640400_1485600# diff_1004400_1479600# diff_1640400_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1732 diff_1660800_1485600# diff_1004400_1479600# diff_1660800_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1733 diff_1681200_1485600# diff_1004400_1479600# diff_1681200_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1734 diff_1701600_1485600# diff_1004400_1479600# diff_1701600_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1735 diff_1722000_1485600# diff_1004400_1479600# diff_1722000_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1736 diff_1742400_1485600# diff_1004400_1479600# diff_1742400_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1737 diff_1762800_1485600# diff_1004400_1479600# diff_1762800_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1738 diff_1783200_1485600# diff_1004400_1479600# diff_1783200_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1739 diff_1803600_1485600# diff_1004400_1479600# diff_1803600_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1740 diff_1824000_1485600# diff_1004400_1479600# diff_1824000_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1741 diff_1844400_1485600# diff_1004400_1479600# diff_1844400_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1742 diff_1864800_1485600# diff_1004400_1479600# diff_1864800_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1743 diff_1885200_1485600# diff_1004400_1479600# diff_1885200_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1744 diff_1905600_1485600# diff_1004400_1479600# diff_1905600_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1745 diff_1926000_1485600# diff_1004400_1479600# diff_1926000_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1746 diff_1946400_1485600# diff_1004400_1479600# diff_1946400_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1747 diff_1966800_1485600# diff_1004400_1479600# diff_1966800_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1748 diff_1987200_1485600# diff_1004400_1479600# diff_1987200_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1749 diff_2007600_1485600# diff_1004400_1479600# diff_2007600_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1750 diff_2028000_1485600# diff_1004400_1479600# diff_2028000_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1751 diff_2048400_1485600# diff_1004400_1479600# diff_2048400_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1752 diff_2068800_1485600# diff_1004400_1479600# diff_2068800_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1753 diff_2089200_1485600# diff_1004400_1479600# diff_2089200_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1754 diff_2109600_1485600# diff_1004400_1479600# diff_2109600_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1755 diff_2130000_1485600# diff_1004400_1479600# diff_2130000_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1756 diff_2150400_1485600# diff_1004400_1479600# diff_2150400_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1757 diff_2170800_1485600# diff_1004400_1479600# diff_2170800_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1758 diff_2191200_1485600# diff_1004400_1479600# diff_2191200_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1759 diff_2211600_1485600# diff_1004400_1479600# diff_2211600_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1760 diff_2232000_1485600# diff_1004400_1479600# diff_2232000_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1761 diff_2252400_1485600# diff_1004400_1479600# diff_2252400_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1762 diff_2272800_1485600# diff_1004400_1479600# diff_2272800_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1763 diff_2293200_1485600# diff_1004400_1479600# diff_2293200_1464000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1764 diff_1004400_1502400# Vdd Vdd GND efet w=6000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M1765 diff_1008000_1464000# diff_1004400_1458000# diff_1008000_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1766 diff_1028400_1464000# diff_1004400_1458000# diff_1028400_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1767 diff_1048800_1464000# diff_1004400_1458000# diff_1048800_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1768 diff_1069200_1464000# diff_1004400_1458000# diff_1069200_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1769 diff_1089600_1464000# diff_1004400_1458000# diff_1089600_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1770 diff_1110000_1464000# diff_1004400_1458000# diff_1110000_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1771 diff_1130400_1464000# diff_1004400_1458000# diff_1130400_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1772 diff_1150800_1464000# diff_1004400_1458000# diff_1150800_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1773 diff_1171200_1464000# diff_1004400_1458000# diff_1171200_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1774 diff_1191600_1464000# diff_1004400_1458000# diff_1191600_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1775 diff_1212000_1464000# diff_1004400_1458000# diff_1212000_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1776 diff_1232400_1464000# diff_1004400_1458000# diff_1232400_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1777 diff_1252800_1464000# diff_1004400_1458000# diff_1252800_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1778 diff_1273200_1464000# diff_1004400_1458000# diff_1273200_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1779 diff_1293600_1464000# diff_1004400_1458000# diff_1293600_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1780 diff_1314000_1464000# diff_1004400_1458000# diff_1314000_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1781 diff_1334400_1464000# diff_1004400_1458000# diff_1334400_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1782 diff_1354800_1464000# diff_1004400_1458000# diff_1354800_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1783 diff_1375200_1464000# diff_1004400_1458000# diff_1375200_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1784 diff_1395600_1464000# diff_1004400_1458000# diff_1395600_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1785 diff_1416000_1464000# diff_1004400_1458000# diff_1416000_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1786 diff_1436400_1464000# diff_1004400_1458000# diff_1436400_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1787 diff_1456800_1464000# diff_1004400_1458000# diff_1456800_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1788 diff_1477200_1464000# diff_1004400_1458000# diff_1477200_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1789 diff_1497600_1464000# diff_1004400_1458000# diff_1497600_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1790 diff_1518000_1464000# diff_1004400_1458000# diff_1518000_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1791 diff_1538400_1464000# diff_1004400_1458000# diff_1538400_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1792 diff_1558800_1464000# diff_1004400_1458000# diff_1558800_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1793 diff_1579200_1464000# diff_1004400_1458000# diff_1579200_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1794 diff_1599600_1464000# diff_1004400_1458000# diff_1599600_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1795 diff_1620000_1464000# diff_1004400_1458000# diff_1620000_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1796 diff_1640400_1464000# diff_1004400_1458000# diff_1640400_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1797 diff_1660800_1464000# diff_1004400_1458000# diff_1660800_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1798 diff_1681200_1464000# diff_1004400_1458000# diff_1681200_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1799 diff_1701600_1464000# diff_1004400_1458000# diff_1701600_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1800 diff_1722000_1464000# diff_1004400_1458000# diff_1722000_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1801 diff_1742400_1464000# diff_1004400_1458000# diff_1742400_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1802 diff_1762800_1464000# diff_1004400_1458000# diff_1762800_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1803 diff_1783200_1464000# diff_1004400_1458000# diff_1783200_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1804 diff_1803600_1464000# diff_1004400_1458000# diff_1803600_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1805 diff_1824000_1464000# diff_1004400_1458000# diff_1824000_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1806 diff_1844400_1464000# diff_1004400_1458000# diff_1844400_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1807 diff_1864800_1464000# diff_1004400_1458000# diff_1864800_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1808 diff_1885200_1464000# diff_1004400_1458000# diff_1885200_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1809 diff_1905600_1464000# diff_1004400_1458000# diff_1905600_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1810 diff_1926000_1464000# diff_1004400_1458000# diff_1926000_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1811 diff_1946400_1464000# diff_1004400_1458000# diff_1946400_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1812 diff_1966800_1464000# diff_1004400_1458000# diff_1966800_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1813 diff_1987200_1464000# diff_1004400_1458000# diff_1987200_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1814 diff_2007600_1464000# diff_1004400_1458000# diff_2007600_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1815 diff_2028000_1464000# diff_1004400_1458000# diff_2028000_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1816 diff_2048400_1464000# diff_1004400_1458000# diff_2048400_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1817 diff_2068800_1464000# diff_1004400_1458000# diff_2068800_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1818 diff_2089200_1464000# diff_1004400_1458000# diff_2089200_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1819 diff_2109600_1464000# diff_1004400_1458000# diff_2109600_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1820 diff_2130000_1464000# diff_1004400_1458000# diff_2130000_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1821 diff_2150400_1464000# diff_1004400_1458000# diff_2150400_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1822 diff_2170800_1464000# diff_1004400_1458000# diff_2170800_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1823 diff_2191200_1464000# diff_1004400_1458000# diff_2191200_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1824 diff_2211600_1464000# diff_1004400_1458000# diff_2211600_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1825 diff_2232000_1464000# diff_1004400_1458000# diff_2232000_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1826 diff_2252400_1464000# diff_1004400_1458000# diff_2252400_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1827 diff_2272800_1464000# diff_1004400_1458000# diff_2272800_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1828 diff_2293200_1464000# diff_1004400_1458000# diff_2293200_1441200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1829 Vdd Vdd diff_1004400_1435200# GND efet w=6000 l=13200
+ ad=0 pd=0 as=8.5104e+08 ps=259200 
M1830 diff_1008000_1441200# diff_1004400_1435200# diff_1008000_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1831 diff_1028400_1441200# diff_1004400_1435200# diff_1028400_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1832 diff_1048800_1441200# diff_1004400_1435200# diff_1048800_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1833 diff_1069200_1441200# diff_1004400_1435200# diff_1069200_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1834 diff_1089600_1441200# diff_1004400_1435200# diff_1089600_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1835 diff_1110000_1441200# diff_1004400_1435200# diff_1110000_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1836 diff_1130400_1441200# diff_1004400_1435200# diff_1130400_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1837 diff_1150800_1441200# diff_1004400_1435200# diff_1150800_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1838 diff_1171200_1441200# diff_1004400_1435200# diff_1171200_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1839 diff_1191600_1441200# diff_1004400_1435200# diff_1191600_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1840 diff_1212000_1441200# diff_1004400_1435200# diff_1212000_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1841 diff_1232400_1441200# diff_1004400_1435200# diff_1232400_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1842 diff_1252800_1441200# diff_1004400_1435200# diff_1252800_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1843 diff_1273200_1441200# diff_1004400_1435200# diff_1273200_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1844 diff_1293600_1441200# diff_1004400_1435200# diff_1293600_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1845 diff_1314000_1441200# diff_1004400_1435200# diff_1314000_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1846 diff_1334400_1441200# diff_1004400_1435200# diff_1334400_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1847 diff_1354800_1441200# diff_1004400_1435200# diff_1354800_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1848 diff_1375200_1441200# diff_1004400_1435200# diff_1375200_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1849 diff_1395600_1441200# diff_1004400_1435200# diff_1395600_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1850 diff_1416000_1441200# diff_1004400_1435200# diff_1416000_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1851 diff_1436400_1441200# diff_1004400_1435200# diff_1436400_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1852 diff_1456800_1441200# diff_1004400_1435200# diff_1456800_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1853 diff_1477200_1441200# diff_1004400_1435200# diff_1477200_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1854 diff_1497600_1441200# diff_1004400_1435200# diff_1497600_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1855 diff_1518000_1441200# diff_1004400_1435200# diff_1518000_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1856 diff_1538400_1441200# diff_1004400_1435200# diff_1538400_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1857 diff_1558800_1441200# diff_1004400_1435200# diff_1558800_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1858 diff_1579200_1441200# diff_1004400_1435200# diff_1579200_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1859 diff_1599600_1441200# diff_1004400_1435200# diff_1599600_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1860 diff_1620000_1441200# diff_1004400_1435200# diff_1620000_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1861 diff_1640400_1441200# diff_1004400_1435200# diff_1640400_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1862 diff_1660800_1441200# diff_1004400_1435200# diff_1660800_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1863 diff_1681200_1441200# diff_1004400_1435200# diff_1681200_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1864 diff_1701600_1441200# diff_1004400_1435200# diff_1701600_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1865 diff_1722000_1441200# diff_1004400_1435200# diff_1722000_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1866 diff_1742400_1441200# diff_1004400_1435200# diff_1742400_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1867 diff_1762800_1441200# diff_1004400_1435200# diff_1762800_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1868 diff_1783200_1441200# diff_1004400_1435200# diff_1783200_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1869 diff_1803600_1441200# diff_1004400_1435200# diff_1803600_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1870 diff_1824000_1441200# diff_1004400_1435200# diff_1824000_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1871 diff_1844400_1441200# diff_1004400_1435200# diff_1844400_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1872 diff_1864800_1441200# diff_1004400_1435200# diff_1864800_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1873 diff_1885200_1441200# diff_1004400_1435200# diff_1885200_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1874 diff_1905600_1441200# diff_1004400_1435200# diff_1905600_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1875 diff_1926000_1441200# diff_1004400_1435200# diff_1926000_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1876 diff_1946400_1441200# diff_1004400_1435200# diff_1946400_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1877 diff_1966800_1441200# diff_1004400_1435200# diff_1966800_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1878 diff_1987200_1441200# diff_1004400_1435200# diff_1987200_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1879 diff_2007600_1441200# diff_1004400_1435200# diff_2007600_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1880 diff_2028000_1441200# diff_1004400_1435200# diff_2028000_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1881 diff_2048400_1441200# diff_1004400_1435200# diff_2048400_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1882 diff_2068800_1441200# diff_1004400_1435200# diff_2068800_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1883 diff_2089200_1441200# diff_1004400_1435200# diff_2089200_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1884 diff_2109600_1441200# diff_1004400_1435200# diff_2109600_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1885 diff_2130000_1441200# diff_1004400_1435200# diff_2130000_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1886 diff_2150400_1441200# diff_1004400_1435200# diff_2150400_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1887 diff_2170800_1441200# diff_1004400_1435200# diff_2170800_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1888 diff_2191200_1441200# diff_1004400_1435200# diff_2191200_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1889 diff_2211600_1441200# diff_1004400_1435200# diff_2211600_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1890 diff_2232000_1441200# diff_1004400_1435200# diff_2232000_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1891 diff_2252400_1441200# diff_1004400_1435200# diff_2252400_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1892 diff_2272800_1441200# diff_1004400_1435200# diff_2272800_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1893 diff_2293200_1441200# diff_1004400_1435200# diff_2293200_1419600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1894 diff_804000_1662000# diff_189600_804000# GND GND efet w=190800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M1895 diff_1004400_1435200# diff_2384400_427200# diff_2367600_1494000# GND efet w=74400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M1896 diff_2367600_1494000# diff_2413200_996000# diff_1004400_1479600# GND efet w=84000 l=6000
+ ad=0 pd=0 as=1.15488e+09 ps=228000 
M1897 diff_1004400_1479600# Vdd Vdd GND efet w=7200 l=10800
+ ad=0 pd=0 as=0 ps=0 
M1898 Vdd Vdd diff_1004400_1458000# GND efet w=7200 l=12000
+ ad=0 pd=0 as=9.4176e+08 ps=247200 
M1899 diff_1008000_1419600# diff_1004400_1413600# diff_1008000_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1900 diff_1028400_1419600# diff_1004400_1413600# diff_1028400_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1901 diff_1048800_1419600# diff_1004400_1413600# diff_1048800_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1902 diff_1069200_1419600# diff_1004400_1413600# diff_1069200_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1903 diff_1089600_1419600# diff_1004400_1413600# diff_1089600_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1904 diff_1110000_1419600# diff_1004400_1413600# diff_1110000_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1905 diff_1130400_1419600# diff_1004400_1413600# diff_1130400_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1906 diff_1150800_1419600# diff_1004400_1413600# diff_1150800_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1907 diff_1171200_1419600# diff_1004400_1413600# diff_1171200_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1908 diff_1191600_1419600# diff_1004400_1413600# diff_1191600_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1909 diff_1212000_1419600# diff_1004400_1413600# diff_1212000_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1910 diff_1232400_1419600# diff_1004400_1413600# diff_1232400_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1911 diff_1252800_1419600# diff_1004400_1413600# diff_1252800_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1912 diff_1273200_1419600# diff_1004400_1413600# diff_1273200_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1913 diff_1293600_1419600# diff_1004400_1413600# diff_1293600_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1914 diff_1314000_1419600# diff_1004400_1413600# diff_1314000_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1915 diff_1334400_1419600# diff_1004400_1413600# diff_1334400_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1916 diff_1354800_1419600# diff_1004400_1413600# diff_1354800_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1917 diff_1375200_1419600# diff_1004400_1413600# diff_1375200_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1918 diff_1395600_1419600# diff_1004400_1413600# diff_1395600_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1919 diff_1416000_1419600# diff_1004400_1413600# diff_1416000_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1920 diff_1436400_1419600# diff_1004400_1413600# diff_1436400_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1921 diff_1456800_1419600# diff_1004400_1413600# diff_1456800_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1922 diff_1477200_1419600# diff_1004400_1413600# diff_1477200_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1923 diff_1497600_1419600# diff_1004400_1413600# diff_1497600_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1924 diff_1518000_1419600# diff_1004400_1413600# diff_1518000_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1925 diff_1538400_1419600# diff_1004400_1413600# diff_1538400_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1926 diff_1558800_1419600# diff_1004400_1413600# diff_1558800_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1927 diff_1579200_1419600# diff_1004400_1413600# diff_1579200_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1928 diff_1599600_1419600# diff_1004400_1413600# diff_1599600_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1929 diff_1620000_1419600# diff_1004400_1413600# diff_1620000_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1930 diff_1640400_1419600# diff_1004400_1413600# diff_1640400_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1931 diff_1660800_1419600# diff_1004400_1413600# diff_1660800_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1932 diff_1681200_1419600# diff_1004400_1413600# diff_1681200_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1933 diff_1701600_1419600# diff_1004400_1413600# diff_1701600_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1934 diff_1722000_1419600# diff_1004400_1413600# diff_1722000_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1935 diff_1742400_1419600# diff_1004400_1413600# diff_1742400_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1936 diff_1762800_1419600# diff_1004400_1413600# diff_1762800_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1937 diff_1783200_1419600# diff_1004400_1413600# diff_1783200_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1938 diff_1803600_1419600# diff_1004400_1413600# diff_1803600_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1939 diff_1824000_1419600# diff_1004400_1413600# diff_1824000_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1940 diff_1844400_1419600# diff_1004400_1413600# diff_1844400_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1941 diff_1864800_1419600# diff_1004400_1413600# diff_1864800_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1942 diff_1885200_1419600# diff_1004400_1413600# diff_1885200_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1943 diff_1905600_1419600# diff_1004400_1413600# diff_1905600_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1944 diff_1926000_1419600# diff_1004400_1413600# diff_1926000_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1945 diff_1946400_1419600# diff_1004400_1413600# diff_1946400_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1946 diff_1966800_1419600# diff_1004400_1413600# diff_1966800_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1947 diff_1987200_1419600# diff_1004400_1413600# diff_1987200_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1948 diff_2007600_1419600# diff_1004400_1413600# diff_2007600_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1949 diff_2028000_1419600# diff_1004400_1413600# diff_2028000_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1950 diff_2048400_1419600# diff_1004400_1413600# diff_2048400_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1951 diff_2068800_1419600# diff_1004400_1413600# diff_2068800_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1952 diff_2089200_1419600# diff_1004400_1413600# diff_2089200_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1953 diff_2109600_1419600# diff_1004400_1413600# diff_2109600_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1954 diff_2130000_1419600# diff_1004400_1413600# diff_2130000_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1955 diff_2150400_1419600# diff_1004400_1413600# diff_2150400_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1956 diff_2170800_1419600# diff_1004400_1413600# diff_2170800_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1957 diff_2191200_1419600# diff_1004400_1413600# diff_2191200_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1958 diff_2211600_1419600# diff_1004400_1413600# diff_2211600_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1959 diff_2232000_1419600# diff_1004400_1413600# diff_2232000_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1960 diff_2252400_1419600# diff_1004400_1413600# diff_2252400_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1961 diff_2272800_1419600# diff_1004400_1413600# diff_2272800_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1962 diff_2293200_1419600# diff_1004400_1413600# diff_2293200_1396800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M1963 diff_2367600_1407600# diff_2361600_427200# diff_1004400_1413600# GND efet w=86400 l=6000
+ ad=-4.68887e+08 pd=729600 as=9.6768e+08 ps=230400 
M1964 diff_1004400_1458000# diff_2431200_979200# diff_2367600_1494000# GND efet w=79200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M1965 diff_1008000_1396800# diff_1004400_1390800# diff_1008000_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1966 diff_1028400_1396800# diff_1004400_1390800# diff_1028400_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1967 diff_1048800_1396800# diff_1004400_1390800# diff_1048800_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1968 diff_1069200_1396800# diff_1004400_1390800# diff_1069200_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1969 diff_1089600_1396800# diff_1004400_1390800# diff_1089600_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1970 diff_1110000_1396800# diff_1004400_1390800# diff_1110000_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1971 diff_1130400_1396800# diff_1004400_1390800# diff_1130400_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1972 diff_1150800_1396800# diff_1004400_1390800# diff_1150800_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1973 diff_1171200_1396800# diff_1004400_1390800# diff_1171200_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1974 diff_1191600_1396800# diff_1004400_1390800# diff_1191600_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1975 diff_1212000_1396800# diff_1004400_1390800# diff_1212000_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1976 diff_1232400_1396800# diff_1004400_1390800# diff_1232400_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1977 diff_1252800_1396800# diff_1004400_1390800# diff_1252800_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1978 diff_1273200_1396800# diff_1004400_1390800# diff_1273200_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1979 diff_1293600_1396800# diff_1004400_1390800# diff_1293600_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1980 diff_1314000_1396800# diff_1004400_1390800# diff_1314000_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1981 diff_1334400_1396800# diff_1004400_1390800# diff_1334400_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1982 diff_1354800_1396800# diff_1004400_1390800# diff_1354800_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1983 diff_1375200_1396800# diff_1004400_1390800# diff_1375200_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1984 diff_1395600_1396800# diff_1004400_1390800# diff_1395600_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1985 diff_1416000_1396800# diff_1004400_1390800# diff_1416000_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1986 diff_1436400_1396800# diff_1004400_1390800# diff_1436400_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1987 diff_1456800_1396800# diff_1004400_1390800# diff_1456800_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1988 diff_1477200_1396800# diff_1004400_1390800# diff_1477200_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1989 diff_1497600_1396800# diff_1004400_1390800# diff_1497600_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1990 diff_1518000_1396800# diff_1004400_1390800# diff_1518000_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1991 diff_1538400_1396800# diff_1004400_1390800# diff_1538400_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1992 diff_1558800_1396800# diff_1004400_1390800# diff_1558800_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1993 diff_1579200_1396800# diff_1004400_1390800# diff_1579200_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1994 diff_1599600_1396800# diff_1004400_1390800# diff_1599600_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1995 diff_1620000_1396800# diff_1004400_1390800# diff_1620000_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1996 diff_1640400_1396800# diff_1004400_1390800# diff_1640400_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1997 diff_1660800_1396800# diff_1004400_1390800# diff_1660800_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1998 diff_1681200_1396800# diff_1004400_1390800# diff_1681200_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M1999 diff_1701600_1396800# diff_1004400_1390800# diff_1701600_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2000 diff_1722000_1396800# diff_1004400_1390800# diff_1722000_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2001 diff_1742400_1396800# diff_1004400_1390800# diff_1742400_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2002 diff_1762800_1396800# diff_1004400_1390800# diff_1762800_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2003 diff_1783200_1396800# diff_1004400_1390800# diff_1783200_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2004 diff_1803600_1396800# diff_1004400_1390800# diff_1803600_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2005 diff_1824000_1396800# diff_1004400_1390800# diff_1824000_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2006 diff_1844400_1396800# diff_1004400_1390800# diff_1844400_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2007 diff_1864800_1396800# diff_1004400_1390800# diff_1864800_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2008 diff_1885200_1396800# diff_1004400_1390800# diff_1885200_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2009 diff_1905600_1396800# diff_1004400_1390800# diff_1905600_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2010 diff_1926000_1396800# diff_1004400_1390800# diff_1926000_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2011 diff_1946400_1396800# diff_1004400_1390800# diff_1946400_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2012 diff_1966800_1396800# diff_1004400_1390800# diff_1966800_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2013 diff_1987200_1396800# diff_1004400_1390800# diff_1987200_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2014 diff_2007600_1396800# diff_1004400_1390800# diff_2007600_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2015 diff_2028000_1396800# diff_1004400_1390800# diff_2028000_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2016 diff_2048400_1396800# diff_1004400_1390800# diff_2048400_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2017 diff_2068800_1396800# diff_1004400_1390800# diff_2068800_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2018 diff_2089200_1396800# diff_1004400_1390800# diff_2089200_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2019 diff_2109600_1396800# diff_1004400_1390800# diff_2109600_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2020 diff_2130000_1396800# diff_1004400_1390800# diff_2130000_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2021 diff_2150400_1396800# diff_1004400_1390800# diff_2150400_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2022 diff_2170800_1396800# diff_1004400_1390800# diff_2170800_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2023 diff_2191200_1396800# diff_1004400_1390800# diff_2191200_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2024 diff_2211600_1396800# diff_1004400_1390800# diff_2211600_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2025 diff_2232000_1396800# diff_1004400_1390800# diff_2232000_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2026 diff_2252400_1396800# diff_1004400_1390800# diff_2252400_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2027 diff_2272800_1396800# diff_1004400_1390800# diff_2272800_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2028 diff_2293200_1396800# diff_1004400_1390800# diff_2293200_1375200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2029 diff_1004400_1413600# Vdd Vdd GND efet w=6000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M2030 diff_1008000_1375200# diff_1004400_1369200# diff_1008000_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2031 diff_1028400_1375200# diff_1004400_1369200# diff_1028400_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2032 diff_1048800_1375200# diff_1004400_1369200# diff_1048800_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2033 diff_1069200_1375200# diff_1004400_1369200# diff_1069200_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2034 diff_1089600_1375200# diff_1004400_1369200# diff_1089600_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2035 diff_1110000_1375200# diff_1004400_1369200# diff_1110000_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2036 diff_1130400_1375200# diff_1004400_1369200# diff_1130400_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2037 diff_1150800_1375200# diff_1004400_1369200# diff_1150800_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2038 diff_1171200_1375200# diff_1004400_1369200# diff_1171200_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2039 diff_1191600_1375200# diff_1004400_1369200# diff_1191600_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2040 diff_1212000_1375200# diff_1004400_1369200# diff_1212000_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2041 diff_1232400_1375200# diff_1004400_1369200# diff_1232400_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2042 diff_1252800_1375200# diff_1004400_1369200# diff_1252800_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2043 diff_1273200_1375200# diff_1004400_1369200# diff_1273200_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2044 diff_1293600_1375200# diff_1004400_1369200# diff_1293600_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2045 diff_1314000_1375200# diff_1004400_1369200# diff_1314000_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2046 diff_1334400_1375200# diff_1004400_1369200# diff_1334400_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2047 diff_1354800_1375200# diff_1004400_1369200# diff_1354800_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2048 diff_1375200_1375200# diff_1004400_1369200# diff_1375200_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2049 diff_1395600_1375200# diff_1004400_1369200# diff_1395600_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2050 diff_1416000_1375200# diff_1004400_1369200# diff_1416000_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2051 diff_1436400_1375200# diff_1004400_1369200# diff_1436400_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2052 diff_1456800_1375200# diff_1004400_1369200# diff_1456800_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2053 diff_1477200_1375200# diff_1004400_1369200# diff_1477200_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2054 diff_1497600_1375200# diff_1004400_1369200# diff_1497600_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2055 diff_1518000_1375200# diff_1004400_1369200# diff_1518000_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2056 diff_1538400_1375200# diff_1004400_1369200# diff_1538400_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2057 diff_1558800_1375200# diff_1004400_1369200# diff_1558800_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2058 diff_1579200_1375200# diff_1004400_1369200# diff_1579200_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2059 diff_1599600_1375200# diff_1004400_1369200# diff_1599600_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2060 diff_1620000_1375200# diff_1004400_1369200# diff_1620000_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2061 diff_1640400_1375200# diff_1004400_1369200# diff_1640400_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2062 diff_1660800_1375200# diff_1004400_1369200# diff_1660800_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2063 diff_1681200_1375200# diff_1004400_1369200# diff_1681200_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2064 diff_1701600_1375200# diff_1004400_1369200# diff_1701600_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2065 diff_1722000_1375200# diff_1004400_1369200# diff_1722000_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2066 diff_1742400_1375200# diff_1004400_1369200# diff_1742400_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2067 diff_1762800_1375200# diff_1004400_1369200# diff_1762800_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2068 diff_1783200_1375200# diff_1004400_1369200# diff_1783200_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2069 diff_1803600_1375200# diff_1004400_1369200# diff_1803600_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2070 diff_1824000_1375200# diff_1004400_1369200# diff_1824000_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2071 diff_1844400_1375200# diff_1004400_1369200# diff_1844400_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2072 diff_1864800_1375200# diff_1004400_1369200# diff_1864800_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2073 diff_1885200_1375200# diff_1004400_1369200# diff_1885200_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2074 diff_1905600_1375200# diff_1004400_1369200# diff_1905600_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2075 diff_1926000_1375200# diff_1004400_1369200# diff_1926000_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2076 diff_1946400_1375200# diff_1004400_1369200# diff_1946400_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2077 diff_1966800_1375200# diff_1004400_1369200# diff_1966800_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2078 diff_1987200_1375200# diff_1004400_1369200# diff_1987200_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2079 diff_2007600_1375200# diff_1004400_1369200# diff_2007600_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2080 diff_2028000_1375200# diff_1004400_1369200# diff_2028000_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2081 diff_2048400_1375200# diff_1004400_1369200# diff_2048400_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2082 diff_2068800_1375200# diff_1004400_1369200# diff_2068800_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2083 diff_2089200_1375200# diff_1004400_1369200# diff_2089200_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2084 diff_2109600_1375200# diff_1004400_1369200# diff_2109600_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2085 diff_2130000_1375200# diff_1004400_1369200# diff_2130000_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2086 diff_2150400_1375200# diff_1004400_1369200# diff_2150400_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2087 diff_2170800_1375200# diff_1004400_1369200# diff_2170800_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2088 diff_2191200_1375200# diff_1004400_1369200# diff_2191200_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2089 diff_2211600_1375200# diff_1004400_1369200# diff_2211600_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2090 diff_2232000_1375200# diff_1004400_1369200# diff_2232000_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2091 diff_2252400_1375200# diff_1004400_1369200# diff_2252400_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2092 diff_2272800_1375200# diff_1004400_1369200# diff_2272800_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2093 diff_2293200_1375200# diff_1004400_1369200# diff_2293200_1352400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2094 d3 clk2 diff_333600_1346400# GND efet w=12000 l=7200
+ ad=0 pd=0 as=1.008e+08 ps=40800 
M2095 d2 clk2 diff_488400_1346400# GND efet w=12000 l=7200
+ ad=0 pd=0 as=1.008e+08 ps=40800 
M2096 d1 clk2 diff_644400_1346400# GND efet w=12000 l=7200
+ ad=0 pd=0 as=1.008e+08 ps=40800 
M2097 d0 clk2 diff_799200_1346400# GND efet w=12000 l=7200
+ ad=0 pd=0 as=1.008e+08 ps=40800 
M2098 Vdd Vdd diff_1004400_1346400# GND efet w=6000 l=13200
+ ad=0 pd=0 as=8.5104e+08 ps=259200 
M2099 diff_333600_1346400# diff_154800_822000# diff_333600_1278000# GND efet w=12000 l=7200
+ ad=0 pd=0 as=1.64736e+09 ps=355200 
M2100 diff_488400_1346400# diff_154800_822000# diff_488400_1276800# GND efet w=12000 l=7200
+ ad=0 pd=0 as=1.61136e+09 ps=352800 
M2101 diff_644400_1346400# diff_154800_822000# diff_644400_1276800# GND efet w=12000 l=7200
+ ad=0 pd=0 as=1.66896e+09 ps=352800 
M2102 diff_799200_1346400# diff_154800_822000# diff_799200_1276800# GND efet w=12000 l=7200
+ ad=0 pd=0 as=1.65888e+09 ps=357600 
M2103 diff_1008000_1352400# diff_1004400_1346400# diff_1008000_1320000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2104 diff_1028400_1352400# diff_1004400_1346400# diff_1024800_1263600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2105 diff_1048800_1352400# diff_1004400_1346400# diff_1048800_1322400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2106 diff_1069200_1352400# diff_1004400_1346400# diff_1069200_1281600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2107 diff_1089600_1352400# diff_1004400_1346400# diff_1089600_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2108 diff_1110000_1352400# diff_1004400_1346400# diff_1110000_1262400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2109 diff_1130400_1352400# diff_1004400_1346400# diff_1130400_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2110 diff_1150800_1352400# diff_1004400_1346400# diff_1150800_1281600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2111 diff_1171200_1352400# diff_1004400_1346400# diff_1171200_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2112 diff_1191600_1352400# diff_1004400_1346400# diff_1191600_1262400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2113 diff_1212000_1352400# diff_1004400_1346400# diff_1212000_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2114 diff_1232400_1352400# diff_1004400_1346400# diff_1232400_1281600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2115 diff_1252800_1352400# diff_1004400_1346400# diff_1252800_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2116 diff_1273200_1352400# diff_1004400_1346400# diff_1273200_1262400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2117 diff_1293600_1352400# diff_1004400_1346400# diff_1293600_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2118 diff_1314000_1352400# diff_1004400_1346400# diff_1314000_1281600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2119 diff_1334400_1352400# diff_1004400_1346400# diff_1334400_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2120 diff_1354800_1352400# diff_1004400_1346400# diff_1354800_1262400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2121 diff_1375200_1352400# diff_1004400_1346400# diff_1375200_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2122 diff_1395600_1352400# diff_1004400_1346400# diff_1395600_1281600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2123 diff_1416000_1352400# diff_1004400_1346400# diff_1416000_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2124 diff_1436400_1352400# diff_1004400_1346400# diff_1436400_1262400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2125 diff_1456800_1352400# diff_1004400_1346400# diff_1456800_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2126 diff_1477200_1352400# diff_1004400_1346400# diff_1477200_1281600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2127 diff_1497600_1352400# diff_1004400_1346400# diff_1497600_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2128 diff_1518000_1352400# diff_1004400_1346400# diff_1518000_1262400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2129 diff_1538400_1352400# diff_1004400_1346400# diff_1538400_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2130 diff_1558800_1352400# diff_1004400_1346400# diff_1558800_1281600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2131 diff_1579200_1352400# diff_1004400_1346400# diff_1579200_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2132 diff_1599600_1352400# diff_1004400_1346400# diff_1599600_1262400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2133 diff_1620000_1352400# diff_1004400_1346400# diff_1620000_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2134 diff_1640400_1352400# diff_1004400_1346400# diff_1640400_1281600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2135 diff_1660800_1352400# diff_1004400_1346400# diff_1660800_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2136 diff_1681200_1352400# diff_1004400_1346400# diff_1681200_1262400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2137 diff_1701600_1352400# diff_1004400_1346400# diff_1701600_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2138 diff_1722000_1352400# diff_1004400_1346400# diff_1722000_1281600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2139 diff_1742400_1352400# diff_1004400_1346400# diff_1742400_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2140 diff_1762800_1352400# diff_1004400_1346400# diff_1762800_1262400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2141 diff_1783200_1352400# diff_1004400_1346400# diff_1783200_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2142 diff_1803600_1352400# diff_1004400_1346400# diff_1803600_1281600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2143 diff_1824000_1352400# diff_1004400_1346400# diff_1824000_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2144 diff_1844400_1352400# diff_1004400_1346400# diff_1844400_1262400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2145 diff_1864800_1352400# diff_1004400_1346400# diff_1864800_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2146 diff_1885200_1352400# diff_1004400_1346400# diff_1885200_1281600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2147 diff_1905600_1352400# diff_1004400_1346400# diff_1905600_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2148 diff_1926000_1352400# diff_1004400_1346400# diff_1926000_1262400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2149 diff_1946400_1352400# diff_1004400_1346400# diff_1946400_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2150 diff_1966800_1352400# diff_1004400_1346400# diff_1966800_1281600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2151 diff_1987200_1352400# diff_1004400_1346400# diff_1987200_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2152 diff_2007600_1352400# diff_1004400_1346400# diff_2007600_1262400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2153 diff_2028000_1352400# diff_1004400_1346400# diff_2028000_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2154 diff_2048400_1352400# diff_1004400_1346400# diff_2048400_1281600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2155 diff_2068800_1352400# diff_1004400_1346400# diff_2068800_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2156 diff_2089200_1352400# diff_1004400_1346400# diff_2089200_1262400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2157 diff_2109600_1352400# diff_1004400_1346400# diff_2109600_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2158 diff_2130000_1352400# diff_1004400_1346400# diff_2130000_1281600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2159 diff_2150400_1352400# diff_1004400_1346400# diff_2150400_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2160 diff_2170800_1352400# diff_1004400_1346400# diff_2170800_1262400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2161 diff_2191200_1352400# diff_1004400_1346400# diff_2191200_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2162 diff_2211600_1352400# diff_1004400_1346400# diff_2211600_1281600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2163 diff_2232000_1352400# diff_1004400_1346400# diff_2232000_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2164 diff_2252400_1352400# diff_1004400_1346400# diff_2252400_1262400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2165 diff_2272800_1352400# diff_1004400_1346400# diff_2272800_1321200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2166 diff_2293200_1352400# diff_1004400_1346400# diff_2293200_1281600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.2672e+08 ps=45600 
M2167 diff_280800_1316400# diff_154800_822000# GND GND efet w=18000 l=7200
+ ad=2.5776e+08 pd=72000 as=0 ps=0 
M2168 diff_333600_1278000# diff_333600_1278000# diff_333600_1278000# GND efet w=3600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2169 Vdd Vdd diff_280800_1316400# GND efet w=4200 l=41400
+ ad=0 pd=0 as=0 ps=0 
M2170 GND GND sync GND efet w=115800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2171 diff_336000_1170000# diff_333600_1278000# GND GND efet w=76800 l=7200
+ ad=7.5168e+08 pd=220800 as=0 ps=0 
M2172 diff_488400_1276800# diff_488400_1276800# diff_488400_1276800# GND efet w=3600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2173 diff_333600_1278000# diff_333600_1278000# diff_333600_1278000# GND efet w=2400 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2174 GND diff_336000_1170000# diff_355200_1299600# GND efet w=50400 l=6000
+ ad=0 pd=0 as=1.3752e+09 ps=345600 
M2175 diff_355200_1299600# diff_280800_1316400# diff_333600_1278000# GND efet w=12000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2176 diff_492000_1170000# diff_488400_1276800# GND GND efet w=76800 l=7200
+ ad=7.4448e+08 pd=220800 as=0 ps=0 
M2177 diff_644400_1276800# diff_644400_1276800# diff_644400_1276800# GND efet w=2400 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2178 diff_488400_1276800# diff_488400_1276800# diff_488400_1276800# GND efet w=2400 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2179 GND diff_492000_1170000# diff_508800_1299600# GND efet w=50400 l=6000
+ ad=0 pd=0 as=1.37664e+09 ps=343200 
M2180 diff_508800_1299600# diff_280800_1316400# diff_488400_1276800# GND efet w=12000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2181 diff_646800_1170000# diff_644400_1276800# GND GND efet w=75600 l=7200
+ ad=7.9488e+08 pd=218400 as=0 ps=0 
M2182 diff_1004400_1346400# diff_2384400_427200# diff_2367600_1407600# GND efet w=74400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2183 diff_2367600_1407600# diff_2413200_996000# diff_1004400_1390800# GND efet w=85200 l=6000
+ ad=0 pd=0 as=1.14768e+09 ps=228000 
M2184 diff_1004400_1390800# Vdd Vdd GND efet w=7200 l=10800
+ ad=0 pd=0 as=0 ps=0 
M2185 Vdd Vdd diff_1004400_1369200# GND efet w=7200 l=13200
+ ad=0 pd=0 as=9.4176e+08 ps=247200 
M2186 diff_799200_1276800# diff_799200_1276800# diff_799200_1276800# GND efet w=3600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2187 diff_644400_1276800# diff_644400_1276800# diff_644400_1276800# GND efet w=1200 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2188 GND diff_646800_1170000# diff_666000_1299600# GND efet w=50400 l=7200
+ ad=0 pd=0 as=1.34208e+09 ps=340800 
M2189 diff_666000_1299600# diff_280800_1316400# diff_644400_1276800# GND efet w=12000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2190 diff_801600_1170000# diff_799200_1276800# GND GND efet w=76800 l=7200
+ ad=7.4448e+08 pd=218400 as=0 ps=0 
M2191 diff_799200_1276800# diff_799200_1276800# diff_799200_1276800# GND efet w=2400 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2192 GND diff_801600_1170000# diff_820800_1299600# GND efet w=50400 l=6000
+ ad=0 pd=0 as=1.368e+09 ps=343200 
M2193 diff_820800_1299600# diff_280800_1316400# diff_799200_1276800# GND efet w=12000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2194 diff_333600_1278000# cl GND GND efet w=36000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2195 GND cl diff_333600_1278000# GND efet w=36000 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2196 diff_333600_1278000# diff_260400_786000# GND GND efet w=47400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2197 diff_336000_1170000# Vdd Vdd GND efet w=6000 l=15600
+ ad=0 pd=0 as=0 ps=0 
M2198 diff_355200_1299600# Vdd Vdd GND efet w=6000 l=14400
+ ad=0 pd=0 as=0 ps=0 
M2199 Vdd Vdd Vdd GND efet w=2400 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2200 Vdd Vdd Vdd GND efet w=1800 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2201 diff_488400_1276800# cl GND GND efet w=36000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2202 GND cl diff_488400_1276800# GND efet w=36000 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2203 GND diff_1008000_1320000# diff_997200_1236000# GND efet w=28800 l=6000
+ ad=0 pd=0 as=7.92e+08 ps=194400 
M2204 diff_1033200_1267200# diff_1024800_1263600# GND GND efet w=46200 l=7200
+ ad=3.6864e+08 pd=105600 as=0 ps=0 
M2205 GND diff_1048800_1322400# diff_1036800_1202400# GND efet w=39600 l=6000
+ ad=0 pd=0 as=7.5456e+08 ps=192000 
M2206 diff_1075200_1284000# diff_1069200_1281600# GND GND efet w=39600 l=6000
+ ad=6.408e+08 pd=187200 as=0 ps=0 
M2207 GND diff_1089600_1321200# diff_1074000_1180800# GND efet w=35400 l=7200
+ ad=0 pd=0 as=6.6816e+08 ps=175200 
M2208 GND diff_1130400_1321200# diff_1116000_1201200# GND efet w=39600 l=6000
+ ad=0 pd=0 as=7.5888e+08 ps=196800 
M2209 diff_1156800_1284000# diff_1150800_1281600# GND GND efet w=39600 l=6000
+ ad=6.6096e+08 pd=187200 as=0 ps=0 
M2210 diff_1116000_1266000# diff_1110000_1262400# GND GND efet w=35400 l=6600
+ ad=3.2976e+08 pd=93600 as=0 ps=0 
M2211 GND diff_1171200_1321200# diff_1155600_1180800# GND efet w=35400 l=7200
+ ad=0 pd=0 as=6.7392e+08 ps=175200 
M2212 GND diff_1212000_1321200# diff_1197600_1202400# GND efet w=39600 l=6000
+ ad=0 pd=0 as=7.7616e+08 ps=196800 
M2213 diff_1238400_1284000# diff_1232400_1281600# GND GND efet w=39600 l=6000
+ ad=6.552e+08 pd=187200 as=0 ps=0 
M2214 diff_1197600_1266000# diff_1191600_1262400# GND GND efet w=35400 l=6600
+ ad=3.2976e+08 pd=93600 as=0 ps=0 
M2215 GND diff_1252800_1321200# diff_1236000_1180800# GND efet w=35400 l=7200
+ ad=0 pd=0 as=7.056e+08 ps=177600 
M2216 GND diff_1293600_1321200# diff_1278000_1202400# GND efet w=39600 l=6000
+ ad=0 pd=0 as=7.9488e+08 ps=196800 
M2217 diff_1320000_1284000# diff_1314000_1281600# GND GND efet w=39600 l=6000
+ ad=6.8688e+08 pd=189600 as=0 ps=0 
M2218 diff_1279200_1266000# diff_1273200_1262400# GND GND efet w=35400 l=6600
+ ad=3.2976e+08 pd=93600 as=0 ps=0 
M2219 GND diff_1334400_1321200# diff_1317600_1180800# GND efet w=35400 l=7200
+ ad=0 pd=0 as=7.1136e+08 ps=177600 
M2220 GND diff_1375200_1321200# diff_1359600_1201200# GND efet w=39600 l=6000
+ ad=0 pd=0 as=8.1504e+08 ps=201600 
M2221 diff_1401600_1284000# diff_1395600_1281600# GND GND efet w=39600 l=6000
+ ad=5.9616e+08 pd=184800 as=0 ps=0 
M2222 diff_1360800_1266000# diff_1354800_1262400# GND GND efet w=35400 l=6600
+ ad=3.2976e+08 pd=93600 as=0 ps=0 
M2223 GND diff_1416000_1321200# diff_1400400_1180800# GND efet w=35400 l=7200
+ ad=0 pd=0 as=6.3072e+08 ps=172800 
M2224 GND diff_1456800_1321200# diff_1442400_1202400# GND efet w=39600 l=6000
+ ad=0 pd=0 as=7.2e+08 ps=192000 
M2225 diff_1483200_1284000# diff_1477200_1281600# GND GND efet w=39600 l=6000
+ ad=6.2064e+08 pd=184800 as=0 ps=0 
M2226 diff_1442400_1266000# diff_1436400_1262400# GND GND efet w=35400 l=6600
+ ad=3.2976e+08 pd=93600 as=0 ps=0 
M2227 GND diff_1497600_1321200# diff_1482000_1180800# GND efet w=35400 l=7200
+ ad=0 pd=0 as=6.3648e+08 ps=172800 
M2228 GND diff_1538400_1321200# diff_1524000_1202400# GND efet w=39600 l=6000
+ ad=0 pd=0 as=7.3872e+08 ps=194400 
M2229 diff_1564800_1284000# diff_1558800_1281600# GND GND efet w=39600 l=6000
+ ad=5.9616e+08 pd=184800 as=0 ps=0 
M2230 diff_1524000_1266000# diff_1518000_1262400# GND GND efet w=35400 l=6600
+ ad=3.2976e+08 pd=93600 as=0 ps=0 
M2231 GND diff_1579200_1321200# diff_1563600_1180800# GND efet w=35400 l=7200
+ ad=0 pd=0 as=6.3072e+08 ps=172800 
M2232 GND diff_1620000_1321200# diff_1605600_1202400# GND efet w=39600 l=6000
+ ad=0 pd=0 as=7.2e+08 ps=192000 
M2233 diff_1646400_1284000# diff_1640400_1281600# GND GND efet w=39600 l=6000
+ ad=6.2496e+08 pd=184800 as=0 ps=0 
M2234 diff_1605600_1266000# diff_1599600_1262400# GND GND efet w=35400 l=6600
+ ad=3.2976e+08 pd=93600 as=0 ps=0 
M2235 GND diff_1660800_1321200# diff_1645200_1180800# GND efet w=35400 l=7200
+ ad=0 pd=0 as=6.3648e+08 ps=172800 
M2236 GND diff_1701600_1321200# diff_1687200_1202400# GND efet w=39600 l=6000
+ ad=0 pd=0 as=7.3872e+08 ps=194400 
M2237 diff_1728000_1284000# diff_1722000_1281600# GND GND efet w=39600 l=6000
+ ad=6.3648e+08 pd=187200 as=0 ps=0 
M2238 diff_1687200_1266000# diff_1681200_1262400# GND GND efet w=35400 l=6600
+ ad=3.2976e+08 pd=93600 as=0 ps=0 
M2239 GND diff_1742400_1321200# diff_1728000_1180800# GND efet w=35400 l=7200
+ ad=0 pd=0 as=6.6816e+08 ps=175200 
M2240 GND diff_1783200_1321200# diff_1770000_1202400# GND efet w=39600 l=6000
+ ad=0 pd=0 as=7.5744e+08 ps=194400 
M2241 diff_1809600_1284000# diff_1803600_1281600# GND GND efet w=39600 l=6000
+ ad=6.6384e+08 pd=187200 as=0 ps=0 
M2242 diff_1768800_1266000# diff_1762800_1262400# GND GND efet w=35400 l=6600
+ ad=3.2976e+08 pd=93600 as=0 ps=0 
M2243 GND diff_1824000_1321200# diff_1809600_1180800# GND efet w=35400 l=7200
+ ad=0 pd=0 as=6.7392e+08 ps=175200 
M2244 GND diff_1864800_1321200# diff_1851600_1202400# GND efet w=39600 l=6000
+ ad=0 pd=0 as=7.7616e+08 ps=196800 
M2245 diff_1891200_1284000# diff_1885200_1281600# GND GND efet w=39600 l=6000
+ ad=6.3504e+08 pd=187200 as=0 ps=0 
M2246 diff_1850400_1266000# diff_1844400_1262400# GND GND efet w=35400 l=6600
+ ad=3.2976e+08 pd=93600 as=0 ps=0 
M2247 GND diff_1905600_1321200# diff_1890000_1180800# GND efet w=35400 l=7200
+ ad=0 pd=0 as=6.6816e+08 ps=175200 
M2248 GND diff_1946400_1321200# diff_1932000_1202400# GND efet w=39600 l=6000
+ ad=0 pd=0 as=7.5744e+08 ps=194400 
M2249 diff_1972800_1284000# diff_1966800_1281600# GND GND efet w=39600 l=6000
+ ad=6.6096e+08 pd=187200 as=0 ps=0 
M2250 diff_1932000_1266000# diff_1926000_1262400# GND GND efet w=35400 l=6600
+ ad=3.2976e+08 pd=93600 as=0 ps=0 
M2251 GND diff_1987200_1321200# diff_1971600_1180800# GND efet w=35400 l=7200
+ ad=0 pd=0 as=6.7392e+08 ps=175200 
M2252 GND diff_2028000_1321200# diff_2013600_1202400# GND efet w=39600 l=6000
+ ad=0 pd=0 as=7.7616e+08 ps=196800 
M2253 diff_2054400_1284000# diff_2048400_1281600# GND GND efet w=39600 l=6000
+ ad=6.3504e+08 pd=187200 as=0 ps=0 
M2254 diff_2013600_1266000# diff_2007600_1262400# GND GND efet w=35400 l=6600
+ ad=3.2976e+08 pd=93600 as=0 ps=0 
M2255 GND diff_2068800_1321200# diff_2053200_1180800# GND efet w=35400 l=7200
+ ad=0 pd=0 as=6.6816e+08 ps=175200 
M2256 GND diff_2109600_1321200# diff_2095200_1202400# GND efet w=39600 l=6000
+ ad=0 pd=0 as=7.5744e+08 ps=194400 
M2257 diff_2136000_1284000# diff_2130000_1281600# GND GND efet w=39600 l=6000
+ ad=6.6096e+08 pd=187200 as=0 ps=0 
M2258 diff_2095200_1266000# diff_2089200_1262400# GND GND efet w=35400 l=6600
+ ad=3.2976e+08 pd=93600 as=0 ps=0 
M2259 GND diff_2150400_1321200# diff_2134800_1180800# GND efet w=35400 l=7200
+ ad=0 pd=0 as=6.7392e+08 ps=175200 
M2260 GND diff_2191200_1321200# diff_2176800_1202400# GND efet w=39600 l=6000
+ ad=0 pd=0 as=7.7616e+08 ps=196800 
M2261 diff_2217600_1284000# diff_2211600_1281600# GND GND efet w=39600 l=6000
+ ad=6.1776e+08 pd=182400 as=0 ps=0 
M2262 diff_2176800_1266000# diff_2170800_1262400# GND GND efet w=35400 l=6600
+ ad=3.2976e+08 pd=93600 as=0 ps=0 
M2263 GND diff_2232000_1321200# diff_2217600_1180800# GND efet w=35400 l=7200
+ ad=0 pd=0 as=6.5952e+08 ps=172800 
M2264 GND diff_2272800_1321200# diff_2259600_1202400# GND efet w=39600 l=6000
+ ad=0 pd=0 as=7.3584e+08 ps=192000 
M2265 diff_2299200_1284000# diff_2293200_1281600# GND GND efet w=39600 l=6000
+ ad=8.0352e+08 pd=249600 as=0 ps=0 
M2266 diff_2258400_1266000# diff_2252400_1262400# GND GND efet w=35400 l=6600
+ ad=3.2976e+08 pd=93600 as=0 ps=0 
M2267 diff_488400_1276800# diff_260400_786000# GND GND efet w=46200 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2268 diff_492000_1170000# Vdd Vdd GND efet w=6000 l=15600
+ ad=0 pd=0 as=0 ps=0 
M2269 diff_508800_1299600# Vdd Vdd GND efet w=6000 l=14400
+ ad=0 pd=0 as=0 ps=0 
M2270 Vdd Vdd Vdd GND efet w=2400 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2271 Vdd Vdd Vdd GND efet w=1200 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2272 diff_644400_1276800# cl GND GND efet w=36000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2273 GND cl diff_644400_1276800# GND efet w=36000 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2274 diff_644400_1276800# diff_260400_786000# GND GND efet w=48600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2275 diff_646800_1170000# Vdd Vdd GND efet w=6000 l=15600
+ ad=0 pd=0 as=0 ps=0 
M2276 diff_666000_1299600# Vdd Vdd GND efet w=6000 l=14400
+ ad=0 pd=0 as=0 ps=0 
M2277 Vdd Vdd Vdd GND efet w=1200 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2278 Vdd Vdd Vdd GND efet w=1200 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2279 diff_799200_1276800# cl GND GND efet w=36000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2280 GND cl diff_799200_1276800# GND efet w=36000 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2281 diff_799200_1276800# diff_260400_786000# GND GND efet w=48600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2282 diff_999600_1216800# diff_1048800_846000# diff_1033200_1267200# GND efet w=31200 l=7200
+ ad=2.03184e+09 pd=480000 as=0 ps=0 
M2283 diff_1077600_1207200# diff_1048800_846000# diff_1116000_1266000# GND efet w=30000 l=6000
+ ad=1.69056e+09 pd=408000 as=0 ps=0 
M2284 diff_1159200_1207200# diff_1048800_846000# diff_1197600_1266000# GND efet w=30000 l=6000
+ ad=1.7568e+09 pd=458400 as=0 ps=0 
M2285 diff_1239600_1208400# diff_1048800_846000# diff_1279200_1266000# GND efet w=30000 l=6000
+ ad=1.62e+09 pd=403200 as=0 ps=0 
M2286 diff_1321200_1208400# diff_1048800_846000# diff_1360800_1266000# GND efet w=30000 l=6000
+ ad=1.79712e+09 pd=468000 as=0 ps=0 
M2287 diff_1404000_1206000# diff_1048800_846000# diff_1442400_1266000# GND efet w=30000 l=6000
+ ad=1.74384e+09 pd=412800 as=0 ps=0 
M2288 diff_1485600_1206000# diff_1048800_846000# diff_1524000_1266000# GND efet w=30000 l=6000
+ ad=1.8576e+09 pd=470400 as=0 ps=0 
M2289 diff_1567200_1206000# diff_1048800_846000# diff_1605600_1266000# GND efet w=30000 l=6000
+ ad=1.74384e+09 pd=412800 as=0 ps=0 
M2290 diff_1648800_1206000# diff_1048800_846000# diff_1687200_1266000# GND efet w=30000 l=6000
+ ad=1.82016e+09 pd=463200 as=0 ps=0 
M2291 diff_1731600_1207200# diff_1048800_846000# diff_1768800_1266000# GND efet w=30000 l=6000
+ ad=1.69344e+09 pd=408000 as=0 ps=0 
M2292 diff_1813200_1207200# diff_1048800_846000# diff_1850400_1266000# GND efet w=30000 l=6000
+ ad=1.8e+09 pd=460800 as=0 ps=0 
M2293 diff_1893600_1207200# diff_1048800_846000# diff_1932000_1266000# GND efet w=30000 l=6000
+ ad=1.68768e+09 pd=408000 as=0 ps=0 
M2294 diff_1975200_1207200# diff_1048800_846000# diff_2013600_1266000# GND efet w=30000 l=6000
+ ad=1.8e+09 pd=463200 as=0 ps=0 
M2295 diff_2056800_1207200# diff_1048800_846000# diff_2095200_1266000# GND efet w=30000 l=6000
+ ad=1.68768e+09 pd=408000 as=0 ps=0 
M2296 diff_2138400_1207200# diff_1048800_846000# diff_2176800_1266000# GND efet w=30000 l=6000
+ ad=1.82304e+09 pd=465600 as=0 ps=0 
M2297 diff_2221200_1206000# diff_1048800_846000# diff_2258400_1266000# GND efet w=30000 l=6000
+ ad=1.77984e+09 pd=424800 as=0 ps=0 
M2298 diff_1004400_1369200# diff_2431200_979200# diff_2367600_1407600# GND efet w=79200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2299 diff_2437200_1698000# diff_2451600_979200# diff_2367600_1407600# GND efet w=154800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2300 diff_2367600_1494000# diff_2469600_912000# diff_2437200_1698000# GND efet w=154800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2301 diff_999600_1216800# diff_994800_1225200# diff_997200_1236000# GND efet w=40800 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2302 diff_801600_1170000# Vdd Vdd GND efet w=6000 l=15600
+ ad=0 pd=0 as=0 ps=0 
M2303 diff_820800_1299600# Vdd Vdd GND efet w=6000 l=14400
+ ad=0 pd=0 as=0 ps=0 
M2304 diff_1320000_1284000# diff_994800_1225200# diff_1321200_1208400# GND efet w=34200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2305 diff_1238400_1284000# diff_994800_1225200# diff_1239600_1208400# GND efet w=31200 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2306 diff_1401600_1284000# diff_994800_1225200# diff_1404000_1206000# GND efet w=31200 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2307 diff_1483200_1284000# diff_994800_1225200# diff_1485600_1206000# GND efet w=32400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2308 diff_1564800_1284000# diff_994800_1225200# diff_1567200_1206000# GND efet w=31200 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2309 diff_1075200_1284000# diff_994800_1225200# diff_1077600_1207200# GND efet w=30600 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2310 diff_1156800_1284000# diff_994800_1225200# diff_1159200_1207200# GND efet w=31200 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2311 diff_1646400_1284000# diff_994800_1225200# diff_1648800_1206000# GND efet w=31200 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2312 diff_1891200_1284000# diff_994800_1225200# diff_1893600_1207200# GND efet w=30600 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2313 diff_1972800_1284000# diff_994800_1225200# diff_1975200_1207200# GND efet w=31200 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2314 diff_2054400_1284000# diff_994800_1225200# diff_2056800_1207200# GND efet w=30600 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2315 diff_2136000_1284000# diff_994800_1225200# diff_2138400_1207200# GND efet w=31200 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2316 Vdd Vdd Vdd GND efet w=1200 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2317 Vdd Vdd Vdd GND efet w=1200 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2318 diff_1036800_1202400# diff_1033200_919200# diff_999600_1216800# GND efet w=28800 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2319 diff_1116000_1201200# diff_1033200_919200# diff_1077600_1207200# GND efet w=34200 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2320 diff_1197600_1202400# diff_1033200_919200# diff_1159200_1207200# GND efet w=33600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2321 diff_1278000_1202400# diff_1033200_919200# diff_1239600_1208400# GND efet w=33600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2322 diff_1359600_1201200# diff_1033200_919200# diff_1321200_1208400# GND efet w=34800 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2323 diff_1442400_1202400# diff_1033200_919200# diff_1404000_1206000# GND efet w=33600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2324 diff_1524000_1202400# diff_1033200_919200# diff_1485600_1206000# GND efet w=34200 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2325 diff_1728000_1284000# diff_994800_1225200# diff_1731600_1207200# GND efet w=30000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2326 diff_1809600_1284000# diff_994800_1225200# diff_1813200_1207200# GND efet w=30600 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2327 diff_1605600_1202400# diff_1033200_919200# diff_1567200_1206000# GND efet w=33600 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2328 diff_1687200_1202400# diff_1033200_919200# diff_1648800_1206000# GND efet w=33600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2329 diff_1770000_1202400# diff_1033200_919200# diff_1731600_1207200# GND efet w=33000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2330 diff_1851600_1202400# diff_1033200_919200# diff_1813200_1207200# GND efet w=33000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2331 diff_1932000_1202400# diff_1033200_919200# diff_1893600_1207200# GND efet w=33600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2332 diff_2013600_1202400# diff_1033200_919200# diff_1975200_1207200# GND efet w=33600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2333 diff_2217600_1284000# diff_994800_1225200# diff_2221200_1206000# GND efet w=28800 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2334 diff_2095200_1202400# diff_1033200_919200# diff_2056800_1207200# GND efet w=33600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2335 diff_2176800_1202400# diff_1033200_919200# diff_2138400_1207200# GND efet w=33600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2336 diff_2259600_1202400# diff_1033200_919200# diff_2221200_1206000# GND efet w=31800 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2337 GND diff_336000_1170000# diff_337200_1087200# GND efet w=56400 l=6000
+ ad=0 pd=0 as=1.11456e+09 ps=259200 
M2338 GND diff_492000_1170000# diff_493200_1087200# GND efet w=56400 l=6000
+ ad=0 pd=0 as=1.11744e+09 ps=254400 
M2339 Vdd Vdd diff_337200_1087200# GND efet w=7200 l=13200
+ ad=0 pd=0 as=0 ps=0 
M2340 GND diff_646800_1170000# diff_648000_1087200# GND efet w=56400 l=6000
+ ad=0 pd=0 as=1.17072e+09 ps=259200 
M2341 diff_337200_1087200# diff_337200_1087200# diff_337200_1087200# GND efet w=1800 l=1800
+ ad=0 pd=0 as=0 ps=0 
M2342 diff_337200_1087200# diff_337200_1087200# diff_337200_1087200# GND efet w=3600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2343 Vdd Vdd diff_493200_1087200# GND efet w=7200 l=10800
+ ad=0 pd=0 as=0 ps=0 
M2344 GND diff_801600_1170000# diff_802800_1087200# GND efet w=56400 l=6000
+ ad=0 pd=0 as=1.17216e+09 ps=266400 
M2345 diff_493200_1087200# diff_493200_1087200# diff_493200_1087200# GND efet w=3600 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2346 Vdd Vdd diff_648000_1087200# GND efet w=7200 l=10800
+ ad=0 pd=0 as=0 ps=0 
M2347 diff_1074000_1180800# diff_1063200_940800# diff_999600_1216800# GND efet w=31200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2348 diff_1155600_1180800# diff_1063200_940800# diff_1077600_1207200# GND efet w=31200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2349 diff_1236000_1180800# diff_1063200_940800# diff_1159200_1207200# GND efet w=31200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2350 diff_1317600_1180800# diff_1063200_940800# diff_1239600_1208400# GND efet w=31200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2351 diff_1400400_1180800# diff_1063200_940800# diff_1321200_1208400# GND efet w=31200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2352 diff_1482000_1180800# diff_1063200_940800# diff_1404000_1206000# GND efet w=31200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2353 diff_1563600_1180800# diff_1063200_940800# diff_1485600_1206000# GND efet w=31200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2354 diff_1645200_1180800# diff_1063200_940800# diff_1567200_1206000# GND efet w=31200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2355 diff_1728000_1180800# diff_1063200_940800# diff_1648800_1206000# GND efet w=31200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2356 diff_1809600_1180800# diff_1063200_940800# diff_1731600_1207200# GND efet w=31200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2357 diff_1890000_1180800# diff_1063200_940800# diff_1813200_1207200# GND efet w=31200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2358 diff_1971600_1180800# diff_1063200_940800# diff_1893600_1207200# GND efet w=31200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2359 diff_2053200_1180800# diff_1063200_940800# diff_1975200_1207200# GND efet w=31200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2360 diff_2134800_1180800# diff_1063200_940800# diff_2056800_1207200# GND efet w=31200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2361 diff_2217600_1180800# diff_1063200_940800# diff_2138400_1207200# GND efet w=30000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2362 diff_2299200_1284000# diff_1063200_940800# diff_2221200_1206000# GND efet w=46200 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2363 diff_648000_1087200# diff_648000_1087200# diff_648000_1087200# GND efet w=4800 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2364 diff_802800_1087200# diff_802800_1087200# diff_802800_1087200# GND efet w=2400 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2365 Vdd Vdd diff_802800_1087200# GND efet w=7200 l=10800
+ ad=0 pd=0 as=0 ps=0 
M2366 diff_802800_1087200# diff_802800_1087200# diff_802800_1087200# GND efet w=4200 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2367 diff_999600_1216800# diff_1011600_1153200# diff_1016400_968400# GND efet w=40800 l=7200
+ ad=0 pd=0 as=-7.52567e+08 ps=691200 
M2368 diff_1077600_1207200# diff_1124400_1153200# diff_1016400_968400# GND efet w=40800 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2369 diff_1239600_1208400# diff_1124400_1153200# diff_1180800_985200# GND efet w=40800 l=6000
+ ad=0 pd=0 as=-9.70007e+08 ps=655200 
M2370 diff_1404000_1206000# diff_1124400_1153200# diff_1342800_1122000# GND efet w=40800 l=6000
+ ad=0 pd=0 as=-5.68247e+08 ps=700800 
M2371 diff_1567200_1206000# diff_1124400_1153200# diff_1507200_984000# GND efet w=40800 l=6000
+ ad=0 pd=0 as=-5.27927e+08 ps=693600 
M2372 diff_1731600_1207200# diff_1124400_1153200# diff_1670400_984000# GND efet w=40800 l=6000
+ ad=0 pd=0 as=-8.36087e+08 ps=660000 
M2373 diff_1893600_1207200# diff_1124400_1153200# diff_1834800_984000# GND efet w=40800 l=6000
+ ad=0 pd=0 as=-9.09527e+08 ps=636000 
M2374 diff_2056800_1207200# diff_1124400_1153200# diff_1996800_984000# GND efet w=40800 l=6000
+ ad=0 pd=0 as=-5.42327e+08 ps=715200 
M2375 diff_2221200_1206000# diff_1124400_1153200# diff_2160000_985200# GND efet w=34800 l=6000
+ ad=0 pd=0 as=-1.33289e+09 ps=576000 
M2376 Vdd diff_337200_1087200# io3 GND efet w=176400 l=7200
+ ad=0 pd=0 as=1.43823e+09 ps=1.9392e+06 
M2377 d3 GND d3 GND efet w=177000 l=112200
+ ad=0 pd=0 as=0 ps=0 
M2378 GND diff_336000_1170000# io3 GND efet w=180600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2379 Vdd diff_493200_1087200# io2 GND efet w=177600 l=7200
+ ad=0 pd=0 as=9.42865e+08 ps=1.9272e+06 
M2380 io2 GND io2 GND efet w=175800 l=107400
+ ad=0 pd=0 as=0 ps=0 
M2381 GND diff_492000_1170000# io2 GND efet w=180600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2382 Vdd diff_648000_1087200# io1 GND efet w=177600 l=7200
+ ad=0 pd=0 as=6.01585e+08 ps=1.8528e+06 
M2383 GND diff_646800_1170000# io1 GND efet w=180600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2384 Vdd diff_802800_1087200# io0 GND efet w=176400 l=7200
+ ad=0 pd=0 as=9.25585e+08 ps=1.9368e+06 
M2385 diff_496800_967200# diff_406800_692400# diff_408000_1448400# GND efet w=22800 l=7200
+ ad=8.9424e+08 pd=230400 as=1.25136e+09 ps=326400 
M2386 diff_543600_1017600# diff_446400_902400# diff_496800_967200# GND efet w=22800 l=7200
+ ad=1.09008e+09 pd=244800 as=0 ps=0 
M2387 diff_648000_967200# diff_406800_692400# diff_562800_1448400# GND efet w=22800 l=7200
+ ad=9.6048e+08 pd=240000 as=1.00656e+09 ps=261600 
M2388 diff_682800_1034400# diff_446400_902400# diff_648000_967200# GND efet w=22800 l=7200
+ ad=1.02528e+09 pd=216000 as=0 ps=0 
M2389 io1 GND io1 GND efet w=167400 l=125400
+ ad=0 pd=0 as=0 ps=0 
M2390 io3 GND io3 GND efet w=149400 l=70200
+ ad=0 pd=0 as=0 ps=0 
M2391 diff_496800_967200# diff_411600_867600# io3 GND efet w=21600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2392 GND diff_801600_1170000# io0 GND efet w=180600 l=8400
+ ad=0 pd=0 as=0 ps=0 
M2393 diff_1159200_1207200# diff_1011600_1153200# diff_1180800_985200# GND efet w=39600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2394 diff_1321200_1208400# diff_1011600_1153200# diff_1342800_1122000# GND efet w=40800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2395 diff_1485600_1206000# diff_1011600_1153200# diff_1507200_984000# GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2396 diff_1648800_1206000# diff_1011600_1153200# diff_1670400_984000# GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2397 diff_1813200_1207200# diff_1011600_1153200# diff_1834800_984000# GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2398 diff_1975200_1207200# diff_1011600_1153200# diff_1996800_984000# GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2399 diff_2138400_1207200# diff_1011600_1153200# diff_2160000_985200# GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2400 diff_901200_968400# diff_406800_692400# diff_873600_1448400# GND efet w=21600 l=7200
+ ad=1.53504e+09 pd=403200 as=2.8224e+08 ps=69600 
M2401 diff_967200_1083600# diff_446400_902400# diff_901200_968400# GND efet w=21600 l=7200
+ ad=7.2432e+08 pd=160800 as=0 ps=0 
M2402 diff_802800_967200# diff_406800_692400# diff_718800_1448400# GND efet w=22800 l=7200
+ ad=1.0368e+09 pd=264000 as=8.8704e+08 ps=232800 
M2403 diff_829200_1039200# diff_446400_902400# diff_802800_967200# GND efet w=22800 l=7200
+ ad=1.6344e+09 pd=343200 as=0 ps=0 
M2404 io0 GND io0 GND efet w=177600 l=129600
+ ad=0 pd=0 as=0 ps=0 
M2405 io3 GND io3 GND efet w=28200 l=34200
+ ad=0 pd=0 as=0 ps=0 
M2406 GND diff_411600_867600# diff_446400_902400# GND efet w=16800 l=7200
+ ad=0 pd=0 as=1.30464e+09 ps=427200 
M2407 diff_494400_889200# io3 GND GND efet w=34800 l=7200
+ ad=8.352e+08 pd=182400 as=0 ps=0 
M2408 GND io3 diff_494400_889200# GND efet w=34800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2409 diff_648000_967200# diff_411600_867600# io2 GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2410 diff_1180800_985200# diff_564000_475200# diff_999600_1087200# GND efet w=22800 l=6000
+ ad=0 pd=0 as=1.57968e+09 ps=331200 
M2411 diff_967200_1083600# diff_999600_1087200# GND GND efet w=50400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2412 diff_999600_1087200# diff_999600_1087200# diff_999600_1087200# GND efet w=1200 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2413 diff_967200_1083600# Vdd Vdd GND efet w=9600 l=25200
+ ad=0 pd=0 as=0 ps=0 
M2414 diff_999600_1087200# diff_999600_1087200# diff_999600_1087200# GND efet w=1200 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2415 diff_1507200_984000# diff_564000_475200# diff_1344000_1008000# GND efet w=24000 l=6000
+ ad=0 pd=0 as=1.4976e+09 ps=316800 
M2416 diff_1834800_984000# diff_564000_475200# diff_1670400_1008000# GND efet w=21600 l=6000
+ ad=0 pd=0 as=1.81296e+09 ps=333600 
M2417 Vdd Vdd Vdd GND efet w=2400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2418 Vdd Vdd Vdd GND efet w=2400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2419 diff_446400_902400# diff_446400_902400# diff_446400_902400# GND efet w=2400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2420 Vdd Vdd Vdd GND efet w=1200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2421 Vdd Vdd diff_1180800_985200# GND efet w=6600 l=64800
+ ad=0 pd=0 as=0 ps=0 
M2422 Vdd Vdd diff_1016400_968400# GND efet w=6000 l=66000
+ ad=0 pd=0 as=0 ps=0 
M2423 Vdd Vdd Vdd GND efet w=1200 l=5400
+ ad=0 pd=0 as=0 ps=0 
M2424 diff_1344000_1008000# diff_1344000_1008000# diff_1344000_1008000# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2425 diff_1344000_1008000# diff_1344000_1008000# diff_1344000_1008000# GND efet w=1200 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2426 diff_1507200_984000# Vdd Vdd GND efet w=6000 l=64800
+ ad=0 pd=0 as=0 ps=0 
M2427 Vdd Vdd diff_829200_1039200# GND efet w=8400 l=24000
+ ad=0 pd=0 as=0 ps=0 
M2428 Vdd Vdd Vdd GND efet w=1200 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2429 Vdd Vdd diff_1342800_1122000# GND efet w=6000 l=64800
+ ad=0 pd=0 as=0 ps=0 
M2430 Vdd Vdd Vdd GND efet w=2400 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2431 diff_829200_1039200# diff_1344000_1008000# GND GND efet w=42000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2432 diff_1670400_984000# Vdd Vdd GND efet w=6600 l=67800
+ ad=0 pd=0 as=0 ps=0 
M2433 Vdd Vdd diff_682800_1034400# GND efet w=8400 l=39600
+ ad=0 pd=0 as=0 ps=0 
M2434 diff_2160000_985200# diff_564000_475200# diff_1996800_1008000# GND efet w=24000 l=7200
+ ad=0 pd=0 as=1.74096e+09 ps=321600 
M2435 diff_1834800_984000# Vdd Vdd GND efet w=5400 l=66600
+ ad=0 pd=0 as=0 ps=0 
M2436 diff_682800_1034400# diff_1670400_1008000# GND GND efet w=50400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2437 Vdd Vdd Vdd GND efet w=1200 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2438 diff_1344000_1008000# diff_624000_475200# diff_1342800_1122000# GND efet w=22800 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2439 diff_1996800_984000# Vdd Vdd GND efet w=7800 l=67800
+ ad=0 pd=0 as=0 ps=0 
M2440 diff_1670400_1008000# diff_624000_475200# diff_1670400_984000# GND efet w=24000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2441 diff_1996800_1008000# diff_624000_475200# diff_1996800_984000# GND efet w=24000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2442 Vdd Vdd diff_543600_1017600# GND efet w=8400 l=25200
+ ad=0 pd=0 as=0 ps=0 
M2443 diff_2160000_985200# Vdd Vdd GND efet w=7200 l=70800
+ ad=0 pd=0 as=0 ps=0 
M2444 diff_543600_1017600# diff_1996800_1008000# GND GND efet w=40800 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2445 Vdd Vdd diff_446400_902400# GND efet w=7200 l=44400
+ ad=0 pd=0 as=0 ps=0 
M2446 diff_446400_902400# diff_446400_902400# diff_446400_902400# GND efet w=1800 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2447 diff_999600_1087200# diff_624000_475200# diff_1016400_968400# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2448 io3 Vdd Vdd GND efet w=8400 l=12000
+ ad=0 pd=0 as=0 ps=0 
M2449 diff_567600_855600# diff_567600_855600# diff_567600_855600# GND efet w=1800 l=3600
+ ad=2.0016e+08 pd=76800 as=0 ps=0 
M2450 diff_411600_867600# diff_411600_867600# diff_411600_867600# GND efet w=600 l=1800
+ ad=1.86192e+09 pd=547200 as=0 ps=0 
M2451 diff_411600_867600# diff_411600_867600# diff_411600_867600# GND efet w=600 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2452 diff_567600_855600# diff_567600_855600# diff_567600_855600# GND efet w=1800 l=5400
+ ad=0 pd=0 as=0 ps=0 
M2453 diff_411600_867600# diff_411600_867600# diff_411600_867600# GND efet w=1200 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2454 diff_646800_888000# io2 GND GND efet w=34800 l=7200
+ ad=8.4384e+08 pd=184800 as=0 ps=0 
M2455 GND io2 diff_646800_888000# GND efet w=34800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2456 diff_802800_967200# diff_411600_867600# io1 GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2457 diff_901200_968400# diff_411600_867600# io0 GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2458 io2 Vdd Vdd GND efet w=8400 l=12000
+ ad=0 pd=0 as=0 ps=0 
M2459 diff_567600_855600# Vdd Vdd GND efet w=7200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2460 diff_411600_867600# clk1 diff_411600_853200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=2.8944e+08 ps=110400 
M2461 diff_411600_853200# diff_411600_853200# diff_411600_853200# GND efet w=1800 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2462 GND diff_411600_853200# diff_446400_902400# GND efet w=36600 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2463 Vdd Vdd diff_494400_889200# GND efet w=7200 l=21600
+ ad=0 pd=0 as=0 ps=0 
M2464 diff_411600_853200# diff_411600_853200# diff_411600_853200# GND efet w=1800 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2465 Vdd Vdd Vdd GND efet w=1200 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2466 Vdd diff_567600_855600# diff_411600_867600# GND efet w=9000 l=21600
+ ad=0 pd=0 as=0 ps=0 
M2467 Vdd Vdd diff_481200_801600# GND efet w=7200 l=14400
+ ad=0 pd=0 as=8.2224e+08 ps=220800 
M2468 diff_411600_867600# diff_567600_855600# diff_411600_867600# GND efet w=46800 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2469 diff_801600_888000# io1 GND GND efet w=34800 l=7200
+ ad=8.352e+08 pd=182400 as=0 ps=0 
M2470 GND io1 diff_801600_888000# GND efet w=34800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2471 diff_1180800_985200# diff_1014000_962400# diff_1159200_908400# GND efet w=39600 l=7200
+ ad=0 pd=0 as=1.69344e+09 ps=453600 
M2472 diff_1342800_1122000# diff_1014000_962400# diff_1321200_904800# GND efet w=39000 l=6600
+ ad=0 pd=0 as=1.71504e+09 ps=460800 
M2473 diff_2160000_985200# diff_1014000_962400# diff_2138400_908400# GND efet w=40800 l=7200
+ ad=0 pd=0 as=1.7136e+09 ps=458400 
M2474 diff_1507200_984000# diff_1014000_962400# diff_1485600_907200# GND efet w=39600 l=6000
+ ad=0 pd=0 as=1.78848e+09 ps=463200 
M2475 diff_1670400_984000# diff_1014000_962400# diff_1648800_908400# GND efet w=39600 l=6000
+ ad=0 pd=0 as=1.7568e+09 ps=458400 
M2476 diff_1016400_968400# diff_1014000_962400# diff_999600_896400# GND efet w=40800 l=7200
+ ad=0 pd=0 as=1.96128e+09 ps=472800 
M2477 diff_1016400_968400# diff_1124400_963600# diff_1077600_907200# GND efet w=40800 l=6000
+ ad=0 pd=0 as=1.62864e+09 ps=403200 
M2478 diff_1180800_985200# diff_1124400_963600# diff_1239600_907200# GND efet w=40800 l=6000
+ ad=0 pd=0 as=1.55808e+09 ps=398400 
M2479 diff_1342800_1122000# diff_1124400_963600# diff_1404000_907200# GND efet w=40800 l=6000
+ ad=0 pd=0 as=1.68192e+09 ps=408000 
M2480 diff_1507200_984000# diff_1124400_963600# diff_1567200_907200# GND efet w=40800 l=6000
+ ad=0 pd=0 as=1.68192e+09 ps=408000 
M2481 diff_1834800_984000# diff_1014000_962400# diff_1813200_908400# GND efet w=39600 l=6000
+ ad=0 pd=0 as=1.73664e+09 ps=456000 
M2482 diff_1670400_984000# diff_1124400_963600# diff_1731600_907200# GND efet w=40800 l=6000
+ ad=0 pd=0 as=1.63152e+09 ps=403200 
M2483 diff_1996800_984000# diff_1014000_962400# diff_1975200_908400# GND efet w=39600 l=6000
+ ad=0 pd=0 as=1.73088e+09 ps=456000 
M2484 diff_1834800_984000# diff_1124400_963600# diff_1893600_907200# GND efet w=40800 l=6000
+ ad=0 pd=0 as=1.62576e+09 ps=403200 
M2485 diff_1996800_984000# diff_1124400_963600# diff_2056800_907200# GND efet w=40800 l=6000
+ ad=0 pd=0 as=1.62576e+09 ps=403200 
M2486 diff_2160000_985200# diff_1124400_963600# diff_2221200_907200# GND efet w=34800 l=4800
+ ad=0 pd=0 as=1.70496e+09 ps=417600 
M2487 diff_2299200_829200# diff_1063200_940800# diff_2221200_907200# GND efet w=43800 l=6600
+ ad=8.5968e+08 pd=249600 as=0 ps=0 
M2488 diff_999600_896400# diff_1063200_940800# diff_1074000_927600# GND efet w=31200 l=6000
+ ad=0 pd=0 as=7.0704e+08 ps=177600 
M2489 diff_1077600_907200# diff_1063200_940800# diff_1155600_927600# GND efet w=31200 l=6000
+ ad=0 pd=0 as=7.128e+08 ps=177600 
M2490 diff_1159200_908400# diff_1063200_940800# diff_1236000_926400# GND efet w=31200 l=6000
+ ad=0 pd=0 as=7.4448e+08 ps=180000 
M2491 diff_1239600_907200# diff_1063200_940800# diff_1317600_926400# GND efet w=31200 l=6000
+ ad=0 pd=0 as=7.5024e+08 ps=180000 
M2492 diff_1321200_904800# diff_1063200_940800# diff_1400400_928800# GND efet w=31200 l=6000
+ ad=0 pd=0 as=6.696e+08 ps=175200 
M2493 diff_1404000_907200# diff_1063200_940800# diff_1482000_928800# GND efet w=31200 l=6000
+ ad=0 pd=0 as=6.7536e+08 ps=175200 
M2494 diff_1485600_907200# diff_1063200_940800# diff_1563600_928800# GND efet w=31200 l=6000
+ ad=0 pd=0 as=6.696e+08 ps=175200 
M2495 diff_1567200_907200# diff_1063200_940800# diff_1645200_928800# GND efet w=31200 l=6000
+ ad=0 pd=0 as=6.7536e+08 ps=175200 
M2496 diff_1648800_908400# diff_1063200_940800# diff_1728000_927600# GND efet w=31200 l=6000
+ ad=0 pd=0 as=7.0704e+08 ps=177600 
M2497 diff_1731600_907200# diff_1063200_940800# diff_1809600_927600# GND efet w=31200 l=6000
+ ad=0 pd=0 as=7.128e+08 ps=177600 
M2498 diff_1813200_908400# diff_1063200_940800# diff_1890000_927600# GND efet w=31200 l=6000
+ ad=0 pd=0 as=7.0704e+08 ps=177600 
M2499 diff_1893600_907200# diff_1063200_940800# diff_1971600_927600# GND efet w=31200 l=6000
+ ad=0 pd=0 as=7.128e+08 ps=177600 
M2500 diff_1975200_908400# diff_1063200_940800# diff_2053200_927600# GND efet w=31200 l=6000
+ ad=0 pd=0 as=7.0704e+08 ps=177600 
M2501 diff_2056800_907200# diff_1063200_940800# diff_2134800_927600# GND efet w=31200 l=6000
+ ad=0 pd=0 as=7.128e+08 ps=177600 
M2502 diff_2138400_908400# diff_1063200_940800# diff_2217600_927600# GND efet w=30000 l=6000
+ ad=0 pd=0 as=6.9696e+08 ps=175200 
M2503 io1 Vdd Vdd GND efet w=8400 l=12000
+ ad=0 pd=0 as=0 ps=0 
M2504 diff_898800_888000# io0 GND GND efet w=34800 l=7200
+ ad=8.4384e+08 pd=184800 as=0 ps=0 
M2505 GND io0 diff_898800_888000# GND efet w=34800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2506 io0 Vdd Vdd GND efet w=8400 l=12000
+ ad=0 pd=0 as=0 ps=0 
M2507 Vdd Vdd diff_646800_888000# GND efet w=7200 l=22800
+ ad=0 pd=0 as=0 ps=0 
M2508 Vdd Vdd diff_801600_888000# GND efet w=7200 l=21600
+ ad=0 pd=0 as=0 ps=0 
M2509 Vdd Vdd diff_898800_888000# GND efet w=7200 l=20400
+ ad=0 pd=0 as=0 ps=0 
M2510 GND diff_496800_798000# diff_481200_801600# GND efet w=61200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2511 diff_481200_801600# diff_406800_692400# diff_447600_771600# GND efet w=12000 l=7200
+ ad=0 pd=0 as=1.6704e+08 ps=52800 
M2512 diff_1077600_907200# diff_1033200_919200# diff_1116000_907200# GND efet w=34200 l=6600
+ ad=0 pd=0 as=7.9056e+08 ps=199200 
M2513 diff_1159200_908400# diff_1033200_919200# diff_1197600_907200# GND efet w=33600 l=8400
+ ad=0 pd=0 as=8.0784e+08 ps=199200 
M2514 diff_1321200_904800# diff_1033200_919200# diff_1359600_906000# GND efet w=34800 l=6000
+ ad=0 pd=0 as=8.4672e+08 ps=204000 
M2515 diff_1239600_907200# diff_1033200_919200# diff_1278000_906000# GND efet w=33600 l=7800
+ ad=0 pd=0 as=8.2656e+08 ps=199200 
M2516 diff_1404000_907200# diff_1033200_919200# diff_1442400_908400# GND efet w=33600 l=7800
+ ad=0 pd=0 as=7.5168e+08 ps=194400 
M2517 diff_1485600_907200# diff_1033200_919200# diff_1524000_908400# GND efet w=34200 l=8400
+ ad=0 pd=0 as=7.704e+08 ps=196800 
M2518 diff_1567200_907200# diff_1033200_919200# diff_1605600_908400# GND efet w=33600 l=7800
+ ad=0 pd=0 as=7.5168e+08 ps=194400 
M2519 diff_1648800_908400# diff_1033200_919200# diff_1687200_908400# GND efet w=33600 l=8400
+ ad=0 pd=0 as=7.704e+08 ps=196800 
M2520 diff_1731600_907200# diff_1033200_919200# diff_1770000_907200# GND efet w=33000 l=7800
+ ad=0 pd=0 as=7.8912e+08 ps=196800 
M2521 diff_1893600_907200# diff_1033200_919200# diff_1932000_907200# GND efet w=33600 l=8400
+ ad=0 pd=0 as=7.8912e+08 ps=196800 
M2522 diff_1813200_908400# diff_1033200_919200# diff_1851600_907200# GND efet w=33000 l=7800
+ ad=0 pd=0 as=8.0784e+08 ps=199200 
M2523 diff_1975200_908400# diff_1033200_919200# diff_2013600_907200# GND efet w=33600 l=8400
+ ad=0 pd=0 as=8.0784e+08 ps=199200 
M2524 diff_2056800_907200# diff_1033200_919200# diff_2095200_907200# GND efet w=33600 l=8400
+ ad=0 pd=0 as=7.8912e+08 ps=196800 
M2525 diff_2138400_908400# diff_1033200_919200# diff_2176800_907200# GND efet w=33600 l=8400
+ ad=0 pd=0 as=8.0784e+08 ps=199200 
M2526 diff_2221200_907200# diff_1033200_919200# diff_2259600_907200# GND efet w=32400 l=8400
+ ad=0 pd=0 as=7.6464e+08 ps=194400 
M2527 diff_411600_867600# diff_411600_867600# diff_411600_867600# GND efet w=1200 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2528 diff_999600_896400# diff_1033200_919200# diff_1036800_903600# GND efet w=28800 l=6000
+ ad=0 pd=0 as=7.8336e+08 ps=194400 
M2529 diff_1077600_907200# diff_994800_1225200# diff_1075200_826800# GND efet w=30600 l=6600
+ ad=0 pd=0 as=6.7104e+08 ps=189600 
M2530 diff_1159200_908400# diff_994800_1225200# diff_1156800_829200# GND efet w=31200 l=6600
+ ad=0 pd=0 as=6.912e+08 ps=189600 
M2531 diff_1321200_904800# diff_994800_1225200# diff_1320000_829200# GND efet w=34200 l=6000
+ ad=0 pd=0 as=7.1712e+08 ps=192000 
M2532 diff_1239600_907200# diff_994800_1225200# diff_1238400_829200# GND efet w=31200 l=6600
+ ad=0 pd=0 as=6.8544e+08 ps=189600 
M2533 diff_1404000_907200# diff_994800_1225200# diff_1401600_829200# GND efet w=31200 l=6600
+ ad=0 pd=0 as=6.264e+08 ps=187200 
M2534 diff_1485600_907200# diff_994800_1225200# diff_1483200_829200# GND efet w=32400 l=6000
+ ad=0 pd=0 as=6.5088e+08 ps=187200 
M2535 diff_1567200_907200# diff_994800_1225200# diff_1564800_829200# GND efet w=31200 l=6600
+ ad=0 pd=0 as=6.264e+08 ps=187200 
M2536 diff_1648800_908400# diff_994800_1225200# diff_1646400_829200# GND efet w=31200 l=6600
+ ad=0 pd=0 as=6.552e+08 ps=187200 
M2537 diff_1731600_907200# diff_994800_1225200# diff_1728000_829200# GND efet w=30000 l=6000
+ ad=0 pd=0 as=6.6672e+08 ps=189600 
M2538 diff_1813200_908400# diff_994800_1225200# diff_1809600_829200# GND efet w=30600 l=6600
+ ad=0 pd=0 as=6.9408e+08 ps=189600 
M2539 diff_1893600_907200# diff_994800_1225200# diff_1891200_829200# GND efet w=30600 l=6600
+ ad=0 pd=0 as=6.6528e+08 ps=189600 
M2540 diff_1975200_908400# diff_994800_1225200# diff_1972800_829200# GND efet w=31200 l=6600
+ ad=0 pd=0 as=6.912e+08 ps=189600 
M2541 diff_2056800_907200# diff_994800_1225200# diff_2054400_829200# GND efet w=30600 l=6600
+ ad=0 pd=0 as=6.6528e+08 ps=189600 
M2542 diff_2138400_908400# diff_994800_1225200# diff_2136000_829200# GND efet w=31200 l=6600
+ ad=0 pd=0 as=6.912e+08 ps=189600 
M2543 diff_2221200_907200# diff_994800_1225200# diff_2217600_829200# GND efet w=28800 l=6000
+ ad=0 pd=0 as=6.4656e+08 ps=184800 
M2544 diff_999600_896400# diff_994800_1225200# diff_997200_836400# GND efet w=38400 l=4800
+ ad=0 pd=0 as=8.3952e+08 ps=194400 
M2545 diff_1033200_850800# diff_1024800_849600# GND GND efet w=46800 l=7200
+ ad=3.6432e+08 pd=105600 as=0 ps=0 
M2546 diff_411600_867600# diff_411600_867600# diff_411600_867600# GND efet w=600 l=1800
+ ad=0 pd=0 as=0 ps=0 
M2547 GND diff_447600_771600# diff_189600_804000# GND efet w=91200 l=7200
+ ad=0 pd=0 as=1.05607e+09 ps=1.1808e+06 
M2548 diff_189600_804000# diff_421200_728400# Vdd GND efet w=83400 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2549 diff_558000_765600# diff_409200_476400# diff_536400_776400# GND efet w=36000 l=7200
+ ad=8.64e+08 pd=228000 as=8.4528e+08 ps=220800 
M2550 diff_536400_776400# diff_339600_532800# diff_496800_798000# GND efet w=39600 l=7200
+ ad=0 pd=0 as=6.0192e+08 ps=151200 
M2551 GND diff_1008000_775200# diff_997200_836400# GND efet w=28800 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2552 diff_999600_896400# diff_1048800_846000# diff_1033200_850800# GND efet w=31200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2553 GND diff_1089600_775200# diff_1074000_927600# GND efet w=35400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2554 diff_1116000_849600# diff_1110000_775200# GND GND efet w=36000 l=7200
+ ad=3.3264e+08 pd=93600 as=0 ps=0 
M2555 diff_1077600_907200# diff_1048800_846000# diff_1116000_849600# GND efet w=30000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2556 GND diff_1171200_775200# diff_1155600_927600# GND efet w=35400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2557 diff_1197600_849600# diff_1191600_775200# GND GND efet w=36000 l=7200
+ ad=3.3264e+08 pd=93600 as=0 ps=0 
M2558 diff_1159200_908400# diff_1048800_846000# diff_1197600_849600# GND efet w=30000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2559 GND diff_1252800_775200# diff_1236000_926400# GND efet w=35400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2560 diff_1279200_849600# diff_1273200_775200# GND GND efet w=36000 l=7200
+ ad=3.3264e+08 pd=93600 as=0 ps=0 
M2561 diff_1239600_907200# diff_1048800_846000# diff_1279200_849600# GND efet w=30000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2562 GND diff_1334400_775200# diff_1317600_926400# GND efet w=35400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2563 diff_1360800_849600# diff_1354800_775200# GND GND efet w=36000 l=7200
+ ad=3.3264e+08 pd=93600 as=0 ps=0 
M2564 diff_1321200_904800# diff_1048800_846000# diff_1360800_849600# GND efet w=30000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2565 GND diff_1416000_775200# diff_1400400_928800# GND efet w=35400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2566 diff_1442400_849600# diff_1436400_775200# GND GND efet w=36000 l=7200
+ ad=3.3264e+08 pd=93600 as=0 ps=0 
M2567 diff_1404000_907200# diff_1048800_846000# diff_1442400_849600# GND efet w=30000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2568 GND diff_1497600_775200# diff_1482000_928800# GND efet w=35400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2569 diff_1524000_849600# diff_1518000_775200# GND GND efet w=36000 l=7200
+ ad=3.3264e+08 pd=93600 as=0 ps=0 
M2570 diff_1485600_907200# diff_1048800_846000# diff_1524000_849600# GND efet w=30000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2571 GND diff_1579200_775200# diff_1563600_928800# GND efet w=35400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2572 diff_1605600_849600# diff_1599600_775200# GND GND efet w=36000 l=7200
+ ad=3.3264e+08 pd=93600 as=0 ps=0 
M2573 diff_1567200_907200# diff_1048800_846000# diff_1605600_849600# GND efet w=30000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2574 GND diff_1660800_775200# diff_1645200_928800# GND efet w=35400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2575 diff_1687200_849600# diff_1681200_775200# GND GND efet w=36000 l=7200
+ ad=3.3264e+08 pd=93600 as=0 ps=0 
M2576 diff_1648800_908400# diff_1048800_846000# diff_1687200_849600# GND efet w=30000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2577 GND diff_1742400_775200# diff_1728000_927600# GND efet w=35400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2578 diff_1768800_849600# diff_1762800_775200# GND GND efet w=36000 l=7200
+ ad=3.3264e+08 pd=93600 as=0 ps=0 
M2579 diff_1731600_907200# diff_1048800_846000# diff_1768800_849600# GND efet w=30000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2580 GND diff_1824000_775200# diff_1809600_927600# GND efet w=35400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2581 diff_1850400_849600# diff_1844400_775200# GND GND efet w=36000 l=7200
+ ad=3.3264e+08 pd=93600 as=0 ps=0 
M2582 diff_1813200_908400# diff_1048800_846000# diff_1850400_849600# GND efet w=30000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2583 GND diff_1905600_775200# diff_1890000_927600# GND efet w=35400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2584 diff_1932000_849600# diff_1926000_775200# GND GND efet w=36000 l=7200
+ ad=3.3264e+08 pd=93600 as=0 ps=0 
M2585 diff_1893600_907200# diff_1048800_846000# diff_1932000_849600# GND efet w=30000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2586 GND diff_1987200_775200# diff_1971600_927600# GND efet w=35400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2587 diff_2013600_849600# diff_2007600_775200# GND GND efet w=36000 l=7200
+ ad=3.3264e+08 pd=93600 as=0 ps=0 
M2588 diff_1975200_908400# diff_1048800_846000# diff_2013600_849600# GND efet w=30000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2589 GND diff_2068800_775200# diff_2053200_927600# GND efet w=35400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2590 diff_2095200_849600# diff_2089200_775200# GND GND efet w=36000 l=7200
+ ad=3.3264e+08 pd=93600 as=0 ps=0 
M2591 diff_2056800_907200# diff_1048800_846000# diff_2095200_849600# GND efet w=30000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2592 GND diff_2150400_775200# diff_2134800_927600# GND efet w=35400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2593 diff_2176800_849600# diff_2170800_775200# GND GND efet w=36000 l=7200
+ ad=3.3264e+08 pd=93600 as=0 ps=0 
M2594 diff_2138400_908400# diff_1048800_846000# diff_2176800_849600# GND efet w=30000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2595 GND diff_2232000_775200# diff_2217600_927600# GND efet w=35400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2596 diff_2258400_849600# diff_2252400_775200# GND GND efet w=36000 l=7200
+ ad=3.3264e+08 pd=93600 as=0 ps=0 
M2597 diff_2221200_907200# diff_1048800_846000# diff_2258400_849600# GND efet w=30000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2598 diff_2592000_1532400# Vdd Vdd GND efet w=13200 l=7200
+ ad=1.5696e+08 pd=57600 as=0 ps=0 
M2599 diff_2592000_1532400# diff_2592000_1532400# diff_2592000_1532400# GND efet w=1800 l=5400
+ ad=0 pd=0 as=0 ps=0 
M2600 diff_2592000_1532400# diff_2592000_1532400# diff_2592000_1532400# GND efet w=1800 l=1800
+ ad=0 pd=0 as=0 ps=0 
M2601 Vdd Vdd Vdd GND efet w=600 l=1800
+ ad=0 pd=0 as=0 ps=0 
M2602 GND diff_2767200_1582800# diff_2649600_1519200# GND efet w=80400 l=6000
+ ad=0 pd=0 as=1.30896e+09 ps=252000 
M2603 Vdd Vdd diff_2649600_1519200# GND efet w=8400 l=16800
+ ad=0 pd=0 as=0 ps=0 
M2604 Vdd Vdd Vdd GND efet w=600 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2605 GND d2 diff_2812800_1003200# GND efet w=195600 l=6000
+ ad=0 pd=0 as=2.04336e+09 ps=396000 
M2606 diff_2812800_1003200# Vdd Vdd GND efet w=8400 l=16800
+ ad=0 pd=0 as=0 ps=0 
M2607 diff_2649600_1519200# clk1 diff_2768400_1540800# GND efet w=13200 l=6000
+ ad=0 pd=0 as=1.6848e+08 ps=55200 
M2608 Vdd Vdd diff_2812800_1134000# GND efet w=8400 l=16800
+ ad=0 pd=0 as=1.09296e+09 ps=228000 
M2609 diff_2768400_1540800# diff_2768400_1540800# diff_2768400_1540800# GND efet w=1800 l=1800
+ ad=0 pd=0 as=0 ps=0 
M2610 GND diff_2768400_1540800# diff_2710800_1356000# GND efet w=44400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2611 Vdd Vdd diff_2710800_1356000# GND efet w=9600 l=19200
+ ad=0 pd=0 as=0 ps=0 
M2612 Vdd Vdd Vdd GND efet w=2400 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2613 Vdd Vdd Vdd GND efet w=2400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2614 diff_2710800_1356000# clk2 diff_2768400_1497600# GND efet w=12000 l=6000
+ ad=0 pd=0 as=1.3824e+08 ps=48000 
M2615 diff_1003200_1702800# diff_2589600_1464000# Vdd GND efet w=15600 l=6000
+ ad=-4.24247e+08 pd=739200 as=0 ps=0 
M2616 GND diff_2649600_1428000# diff_1003200_1702800# GND efet w=296400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2617 diff_1003200_1702800# diff_2589600_1464000# diff_1003200_1702800# GND efet w=40800 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2618 diff_2589600_1464000# Vdd Vdd GND efet w=12000 l=6000
+ ad=1.7424e+08 pd=60000 as=0 ps=0 
M2619 diff_2589600_1464000# diff_2589600_1464000# diff_2589600_1464000# GND efet w=1200 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2620 diff_2589600_1464000# diff_2589600_1464000# diff_2589600_1464000# GND efet w=1800 l=1800
+ ad=0 pd=0 as=0 ps=0 
M2621 diff_2768400_1497600# diff_2768400_1497600# diff_2768400_1497600# GND efet w=1200 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2622 GND diff_2768400_1497600# diff_2664000_1422000# GND efet w=44400 l=7200
+ ad=0 pd=0 as=1.56816e+09 ps=336000 
M2623 Vdd Vdd diff_2664000_1422000# GND efet w=8400 l=18000
+ ad=0 pd=0 as=0 ps=0 
M2624 Vdd Vdd Vdd GND efet w=600 l=1800
+ ad=0 pd=0 as=0 ps=0 
M2625 GND diff_2812800_1003200# diff_2812800_1134000# GND efet w=44400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2626 diff_2664000_1422000# clk1 diff_2767200_1456800# GND efet w=14400 l=6000
+ ad=0 pd=0 as=1.6704e+08 ps=52800 
M2627 GND diff_2767200_1456800# diff_2722800_844800# GND efet w=44400 l=6000
+ ad=0 pd=0 as=1.13616e+09 ps=225600 
M2628 Vdd Vdd diff_2722800_844800# GND efet w=8400 l=16800
+ ad=0 pd=0 as=0 ps=0 
M2629 Vdd Vdd Vdd GND efet w=1200 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2630 Vdd Vdd Vdd GND efet w=1200 l=1800
+ ad=0 pd=0 as=0 ps=0 
M2631 GND diff_2664000_1422000# diff_2626800_1411200# GND efet w=13200 l=6000
+ ad=0 pd=0 as=4.824e+08 ps=139200 
M2632 diff_2626800_1411200# Vdd Vdd GND efet w=7200 l=36000
+ ad=0 pd=0 as=0 ps=0 
M2633 diff_2605200_1372800# Vdd Vdd GND efet w=7200 l=18000
+ ad=7.1568e+08 pd=175200 as=0 ps=0 
M2634 diff_2708400_1392000# diff_2664000_1422000# diff_2601600_1368000# GND efet w=15600 l=6000
+ ad=2.8368e+08 pd=88800 as=5.1552e+08 ps=136800 
M2635 diff_2605200_1372800# diff_2601600_1368000# GND GND efet w=61200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2636 diff_2601600_1368000# diff_2601600_1368000# diff_2601600_1368000# GND efet w=3000 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2637 diff_2601600_1368000# diff_2601600_1368000# diff_2601600_1368000# GND efet w=1800 l=1800
+ ad=0 pd=0 as=0 ps=0 
M2638 diff_2708400_1392000# diff_2613600_1719600# diff_2710800_1356000# GND efet w=13200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2639 diff_2601600_1368000# diff_2626800_1411200# GND GND efet w=12000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2640 diff_2738400_1274400# diff_2710800_1356000# diff_2526000_1243200# GND efet w=20400 l=6000
+ ad=5.688e+08 pd=136800 as=2.9088e+08 ps=69600 
M2641 diff_2774400_1308000# clk2 diff_2738400_1274400# GND efet w=20400 l=6000
+ ad=9.9216e+08 pd=163200 as=0 ps=0 
M2642 GND diff_2568000_1281600# diff_1124400_1153200# GND efet w=140400 l=6000
+ ad=0 pd=0 as=1.95408e+09 ps=396000 
M2643 diff_2738400_1274400# diff_2722800_844800# diff_2568000_1281600# GND efet w=19200 l=6000
+ ad=0 pd=0 as=2.5056e+08 ps=64800 
M2644 GND diff_411600_867600# diff_536400_776400# GND efet w=27000 l=7800
+ ad=0 pd=0 as=0 ps=0 
M2645 diff_558000_765600# diff_564000_475200# GND GND efet w=37200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2646 GND diff_624000_475200# diff_558000_765600# GND efet w=36000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2647 diff_825600_782400# d3 GND GND efet w=36600 l=6600
+ ad=8.8704e+08 pd=211200 as=0 ps=0 
M2648 GND diff_700800_679200# diff_696000_782400# GND efet w=21600 l=7200
+ ad=0 pd=0 as=3.4272e+08 ps=81600 
M2649 GND diff_696000_782400# diff_154800_822000# GND efet w=16800 l=7200
+ ad=0 pd=0 as=-1.96505e+09 ps=736800 
M2650 diff_816000_787200# clk2 diff_700800_679200# GND efet w=10800 l=7200
+ ad=1.0368e+08 pd=40800 as=3.4272e+08 ps=110400 
M2651 Vdd diff_825600_782400# diff_816000_787200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2652 diff_825600_782400# Vdd Vdd GND efet w=7200 l=33600
+ ad=0 pd=0 as=0 ps=0 
M2653 GND diff_694800_556800# diff_825600_782400# GND efet w=18000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2654 GND diff_919200_421200# diff_825600_782400# GND efet w=18000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2655 GND diff_1048800_775200# diff_1036800_903600# GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2656 diff_1075200_826800# diff_1069200_775200# GND GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2657 GND diff_1130400_775200# diff_1116000_907200# GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2658 diff_1156800_829200# diff_1150800_775200# GND GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2659 GND diff_1212000_775200# diff_1197600_907200# GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2660 diff_1238400_829200# diff_1232400_775200# GND GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2661 GND diff_1293600_775200# diff_1278000_906000# GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2662 diff_1320000_829200# diff_1314000_775200# GND GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2663 GND diff_1375200_775200# diff_1359600_906000# GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2664 diff_1401600_829200# diff_1395600_775200# GND GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2665 GND diff_1456800_775200# diff_1442400_908400# GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2666 diff_1483200_829200# diff_1477200_775200# GND GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2667 GND diff_1538400_775200# diff_1524000_908400# GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2668 diff_1564800_829200# diff_1558800_775200# GND GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2669 GND diff_1620000_775200# diff_1605600_908400# GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2670 diff_1646400_829200# diff_1640400_775200# GND GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2671 GND diff_1701600_775200# diff_1687200_908400# GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2672 diff_1728000_829200# diff_1722000_775200# GND GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2673 GND diff_1783200_775200# diff_1770000_907200# GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2674 diff_1809600_829200# diff_1803600_775200# GND GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2675 GND diff_1864800_775200# diff_1851600_907200# GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2676 diff_1891200_829200# diff_1885200_775200# GND GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2677 GND diff_1946400_775200# diff_1932000_907200# GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2678 diff_1972800_829200# diff_1966800_775200# GND GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2679 GND diff_2028000_775200# diff_2013600_907200# GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2680 diff_2054400_829200# diff_2048400_775200# GND GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2681 GND diff_2109600_775200# diff_2095200_907200# GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2682 diff_2136000_829200# diff_2130000_775200# GND GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2683 GND diff_2191200_775200# diff_2176800_907200# GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2684 diff_2217600_829200# diff_2211600_775200# GND GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2685 GND diff_2272800_775200# diff_2259600_907200# GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2686 diff_2299200_829200# diff_2293200_775200# GND GND efet w=39600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2687 GND diff_481200_801600# diff_498000_715200# GND efet w=48600 l=6600
+ ad=0 pd=0 as=3.9024e+08 ps=124800 
M2688 diff_498000_715200# diff_406800_692400# diff_421200_728400# GND efet w=10800 l=6000
+ ad=0 pd=0 as=3.1248e+08 ps=100800 
M2689 diff_498000_715200# Vdd Vdd GND efet w=7200 l=15600
+ ad=0 pd=0 as=0 ps=0 
M2690 Vdd Vdd Vdd GND efet w=1200 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2691 Vdd Vdd Vdd GND efet w=1800 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2692 Vdd Vdd diff_496800_798000# GND efet w=7200 l=67200
+ ad=0 pd=0 as=0 ps=0 
M2693 Vdd Vdd Vdd GND efet w=1800 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2694 Vdd Vdd Vdd GND efet w=1800 l=5400
+ ad=0 pd=0 as=0 ps=0 
M2695 diff_260400_786000# Vdd Vdd GND efet w=9600 l=18000
+ ad=9.5184e+08 pd=213600 as=0 ps=0 
M2696 diff_406800_692400# diff_480000_614400# Vdd GND efet w=8400 l=8400
+ ad=9.8352e+08 pd=240000 as=0 ps=0 
M2697 diff_406800_692400# diff_480000_614400# diff_406800_692400# GND efet w=46200 l=23400
+ ad=0 pd=0 as=0 ps=0 
M2698 diff_480000_614400# Vdd Vdd GND efet w=8400 l=7200
+ ad=1.8e+08 pd=57600 as=0 ps=0 
M2699 Vdd Vdd diff_339600_532800# GND efet w=8400 l=18000
+ ad=0 pd=0 as=1.39104e+09 ps=292800 
M2700 diff_260400_786000# diff_339600_532800# GND GND efet w=86400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2701 GND clk2 diff_406800_692400# GND efet w=45600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2702 Vdd Vdd Vdd GND efet w=3000 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2703 reset GND reset GND efet w=182400 l=112800
+ ad=-7.16567e+08 pd=873600 as=0 ps=0 
M2704 diff_339600_532800# reset GND GND efet w=144600 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2705 Vdd Vdd Vdd GND efet w=1800 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2706 sync clk2 diff_284400_465600# GND efet w=12000 l=7200
+ ad=0 pd=0 as=1.8144e+08 ps=60000 
M2707 diff_284400_465600# diff_284400_465600# diff_284400_465600# GND efet w=2400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2708 diff_284400_465600# diff_284400_465600# diff_284400_465600# GND efet w=1200 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2709 GND diff_284400_465600# diff_289200_457200# GND efet w=40200 l=6600
+ ad=0 pd=0 as=1.11456e+09 ps=295200 
M2710 Vdd Vdd Vdd GND efet w=600 l=1800
+ ad=0 pd=0 as=0 ps=0 
M2711 Vdd Vdd diff_409200_476400# GND efet w=9000 l=35400
+ ad=0 pd=0 as=3.7584e+08 ps=100800 
M2712 Vdd Vdd diff_490800_500400# GND efet w=8400 l=64800
+ ad=0 pd=0 as=4.1904e+08 ps=98400 
M2713 diff_154800_822000# diff_694800_762000# GND GND efet w=16800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2714 diff_154800_822000# Vdd Vdd GND efet w=7200 l=33600
+ ad=0 pd=0 as=0 ps=0 
M2715 Vdd Vdd Vdd GND efet w=1200 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2716 Vdd Vdd Vdd GND efet w=1200 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2717 diff_696000_782400# Vdd Vdd GND efet w=7200 l=50400
+ ad=0 pd=0 as=0 ps=0 
M2718 diff_700800_679200# diff_338400_375600# GND GND efet w=12000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2719 diff_700800_679200# diff_700800_679200# diff_700800_679200# GND efet w=1800 l=1800
+ ad=0 pd=0 as=0 ps=0 
M2720 diff_700800_679200# diff_700800_679200# diff_700800_679200# GND efet w=600 l=1800
+ ad=0 pd=0 as=0 ps=0 
M2721 diff_904800_769200# Vdd Vdd GND efet w=7200 l=51600
+ ad=5.8464e+08 pd=175200 as=0 ps=0 
M2722 GND d3 diff_904800_769200# GND efet w=28800 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2723 diff_1008000_775200# diff_1004400_769200# diff_1008000_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2724 diff_1024800_849600# diff_1004400_769200# diff_1028400_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2725 diff_1048800_775200# diff_1004400_769200# diff_1048800_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2726 diff_1069200_775200# diff_1004400_769200# diff_1069200_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2727 diff_1089600_775200# diff_1004400_769200# diff_1089600_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2728 diff_1110000_775200# diff_1004400_769200# diff_1110000_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2729 diff_1130400_775200# diff_1004400_769200# diff_1130400_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2730 diff_1150800_775200# diff_1004400_769200# diff_1150800_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2731 diff_1171200_775200# diff_1004400_769200# diff_1171200_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2732 diff_1191600_775200# diff_1004400_769200# diff_1191600_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2733 diff_1212000_775200# diff_1004400_769200# diff_1212000_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2734 diff_1232400_775200# diff_1004400_769200# diff_1232400_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2735 diff_1252800_775200# diff_1004400_769200# diff_1252800_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2736 diff_1273200_775200# diff_1004400_769200# diff_1273200_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2737 diff_1293600_775200# diff_1004400_769200# diff_1293600_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2738 diff_1314000_775200# diff_1004400_769200# diff_1314000_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2739 diff_1334400_775200# diff_1004400_769200# diff_1334400_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2740 diff_1354800_775200# diff_1004400_769200# diff_1354800_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2741 diff_1375200_775200# diff_1004400_769200# diff_1375200_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2742 diff_1395600_775200# diff_1004400_769200# diff_1395600_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2743 diff_1416000_775200# diff_1004400_769200# diff_1416000_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2744 diff_1436400_775200# diff_1004400_769200# diff_1436400_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2745 diff_1456800_775200# diff_1004400_769200# diff_1456800_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2746 diff_1477200_775200# diff_1004400_769200# diff_1477200_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2747 diff_1497600_775200# diff_1004400_769200# diff_1497600_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2748 diff_1518000_775200# diff_1004400_769200# diff_1518000_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2749 diff_1538400_775200# diff_1004400_769200# diff_1538400_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2750 diff_1558800_775200# diff_1004400_769200# diff_1558800_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2751 diff_1579200_775200# diff_1004400_769200# diff_1579200_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2752 diff_1599600_775200# diff_1004400_769200# diff_1599600_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2753 diff_1620000_775200# diff_1004400_769200# diff_1620000_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2754 diff_1640400_775200# diff_1004400_769200# diff_1640400_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2755 diff_1660800_775200# diff_1004400_769200# diff_1660800_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2756 diff_1681200_775200# diff_1004400_769200# diff_1681200_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2757 diff_1701600_775200# diff_1004400_769200# diff_1701600_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2758 diff_1722000_775200# diff_1004400_769200# diff_1722000_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2759 diff_1742400_775200# diff_1004400_769200# diff_1742400_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2760 diff_1762800_775200# diff_1004400_769200# diff_1762800_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2761 diff_1783200_775200# diff_1004400_769200# diff_1783200_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2762 diff_1803600_775200# diff_1004400_769200# diff_1803600_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2763 diff_1824000_775200# diff_1004400_769200# diff_1824000_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2764 diff_1844400_775200# diff_1004400_769200# diff_1844400_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2765 diff_1864800_775200# diff_1004400_769200# diff_1864800_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2766 diff_1885200_775200# diff_1004400_769200# diff_1885200_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2767 diff_1905600_775200# diff_1004400_769200# diff_1905600_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2768 diff_1926000_775200# diff_1004400_769200# diff_1926000_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2769 diff_1946400_775200# diff_1004400_769200# diff_1946400_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2770 diff_1966800_775200# diff_1004400_769200# diff_1966800_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2771 diff_1987200_775200# diff_1004400_769200# diff_1987200_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2772 diff_2007600_775200# diff_1004400_769200# diff_2007600_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2773 diff_2028000_775200# diff_1004400_769200# diff_2028000_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2774 diff_2048400_775200# diff_1004400_769200# diff_2048400_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2775 diff_2068800_775200# diff_1004400_769200# diff_2068800_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2776 diff_2089200_775200# diff_1004400_769200# diff_2089200_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2777 diff_2109600_775200# diff_1004400_769200# diff_2109600_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2778 diff_2130000_775200# diff_1004400_769200# diff_2130000_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2779 diff_2150400_775200# diff_1004400_769200# diff_2150400_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2780 diff_2170800_775200# diff_1004400_769200# diff_2170800_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2781 diff_2191200_775200# diff_1004400_769200# diff_2191200_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2782 diff_2211600_775200# diff_1004400_769200# diff_2211600_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2783 diff_2232000_775200# diff_1004400_769200# diff_2232000_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2784 diff_2252400_775200# diff_1004400_769200# diff_2252400_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2785 diff_2272800_775200# diff_1004400_769200# diff_2272800_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2786 diff_2293200_775200# diff_1004400_769200# diff_2293200_752400# GND efet w=10800 l=7200
+ ad=1.1376e+08 pd=43200 as=1.6848e+08 ps=52800 
M2787 GND diff_2526000_1243200# diff_2431200_979200# GND efet w=122400 l=6000
+ ad=0 pd=0 as=1.69776e+09 ps=331200 
M2788 Vdd Vdd diff_1124400_1153200# GND efet w=7200 l=14400
+ ad=0 pd=0 as=0 ps=0 
M2789 Vdd Vdd diff_2431200_979200# GND efet w=7200 l=14400
+ ad=0 pd=0 as=0 ps=0 
M2790 diff_2738400_1228800# diff_2722800_844800# diff_2530800_1201200# GND efet w=19200 l=6000
+ ad=5.8752e+08 pd=139200 as=2.736e+08 ps=67200 
M2791 Vdd Vdd diff_1124400_963600# GND efet w=7200 l=14400
+ ad=0 pd=0 as=1.77552e+09 ps=321600 
M2792 diff_1124400_963600# diff_2530800_1201200# GND GND efet w=122400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2793 GND diff_2530800_1178400# diff_2361600_427200# GND efet w=122400 l=6000
+ ad=0 pd=0 as=2.0016e+09 ps=331200 
M2794 Vdd Vdd diff_2361600_427200# GND efet w=7200 l=14400
+ ad=0 pd=0 as=0 ps=0 
M2795 Vdd Vdd diff_2384400_427200# GND efet w=7200 l=14400
+ ad=0 pd=0 as=1.99008e+09 ps=326400 
M2796 diff_2774400_1308000# Vdd Vdd GND efet w=8400 l=33600
+ ad=0 pd=0 as=0 ps=0 
M2797 diff_2818800_1292400# diff_2812800_1134000# diff_2774400_1308000# GND efet w=36000 l=6000
+ ad=3.456e+08 pd=91200 as=0 ps=0 
M2798 GND diff_2828400_1273200# diff_2818800_1292400# GND efet w=36000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2799 Vdd Vdd Vdd GND efet w=1200 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2800 Vdd Vdd Vdd GND efet w=1200 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2801 Vdd Vdd diff_2774400_1189200# GND efet w=8400 l=33600
+ ad=0 pd=0 as=1.1808e+09 ps=211200 
M2802 diff_2738400_1228800# diff_2710800_1356000# diff_2530800_1178400# GND efet w=21600 l=6000
+ ad=0 pd=0 as=3.3408e+08 ps=74400 
M2803 diff_2774400_1189200# clk2 diff_2738400_1228800# GND efet w=21600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2804 diff_2841600_1227600# diff_2828400_1273200# diff_2774400_1189200# GND efet w=34800 l=6000
+ ad=3.3408e+08 pd=88800 as=0 ps=0 
M2805 GND diff_2812800_1003200# diff_2841600_1227600# GND efet w=34800 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2806 GND diff_2828400_1086000# diff_2818800_1136400# GND efet w=36000 l=6000
+ ad=0 pd=0 as=9.8784e+08 ps=199200 
M2807 diff_2738400_1114800# diff_2710800_1356000# diff_2530800_1132800# GND efet w=19200 l=6000
+ ad=5.6592e+08 pd=136800 as=2.736e+08 ps=67200 
M2808 diff_2774400_1153200# clk2 diff_2738400_1114800# GND efet w=19200 l=6000
+ ad=8.9568e+08 pd=153600 as=0 ps=0 
M2809 diff_2384400_427200# diff_2530800_1132800# GND GND efet w=122400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2810 GND diff_2532000_1111200# diff_1011600_1153200# GND efet w=122400 l=6000
+ ad=0 pd=0 as=1.88064e+09 ps=324000 
M2811 diff_2738400_1114800# diff_2722800_844800# diff_2532000_1111200# GND efet w=20400 l=6000
+ ad=0 pd=0 as=2.9088e+08 ps=69600 
M2812 Vdd Vdd diff_1011600_1153200# GND efet w=7200 l=14400
+ ad=0 pd=0 as=0 ps=0 
M2813 diff_2738400_1077600# diff_2722800_844800# diff_2530800_1058400# GND efet w=19200 l=6000
+ ad=5.5008e+08 pd=134400 as=2.736e+08 ps=67200 
M2814 Vdd Vdd diff_1014000_962400# GND efet w=7200 l=14400
+ ad=0 pd=0 as=1.90944e+09 ps=324000 
M2815 diff_1014000_962400# diff_2530800_1058400# GND GND efet w=122400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2816 GND diff_2530800_1035600# diff_2413200_996000# GND efet w=122400 l=6000
+ ad=0 pd=0 as=1.94256e+09 ps=324000 
M2817 Vdd Vdd diff_2413200_996000# GND efet w=7200 l=14400
+ ad=0 pd=0 as=0 ps=0 
M2818 Vdd Vdd diff_2469600_912000# GND efet w=7200 l=14400
+ ad=0 pd=0 as=1.9512e+09 ps=326400 
M2819 diff_2469600_912000# diff_2530800_991200# GND GND efet w=122400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2820 GND diff_2530800_968400# diff_1033200_919200# GND efet w=122400 l=6000
+ ad=0 pd=0 as=1.85184e+09 ps=326400 
M2821 diff_2774400_1153200# Vdd Vdd GND efet w=7200 l=33600
+ ad=0 pd=0 as=0 ps=0 
M2822 diff_2818800_1136400# diff_2812800_1134000# diff_2774400_1153200# GND efet w=36000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2823 diff_2865600_1124400# diff_2812800_1003200# diff_2774400_1040400# GND efet w=37200 l=6000
+ ad=4.0176e+08 pd=96000 as=1.18656e+09 ps=216000 
M2824 GND diff_2828400_1086000# diff_2865600_1124400# GND efet w=37200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2825 Vdd Vdd Vdd GND efet w=1800 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2826 Vdd Vdd Vdd GND efet w=1800 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2827 Vdd Vdd diff_2774400_1040400# GND efet w=7200 l=33600
+ ad=0 pd=0 as=0 ps=0 
M2828 diff_2738400_1077600# diff_2710800_1356000# diff_2530800_1035600# GND efet w=19200 l=6000
+ ad=0 pd=0 as=2.736e+08 ps=67200 
M2829 diff_2774400_1040400# clk2 diff_2738400_1077600# GND efet w=19200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2830 diff_2738400_964800# diff_2710800_1356000# diff_2530800_991200# GND efet w=20400 l=6000
+ ad=5.8464e+08 pd=139200 as=2.9088e+08 ps=69600 
M2831 diff_2774400_1002000# clk2 diff_2738400_964800# GND efet w=20400 l=6000
+ ad=1.188e+09 pd=216000 as=0 ps=0 
M2832 d1 GND d1 GND efet w=177600 l=111600
+ ad=0 pd=0 as=0 ps=0 
M2833 GND diff_2828400_1086000# diff_2832000_1075200# GND efet w=63600 l=6000
+ ad=0 pd=0 as=6.1056e+08 ps=146400 
M2834 diff_2832000_1075200# diff_2812800_1003200# diff_2832000_1056000# GND efet w=63600 l=6000
+ ad=0 pd=0 as=1.92528e+09 ps=350400 
M2835 diff_919200_421200# diff_2812800_1003200# diff_2848800_992400# GND efet w=46800 l=6000
+ ad=-1.43801e+09 pd=600000 as=4.4928e+08 ps=112800 
M2836 diff_2738400_964800# diff_2722800_844800# diff_2530800_968400# GND efet w=20400 l=6000
+ ad=0 pd=0 as=2.9088e+08 ps=69600 
M2837 Vdd Vdd diff_1033200_919200# GND efet w=6000 l=14400
+ ad=0 pd=0 as=0 ps=0 
M2838 Vdd Vdd diff_1063200_940800# GND efet w=6000 l=14400
+ ad=0 pd=0 as=1.764e+09 ps=324000 
M2839 diff_2738400_926400# diff_2722800_844800# diff_2529600_915600# GND efet w=21600 l=6000
+ ad=6.0048e+08 pd=141600 as=3.0816e+08 ps=72000 
M2840 diff_1063200_940800# diff_2529600_915600# GND GND efet w=121200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2841 GND diff_2529600_894000# diff_2451600_979200# GND efet w=121200 l=6000
+ ad=0 pd=0 as=1.96272e+09 ps=324000 
M2842 Vdd Vdd diff_2451600_979200# GND efet w=8400 l=14400
+ ad=0 pd=0 as=0 ps=0 
M2843 Vdd Vdd Vdd GND efet w=6000 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2844 diff_1008000_752400# diff_1004400_746400# diff_1008000_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2845 diff_1028400_752400# diff_1004400_746400# diff_1028400_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2846 diff_1048800_752400# diff_1004400_746400# diff_1048800_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2847 diff_1069200_752400# diff_1004400_746400# diff_1069200_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2848 diff_1089600_752400# diff_1004400_746400# diff_1089600_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2849 diff_1110000_752400# diff_1004400_746400# diff_1110000_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2850 diff_1130400_752400# diff_1004400_746400# diff_1130400_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2851 diff_1150800_752400# diff_1004400_746400# diff_1150800_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2852 diff_1171200_752400# diff_1004400_746400# diff_1171200_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2853 diff_1191600_752400# diff_1004400_746400# diff_1191600_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2854 diff_1212000_752400# diff_1004400_746400# diff_1212000_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2855 diff_1232400_752400# diff_1004400_746400# diff_1232400_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2856 diff_1252800_752400# diff_1004400_746400# diff_1252800_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2857 diff_1273200_752400# diff_1004400_746400# diff_1273200_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2858 diff_1293600_752400# diff_1004400_746400# diff_1293600_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2859 diff_1314000_752400# diff_1004400_746400# diff_1314000_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2860 diff_1334400_752400# diff_1004400_746400# diff_1334400_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2861 diff_1354800_752400# diff_1004400_746400# diff_1354800_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2862 diff_1375200_752400# diff_1004400_746400# diff_1375200_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2863 diff_1395600_752400# diff_1004400_746400# diff_1395600_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2864 diff_1416000_752400# diff_1004400_746400# diff_1416000_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2865 diff_1436400_752400# diff_1004400_746400# diff_1436400_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2866 diff_1456800_752400# diff_1004400_746400# diff_1456800_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2867 diff_1477200_752400# diff_1004400_746400# diff_1477200_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2868 diff_1497600_752400# diff_1004400_746400# diff_1497600_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2869 diff_1518000_752400# diff_1004400_746400# diff_1518000_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2870 diff_1538400_752400# diff_1004400_746400# diff_1538400_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2871 diff_1558800_752400# diff_1004400_746400# diff_1558800_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2872 diff_1579200_752400# diff_1004400_746400# diff_1579200_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2873 diff_1599600_752400# diff_1004400_746400# diff_1599600_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2874 diff_1620000_752400# diff_1004400_746400# diff_1620000_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2875 diff_1640400_752400# diff_1004400_746400# diff_1640400_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2876 diff_1660800_752400# diff_1004400_746400# diff_1660800_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2877 diff_1681200_752400# diff_1004400_746400# diff_1681200_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2878 diff_1701600_752400# diff_1004400_746400# diff_1701600_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2879 diff_1722000_752400# diff_1004400_746400# diff_1722000_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2880 diff_1742400_752400# diff_1004400_746400# diff_1742400_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2881 diff_1762800_752400# diff_1004400_746400# diff_1762800_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2882 diff_1783200_752400# diff_1004400_746400# diff_1783200_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2883 diff_1803600_752400# diff_1004400_746400# diff_1803600_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2884 diff_1824000_752400# diff_1004400_746400# diff_1824000_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2885 diff_1844400_752400# diff_1004400_746400# diff_1844400_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2886 diff_1864800_752400# diff_1004400_746400# diff_1864800_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2887 diff_1885200_752400# diff_1004400_746400# diff_1885200_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2888 diff_1905600_752400# diff_1004400_746400# diff_1905600_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2889 diff_1926000_752400# diff_1004400_746400# diff_1926000_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2890 diff_1946400_752400# diff_1004400_746400# diff_1946400_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2891 diff_1966800_752400# diff_1004400_746400# diff_1966800_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2892 diff_1987200_752400# diff_1004400_746400# diff_1987200_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2893 diff_2007600_752400# diff_1004400_746400# diff_2007600_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2894 diff_2028000_752400# diff_1004400_746400# diff_2028000_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2895 diff_2048400_752400# diff_1004400_746400# diff_2048400_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2896 diff_2068800_752400# diff_1004400_746400# diff_2068800_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2897 diff_2089200_752400# diff_1004400_746400# diff_2089200_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2898 diff_2109600_752400# diff_1004400_746400# diff_2109600_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2899 diff_2130000_752400# diff_1004400_746400# diff_2130000_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2900 diff_2150400_752400# diff_1004400_746400# diff_2150400_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2901 diff_2170800_752400# diff_1004400_746400# diff_2170800_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2902 diff_2191200_752400# diff_1004400_746400# diff_2191200_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2903 diff_2211600_752400# diff_1004400_746400# diff_2211600_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2904 diff_2232000_752400# diff_1004400_746400# diff_2232000_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2905 diff_2252400_752400# diff_1004400_746400# diff_2252400_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2906 diff_2272800_752400# diff_1004400_746400# diff_2272800_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2907 diff_2293200_752400# diff_1004400_746400# diff_2293200_730800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2908 diff_1004400_769200# Vdd Vdd GND efet w=6000 l=13200
+ ad=9.4032e+08 pd=261600 as=0 ps=0 
M2909 Vdd Vdd Vdd GND efet w=2400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2910 Vdd Vdd Vdd GND efet w=1200 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2911 diff_866400_691200# Vdd Vdd GND efet w=7200 l=50400
+ ad=6.2064e+08 pd=148800 as=0 ps=0 
M2912 diff_411600_867600# diff_840000_375600# GND GND efet w=21600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2913 GND diff_866400_691200# diff_411600_867600# GND efet w=22800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2914 diff_1008000_730800# diff_1004400_724800# diff_1008000_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2915 diff_1028400_730800# diff_1004400_724800# diff_1028400_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2916 diff_1048800_730800# diff_1004400_724800# diff_1048800_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2917 diff_1069200_730800# diff_1004400_724800# diff_1069200_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2918 diff_1089600_730800# diff_1004400_724800# diff_1089600_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2919 diff_1110000_730800# diff_1004400_724800# diff_1110000_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2920 diff_1130400_730800# diff_1004400_724800# diff_1130400_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2921 diff_1150800_730800# diff_1004400_724800# diff_1150800_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2922 diff_1171200_730800# diff_1004400_724800# diff_1171200_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2923 diff_1191600_730800# diff_1004400_724800# diff_1191600_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2924 diff_1212000_730800# diff_1004400_724800# diff_1212000_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2925 diff_1232400_730800# diff_1004400_724800# diff_1232400_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2926 diff_1252800_730800# diff_1004400_724800# diff_1252800_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2927 diff_1273200_730800# diff_1004400_724800# diff_1273200_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2928 diff_1293600_730800# diff_1004400_724800# diff_1293600_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2929 diff_1314000_730800# diff_1004400_724800# diff_1314000_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2930 diff_1334400_730800# diff_1004400_724800# diff_1334400_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2931 diff_1354800_730800# diff_1004400_724800# diff_1354800_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2932 diff_1375200_730800# diff_1004400_724800# diff_1375200_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2933 diff_1395600_730800# diff_1004400_724800# diff_1395600_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2934 diff_1416000_730800# diff_1004400_724800# diff_1416000_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2935 diff_1436400_730800# diff_1004400_724800# diff_1436400_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2936 diff_1456800_730800# diff_1004400_724800# diff_1456800_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2937 diff_1477200_730800# diff_1004400_724800# diff_1477200_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2938 diff_1497600_730800# diff_1004400_724800# diff_1497600_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2939 diff_1518000_730800# diff_1004400_724800# diff_1518000_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2940 diff_1538400_730800# diff_1004400_724800# diff_1538400_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2941 diff_1558800_730800# diff_1004400_724800# diff_1558800_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2942 diff_1579200_730800# diff_1004400_724800# diff_1579200_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2943 diff_1599600_730800# diff_1004400_724800# diff_1599600_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2944 diff_1620000_730800# diff_1004400_724800# diff_1620000_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2945 diff_1640400_730800# diff_1004400_724800# diff_1640400_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2946 diff_1660800_730800# diff_1004400_724800# diff_1660800_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2947 diff_1681200_730800# diff_1004400_724800# diff_1681200_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2948 diff_1701600_730800# diff_1004400_724800# diff_1701600_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2949 diff_1722000_730800# diff_1004400_724800# diff_1722000_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2950 diff_1742400_730800# diff_1004400_724800# diff_1742400_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2951 diff_1762800_730800# diff_1004400_724800# diff_1762800_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2952 diff_1783200_730800# diff_1004400_724800# diff_1783200_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2953 diff_1803600_730800# diff_1004400_724800# diff_1803600_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2954 diff_1824000_730800# diff_1004400_724800# diff_1824000_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2955 diff_1844400_730800# diff_1004400_724800# diff_1844400_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2956 diff_1864800_730800# diff_1004400_724800# diff_1864800_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2957 diff_1885200_730800# diff_1004400_724800# diff_1885200_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2958 diff_1905600_730800# diff_1004400_724800# diff_1905600_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2959 diff_1926000_730800# diff_1004400_724800# diff_1926000_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2960 diff_1946400_730800# diff_1004400_724800# diff_1946400_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2961 diff_1966800_730800# diff_1004400_724800# diff_1966800_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2962 diff_1987200_730800# diff_1004400_724800# diff_1987200_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2963 diff_2007600_730800# diff_1004400_724800# diff_2007600_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2964 diff_2028000_730800# diff_1004400_724800# diff_2028000_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2965 diff_2048400_730800# diff_1004400_724800# diff_2048400_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2966 diff_2068800_730800# diff_1004400_724800# diff_2068800_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2967 diff_2089200_730800# diff_1004400_724800# diff_2089200_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2968 diff_2109600_730800# diff_1004400_724800# diff_2109600_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2969 diff_2130000_730800# diff_1004400_724800# diff_2130000_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2970 diff_2150400_730800# diff_1004400_724800# diff_2150400_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2971 diff_2170800_730800# diff_1004400_724800# diff_2170800_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2972 diff_2191200_730800# diff_1004400_724800# diff_2191200_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2973 diff_2211600_730800# diff_1004400_724800# diff_2211600_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2974 diff_2232000_730800# diff_1004400_724800# diff_2232000_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2975 diff_2252400_730800# diff_1004400_724800# diff_2252400_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2976 diff_2272800_730800# diff_1004400_724800# diff_2272800_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2977 diff_2293200_730800# diff_1004400_724800# diff_2293200_708000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M2978 Vdd Vdd diff_1004400_702000# GND efet w=6000 l=12000
+ ad=0 pd=0 as=8.7264e+08 ps=228000 
M2979 diff_2367600_696000# diff_2361600_427200# diff_1004400_702000# GND efet w=86400 l=6000
+ ad=-6.48887e+08 pd=727200 as=0 ps=0 
M2980 diff_866400_691200# diff_866400_691200# diff_866400_691200# GND efet w=1800 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2981 diff_866400_691200# diff_866400_691200# diff_866400_691200# GND efet w=2400 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2982 GND diff_904800_656400# diff_866400_691200# GND efet w=20400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2983 diff_1008000_708000# diff_1004400_702000# diff_1008000_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2984 diff_1028400_708000# diff_1004400_702000# diff_1028400_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2985 diff_1048800_708000# diff_1004400_702000# diff_1048800_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2986 diff_1069200_708000# diff_1004400_702000# diff_1069200_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2987 diff_1089600_708000# diff_1004400_702000# diff_1089600_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2988 diff_1110000_708000# diff_1004400_702000# diff_1110000_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2989 diff_1130400_708000# diff_1004400_702000# diff_1130400_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2990 diff_1150800_708000# diff_1004400_702000# diff_1150800_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2991 diff_1171200_708000# diff_1004400_702000# diff_1171200_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2992 diff_1191600_708000# diff_1004400_702000# diff_1191600_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2993 diff_1212000_708000# diff_1004400_702000# diff_1212000_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2994 diff_1232400_708000# diff_1004400_702000# diff_1232400_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2995 diff_1252800_708000# diff_1004400_702000# diff_1252800_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2996 diff_1273200_708000# diff_1004400_702000# diff_1273200_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2997 diff_1293600_708000# diff_1004400_702000# diff_1293600_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2998 diff_1314000_708000# diff_1004400_702000# diff_1314000_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M2999 diff_1334400_708000# diff_1004400_702000# diff_1334400_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3000 diff_1354800_708000# diff_1004400_702000# diff_1354800_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3001 diff_1375200_708000# diff_1004400_702000# diff_1375200_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3002 diff_1395600_708000# diff_1004400_702000# diff_1395600_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3003 diff_1416000_708000# diff_1004400_702000# diff_1416000_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3004 diff_1436400_708000# diff_1004400_702000# diff_1436400_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3005 diff_1456800_708000# diff_1004400_702000# diff_1456800_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3006 diff_1477200_708000# diff_1004400_702000# diff_1477200_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3007 diff_1497600_708000# diff_1004400_702000# diff_1497600_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3008 diff_1518000_708000# diff_1004400_702000# diff_1518000_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3009 diff_1538400_708000# diff_1004400_702000# diff_1538400_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3010 diff_1558800_708000# diff_1004400_702000# diff_1558800_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3011 diff_1579200_708000# diff_1004400_702000# diff_1579200_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3012 diff_1599600_708000# diff_1004400_702000# diff_1599600_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3013 diff_1620000_708000# diff_1004400_702000# diff_1620000_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3014 diff_1640400_708000# diff_1004400_702000# diff_1640400_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3015 diff_1660800_708000# diff_1004400_702000# diff_1660800_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3016 diff_1681200_708000# diff_1004400_702000# diff_1681200_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3017 diff_1701600_708000# diff_1004400_702000# diff_1701600_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3018 diff_1722000_708000# diff_1004400_702000# diff_1722000_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3019 diff_1742400_708000# diff_1004400_702000# diff_1742400_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3020 diff_1762800_708000# diff_1004400_702000# diff_1762800_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3021 diff_1783200_708000# diff_1004400_702000# diff_1783200_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3022 diff_1803600_708000# diff_1004400_702000# diff_1803600_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3023 diff_1824000_708000# diff_1004400_702000# diff_1824000_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3024 diff_1844400_708000# diff_1004400_702000# diff_1844400_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3025 diff_1864800_708000# diff_1004400_702000# diff_1864800_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3026 diff_1885200_708000# diff_1004400_702000# diff_1885200_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3027 diff_1905600_708000# diff_1004400_702000# diff_1905600_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3028 diff_1926000_708000# diff_1004400_702000# diff_1926000_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3029 diff_1946400_708000# diff_1004400_702000# diff_1946400_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3030 diff_1966800_708000# diff_1004400_702000# diff_1966800_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3031 diff_1987200_708000# diff_1004400_702000# diff_1987200_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3032 diff_2007600_708000# diff_1004400_702000# diff_2007600_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3033 diff_2028000_708000# diff_1004400_702000# diff_2028000_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3034 diff_2048400_708000# diff_1004400_702000# diff_2048400_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3035 diff_2068800_708000# diff_1004400_702000# diff_2068800_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3036 diff_2089200_708000# diff_1004400_702000# diff_2089200_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3037 diff_2109600_708000# diff_1004400_702000# diff_2109600_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3038 diff_2130000_708000# diff_1004400_702000# diff_2130000_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3039 diff_2150400_708000# diff_1004400_702000# diff_2150400_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3040 diff_2170800_708000# diff_1004400_702000# diff_2170800_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3041 diff_2191200_708000# diff_1004400_702000# diff_2191200_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3042 diff_2211600_708000# diff_1004400_702000# diff_2211600_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3043 diff_2232000_708000# diff_1004400_702000# diff_2232000_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3044 diff_2252400_708000# diff_1004400_702000# diff_2252400_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3045 diff_2272800_708000# diff_1004400_702000# diff_2272800_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3046 diff_2293200_708000# diff_1004400_702000# diff_2293200_686400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3047 diff_1004400_769200# diff_2384400_427200# diff_2367600_696000# GND efet w=74400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3048 diff_1004400_746400# Vdd Vdd GND efet w=7200 l=13200
+ ad=1.0368e+09 pd=249600 as=0 ps=0 
M3049 Vdd Vdd diff_1004400_724800# GND efet w=7200 l=10800
+ ad=0 pd=0 as=1.05264e+09 ps=225600 
M3050 diff_2367600_696000# diff_2413200_996000# diff_1004400_724800# GND efet w=85200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3051 diff_1008000_686400# diff_1004400_680400# diff_1008000_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3052 diff_1028400_686400# diff_1004400_680400# diff_1028400_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3053 diff_1048800_686400# diff_1004400_680400# diff_1048800_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3054 diff_1069200_686400# diff_1004400_680400# diff_1069200_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3055 diff_1089600_686400# diff_1004400_680400# diff_1089600_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3056 diff_1110000_686400# diff_1004400_680400# diff_1110000_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3057 diff_1130400_686400# diff_1004400_680400# diff_1130400_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3058 diff_1150800_686400# diff_1004400_680400# diff_1150800_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3059 diff_1171200_686400# diff_1004400_680400# diff_1171200_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3060 diff_1191600_686400# diff_1004400_680400# diff_1191600_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3061 diff_1212000_686400# diff_1004400_680400# diff_1212000_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3062 diff_1232400_686400# diff_1004400_680400# diff_1232400_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3063 diff_1252800_686400# diff_1004400_680400# diff_1252800_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3064 diff_1273200_686400# diff_1004400_680400# diff_1273200_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3065 diff_1293600_686400# diff_1004400_680400# diff_1293600_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3066 diff_1314000_686400# diff_1004400_680400# diff_1314000_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3067 diff_1334400_686400# diff_1004400_680400# diff_1334400_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3068 diff_1354800_686400# diff_1004400_680400# diff_1354800_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3069 diff_1375200_686400# diff_1004400_680400# diff_1375200_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3070 diff_1395600_686400# diff_1004400_680400# diff_1395600_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3071 diff_1416000_686400# diff_1004400_680400# diff_1416000_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3072 diff_1436400_686400# diff_1004400_680400# diff_1436400_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3073 diff_1456800_686400# diff_1004400_680400# diff_1456800_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3074 diff_1477200_686400# diff_1004400_680400# diff_1477200_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3075 diff_1497600_686400# diff_1004400_680400# diff_1497600_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3076 diff_1518000_686400# diff_1004400_680400# diff_1518000_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3077 diff_1538400_686400# diff_1004400_680400# diff_1538400_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3078 diff_1558800_686400# diff_1004400_680400# diff_1558800_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3079 diff_1579200_686400# diff_1004400_680400# diff_1579200_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3080 diff_1599600_686400# diff_1004400_680400# diff_1599600_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3081 diff_1620000_686400# diff_1004400_680400# diff_1620000_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3082 diff_1640400_686400# diff_1004400_680400# diff_1640400_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3083 diff_1660800_686400# diff_1004400_680400# diff_1660800_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3084 diff_1681200_686400# diff_1004400_680400# diff_1681200_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3085 diff_1701600_686400# diff_1004400_680400# diff_1701600_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3086 diff_1722000_686400# diff_1004400_680400# diff_1722000_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3087 diff_1742400_686400# diff_1004400_680400# diff_1742400_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3088 diff_1762800_686400# diff_1004400_680400# diff_1762800_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3089 diff_1783200_686400# diff_1004400_680400# diff_1783200_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3090 diff_1803600_686400# diff_1004400_680400# diff_1803600_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3091 diff_1824000_686400# diff_1004400_680400# diff_1824000_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3092 diff_1844400_686400# diff_1004400_680400# diff_1844400_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3093 diff_1864800_686400# diff_1004400_680400# diff_1864800_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3094 diff_1885200_686400# diff_1004400_680400# diff_1885200_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3095 diff_1905600_686400# diff_1004400_680400# diff_1905600_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3096 diff_1926000_686400# diff_1004400_680400# diff_1926000_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3097 diff_1946400_686400# diff_1004400_680400# diff_1946400_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3098 diff_1966800_686400# diff_1004400_680400# diff_1966800_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3099 diff_1987200_686400# diff_1004400_680400# diff_1987200_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3100 diff_2007600_686400# diff_1004400_680400# diff_2007600_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3101 diff_2028000_686400# diff_1004400_680400# diff_2028000_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3102 diff_2048400_686400# diff_1004400_680400# diff_2048400_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3103 diff_2068800_686400# diff_1004400_680400# diff_2068800_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3104 diff_2089200_686400# diff_1004400_680400# diff_2089200_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3105 diff_2109600_686400# diff_1004400_680400# diff_2109600_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3106 diff_2130000_686400# diff_1004400_680400# diff_2130000_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3107 diff_2150400_686400# diff_1004400_680400# diff_2150400_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3108 diff_2170800_686400# diff_1004400_680400# diff_2170800_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3109 diff_2191200_686400# diff_1004400_680400# diff_2191200_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3110 diff_2211600_686400# diff_1004400_680400# diff_2211600_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3111 diff_2232000_686400# diff_1004400_680400# diff_2232000_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3112 diff_2252400_686400# diff_1004400_680400# diff_2252400_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3113 diff_2272800_686400# diff_1004400_680400# diff_2272800_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3114 diff_2293200_686400# diff_1004400_680400# diff_2293200_663600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3115 diff_1004400_746400# diff_2431200_979200# diff_2367600_696000# GND efet w=79200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3116 diff_2367600_607200# diff_2361600_427200# diff_1004400_613200# GND efet w=88200 l=7200
+ ad=-2.41367e+08 pd=720000 as=8.4672e+08 ps=228000 
M3117 diff_891600_656400# clk2 Vdd GND efet w=12000 l=7200
+ ad=7.2e+07 pd=36000 as=0 ps=0 
M3118 diff_904800_656400# diff_897600_638400# diff_891600_656400# GND efet w=12000 l=7200
+ ad=4.608e+08 pd=100800 as=0 ps=0 
M3119 GND diff_338400_375600# diff_904800_656400# GND efet w=12000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3120 diff_1008000_663600# diff_1004400_657600# diff_1008000_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3121 diff_1028400_663600# diff_1004400_657600# diff_1028400_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3122 diff_1048800_663600# diff_1004400_657600# diff_1048800_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3123 diff_1069200_663600# diff_1004400_657600# diff_1069200_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3124 diff_1089600_663600# diff_1004400_657600# diff_1089600_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3125 diff_1110000_663600# diff_1004400_657600# diff_1110000_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3126 diff_1130400_663600# diff_1004400_657600# diff_1130400_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3127 diff_1150800_663600# diff_1004400_657600# diff_1150800_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3128 diff_1171200_663600# diff_1004400_657600# diff_1171200_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3129 diff_1191600_663600# diff_1004400_657600# diff_1191600_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3130 diff_1212000_663600# diff_1004400_657600# diff_1212000_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3131 diff_1232400_663600# diff_1004400_657600# diff_1232400_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3132 diff_1252800_663600# diff_1004400_657600# diff_1252800_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3133 diff_1273200_663600# diff_1004400_657600# diff_1273200_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3134 diff_1293600_663600# diff_1004400_657600# diff_1293600_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3135 diff_1314000_663600# diff_1004400_657600# diff_1314000_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3136 diff_1334400_663600# diff_1004400_657600# diff_1334400_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3137 diff_1354800_663600# diff_1004400_657600# diff_1354800_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3138 diff_1375200_663600# diff_1004400_657600# diff_1375200_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3139 diff_1395600_663600# diff_1004400_657600# diff_1395600_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3140 diff_1416000_663600# diff_1004400_657600# diff_1416000_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3141 diff_1436400_663600# diff_1004400_657600# diff_1436400_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3142 diff_1456800_663600# diff_1004400_657600# diff_1456800_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3143 diff_1477200_663600# diff_1004400_657600# diff_1477200_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3144 diff_1497600_663600# diff_1004400_657600# diff_1497600_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3145 diff_1518000_663600# diff_1004400_657600# diff_1518000_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3146 diff_1538400_663600# diff_1004400_657600# diff_1538400_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3147 diff_1558800_663600# diff_1004400_657600# diff_1558800_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3148 diff_1579200_663600# diff_1004400_657600# diff_1579200_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3149 diff_1599600_663600# diff_1004400_657600# diff_1599600_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3150 diff_1620000_663600# diff_1004400_657600# diff_1620000_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3151 diff_1640400_663600# diff_1004400_657600# diff_1640400_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3152 diff_1660800_663600# diff_1004400_657600# diff_1660800_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3153 diff_1681200_663600# diff_1004400_657600# diff_1681200_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3154 diff_1701600_663600# diff_1004400_657600# diff_1701600_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3155 diff_1722000_663600# diff_1004400_657600# diff_1722000_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3156 diff_1742400_663600# diff_1004400_657600# diff_1742400_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3157 diff_1762800_663600# diff_1004400_657600# diff_1762800_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3158 diff_1783200_663600# diff_1004400_657600# diff_1783200_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3159 diff_1803600_663600# diff_1004400_657600# diff_1803600_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3160 diff_1824000_663600# diff_1004400_657600# diff_1824000_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3161 diff_1844400_663600# diff_1004400_657600# diff_1844400_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3162 diff_1864800_663600# diff_1004400_657600# diff_1864800_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3163 diff_1885200_663600# diff_1004400_657600# diff_1885200_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3164 diff_1905600_663600# diff_1004400_657600# diff_1905600_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3165 diff_1926000_663600# diff_1004400_657600# diff_1926000_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3166 diff_1946400_663600# diff_1004400_657600# diff_1946400_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3167 diff_1966800_663600# diff_1004400_657600# diff_1966800_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3168 diff_1987200_663600# diff_1004400_657600# diff_1987200_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3169 diff_2007600_663600# diff_1004400_657600# diff_2007600_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3170 diff_2028000_663600# diff_1004400_657600# diff_2028000_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3171 diff_2048400_663600# diff_1004400_657600# diff_2048400_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3172 diff_2068800_663600# diff_1004400_657600# diff_2068800_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3173 diff_2089200_663600# diff_1004400_657600# diff_2089200_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3174 diff_2109600_663600# diff_1004400_657600# diff_2109600_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3175 diff_2130000_663600# diff_1004400_657600# diff_2130000_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3176 diff_2150400_663600# diff_1004400_657600# diff_2150400_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3177 diff_2170800_663600# diff_1004400_657600# diff_2170800_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3178 diff_2191200_663600# diff_1004400_657600# diff_2191200_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3179 diff_2211600_663600# diff_1004400_657600# diff_2211600_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3180 diff_2232000_663600# diff_1004400_657600# diff_2232000_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3181 diff_2252400_663600# diff_1004400_657600# diff_2252400_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3182 diff_2272800_663600# diff_1004400_657600# diff_2272800_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3183 diff_2293200_663600# diff_1004400_657600# diff_2293200_642000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3184 diff_1004400_680400# Vdd Vdd GND efet w=6000 l=13200
+ ad=9.4032e+08 pd=261600 as=0 ps=0 
M3185 diff_694800_762000# diff_746400_625200# GND GND efet w=12000 l=7200
+ ad=2.4768e+08 pd=69600 as=0 ps=0 
M3186 Vdd Vdd diff_694800_762000# GND efet w=7800 l=51000
+ ad=0 pd=0 as=0 ps=0 
M3187 diff_564000_475200# diff_564000_475200# diff_564000_475200# GND efet w=3000 l=3600
+ ad=1.12032e+09 pd=256800 as=0 ps=0 
M3188 diff_564000_475200# diff_564000_475200# diff_564000_475200# GND efet w=3000 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3189 Vdd Vdd diff_564000_475200# GND efet w=9600 l=16800
+ ad=0 pd=0 as=0 ps=0 
M3190 diff_1008000_642000# diff_1004400_636000# diff_1008000_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3191 diff_1028400_642000# diff_1004400_636000# diff_1028400_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3192 diff_1048800_642000# diff_1004400_636000# diff_1048800_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3193 diff_1069200_642000# diff_1004400_636000# diff_1069200_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3194 diff_1089600_642000# diff_1004400_636000# diff_1089600_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3195 diff_1110000_642000# diff_1004400_636000# diff_1110000_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3196 diff_1130400_642000# diff_1004400_636000# diff_1130400_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3197 diff_1150800_642000# diff_1004400_636000# diff_1150800_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3198 diff_1171200_642000# diff_1004400_636000# diff_1171200_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3199 diff_1191600_642000# diff_1004400_636000# diff_1191600_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3200 diff_1212000_642000# diff_1004400_636000# diff_1212000_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3201 diff_1232400_642000# diff_1004400_636000# diff_1232400_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3202 diff_1252800_642000# diff_1004400_636000# diff_1252800_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3203 diff_1273200_642000# diff_1004400_636000# diff_1273200_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3204 diff_1293600_642000# diff_1004400_636000# diff_1293600_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3205 diff_1314000_642000# diff_1004400_636000# diff_1314000_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3206 diff_1334400_642000# diff_1004400_636000# diff_1334400_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3207 diff_1354800_642000# diff_1004400_636000# diff_1354800_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3208 diff_1375200_642000# diff_1004400_636000# diff_1375200_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3209 diff_1395600_642000# diff_1004400_636000# diff_1395600_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3210 diff_1416000_642000# diff_1004400_636000# diff_1416000_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3211 diff_1436400_642000# diff_1004400_636000# diff_1436400_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3212 diff_1456800_642000# diff_1004400_636000# diff_1456800_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3213 diff_1477200_642000# diff_1004400_636000# diff_1477200_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3214 diff_1497600_642000# diff_1004400_636000# diff_1497600_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3215 diff_1518000_642000# diff_1004400_636000# diff_1518000_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3216 diff_1538400_642000# diff_1004400_636000# diff_1538400_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3217 diff_1558800_642000# diff_1004400_636000# diff_1558800_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3218 diff_1579200_642000# diff_1004400_636000# diff_1579200_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3219 diff_1599600_642000# diff_1004400_636000# diff_1599600_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3220 diff_1620000_642000# diff_1004400_636000# diff_1620000_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3221 diff_1640400_642000# diff_1004400_636000# diff_1640400_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3222 diff_1660800_642000# diff_1004400_636000# diff_1660800_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3223 diff_1681200_642000# diff_1004400_636000# diff_1681200_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3224 diff_1701600_642000# diff_1004400_636000# diff_1701600_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3225 diff_1722000_642000# diff_1004400_636000# diff_1722000_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3226 diff_1742400_642000# diff_1004400_636000# diff_1742400_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3227 diff_1762800_642000# diff_1004400_636000# diff_1762800_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3228 diff_1783200_642000# diff_1004400_636000# diff_1783200_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3229 diff_1803600_642000# diff_1004400_636000# diff_1803600_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3230 diff_1824000_642000# diff_1004400_636000# diff_1824000_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3231 diff_1844400_642000# diff_1004400_636000# diff_1844400_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3232 diff_1864800_642000# diff_1004400_636000# diff_1864800_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3233 diff_1885200_642000# diff_1004400_636000# diff_1885200_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3234 diff_1905600_642000# diff_1004400_636000# diff_1905600_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3235 diff_1926000_642000# diff_1004400_636000# diff_1926000_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3236 diff_1946400_642000# diff_1004400_636000# diff_1946400_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3237 diff_1966800_642000# diff_1004400_636000# diff_1966800_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3238 diff_1987200_642000# diff_1004400_636000# diff_1987200_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3239 diff_2007600_642000# diff_1004400_636000# diff_2007600_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3240 diff_2028000_642000# diff_1004400_636000# diff_2028000_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3241 diff_2048400_642000# diff_1004400_636000# diff_2048400_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3242 diff_2068800_642000# diff_1004400_636000# diff_2068800_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3243 diff_2089200_642000# diff_1004400_636000# diff_2089200_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3244 diff_2109600_642000# diff_1004400_636000# diff_2109600_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3245 diff_2130000_642000# diff_1004400_636000# diff_2130000_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3246 diff_2150400_642000# diff_1004400_636000# diff_2150400_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3247 diff_2170800_642000# diff_1004400_636000# diff_2170800_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3248 diff_2191200_642000# diff_1004400_636000# diff_2191200_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3249 diff_2211600_642000# diff_1004400_636000# diff_2211600_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3250 diff_2232000_642000# diff_1004400_636000# diff_2232000_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3251 diff_2252400_642000# diff_1004400_636000# diff_2252400_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3252 diff_2272800_642000# diff_1004400_636000# diff_2272800_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3253 diff_2293200_642000# diff_1004400_636000# diff_2293200_619200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3254 Vdd Vdd diff_1004400_613200# GND efet w=6000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M3255 Vdd Vdd diff_624000_475200# GND efet w=9600 l=16800
+ ad=0 pd=0 as=8.5104e+08 ps=189600 
M3256 Vdd Vdd Vdd GND efet w=4200 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3257 Vdd Vdd diff_694800_556800# GND efet w=7200 l=63600
+ ad=0 pd=0 as=8.6256e+08 ps=208800 
M3258 diff_694800_556800# cm diff_694800_493200# GND efet w=78000 l=7200
+ ad=0 pd=0 as=7.1424e+08 ps=172800 
M3259 diff_404400_470400# diff_338400_375600# Vdd GND efet w=13200 l=6000
+ ad=2.5344e+08 pd=64800 as=0 ps=0 
M3260 diff_475200_500400# clk2 diff_404400_470400# GND efet w=13200 l=7200
+ ad=1.1088e+08 pd=43200 as=0 ps=0 
M3261 diff_490800_500400# diff_478800_470400# diff_475200_500400# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3262 Vdd Vdd diff_691200_487200# GND efet w=8400 l=50400
+ ad=0 pd=0 as=1.02096e+09 ps=220800 
M3263 Vdd Vdd diff_756000_454800# GND efet w=7200 l=50400
+ ad=0 pd=0 as=4.7808e+08 ps=129600 
M3264 Vdd Vdd Vdd GND efet w=3600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3265 diff_897600_638400# Vdd Vdd GND efet w=7200 l=34800
+ ad=6.3792e+08 pd=163200 as=0 ps=0 
M3266 GND diff_694800_556800# diff_897600_638400# GND efet w=18000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3267 diff_897600_638400# diff_904800_769200# GND GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3268 GND diff_919200_421200# diff_897600_638400# GND efet w=18000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3269 diff_1008000_619200# diff_1004400_613200# diff_1008000_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3270 diff_1028400_619200# diff_1004400_613200# diff_1028400_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3271 diff_1048800_619200# diff_1004400_613200# diff_1048800_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3272 diff_1069200_619200# diff_1004400_613200# diff_1069200_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3273 diff_1089600_619200# diff_1004400_613200# diff_1089600_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3274 diff_1110000_619200# diff_1004400_613200# diff_1110000_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3275 diff_1130400_619200# diff_1004400_613200# diff_1130400_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3276 diff_1150800_619200# diff_1004400_613200# diff_1150800_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3277 diff_1171200_619200# diff_1004400_613200# diff_1171200_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3278 diff_1191600_619200# diff_1004400_613200# diff_1191600_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3279 diff_1212000_619200# diff_1004400_613200# diff_1212000_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3280 diff_1232400_619200# diff_1004400_613200# diff_1232400_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3281 diff_1252800_619200# diff_1004400_613200# diff_1252800_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3282 diff_1273200_619200# diff_1004400_613200# diff_1273200_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3283 diff_1293600_619200# diff_1004400_613200# diff_1293600_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3284 diff_1314000_619200# diff_1004400_613200# diff_1314000_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3285 diff_1334400_619200# diff_1004400_613200# diff_1334400_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3286 diff_1354800_619200# diff_1004400_613200# diff_1354800_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3287 diff_1375200_619200# diff_1004400_613200# diff_1375200_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3288 diff_1395600_619200# diff_1004400_613200# diff_1395600_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3289 diff_1416000_619200# diff_1004400_613200# diff_1416000_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3290 diff_1436400_619200# diff_1004400_613200# diff_1436400_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3291 diff_1456800_619200# diff_1004400_613200# diff_1456800_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3292 diff_1477200_619200# diff_1004400_613200# diff_1477200_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3293 diff_1497600_619200# diff_1004400_613200# diff_1497600_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3294 diff_1518000_619200# diff_1004400_613200# diff_1518000_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3295 diff_1538400_619200# diff_1004400_613200# diff_1538400_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3296 diff_1558800_619200# diff_1004400_613200# diff_1558800_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3297 diff_1579200_619200# diff_1004400_613200# diff_1579200_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3298 diff_1599600_619200# diff_1004400_613200# diff_1599600_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3299 diff_1620000_619200# diff_1004400_613200# diff_1620000_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3300 diff_1640400_619200# diff_1004400_613200# diff_1640400_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3301 diff_1660800_619200# diff_1004400_613200# diff_1660800_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3302 diff_1681200_619200# diff_1004400_613200# diff_1681200_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3303 diff_1701600_619200# diff_1004400_613200# diff_1701600_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3304 diff_1722000_619200# diff_1004400_613200# diff_1722000_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3305 diff_1742400_619200# diff_1004400_613200# diff_1742400_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3306 diff_1762800_619200# diff_1004400_613200# diff_1762800_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3307 diff_1783200_619200# diff_1004400_613200# diff_1783200_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3308 diff_1803600_619200# diff_1004400_613200# diff_1803600_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3309 diff_1824000_619200# diff_1004400_613200# diff_1824000_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3310 diff_1844400_619200# diff_1004400_613200# diff_1844400_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3311 diff_1864800_619200# diff_1004400_613200# diff_1864800_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3312 diff_1885200_619200# diff_1004400_613200# diff_1885200_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3313 diff_1905600_619200# diff_1004400_613200# diff_1905600_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3314 diff_1926000_619200# diff_1004400_613200# diff_1926000_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3315 diff_1946400_619200# diff_1004400_613200# diff_1946400_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3316 diff_1966800_619200# diff_1004400_613200# diff_1966800_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3317 diff_1987200_619200# diff_1004400_613200# diff_1987200_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3318 diff_2007600_619200# diff_1004400_613200# diff_2007600_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3319 diff_2028000_619200# diff_1004400_613200# diff_2028000_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3320 diff_2048400_619200# diff_1004400_613200# diff_2048400_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3321 diff_2068800_619200# diff_1004400_613200# diff_2068800_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3322 diff_2089200_619200# diff_1004400_613200# diff_2089200_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3323 diff_2109600_619200# diff_1004400_613200# diff_2109600_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3324 diff_2130000_619200# diff_1004400_613200# diff_2130000_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3325 diff_2150400_619200# diff_1004400_613200# diff_2150400_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3326 diff_2170800_619200# diff_1004400_613200# diff_2170800_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3327 diff_2191200_619200# diff_1004400_613200# diff_2191200_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3328 diff_2211600_619200# diff_1004400_613200# diff_2211600_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3329 diff_2232000_619200# diff_1004400_613200# diff_2232000_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3330 diff_2252400_619200# diff_1004400_613200# diff_2252400_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3331 diff_2272800_619200# diff_1004400_613200# diff_2272800_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3332 diff_2293200_619200# diff_1004400_613200# diff_2293200_597600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3333 Vdd Vdd diff_810000_510000# GND efet w=7200 l=51600
+ ad=0 pd=0 as=6.4368e+08 ps=172800 
M3334 diff_1004400_680400# diff_2384400_427200# diff_2367600_607200# GND efet w=74400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3335 diff_1004400_657600# Vdd Vdd GND efet w=7200 l=12000
+ ad=1.0368e+09 pd=249600 as=0 ps=0 
M3336 Vdd Vdd diff_1004400_636000# GND efet w=7200 l=10800
+ ad=0 pd=0 as=1.05984e+09 ps=225600 
M3337 diff_2367600_607200# diff_2413200_996000# diff_1004400_636000# GND efet w=84000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3338 diff_1008000_597600# diff_1004400_591600# diff_1008000_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3339 diff_1028400_597600# diff_1004400_591600# diff_1028400_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3340 diff_1048800_597600# diff_1004400_591600# diff_1048800_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3341 diff_1069200_597600# diff_1004400_591600# diff_1069200_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3342 diff_1089600_597600# diff_1004400_591600# diff_1089600_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3343 diff_1110000_597600# diff_1004400_591600# diff_1110000_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3344 diff_1130400_597600# diff_1004400_591600# diff_1130400_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3345 diff_1150800_597600# diff_1004400_591600# diff_1150800_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3346 diff_1171200_597600# diff_1004400_591600# diff_1171200_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3347 diff_1191600_597600# diff_1004400_591600# diff_1191600_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3348 diff_1212000_597600# diff_1004400_591600# diff_1212000_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3349 diff_1232400_597600# diff_1004400_591600# diff_1232400_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3350 diff_1252800_597600# diff_1004400_591600# diff_1252800_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3351 diff_1273200_597600# diff_1004400_591600# diff_1273200_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3352 diff_1293600_597600# diff_1004400_591600# diff_1293600_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3353 diff_1314000_597600# diff_1004400_591600# diff_1314000_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3354 diff_1334400_597600# diff_1004400_591600# diff_1334400_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3355 diff_1354800_597600# diff_1004400_591600# diff_1354800_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3356 diff_1375200_597600# diff_1004400_591600# diff_1375200_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3357 diff_1395600_597600# diff_1004400_591600# diff_1395600_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3358 diff_1416000_597600# diff_1004400_591600# diff_1416000_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3359 diff_1436400_597600# diff_1004400_591600# diff_1436400_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3360 diff_1456800_597600# diff_1004400_591600# diff_1456800_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3361 diff_1477200_597600# diff_1004400_591600# diff_1477200_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3362 diff_1497600_597600# diff_1004400_591600# diff_1497600_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3363 diff_1518000_597600# diff_1004400_591600# diff_1518000_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3364 diff_1538400_597600# diff_1004400_591600# diff_1538400_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3365 diff_1558800_597600# diff_1004400_591600# diff_1558800_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3366 diff_1579200_597600# diff_1004400_591600# diff_1579200_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3367 diff_1599600_597600# diff_1004400_591600# diff_1599600_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3368 diff_1620000_597600# diff_1004400_591600# diff_1620000_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3369 diff_1640400_597600# diff_1004400_591600# diff_1640400_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3370 diff_1660800_597600# diff_1004400_591600# diff_1660800_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3371 diff_1681200_597600# diff_1004400_591600# diff_1681200_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3372 diff_1701600_597600# diff_1004400_591600# diff_1701600_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3373 diff_1722000_597600# diff_1004400_591600# diff_1722000_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3374 diff_1742400_597600# diff_1004400_591600# diff_1742400_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3375 diff_1762800_597600# diff_1004400_591600# diff_1762800_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3376 diff_1783200_597600# diff_1004400_591600# diff_1783200_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3377 diff_1803600_597600# diff_1004400_591600# diff_1803600_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3378 diff_1824000_597600# diff_1004400_591600# diff_1824000_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3379 diff_1844400_597600# diff_1004400_591600# diff_1844400_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3380 diff_1864800_597600# diff_1004400_591600# diff_1864800_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3381 diff_1885200_597600# diff_1004400_591600# diff_1885200_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3382 diff_1905600_597600# diff_1004400_591600# diff_1905600_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3383 diff_1926000_597600# diff_1004400_591600# diff_1926000_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3384 diff_1946400_597600# diff_1004400_591600# diff_1946400_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3385 diff_1966800_597600# diff_1004400_591600# diff_1966800_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3386 diff_1987200_597600# diff_1004400_591600# diff_1987200_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3387 diff_2007600_597600# diff_1004400_591600# diff_2007600_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3388 diff_2028000_597600# diff_1004400_591600# diff_2028000_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3389 diff_2048400_597600# diff_1004400_591600# diff_2048400_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3390 diff_2068800_597600# diff_1004400_591600# diff_2068800_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3391 diff_2089200_597600# diff_1004400_591600# diff_2089200_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3392 diff_2109600_597600# diff_1004400_591600# diff_2109600_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3393 diff_2130000_597600# diff_1004400_591600# diff_2130000_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3394 diff_2150400_597600# diff_1004400_591600# diff_2150400_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3395 diff_2170800_597600# diff_1004400_591600# diff_2170800_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3396 diff_2191200_597600# diff_1004400_591600# diff_2191200_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3397 diff_2211600_597600# diff_1004400_591600# diff_2211600_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3398 diff_2232000_597600# diff_1004400_591600# diff_2232000_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3399 diff_2252400_597600# diff_1004400_591600# diff_2252400_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3400 diff_2272800_597600# diff_1004400_591600# diff_2272800_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3401 diff_2293200_597600# diff_1004400_591600# diff_2293200_574800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3402 diff_1004400_657600# diff_2431200_979200# diff_2367600_607200# GND efet w=79200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3403 diff_2508000_430800# diff_2451600_979200# diff_2367600_696000# GND efet w=154800 l=7200
+ ad=-1.40721e+09 pd=1.1256e+06 as=0 ps=0 
M3404 diff_2367600_607200# diff_2469600_912000# diff_2508000_430800# GND efet w=154800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3405 diff_2367600_519600# diff_2361600_427200# diff_1004400_524400# GND efet w=87600 l=6600
+ ad=-6.51767e+08 pd=729600 as=7.9488e+08 ps=223200 
M3406 diff_1008000_574800# diff_1004400_568800# diff_1008000_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3407 diff_1028400_574800# diff_1004400_568800# diff_1028400_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3408 diff_1048800_574800# diff_1004400_568800# diff_1048800_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3409 diff_1069200_574800# diff_1004400_568800# diff_1069200_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3410 diff_1089600_574800# diff_1004400_568800# diff_1089600_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3411 diff_1110000_574800# diff_1004400_568800# diff_1110000_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3412 diff_1130400_574800# diff_1004400_568800# diff_1130400_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3413 diff_1150800_574800# diff_1004400_568800# diff_1150800_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3414 diff_1171200_574800# diff_1004400_568800# diff_1171200_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3415 diff_1191600_574800# diff_1004400_568800# diff_1191600_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3416 diff_1212000_574800# diff_1004400_568800# diff_1212000_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3417 diff_1232400_574800# diff_1004400_568800# diff_1232400_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3418 diff_1252800_574800# diff_1004400_568800# diff_1252800_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3419 diff_1273200_574800# diff_1004400_568800# diff_1273200_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3420 diff_1293600_574800# diff_1004400_568800# diff_1293600_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3421 diff_1314000_574800# diff_1004400_568800# diff_1314000_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3422 diff_1334400_574800# diff_1004400_568800# diff_1334400_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3423 diff_1354800_574800# diff_1004400_568800# diff_1354800_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3424 diff_1375200_574800# diff_1004400_568800# diff_1375200_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3425 diff_1395600_574800# diff_1004400_568800# diff_1395600_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3426 diff_1416000_574800# diff_1004400_568800# diff_1416000_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3427 diff_1436400_574800# diff_1004400_568800# diff_1436400_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3428 diff_1456800_574800# diff_1004400_568800# diff_1456800_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3429 diff_1477200_574800# diff_1004400_568800# diff_1477200_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3430 diff_1497600_574800# diff_1004400_568800# diff_1497600_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3431 diff_1518000_574800# diff_1004400_568800# diff_1518000_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3432 diff_1538400_574800# diff_1004400_568800# diff_1538400_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3433 diff_1558800_574800# diff_1004400_568800# diff_1558800_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3434 diff_1579200_574800# diff_1004400_568800# diff_1579200_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3435 diff_1599600_574800# diff_1004400_568800# diff_1599600_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3436 diff_1620000_574800# diff_1004400_568800# diff_1620000_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3437 diff_1640400_574800# diff_1004400_568800# diff_1640400_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3438 diff_1660800_574800# diff_1004400_568800# diff_1660800_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3439 diff_1681200_574800# diff_1004400_568800# diff_1681200_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3440 diff_1701600_574800# diff_1004400_568800# diff_1701600_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3441 diff_1722000_574800# diff_1004400_568800# diff_1722000_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3442 diff_1742400_574800# diff_1004400_568800# diff_1742400_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3443 diff_1762800_574800# diff_1004400_568800# diff_1762800_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3444 diff_1783200_574800# diff_1004400_568800# diff_1783200_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3445 diff_1803600_574800# diff_1004400_568800# diff_1803600_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3446 diff_1824000_574800# diff_1004400_568800# diff_1824000_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3447 diff_1844400_574800# diff_1004400_568800# diff_1844400_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3448 diff_1864800_574800# diff_1004400_568800# diff_1864800_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3449 diff_1885200_574800# diff_1004400_568800# diff_1885200_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3450 diff_1905600_574800# diff_1004400_568800# diff_1905600_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3451 diff_1926000_574800# diff_1004400_568800# diff_1926000_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3452 diff_1946400_574800# diff_1004400_568800# diff_1946400_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3453 diff_1966800_574800# diff_1004400_568800# diff_1966800_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3454 diff_1987200_574800# diff_1004400_568800# diff_1987200_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3455 diff_2007600_574800# diff_1004400_568800# diff_2007600_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3456 diff_2028000_574800# diff_1004400_568800# diff_2028000_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3457 diff_2048400_574800# diff_1004400_568800# diff_2048400_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3458 diff_2068800_574800# diff_1004400_568800# diff_2068800_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3459 diff_2089200_574800# diff_1004400_568800# diff_2089200_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3460 diff_2109600_574800# diff_1004400_568800# diff_2109600_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3461 diff_2130000_574800# diff_1004400_568800# diff_2130000_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3462 diff_2150400_574800# diff_1004400_568800# diff_2150400_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3463 diff_2170800_574800# diff_1004400_568800# diff_2170800_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3464 diff_2191200_574800# diff_1004400_568800# diff_2191200_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3465 diff_2211600_574800# diff_1004400_568800# diff_2211600_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3466 diff_2232000_574800# diff_1004400_568800# diff_2232000_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3467 diff_2252400_574800# diff_1004400_568800# diff_2252400_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3468 diff_2272800_574800# diff_1004400_568800# diff_2272800_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3469 diff_2293200_574800# diff_1004400_568800# diff_2293200_553200# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3470 diff_1004400_591600# Vdd Vdd GND efet w=6000 l=13200
+ ad=9.4032e+08 pd=261600 as=0 ps=0 
M3471 diff_776400_488400# Vdd Vdd GND efet w=7800 l=87000
+ ad=3.6288e+08 pd=108000 as=0 ps=0 
M3472 diff_1008000_553200# diff_1004400_547200# diff_1008000_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3473 diff_1028400_553200# diff_1004400_547200# diff_1028400_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3474 diff_1048800_553200# diff_1004400_547200# diff_1048800_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3475 diff_1069200_553200# diff_1004400_547200# diff_1069200_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3476 diff_1089600_553200# diff_1004400_547200# diff_1089600_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3477 diff_1110000_553200# diff_1004400_547200# diff_1110000_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3478 diff_1130400_553200# diff_1004400_547200# diff_1130400_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3479 diff_1150800_553200# diff_1004400_547200# diff_1150800_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3480 diff_1171200_553200# diff_1004400_547200# diff_1171200_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3481 diff_1191600_553200# diff_1004400_547200# diff_1191600_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3482 diff_1212000_553200# diff_1004400_547200# diff_1212000_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3483 diff_1232400_553200# diff_1004400_547200# diff_1232400_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3484 diff_1252800_553200# diff_1004400_547200# diff_1252800_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3485 diff_1273200_553200# diff_1004400_547200# diff_1273200_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3486 diff_1293600_553200# diff_1004400_547200# diff_1293600_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3487 diff_1314000_553200# diff_1004400_547200# diff_1314000_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3488 diff_1334400_553200# diff_1004400_547200# diff_1334400_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3489 diff_1354800_553200# diff_1004400_547200# diff_1354800_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3490 diff_1375200_553200# diff_1004400_547200# diff_1375200_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3491 diff_1395600_553200# diff_1004400_547200# diff_1395600_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3492 diff_1416000_553200# diff_1004400_547200# diff_1416000_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3493 diff_1436400_553200# diff_1004400_547200# diff_1436400_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3494 diff_1456800_553200# diff_1004400_547200# diff_1456800_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3495 diff_1477200_553200# diff_1004400_547200# diff_1477200_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3496 diff_1497600_553200# diff_1004400_547200# diff_1497600_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3497 diff_1518000_553200# diff_1004400_547200# diff_1518000_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3498 diff_1538400_553200# diff_1004400_547200# diff_1538400_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3499 diff_1558800_553200# diff_1004400_547200# diff_1558800_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3500 diff_1579200_553200# diff_1004400_547200# diff_1579200_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3501 diff_1599600_553200# diff_1004400_547200# diff_1599600_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3502 diff_1620000_553200# diff_1004400_547200# diff_1620000_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3503 diff_1640400_553200# diff_1004400_547200# diff_1640400_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3504 diff_1660800_553200# diff_1004400_547200# diff_1660800_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3505 diff_1681200_553200# diff_1004400_547200# diff_1681200_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3506 diff_1701600_553200# diff_1004400_547200# diff_1701600_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3507 diff_1722000_553200# diff_1004400_547200# diff_1722000_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3508 diff_1742400_553200# diff_1004400_547200# diff_1742400_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3509 diff_1762800_553200# diff_1004400_547200# diff_1762800_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3510 diff_1783200_553200# diff_1004400_547200# diff_1783200_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3511 diff_1803600_553200# diff_1004400_547200# diff_1803600_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3512 diff_1824000_553200# diff_1004400_547200# diff_1824000_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3513 diff_1844400_553200# diff_1004400_547200# diff_1844400_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3514 diff_1864800_553200# diff_1004400_547200# diff_1864800_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3515 diff_1885200_553200# diff_1004400_547200# diff_1885200_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3516 diff_1905600_553200# diff_1004400_547200# diff_1905600_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3517 diff_1926000_553200# diff_1004400_547200# diff_1926000_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3518 diff_1946400_553200# diff_1004400_547200# diff_1946400_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3519 diff_1966800_553200# diff_1004400_547200# diff_1966800_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3520 diff_1987200_553200# diff_1004400_547200# diff_1987200_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3521 diff_2007600_553200# diff_1004400_547200# diff_2007600_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3522 diff_2028000_553200# diff_1004400_547200# diff_2028000_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3523 diff_2048400_553200# diff_1004400_547200# diff_2048400_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3524 diff_2068800_553200# diff_1004400_547200# diff_2068800_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3525 diff_2089200_553200# diff_1004400_547200# diff_2089200_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3526 diff_2109600_553200# diff_1004400_547200# diff_2109600_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3527 diff_2130000_553200# diff_1004400_547200# diff_2130000_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3528 diff_2150400_553200# diff_1004400_547200# diff_2150400_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3529 diff_2170800_553200# diff_1004400_547200# diff_2170800_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3530 diff_2191200_553200# diff_1004400_547200# diff_2191200_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3531 diff_2211600_553200# diff_1004400_547200# diff_2211600_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3532 diff_2232000_553200# diff_1004400_547200# diff_2232000_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3533 diff_2252400_553200# diff_1004400_547200# diff_2252400_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3534 diff_2272800_553200# diff_1004400_547200# diff_2272800_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3535 diff_2293200_553200# diff_1004400_547200# diff_2293200_530400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3536 diff_409200_476400# diff_404400_470400# GND GND efet w=32400 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3537 diff_490800_500400# diff_496800_492000# diff_500400_480000# GND efet w=19200 l=7200
+ ad=0 pd=0 as=3.096e+08 ps=88800 
M3538 diff_780000_446400# diff_776400_488400# diff_691200_487200# GND efet w=13200 l=7200
+ ad=8.7552e+08 pd=196800 as=0 ps=0 
M3539 diff_496800_492000# diff_810000_510000# diff_780000_446400# GND efet w=13200 l=7200
+ ad=1.04688e+09 pd=240000 as=0 ps=0 
M3540 diff_500400_480000# cm GND GND efet w=33600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3541 diff_694800_493200# diff_691200_487200# diff_694800_478800# GND efet w=30000 l=7200
+ ad=0 pd=0 as=2.3184e+08 ps=84000 
M3542 diff_691200_487200# diff_691200_487200# diff_691200_487200# GND efet w=1200 l=1200
+ ad=0 pd=0 as=0 ps=0 
M3543 diff_691200_487200# diff_691200_487200# diff_691200_487200# GND efet w=1800 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3544 diff_694800_478800# diff_691200_472800# GND GND efet w=34800 l=6600
+ ad=0 pd=0 as=0 ps=0 
M3545 diff_564000_475200# diff_550800_454800# GND GND efet w=45600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3546 diff_624000_475200# diff_621600_469200# GND GND efet w=45600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3547 diff_338400_375600# diff_321600_398400# GND GND efet w=20400 l=7200
+ ad=8.856e+08 pd=204000 as=0 ps=0 
M3548 diff_382800_375600# diff_367200_398400# GND GND efet w=19200 l=7200
+ ad=7.488e+08 pd=192000 as=0 ps=0 
M3549 diff_429600_375600# diff_414000_398400# GND GND efet w=20400 l=7200
+ ad=6.8544e+08 pd=187200 as=0 ps=0 
M3550 diff_321600_398400# clk1 diff_289200_457200# GND efet w=10800 l=7200
+ ad=1.3824e+08 pd=55200 as=0 ps=0 
M3551 diff_321600_398400# diff_321600_398400# diff_321600_398400# GND efet w=1200 l=5400
+ ad=0 pd=0 as=0 ps=0 
M3552 diff_321600_398400# diff_321600_398400# diff_321600_398400# GND efet w=1800 l=2400
+ ad=0 pd=0 as=0 ps=0 
M3553 diff_367200_398400# clk2 diff_338400_375600# GND efet w=12000 l=7200
+ ad=1.4832e+08 pd=52800 as=0 ps=0 
M3554 diff_367200_398400# diff_367200_398400# diff_367200_398400# GND efet w=1800 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3555 diff_367200_398400# diff_367200_398400# diff_367200_398400# GND efet w=600 l=1200
+ ad=0 pd=0 as=0 ps=0 
M3556 diff_414000_398400# clk1 diff_382800_375600# GND efet w=12000 l=7200
+ ad=1.4256e+08 pd=55200 as=0 ps=0 
M3557 diff_414000_398400# diff_414000_398400# diff_414000_398400# GND efet w=2400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3558 GND diff_756000_454800# diff_691200_487200# GND efet w=13200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3559 diff_474000_375600# diff_459600_398400# GND GND efet w=19200 l=7200
+ ad=7.4016e+08 pd=192000 as=0 ps=0 
M3560 diff_478800_470400# diff_506400_398400# GND GND efet w=20400 l=7200
+ ad=8.5824e+08 pd=211200 as=0 ps=0 
M3561 diff_550800_454800# diff_550800_398400# GND GND efet w=19200 l=7200
+ ad=8.7408e+08 pd=211200 as=0 ps=0 
M3562 diff_613200_375600# diff_597600_398400# GND GND efet w=20400 l=7200
+ ad=6.8544e+08 pd=187200 as=0 ps=0 
M3563 diff_621600_469200# diff_643200_398400# GND GND efet w=19200 l=7200
+ ad=8.5392e+08 pd=211200 as=0 ps=0 
M3564 diff_756000_454800# diff_780000_446400# GND GND efet w=21600 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3565 diff_776400_488400# diff_776400_488400# diff_776400_488400# GND efet w=600 l=1800
+ ad=0 pd=0 as=0 ps=0 
M3566 diff_810000_510000# diff_776400_488400# GND GND efet w=12000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3567 diff_776400_488400# diff_776400_488400# diff_776400_488400# GND efet w=1200 l=1200
+ ad=0 pd=0 as=0 ps=0 
M3568 diff_780000_446400# diff_780000_446400# diff_780000_446400# GND efet w=1800 l=5400
+ ad=0 pd=0 as=0 ps=0 
M3569 diff_780000_446400# diff_780000_446400# diff_780000_446400# GND efet w=1800 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3570 diff_904800_464400# clk2 diff_776400_488400# GND efet w=22800 l=7200
+ ad=2.8944e+08 pd=79200 as=0 ps=0 
M3571 diff_922800_458400# diff_746400_625200# diff_904800_464400# GND efet w=28800 l=7200
+ ad=9.3024e+08 pd=199200 as=0 ps=0 
M3572 Vdd Vdd diff_1004400_524400# GND efet w=6000 l=13200
+ ad=0 pd=0 as=0 ps=0 
M3573 diff_1008000_530400# diff_1004400_524400# diff_1008000_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3574 diff_1028400_530400# diff_1004400_524400# diff_1028400_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3575 diff_1048800_530400# diff_1004400_524400# diff_1048800_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3576 diff_1069200_530400# diff_1004400_524400# diff_1069200_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3577 diff_1089600_530400# diff_1004400_524400# diff_1089600_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3578 diff_1110000_530400# diff_1004400_524400# diff_1110000_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3579 diff_1130400_530400# diff_1004400_524400# diff_1130400_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3580 diff_1150800_530400# diff_1004400_524400# diff_1150800_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3581 diff_1171200_530400# diff_1004400_524400# diff_1171200_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3582 diff_1191600_530400# diff_1004400_524400# diff_1191600_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3583 diff_1212000_530400# diff_1004400_524400# diff_1212000_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3584 diff_1232400_530400# diff_1004400_524400# diff_1232400_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3585 diff_1252800_530400# diff_1004400_524400# diff_1252800_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3586 diff_1273200_530400# diff_1004400_524400# diff_1273200_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3587 diff_1293600_530400# diff_1004400_524400# diff_1293600_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3588 diff_1314000_530400# diff_1004400_524400# diff_1314000_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3589 diff_1334400_530400# diff_1004400_524400# diff_1334400_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3590 diff_1354800_530400# diff_1004400_524400# diff_1354800_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3591 diff_1375200_530400# diff_1004400_524400# diff_1375200_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3592 diff_1395600_530400# diff_1004400_524400# diff_1395600_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3593 diff_1416000_530400# diff_1004400_524400# diff_1416000_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3594 diff_1436400_530400# diff_1004400_524400# diff_1436400_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3595 diff_1456800_530400# diff_1004400_524400# diff_1456800_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3596 diff_1477200_530400# diff_1004400_524400# diff_1477200_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3597 diff_1497600_530400# diff_1004400_524400# diff_1497600_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3598 diff_1518000_530400# diff_1004400_524400# diff_1518000_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3599 diff_1538400_530400# diff_1004400_524400# diff_1538400_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3600 diff_1558800_530400# diff_1004400_524400# diff_1558800_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3601 diff_1579200_530400# diff_1004400_524400# diff_1579200_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3602 diff_1599600_530400# diff_1004400_524400# diff_1599600_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3603 diff_1620000_530400# diff_1004400_524400# diff_1620000_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3604 diff_1640400_530400# diff_1004400_524400# diff_1640400_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3605 diff_1660800_530400# diff_1004400_524400# diff_1660800_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3606 diff_1681200_530400# diff_1004400_524400# diff_1681200_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3607 diff_1701600_530400# diff_1004400_524400# diff_1701600_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3608 diff_1722000_530400# diff_1004400_524400# diff_1722000_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3609 diff_1742400_530400# diff_1004400_524400# diff_1742400_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3610 diff_1762800_530400# diff_1004400_524400# diff_1762800_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3611 diff_1783200_530400# diff_1004400_524400# diff_1783200_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3612 diff_1803600_530400# diff_1004400_524400# diff_1803600_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3613 diff_1824000_530400# diff_1004400_524400# diff_1824000_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3614 diff_1844400_530400# diff_1004400_524400# diff_1844400_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3615 diff_1864800_530400# diff_1004400_524400# diff_1864800_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3616 diff_1885200_530400# diff_1004400_524400# diff_1885200_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3617 diff_1905600_530400# diff_1004400_524400# diff_1905600_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3618 diff_1926000_530400# diff_1004400_524400# diff_1926000_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3619 diff_1946400_530400# diff_1004400_524400# diff_1946400_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3620 diff_1966800_530400# diff_1004400_524400# diff_1966800_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3621 diff_1987200_530400# diff_1004400_524400# diff_1987200_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3622 diff_2007600_530400# diff_1004400_524400# diff_2007600_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3623 diff_2028000_530400# diff_1004400_524400# diff_2028000_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3624 diff_2048400_530400# diff_1004400_524400# diff_2048400_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3625 diff_2068800_530400# diff_1004400_524400# diff_2068800_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3626 diff_2089200_530400# diff_1004400_524400# diff_2089200_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3627 diff_2109600_530400# diff_1004400_524400# diff_2109600_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3628 diff_2130000_530400# diff_1004400_524400# diff_2130000_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3629 diff_2150400_530400# diff_1004400_524400# diff_2150400_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3630 diff_2170800_530400# diff_1004400_524400# diff_2170800_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3631 diff_2191200_530400# diff_1004400_524400# diff_2191200_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3632 diff_2211600_530400# diff_1004400_524400# diff_2211600_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3633 diff_2232000_530400# diff_1004400_524400# diff_2232000_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3634 diff_2252400_530400# diff_1004400_524400# diff_2252400_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3635 diff_2272800_530400# diff_1004400_524400# diff_2272800_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3636 diff_2293200_530400# diff_1004400_524400# diff_2293200_508800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3637 diff_1004400_591600# diff_2384400_427200# diff_2367600_519600# GND efet w=74400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3638 diff_1004400_568800# Vdd Vdd GND efet w=7200 l=13200
+ ad=1.0368e+09 pd=249600 as=0 ps=0 
M3639 Vdd Vdd diff_1004400_547200# GND efet w=7200 l=14400
+ ad=0 pd=0 as=1.02816e+09 ps=220800 
M3640 diff_2367600_519600# diff_2413200_996000# diff_1004400_547200# GND efet w=84600 l=6600
+ ad=0 pd=0 as=0 ps=0 
M3641 diff_1008000_508800# diff_1004400_502800# diff_1008000_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3642 diff_1028400_508800# diff_1004400_502800# diff_1028400_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3643 diff_1048800_508800# diff_1004400_502800# diff_1048800_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3644 diff_1069200_508800# diff_1004400_502800# diff_1069200_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3645 diff_1089600_508800# diff_1004400_502800# diff_1089600_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3646 diff_1110000_508800# diff_1004400_502800# diff_1110000_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3647 diff_1130400_508800# diff_1004400_502800# diff_1130400_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3648 diff_1150800_508800# diff_1004400_502800# diff_1150800_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3649 diff_1171200_508800# diff_1004400_502800# diff_1171200_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3650 diff_1191600_508800# diff_1004400_502800# diff_1191600_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3651 diff_1212000_508800# diff_1004400_502800# diff_1212000_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3652 diff_1232400_508800# diff_1004400_502800# diff_1232400_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3653 diff_1252800_508800# diff_1004400_502800# diff_1252800_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3654 diff_1273200_508800# diff_1004400_502800# diff_1273200_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3655 diff_1293600_508800# diff_1004400_502800# diff_1293600_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3656 diff_1314000_508800# diff_1004400_502800# diff_1314000_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3657 diff_1334400_508800# diff_1004400_502800# diff_1334400_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3658 diff_1354800_508800# diff_1004400_502800# diff_1354800_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3659 diff_1375200_508800# diff_1004400_502800# diff_1375200_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3660 diff_1395600_508800# diff_1004400_502800# diff_1395600_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3661 diff_1416000_508800# diff_1004400_502800# diff_1416000_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3662 diff_1436400_508800# diff_1004400_502800# diff_1436400_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3663 diff_1456800_508800# diff_1004400_502800# diff_1456800_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3664 diff_1477200_508800# diff_1004400_502800# diff_1477200_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3665 diff_1497600_508800# diff_1004400_502800# diff_1497600_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3666 diff_1518000_508800# diff_1004400_502800# diff_1518000_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3667 diff_1538400_508800# diff_1004400_502800# diff_1538400_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3668 diff_1558800_508800# diff_1004400_502800# diff_1558800_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3669 diff_1579200_508800# diff_1004400_502800# diff_1579200_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3670 diff_1599600_508800# diff_1004400_502800# diff_1599600_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3671 diff_1620000_508800# diff_1004400_502800# diff_1620000_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3672 diff_1640400_508800# diff_1004400_502800# diff_1640400_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3673 diff_1660800_508800# diff_1004400_502800# diff_1660800_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3674 diff_1681200_508800# diff_1004400_502800# diff_1681200_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3675 diff_1701600_508800# diff_1004400_502800# diff_1701600_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3676 diff_1722000_508800# diff_1004400_502800# diff_1722000_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3677 diff_1742400_508800# diff_1004400_502800# diff_1742400_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3678 diff_1762800_508800# diff_1004400_502800# diff_1762800_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3679 diff_1783200_508800# diff_1004400_502800# diff_1783200_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3680 diff_1803600_508800# diff_1004400_502800# diff_1803600_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3681 diff_1824000_508800# diff_1004400_502800# diff_1824000_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3682 diff_1844400_508800# diff_1004400_502800# diff_1844400_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3683 diff_1864800_508800# diff_1004400_502800# diff_1864800_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3684 diff_1885200_508800# diff_1004400_502800# diff_1885200_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3685 diff_1905600_508800# diff_1004400_502800# diff_1905600_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3686 diff_1926000_508800# diff_1004400_502800# diff_1926000_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3687 diff_1946400_508800# diff_1004400_502800# diff_1946400_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3688 diff_1966800_508800# diff_1004400_502800# diff_1966800_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3689 diff_1987200_508800# diff_1004400_502800# diff_1987200_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3690 diff_2007600_508800# diff_1004400_502800# diff_2007600_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3691 diff_2028000_508800# diff_1004400_502800# diff_2028000_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3692 diff_2048400_508800# diff_1004400_502800# diff_2048400_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3693 diff_2068800_508800# diff_1004400_502800# diff_2068800_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3694 diff_2089200_508800# diff_1004400_502800# diff_2089200_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3695 diff_2109600_508800# diff_1004400_502800# diff_2109600_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3696 diff_2130000_508800# diff_1004400_502800# diff_2130000_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3697 diff_2150400_508800# diff_1004400_502800# diff_2150400_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3698 diff_2170800_508800# diff_1004400_502800# diff_2170800_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3699 diff_2191200_508800# diff_1004400_502800# diff_2191200_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3700 diff_2211600_508800# diff_1004400_502800# diff_2211600_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3701 diff_2232000_508800# diff_1004400_502800# diff_2232000_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3702 diff_2252400_508800# diff_1004400_502800# diff_2252400_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3703 diff_2272800_508800# diff_1004400_502800# diff_2272800_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3704 diff_2293200_508800# diff_1004400_502800# diff_2293200_486000# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3705 diff_1004400_568800# diff_2431200_979200# diff_2367600_519600# GND efet w=79200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3706 Vdd Vdd Vdd GND efet w=5400 l=7800
+ ad=0 pd=0 as=0 ps=0 
M3707 Vdd Vdd diff_2488800_853200# GND efet w=7200 l=14400
+ ad=0 pd=0 as=-1.86569e+09 ps=422400 
M3708 diff_2774400_1002000# Vdd Vdd GND efet w=7200 l=32400
+ ad=0 pd=0 as=0 ps=0 
M3709 diff_2848800_992400# diff_2779200_486000# diff_2848800_976800# GND efet w=46800 l=6000
+ ad=0 pd=0 as=4.4928e+08 ps=112800 
M3710 Vdd Vdd Vdd GND efet w=2400 l=4800
+ ad=0 pd=0 as=0 ps=0 
M3711 Vdd Vdd Vdd GND efet w=1800 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3712 Vdd Vdd diff_2774400_889200# GND efet w=7200 l=32400
+ ad=0 pd=0 as=9.7776e+08 ps=160800 
M3713 diff_2848800_976800# diff_2732400_549600# GND GND efet w=46800 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3714 diff_2738400_926400# diff_2710800_1356000# diff_2529600_894000# GND efet w=20400 l=6000
+ ad=0 pd=0 as=3.1536e+08 ps=72000 
M3715 diff_2774400_889200# clk2 diff_2738400_926400# GND efet w=20400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3716 diff_2818800_889200# diff_2738400_552000# diff_2774400_889200# GND efet w=37200 l=6000
+ ad=9.6048e+08 pd=199200 as=0 ps=0 
M3717 diff_2738400_813600# diff_2710800_1356000# diff_2598000_656400# GND efet w=20400 l=6000
+ ad=5.8464e+08 pd=139200 as=2.9088e+08 ps=69600 
M3718 diff_2774400_852000# clk2 diff_2738400_813600# GND efet w=20400 l=6000
+ ad=1.15632e+09 pd=211200 as=0 ps=0 
M3719 Vdd Vdd diff_1048800_846000# GND efet w=7200 l=13200
+ ad=0 pd=0 as=1.81152e+09 ps=324000 
M3720 Vdd Vdd diff_994800_1225200# GND efet w=7200 l=13200
+ ad=0 pd=0 as=2.10816e+09 ps=328800 
M3721 Vdd Vdd diff_2505600_919200# GND efet w=8400 l=13200
+ ad=0 pd=0 as=1.99008e+09 ps=326400 
M3722 diff_2738400_813600# diff_2722800_844800# diff_2617200_789600# GND efet w=20400 l=6000
+ ad=0 pd=0 as=2.9088e+08 ps=69600 
M3723 GND diff_2598000_656400# diff_2488800_853200# GND efet w=123600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3724 diff_1048800_846000# diff_2617200_789600# GND GND efet w=123600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3725 GND diff_2665200_789600# diff_994800_1225200# GND efet w=123600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3726 diff_2505600_919200# diff_2686800_789600# GND GND efet w=123600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3727 diff_2738400_776400# diff_2722800_844800# diff_2665200_789600# GND efet w=20400 l=6000
+ ad=6.0336e+08 pd=141600 as=2.9088e+08 ps=69600 
M3728 diff_2774400_852000# Vdd Vdd GND efet w=7200 l=33600
+ ad=0 pd=0 as=0 ps=0 
M3729 Vdd Vdd Vdd GND efet w=3000 l=6600
+ ad=0 pd=0 as=0 ps=0 
M3730 Vdd Vdd Vdd GND efet w=1200 l=4800
+ ad=0 pd=0 as=0 ps=0 
M3731 Vdd Vdd diff_2774400_738000# GND efet w=7200 l=32400
+ ad=0 pd=0 as=1.0152e+09 ps=160800 
M3732 diff_2865600_900000# diff_2732400_549600# diff_2774400_1002000# GND efet w=38400 l=6000
+ ad=3.6864e+08 pd=96000 as=0 ps=0 
M3733 GND diff_2751600_452400# diff_2865600_900000# GND efet w=38400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3734 d0 GND d0 GND efet w=179400 l=112200
+ ad=0 pd=0 as=0 ps=0 
M3735 GND diff_2751600_452400# diff_2818800_889200# GND efet w=36000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3736 diff_2841600_799200# diff_2779200_486000# diff_2774400_852000# GND efet w=36000 l=6000
+ ad=3.456e+08 pd=91200 as=0 ps=0 
M3737 GND diff_2732400_549600# diff_2841600_799200# GND efet w=36000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3738 diff_2738400_776400# diff_2710800_1356000# diff_2686800_789600# GND efet w=21600 l=6000
+ ad=0 pd=0 as=3.312e+08 ps=74400 
M3739 diff_2774400_738000# clk2 diff_2738400_776400# GND efet w=21600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3740 diff_2818800_738000# diff_2738400_552000# diff_2774400_738000# GND efet w=38400 l=6000
+ ad=3.6864e+08 pd=96000 as=0 ps=0 
M3741 GND diff_2779200_486000# diff_2818800_738000# GND efet w=38400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3742 Vdd Vdd Vdd GND efet w=2400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3743 Vdd Vdd Vdd GND efet w=2400 l=4800
+ ad=0 pd=0 as=0 ps=0 
M3744 diff_2732400_549600# Vdd Vdd GND efet w=10800 l=16800
+ ad=1.73808e+09 pd=338400 as=0 ps=0 
M3745 GND diff_2433600_1742400# diff_2508000_430800# GND efet w=301200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3746 diff_2367600_430800# diff_2361600_427200# diff_1004400_435600# GND efet w=89400 l=7200
+ ad=-4.99127e+08 pd=691200 as=8.6112e+08 ps=228000 
M3747 diff_1008000_486000# diff_1004400_480000# diff_1008000_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3748 diff_1028400_486000# diff_1004400_480000# diff_1028400_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3749 diff_1048800_486000# diff_1004400_480000# diff_1048800_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3750 diff_1069200_486000# diff_1004400_480000# diff_1069200_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3751 diff_1089600_486000# diff_1004400_480000# diff_1089600_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3752 diff_1110000_486000# diff_1004400_480000# diff_1110000_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3753 diff_1130400_486000# diff_1004400_480000# diff_1130400_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3754 diff_1150800_486000# diff_1004400_480000# diff_1150800_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3755 diff_1171200_486000# diff_1004400_480000# diff_1171200_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3756 diff_1191600_486000# diff_1004400_480000# diff_1191600_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3757 diff_1212000_486000# diff_1004400_480000# diff_1212000_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3758 diff_1232400_486000# diff_1004400_480000# diff_1232400_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3759 diff_1252800_486000# diff_1004400_480000# diff_1252800_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3760 diff_1273200_486000# diff_1004400_480000# diff_1273200_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3761 diff_1293600_486000# diff_1004400_480000# diff_1293600_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3762 diff_1314000_486000# diff_1004400_480000# diff_1314000_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3763 diff_1334400_486000# diff_1004400_480000# diff_1334400_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3764 diff_1354800_486000# diff_1004400_480000# diff_1354800_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3765 diff_1375200_486000# diff_1004400_480000# diff_1375200_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3766 diff_1395600_486000# diff_1004400_480000# diff_1395600_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3767 diff_1416000_486000# diff_1004400_480000# diff_1416000_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3768 diff_1436400_486000# diff_1004400_480000# diff_1436400_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3769 diff_1456800_486000# diff_1004400_480000# diff_1456800_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3770 diff_1477200_486000# diff_1004400_480000# diff_1477200_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3771 diff_1497600_486000# diff_1004400_480000# diff_1497600_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3772 diff_1518000_486000# diff_1004400_480000# diff_1518000_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3773 diff_1538400_486000# diff_1004400_480000# diff_1538400_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3774 diff_1558800_486000# diff_1004400_480000# diff_1558800_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3775 diff_1579200_486000# diff_1004400_480000# diff_1579200_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3776 diff_1599600_486000# diff_1004400_480000# diff_1599600_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3777 diff_1620000_486000# diff_1004400_480000# diff_1620000_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3778 diff_1640400_486000# diff_1004400_480000# diff_1640400_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3779 diff_1660800_486000# diff_1004400_480000# diff_1660800_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3780 diff_1681200_486000# diff_1004400_480000# diff_1681200_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3781 diff_1701600_486000# diff_1004400_480000# diff_1701600_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3782 diff_1722000_486000# diff_1004400_480000# diff_1722000_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3783 diff_1742400_486000# diff_1004400_480000# diff_1742400_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3784 diff_1762800_486000# diff_1004400_480000# diff_1762800_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3785 diff_1783200_486000# diff_1004400_480000# diff_1783200_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3786 diff_1803600_486000# diff_1004400_480000# diff_1803600_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3787 diff_1824000_486000# diff_1004400_480000# diff_1824000_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3788 diff_1844400_486000# diff_1004400_480000# diff_1844400_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3789 diff_1864800_486000# diff_1004400_480000# diff_1864800_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3790 diff_1885200_486000# diff_1004400_480000# diff_1885200_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3791 diff_1905600_486000# diff_1004400_480000# diff_1905600_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3792 diff_1926000_486000# diff_1004400_480000# diff_1926000_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3793 diff_1946400_486000# diff_1004400_480000# diff_1946400_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3794 diff_1966800_486000# diff_1004400_480000# diff_1966800_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3795 diff_1987200_486000# diff_1004400_480000# diff_1987200_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3796 diff_2007600_486000# diff_1004400_480000# diff_2007600_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3797 diff_2028000_486000# diff_1004400_480000# diff_2028000_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3798 diff_2048400_486000# diff_1004400_480000# diff_2048400_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3799 diff_2068800_486000# diff_1004400_480000# diff_2068800_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3800 diff_2089200_486000# diff_1004400_480000# diff_2089200_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3801 diff_2109600_486000# diff_1004400_480000# diff_2109600_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3802 diff_2130000_486000# diff_1004400_480000# diff_2130000_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3803 diff_2150400_486000# diff_1004400_480000# diff_2150400_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3804 diff_2170800_486000# diff_1004400_480000# diff_2170800_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3805 diff_2191200_486000# diff_1004400_480000# diff_2191200_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3806 diff_2211600_486000# diff_1004400_480000# diff_2211600_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3807 diff_2232000_486000# diff_1004400_480000# diff_2232000_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3808 diff_2252400_486000# diff_1004400_480000# diff_2252400_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3809 diff_2272800_486000# diff_1004400_480000# diff_2272800_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3810 diff_2293200_486000# diff_1004400_480000# diff_2293200_464400# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.5552e+08 ps=50400 
M3811 diff_1004400_502800# Vdd Vdd GND efet w=6000 l=12000
+ ad=9.4032e+08 pd=261600 as=0 ps=0 
M3812 GND cm diff_922800_458400# GND efet w=67200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3813 diff_691200_472800# clk1 GND GND efet w=20400 l=7200
+ ad=8.3088e+08 pd=206400 as=0 ps=0 
M3814 diff_748800_375600# diff_733200_398400# GND GND efet w=19200 l=7200
+ ad=7.488e+08 pd=192000 as=0 ps=0 
M3815 diff_795600_375600# diff_780000_398400# GND GND efet w=20400 l=7200
+ ad=6.8544e+08 pd=187200 as=0 ps=0 
M3816 diff_414000_398400# diff_414000_398400# diff_414000_398400# GND efet w=1200 l=1800
+ ad=0 pd=0 as=0 ps=0 
M3817 diff_459600_398400# clk2 diff_429600_375600# GND efet w=12000 l=7200
+ ad=1.3824e+08 pd=48000 as=0 ps=0 
M3818 diff_459600_398400# diff_459600_398400# diff_459600_398400# GND efet w=1200 l=1800
+ ad=0 pd=0 as=0 ps=0 
M3819 diff_506400_398400# clk1 diff_474000_375600# GND efet w=12000 l=7200
+ ad=1.2816e+08 pd=52800 as=0 ps=0 
M3820 diff_506400_398400# diff_506400_398400# diff_506400_398400# GND efet w=2400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3821 diff_506400_398400# diff_506400_398400# diff_506400_398400# GND efet w=1200 l=1800
+ ad=0 pd=0 as=0 ps=0 
M3822 diff_550800_398400# clk2 diff_478800_470400# GND efet w=12000 l=7200
+ ad=1.4832e+08 pd=52800 as=0 ps=0 
M3823 diff_550800_398400# diff_550800_398400# diff_550800_398400# GND efet w=1800 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3824 diff_550800_398400# diff_550800_398400# diff_550800_398400# GND efet w=600 l=1200
+ ad=0 pd=0 as=0 ps=0 
M3825 diff_597600_398400# clk1 diff_550800_454800# GND efet w=12000 l=7200
+ ad=1.4256e+08 pd=55200 as=0 ps=0 
M3826 diff_597600_398400# diff_597600_398400# diff_597600_398400# GND efet w=2400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3827 diff_597600_398400# diff_597600_398400# diff_597600_398400# GND efet w=1200 l=1800
+ ad=0 pd=0 as=0 ps=0 
M3828 diff_643200_398400# clk2 diff_613200_375600# GND efet w=12000 l=7200
+ ad=1.3824e+08 pd=48000 as=0 ps=0 
M3829 diff_643200_398400# diff_643200_398400# diff_643200_398400# GND efet w=1200 l=1800
+ ad=0 pd=0 as=0 ps=0 
M3830 clk1 clk1 diff_621600_469200# GND efet w=10200 l=9000
+ ad=0 pd=0 as=0 ps=0 
M3831 clk1 clk1 clk1 GND efet w=2400 l=4800
+ ad=0 pd=0 as=0 ps=0 
M3832 clk1 clk1 clk1 GND efet w=1800 l=2400
+ ad=0 pd=0 as=0 ps=0 
M3833 diff_733200_398400# clk2 diff_691200_472800# GND efet w=12000 l=7200
+ ad=1.4832e+08 pd=52800 as=0 ps=0 
M3834 diff_733200_398400# diff_733200_398400# diff_733200_398400# GND efet w=1800 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3835 diff_733200_398400# diff_733200_398400# diff_733200_398400# GND efet w=600 l=1200
+ ad=0 pd=0 as=0 ps=0 
M3836 diff_780000_398400# clk1 diff_748800_375600# GND efet w=12000 l=7200
+ ad=1.4256e+08 pd=55200 as=0 ps=0 
M3837 diff_780000_398400# diff_780000_398400# diff_780000_398400# GND efet w=2400 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3838 diff_840000_375600# diff_825600_398400# GND GND efet w=19200 l=7200
+ ad=8.2944e+08 pd=208800 as=0 ps=0 
M3839 diff_746400_625200# diff_872400_398400# GND GND efet w=20400 l=6000
+ ad=7.5456e+08 pd=199200 as=0 ps=0 
M3840 diff_1008000_464400# diff_1004400_458400# diff_1008000_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3841 diff_1028400_464400# diff_1004400_458400# diff_1028400_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3842 diff_1048800_464400# diff_1004400_458400# diff_1048800_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3843 diff_1069200_464400# diff_1004400_458400# diff_1069200_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3844 diff_1089600_464400# diff_1004400_458400# diff_1089600_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3845 diff_1110000_464400# diff_1004400_458400# diff_1110000_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3846 diff_1130400_464400# diff_1004400_458400# diff_1130400_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3847 diff_1150800_464400# diff_1004400_458400# diff_1150800_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3848 diff_1171200_464400# diff_1004400_458400# diff_1171200_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3849 diff_1191600_464400# diff_1004400_458400# diff_1191600_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3850 diff_1212000_464400# diff_1004400_458400# diff_1212000_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3851 diff_1232400_464400# diff_1004400_458400# diff_1232400_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3852 diff_1252800_464400# diff_1004400_458400# diff_1252800_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3853 diff_1273200_464400# diff_1004400_458400# diff_1273200_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3854 diff_1293600_464400# diff_1004400_458400# diff_1293600_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3855 diff_1314000_464400# diff_1004400_458400# diff_1314000_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3856 diff_1334400_464400# diff_1004400_458400# diff_1334400_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3857 diff_1354800_464400# diff_1004400_458400# diff_1354800_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3858 diff_1375200_464400# diff_1004400_458400# diff_1375200_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3859 diff_1395600_464400# diff_1004400_458400# diff_1395600_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3860 diff_1416000_464400# diff_1004400_458400# diff_1416000_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3861 diff_1436400_464400# diff_1004400_458400# diff_1436400_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3862 diff_1456800_464400# diff_1004400_458400# diff_1456800_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3863 diff_1477200_464400# diff_1004400_458400# diff_1477200_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3864 diff_1497600_464400# diff_1004400_458400# diff_1497600_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3865 diff_1518000_464400# diff_1004400_458400# diff_1518000_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3866 diff_1538400_464400# diff_1004400_458400# diff_1538400_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3867 diff_1558800_464400# diff_1004400_458400# diff_1558800_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3868 diff_1579200_464400# diff_1004400_458400# diff_1579200_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3869 diff_1599600_464400# diff_1004400_458400# diff_1599600_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3870 diff_1620000_464400# diff_1004400_458400# diff_1620000_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3871 diff_1640400_464400# diff_1004400_458400# diff_1640400_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3872 diff_1660800_464400# diff_1004400_458400# diff_1660800_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3873 diff_1681200_464400# diff_1004400_458400# diff_1681200_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3874 diff_1701600_464400# diff_1004400_458400# diff_1701600_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3875 diff_1722000_464400# diff_1004400_458400# diff_1722000_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3876 diff_1742400_464400# diff_1004400_458400# diff_1742400_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3877 diff_1762800_464400# diff_1004400_458400# diff_1762800_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3878 diff_1783200_464400# diff_1004400_458400# diff_1783200_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3879 diff_1803600_464400# diff_1004400_458400# diff_1803600_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3880 diff_1824000_464400# diff_1004400_458400# diff_1824000_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3881 diff_1844400_464400# diff_1004400_458400# diff_1844400_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3882 diff_1864800_464400# diff_1004400_458400# diff_1864800_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3883 diff_1885200_464400# diff_1004400_458400# diff_1885200_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3884 diff_1905600_464400# diff_1004400_458400# diff_1905600_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3885 diff_1926000_464400# diff_1004400_458400# diff_1926000_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3886 diff_1946400_464400# diff_1004400_458400# diff_1946400_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3887 diff_1966800_464400# diff_1004400_458400# diff_1966800_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3888 diff_1987200_464400# diff_1004400_458400# diff_1987200_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3889 diff_2007600_464400# diff_1004400_458400# diff_2007600_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3890 diff_2028000_464400# diff_1004400_458400# diff_2028000_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3891 diff_2048400_464400# diff_1004400_458400# diff_2048400_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3892 diff_2068800_464400# diff_1004400_458400# diff_2068800_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3893 diff_2089200_464400# diff_1004400_458400# diff_2089200_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3894 diff_2109600_464400# diff_1004400_458400# diff_2109600_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3895 diff_2130000_464400# diff_1004400_458400# diff_2130000_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3896 diff_2150400_464400# diff_1004400_458400# diff_2150400_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3897 diff_2170800_464400# diff_1004400_458400# diff_2170800_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3898 diff_2191200_464400# diff_1004400_458400# diff_2191200_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3899 diff_2211600_464400# diff_1004400_458400# diff_2211600_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3900 diff_2232000_464400# diff_1004400_458400# diff_2232000_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3901 diff_2252400_464400# diff_1004400_458400# diff_2252400_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3902 diff_2272800_464400# diff_1004400_458400# diff_2272800_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3903 diff_2293200_464400# diff_1004400_458400# diff_2293200_441600# GND efet w=10800 l=7200
+ ad=0 pd=0 as=1.6848e+08 ps=52800 
M3904 diff_780000_398400# diff_780000_398400# diff_780000_398400# GND efet w=1200 l=1800
+ ad=0 pd=0 as=0 ps=0 
M3905 diff_825600_398400# clk2 diff_795600_375600# GND efet w=12000 l=7200
+ ad=1.3824e+08 pd=48000 as=0 ps=0 
M3906 diff_825600_398400# diff_825600_398400# diff_825600_398400# GND efet w=1200 l=1800
+ ad=0 pd=0 as=0 ps=0 
M3907 diff_872400_398400# clk1 diff_840000_375600# GND efet w=12000 l=7200
+ ad=1.3104e+08 pd=55200 as=0 ps=0 
M3908 diff_872400_398400# diff_872400_398400# diff_872400_398400# GND efet w=2400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3909 diff_872400_398400# diff_872400_398400# diff_872400_398400# GND efet w=1200 l=1800
+ ad=0 pd=0 as=0 ps=0 
M3910 Vdd Vdd diff_289200_457200# GND efet w=7800 l=35400
+ ad=0 pd=0 as=0 ps=0 
M3911 diff_338400_375600# Vdd Vdd GND efet w=7200 l=34800
+ ad=0 pd=0 as=0 ps=0 
M3912 Vdd Vdd diff_382800_375600# GND efet w=7800 l=36600
+ ad=0 pd=0 as=0 ps=0 
M3913 diff_429600_375600# Vdd Vdd GND efet w=7200 l=33600
+ ad=0 pd=0 as=0 ps=0 
M3914 Vdd Vdd diff_474000_375600# GND efet w=7800 l=37800
+ ad=0 pd=0 as=0 ps=0 
M3915 diff_478800_470400# Vdd Vdd GND efet w=7200 l=33600
+ ad=0 pd=0 as=0 ps=0 
M3916 Vdd Vdd diff_550800_454800# GND efet w=7800 l=36600
+ ad=0 pd=0 as=0 ps=0 
M3917 diff_613200_375600# Vdd Vdd GND efet w=7200 l=33600
+ ad=0 pd=0 as=0 ps=0 
M3918 Vdd Vdd diff_621600_469200# GND efet w=7800 l=37800
+ ad=0 pd=0 as=0 ps=0 
M3919 diff_691200_472800# Vdd Vdd GND efet w=7200 l=34800
+ ad=0 pd=0 as=0 ps=0 
M3920 Vdd Vdd diff_748800_375600# GND efet w=7800 l=36600
+ ad=0 pd=0 as=0 ps=0 
M3921 diff_795600_375600# Vdd Vdd GND efet w=7200 l=33600
+ ad=0 pd=0 as=0 ps=0 
M3922 Vdd Vdd diff_840000_375600# GND efet w=7800 l=37800
+ ad=0 pd=0 as=0 ps=0 
M3923 diff_746400_625200# Vdd Vdd GND efet w=7200 l=33600
+ ad=0 pd=0 as=0 ps=0 
M3924 cl GND GND GND efet w=98400 l=7200
+ ad=-1.98167e+08 pd=967200 as=0 ps=0 
M3925 Vdd Vdd diff_1004400_435600# GND efet w=6000 l=12000
+ ad=0 pd=0 as=0 ps=0 
M3926 diff_1008000_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=-2.02332e+09 ps=2.7768e+06 
M3927 diff_1028400_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3928 diff_1048800_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3929 diff_1069200_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3930 diff_1089600_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3931 diff_1110000_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3932 diff_1130400_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3933 diff_1150800_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3934 diff_1171200_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3935 diff_1191600_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3936 diff_1212000_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3937 diff_1232400_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3938 diff_1252800_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3939 diff_1273200_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3940 diff_1293600_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3941 diff_1314000_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3942 diff_1334400_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3943 diff_1354800_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3944 diff_1375200_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3945 diff_1395600_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3946 diff_1416000_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3947 diff_1436400_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3948 diff_1456800_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3949 diff_1477200_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3950 diff_1497600_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3951 diff_1518000_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3952 diff_1538400_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3953 diff_1558800_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3954 diff_1579200_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3955 diff_1599600_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3956 diff_1620000_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3957 diff_1640400_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3958 diff_1660800_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3959 diff_1681200_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3960 diff_1701600_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3961 diff_1722000_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3962 diff_1742400_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3963 diff_1762800_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3964 diff_1783200_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3965 diff_1803600_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3966 diff_1824000_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3967 diff_1844400_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3968 diff_1864800_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3969 diff_1885200_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3970 diff_1905600_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3971 diff_1926000_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3972 diff_1946400_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3973 diff_1966800_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3974 diff_1987200_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3975 diff_2007600_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3976 diff_2028000_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3977 diff_2048400_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3978 diff_2068800_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3979 diff_2089200_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3980 diff_2109600_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3981 diff_2130000_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3982 diff_2150400_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3983 diff_2170800_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3984 diff_2191200_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3985 diff_2211600_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3986 diff_2232000_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3987 diff_2252400_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3988 diff_2272800_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3989 diff_2293200_441600# diff_1004400_435600# diff_1008000_418800# GND efet w=10800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3990 diff_1004400_502800# diff_2384400_427200# diff_2367600_430800# GND efet w=74400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3991 diff_1004400_480000# Vdd Vdd GND efet w=7200 l=12000
+ ad=1.0368e+09 pd=249600 as=0 ps=0 
M3992 Vdd Vdd diff_1004400_458400# GND efet w=7200 l=12000
+ ad=0 pd=0 as=9.8496e+08 ps=220800 
M3993 diff_2367600_430800# diff_2413200_996000# diff_1004400_458400# GND efet w=82800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3994 diff_1004400_480000# diff_2431200_979200# diff_2367600_430800# GND efet w=79200 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3995 diff_2508000_430800# diff_2488800_853200# diff_2367600_519600# GND efet w=154800 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3996 diff_2367600_430800# diff_2505600_919200# diff_2508000_430800# GND efet w=162000 l=7200
+ ad=0 pd=0 as=0 ps=0 
M3997 diff_2732400_549600# d0 GND GND efet w=171600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M3998 diff_2859600_612000# diff_2732400_549600# diff_951600_436800# GND efet w=82800 l=6000
+ ad=8.3088e+08 pd=187200 as=-9.88727e+08 ps=703200 
M3999 diff_2832000_1056000# diff_2751600_452400# diff_2859600_612000# GND efet w=84000 l=6000
+ ad=0 pd=0 as=0 ps=0 
M4000 diff_2738400_552000# diff_2732400_549600# GND GND efet w=44400 l=6000
+ ad=7.2432e+08 pd=153600 as=0 ps=0 
M4001 diff_2738400_552000# Vdd Vdd GND efet w=7200 l=16800
+ ad=0 pd=0 as=0 ps=0 
M4002 diff_2779200_486000# Vdd Vdd GND efet w=9600 l=16800
+ ad=5.8032e+08 pd=124800 as=0 ps=0 
M4003 Vdd Vdd diff_2751600_452400# GND efet w=7200 l=18000
+ ad=0 pd=0 as=-2.13785e+09 ps=518400 
M4004 GND diff_2751600_452400# diff_2779200_486000# GND efet w=44400 l=6000
+ ad=0 pd=0 as=0 ps=0 
M4005 diff_2751600_452400# d1 GND GND efet w=171600 l=6000
+ ad=0 pd=0 as=0 ps=0 
M4006 GND diff_951600_436800# diff_496800_492000# GND efet w=19200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M4007 diff_1008000_418800# diff_1003200_1702800# GND GND efet w=619200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M4008 diff_1008000_418800# diff_1657200_1702800# Vdd GND efet w=643200 l=7200
+ ad=0 pd=0 as=0 ps=0 
M4009 Vdd Vdd Vdd GND efet w=3000 l=4800
+ ad=0 pd=0 as=0 ps=0 
M4010 Vdd Vdd Vdd GND efet w=2400 l=6600
+ ad=0 pd=0 as=0 ps=0 
M4011 Vdd Vdd diff_496800_492000# GND efet w=8400 l=33600
+ ad=0 pd=0 as=0 ps=0 
M4012 Vdd Vdd Vdd GND efet w=600 l=1800
+ ad=0 pd=0 as=0 ps=0 
M4013 Vdd Vdd Vdd GND efet w=2400 l=3000
+ ad=0 pd=0 as=0 ps=0 
M4014 diff_919200_421200# Vdd Vdd GND efet w=7800 l=41400
+ ad=0 pd=0 as=0 ps=0 
M4015 Vdd Vdd diff_951600_436800# GND efet w=9000 l=34200
+ ad=0 pd=0 as=0 ps=0 
M4016 cm GND GND GND efet w=99600 l=7200
+ ad=-7.79927e+08 pd=770400 as=0 ps=0 
C0 metal_1828800_184800# gnd! 5.9fF ;**FLOATING
C1 metal_1810800_188400# gnd! 7.5fF ;**FLOATING
C2 metal_1708800_156000# gnd! 7.1fF ;**FLOATING
C3 metal_1702800_156000# gnd! 3.0fF ;**FLOATING
C4 metal_1729200_178800# gnd! 21.1fF ;**FLOATING
C5 metal_1657200_166800# gnd! 8.3fF ;**FLOATING
C6 metal_1794000_157200# gnd! 10.6fF ;**FLOATING
C7 metal_1783200_184800# gnd! 5.9fF ;**FLOATING
C8 metal_1648800_163200# gnd! 18.4fF ;**FLOATING
C9 metal_411600_163200# gnd! 18.8fF ;**FLOATING
C10 metal_361200_170400# gnd! 39.8fF ;**FLOATING
C11 metal_312000_172800# gnd! 41.6fF ;**FLOATING
C12 metal_265200_181200# gnd! 37.8fF ;**FLOATING
C13 diff_2622000_69600# gnd! 1328.1fF ;**FLOATING
C14 diff_2859600_612000# gnd! 101.8fF
C15 diff_1008000_418800# gnd! 1748.0fF
C16 diff_951600_436800# gnd! 734.5fF
C17 diff_2293200_441600# gnd! 26.2fF
C18 diff_2272800_441600# gnd! 26.2fF
C19 diff_2252400_441600# gnd! 26.2fF
C20 diff_2232000_441600# gnd! 26.2fF
C21 diff_2211600_441600# gnd! 26.2fF
C22 diff_2191200_441600# gnd! 26.2fF
C23 diff_2170800_441600# gnd! 26.2fF
C24 diff_2150400_441600# gnd! 26.2fF
C25 diff_2130000_441600# gnd! 26.2fF
C26 diff_2109600_441600# gnd! 26.2fF
C27 diff_2089200_441600# gnd! 26.2fF
C28 diff_2068800_441600# gnd! 26.2fF
C29 diff_2048400_441600# gnd! 26.2fF
C30 diff_2028000_441600# gnd! 26.2fF
C31 diff_2007600_441600# gnd! 26.2fF
C32 diff_1987200_441600# gnd! 26.2fF
C33 diff_1966800_441600# gnd! 26.2fF
C34 diff_1946400_441600# gnd! 26.2fF
C35 diff_1926000_441600# gnd! 26.2fF
C36 diff_1905600_441600# gnd! 26.2fF
C37 diff_1885200_441600# gnd! 26.2fF
C38 diff_1864800_441600# gnd! 26.2fF
C39 diff_1844400_441600# gnd! 26.2fF
C40 diff_1824000_441600# gnd! 26.2fF
C41 diff_1803600_441600# gnd! 26.2fF
C42 diff_1783200_441600# gnd! 26.2fF
C43 diff_1762800_441600# gnd! 26.2fF
C44 diff_1742400_441600# gnd! 26.2fF
C45 diff_1722000_441600# gnd! 26.2fF
C46 diff_1701600_441600# gnd! 26.2fF
C47 diff_1681200_441600# gnd! 26.2fF
C48 diff_1660800_441600# gnd! 26.2fF
C49 diff_1640400_441600# gnd! 26.2fF
C50 diff_1620000_441600# gnd! 26.2fF
C51 diff_1599600_441600# gnd! 26.2fF
C52 diff_1579200_441600# gnd! 26.2fF
C53 diff_1558800_441600# gnd! 26.2fF
C54 diff_1538400_441600# gnd! 26.2fF
C55 diff_1518000_441600# gnd! 26.2fF
C56 diff_1497600_441600# gnd! 26.2fF
C57 diff_1477200_441600# gnd! 26.2fF
C58 diff_1456800_441600# gnd! 26.2fF
C59 diff_1436400_441600# gnd! 26.2fF
C60 diff_1416000_441600# gnd! 26.2fF
C61 diff_1395600_441600# gnd! 26.2fF
C62 diff_1375200_441600# gnd! 26.2fF
C63 diff_1354800_441600# gnd! 26.2fF
C64 diff_1334400_441600# gnd! 26.2fF
C65 diff_1314000_441600# gnd! 26.2fF
C66 diff_1293600_441600# gnd! 26.2fF
C67 diff_1273200_441600# gnd! 26.2fF
C68 diff_1252800_441600# gnd! 26.2fF
C69 diff_1232400_441600# gnd! 26.2fF
C70 diff_1212000_441600# gnd! 26.2fF
C71 diff_1191600_441600# gnd! 26.2fF
C72 diff_1171200_441600# gnd! 26.2fF
C73 diff_1150800_441600# gnd! 26.2fF
C74 diff_1130400_441600# gnd! 26.2fF
C75 diff_1110000_441600# gnd! 26.2fF
C76 diff_1089600_441600# gnd! 26.2fF
C77 diff_1069200_441600# gnd! 26.2fF
C78 diff_1048800_441600# gnd! 26.2fF
C79 diff_1028400_441600# gnd! 26.2fF
C80 diff_1008000_441600# gnd! 26.2fF
C81 diff_1004400_458400# gnd! 631.7fF
C82 diff_2293200_464400# gnd! 24.7fF
C83 diff_2272800_464400# gnd! 24.7fF
C84 diff_2252400_464400# gnd! 24.7fF
C85 diff_2232000_464400# gnd! 24.7fF
C86 diff_2211600_464400# gnd! 24.7fF
C87 diff_2191200_464400# gnd! 24.7fF
C88 diff_2170800_464400# gnd! 24.7fF
C89 diff_2150400_464400# gnd! 24.7fF
C90 diff_2130000_464400# gnd! 24.7fF
C91 diff_2109600_464400# gnd! 24.7fF
C92 diff_2089200_464400# gnd! 24.7fF
C93 diff_2068800_464400# gnd! 24.7fF
C94 diff_2048400_464400# gnd! 24.7fF
C95 diff_2028000_464400# gnd! 24.7fF
C96 diff_2007600_464400# gnd! 24.7fF
C97 diff_1987200_464400# gnd! 24.7fF
C98 diff_1966800_464400# gnd! 24.7fF
C99 diff_1946400_464400# gnd! 24.7fF
C100 diff_1926000_464400# gnd! 24.7fF
C101 diff_1905600_464400# gnd! 24.7fF
C102 diff_1885200_464400# gnd! 24.7fF
C103 diff_1864800_464400# gnd! 24.7fF
C104 diff_1844400_464400# gnd! 24.7fF
C105 diff_1824000_464400# gnd! 24.7fF
C106 diff_1803600_464400# gnd! 24.7fF
C107 diff_1783200_464400# gnd! 24.7fF
C108 diff_1762800_464400# gnd! 24.7fF
C109 diff_1742400_464400# gnd! 24.7fF
C110 diff_1722000_464400# gnd! 24.7fF
C111 diff_1701600_464400# gnd! 24.7fF
C112 diff_1681200_464400# gnd! 24.7fF
C113 diff_1660800_464400# gnd! 24.7fF
C114 diff_1640400_464400# gnd! 24.7fF
C115 diff_1620000_464400# gnd! 24.7fF
C116 diff_1599600_464400# gnd! 24.7fF
C117 diff_1579200_464400# gnd! 24.7fF
C118 diff_1558800_464400# gnd! 24.7fF
C119 diff_1538400_464400# gnd! 24.7fF
C120 diff_1518000_464400# gnd! 24.7fF
C121 diff_1497600_464400# gnd! 24.7fF
C122 diff_1477200_464400# gnd! 24.7fF
C123 diff_1456800_464400# gnd! 24.7fF
C124 diff_1436400_464400# gnd! 24.7fF
C125 diff_1416000_464400# gnd! 24.7fF
C126 diff_1395600_464400# gnd! 24.7fF
C127 diff_1375200_464400# gnd! 24.7fF
C128 diff_1354800_464400# gnd! 24.7fF
C129 diff_1334400_464400# gnd! 24.7fF
C130 diff_1314000_464400# gnd! 24.7fF
C131 diff_1293600_464400# gnd! 24.7fF
C132 diff_1273200_464400# gnd! 24.7fF
C133 diff_1252800_464400# gnd! 24.7fF
C134 diff_1232400_464400# gnd! 24.7fF
C135 diff_1212000_464400# gnd! 24.7fF
C136 diff_1191600_464400# gnd! 24.7fF
C137 diff_1171200_464400# gnd! 24.7fF
C138 diff_1150800_464400# gnd! 24.7fF
C139 diff_1130400_464400# gnd! 24.7fF
C140 diff_1110000_464400# gnd! 24.7fF
C141 diff_1089600_464400# gnd! 24.7fF
C142 diff_1069200_464400# gnd! 24.7fF
C143 diff_1048800_464400# gnd! 24.7fF
C144 diff_1028400_464400# gnd! 24.7fF
C145 diff_795600_375600# gnd! 87.3fF
C146 diff_748800_375600# gnd! 94.1fF
C147 diff_872400_398400# gnd! 37.8fF
C148 diff_825600_398400# gnd! 41.1fF
C149 diff_780000_398400# gnd! 42.1fF
C150 diff_733200_398400# gnd! 42.2fF
C151 diff_1008000_464400# gnd! 24.7fF
C152 diff_1004400_480000# gnd! 653.0fF
C153 diff_2293200_486000# gnd! 26.2fF
C154 diff_2272800_486000# gnd! 26.2fF
C155 diff_2252400_486000# gnd! 26.2fF
C156 diff_2232000_486000# gnd! 26.2fF
C157 diff_2211600_486000# gnd! 26.2fF
C158 diff_2191200_486000# gnd! 26.2fF
C159 diff_2170800_486000# gnd! 26.2fF
C160 diff_2150400_486000# gnd! 26.2fF
C161 diff_2130000_486000# gnd! 26.2fF
C162 diff_2109600_486000# gnd! 26.2fF
C163 diff_2089200_486000# gnd! 26.2fF
C164 diff_2068800_486000# gnd! 26.2fF
C165 diff_2048400_486000# gnd! 26.2fF
C166 diff_2028000_486000# gnd! 26.2fF
C167 diff_2007600_486000# gnd! 26.2fF
C168 diff_1987200_486000# gnd! 26.2fF
C169 diff_1966800_486000# gnd! 26.2fF
C170 diff_1946400_486000# gnd! 26.2fF
C171 diff_1926000_486000# gnd! 26.2fF
C172 diff_1905600_486000# gnd! 26.2fF
C173 diff_1885200_486000# gnd! 26.2fF
C174 diff_1864800_486000# gnd! 26.2fF
C175 diff_1844400_486000# gnd! 26.2fF
C176 diff_1824000_486000# gnd! 26.2fF
C177 diff_1803600_486000# gnd! 26.2fF
C178 diff_1783200_486000# gnd! 26.2fF
C179 diff_1762800_486000# gnd! 26.2fF
C180 diff_1742400_486000# gnd! 26.2fF
C181 diff_1722000_486000# gnd! 26.2fF
C182 diff_1701600_486000# gnd! 26.2fF
C183 diff_1681200_486000# gnd! 26.2fF
C184 diff_1660800_486000# gnd! 26.2fF
C185 diff_1640400_486000# gnd! 26.2fF
C186 diff_1620000_486000# gnd! 26.2fF
C187 diff_1599600_486000# gnd! 26.2fF
C188 diff_1579200_486000# gnd! 26.2fF
C189 diff_1558800_486000# gnd! 26.2fF
C190 diff_1538400_486000# gnd! 26.2fF
C191 diff_1518000_486000# gnd! 26.2fF
C192 diff_1497600_486000# gnd! 26.2fF
C193 diff_1477200_486000# gnd! 26.2fF
C194 diff_1456800_486000# gnd! 26.2fF
C195 diff_1436400_486000# gnd! 26.2fF
C196 diff_1416000_486000# gnd! 26.2fF
C197 diff_1395600_486000# gnd! 26.2fF
C198 diff_1375200_486000# gnd! 26.2fF
C199 diff_1354800_486000# gnd! 26.2fF
C200 diff_1334400_486000# gnd! 26.2fF
C201 diff_1314000_486000# gnd! 26.2fF
C202 diff_1293600_486000# gnd! 26.2fF
C203 diff_1273200_486000# gnd! 26.2fF
C204 diff_1252800_486000# gnd! 26.2fF
C205 diff_1232400_486000# gnd! 26.2fF
C206 diff_1212000_486000# gnd! 26.2fF
C207 diff_1191600_486000# gnd! 26.2fF
C208 diff_1171200_486000# gnd! 26.2fF
C209 diff_1150800_486000# gnd! 26.2fF
C210 diff_1130400_486000# gnd! 26.2fF
C211 diff_1110000_486000# gnd! 26.2fF
C212 diff_1089600_486000# gnd! 26.2fF
C213 diff_1069200_486000# gnd! 26.2fF
C214 diff_1048800_486000# gnd! 26.2fF
C215 diff_1028400_486000# gnd! 26.2fF
C216 diff_1008000_486000# gnd! 26.2fF
C217 diff_2367600_430800# gnd! 519.2fF
C218 diff_1004400_435600# gnd! 598.0fF
C219 diff_2818800_738000# gnd! 46.5fF
C220 diff_2774400_738000# gnd! 117.6fF
C221 diff_2841600_799200# gnd! 43.7fF
C222 diff_2865600_900000# gnd! 46.5fF
C223 diff_2738400_776400# gnd! 92.4fF
C224 diff_2686800_789600# gnd! 113.8fF
C225 diff_2665200_789600# gnd! 110.7fF
C226 diff_2617200_789600# gnd! 122.4fF
C227 diff_2774400_852000# gnd! 164.5fF
C228 diff_2738400_813600# gnd! 90.0fF
C229 diff_2598000_656400# gnd! 138.3fF
C230 diff_2818800_889200# gnd! 145.9fF
C231 diff_2774400_889200# gnd! 113.9fF
C232 diff_2738400_552000# gnd! 217.4fF
C233 diff_2751600_452400# gnd! 542.6fF
C234 diff_2732400_549600# gnd! 457.7fF
C235 diff_2848800_976800# gnd! 56.2fF
C236 diff_2779200_486000# gnd! 326.9fF
C237 diff_2848800_992400# gnd! 56.2fF
C238 diff_1004400_502800# gnd! 622.9fF
C239 diff_2293200_508800# gnd! 24.7fF
C240 diff_2272800_508800# gnd! 24.7fF
C241 diff_2252400_508800# gnd! 24.7fF
C242 diff_2232000_508800# gnd! 24.7fF
C243 diff_2211600_508800# gnd! 24.7fF
C244 diff_2191200_508800# gnd! 24.7fF
C245 diff_2170800_508800# gnd! 24.7fF
C246 diff_2150400_508800# gnd! 24.7fF
C247 diff_2130000_508800# gnd! 24.7fF
C248 diff_2109600_508800# gnd! 24.7fF
C249 diff_2089200_508800# gnd! 24.7fF
C250 diff_2068800_508800# gnd! 24.7fF
C251 diff_2048400_508800# gnd! 24.7fF
C252 diff_2028000_508800# gnd! 24.7fF
C253 diff_2007600_508800# gnd! 24.7fF
C254 diff_1987200_508800# gnd! 24.7fF
C255 diff_1966800_508800# gnd! 24.7fF
C256 diff_1946400_508800# gnd! 24.7fF
C257 diff_1926000_508800# gnd! 24.7fF
C258 diff_1905600_508800# gnd! 24.7fF
C259 diff_1885200_508800# gnd! 24.7fF
C260 diff_1864800_508800# gnd! 24.7fF
C261 diff_1844400_508800# gnd! 24.7fF
C262 diff_1824000_508800# gnd! 24.7fF
C263 diff_1803600_508800# gnd! 24.7fF
C264 diff_1783200_508800# gnd! 24.7fF
C265 diff_1762800_508800# gnd! 24.7fF
C266 diff_1742400_508800# gnd! 24.7fF
C267 diff_1722000_508800# gnd! 24.7fF
C268 diff_1701600_508800# gnd! 24.7fF
C269 diff_1681200_508800# gnd! 24.7fF
C270 diff_1660800_508800# gnd! 24.7fF
C271 diff_1640400_508800# gnd! 24.7fF
C272 diff_1620000_508800# gnd! 24.7fF
C273 diff_1599600_508800# gnd! 24.7fF
C274 diff_1579200_508800# gnd! 24.7fF
C275 diff_1558800_508800# gnd! 24.7fF
C276 diff_1538400_508800# gnd! 24.7fF
C277 diff_1518000_508800# gnd! 24.7fF
C278 diff_1497600_508800# gnd! 24.7fF
C279 diff_1477200_508800# gnd! 24.7fF
C280 diff_1456800_508800# gnd! 24.7fF
C281 diff_1436400_508800# gnd! 24.7fF
C282 diff_1416000_508800# gnd! 24.7fF
C283 diff_1395600_508800# gnd! 24.7fF
C284 diff_1375200_508800# gnd! 24.7fF
C285 diff_1354800_508800# gnd! 24.7fF
C286 diff_1334400_508800# gnd! 24.7fF
C287 diff_1314000_508800# gnd! 24.7fF
C288 diff_1293600_508800# gnd! 24.7fF
C289 diff_1273200_508800# gnd! 24.7fF
C290 diff_1252800_508800# gnd! 24.7fF
C291 diff_1232400_508800# gnd! 24.7fF
C292 diff_1212000_508800# gnd! 24.7fF
C293 diff_1191600_508800# gnd! 24.7fF
C294 diff_1171200_508800# gnd! 24.7fF
C295 diff_1150800_508800# gnd! 24.7fF
C296 diff_1130400_508800# gnd! 24.7fF
C297 diff_1110000_508800# gnd! 24.7fF
C298 diff_1089600_508800# gnd! 24.7fF
C299 diff_1069200_508800# gnd! 24.7fF
C300 diff_1048800_508800# gnd! 24.7fF
C301 diff_1028400_508800# gnd! 24.7fF
C302 diff_1008000_508800# gnd! 24.7fF
C303 diff_2293200_530400# gnd! 26.2fF
C304 diff_2272800_530400# gnd! 26.2fF
C305 diff_2252400_530400# gnd! 26.2fF
C306 diff_2232000_530400# gnd! 26.2fF
C307 diff_2211600_530400# gnd! 26.2fF
C308 diff_2191200_530400# gnd! 26.2fF
C309 diff_2170800_530400# gnd! 26.2fF
C310 diff_2150400_530400# gnd! 26.2fF
C311 diff_2130000_530400# gnd! 26.2fF
C312 diff_2109600_530400# gnd! 26.2fF
C313 diff_2089200_530400# gnd! 26.2fF
C314 diff_2068800_530400# gnd! 26.2fF
C315 diff_2048400_530400# gnd! 26.2fF
C316 diff_2028000_530400# gnd! 26.2fF
C317 diff_2007600_530400# gnd! 26.2fF
C318 diff_1987200_530400# gnd! 26.2fF
C319 diff_1966800_530400# gnd! 26.2fF
C320 diff_1946400_530400# gnd! 26.2fF
C321 diff_1926000_530400# gnd! 26.2fF
C322 diff_1905600_530400# gnd! 26.2fF
C323 diff_1885200_530400# gnd! 26.2fF
C324 diff_1864800_530400# gnd! 26.2fF
C325 diff_1844400_530400# gnd! 26.2fF
C326 diff_1824000_530400# gnd! 26.2fF
C327 diff_1803600_530400# gnd! 26.2fF
C328 diff_1783200_530400# gnd! 26.2fF
C329 diff_1762800_530400# gnd! 26.2fF
C330 diff_1742400_530400# gnd! 26.2fF
C331 diff_1722000_530400# gnd! 26.2fF
C332 diff_1701600_530400# gnd! 26.2fF
C333 diff_1681200_530400# gnd! 26.2fF
C334 diff_1660800_530400# gnd! 26.2fF
C335 diff_1640400_530400# gnd! 26.2fF
C336 diff_1620000_530400# gnd! 26.2fF
C337 diff_1599600_530400# gnd! 26.2fF
C338 diff_1579200_530400# gnd! 26.2fF
C339 diff_1558800_530400# gnd! 26.2fF
C340 diff_1538400_530400# gnd! 26.2fF
C341 diff_1518000_530400# gnd! 26.2fF
C342 diff_1497600_530400# gnd! 26.2fF
C343 diff_1477200_530400# gnd! 26.2fF
C344 diff_1456800_530400# gnd! 26.2fF
C345 diff_1436400_530400# gnd! 26.2fF
C346 diff_1416000_530400# gnd! 26.2fF
C347 diff_1395600_530400# gnd! 26.2fF
C348 diff_1375200_530400# gnd! 26.2fF
C349 diff_1354800_530400# gnd! 26.2fF
C350 diff_1334400_530400# gnd! 26.2fF
C351 diff_1314000_530400# gnd! 26.2fF
C352 diff_1293600_530400# gnd! 26.2fF
C353 diff_1273200_530400# gnd! 26.2fF
C354 diff_1252800_530400# gnd! 26.2fF
C355 diff_1232400_530400# gnd! 26.2fF
C356 diff_1212000_530400# gnd! 26.2fF
C357 diff_1191600_530400# gnd! 26.2fF
C358 diff_1171200_530400# gnd! 26.2fF
C359 diff_1150800_530400# gnd! 26.2fF
C360 diff_1130400_530400# gnd! 26.2fF
C361 diff_1110000_530400# gnd! 26.2fF
C362 diff_1089600_530400# gnd! 26.2fF
C363 diff_1069200_530400# gnd! 26.2fF
C364 diff_1048800_530400# gnd! 26.2fF
C365 diff_1028400_530400# gnd! 26.2fF
C366 diff_922800_458400# gnd! 112.9fF
C367 diff_904800_464400# gnd! 36.9fF
C368 diff_613200_375600# gnd! 87.3fF
C369 diff_474000_375600# gnd! 93.2fF
C370 diff_643200_398400# gnd! 41.5fF
C371 diff_597600_398400# gnd! 41.7fF
C372 diff_550800_398400# gnd! 42.6fF
C373 diff_506400_398400# gnd! 40.0fF
C374 diff_459600_398400# gnd! 41.5fF
C375 diff_429600_375600# gnd! 87.3fF
C376 diff_382800_375600# gnd! 94.1fF
C377 diff_414000_398400# gnd! 41.7fF
C378 diff_367200_398400# gnd! 42.6fF
C379 diff_321600_398400# gnd! 40.9fF
C380 diff_621600_469200# gnd! 145.3fF
C381 diff_550800_454800# gnd! 153.6fF
C382 diff_691200_472800# gnd! 138.8fF
C383 diff_694800_478800# gnd! 31.6fF
C384 diff_500400_480000# gnd! 39.8fF
C385 diff_780000_446400# gnd! 140.2fF
C386 diff_289200_457200# gnd! 141.0fF
C387 diff_810000_510000# gnd! 108.7fF
C388 diff_1008000_530400# gnd! 26.2fF
C389 diff_1004400_547200# gnd! 636.7fF
C390 diff_2293200_553200# gnd! 24.7fF
C391 diff_2272800_553200# gnd! 24.7fF
C392 diff_2252400_553200# gnd! 24.7fF
C393 diff_2232000_553200# gnd! 24.7fF
C394 diff_2211600_553200# gnd! 24.7fF
C395 diff_2191200_553200# gnd! 24.7fF
C396 diff_2170800_553200# gnd! 24.7fF
C397 diff_2150400_553200# gnd! 24.7fF
C398 diff_2130000_553200# gnd! 24.7fF
C399 diff_2109600_553200# gnd! 24.7fF
C400 diff_2089200_553200# gnd! 24.7fF
C401 diff_2068800_553200# gnd! 24.7fF
C402 diff_2048400_553200# gnd! 24.7fF
C403 diff_2028000_553200# gnd! 24.7fF
C404 diff_2007600_553200# gnd! 24.7fF
C405 diff_1987200_553200# gnd! 24.7fF
C406 diff_1966800_553200# gnd! 24.7fF
C407 diff_1946400_553200# gnd! 24.7fF
C408 diff_1926000_553200# gnd! 24.7fF
C409 diff_1905600_553200# gnd! 24.7fF
C410 diff_1885200_553200# gnd! 24.7fF
C411 diff_1864800_553200# gnd! 24.7fF
C412 diff_1844400_553200# gnd! 24.7fF
C413 diff_1824000_553200# gnd! 24.7fF
C414 diff_1803600_553200# gnd! 24.7fF
C415 diff_1783200_553200# gnd! 24.7fF
C416 diff_1762800_553200# gnd! 24.7fF
C417 diff_1742400_553200# gnd! 24.7fF
C418 diff_1722000_553200# gnd! 24.7fF
C419 diff_1701600_553200# gnd! 24.7fF
C420 diff_1681200_553200# gnd! 24.7fF
C421 diff_1660800_553200# gnd! 24.7fF
C422 diff_1640400_553200# gnd! 24.7fF
C423 diff_1620000_553200# gnd! 24.7fF
C424 diff_1599600_553200# gnd! 24.7fF
C425 diff_1579200_553200# gnd! 24.7fF
C426 diff_1558800_553200# gnd! 24.7fF
C427 diff_1538400_553200# gnd! 24.7fF
C428 diff_1518000_553200# gnd! 24.7fF
C429 diff_1497600_553200# gnd! 24.7fF
C430 diff_1477200_553200# gnd! 24.7fF
C431 diff_1456800_553200# gnd! 24.7fF
C432 diff_1436400_553200# gnd! 24.7fF
C433 diff_1416000_553200# gnd! 24.7fF
C434 diff_1395600_553200# gnd! 24.7fF
C435 diff_1375200_553200# gnd! 24.7fF
C436 diff_1354800_553200# gnd! 24.7fF
C437 diff_1334400_553200# gnd! 24.7fF
C438 diff_1314000_553200# gnd! 24.7fF
C439 diff_1293600_553200# gnd! 24.7fF
C440 diff_1273200_553200# gnd! 24.7fF
C441 diff_1252800_553200# gnd! 24.7fF
C442 diff_1232400_553200# gnd! 24.7fF
C443 diff_1212000_553200# gnd! 24.7fF
C444 diff_1191600_553200# gnd! 24.7fF
C445 diff_1171200_553200# gnd! 24.7fF
C446 diff_1150800_553200# gnd! 24.7fF
C447 diff_1130400_553200# gnd! 24.7fF
C448 diff_1110000_553200# gnd! 24.7fF
C449 diff_1089600_553200# gnd! 24.7fF
C450 diff_1069200_553200# gnd! 24.7fF
C451 diff_1048800_553200# gnd! 24.7fF
C452 diff_1028400_553200# gnd! 24.7fF
C453 diff_1008000_553200# gnd! 24.7fF
C454 diff_1004400_568800# gnd! 652.0fF
C455 diff_2293200_574800# gnd! 26.2fF
C456 diff_2272800_574800# gnd! 26.2fF
C457 diff_2252400_574800# gnd! 26.2fF
C458 diff_2232000_574800# gnd! 26.2fF
C459 diff_2211600_574800# gnd! 26.2fF
C460 diff_2191200_574800# gnd! 26.2fF
C461 diff_2170800_574800# gnd! 26.2fF
C462 diff_2150400_574800# gnd! 26.2fF
C463 diff_2130000_574800# gnd! 26.2fF
C464 diff_2109600_574800# gnd! 26.2fF
C465 diff_2089200_574800# gnd! 26.2fF
C466 diff_2068800_574800# gnd! 26.2fF
C467 diff_2048400_574800# gnd! 26.2fF
C468 diff_2028000_574800# gnd! 26.2fF
C469 diff_2007600_574800# gnd! 26.2fF
C470 diff_1987200_574800# gnd! 26.2fF
C471 diff_1966800_574800# gnd! 26.2fF
C472 diff_1946400_574800# gnd! 26.2fF
C473 diff_1926000_574800# gnd! 26.2fF
C474 diff_1905600_574800# gnd! 26.2fF
C475 diff_1885200_574800# gnd! 26.2fF
C476 diff_1864800_574800# gnd! 26.2fF
C477 diff_1844400_574800# gnd! 26.2fF
C478 diff_1824000_574800# gnd! 26.2fF
C479 diff_1803600_574800# gnd! 26.2fF
C480 diff_1783200_574800# gnd! 26.2fF
C481 diff_1762800_574800# gnd! 26.2fF
C482 diff_1742400_574800# gnd! 26.2fF
C483 diff_1722000_574800# gnd! 26.2fF
C484 diff_1701600_574800# gnd! 26.2fF
C485 diff_1681200_574800# gnd! 26.2fF
C486 diff_1660800_574800# gnd! 26.2fF
C487 diff_1640400_574800# gnd! 26.2fF
C488 diff_1620000_574800# gnd! 26.2fF
C489 diff_1599600_574800# gnd! 26.2fF
C490 diff_1579200_574800# gnd! 26.2fF
C491 diff_1558800_574800# gnd! 26.2fF
C492 diff_1538400_574800# gnd! 26.2fF
C493 diff_1518000_574800# gnd! 26.2fF
C494 diff_1497600_574800# gnd! 26.2fF
C495 diff_1477200_574800# gnd! 26.2fF
C496 diff_1456800_574800# gnd! 26.2fF
C497 diff_1436400_574800# gnd! 26.2fF
C498 diff_1416000_574800# gnd! 26.2fF
C499 diff_1395600_574800# gnd! 26.2fF
C500 diff_1375200_574800# gnd! 26.2fF
C501 diff_1354800_574800# gnd! 26.2fF
C502 diff_1334400_574800# gnd! 26.2fF
C503 diff_1314000_574800# gnd! 26.2fF
C504 diff_1293600_574800# gnd! 26.2fF
C505 diff_1273200_574800# gnd! 26.2fF
C506 diff_1252800_574800# gnd! 26.2fF
C507 diff_1232400_574800# gnd! 26.2fF
C508 diff_1212000_574800# gnd! 26.2fF
C509 diff_1191600_574800# gnd! 26.2fF
C510 diff_1171200_574800# gnd! 26.2fF
C511 diff_1150800_574800# gnd! 26.2fF
C512 diff_1130400_574800# gnd! 26.2fF
C513 diff_1110000_574800# gnd! 26.2fF
C514 diff_1089600_574800# gnd! 26.2fF
C515 diff_1069200_574800# gnd! 26.2fF
C516 diff_1048800_574800# gnd! 26.2fF
C517 diff_1028400_574800# gnd! 26.2fF
C518 diff_1008000_574800# gnd! 26.2fF
C519 diff_2367600_519600# gnd! 482.7fF
C520 diff_1004400_524400# gnd! 592.4fF
C521 diff_2508000_430800# gnd! 973.1fF
C522 diff_1004400_591600# gnd! 621.9fF
C523 diff_2293200_597600# gnd! 24.7fF
C524 diff_2272800_597600# gnd! 24.7fF
C525 diff_2252400_597600# gnd! 24.7fF
C526 diff_2232000_597600# gnd! 24.7fF
C527 diff_2211600_597600# gnd! 24.7fF
C528 diff_2191200_597600# gnd! 24.7fF
C529 diff_2170800_597600# gnd! 24.7fF
C530 diff_2150400_597600# gnd! 24.7fF
C531 diff_2130000_597600# gnd! 24.7fF
C532 diff_2109600_597600# gnd! 24.7fF
C533 diff_2089200_597600# gnd! 24.7fF
C534 diff_2068800_597600# gnd! 24.7fF
C535 diff_2048400_597600# gnd! 24.7fF
C536 diff_2028000_597600# gnd! 24.7fF
C537 diff_2007600_597600# gnd! 24.7fF
C538 diff_1987200_597600# gnd! 24.7fF
C539 diff_1966800_597600# gnd! 24.7fF
C540 diff_1946400_597600# gnd! 24.7fF
C541 diff_1926000_597600# gnd! 24.7fF
C542 diff_1905600_597600# gnd! 24.7fF
C543 diff_1885200_597600# gnd! 24.7fF
C544 diff_1864800_597600# gnd! 24.7fF
C545 diff_1844400_597600# gnd! 24.7fF
C546 diff_1824000_597600# gnd! 24.7fF
C547 diff_1803600_597600# gnd! 24.7fF
C548 diff_1783200_597600# gnd! 24.7fF
C549 diff_1762800_597600# gnd! 24.7fF
C550 diff_1742400_597600# gnd! 24.7fF
C551 diff_1722000_597600# gnd! 24.7fF
C552 diff_1701600_597600# gnd! 24.7fF
C553 diff_1681200_597600# gnd! 24.7fF
C554 diff_1660800_597600# gnd! 24.7fF
C555 diff_1640400_597600# gnd! 24.7fF
C556 diff_1620000_597600# gnd! 24.7fF
C557 diff_1599600_597600# gnd! 24.7fF
C558 diff_1579200_597600# gnd! 24.7fF
C559 diff_1558800_597600# gnd! 24.7fF
C560 diff_1538400_597600# gnd! 24.7fF
C561 diff_1518000_597600# gnd! 24.7fF
C562 diff_1497600_597600# gnd! 24.7fF
C563 diff_1477200_597600# gnd! 24.7fF
C564 diff_1456800_597600# gnd! 24.7fF
C565 diff_1436400_597600# gnd! 24.7fF
C566 diff_1416000_597600# gnd! 24.7fF
C567 diff_1395600_597600# gnd! 24.7fF
C568 diff_1375200_597600# gnd! 24.7fF
C569 diff_1354800_597600# gnd! 24.7fF
C570 diff_1334400_597600# gnd! 24.7fF
C571 diff_1314000_597600# gnd! 24.7fF
C572 diff_1293600_597600# gnd! 24.7fF
C573 diff_1273200_597600# gnd! 24.7fF
C574 diff_1252800_597600# gnd! 24.7fF
C575 diff_1232400_597600# gnd! 24.7fF
C576 diff_1212000_597600# gnd! 24.7fF
C577 diff_1191600_597600# gnd! 24.7fF
C578 diff_1171200_597600# gnd! 24.7fF
C579 diff_1150800_597600# gnd! 24.7fF
C580 diff_1130400_597600# gnd! 24.7fF
C581 diff_1110000_597600# gnd! 24.7fF
C582 diff_1089600_597600# gnd! 24.7fF
C583 diff_1069200_597600# gnd! 24.7fF
C584 diff_1048800_597600# gnd! 24.7fF
C585 diff_1028400_597600# gnd! 24.7fF
C586 diff_776400_488400# gnd! 105.8fF
C587 diff_691200_487200# gnd! 146.6fF
C588 diff_756000_454800# gnd! 104.1fF
C589 diff_1008000_597600# gnd! 24.7fF
C590 diff_694800_493200# gnd! 88.7fF
C591 diff_475200_500400# gnd! 15.4fF
C592 diff_404400_470400# gnd! 67.7fF
C593 diff_490800_500400# gnd! 51.7fF
C594 diff_478800_470400# gnd! 150.8fF
C595 diff_496800_492000# gnd! 357.1fF
C596 cm gnd! 1181.1fF
C597 diff_2367600_607200# gnd! 544.8fF
C598 diff_2293200_619200# gnd! 26.2fF
C599 diff_2272800_619200# gnd! 26.2fF
C600 diff_2252400_619200# gnd! 26.2fF
C601 diff_2232000_619200# gnd! 26.2fF
C602 diff_2211600_619200# gnd! 26.2fF
C603 diff_2191200_619200# gnd! 26.2fF
C604 diff_2170800_619200# gnd! 26.2fF
C605 diff_2150400_619200# gnd! 26.2fF
C606 diff_2130000_619200# gnd! 26.2fF
C607 diff_2109600_619200# gnd! 26.2fF
C608 diff_2089200_619200# gnd! 26.2fF
C609 diff_2068800_619200# gnd! 26.2fF
C610 diff_2048400_619200# gnd! 26.2fF
C611 diff_2028000_619200# gnd! 26.2fF
C612 diff_2007600_619200# gnd! 26.2fF
C613 diff_1987200_619200# gnd! 26.2fF
C614 diff_1966800_619200# gnd! 26.2fF
C615 diff_1946400_619200# gnd! 26.2fF
C616 diff_1926000_619200# gnd! 26.2fF
C617 diff_1905600_619200# gnd! 26.2fF
C618 diff_1885200_619200# gnd! 26.2fF
C619 diff_1864800_619200# gnd! 26.2fF
C620 diff_1844400_619200# gnd! 26.2fF
C621 diff_1824000_619200# gnd! 26.2fF
C622 diff_1803600_619200# gnd! 26.2fF
C623 diff_1783200_619200# gnd! 26.2fF
C624 diff_1762800_619200# gnd! 26.2fF
C625 diff_1742400_619200# gnd! 26.2fF
C626 diff_1722000_619200# gnd! 26.2fF
C627 diff_1701600_619200# gnd! 26.2fF
C628 diff_1681200_619200# gnd! 26.2fF
C629 diff_1660800_619200# gnd! 26.2fF
C630 diff_1640400_619200# gnd! 26.2fF
C631 diff_1620000_619200# gnd! 26.2fF
C632 diff_1599600_619200# gnd! 26.2fF
C633 diff_1579200_619200# gnd! 26.2fF
C634 diff_1558800_619200# gnd! 26.2fF
C635 diff_1538400_619200# gnd! 26.2fF
C636 diff_1518000_619200# gnd! 26.2fF
C637 diff_1497600_619200# gnd! 26.2fF
C638 diff_1477200_619200# gnd! 26.2fF
C639 diff_1456800_619200# gnd! 26.2fF
C640 diff_1436400_619200# gnd! 26.2fF
C641 diff_1416000_619200# gnd! 26.2fF
C642 diff_1395600_619200# gnd! 26.2fF
C643 diff_1375200_619200# gnd! 26.2fF
C644 diff_1354800_619200# gnd! 26.2fF
C645 diff_1334400_619200# gnd! 26.2fF
C646 diff_1314000_619200# gnd! 26.2fF
C647 diff_1293600_619200# gnd! 26.2fF
C648 diff_1273200_619200# gnd! 26.2fF
C649 diff_1252800_619200# gnd! 26.2fF
C650 diff_1232400_619200# gnd! 26.2fF
C651 diff_1212000_619200# gnd! 26.2fF
C652 diff_1191600_619200# gnd! 26.2fF
C653 diff_1171200_619200# gnd! 26.2fF
C654 diff_1150800_619200# gnd! 26.2fF
C655 diff_1130400_619200# gnd! 26.2fF
C656 diff_1110000_619200# gnd! 26.2fF
C657 diff_1089600_619200# gnd! 26.2fF
C658 diff_1069200_619200# gnd! 26.2fF
C659 diff_1048800_619200# gnd! 26.2fF
C660 diff_1028400_619200# gnd! 26.2fF
C661 diff_1008000_619200# gnd! 26.2fF
C662 diff_1004400_636000# gnd! 641.1fF
C663 diff_2293200_642000# gnd! 24.7fF
C664 diff_2272800_642000# gnd! 24.7fF
C665 diff_2252400_642000# gnd! 24.7fF
C666 diff_2232000_642000# gnd! 24.7fF
C667 diff_2211600_642000# gnd! 24.7fF
C668 diff_2191200_642000# gnd! 24.7fF
C669 diff_2170800_642000# gnd! 24.7fF
C670 diff_2150400_642000# gnd! 24.7fF
C671 diff_2130000_642000# gnd! 24.7fF
C672 diff_2109600_642000# gnd! 24.7fF
C673 diff_2089200_642000# gnd! 24.7fF
C674 diff_2068800_642000# gnd! 24.7fF
C675 diff_2048400_642000# gnd! 24.7fF
C676 diff_2028000_642000# gnd! 24.7fF
C677 diff_2007600_642000# gnd! 24.7fF
C678 diff_1987200_642000# gnd! 24.7fF
C679 diff_1966800_642000# gnd! 24.7fF
C680 diff_1946400_642000# gnd! 24.7fF
C681 diff_1926000_642000# gnd! 24.7fF
C682 diff_1905600_642000# gnd! 24.7fF
C683 diff_1885200_642000# gnd! 24.7fF
C684 diff_1864800_642000# gnd! 24.7fF
C685 diff_1844400_642000# gnd! 24.7fF
C686 diff_1824000_642000# gnd! 24.7fF
C687 diff_1803600_642000# gnd! 24.7fF
C688 diff_1783200_642000# gnd! 24.7fF
C689 diff_1762800_642000# gnd! 24.7fF
C690 diff_1742400_642000# gnd! 24.7fF
C691 diff_1722000_642000# gnd! 24.7fF
C692 diff_1701600_642000# gnd! 24.7fF
C693 diff_1681200_642000# gnd! 24.7fF
C694 diff_1660800_642000# gnd! 24.7fF
C695 diff_1640400_642000# gnd! 24.7fF
C696 diff_1620000_642000# gnd! 24.7fF
C697 diff_1599600_642000# gnd! 24.7fF
C698 diff_1579200_642000# gnd! 24.7fF
C699 diff_1558800_642000# gnd! 24.7fF
C700 diff_1538400_642000# gnd! 24.7fF
C701 diff_1518000_642000# gnd! 24.7fF
C702 diff_1497600_642000# gnd! 24.7fF
C703 diff_1477200_642000# gnd! 24.7fF
C704 diff_1456800_642000# gnd! 24.7fF
C705 diff_1436400_642000# gnd! 24.7fF
C706 diff_1416000_642000# gnd! 24.7fF
C707 diff_1395600_642000# gnd! 24.7fF
C708 diff_1375200_642000# gnd! 24.7fF
C709 diff_1354800_642000# gnd! 24.7fF
C710 diff_1334400_642000# gnd! 24.7fF
C711 diff_1314000_642000# gnd! 24.7fF
C712 diff_1293600_642000# gnd! 24.7fF
C713 diff_1273200_642000# gnd! 24.7fF
C714 diff_1252800_642000# gnd! 24.7fF
C715 diff_1232400_642000# gnd! 24.7fF
C716 diff_1212000_642000# gnd! 24.7fF
C717 diff_1191600_642000# gnd! 24.7fF
C718 diff_1171200_642000# gnd! 24.7fF
C719 diff_1150800_642000# gnd! 24.7fF
C720 diff_1130400_642000# gnd! 24.7fF
C721 diff_1110000_642000# gnd! 24.7fF
C722 diff_1089600_642000# gnd! 24.7fF
C723 diff_1069200_642000# gnd! 24.7fF
C724 diff_1048800_642000# gnd! 24.7fF
C725 diff_1028400_642000# gnd! 24.7fF
C726 diff_1008000_642000# gnd! 24.7fF
C727 diff_746400_625200# gnd! 237.2fF
C728 diff_1004400_657600# gnd! 652.7fF
C729 diff_2293200_663600# gnd! 26.2fF
C730 diff_2272800_663600# gnd! 26.2fF
C731 diff_2252400_663600# gnd! 26.2fF
C732 diff_2232000_663600# gnd! 26.2fF
C733 diff_2211600_663600# gnd! 26.2fF
C734 diff_2191200_663600# gnd! 26.2fF
C735 diff_2170800_663600# gnd! 26.2fF
C736 diff_2150400_663600# gnd! 26.2fF
C737 diff_2130000_663600# gnd! 26.2fF
C738 diff_2109600_663600# gnd! 26.2fF
C739 diff_2089200_663600# gnd! 26.2fF
C740 diff_2068800_663600# gnd! 26.2fF
C741 diff_2048400_663600# gnd! 26.2fF
C742 diff_2028000_663600# gnd! 26.2fF
C743 diff_2007600_663600# gnd! 26.2fF
C744 diff_1987200_663600# gnd! 26.2fF
C745 diff_1966800_663600# gnd! 26.2fF
C746 diff_1946400_663600# gnd! 26.2fF
C747 diff_1926000_663600# gnd! 26.2fF
C748 diff_1905600_663600# gnd! 26.2fF
C749 diff_1885200_663600# gnd! 26.2fF
C750 diff_1864800_663600# gnd! 26.2fF
C751 diff_1844400_663600# gnd! 26.2fF
C752 diff_1824000_663600# gnd! 26.2fF
C753 diff_1803600_663600# gnd! 26.2fF
C754 diff_1783200_663600# gnd! 26.2fF
C755 diff_1762800_663600# gnd! 26.2fF
C756 diff_1742400_663600# gnd! 26.2fF
C757 diff_1722000_663600# gnd! 26.2fF
C758 diff_1701600_663600# gnd! 26.2fF
C759 diff_1681200_663600# gnd! 26.2fF
C760 diff_1660800_663600# gnd! 26.2fF
C761 diff_1640400_663600# gnd! 26.2fF
C762 diff_1620000_663600# gnd! 26.2fF
C763 diff_1599600_663600# gnd! 26.2fF
C764 diff_1579200_663600# gnd! 26.2fF
C765 diff_1558800_663600# gnd! 26.2fF
C766 diff_1538400_663600# gnd! 26.2fF
C767 diff_1518000_663600# gnd! 26.2fF
C768 diff_1497600_663600# gnd! 26.2fF
C769 diff_1477200_663600# gnd! 26.2fF
C770 diff_1456800_663600# gnd! 26.2fF
C771 diff_1436400_663600# gnd! 26.2fF
C772 diff_1416000_663600# gnd! 26.2fF
C773 diff_1395600_663600# gnd! 26.2fF
C774 diff_1375200_663600# gnd! 26.2fF
C775 diff_1354800_663600# gnd! 26.2fF
C776 diff_1334400_663600# gnd! 26.2fF
C777 diff_1314000_663600# gnd! 26.2fF
C778 diff_1293600_663600# gnd! 26.2fF
C779 diff_1273200_663600# gnd! 26.2fF
C780 diff_1252800_663600# gnd! 26.2fF
C781 diff_1232400_663600# gnd! 26.2fF
C782 diff_1212000_663600# gnd! 26.2fF
C783 diff_1191600_663600# gnd! 26.2fF
C784 diff_1171200_663600# gnd! 26.2fF
C785 diff_1150800_663600# gnd! 26.2fF
C786 diff_1130400_663600# gnd! 26.2fF
C787 diff_1110000_663600# gnd! 26.2fF
C788 diff_1089600_663600# gnd! 26.2fF
C789 diff_1069200_663600# gnd! 26.2fF
C790 diff_1048800_663600# gnd! 26.2fF
C791 diff_1028400_663600# gnd! 26.2fF
C792 diff_891600_656400# gnd! 10.8fF
C793 diff_897600_638400# gnd! 124.6fF
C794 diff_1008000_663600# gnd! 26.2fF
C795 diff_1004400_613200# gnd! 597.6fF
C796 diff_1004400_680400# gnd! 622.9fF
C797 diff_2293200_686400# gnd! 24.7fF
C798 diff_2272800_686400# gnd! 24.7fF
C799 diff_2252400_686400# gnd! 24.7fF
C800 diff_2232000_686400# gnd! 24.7fF
C801 diff_2211600_686400# gnd! 24.7fF
C802 diff_2191200_686400# gnd! 24.7fF
C803 diff_2170800_686400# gnd! 24.7fF
C804 diff_2150400_686400# gnd! 24.7fF
C805 diff_2130000_686400# gnd! 24.7fF
C806 diff_2109600_686400# gnd! 24.7fF
C807 diff_2089200_686400# gnd! 24.7fF
C808 diff_2068800_686400# gnd! 24.7fF
C809 diff_2048400_686400# gnd! 24.7fF
C810 diff_2028000_686400# gnd! 24.7fF
C811 diff_2007600_686400# gnd! 24.7fF
C812 diff_1987200_686400# gnd! 24.7fF
C813 diff_1966800_686400# gnd! 24.7fF
C814 diff_1946400_686400# gnd! 24.7fF
C815 diff_1926000_686400# gnd! 24.7fF
C816 diff_1905600_686400# gnd! 24.7fF
C817 diff_1885200_686400# gnd! 24.7fF
C818 diff_1864800_686400# gnd! 24.7fF
C819 diff_1844400_686400# gnd! 24.7fF
C820 diff_1824000_686400# gnd! 24.7fF
C821 diff_1803600_686400# gnd! 24.7fF
C822 diff_1783200_686400# gnd! 24.7fF
C823 diff_1762800_686400# gnd! 24.7fF
C824 diff_1742400_686400# gnd! 24.7fF
C825 diff_1722000_686400# gnd! 24.7fF
C826 diff_1701600_686400# gnd! 24.7fF
C827 diff_1681200_686400# gnd! 24.7fF
C828 diff_1660800_686400# gnd! 24.7fF
C829 diff_1640400_686400# gnd! 24.7fF
C830 diff_1620000_686400# gnd! 24.7fF
C831 diff_1599600_686400# gnd! 24.7fF
C832 diff_1579200_686400# gnd! 24.7fF
C833 diff_1558800_686400# gnd! 24.7fF
C834 diff_1538400_686400# gnd! 24.7fF
C835 diff_1518000_686400# gnd! 24.7fF
C836 diff_1497600_686400# gnd! 24.7fF
C837 diff_1477200_686400# gnd! 24.7fF
C838 diff_1456800_686400# gnd! 24.7fF
C839 diff_1436400_686400# gnd! 24.7fF
C840 diff_1416000_686400# gnd! 24.7fF
C841 diff_1395600_686400# gnd! 24.7fF
C842 diff_1375200_686400# gnd! 24.7fF
C843 diff_1354800_686400# gnd! 24.7fF
C844 diff_1334400_686400# gnd! 24.7fF
C845 diff_1314000_686400# gnd! 24.7fF
C846 diff_1293600_686400# gnd! 24.7fF
C847 diff_1273200_686400# gnd! 24.7fF
C848 diff_1252800_686400# gnd! 24.7fF
C849 diff_1232400_686400# gnd! 24.7fF
C850 diff_1212000_686400# gnd! 24.7fF
C851 diff_1191600_686400# gnd! 24.7fF
C852 diff_1171200_686400# gnd! 24.7fF
C853 diff_1150800_686400# gnd! 24.7fF
C854 diff_1130400_686400# gnd! 24.7fF
C855 diff_1110000_686400# gnd! 24.7fF
C856 diff_1089600_686400# gnd! 24.7fF
C857 diff_1069200_686400# gnd! 24.7fF
C858 diff_1048800_686400# gnd! 24.7fF
C859 diff_1028400_686400# gnd! 24.7fF
C860 diff_1008000_686400# gnd! 24.7fF
C861 diff_2367600_696000# gnd! 481.1fF
C862 diff_2293200_708000# gnd! 26.2fF
C863 diff_2272800_708000# gnd! 26.2fF
C864 diff_2252400_708000# gnd! 26.2fF
C865 diff_2232000_708000# gnd! 26.2fF
C866 diff_2211600_708000# gnd! 26.2fF
C867 diff_2191200_708000# gnd! 26.2fF
C868 diff_2170800_708000# gnd! 26.2fF
C869 diff_2150400_708000# gnd! 26.2fF
C870 diff_2130000_708000# gnd! 26.2fF
C871 diff_2109600_708000# gnd! 26.2fF
C872 diff_2089200_708000# gnd! 26.2fF
C873 diff_2068800_708000# gnd! 26.2fF
C874 diff_2048400_708000# gnd! 26.2fF
C875 diff_2028000_708000# gnd! 26.2fF
C876 diff_2007600_708000# gnd! 26.2fF
C877 diff_1987200_708000# gnd! 26.2fF
C878 diff_1966800_708000# gnd! 26.2fF
C879 diff_1946400_708000# gnd! 26.2fF
C880 diff_1926000_708000# gnd! 26.2fF
C881 diff_1905600_708000# gnd! 26.2fF
C882 diff_1885200_708000# gnd! 26.2fF
C883 diff_1864800_708000# gnd! 26.2fF
C884 diff_1844400_708000# gnd! 26.2fF
C885 diff_1824000_708000# gnd! 26.2fF
C886 diff_1803600_708000# gnd! 26.2fF
C887 diff_1783200_708000# gnd! 26.2fF
C888 diff_1762800_708000# gnd! 26.2fF
C889 diff_1742400_708000# gnd! 26.2fF
C890 diff_1722000_708000# gnd! 26.2fF
C891 diff_1701600_708000# gnd! 26.2fF
C892 diff_1681200_708000# gnd! 26.2fF
C893 diff_1660800_708000# gnd! 26.2fF
C894 diff_1640400_708000# gnd! 26.2fF
C895 diff_1620000_708000# gnd! 26.2fF
C896 diff_1599600_708000# gnd! 26.2fF
C897 diff_1579200_708000# gnd! 26.2fF
C898 diff_1558800_708000# gnd! 26.2fF
C899 diff_1538400_708000# gnd! 26.2fF
C900 diff_1518000_708000# gnd! 26.2fF
C901 diff_1497600_708000# gnd! 26.2fF
C902 diff_1477200_708000# gnd! 26.2fF
C903 diff_1456800_708000# gnd! 26.2fF
C904 diff_1436400_708000# gnd! 26.2fF
C905 diff_1416000_708000# gnd! 26.2fF
C906 diff_1395600_708000# gnd! 26.2fF
C907 diff_1375200_708000# gnd! 26.2fF
C908 diff_1354800_708000# gnd! 26.2fF
C909 diff_1334400_708000# gnd! 26.2fF
C910 diff_1314000_708000# gnd! 26.2fF
C911 diff_1293600_708000# gnd! 26.2fF
C912 diff_1273200_708000# gnd! 26.2fF
C913 diff_1252800_708000# gnd! 26.2fF
C914 diff_1232400_708000# gnd! 26.2fF
C915 diff_1212000_708000# gnd! 26.2fF
C916 diff_1191600_708000# gnd! 26.2fF
C917 diff_1171200_708000# gnd! 26.2fF
C918 diff_1150800_708000# gnd! 26.2fF
C919 diff_1130400_708000# gnd! 26.2fF
C920 diff_1110000_708000# gnd! 26.2fF
C921 diff_1089600_708000# gnd! 26.2fF
C922 diff_1069200_708000# gnd! 26.2fF
C923 diff_1048800_708000# gnd! 26.2fF
C924 diff_1028400_708000# gnd! 26.2fF
C925 diff_904800_656400# gnd! 78.3fF
C926 diff_1008000_708000# gnd! 26.2fF
C927 diff_1004400_724800# gnd! 639.6fF
C928 diff_2293200_730800# gnd! 24.7fF
C929 diff_2272800_730800# gnd! 24.7fF
C930 diff_2252400_730800# gnd! 24.7fF
C931 diff_2232000_730800# gnd! 24.7fF
C932 diff_2211600_730800# gnd! 24.7fF
C933 diff_2191200_730800# gnd! 24.7fF
C934 diff_2170800_730800# gnd! 24.7fF
C935 diff_2150400_730800# gnd! 24.7fF
C936 diff_2130000_730800# gnd! 24.7fF
C937 diff_2109600_730800# gnd! 24.7fF
C938 diff_2089200_730800# gnd! 24.7fF
C939 diff_2068800_730800# gnd! 24.7fF
C940 diff_2048400_730800# gnd! 24.7fF
C941 diff_2028000_730800# gnd! 24.7fF
C942 diff_2007600_730800# gnd! 24.7fF
C943 diff_1987200_730800# gnd! 24.7fF
C944 diff_1966800_730800# gnd! 24.7fF
C945 diff_1946400_730800# gnd! 24.7fF
C946 diff_1926000_730800# gnd! 24.7fF
C947 diff_1905600_730800# gnd! 24.7fF
C948 diff_1885200_730800# gnd! 24.7fF
C949 diff_1864800_730800# gnd! 24.7fF
C950 diff_1844400_730800# gnd! 24.7fF
C951 diff_1824000_730800# gnd! 24.7fF
C952 diff_1803600_730800# gnd! 24.7fF
C953 diff_1783200_730800# gnd! 24.7fF
C954 diff_1762800_730800# gnd! 24.7fF
C955 diff_1742400_730800# gnd! 24.7fF
C956 diff_1722000_730800# gnd! 24.7fF
C957 diff_1701600_730800# gnd! 24.7fF
C958 diff_1681200_730800# gnd! 24.7fF
C959 diff_1660800_730800# gnd! 24.7fF
C960 diff_1640400_730800# gnd! 24.7fF
C961 diff_1620000_730800# gnd! 24.7fF
C962 diff_1599600_730800# gnd! 24.7fF
C963 diff_1579200_730800# gnd! 24.7fF
C964 diff_1558800_730800# gnd! 24.7fF
C965 diff_1538400_730800# gnd! 24.7fF
C966 diff_1518000_730800# gnd! 24.7fF
C967 diff_1497600_730800# gnd! 24.7fF
C968 diff_1477200_730800# gnd! 24.7fF
C969 diff_1456800_730800# gnd! 24.7fF
C970 diff_1436400_730800# gnd! 24.7fF
C971 diff_1416000_730800# gnd! 24.7fF
C972 diff_1395600_730800# gnd! 24.7fF
C973 diff_1375200_730800# gnd! 24.7fF
C974 diff_1354800_730800# gnd! 24.7fF
C975 diff_1334400_730800# gnd! 24.7fF
C976 diff_1314000_730800# gnd! 24.7fF
C977 diff_1293600_730800# gnd! 24.7fF
C978 diff_1273200_730800# gnd! 24.7fF
C979 diff_1252800_730800# gnd! 24.7fF
C980 diff_1232400_730800# gnd! 24.7fF
C981 diff_1212000_730800# gnd! 24.7fF
C982 diff_1191600_730800# gnd! 24.7fF
C983 diff_1171200_730800# gnd! 24.7fF
C984 diff_1150800_730800# gnd! 24.7fF
C985 diff_1130400_730800# gnd! 24.7fF
C986 diff_1110000_730800# gnd! 24.7fF
C987 diff_1089600_730800# gnd! 24.7fF
C988 diff_1069200_730800# gnd! 24.7fF
C989 diff_1048800_730800# gnd! 24.7fF
C990 diff_1028400_730800# gnd! 24.7fF
C991 diff_1008000_730800# gnd! 24.7fF
C992 diff_1004400_746400# gnd! 652.7fF
C993 diff_2293200_752400# gnd! 26.2fF
C994 diff_2272800_752400# gnd! 26.2fF
C995 diff_2252400_752400# gnd! 26.2fF
C996 diff_2232000_752400# gnd! 26.2fF
C997 diff_2211600_752400# gnd! 26.2fF
C998 diff_2191200_752400# gnd! 26.2fF
C999 diff_2170800_752400# gnd! 26.2fF
C1000 diff_2150400_752400# gnd! 26.2fF
C1001 diff_2130000_752400# gnd! 26.2fF
C1002 diff_2109600_752400# gnd! 26.2fF
C1003 diff_2089200_752400# gnd! 26.2fF
C1004 diff_2068800_752400# gnd! 26.2fF
C1005 diff_2048400_752400# gnd! 26.2fF
C1006 diff_2028000_752400# gnd! 26.2fF
C1007 diff_2007600_752400# gnd! 26.2fF
C1008 diff_1987200_752400# gnd! 26.2fF
C1009 diff_1966800_752400# gnd! 26.2fF
C1010 diff_1946400_752400# gnd! 26.2fF
C1011 diff_1926000_752400# gnd! 26.2fF
C1012 diff_1905600_752400# gnd! 26.2fF
C1013 diff_1885200_752400# gnd! 26.2fF
C1014 diff_1864800_752400# gnd! 26.2fF
C1015 diff_1844400_752400# gnd! 26.2fF
C1016 diff_1824000_752400# gnd! 26.2fF
C1017 diff_1803600_752400# gnd! 26.2fF
C1018 diff_1783200_752400# gnd! 26.2fF
C1019 diff_1762800_752400# gnd! 26.2fF
C1020 diff_1742400_752400# gnd! 26.2fF
C1021 diff_1722000_752400# gnd! 26.2fF
C1022 diff_1701600_752400# gnd! 26.2fF
C1023 diff_1681200_752400# gnd! 26.2fF
C1024 diff_1660800_752400# gnd! 26.2fF
C1025 diff_1640400_752400# gnd! 26.2fF
C1026 diff_1620000_752400# gnd! 26.2fF
C1027 diff_1599600_752400# gnd! 26.2fF
C1028 diff_1579200_752400# gnd! 26.2fF
C1029 diff_1558800_752400# gnd! 26.2fF
C1030 diff_1538400_752400# gnd! 26.2fF
C1031 diff_1518000_752400# gnd! 26.2fF
C1032 diff_1497600_752400# gnd! 26.2fF
C1033 diff_1477200_752400# gnd! 26.2fF
C1034 diff_1456800_752400# gnd! 26.2fF
C1035 diff_1436400_752400# gnd! 26.2fF
C1036 diff_1416000_752400# gnd! 26.2fF
C1037 diff_1395600_752400# gnd! 26.2fF
C1038 diff_1375200_752400# gnd! 26.2fF
C1039 diff_1354800_752400# gnd! 26.2fF
C1040 diff_1334400_752400# gnd! 26.2fF
C1041 diff_1314000_752400# gnd! 26.2fF
C1042 diff_1293600_752400# gnd! 26.2fF
C1043 diff_1273200_752400# gnd! 26.2fF
C1044 diff_1252800_752400# gnd! 26.2fF
C1045 diff_1232400_752400# gnd! 26.2fF
C1046 diff_1212000_752400# gnd! 26.2fF
C1047 diff_1191600_752400# gnd! 26.2fF
C1048 diff_1171200_752400# gnd! 26.2fF
C1049 diff_1150800_752400# gnd! 26.2fF
C1050 diff_1130400_752400# gnd! 26.2fF
C1051 diff_1110000_752400# gnd! 26.2fF
C1052 diff_1089600_752400# gnd! 26.2fF
C1053 diff_1069200_752400# gnd! 26.2fF
C1054 diff_1048800_752400# gnd! 26.2fF
C1055 diff_1028400_752400# gnd! 26.2fF
C1056 diff_1008000_752400# gnd! 26.2fF
C1057 diff_866400_691200# gnd! 97.8fF
C1058 diff_840000_375600# gnd! 212.4fF
C1059 diff_1004400_702000# gnd! 600.3fF
C1060 diff_2529600_894000# gnd! 107.9fF
C1061 diff_2738400_926400# gnd! 91.8fF
C1062 diff_2529600_915600# gnd! 106.8fF
C1063 diff_2832000_1056000# gnd! 244.8fF
C1064 diff_2832000_1075200# gnd! 75.7fF
C1065 diff_2774400_1002000# gnd! 185.6fF
C1066 diff_2738400_964800# gnd! 92.6fF
C1067 diff_2865600_1124400# gnd! 49.8fF
C1068 diff_2774400_1040400# gnd! 182.7fF
C1069 diff_2530800_968400# gnd! 101.7fF
C1070 diff_2530800_991200# gnd! 109.8fF
C1071 diff_2530800_1035600# gnd! 104.8fF
C1072 diff_2738400_1077600# gnd! 86.6fF
C1073 diff_2530800_1058400# gnd! 104.0fF
C1074 diff_2532000_1111200# gnd! 101.9fF
C1075 diff_2774400_1153200# gnd! 104.9fF
C1076 diff_2738400_1114800# gnd! 85.9fF
C1077 diff_2530800_1132800# gnd! 108.9fF
C1078 diff_2818800_1136400# gnd! 148.5fF
C1079 diff_2841600_1227600# gnd! 42.3fF
C1080 diff_2774400_1189200# gnd! 165.5fF
C1081 diff_2818800_1292400# gnd! 43.7fF
C1082 diff_2530800_1178400# gnd! 114.0fF
C1083 diff_2738400_1228800# gnd! 91.0fF
C1084 diff_2530800_1201200# gnd! 107.1fF
C1085 diff_1004400_769200# gnd! 622.9fF
C1086 diff_904800_769200# gnd! 128.8fF
C1087 diff_284400_465600# gnd! 58.9fF
C1088 diff_338400_375600# gnd! 430.5fF
C1089 reset gnd! 751.2fF
C1090 diff_480000_614400# gnd! 91.6fF
C1091 diff_498000_715200# gnd! 51.5fF
C1092 diff_694800_762000# gnd! 135.1fF
C1093 diff_2293200_775200# gnd! 41.3fF
C1094 diff_2272800_775200# gnd! 41.9fF
C1095 diff_2211600_775200# gnd! 41.3fF
C1096 diff_2191200_775200# gnd! 41.9fF
C1097 diff_2130000_775200# gnd! 41.3fF
C1098 diff_2109600_775200# gnd! 41.9fF
C1099 diff_2048400_775200# gnd! 41.3fF
C1100 diff_2028000_775200# gnd! 41.9fF
C1101 diff_1966800_775200# gnd! 41.3fF
C1102 diff_1946400_775200# gnd! 41.9fF
C1103 diff_1885200_775200# gnd! 41.3fF
C1104 diff_1864800_775200# gnd! 41.9fF
C1105 diff_1803600_775200# gnd! 41.3fF
C1106 diff_1783200_775200# gnd! 41.9fF
C1107 diff_1722000_775200# gnd! 41.3fF
C1108 diff_1701600_775200# gnd! 41.9fF
C1109 diff_1640400_775200# gnd! 41.3fF
C1110 diff_1620000_775200# gnd! 41.9fF
C1111 diff_1558800_775200# gnd! 41.3fF
C1112 diff_1538400_775200# gnd! 41.9fF
C1113 diff_1477200_775200# gnd! 41.3fF
C1114 diff_1456800_775200# gnd! 41.9fF
C1115 diff_1395600_775200# gnd! 41.3fF
C1116 diff_1375200_775200# gnd! 41.9fF
C1117 diff_1314000_775200# gnd! 41.3fF
C1118 diff_1293600_775200# gnd! 41.9fF
C1119 diff_1232400_775200# gnd! 41.3fF
C1120 diff_1212000_775200# gnd! 41.9fF
C1121 diff_1150800_775200# gnd! 41.3fF
C1122 diff_1130400_775200# gnd! 41.9fF
C1123 diff_1069200_775200# gnd! 40.3fF
C1124 diff_1048800_775200# gnd! 41.1fF
C1125 diff_816000_787200# gnd! 14.4fF
C1126 diff_696000_782400# gnd! 69.5fF
C1127 diff_700800_679200# gnd! 147.1fF
C1128 diff_694800_556800# gnd! 265.6fF
C1129 diff_919200_421200# gnd! 697.3fF
C1130 diff_825600_782400# gnd! 167.2fF
C1131 diff_2774400_1308000# gnd! 115.5fF
C1132 diff_2738400_1274400# gnd! 89.4fF
C1133 diff_2526000_1243200# gnd! 141.7fF
C1134 diff_2568000_1281600# gnd! 88.2fF
C1135 diff_2708400_1392000# gnd! 37.2fF
C1136 diff_2605200_1372800# gnd! 92.6fF
C1137 diff_2601600_1368000# gnd! 97.9fF
C1138 diff_2626800_1411200# gnd! 91.0fF
C1139 diff_2722800_844800# gnd! 365.9fF
C1140 diff_2767200_1456800# gnd! 49.5fF
C1141 diff_2589600_1464000# gnd! 78.8fF
C1142 diff_2812800_1134000# gnd! 303.0fF
C1143 diff_2768400_1497600# gnd! 49.5fF
C1144 diff_2768400_1540800# gnd! 48.3fF
C1145 diff_2252400_775200# gnd! 53.1fF
C1146 diff_2232000_775200# gnd! 53.0fF
C1147 diff_2258400_849600# gnd! 42.5fF
C1148 diff_2170800_775200# gnd! 53.1fF
C1149 diff_2150400_775200# gnd! 53.0fF
C1150 diff_2176800_849600# gnd! 42.5fF
C1151 diff_2089200_775200# gnd! 53.1fF
C1152 diff_2068800_775200# gnd! 53.0fF
C1153 diff_2095200_849600# gnd! 42.5fF
C1154 diff_2007600_775200# gnd! 53.1fF
C1155 diff_1987200_775200# gnd! 53.0fF
C1156 diff_2013600_849600# gnd! 42.5fF
C1157 diff_1926000_775200# gnd! 53.1fF
C1158 diff_1905600_775200# gnd! 53.0fF
C1159 diff_1932000_849600# gnd! 42.5fF
C1160 diff_1844400_775200# gnd! 53.1fF
C1161 diff_1824000_775200# gnd! 53.0fF
C1162 diff_1850400_849600# gnd! 42.5fF
C1163 diff_1762800_775200# gnd! 53.1fF
C1164 diff_1742400_775200# gnd! 53.0fF
C1165 diff_1768800_849600# gnd! 42.5fF
C1166 diff_1681200_775200# gnd! 53.1fF
C1167 diff_1660800_775200# gnd! 53.0fF
C1168 diff_1687200_849600# gnd! 42.5fF
C1169 diff_1599600_775200# gnd! 53.1fF
C1170 diff_1579200_775200# gnd! 53.0fF
C1171 diff_1605600_849600# gnd! 42.5fF
C1172 diff_1518000_775200# gnd! 53.1fF
C1173 diff_1497600_775200# gnd! 53.0fF
C1174 diff_1524000_849600# gnd! 42.5fF
C1175 diff_1436400_775200# gnd! 53.1fF
C1176 diff_1416000_775200# gnd! 53.0fF
C1177 diff_1442400_849600# gnd! 42.5fF
C1178 diff_1354800_775200# gnd! 53.1fF
C1179 diff_1334400_775200# gnd! 53.0fF
C1180 diff_1360800_849600# gnd! 42.5fF
C1181 diff_1273200_775200# gnd! 53.1fF
C1182 diff_1252800_775200# gnd! 53.0fF
C1183 diff_1279200_849600# gnd! 42.5fF
C1184 diff_1191600_775200# gnd! 53.1fF
C1185 diff_1171200_775200# gnd! 53.0fF
C1186 diff_1197600_849600# gnd! 42.5fF
C1187 diff_1110000_775200# gnd! 53.1fF
C1188 diff_1089600_775200# gnd! 53.0fF
C1189 diff_1116000_849600# gnd! 42.5fF
C1190 diff_558000_765600# gnd! 136.6fF
C1191 diff_421200_728400# gnd! 98.6fF
C1192 diff_536400_776400# gnd! 127.9fF
C1193 diff_339600_532800# gnd! 392.4fF
C1194 diff_409200_476400# gnd! 209.4fF
C1195 diff_1008000_775200# gnd! 47.9fF
C1196 diff_1033200_850800# gnd! 46.8fF
C1197 diff_1024800_849600# gnd! 55.4fF
C1198 diff_997200_836400# gnd! 103.4fF
C1199 diff_2217600_829200# gnd! 109.8fF
C1200 diff_2054400_829200# gnd! 112.1fF
C1201 diff_1891200_829200# gnd! 112.1fF
C1202 diff_1728000_829200# gnd! 112.3fF
C1203 diff_1564800_829200# gnd! 108.0fF
C1204 diff_1401600_829200# gnd! 108.0fF
C1205 diff_1238400_829200# gnd! 114.1fF
C1206 diff_1075200_826800# gnd! 112.7fF
C1207 diff_2136000_829200# gnd! 114.7fF
C1208 diff_2259600_907200# gnd! 122.5fF
C1209 diff_1972800_829200# gnd! 114.7fF
C1210 diff_2176800_907200# gnd! 127.3fF
C1211 diff_2095200_907200# gnd! 125.2fF
C1212 diff_2013600_907200# gnd! 127.3fF
C1213 diff_1809600_829200# gnd! 115.0fF
C1214 diff_1932000_907200# gnd! 125.2fF
C1215 diff_1851600_907200# gnd! 127.3fF
C1216 diff_1646400_829200# gnd! 110.9fF
C1217 diff_1770000_907200# gnd! 125.2fF
C1218 diff_1687200_908400# gnd! 123.3fF
C1219 diff_1483200_829200# gnd! 110.4fF
C1220 diff_1605600_908400# gnd! 121.2fF
C1221 diff_1524000_908400# gnd! 123.3fF
C1222 diff_1320000_829200# gnd! 117.5fF
C1223 diff_1442400_908400# gnd! 121.2fF
C1224 diff_1156800_829200# gnd! 114.7fF
C1225 diff_1278000_906000# gnd! 129.2fF
C1226 diff_1197600_907200# gnd! 127.3fF
C1227 diff_1036800_903600# gnd! 124.5fF
C1228 diff_1359600_906000# gnd! 129.6fF
C1229 diff_1116000_907200# gnd! 125.6fF
C1230 diff_2217600_927600# gnd! 111.9fF
C1231 diff_2134800_927600# gnd! 113.7fF
C1232 diff_2053200_927600# gnd! 113.1fF
C1233 diff_1971600_927600# gnd! 113.7fF
C1234 diff_1890000_927600# gnd! 113.1fF
C1235 diff_1809600_927600# gnd! 113.7fF
C1236 diff_1728000_927600# gnd! 113.1fF
C1237 diff_1645200_928800# gnd! 109.7fF
C1238 diff_1563600_928800# gnd! 109.2fF
C1239 diff_1482000_928800# gnd! 109.7fF
C1240 diff_1400400_928800# gnd! 109.2fF
C1241 diff_1317600_926400# gnd! 116.6fF
C1242 diff_1236000_926400# gnd! 117.1fF
C1243 diff_447600_771600# gnd! 78.1fF
C1244 diff_496800_798000# gnd! 136.7fF
C1245 diff_898800_888000# gnd! 111.5fF
C1246 diff_1155600_927600# gnd! 113.7fF
C1247 diff_1074000_927600# gnd! 113.1fF
C1248 diff_2299200_829200# gnd! 137.1fF
C1249 diff_2056800_907200# gnd! 259.2fF
C1250 diff_1893600_907200# gnd! 259.6fF
C1251 diff_1731600_907200# gnd! 260.2fF
C1252 diff_1567200_907200# gnd! 264.9fF
C1253 diff_1404000_907200# gnd! 263.6fF
C1254 diff_1239600_907200# gnd! 250.6fF
C1255 diff_1077600_907200# gnd! 257.7fF
C1256 diff_999600_896400# gnd! 314.6fF
C1257 diff_2221200_907200# gnd! 265.1fF
C1258 diff_2138400_908400# gnd! 288.9fF
C1259 diff_1975200_908400# gnd! 287.2fF
C1260 diff_1813200_908400# gnd! 289.6fF
C1261 diff_1648800_908400# gnd! 289.1fF
C1262 diff_1485600_907200# gnd! 293.2fF
C1263 diff_1321200_904800# gnd! 285.3fF
C1264 diff_1159200_908400# gnd! 282.6fF
C1265 diff_1124400_963600# gnd! 757.2fF
C1266 diff_801600_888000# gnd! 110.4fF
C1267 diff_481200_801600# gnd! 151.9fF
C1268 diff_646800_888000# gnd! 111.5fF
C1269 diff_411600_853200# gnd! 61.3fF
C1270 diff_567600_855600# gnd! 100.9fF
C1271 diff_1014000_962400# gnd! 823.9fF
C1272 diff_1996800_1008000# gnd! 296.7fF
C1273 diff_1670400_1008000# gnd! 331.5fF
C1274 diff_624000_475200# gnd! 849.3fF
C1275 diff_1344000_1008000# gnd! 290.6fF
C1276 diff_999600_1087200# gnd! 267.7fF
C1277 diff_494400_889200# gnd! 110.4fF
C1278 diff_829200_1039200# gnd! 391.8fF
C1279 diff_802800_967200# gnd! 130.1fF
C1280 diff_967200_1083600# gnd! 107.7fF
C1281 diff_901200_968400# gnd! 193.8fF
C1282 diff_2160000_985200# gnd! 470.1fF
C1283 diff_1996800_984000# gnd! 559.2fF
C1284 diff_564000_475200# gnd! 986.9fF
C1285 diff_1834800_984000# gnd! 529.8fF
C1286 diff_1670400_984000# gnd! 532.3fF
C1287 diff_1507200_984000# gnd! 574.9fF
C1288 diff_1342800_1122000# gnd! 548.7fF
C1289 diff_1180800_985200# gnd! 507.2fF
C1290 diff_411600_867600# gnd! 680.4fF
C1291 diff_682800_1034400# gnd! 407.4fF
C1292 diff_648000_967200# gnd! 120.0fF
C1293 diff_543600_1017600# gnd! 558.4fF
C1294 diff_496800_967200# gnd! 112.5fF
C1295 io0 gnd! 1985.2fF
C1296 diff_446400_902400# gnd! 452.9fF
C1297 diff_406800_692400# gnd! 589.3fF
C1298 io1 gnd! 2019.9fF
C1299 io2 gnd! 1863.1fF
C1300 io3 gnd! 1883.2fF
C1301 diff_1016400_968400# gnd! 534.7fF
C1302 diff_1011600_1153200# gnd! 800.4fF
C1303 diff_802800_1087200# gnd! 222.6fF
C1304 diff_648000_1087200# gnd! 221.8fF
C1305 diff_493200_1087200# gnd! 216.4fF
C1306 diff_337200_1087200# gnd! 216.7fF
C1307 diff_1063200_940800# gnd! 1157.4fF
C1308 diff_1033200_919200# gnd! 1257.7fF
C1309 diff_994800_1225200# gnd! 1372.5fF
C1310 diff_2221200_1206000# gnd! 269.5fF
C1311 diff_2258400_1266000# gnd! 42.2fF
C1312 diff_2138400_1207200# gnd! 294.8fF
C1313 diff_2217600_1180800# gnd! 105.1fF
C1314 diff_2176800_1266000# gnd! 42.2fF
C1315 diff_2056800_1207200# gnd! 257.9fF
C1316 diff_2134800_1180800# gnd! 106.6fF
C1317 diff_2095200_1266000# gnd! 42.2fF
C1318 diff_1975200_1207200# gnd! 291.9fF
C1319 diff_2053200_1180800# gnd! 106.2fF
C1320 diff_2013600_1266000# gnd! 42.2fF
C1321 diff_1893600_1207200# gnd! 257.9fF
C1322 diff_1971600_1180800# gnd! 106.6fF
C1323 diff_1932000_1266000# gnd! 42.2fF
C1324 diff_1813200_1207200# gnd! 290.2fF
C1325 diff_1890000_1180800# gnd! 106.2fF
C1326 diff_1850400_1266000# gnd! 42.2fF
C1327 diff_1731600_1207200# gnd! 258.3fF
C1328 diff_1809600_1180800# gnd! 106.6fF
C1329 diff_1768800_1266000# gnd! 42.2fF
C1330 diff_1648800_1206000# gnd! 292.5fF
C1331 diff_1728000_1180800# gnd! 106.2fF
C1332 diff_1687200_1266000# gnd! 42.2fF
C1333 diff_1567200_1206000# gnd! 264.0fF
C1334 diff_1645200_1180800# gnd! 102.6fF
C1335 diff_1605600_1266000# gnd! 42.2fF
C1336 diff_1485600_1206000# gnd! 296.4fF
C1337 diff_1563600_1180800# gnd! 102.2fF
C1338 diff_1524000_1266000# gnd! 42.2fF
C1339 diff_1404000_1206000# gnd! 264.0fF
C1340 diff_1482000_1180800# gnd! 102.6fF
C1341 diff_1442400_1266000# gnd! 42.2fF
C1342 diff_1321200_1208400# gnd! 290.3fF
C1343 diff_1400400_1180800# gnd! 102.2fF
C1344 diff_1360800_1266000# gnd! 42.2fF
C1345 diff_1239600_1208400# gnd! 250.3fF
C1346 diff_1317600_1180800# gnd! 107.6fF
C1347 diff_1279200_1266000# gnd! 42.2fF
C1348 diff_1159200_1207200# gnd! 285.7fF
C1349 diff_1236000_1180800# gnd! 110.2fF
C1350 diff_1197600_1266000# gnd! 42.2fF
C1351 diff_1077600_1207200# gnd! 258.2fF
C1352 diff_1155600_1180800# gnd! 106.6fF
C1353 diff_1116000_1266000# gnd! 42.2fF
C1354 diff_1074000_1180800# gnd! 106.2fF
C1355 diff_999600_1216800# gnd! 312.8fF
C1356 diff_1033200_1267200# gnd! 47.3fF
C1357 diff_1048800_846000# gnd! 1177.0fF
C1358 diff_2299200_1284000# gnd! 131.7fF
C1359 diff_2259600_1202400# gnd! 117.6fF
C1360 diff_2217600_1284000# gnd! 103.0fF
C1361 diff_2176800_1202400# gnd! 122.4fF
C1362 diff_2136000_1284000# gnd! 108.7fF
C1363 diff_2095200_1202400# gnd! 120.2fF
C1364 diff_2054400_1284000# gnd! 105.2fF
C1365 diff_2013600_1202400# gnd! 122.4fF
C1366 diff_1972800_1284000# gnd! 108.7fF
C1367 diff_1932000_1202400# gnd! 120.2fF
C1368 diff_1891200_1284000# gnd! 105.2fF
C1369 diff_1851600_1202400# gnd! 122.4fF
C1370 diff_1809600_1284000# gnd! 109.0fF
C1371 diff_1770000_1202400# gnd! 120.2fF
C1372 diff_1728000_1284000# gnd! 105.4fF
C1373 diff_1687200_1202400# gnd! 118.5fF
C1374 diff_1646400_1284000# gnd! 104.8fF
C1375 diff_1605600_1202400# gnd! 116.2fF
C1376 diff_1564800_1284000# gnd! 101.1fF
C1377 diff_1524000_1202400# gnd! 118.5fF
C1378 diff_1483200_1284000# gnd! 104.1fF
C1379 diff_1442400_1202400# gnd! 116.2fF
C1380 diff_1401600_1284000# gnd! 101.1fF
C1381 diff_1359600_1201200# gnd! 126.8fF
C1382 diff_1320000_1284000# gnd! 111.6fF
C1383 diff_1278000_1202400# gnd! 124.1fF
C1384 diff_1238400_1284000# gnd! 107.2fF
C1385 diff_1197600_1202400# gnd! 122.4fF
C1386 diff_1156800_1284000# gnd! 109.0fF
C1387 diff_1116000_1201200# gnd! 120.5fF
C1388 diff_1075200_1284000# gnd! 105.8fF
C1389 diff_1036800_1202400# gnd! 119.6fF
C1390 diff_1124400_1153200# gnd! 787.8fF
C1391 diff_260400_786000# gnd! 536.7fF
C1392 cl gnd! 1201.9fF
C1393 diff_997200_1236000# gnd! 98.6fF
C1394 diff_820800_1299600# gnd! 206.4fF
C1395 diff_936000_1282800# gnd! 24.3fF ;**FLOATING
C1396 diff_666000_1299600# gnd! 203.3fF
C1397 diff_801600_1170000# gnd! 309.1fF
C1398 diff_2293200_1281600# gnd! 42.9fF
C1399 diff_2272800_1321200# gnd! 43.5fF
C1400 diff_2252400_1262400# gnd! 54.6fF
C1401 diff_2232000_1321200# gnd! 54.5fF
C1402 diff_2211600_1281600# gnd! 42.9fF
C1403 diff_2191200_1321200# gnd! 43.5fF
C1404 diff_2170800_1262400# gnd! 54.6fF
C1405 diff_2150400_1321200# gnd! 54.5fF
C1406 diff_2130000_1281600# gnd! 42.9fF
C1407 diff_2109600_1321200# gnd! 43.5fF
C1408 diff_2089200_1262400# gnd! 54.6fF
C1409 diff_2068800_1321200# gnd! 54.5fF
C1410 diff_2048400_1281600# gnd! 42.9fF
C1411 diff_2028000_1321200# gnd! 43.5fF
C1412 diff_2007600_1262400# gnd! 54.6fF
C1413 diff_1987200_1321200# gnd! 54.5fF
C1414 diff_1966800_1281600# gnd! 42.9fF
C1415 diff_1946400_1321200# gnd! 43.5fF
C1416 diff_1926000_1262400# gnd! 54.6fF
C1417 diff_1905600_1321200# gnd! 54.5fF
C1418 diff_1885200_1281600# gnd! 42.9fF
C1419 diff_1864800_1321200# gnd! 43.5fF
C1420 diff_1844400_1262400# gnd! 54.6fF
C1421 diff_1824000_1321200# gnd! 54.5fF
C1422 diff_1803600_1281600# gnd! 42.9fF
C1423 diff_1783200_1321200# gnd! 43.5fF
C1424 diff_1762800_1262400# gnd! 54.6fF
C1425 diff_1742400_1321200# gnd! 54.5fF
C1426 diff_1722000_1281600# gnd! 42.9fF
C1427 diff_1701600_1321200# gnd! 43.5fF
C1428 diff_1681200_1262400# gnd! 54.6fF
C1429 diff_1660800_1321200# gnd! 54.5fF
C1430 diff_1640400_1281600# gnd! 42.9fF
C1431 diff_1620000_1321200# gnd! 43.5fF
C1432 diff_1599600_1262400# gnd! 54.6fF
C1433 diff_1579200_1321200# gnd! 54.5fF
C1434 diff_1558800_1281600# gnd! 42.9fF
C1435 diff_1538400_1321200# gnd! 43.5fF
C1436 diff_1518000_1262400# gnd! 54.6fF
C1437 diff_1497600_1321200# gnd! 54.5fF
C1438 diff_1477200_1281600# gnd! 42.9fF
C1439 diff_1456800_1321200# gnd! 43.5fF
C1440 diff_1436400_1262400# gnd! 54.6fF
C1441 diff_1416000_1321200# gnd! 54.5fF
C1442 diff_1395600_1281600# gnd! 42.9fF
C1443 diff_1375200_1321200# gnd! 43.5fF
C1444 diff_1354800_1262400# gnd! 54.6fF
C1445 diff_1334400_1321200# gnd! 54.5fF
C1446 diff_1314000_1281600# gnd! 42.9fF
C1447 diff_1293600_1321200# gnd! 43.5fF
C1448 diff_1273200_1262400# gnd! 54.6fF
C1449 diff_1252800_1321200# gnd! 54.5fF
C1450 diff_1232400_1281600# gnd! 42.9fF
C1451 diff_1212000_1321200# gnd! 43.5fF
C1452 diff_1191600_1262400# gnd! 54.6fF
C1453 diff_1171200_1321200# gnd! 54.5fF
C1454 diff_1150800_1281600# gnd! 42.9fF
C1455 diff_1130400_1321200# gnd! 43.5fF
C1456 diff_1110000_1262400# gnd! 54.6fF
C1457 diff_1089600_1321200# gnd! 54.5fF
C1458 diff_1069200_1281600# gnd! 41.8fF
C1459 diff_1048800_1322400# gnd! 42.6fF
C1460 diff_1024800_1263600# gnd! 56.9fF
C1461 diff_799200_1276800# gnd! 305.3fF
C1462 diff_508800_1299600# gnd! 206.6fF
C1463 diff_646800_1170000# gnd! 318.7fF
C1464 diff_644400_1276800# gnd! 304.3fF
C1465 diff_355200_1299600# gnd! 207.4fF
C1466 diff_492000_1170000# gnd! 308.5fF
C1467 diff_488400_1276800# gnd! 297.6fF
C1468 diff_336000_1170000# gnd! 309.9fF
C1469 diff_333600_1278000# gnd! 303.1fF
C1470 diff_280800_1316400# gnd! 63.5fF
C1471 diff_1008000_1320000# gnd! 50.4fF
C1472 diff_1004400_1346400# gnd! 613.8fF
C1473 diff_2293200_1352400# gnd! 26.2fF
C1474 diff_2272800_1352400# gnd! 26.2fF
C1475 diff_2252400_1352400# gnd! 26.2fF
C1476 diff_2232000_1352400# gnd! 26.2fF
C1477 diff_2211600_1352400# gnd! 26.2fF
C1478 diff_2191200_1352400# gnd! 26.2fF
C1479 diff_2170800_1352400# gnd! 26.2fF
C1480 diff_2150400_1352400# gnd! 26.2fF
C1481 diff_2130000_1352400# gnd! 26.2fF
C1482 diff_2109600_1352400# gnd! 26.2fF
C1483 diff_2089200_1352400# gnd! 26.2fF
C1484 diff_2068800_1352400# gnd! 26.2fF
C1485 diff_2048400_1352400# gnd! 26.2fF
C1486 diff_2028000_1352400# gnd! 26.2fF
C1487 diff_2007600_1352400# gnd! 26.2fF
C1488 diff_1987200_1352400# gnd! 26.2fF
C1489 diff_1966800_1352400# gnd! 26.2fF
C1490 diff_1946400_1352400# gnd! 26.2fF
C1491 diff_1926000_1352400# gnd! 26.2fF
C1492 diff_1905600_1352400# gnd! 26.2fF
C1493 diff_1885200_1352400# gnd! 26.2fF
C1494 diff_1864800_1352400# gnd! 26.2fF
C1495 diff_1844400_1352400# gnd! 26.2fF
C1496 diff_1824000_1352400# gnd! 26.2fF
C1497 diff_1803600_1352400# gnd! 26.2fF
C1498 diff_1783200_1352400# gnd! 26.2fF
C1499 diff_1762800_1352400# gnd! 26.2fF
C1500 diff_1742400_1352400# gnd! 26.2fF
C1501 diff_1722000_1352400# gnd! 26.2fF
C1502 diff_1701600_1352400# gnd! 26.2fF
C1503 diff_1681200_1352400# gnd! 26.2fF
C1504 diff_1660800_1352400# gnd! 26.2fF
C1505 diff_1640400_1352400# gnd! 26.2fF
C1506 diff_1620000_1352400# gnd! 26.2fF
C1507 diff_1599600_1352400# gnd! 26.2fF
C1508 diff_1579200_1352400# gnd! 26.2fF
C1509 diff_1558800_1352400# gnd! 26.2fF
C1510 diff_1538400_1352400# gnd! 26.2fF
C1511 diff_1518000_1352400# gnd! 26.2fF
C1512 diff_1497600_1352400# gnd! 26.2fF
C1513 diff_1477200_1352400# gnd! 26.2fF
C1514 diff_1456800_1352400# gnd! 26.2fF
C1515 diff_1436400_1352400# gnd! 26.2fF
C1516 diff_1416000_1352400# gnd! 26.2fF
C1517 diff_1395600_1352400# gnd! 26.2fF
C1518 diff_1375200_1352400# gnd! 26.2fF
C1519 diff_1354800_1352400# gnd! 26.2fF
C1520 diff_1334400_1352400# gnd! 26.2fF
C1521 diff_1314000_1352400# gnd! 26.2fF
C1522 diff_1293600_1352400# gnd! 26.2fF
C1523 diff_1273200_1352400# gnd! 26.2fF
C1524 diff_1252800_1352400# gnd! 26.2fF
C1525 diff_1232400_1352400# gnd! 26.2fF
C1526 diff_1212000_1352400# gnd! 26.2fF
C1527 diff_1191600_1352400# gnd! 26.2fF
C1528 diff_1171200_1352400# gnd! 26.2fF
C1529 diff_1150800_1352400# gnd! 26.2fF
C1530 diff_1130400_1352400# gnd! 26.2fF
C1531 diff_1110000_1352400# gnd! 26.2fF
C1532 diff_1089600_1352400# gnd! 26.2fF
C1533 diff_1069200_1352400# gnd! 26.2fF
C1534 diff_1048800_1352400# gnd! 26.2fF
C1535 diff_1028400_1352400# gnd! 26.2fF
C1536 diff_799200_1346400# gnd! 14.2fF
C1537 diff_644400_1346400# gnd! 14.2fF
C1538 diff_488400_1346400# gnd! 14.2fF
C1539 diff_333600_1346400# gnd! 14.2fF
C1540 diff_154800_822000# gnd! 664.1fF
C1541 diff_1008000_1352400# gnd! 26.2fF
C1542 diff_1004400_1369200# gnd! 644.8fF
C1543 diff_2293200_1375200# gnd! 24.7fF
C1544 diff_2272800_1375200# gnd! 24.7fF
C1545 diff_2252400_1375200# gnd! 24.7fF
C1546 diff_2232000_1375200# gnd! 24.7fF
C1547 diff_2211600_1375200# gnd! 24.7fF
C1548 diff_2191200_1375200# gnd! 24.7fF
C1549 diff_2170800_1375200# gnd! 24.7fF
C1550 diff_2150400_1375200# gnd! 24.7fF
C1551 diff_2130000_1375200# gnd! 24.7fF
C1552 diff_2109600_1375200# gnd! 24.7fF
C1553 diff_2089200_1375200# gnd! 24.7fF
C1554 diff_2068800_1375200# gnd! 24.7fF
C1555 diff_2048400_1375200# gnd! 24.7fF
C1556 diff_2028000_1375200# gnd! 24.7fF
C1557 diff_2007600_1375200# gnd! 24.7fF
C1558 diff_1987200_1375200# gnd! 24.7fF
C1559 diff_1966800_1375200# gnd! 24.7fF
C1560 diff_1946400_1375200# gnd! 24.7fF
C1561 diff_1926000_1375200# gnd! 24.7fF
C1562 diff_1905600_1375200# gnd! 24.7fF
C1563 diff_1885200_1375200# gnd! 24.7fF
C1564 diff_1864800_1375200# gnd! 24.7fF
C1565 diff_1844400_1375200# gnd! 24.7fF
C1566 diff_1824000_1375200# gnd! 24.7fF
C1567 diff_1803600_1375200# gnd! 24.7fF
C1568 diff_1783200_1375200# gnd! 24.7fF
C1569 diff_1762800_1375200# gnd! 24.7fF
C1570 diff_1742400_1375200# gnd! 24.7fF
C1571 diff_1722000_1375200# gnd! 24.7fF
C1572 diff_1701600_1375200# gnd! 24.7fF
C1573 diff_1681200_1375200# gnd! 24.7fF
C1574 diff_1660800_1375200# gnd! 24.7fF
C1575 diff_1640400_1375200# gnd! 24.7fF
C1576 diff_1620000_1375200# gnd! 24.7fF
C1577 diff_1599600_1375200# gnd! 24.7fF
C1578 diff_1579200_1375200# gnd! 24.7fF
C1579 diff_1558800_1375200# gnd! 24.7fF
C1580 diff_1538400_1375200# gnd! 24.7fF
C1581 diff_1518000_1375200# gnd! 24.7fF
C1582 diff_1497600_1375200# gnd! 24.7fF
C1583 diff_1477200_1375200# gnd! 24.7fF
C1584 diff_1456800_1375200# gnd! 24.7fF
C1585 diff_1436400_1375200# gnd! 24.7fF
C1586 diff_1416000_1375200# gnd! 24.7fF
C1587 diff_1395600_1375200# gnd! 24.7fF
C1588 diff_1375200_1375200# gnd! 24.7fF
C1589 diff_1354800_1375200# gnd! 24.7fF
C1590 diff_1334400_1375200# gnd! 24.7fF
C1591 diff_1314000_1375200# gnd! 24.7fF
C1592 diff_1293600_1375200# gnd! 24.7fF
C1593 diff_1273200_1375200# gnd! 24.7fF
C1594 diff_1252800_1375200# gnd! 24.7fF
C1595 diff_1232400_1375200# gnd! 24.7fF
C1596 diff_1212000_1375200# gnd! 24.7fF
C1597 diff_1191600_1375200# gnd! 24.7fF
C1598 diff_1171200_1375200# gnd! 24.7fF
C1599 diff_1150800_1375200# gnd! 24.7fF
C1600 diff_1130400_1375200# gnd! 24.7fF
C1601 diff_1110000_1375200# gnd! 24.7fF
C1602 diff_1089600_1375200# gnd! 24.7fF
C1603 diff_1069200_1375200# gnd! 24.7fF
C1604 diff_1048800_1375200# gnd! 24.7fF
C1605 diff_1028400_1375200# gnd! 24.7fF
C1606 diff_1008000_1375200# gnd! 24.7fF
C1607 diff_1004400_1390800# gnd! 649.5fF
C1608 diff_2367600_1407600# gnd! 500.4fF
C1609 diff_2293200_1396800# gnd! 26.2fF
C1610 diff_2272800_1396800# gnd! 26.2fF
C1611 diff_2252400_1396800# gnd! 26.2fF
C1612 diff_2232000_1396800# gnd! 26.2fF
C1613 diff_2211600_1396800# gnd! 26.2fF
C1614 diff_2191200_1396800# gnd! 26.2fF
C1615 diff_2170800_1396800# gnd! 26.2fF
C1616 diff_2150400_1396800# gnd! 26.2fF
C1617 diff_2130000_1396800# gnd! 26.2fF
C1618 diff_2109600_1396800# gnd! 26.2fF
C1619 diff_2089200_1396800# gnd! 26.2fF
C1620 diff_2068800_1396800# gnd! 26.2fF
C1621 diff_2048400_1396800# gnd! 26.2fF
C1622 diff_2028000_1396800# gnd! 26.2fF
C1623 diff_2007600_1396800# gnd! 26.2fF
C1624 diff_1987200_1396800# gnd! 26.2fF
C1625 diff_1966800_1396800# gnd! 26.2fF
C1626 diff_1946400_1396800# gnd! 26.2fF
C1627 diff_1926000_1396800# gnd! 26.2fF
C1628 diff_1905600_1396800# gnd! 26.2fF
C1629 diff_1885200_1396800# gnd! 26.2fF
C1630 diff_1864800_1396800# gnd! 26.2fF
C1631 diff_1844400_1396800# gnd! 26.2fF
C1632 diff_1824000_1396800# gnd! 26.2fF
C1633 diff_1803600_1396800# gnd! 26.2fF
C1634 diff_1783200_1396800# gnd! 26.2fF
C1635 diff_1762800_1396800# gnd! 26.2fF
C1636 diff_1742400_1396800# gnd! 26.2fF
C1637 diff_1722000_1396800# gnd! 26.2fF
C1638 diff_1701600_1396800# gnd! 26.2fF
C1639 diff_1681200_1396800# gnd! 26.2fF
C1640 diff_1660800_1396800# gnd! 26.2fF
C1641 diff_1640400_1396800# gnd! 26.2fF
C1642 diff_1620000_1396800# gnd! 26.2fF
C1643 diff_1599600_1396800# gnd! 26.2fF
C1644 diff_1579200_1396800# gnd! 26.2fF
C1645 diff_1558800_1396800# gnd! 26.2fF
C1646 diff_1538400_1396800# gnd! 26.2fF
C1647 diff_1518000_1396800# gnd! 26.2fF
C1648 diff_1497600_1396800# gnd! 26.2fF
C1649 diff_1477200_1396800# gnd! 26.2fF
C1650 diff_1456800_1396800# gnd! 26.2fF
C1651 diff_1436400_1396800# gnd! 26.2fF
C1652 diff_1416000_1396800# gnd! 26.2fF
C1653 diff_1395600_1396800# gnd! 26.2fF
C1654 diff_1375200_1396800# gnd! 26.2fF
C1655 diff_1354800_1396800# gnd! 26.2fF
C1656 diff_1334400_1396800# gnd! 26.2fF
C1657 diff_1314000_1396800# gnd! 26.2fF
C1658 diff_1293600_1396800# gnd! 26.2fF
C1659 diff_1273200_1396800# gnd! 26.2fF
C1660 diff_1252800_1396800# gnd! 26.2fF
C1661 diff_1232400_1396800# gnd! 26.2fF
C1662 diff_1212000_1396800# gnd! 26.2fF
C1663 diff_1191600_1396800# gnd! 26.2fF
C1664 diff_1171200_1396800# gnd! 26.2fF
C1665 diff_1150800_1396800# gnd! 26.2fF
C1666 diff_1130400_1396800# gnd! 26.2fF
C1667 diff_1110000_1396800# gnd! 26.2fF
C1668 diff_1089600_1396800# gnd! 26.2fF
C1669 diff_1069200_1396800# gnd! 26.2fF
C1670 diff_1048800_1396800# gnd! 26.2fF
C1671 diff_1028400_1396800# gnd! 26.2fF
C1672 diff_1008000_1396800# gnd! 26.2fF
C1673 diff_1004400_1413600# gnd! 609.5fF
C1674 diff_2293200_1419600# gnd! 24.7fF
C1675 diff_2272800_1419600# gnd! 24.7fF
C1676 diff_2252400_1419600# gnd! 24.7fF
C1677 diff_2232000_1419600# gnd! 24.7fF
C1678 diff_2211600_1419600# gnd! 24.7fF
C1679 diff_2191200_1419600# gnd! 24.7fF
C1680 diff_2170800_1419600# gnd! 24.7fF
C1681 diff_2150400_1419600# gnd! 24.7fF
C1682 diff_2130000_1419600# gnd! 24.7fF
C1683 diff_2109600_1419600# gnd! 24.7fF
C1684 diff_2089200_1419600# gnd! 24.7fF
C1685 diff_2068800_1419600# gnd! 24.7fF
C1686 diff_2048400_1419600# gnd! 24.7fF
C1687 diff_2028000_1419600# gnd! 24.7fF
C1688 diff_2007600_1419600# gnd! 24.7fF
C1689 diff_1987200_1419600# gnd! 24.7fF
C1690 diff_1966800_1419600# gnd! 24.7fF
C1691 diff_1946400_1419600# gnd! 24.7fF
C1692 diff_1926000_1419600# gnd! 24.7fF
C1693 diff_1905600_1419600# gnd! 24.7fF
C1694 diff_1885200_1419600# gnd! 24.7fF
C1695 diff_1864800_1419600# gnd! 24.7fF
C1696 diff_1844400_1419600# gnd! 24.7fF
C1697 diff_1824000_1419600# gnd! 24.7fF
C1698 diff_1803600_1419600# gnd! 24.7fF
C1699 diff_1783200_1419600# gnd! 24.7fF
C1700 diff_1762800_1419600# gnd! 24.7fF
C1701 diff_1742400_1419600# gnd! 24.7fF
C1702 diff_1722000_1419600# gnd! 24.7fF
C1703 diff_1701600_1419600# gnd! 24.7fF
C1704 diff_1681200_1419600# gnd! 24.7fF
C1705 diff_1660800_1419600# gnd! 24.7fF
C1706 diff_1640400_1419600# gnd! 24.7fF
C1707 diff_1620000_1419600# gnd! 24.7fF
C1708 diff_1599600_1419600# gnd! 24.7fF
C1709 diff_1579200_1419600# gnd! 24.7fF
C1710 diff_1558800_1419600# gnd! 24.7fF
C1711 diff_1538400_1419600# gnd! 24.7fF
C1712 diff_1518000_1419600# gnd! 24.7fF
C1713 diff_1497600_1419600# gnd! 24.7fF
C1714 diff_1477200_1419600# gnd! 24.7fF
C1715 diff_1456800_1419600# gnd! 24.7fF
C1716 diff_1436400_1419600# gnd! 24.7fF
C1717 diff_1416000_1419600# gnd! 24.7fF
C1718 diff_1395600_1419600# gnd! 24.7fF
C1719 diff_1375200_1419600# gnd! 24.7fF
C1720 diff_1354800_1419600# gnd! 24.7fF
C1721 diff_1334400_1419600# gnd! 24.7fF
C1722 diff_1314000_1419600# gnd! 24.7fF
C1723 diff_1293600_1419600# gnd! 24.7fF
C1724 diff_1273200_1419600# gnd! 24.7fF
C1725 diff_1252800_1419600# gnd! 24.7fF
C1726 diff_1232400_1419600# gnd! 24.7fF
C1727 diff_1212000_1419600# gnd! 24.7fF
C1728 diff_1191600_1419600# gnd! 24.7fF
C1729 diff_1171200_1419600# gnd! 24.7fF
C1730 diff_1150800_1419600# gnd! 24.7fF
C1731 diff_1130400_1419600# gnd! 24.7fF
C1732 diff_1110000_1419600# gnd! 24.7fF
C1733 diff_1089600_1419600# gnd! 24.7fF
C1734 diff_1069200_1419600# gnd! 24.7fF
C1735 diff_1048800_1419600# gnd! 24.7fF
C1736 diff_1028400_1419600# gnd! 24.7fF
C1737 diff_1008000_1419600# gnd! 24.7fF
C1738 diff_1004400_1435200# gnd! 614.5fF
C1739 diff_2293200_1441200# gnd! 26.2fF
C1740 diff_2272800_1441200# gnd! 26.2fF
C1741 diff_2252400_1441200# gnd! 26.2fF
C1742 diff_2232000_1441200# gnd! 26.2fF
C1743 diff_2211600_1441200# gnd! 26.2fF
C1744 diff_2191200_1441200# gnd! 26.2fF
C1745 diff_2170800_1441200# gnd! 26.2fF
C1746 diff_2150400_1441200# gnd! 26.2fF
C1747 diff_2130000_1441200# gnd! 26.2fF
C1748 diff_2109600_1441200# gnd! 26.2fF
C1749 diff_2089200_1441200# gnd! 26.2fF
C1750 diff_2068800_1441200# gnd! 26.2fF
C1751 diff_2048400_1441200# gnd! 26.2fF
C1752 diff_2028000_1441200# gnd! 26.2fF
C1753 diff_2007600_1441200# gnd! 26.2fF
C1754 diff_1987200_1441200# gnd! 26.2fF
C1755 diff_1966800_1441200# gnd! 26.2fF
C1756 diff_1946400_1441200# gnd! 26.2fF
C1757 diff_1926000_1441200# gnd! 26.2fF
C1758 diff_1905600_1441200# gnd! 26.2fF
C1759 diff_1885200_1441200# gnd! 26.2fF
C1760 diff_1864800_1441200# gnd! 26.2fF
C1761 diff_1844400_1441200# gnd! 26.2fF
C1762 diff_1824000_1441200# gnd! 26.2fF
C1763 diff_1803600_1441200# gnd! 26.2fF
C1764 diff_1783200_1441200# gnd! 26.2fF
C1765 diff_1762800_1441200# gnd! 26.2fF
C1766 diff_1742400_1441200# gnd! 26.2fF
C1767 diff_1722000_1441200# gnd! 26.2fF
C1768 diff_1701600_1441200# gnd! 26.2fF
C1769 diff_1681200_1441200# gnd! 26.2fF
C1770 diff_1660800_1441200# gnd! 26.2fF
C1771 diff_1640400_1441200# gnd! 26.2fF
C1772 diff_1620000_1441200# gnd! 26.2fF
C1773 diff_1599600_1441200# gnd! 26.2fF
C1774 diff_1579200_1441200# gnd! 26.2fF
C1775 diff_1558800_1441200# gnd! 26.2fF
C1776 diff_1538400_1441200# gnd! 26.2fF
C1777 diff_1518000_1441200# gnd! 26.2fF
C1778 diff_1497600_1441200# gnd! 26.2fF
C1779 diff_1477200_1441200# gnd! 26.2fF
C1780 diff_1456800_1441200# gnd! 26.2fF
C1781 diff_1436400_1441200# gnd! 26.2fF
C1782 diff_1416000_1441200# gnd! 26.2fF
C1783 diff_1395600_1441200# gnd! 26.2fF
C1784 diff_1375200_1441200# gnd! 26.2fF
C1785 diff_1354800_1441200# gnd! 26.2fF
C1786 diff_1334400_1441200# gnd! 26.2fF
C1787 diff_1314000_1441200# gnd! 26.2fF
C1788 diff_1293600_1441200# gnd! 26.2fF
C1789 diff_1273200_1441200# gnd! 26.2fF
C1790 diff_1252800_1441200# gnd! 26.2fF
C1791 diff_1232400_1441200# gnd! 26.2fF
C1792 diff_1212000_1441200# gnd! 26.2fF
C1793 diff_1191600_1441200# gnd! 26.2fF
C1794 diff_1171200_1441200# gnd! 26.2fF
C1795 diff_1150800_1441200# gnd! 26.2fF
C1796 diff_1130400_1441200# gnd! 26.2fF
C1797 diff_1110000_1441200# gnd! 26.2fF
C1798 diff_1089600_1441200# gnd! 26.2fF
C1799 diff_1069200_1441200# gnd! 26.2fF
C1800 diff_1048800_1441200# gnd! 26.2fF
C1801 diff_1028400_1441200# gnd! 26.2fF
C1802 diff_1008000_1441200# gnd! 26.2fF
C1803 diff_1004400_1458000# gnd! 646.1fF
C1804 diff_2293200_1464000# gnd! 24.7fF
C1805 diff_2272800_1464000# gnd! 24.7fF
C1806 diff_2252400_1464000# gnd! 24.7fF
C1807 diff_2232000_1464000# gnd! 24.7fF
C1808 diff_2211600_1464000# gnd! 24.7fF
C1809 diff_2191200_1464000# gnd! 24.7fF
C1810 diff_2170800_1464000# gnd! 24.7fF
C1811 diff_2150400_1464000# gnd! 24.7fF
C1812 diff_2130000_1464000# gnd! 24.7fF
C1813 diff_2109600_1464000# gnd! 24.7fF
C1814 diff_2089200_1464000# gnd! 24.7fF
C1815 diff_2068800_1464000# gnd! 24.7fF
C1816 diff_2048400_1464000# gnd! 24.7fF
C1817 diff_2028000_1464000# gnd! 24.7fF
C1818 diff_2007600_1464000# gnd! 24.7fF
C1819 diff_1987200_1464000# gnd! 24.7fF
C1820 diff_1966800_1464000# gnd! 24.7fF
C1821 diff_1946400_1464000# gnd! 24.7fF
C1822 diff_1926000_1464000# gnd! 24.7fF
C1823 diff_1905600_1464000# gnd! 24.7fF
C1824 diff_1885200_1464000# gnd! 24.7fF
C1825 diff_1864800_1464000# gnd! 24.7fF
C1826 diff_1844400_1464000# gnd! 24.7fF
C1827 diff_1824000_1464000# gnd! 24.7fF
C1828 diff_1803600_1464000# gnd! 24.7fF
C1829 diff_1783200_1464000# gnd! 24.7fF
C1830 diff_1762800_1464000# gnd! 24.7fF
C1831 diff_1742400_1464000# gnd! 24.7fF
C1832 diff_1722000_1464000# gnd! 24.7fF
C1833 diff_1701600_1464000# gnd! 24.7fF
C1834 diff_1681200_1464000# gnd! 24.7fF
C1835 diff_1660800_1464000# gnd! 24.7fF
C1836 diff_1640400_1464000# gnd! 24.7fF
C1837 diff_1620000_1464000# gnd! 24.7fF
C1838 diff_1599600_1464000# gnd! 24.7fF
C1839 diff_1579200_1464000# gnd! 24.7fF
C1840 diff_1558800_1464000# gnd! 24.7fF
C1841 diff_1538400_1464000# gnd! 24.7fF
C1842 diff_1518000_1464000# gnd! 24.7fF
C1843 diff_1497600_1464000# gnd! 24.7fF
C1844 diff_1477200_1464000# gnd! 24.7fF
C1845 diff_1456800_1464000# gnd! 24.7fF
C1846 diff_1436400_1464000# gnd! 24.7fF
C1847 diff_1416000_1464000# gnd! 24.7fF
C1848 diff_1395600_1464000# gnd! 24.7fF
C1849 diff_1375200_1464000# gnd! 24.7fF
C1850 diff_1354800_1464000# gnd! 24.7fF
C1851 diff_1334400_1464000# gnd! 24.7fF
C1852 diff_1314000_1464000# gnd! 24.7fF
C1853 diff_1293600_1464000# gnd! 24.7fF
C1854 diff_1273200_1464000# gnd! 24.7fF
C1855 diff_1252800_1464000# gnd! 24.7fF
C1856 diff_1232400_1464000# gnd! 24.7fF
C1857 diff_1212000_1464000# gnd! 24.7fF
C1858 diff_1191600_1464000# gnd! 24.7fF
C1859 diff_1171200_1464000# gnd! 24.7fF
C1860 diff_1150800_1464000# gnd! 24.7fF
C1861 diff_1130400_1464000# gnd! 24.7fF
C1862 diff_1110000_1464000# gnd! 24.7fF
C1863 diff_1089600_1464000# gnd! 24.7fF
C1864 diff_1069200_1464000# gnd! 24.7fF
C1865 diff_1048800_1464000# gnd! 24.7fF
C1866 diff_1028400_1464000# gnd! 24.7fF
C1867 diff_1008000_1464000# gnd! 24.7fF
C1868 diff_1004400_1479600# gnd! 650.3fF
C1869 diff_2451600_979200# gnd! 624.8fF
C1870 diff_2469600_912000# gnd! 639.2fF
C1871 diff_2592000_1532400# gnd! 78.7fF
C1872 diff_2812800_1003200# gnd! 664.5fF
C1873 diff_2767200_1582800# gnd! 54.0fF
C1874 diff_2710800_1356000# gnd! 535.5fF
C1875 diff_2828400_1273200# gnd! 309.1fF
C1876 diff_2828400_1086000# gnd! 573.8fF
C1877 diff_2682000_1690800# gnd! 53.5fF
C1878 diff_2649600_1519200# gnd! 381.4fF
C1879 diff_2743200_1702800# gnd! 55.8fF
C1880 diff_2664000_1422000# gnd! 332.6fF
C1881 diff_2743200_1714800# gnd! 49.2fF
C1882 diff_2367600_1494000# gnd! 529.2fF
C1883 diff_2293200_1485600# gnd! 26.2fF
C1884 diff_2272800_1485600# gnd! 26.2fF
C1885 diff_2252400_1485600# gnd! 26.2fF
C1886 diff_2232000_1485600# gnd! 26.2fF
C1887 diff_2211600_1485600# gnd! 26.2fF
C1888 diff_2191200_1485600# gnd! 26.2fF
C1889 diff_2170800_1485600# gnd! 26.2fF
C1890 diff_2150400_1485600# gnd! 26.2fF
C1891 diff_2130000_1485600# gnd! 26.2fF
C1892 diff_2109600_1485600# gnd! 26.2fF
C1893 diff_2089200_1485600# gnd! 26.2fF
C1894 diff_2068800_1485600# gnd! 26.2fF
C1895 diff_2048400_1485600# gnd! 26.2fF
C1896 diff_2028000_1485600# gnd! 26.2fF
C1897 diff_2007600_1485600# gnd! 26.2fF
C1898 diff_1987200_1485600# gnd! 26.2fF
C1899 diff_1966800_1485600# gnd! 26.2fF
C1900 diff_1946400_1485600# gnd! 26.2fF
C1901 diff_1926000_1485600# gnd! 26.2fF
C1902 diff_1905600_1485600# gnd! 26.2fF
C1903 diff_1885200_1485600# gnd! 26.2fF
C1904 diff_1864800_1485600# gnd! 26.2fF
C1905 diff_1844400_1485600# gnd! 26.2fF
C1906 diff_1824000_1485600# gnd! 26.2fF
C1907 diff_1803600_1485600# gnd! 26.2fF
C1908 diff_1783200_1485600# gnd! 26.2fF
C1909 diff_1762800_1485600# gnd! 26.2fF
C1910 diff_1742400_1485600# gnd! 26.2fF
C1911 diff_1722000_1485600# gnd! 26.2fF
C1912 diff_1701600_1485600# gnd! 26.2fF
C1913 diff_1681200_1485600# gnd! 26.2fF
C1914 diff_1660800_1485600# gnd! 26.2fF
C1915 diff_1640400_1485600# gnd! 26.2fF
C1916 diff_1620000_1485600# gnd! 26.2fF
C1917 diff_1599600_1485600# gnd! 26.2fF
C1918 diff_1579200_1485600# gnd! 26.2fF
C1919 diff_1558800_1485600# gnd! 26.2fF
C1920 diff_1538400_1485600# gnd! 26.2fF
C1921 diff_1518000_1485600# gnd! 26.2fF
C1922 diff_1497600_1485600# gnd! 26.2fF
C1923 diff_1477200_1485600# gnd! 26.2fF
C1924 diff_1456800_1485600# gnd! 26.2fF
C1925 diff_1436400_1485600# gnd! 26.2fF
C1926 diff_1416000_1485600# gnd! 26.2fF
C1927 diff_1395600_1485600# gnd! 26.2fF
C1928 diff_1375200_1485600# gnd! 26.2fF
C1929 diff_1354800_1485600# gnd! 26.2fF
C1930 diff_1334400_1485600# gnd! 26.2fF
C1931 diff_1314000_1485600# gnd! 26.2fF
C1932 diff_1293600_1485600# gnd! 26.2fF
C1933 diff_1273200_1485600# gnd! 26.2fF
C1934 diff_1252800_1485600# gnd! 26.2fF
C1935 diff_1232400_1485600# gnd! 26.2fF
C1936 diff_1212000_1485600# gnd! 26.2fF
C1937 diff_1191600_1485600# gnd! 26.2fF
C1938 diff_1171200_1485600# gnd! 26.2fF
C1939 diff_1150800_1485600# gnd! 26.2fF
C1940 diff_1130400_1485600# gnd! 26.2fF
C1941 diff_1110000_1485600# gnd! 26.2fF
C1942 diff_1089600_1485600# gnd! 26.2fF
C1943 diff_1069200_1485600# gnd! 26.2fF
C1944 diff_1048800_1485600# gnd! 26.2fF
C1945 diff_1028400_1485600# gnd! 26.2fF
C1946 diff_873600_1448400# gnd! 106.6fF
C1947 diff_1008000_1485600# gnd! 26.2fF
C1948 diff_718800_1448400# gnd! 309.7fF
C1949 diff_1004400_1502400# gnd! 606.7fF
C1950 diff_2293200_1508400# gnd! 24.7fF
C1951 diff_2272800_1508400# gnd! 24.7fF
C1952 diff_2252400_1508400# gnd! 24.7fF
C1953 diff_2232000_1508400# gnd! 24.7fF
C1954 diff_2211600_1508400# gnd! 24.7fF
C1955 diff_2191200_1508400# gnd! 24.7fF
C1956 diff_2170800_1508400# gnd! 24.7fF
C1957 diff_2150400_1508400# gnd! 24.7fF
C1958 diff_2130000_1508400# gnd! 24.7fF
C1959 diff_2109600_1508400# gnd! 24.7fF
C1960 diff_2089200_1508400# gnd! 24.7fF
C1961 diff_2068800_1508400# gnd! 24.7fF
C1962 diff_2048400_1508400# gnd! 24.7fF
C1963 diff_2028000_1508400# gnd! 24.7fF
C1964 diff_2007600_1508400# gnd! 24.7fF
C1965 diff_1987200_1508400# gnd! 24.7fF
C1966 diff_1966800_1508400# gnd! 24.7fF
C1967 diff_1946400_1508400# gnd! 24.7fF
C1968 diff_1926000_1508400# gnd! 24.7fF
C1969 diff_1905600_1508400# gnd! 24.7fF
C1970 diff_1885200_1508400# gnd! 24.7fF
C1971 diff_1864800_1508400# gnd! 24.7fF
C1972 diff_1844400_1508400# gnd! 24.7fF
C1973 diff_1824000_1508400# gnd! 24.7fF
C1974 diff_1803600_1508400# gnd! 24.7fF
C1975 diff_1783200_1508400# gnd! 24.7fF
C1976 diff_1762800_1508400# gnd! 24.7fF
C1977 diff_1742400_1508400# gnd! 24.7fF
C1978 diff_1722000_1508400# gnd! 24.7fF
C1979 diff_1701600_1508400# gnd! 24.7fF
C1980 diff_1681200_1508400# gnd! 24.7fF
C1981 diff_1660800_1508400# gnd! 24.7fF
C1982 diff_1640400_1508400# gnd! 24.7fF
C1983 diff_1620000_1508400# gnd! 24.7fF
C1984 diff_1599600_1508400# gnd! 24.7fF
C1985 diff_1579200_1508400# gnd! 24.7fF
C1986 diff_1558800_1508400# gnd! 24.7fF
C1987 diff_1538400_1508400# gnd! 24.7fF
C1988 diff_1518000_1508400# gnd! 24.7fF
C1989 diff_1497600_1508400# gnd! 24.7fF
C1990 diff_1477200_1508400# gnd! 24.7fF
C1991 diff_1456800_1508400# gnd! 24.7fF
C1992 diff_1436400_1508400# gnd! 24.7fF
C1993 diff_1416000_1508400# gnd! 24.7fF
C1994 diff_1395600_1508400# gnd! 24.7fF
C1995 diff_1375200_1508400# gnd! 24.7fF
C1996 diff_1354800_1508400# gnd! 24.7fF
C1997 diff_1334400_1508400# gnd! 24.7fF
C1998 diff_1314000_1508400# gnd! 24.7fF
C1999 diff_1293600_1508400# gnd! 24.7fF
C2000 diff_1273200_1508400# gnd! 24.7fF
C2001 diff_1252800_1508400# gnd! 24.7fF
C2002 diff_1232400_1508400# gnd! 24.7fF
C2003 diff_1212000_1508400# gnd! 24.7fF
C2004 diff_1191600_1508400# gnd! 24.7fF
C2005 diff_1171200_1508400# gnd! 24.7fF
C2006 diff_1150800_1508400# gnd! 24.7fF
C2007 diff_1130400_1508400# gnd! 24.7fF
C2008 diff_1110000_1508400# gnd! 24.7fF
C2009 diff_1089600_1508400# gnd! 24.7fF
C2010 diff_1069200_1508400# gnd! 24.7fF
C2011 diff_1048800_1508400# gnd! 24.7fF
C2012 diff_1028400_1508400# gnd! 24.7fF
C2013 diff_1008000_1508400# gnd! 24.7fF
C2014 diff_1004400_1524000# gnd! 614.7fF
C2015 diff_2293200_1530000# gnd! 26.2fF
C2016 diff_2272800_1530000# gnd! 26.2fF
C2017 diff_2252400_1530000# gnd! 26.2fF
C2018 diff_2232000_1530000# gnd! 26.2fF
C2019 diff_2211600_1530000# gnd! 26.2fF
C2020 diff_2191200_1530000# gnd! 26.2fF
C2021 diff_2170800_1530000# gnd! 26.2fF
C2022 diff_2150400_1530000# gnd! 26.2fF
C2023 diff_2130000_1530000# gnd! 26.2fF
C2024 diff_2109600_1530000# gnd! 26.2fF
C2025 diff_2089200_1530000# gnd! 26.2fF
C2026 diff_2068800_1530000# gnd! 26.2fF
C2027 diff_2048400_1530000# gnd! 26.2fF
C2028 diff_2028000_1530000# gnd! 26.2fF
C2029 diff_2007600_1530000# gnd! 26.2fF
C2030 diff_1987200_1530000# gnd! 26.2fF
C2031 diff_1966800_1530000# gnd! 26.2fF
C2032 diff_1946400_1530000# gnd! 26.2fF
C2033 diff_1926000_1530000# gnd! 26.2fF
C2034 diff_1905600_1530000# gnd! 26.2fF
C2035 diff_1885200_1530000# gnd! 26.2fF
C2036 diff_1864800_1530000# gnd! 26.2fF
C2037 diff_1844400_1530000# gnd! 26.2fF
C2038 diff_1824000_1530000# gnd! 26.2fF
C2039 diff_1803600_1530000# gnd! 26.2fF
C2040 diff_1783200_1530000# gnd! 26.2fF
C2041 diff_1762800_1530000# gnd! 26.2fF
C2042 diff_1742400_1530000# gnd! 26.2fF
C2043 diff_1722000_1530000# gnd! 26.2fF
C2044 diff_1701600_1530000# gnd! 26.2fF
C2045 diff_1681200_1530000# gnd! 26.2fF
C2046 diff_1660800_1530000# gnd! 26.2fF
C2047 diff_1640400_1530000# gnd! 26.2fF
C2048 diff_1620000_1530000# gnd! 26.2fF
C2049 diff_1599600_1530000# gnd! 26.2fF
C2050 diff_1579200_1530000# gnd! 26.2fF
C2051 diff_1558800_1530000# gnd! 26.2fF
C2052 diff_1538400_1530000# gnd! 26.2fF
C2053 diff_1518000_1530000# gnd! 26.2fF
C2054 diff_1497600_1530000# gnd! 26.2fF
C2055 diff_1477200_1530000# gnd! 26.2fF
C2056 diff_1456800_1530000# gnd! 26.2fF
C2057 diff_1436400_1530000# gnd! 26.2fF
C2058 diff_1416000_1530000# gnd! 26.2fF
C2059 diff_1395600_1530000# gnd! 26.2fF
C2060 diff_1375200_1530000# gnd! 26.2fF
C2061 diff_1354800_1530000# gnd! 26.2fF
C2062 diff_1334400_1530000# gnd! 26.2fF
C2063 diff_1314000_1530000# gnd! 26.2fF
C2064 diff_1293600_1530000# gnd! 26.2fF
C2065 diff_1273200_1530000# gnd! 26.2fF
C2066 diff_1252800_1530000# gnd! 26.2fF
C2067 diff_1232400_1530000# gnd! 26.2fF
C2068 diff_1212000_1530000# gnd! 26.2fF
C2069 diff_1191600_1530000# gnd! 26.2fF
C2070 diff_1171200_1530000# gnd! 26.2fF
C2071 diff_1150800_1530000# gnd! 26.2fF
C2072 diff_1130400_1530000# gnd! 26.2fF
C2073 diff_1110000_1530000# gnd! 26.2fF
C2074 diff_1089600_1530000# gnd! 26.2fF
C2075 diff_1069200_1530000# gnd! 26.2fF
C2076 diff_1048800_1530000# gnd! 26.2fF
C2077 diff_1028400_1530000# gnd! 26.2fF
C2078 diff_1008000_1530000# gnd! 26.2fF
C2079 diff_1004400_1546800# gnd! 645.4fF
C2080 diff_2293200_1552800# gnd! 24.7fF
C2081 diff_2272800_1552800# gnd! 24.7fF
C2082 diff_2252400_1552800# gnd! 24.7fF
C2083 diff_2232000_1552800# gnd! 24.7fF
C2084 diff_2211600_1552800# gnd! 24.7fF
C2085 diff_2191200_1552800# gnd! 24.7fF
C2086 diff_2170800_1552800# gnd! 24.7fF
C2087 diff_2150400_1552800# gnd! 24.7fF
C2088 diff_2130000_1552800# gnd! 24.7fF
C2089 diff_2109600_1552800# gnd! 24.7fF
C2090 diff_2089200_1552800# gnd! 24.7fF
C2091 diff_2068800_1552800# gnd! 24.7fF
C2092 diff_2048400_1552800# gnd! 24.7fF
C2093 diff_2028000_1552800# gnd! 24.7fF
C2094 diff_2007600_1552800# gnd! 24.7fF
C2095 diff_1987200_1552800# gnd! 24.7fF
C2096 diff_1966800_1552800# gnd! 24.7fF
C2097 diff_1946400_1552800# gnd! 24.7fF
C2098 diff_1926000_1552800# gnd! 24.7fF
C2099 diff_1905600_1552800# gnd! 24.7fF
C2100 diff_1885200_1552800# gnd! 24.7fF
C2101 diff_1864800_1552800# gnd! 24.7fF
C2102 diff_1844400_1552800# gnd! 24.7fF
C2103 diff_1824000_1552800# gnd! 24.7fF
C2104 diff_1803600_1552800# gnd! 24.7fF
C2105 diff_1783200_1552800# gnd! 24.7fF
C2106 diff_1762800_1552800# gnd! 24.7fF
C2107 diff_1742400_1552800# gnd! 24.7fF
C2108 diff_1722000_1552800# gnd! 24.7fF
C2109 diff_1701600_1552800# gnd! 24.7fF
C2110 diff_1681200_1552800# gnd! 24.7fF
C2111 diff_1660800_1552800# gnd! 24.7fF
C2112 diff_1640400_1552800# gnd! 24.7fF
C2113 diff_1620000_1552800# gnd! 24.7fF
C2114 diff_1599600_1552800# gnd! 24.7fF
C2115 diff_1579200_1552800# gnd! 24.7fF
C2116 diff_1558800_1552800# gnd! 24.7fF
C2117 diff_1538400_1552800# gnd! 24.7fF
C2118 diff_1518000_1552800# gnd! 24.7fF
C2119 diff_1497600_1552800# gnd! 24.7fF
C2120 diff_1477200_1552800# gnd! 24.7fF
C2121 diff_1456800_1552800# gnd! 24.7fF
C2122 diff_1436400_1552800# gnd! 24.7fF
C2123 diff_1416000_1552800# gnd! 24.7fF
C2124 diff_1395600_1552800# gnd! 24.7fF
C2125 diff_1375200_1552800# gnd! 24.7fF
C2126 diff_1354800_1552800# gnd! 24.7fF
C2127 diff_1334400_1552800# gnd! 24.7fF
C2128 diff_1314000_1552800# gnd! 24.7fF
C2129 diff_1293600_1552800# gnd! 24.7fF
C2130 diff_1273200_1552800# gnd! 24.7fF
C2131 diff_1252800_1552800# gnd! 24.7fF
C2132 diff_1232400_1552800# gnd! 24.7fF
C2133 diff_1212000_1552800# gnd! 24.7fF
C2134 diff_1191600_1552800# gnd! 24.7fF
C2135 diff_1171200_1552800# gnd! 24.7fF
C2136 diff_1150800_1552800# gnd! 24.7fF
C2137 diff_1130400_1552800# gnd! 24.7fF
C2138 diff_1110000_1552800# gnd! 24.7fF
C2139 diff_1089600_1552800# gnd! 24.7fF
C2140 diff_1069200_1552800# gnd! 24.7fF
C2141 diff_1048800_1552800# gnd! 24.7fF
C2142 diff_1028400_1552800# gnd! 24.7fF
C2143 diff_1008000_1552800# gnd! 24.7fF
C2144 diff_562800_1448400# gnd! 324.8fF
C2145 diff_408000_1448400# gnd! 356.5fF
C2146 diff_1004400_1568400# gnd! 646.5fF
C2147 diff_2367600_1585200# gnd! 505.2fF
C2148 diff_2293200_1574400# gnd! 26.2fF
C2149 diff_2272800_1574400# gnd! 26.2fF
C2150 diff_2252400_1574400# gnd! 26.2fF
C2151 diff_2232000_1574400# gnd! 26.2fF
C2152 diff_2211600_1574400# gnd! 26.2fF
C2153 diff_2191200_1574400# gnd! 26.2fF
C2154 diff_2170800_1574400# gnd! 26.2fF
C2155 diff_2150400_1574400# gnd! 26.2fF
C2156 diff_2130000_1574400# gnd! 26.2fF
C2157 diff_2109600_1574400# gnd! 26.2fF
C2158 diff_2089200_1574400# gnd! 26.2fF
C2159 diff_2068800_1574400# gnd! 26.2fF
C2160 diff_2048400_1574400# gnd! 26.2fF
C2161 diff_2028000_1574400# gnd! 26.2fF
C2162 diff_2007600_1574400# gnd! 26.2fF
C2163 diff_1987200_1574400# gnd! 26.2fF
C2164 diff_1966800_1574400# gnd! 26.2fF
C2165 diff_1946400_1574400# gnd! 26.2fF
C2166 diff_1926000_1574400# gnd! 26.2fF
C2167 diff_1905600_1574400# gnd! 26.2fF
C2168 diff_1885200_1574400# gnd! 26.2fF
C2169 diff_1864800_1574400# gnd! 26.2fF
C2170 diff_1844400_1574400# gnd! 26.2fF
C2171 diff_1824000_1574400# gnd! 26.2fF
C2172 diff_1803600_1574400# gnd! 26.2fF
C2173 diff_1783200_1574400# gnd! 26.2fF
C2174 diff_1762800_1574400# gnd! 26.2fF
C2175 diff_1742400_1574400# gnd! 26.2fF
C2176 diff_1722000_1574400# gnd! 26.2fF
C2177 diff_1701600_1574400# gnd! 26.2fF
C2178 diff_1681200_1574400# gnd! 26.2fF
C2179 diff_1660800_1574400# gnd! 26.2fF
C2180 diff_1640400_1574400# gnd! 26.2fF
C2181 diff_1620000_1574400# gnd! 26.2fF
C2182 diff_1599600_1574400# gnd! 26.2fF
C2183 diff_1579200_1574400# gnd! 26.2fF
C2184 diff_1558800_1574400# gnd! 26.2fF
C2185 diff_1538400_1574400# gnd! 26.2fF
C2186 diff_1518000_1574400# gnd! 26.2fF
C2187 diff_1497600_1574400# gnd! 26.2fF
C2188 diff_1477200_1574400# gnd! 26.2fF
C2189 diff_1456800_1574400# gnd! 26.2fF
C2190 diff_1436400_1574400# gnd! 26.2fF
C2191 diff_1416000_1574400# gnd! 26.2fF
C2192 diff_1395600_1574400# gnd! 26.2fF
C2193 diff_1375200_1574400# gnd! 26.2fF
C2194 diff_1354800_1574400# gnd! 26.2fF
C2195 diff_1334400_1574400# gnd! 26.2fF
C2196 diff_1314000_1574400# gnd! 26.2fF
C2197 diff_1293600_1574400# gnd! 26.2fF
C2198 diff_1273200_1574400# gnd! 26.2fF
C2199 diff_1252800_1574400# gnd! 26.2fF
C2200 diff_1232400_1574400# gnd! 26.2fF
C2201 diff_1212000_1574400# gnd! 26.2fF
C2202 diff_1191600_1574400# gnd! 26.2fF
C2203 diff_1171200_1574400# gnd! 26.2fF
C2204 diff_1150800_1574400# gnd! 26.2fF
C2205 diff_1130400_1574400# gnd! 26.2fF
C2206 diff_1110000_1574400# gnd! 26.2fF
C2207 diff_1089600_1574400# gnd! 26.2fF
C2208 diff_1069200_1574400# gnd! 26.2fF
C2209 diff_1048800_1574400# gnd! 26.2fF
C2210 diff_1028400_1574400# gnd! 26.2fF
C2211 diff_1008000_1574400# gnd! 26.2fF
C2212 diff_1004400_1591200# gnd! 600.9fF
C2213 diff_2293200_1597200# gnd! 24.7fF
C2214 diff_2272800_1597200# gnd! 24.7fF
C2215 diff_2252400_1597200# gnd! 24.7fF
C2216 diff_2232000_1597200# gnd! 24.7fF
C2217 diff_2211600_1597200# gnd! 24.7fF
C2218 diff_2191200_1597200# gnd! 24.7fF
C2219 diff_2170800_1597200# gnd! 24.7fF
C2220 diff_2150400_1597200# gnd! 24.7fF
C2221 diff_2130000_1597200# gnd! 24.7fF
C2222 diff_2109600_1597200# gnd! 24.7fF
C2223 diff_2089200_1597200# gnd! 24.7fF
C2224 diff_2068800_1597200# gnd! 24.7fF
C2225 diff_2048400_1597200# gnd! 24.7fF
C2226 diff_2028000_1597200# gnd! 24.7fF
C2227 diff_2007600_1597200# gnd! 24.7fF
C2228 diff_1987200_1597200# gnd! 24.7fF
C2229 diff_1966800_1597200# gnd! 24.7fF
C2230 diff_1946400_1597200# gnd! 24.7fF
C2231 diff_1926000_1597200# gnd! 24.7fF
C2232 diff_1905600_1597200# gnd! 24.7fF
C2233 diff_1885200_1597200# gnd! 24.7fF
C2234 diff_1864800_1597200# gnd! 24.7fF
C2235 diff_1844400_1597200# gnd! 24.7fF
C2236 diff_1824000_1597200# gnd! 24.7fF
C2237 diff_1803600_1597200# gnd! 24.7fF
C2238 diff_1783200_1597200# gnd! 24.7fF
C2239 diff_1762800_1597200# gnd! 24.7fF
C2240 diff_1742400_1597200# gnd! 24.7fF
C2241 diff_1722000_1597200# gnd! 24.7fF
C2242 diff_1701600_1597200# gnd! 24.7fF
C2243 diff_1681200_1597200# gnd! 24.7fF
C2244 diff_1660800_1597200# gnd! 24.7fF
C2245 diff_1640400_1597200# gnd! 24.7fF
C2246 diff_1620000_1597200# gnd! 24.7fF
C2247 diff_1599600_1597200# gnd! 24.7fF
C2248 diff_1579200_1597200# gnd! 24.7fF
C2249 diff_1558800_1597200# gnd! 24.7fF
C2250 diff_1538400_1597200# gnd! 24.7fF
C2251 diff_1518000_1597200# gnd! 24.7fF
C2252 diff_1497600_1597200# gnd! 24.7fF
C2253 diff_1477200_1597200# gnd! 24.7fF
C2254 diff_1456800_1597200# gnd! 24.7fF
C2255 diff_1436400_1597200# gnd! 24.7fF
C2256 diff_1416000_1597200# gnd! 24.7fF
C2257 diff_1395600_1597200# gnd! 24.7fF
C2258 diff_1375200_1597200# gnd! 24.7fF
C2259 diff_1354800_1597200# gnd! 24.7fF
C2260 diff_1334400_1597200# gnd! 24.7fF
C2261 diff_1314000_1597200# gnd! 24.7fF
C2262 diff_1293600_1597200# gnd! 24.7fF
C2263 diff_1273200_1597200# gnd! 24.7fF
C2264 diff_1252800_1597200# gnd! 24.7fF
C2265 diff_1232400_1597200# gnd! 24.7fF
C2266 diff_1212000_1597200# gnd! 24.7fF
C2267 diff_1191600_1597200# gnd! 24.7fF
C2268 diff_1171200_1597200# gnd! 24.7fF
C2269 diff_1150800_1597200# gnd! 24.7fF
C2270 diff_1130400_1597200# gnd! 24.7fF
C2271 diff_1110000_1597200# gnd! 24.7fF
C2272 diff_1089600_1597200# gnd! 24.7fF
C2273 diff_1069200_1597200# gnd! 24.7fF
C2274 diff_1048800_1597200# gnd! 24.7fF
C2275 diff_1028400_1597200# gnd! 24.7fF
C2276 diff_1008000_1597200# gnd! 24.7fF
C2277 diff_1004400_1612800# gnd! 613.3fF
C2278 diff_2293200_1618800# gnd! 26.2fF
C2279 diff_2272800_1618800# gnd! 26.2fF
C2280 diff_2252400_1618800# gnd! 26.2fF
C2281 diff_2232000_1618800# gnd! 26.2fF
C2282 diff_2211600_1618800# gnd! 26.2fF
C2283 diff_2191200_1618800# gnd! 26.2fF
C2284 diff_2170800_1618800# gnd! 26.2fF
C2285 diff_2150400_1618800# gnd! 26.2fF
C2286 diff_2130000_1618800# gnd! 26.2fF
C2287 diff_2109600_1618800# gnd! 26.2fF
C2288 diff_2089200_1618800# gnd! 26.2fF
C2289 diff_2068800_1618800# gnd! 26.2fF
C2290 diff_2048400_1618800# gnd! 26.2fF
C2291 diff_2028000_1618800# gnd! 26.2fF
C2292 diff_2007600_1618800# gnd! 26.2fF
C2293 diff_1987200_1618800# gnd! 26.2fF
C2294 diff_1966800_1618800# gnd! 26.2fF
C2295 diff_1946400_1618800# gnd! 26.2fF
C2296 diff_1926000_1618800# gnd! 26.2fF
C2297 diff_1905600_1618800# gnd! 26.2fF
C2298 diff_1885200_1618800# gnd! 26.2fF
C2299 diff_1864800_1618800# gnd! 26.2fF
C2300 diff_1844400_1618800# gnd! 26.2fF
C2301 diff_1824000_1618800# gnd! 26.2fF
C2302 diff_1803600_1618800# gnd! 26.2fF
C2303 diff_1783200_1618800# gnd! 26.2fF
C2304 diff_1762800_1618800# gnd! 26.2fF
C2305 diff_1742400_1618800# gnd! 26.2fF
C2306 diff_1722000_1618800# gnd! 26.2fF
C2307 diff_1701600_1618800# gnd! 26.2fF
C2308 diff_1681200_1618800# gnd! 26.2fF
C2309 diff_1660800_1618800# gnd! 26.2fF
C2310 diff_1640400_1618800# gnd! 26.2fF
C2311 diff_1620000_1618800# gnd! 26.2fF
C2312 diff_1599600_1618800# gnd! 26.2fF
C2313 diff_1579200_1618800# gnd! 26.2fF
C2314 diff_1558800_1618800# gnd! 26.2fF
C2315 diff_1538400_1618800# gnd! 26.2fF
C2316 diff_1518000_1618800# gnd! 26.2fF
C2317 diff_1497600_1618800# gnd! 26.2fF
C2318 diff_1477200_1618800# gnd! 26.2fF
C2319 diff_1456800_1618800# gnd! 26.2fF
C2320 diff_1436400_1618800# gnd! 26.2fF
C2321 diff_1416000_1618800# gnd! 26.2fF
C2322 diff_1395600_1618800# gnd! 26.2fF
C2323 diff_1375200_1618800# gnd! 26.2fF
C2324 diff_1354800_1618800# gnd! 26.2fF
C2325 diff_1334400_1618800# gnd! 26.2fF
C2326 diff_1314000_1618800# gnd! 26.2fF
C2327 diff_1293600_1618800# gnd! 26.2fF
C2328 diff_1273200_1618800# gnd! 26.2fF
C2329 diff_1252800_1618800# gnd! 26.2fF
C2330 diff_1232400_1618800# gnd! 26.2fF
C2331 diff_1212000_1618800# gnd! 26.2fF
C2332 diff_1191600_1618800# gnd! 26.2fF
C2333 diff_1171200_1618800# gnd! 26.2fF
C2334 diff_1150800_1618800# gnd! 26.2fF
C2335 diff_1130400_1618800# gnd! 26.2fF
C2336 diff_1110000_1618800# gnd! 26.2fF
C2337 diff_1089600_1618800# gnd! 26.2fF
C2338 diff_1069200_1618800# gnd! 26.2fF
C2339 diff_1048800_1618800# gnd! 26.2fF
C2340 diff_1028400_1618800# gnd! 26.2fF
C2341 diff_1008000_1618800# gnd! 26.2fF
C2342 diff_1004400_1635600# gnd! 644.8fF
C2343 diff_2293200_1641600# gnd! 24.7fF
C2344 diff_2272800_1641600# gnd! 24.7fF
C2345 diff_2252400_1641600# gnd! 24.7fF
C2346 diff_2232000_1641600# gnd! 24.7fF
C2347 diff_2211600_1641600# gnd! 24.7fF
C2348 diff_2191200_1641600# gnd! 24.7fF
C2349 diff_2170800_1641600# gnd! 24.7fF
C2350 diff_2150400_1641600# gnd! 24.7fF
C2351 diff_2130000_1641600# gnd! 24.7fF
C2352 diff_2109600_1641600# gnd! 24.7fF
C2353 diff_2089200_1641600# gnd! 24.7fF
C2354 diff_2068800_1641600# gnd! 24.7fF
C2355 diff_2048400_1641600# gnd! 24.7fF
C2356 diff_2028000_1641600# gnd! 24.7fF
C2357 diff_2007600_1641600# gnd! 24.7fF
C2358 diff_1987200_1641600# gnd! 24.7fF
C2359 diff_1966800_1641600# gnd! 24.7fF
C2360 diff_1946400_1641600# gnd! 24.7fF
C2361 diff_1926000_1641600# gnd! 24.7fF
C2362 diff_1905600_1641600# gnd! 24.7fF
C2363 diff_1885200_1641600# gnd! 24.7fF
C2364 diff_1864800_1641600# gnd! 24.7fF
C2365 diff_1844400_1641600# gnd! 24.7fF
C2366 diff_1824000_1641600# gnd! 24.7fF
C2367 diff_1803600_1641600# gnd! 24.7fF
C2368 diff_1783200_1641600# gnd! 24.7fF
C2369 diff_1762800_1641600# gnd! 24.7fF
C2370 diff_1742400_1641600# gnd! 24.7fF
C2371 diff_1722000_1641600# gnd! 24.7fF
C2372 diff_1701600_1641600# gnd! 24.7fF
C2373 diff_1681200_1641600# gnd! 24.7fF
C2374 diff_1660800_1641600# gnd! 24.7fF
C2375 diff_1640400_1641600# gnd! 24.7fF
C2376 diff_1620000_1641600# gnd! 24.7fF
C2377 diff_1599600_1641600# gnd! 24.7fF
C2378 diff_1579200_1641600# gnd! 24.7fF
C2379 diff_1558800_1641600# gnd! 24.7fF
C2380 diff_1538400_1641600# gnd! 24.7fF
C2381 diff_1518000_1641600# gnd! 24.7fF
C2382 diff_1497600_1641600# gnd! 24.7fF
C2383 diff_1477200_1641600# gnd! 24.7fF
C2384 diff_1456800_1641600# gnd! 24.7fF
C2385 diff_1436400_1641600# gnd! 24.7fF
C2386 diff_1416000_1641600# gnd! 24.7fF
C2387 diff_1395600_1641600# gnd! 24.7fF
C2388 diff_1375200_1641600# gnd! 24.7fF
C2389 diff_1354800_1641600# gnd! 24.7fF
C2390 diff_1334400_1641600# gnd! 24.7fF
C2391 diff_1314000_1641600# gnd! 24.7fF
C2392 diff_1293600_1641600# gnd! 24.7fF
C2393 diff_1273200_1641600# gnd! 24.7fF
C2394 diff_1252800_1641600# gnd! 24.7fF
C2395 diff_1232400_1641600# gnd! 24.7fF
C2396 diff_1212000_1641600# gnd! 24.7fF
C2397 diff_1191600_1641600# gnd! 24.7fF
C2398 diff_1171200_1641600# gnd! 24.7fF
C2399 diff_1150800_1641600# gnd! 24.7fF
C2400 diff_1130400_1641600# gnd! 24.7fF
C2401 diff_1110000_1641600# gnd! 24.7fF
C2402 diff_1089600_1641600# gnd! 24.7fF
C2403 diff_1069200_1641600# gnd! 24.7fF
C2404 diff_1048800_1641600# gnd! 24.7fF
C2405 diff_1028400_1641600# gnd! 24.7fF
C2406 diff_1008000_1641600# gnd! 24.7fF
C2407 diff_886800_1546800# gnd! 88.0fF
C2408 diff_831600_1504800# gnd! 90.3fF
C2409 diff_820800_1365600# gnd! 612.4fF
C2410 diff_738000_1506000# gnd! 88.4fF
C2411 diff_673200_1506000# gnd! 97.3fF
C2412 diff_664800_1365600# gnd! 604.0fF
C2413 diff_189600_804000# gnd! 1761.5fF
C2414 diff_583200_1506000# gnd! 94.7fF
C2415 diff_520800_1503600# gnd! 89.9fF
C2416 diff_510000_1366800# gnd! 615.1fF
C2417 diff_428400_1507200# gnd! 90.8fF
C2418 diff_366000_1504800# gnd! 94.2fF
C2419 diff_1004400_1657200# gnd! 642.3fF
C2420 diff_2505600_919200# gnd! 629.7fF
C2421 diff_2488800_853200# gnd! 640.2fF
C2422 diff_2367600_1674000# gnd! 499.8fF
C2423 diff_2293200_1663200# gnd! 26.2fF
C2424 diff_2272800_1663200# gnd! 26.2fF
C2425 diff_2252400_1663200# gnd! 26.2fF
C2426 diff_2232000_1663200# gnd! 26.2fF
C2427 diff_2211600_1663200# gnd! 26.2fF
C2428 diff_2191200_1663200# gnd! 26.2fF
C2429 diff_2170800_1663200# gnd! 26.2fF
C2430 diff_2150400_1663200# gnd! 26.2fF
C2431 diff_2130000_1663200# gnd! 26.2fF
C2432 diff_2109600_1663200# gnd! 26.2fF
C2433 diff_2089200_1663200# gnd! 26.2fF
C2434 diff_2068800_1663200# gnd! 26.2fF
C2435 diff_2048400_1663200# gnd! 26.2fF
C2436 diff_2028000_1663200# gnd! 26.2fF
C2437 diff_2007600_1663200# gnd! 26.2fF
C2438 diff_1987200_1663200# gnd! 26.2fF
C2439 diff_1966800_1663200# gnd! 26.2fF
C2440 diff_1946400_1663200# gnd! 26.2fF
C2441 diff_1926000_1663200# gnd! 26.2fF
C2442 diff_1905600_1663200# gnd! 26.2fF
C2443 diff_1885200_1663200# gnd! 26.2fF
C2444 diff_1864800_1663200# gnd! 26.2fF
C2445 diff_1844400_1663200# gnd! 26.2fF
C2446 diff_1824000_1663200# gnd! 26.2fF
C2447 diff_1803600_1663200# gnd! 26.2fF
C2448 diff_1783200_1663200# gnd! 26.2fF
C2449 diff_1762800_1663200# gnd! 26.2fF
C2450 diff_1742400_1663200# gnd! 26.2fF
C2451 diff_1722000_1663200# gnd! 26.2fF
C2452 diff_1701600_1663200# gnd! 26.2fF
C2453 diff_1681200_1663200# gnd! 26.2fF
C2454 diff_1660800_1663200# gnd! 26.2fF
C2455 diff_1640400_1663200# gnd! 26.2fF
C2456 diff_1620000_1663200# gnd! 26.2fF
C2457 diff_1599600_1663200# gnd! 26.2fF
C2458 diff_1579200_1663200# gnd! 26.2fF
C2459 diff_1558800_1663200# gnd! 26.2fF
C2460 diff_1538400_1663200# gnd! 26.2fF
C2461 diff_1518000_1663200# gnd! 26.2fF
C2462 diff_1497600_1663200# gnd! 26.2fF
C2463 diff_1477200_1663200# gnd! 26.2fF
C2464 diff_1456800_1663200# gnd! 26.2fF
C2465 diff_1436400_1663200# gnd! 26.2fF
C2466 diff_1416000_1663200# gnd! 26.2fF
C2467 diff_1395600_1663200# gnd! 26.2fF
C2468 diff_1375200_1663200# gnd! 26.2fF
C2469 diff_1354800_1663200# gnd! 26.2fF
C2470 diff_1334400_1663200# gnd! 26.2fF
C2471 diff_1314000_1663200# gnd! 26.2fF
C2472 diff_1293600_1663200# gnd! 26.2fF
C2473 diff_1273200_1663200# gnd! 26.2fF
C2474 diff_1252800_1663200# gnd! 26.2fF
C2475 diff_1232400_1663200# gnd! 26.2fF
C2476 diff_1212000_1663200# gnd! 26.2fF
C2477 diff_1191600_1663200# gnd! 26.2fF
C2478 diff_1171200_1663200# gnd! 26.2fF
C2479 diff_1150800_1663200# gnd! 26.2fF
C2480 diff_1130400_1663200# gnd! 26.2fF
C2481 diff_1110000_1663200# gnd! 26.2fF
C2482 diff_1089600_1663200# gnd! 26.2fF
C2483 diff_1069200_1663200# gnd! 26.2fF
C2484 diff_1048800_1663200# gnd! 26.2fF
C2485 diff_1028400_1663200# gnd! 26.2fF
C2486 diff_1008000_1663200# gnd! 26.2fF
C2487 diff_1004400_1680000# gnd! 607.3fF
C2488 diff_2431200_979200# gnd! 701.5fF
C2489 diff_2413200_996000# gnd! 740.5fF
C2490 diff_2384400_427200# gnd! 721.5fF
C2491 diff_2361600_427200# gnd! 533.5fF
C2492 diff_1008000_1686000# gnd! 1615.4fF
C2493 diff_1657200_1702800# gnd! 1099.3fF
C2494 diff_2664000_1686000# gnd! 153.5fF
C2495 diff_2649600_1428000# gnd! 296.5fF
C2496 diff_2613600_1719600# gnd! 236.2fF
C2497 diff_2437200_1698000# gnd! 1171.5fF
C2498 diff_1003200_1702800# gnd! 784.0fF
C2499 diff_2433600_1742400# gnd! 897.8fF
C2500 diff_2751600_1686000# gnd! 129.0fF
C2501 diff_2802000_1732800# gnd! 101.5fF
C2502 diff_804000_1662000# gnd! 965.5fF
C2503 diff_649200_1662000# gnd! 967.9fF
C2504 Vdd gnd! 17173.4fF
C2505 diff_355200_1366800# gnd! 615.1fF
C2506 diff_494400_1662000# gnd! 978.3fF
C2507 diff_338400_1662000# gnd! 977.5fF
C2508 d0 gnd! 2086.6fF
C2509 d1 gnd! 1942.9fF
C2510 d3 gnd! 3676.4fF
C2511 sync gnd! 2261.0fF
C2512 d2 gnd! 2260.5fF
C2513 clk1 gnd! 2051.4fF
C2514 clk2 gnd! 3136.5fF
