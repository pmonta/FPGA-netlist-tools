* SPICE3 netlist

M0 pcl0 dpc39_PCLPCL pclp0 GND efet
M1 pcl3 dpc39_PCLPCL pclp3 GND efet
M2 pcl4 dpc39_PCLPCL pclp4 GND efet
M3 pcl7 dpc39_PCLPCL pclp7 GND efet
M4 pcl6 dpc39_PCLPCL pclp6 GND efet
M5 pcl1 dpc39_PCLPCL pclp1 GND efet
M6 DA_C01 n_A_B_0 GND GND efet
M7 n_1347 n_782 GND GND efet
M8 op_SRS n_366 GND GND efet
M9 pcl5 dpc39_PCLPCL pclp5 GND efet
M10 op_T__dex notir1 GND GND efet
M11 n_1347 n_979 GND GND efet
M12 n_1103 op_T2_idx_x_xy n_1106 GND efet
M13 GND pd2 pd2_clearIR GND efet
M14 GND op_T5_brk n_1464 GND efet
M15 GND n_790 op_rmw GND efet
M16 n_911 n_1343 GND GND efet
M17 GND x_op_T0_txa n_1106 GND efet
M18 GND n_1054 n_70 GND efet
M19 idb0 dpc37_PCLDB pclp0 GND efet
M20 n_320 sb1 GND GND efet
M21 n_253 pipeUNK42 GND GND efet
M22 dpc14_SRS n_1552 GND GND efet
M23 GND n_71 dpc7_SS GND efet
M24 x7 dpc3_SBX sb7 GND efet
M25 GND n_1629 dasb5 GND efet
M26 GND nABL2 abl2 GND efet
M27 Vdd n_520 db2 GND efet
M28 Vdd n_520 db2 GND efet
M29 n_1719 a5 GND GND efet
M30 n_1717 op_T3_ind_y GND GND efet
M31 n_524 ADL_ABL nABL6 GND efet
M32 n_886 cclk GND GND efet
M33 n_738 ADL_ABL nABL4 GND efet
M34 n_577 ADL_ABL nABL7 GND efet
M35 n_1094 adl5 GND GND efet
M36 n_463 ADL_ABL nABL5 GND efet
M37 n_261 x_op_T4_ind_y GND GND efet
M38 GND nNMIG n_1712 GND efet
M39 n_380 fetch clearIR GND efet
M40 n_726 x_op_T4_ind_y GND GND efet
M41 Vdd dor5 n_373 GND efet
M42 Vdd n_1296 ab11 GND efet
M43 n_711 n_761 n_739 GND efet
M44 n_914 n_715 GND GND efet
M45 n_426 n_715 GND GND efet
M46 n_952 n_272 GND GND efet
M47 n_1366 pipeT3out GND GND efet
M48 GND nVEC n_70 GND efet
M49 GND n_646 n_812 GND efet
M50 GND n_1312 nNMIG GND efet
M51 n_658 cclk y4 GND efet
M52 n_1056 n_761 GND GND efet
M53 ab15 n_659 GND GND efet
M54 sb0 dpc24_ACSB n_146 GND efet
M55 ab15 n_659 GND GND efet
M56 GND n_659 ab15 GND efet
M57 sb3 dpc24_ACSB n_1654 GND efet
M58 sb4 dpc24_ACSB n_1344 GND efet
M59 sb1 dpc24_ACSB n_929 GND efet
M60 n_1618 dpc24_ACSB sb2 GND efet
M61 sb5 dpc24_ACSB n_831 GND efet
M62 n_326 dpc24_ACSB sb6 GND efet
M63 Vdd n_772 dpc17_SUMS GND efet
M64 GND s5 n_496 GND efet
M65 pclp2 npclp2 GND GND efet
M66 dpc23_SBAC cclk GND GND efet
M67 n_625 n_459 GND GND efet
M68 n_830 n_43 GND GND efet
M69 irq GND GND GND efet
M70 n_566 n_755 n_580 GND efet
M71 n_520 dor2 Vdd GND efet
M72 GND n_732 n_17 GND efet
M73 GND n_743 n_1547 GND efet
M74 GND notx2 n_1694 GND efet
M75 GND n_743 n_875 GND efet
M76 n_545 n_743 n_609 GND efet
M77 n_1194 p3 GND GND efet
M78 n_988 nA_B3 GND GND efet
M79 n_620 n_1293 GND GND efet
M80 nC12 n_936 GND GND efet
M81 n_321 n_398 GND GND efet
M82 n_692 n_43 GND GND efet
M83 op_T3_branch irline3 GND GND efet
M84 GND irline3 op_brk_rti GND efet
M85 op_T0_brk_rti irline3 GND GND efet
M86 op_T0_jmp irline3 GND GND efet
M87 op_T2_branch irline3 GND GND efet
M88 op_T5_rts irline3 GND GND efet
M89 GND irline3 op_T2_brk GND efet
M90 GND irline3 op_T3_jsr GND efet
M91 GND irline3 op_jsr GND efet
M92 GND irline3 x_op_jmp GND efet
M93 GND n_1033 dpc21_ADDADL GND efet
M94 n_457 idb3 GND GND efet
M95 GND n_1274 n_1069 GND efet
M96 n_11 cclk n_55 GND efet
M97 n_306 dpc22_nDSA GND GND efet
M98 GND n_882 NMIL GND efet
M99 PD_1xx000x0 pd0_clearIR GND GND efet
M100 GND pd0_clearIR PD_xxxx10x0 GND efet
M101 n_269 n_1038 GND GND efet
M102 n_1365 n_862 GND GND efet
M103 GND op_T0_txa n_1455 GND efet
M104 GND n_526 npclp0 GND efet
M105 GND n_1392 n_284 GND efet
M106 x1 cclk n_1709 GND efet
M107 GND abl1 n_842 GND efet
M108 n_66 abl1 GND GND efet
M109 nNMIP n_1392 n_346 GND efet
M110 n_1705 n_467 GND GND efet
M111 n_562 cp1 n_645 GND efet
M112 GND n_0_ADL1 adl1 GND efet
M113 adh4 dpc27_SBADH sb4 GND efet
M114 GND notRdy0 notRnWprepad GND efet
M115 GND n_869 ab13 GND efet
M116 ab13 n_869 GND GND efet
M117 adl0 dpc10_ADLADD alub0 GND efet
M118 GND C1x5Reset n_1054 GND efet
M119 n_424 n_198 GND GND efet
M120 n_1717 n_335 n_1604 GND efet
M121 GND n_869 ab13 GND efet
M122 ab13 n_869 GND GND efet
M123 n_694 dpc4_SSB sb1 GND efet
M124 GND n_869 ab13 GND efet
M125 pclp5 dpc38_PCLADL adl5 GND efet
M126 adl6 dpc38_PCLADL pclp6 GND efet
M127 n_1694 dpc2_XSB sb2 GND efet
M128 n_242 dpc2_XSB sb3 GND efet
M129 n_1159 n_1580 GND GND efet
M130 n_845 n_1573 n_1550 GND efet
M131 GND n_236 n_506 GND efet
M132 n_1656 n_1580 GND GND efet
M133 n_1724 dpc2_XSB sb6 GND efet
M134 GND n_1256 dpc15_ANDS GND efet
M135 n_959 short_circuit_branch_add GND GND efet
M136 n_578 dpc2_XSB sb5 GND efet
M137 GND notidl3 idl3 GND efet
M138 GND n_646 n_1172 GND efet
M139 GND notidl3 idl3 GND efet
M140 GND notidl3 idl3 GND efet
M141 GND idb2 n_1573 GND efet
M142 GND notalu5 alu5 GND efet
M143 Vdd n_625 dpc3_SBX GND efet
M144 n_319 DA_C01 n_1707 GND efet
M145 n_218 n_368 GND GND efet
M146 DBZ idb6 GND GND efet
M147 clk0 GND GND GND efet
M148 GND n_1120 n_137 GND efet
M149 sb0 dpc6_SBS s0 GND efet
M150 n_1694 cclk x2 GND efet
M151 idb3 cclk Vdd GND efet
M152 GND clock2 op_T__cpx_cpy_imm_zp GND efet
M153 GND npchp2 pchp2 GND efet
M154 GND RnWstretched n_37 GND efet
M155 nA_B3 alub3 n_313 GND efet
M156 GND op_T0_jsr n_1464 GND efet
M157 n_279 n_954 GND GND efet
M158 Vdd n_288 n_794 GND efet
M159 n_826 abh0 Vdd GND efet
M160 n_625 n_43 GND GND efet
M161 GND s3 n_34 GND efet
M162 GND npchp6 pchp6 GND efet
M163 GND adl4 n_1519 GND efet
M164 n_262 cp1 n_1447 GND efet
M165 n_717 pipephi2Reset0x GND GND efet
M166 GND notx5 n_578 GND efet
M167 GND n_906 dpc19_ADDSB7 GND efet
M168 n_1341 cclk n_695 GND efet
M169 GND nots6 n_618 GND efet
M170 n_1260 n_598 GND GND efet
M171 noty5 y5 GND GND efet
M172 sb7 dpc11_SBADD alua7 GND efet
M173 GND pipeUNK08 n_954 GND efet
M174 GND n_1049 n_507 GND efet
M175 GND cp1 n_839 GND efet
M176 GND cp1 n_43 GND efet
M177 n_1095 cp1 idl4 GND efet
M178 n_548 cclk nots7 GND efet
M179 sb5 cclk Vdd GND efet
M180 Vdd n_154 dpc20_ADDSB06 GND efet
M181 GND n_154 n_75 GND efet
M182 n_789 idb7 GND GND efet
M183 n_397 op_T0_lda GND GND efet
M184 GND idb0 n_624 GND efet
M185 n_AxB_3 AxB3 GND GND efet
M186 GND x5 notx5 GND efet
M187 n_1590 cp1 n_1083 GND efet
M188 n_1455 op_T0_lda GND GND efet
M189 n_1424 cp1 idl2 GND efet
M190 n_795 cclk n_360 GND efet
M191 dasb6 n_739 n_1554 GND efet
M192 rw n_1696 GND GND efet
M193 rw n_1696 GND GND efet
M194 naluresult2 cclk notalu2 GND efet
M195 GND op_rol_ror n_1000 GND efet
M196 n_753 n_1257 GND GND efet
M197 n_711 n_1257 GND GND efet
M198 GND n_1257 n_569 GND efet
M199 n_152 n_630 GND GND efet
M200 noty0 y0 GND GND efet
M201 GND op_T3_abs_idx n_1107 GND efet
M202 op_T2_jsr ir3 GND GND efet
M203 GND op_T2_mem_zp n_347 GND efet
M204 Vdd abh2 n_1545 GND efet
M205 GND abh2 n_1034 GND efet
M206 n_1584 n_8 n_345 GND efet
M207 GND dor2 n_37 GND efet
M208 n_718 cclk notidl0 GND efet
M209 n_165 A_B5 GND GND efet
M210 GND n_1417 clk1out GND efet
M211 clk1out n_1417 GND GND efet
M212 GND n_1417 clk1out GND efet
M213 clk1out n_1417 GND GND efet
M214 n_1130 n_1109 GND GND efet
M215 clk1out n_1417 GND GND efet
M216 sb1 dpc27_SBADH adh1 GND efet
M217 GND dpc12_0ADD alua2 GND efet
M218 n_1275 cp1 n_1581 GND efet
M219 D1x1 cp1 n_1472 GND efet
M220 D1x1 INTG GND GND efet
M221 GND op_T2_pha n_1037 GND efet
M222 GND n_445 n_417 GND efet
M223 n_127 cp1 GND GND efet
M224 sync n_445 GND GND efet
M225 GND n_445 sync GND efet
M226 sync n_445 GND GND efet
M227 GND n_445 sync GND efet
M228 GND n_445 sync GND efet
M229 abh2 nABH2 GND GND efet
M230 n_1215 brk_done GND GND efet
M231 GND AxB5 n_547 GND efet
M232 op_T3_branch ir2 GND GND efet
M233 op_brk_rti ir2 GND GND efet
M234 op_T2_branch ir2 GND GND efet
M235 op_T2_ind ir2 GND GND efet
M236 op_T2_brk ir2 GND GND efet
M237 op_T3_jsr ir2 GND GND efet
M238 op_T5_ind_x ir2 GND GND efet
M239 x_op_T4_ind_y ir2 GND GND efet
M240 op_T5_rts ir2 GND GND efet
M241 op_T0_brk_rti ir2 GND GND efet
M242 n_1391 cclk pipeUNK15 GND efet
M243 GND n_531 n_1255 GND efet
M244 Vdd n_531 dpc13_ORS GND efet
M245 Vdd dor7 n_298 GND efet
M246 nABH4 cclk n_999 GND efet
M247 n_1298 ADH_ABH nABH1 GND efet
M248 n_1106 cclk n_1404 GND efet
M249 GND notidl5 idl5 GND efet
M250 GND notidl5 idl5 GND efet
M251 GND notidl5 idl5 GND efet
M252 n_368 op_T2_php_pha GND GND efet
M253 n_556 a4 GND GND efet
M254 n_1194 cclk pipeUNK04 GND efet
M255 n_470 n_646 GND GND efet
M256 db0 GND GND GND efet
M257 pipeUNK30 cclk n_385 GND efet
M258 GND VEC1 n_912 GND efet
M259 GND n_781 n_160 GND efet
M260 n_291 n_1121 GND GND efet
M261 GND op_T2_php_pha nWR GND efet
M262 GND pd5_clearIR n_928 GND efet
M263 n_891 n_284 NMIP GND efet
M264 n_1070 pch1 GND GND efet
M265 op_T3_ind_y notir4 GND GND efet
M266 op_T2_abs_y notir4 GND GND efet
M267 x_op_T0_tya notir4 GND GND efet
M268 op_T2_idx_x_xy notir4 GND GND efet
M269 op_T0_txs notir4 GND GND efet
M270 op_T0_tsx notir4 GND GND efet
M271 op_T4_ind_y notir4 GND GND efet
M272 n_1558 n_16 n_428 GND efet
M273 GND op_T4 n_256 GND efet
M274 GND GND so GND efet
M275 nop_set_C op_asl_rol n_591 GND efet
M276 n_AxB_5 dpc16_EORS naluresult5 GND efet
M277 n_AxB_4 dpc16_EORS naluresult4 GND efet
M278 naluresult7 dpc16_EORS n_AxB_7 GND efet
M279 n_AxB_6 dpc16_EORS naluresult6 GND efet
M280 GND clock2 op_T__dex GND efet
M281 n_1053 Pout3 GND GND efet
M282 ab11 n_359 GND GND efet
M283 GND n_359 ab11 GND efet
M284 ab11 n_359 GND GND efet
M285 GND n_359 ab11 GND efet
M286 n_1107 op_T2_ind_y GND GND efet
M287 GND ir4 notir4 GND efet
M288 n_811 n_838 GND GND efet
M289 GND clearIR pd6_clearIR GND efet
M290 pd2_clearIR clearIR GND GND efet
M291 GND n_1184 n_410 GND efet
M292 n_474 n_1184 n_766 GND efet
M293 short_circuit_branch_add n_771 n_465 GND efet
M294 GND n_771 n_1446 GND efet
M295 GND n_745 n_241 GND efet
M296 GND op_T__cmp nop_set_C GND efet
M297 op_T__cpx_cpy_abs notir2 GND GND efet
M298 GND notir2 op_T3_mem_abs GND efet
M299 op_T2_jmp_abs notir2 GND GND efet
M300 op_T__bit notir2 GND GND efet
M301 op_T3_mem_zp_idx notir2 GND GND efet
M302 x_op_T0_bit notir2 GND GND efet
M303 op_T2_zp_zp_idx notir2 GND GND efet
M304 op_T0_jmp notir2 GND GND efet
M305 x_op_jmp notir2 GND GND efet
M306 op_T4_jmp notir2 GND GND efet
M307 n_1388 AxB1 GND GND efet
M308 n_1517 n_853 GND GND efet
M309 n_1584 n_876 GND GND efet
M310 ab7 n_322 Vdd GND efet
M311 ab7 n_322 Vdd GND efet
M312 op_T5_brk ir4 GND GND efet
M313 op_T0_php_pha ir4 GND GND efet
M314 op_T0_tay_ldy_not_idx ir4 GND GND efet
M315 op_T0_jsr ir4 GND GND efet
M316 n_676 cclk nABH1 GND efet
M317 op_T5_rti ir4 GND GND efet
M318 op_jmp ir4 GND GND efet
M319 op_T4_rts ir4 GND GND efet
M320 n_239 n_595 GND GND efet
M321 op_T3_plp_pla ir4 GND GND efet
M322 GND n_339 n_543 GND efet
M323 Vdd n_91 dpc15_ANDS GND efet
M324 n_442 cclk n_509 GND efet
M325 GND n_126 npchp1 GND efet
M326 GND notir7 op_sty_cpy_mem GND efet
M327 GND noty0 n_564 GND efet
M328 n_1368 cp1 n_1149 GND efet
M329 GND n_402 n_834 GND efet
M330 GND n_1369 n_1462 GND efet
M331 n_1389 dpc4_SSB sb2 GND efet
M332 nABH7 ADH_ABH n_514 GND efet
M333 n_1358 n_917 GND GND efet
M334 GND npclp7 pclp7 GND efet
M335 n_692 n_460 GND GND efet
M336 n_998 dpc4_SSB sb3 GND efet
M337 n_1179 cclk n_393 GND efet
M338 short_circuit_branch_add cp1 n_1570 GND efet
M339 GND DBZ nDBZ GND efet
M340 op_T0_clc_sec notir3 GND GND efet
M341 op_T0_plp notir3 GND GND efet
M342 op_implied notir3 GND GND efet
M343 op_clv notir3 GND GND efet
M344 op_T4_jmp notir3 GND GND efet
M345 op_T2_jmp_abs notir3 GND GND efet
M346 x_op_T3_plp_pla notir3 GND GND efet
M347 op_T0_cli_sei notir3 GND GND efet
M348 op_T__cpx_cpy_abs notir3 GND GND efet
M349 op_T4_mem_abs_idx notir3 GND GND efet
M350 GND clock1 op_T0_tax GND efet
M351 n_1631 n_1184 n_903 GND efet
M352 n_924 A_B3 GND GND efet
M353 GND op_T0_brk_rti n_256 GND efet
M354 GND n_1105 cp1 GND efet
M355 GND n_1105 cp1 GND efet
M356 n_643 dor3 GND GND efet
M357 GND op_T4_abs_idx n_595 GND efet
M358 pipenVEC cclk nVEC GND efet
M359 n_1613 dor3 GND GND efet
M360 GND n_1105 cp1 GND efet
M361 cp1 n_1105 GND GND efet
M362 adl3 dpc5_SADL n_998 GND efet
M363 adl4 dpc5_SADL n_3 GND efet
M364 adl5 dpc5_SADL n_280 GND efet
M365 n_503 notir5 GND GND efet
M366 n_721 dpc5_SADL adl7 GND efet
M367 n_553 n_1662 GND GND efet
M368 adl2 dpc5_SADL n_1389 GND efet
M369 GND nABL1 abl1 GND efet
M370 pclp0 npclp0 GND GND efet
M371 n_182 op_T5_rts GND GND efet
M372 n_1183 cp1 n_1605 GND efet
M373 n_1181 n_1595 n_793 GND efet
M374 n_261 cclk pipeUNK36 GND efet
M375 n_959 cp1 n_323 GND efet
M376 n_442 n_182 GND GND efet
M377 Vdd dor1 n_798 GND efet
M378 n_335 n_347 GND GND efet
M379 n_1215 n_238 GND GND efet
M380 n_1578 pipenVEC GND GND efet
M381 GND n_785 n_267 GND efet
M382 ab11 n_1296 Vdd GND efet
M383 GND n_1159 dasb2 GND efet
M384 RnWstretched n_1028 Vdd GND efet
M385 GND n_676 ab9 GND efet
M386 GND n_676 ab9 GND efet
M387 GND n_748 AxB7 GND efet
M388 GND n_676 ab9 GND efet
M389 n_1103 n_1244 GND GND efet
M390 n_620 n_1433 GND GND efet
M391 pipeUNK29 cclk n_169 GND efet
M392 n_1714 pipeUNK26 GND GND efet
M393 n_1687 cp1 notdor0 GND efet
M394 n_299 cp1 n_1625 GND efet
M395 ir3 n_1620 GND GND efet
M396 pipeUNK11 cclk n_862 GND efet
M397 n_1498 n_163 GND GND efet
M398 n_903 n_163 GND GND efet
M399 GND pch6 n_278 GND efet
M400 GND notRdy0 n_372 GND efet
M401 GND n_221 n_251 GND efet
M402 n_171 abl7 GND GND efet
M403 GND n_551 n_8 GND efet
M404 Vdd abl7 n_322 GND efet
M405 nmi GND GND GND efet
M406 n_1620 cclk notir3 GND efet
M407 dpc10_ADLADD n_491 GND GND efet
M408 n_1275 pipeBRtaken GND GND efet
M409 dor2 notdor2 GND GND efet
M410 ab9 n_1140 Vdd GND efet
M411 n_656 n_779 n_1594 GND efet
M412 op_implied x_op_push_pull GND GND efet
M413 n_862 cclk pipeT_SYNC GND efet
M414 n_213 cclk notidl1 GND efet
M415 n_1685 n_1166 GND GND efet
M416 n_789 cp1 notdor7 GND efet
M417 GND n_1660 n_855 GND efet
M418 n_1568 n_1166 GND GND efet
M419 GND nVEC n_1712 GND efet
M420 n_1100 n_1660 Vdd GND efet
M421 notRdy0 cp1 n_902 GND efet
M422 notir2 ir2 GND GND efet
M423 n_AxB1__C01 nC01 GND GND efet
M424 GND RnWstretched n_7 GND efet
M425 n_771 n_1110 GND GND efet
M426 n_AxBxC_1 nC01 n_1388 GND efet
M427 n_920 pipeUNK27 GND GND efet
M428 n_AxBxC_4 _AxB_4_nC34 GND GND efet
M429 GND n_810 n_207 GND efet
M430 n_AxBxC_0 _AxB_0_nC0in GND GND efet
M431 n_202 nnT2BR GND GND efet
M432 Vdd n_963 ab14 GND efet
M433 n_1563 op_T0_acc GND GND efet
M434 Vdd abh3 n_1296 GND efet
M435 n_844 op_T__dex GND GND efet
M436 GND db4 n_1075 GND efet
M437 GND dpc34_PCLC n_1007 GND efet
M438 notx0 x0 GND GND efet
M439 GND n_318 n_1293 GND efet
M440 pch7 dpc31_PCHPCH pchp7 GND efet
M441 pch4 dpc31_PCHPCH pchp4 GND efet
M442 n_176 n_236 GND GND efet
M443 pch6 dpc31_PCHPCH pchp6 GND efet
M444 pch5 dpc31_PCHPCH pchp5 GND efet
M445 pch2 dpc31_PCHPCH pchp2 GND efet
M446 GND db2 n_1199 GND efet
M447 n_524 cp1 n_1548 GND efet
M448 nABH6 ADH_ABH n_1514 GND efet
M449 GND GND clk0 GND efet
M450 ab8 n_826 Vdd GND efet
M451 GND db1 n_1319 GND efet
M452 GND notalucout alucout GND efet
M453 GND GND cclk GND efet
M454 GND pipeVectorA0 n_0_ADL0 GND efet
M455 Vdd n_1608 ab13 GND efet
M456 GND notir5 op_T0_jsr GND efet
M457 GND notir5 op_ror GND efet
M458 GND notir5 op_T3_plp_pla GND efet
M459 GND notir5 op_T0_tsx GND efet
M460 GND notir5 op_T__inx GND efet
M461 GND notir5 op_T0_tay_ldy_not_idx GND efet
M462 GND notir5 op_T0_ldy_mem GND efet
M463 GND notir5 op_inc_nop GND efet
M464 GND notir5 op_plp_pla GND efet
M465 op_T0_cmp notir6 GND GND efet
M466 op_T0_sbc notir6 GND GND efet
M467 op_rti_rts notir6 GND GND efet
M468 GND notir6 op_T0_cpx_cpy_inx_iny GND efet
M469 op_T4_rti notir6 GND GND efet
M470 op_inc_nop notir6 GND GND efet
M471 op_T0_eor notir6 GND GND efet
M472 GND notir6 op_jmp GND efet
M473 GND notir6 op_T0_adc_sbc GND efet
M474 GND notir6 op_T3_jmp GND efet
M475 n_1499 n_1450 GND GND efet
M476 ir5 n_1609 GND GND efet
M477 Vdd n_1152 ab2 GND efet
M478 Vdd n_1152 ab2 GND efet
M479 n_1081 n_1560 GND GND efet
M480 ab2 n_1152 Vdd GND efet
M481 n_299 n_1245 n_1723 GND efet
M482 GND alu1 nDA_ADD1 GND efet
M483 ab2 n_1152 Vdd GND efet
M484 ab2 n_1152 Vdd GND efet
M485 GND n_994 ab10 GND efet
M486 GND n_994 ab10 GND efet
M487 ab10 n_994 GND GND efet
M488 GND n_994 ab10 GND efet
M489 GND n_781 n_1170 GND efet
M490 n_1417 n_670 Vdd GND efet
M491 GND n_994 ab10 GND efet
M492 ab10 n_994 GND GND efet
M493 ab10 n_994 GND GND efet
M494 GND noty6 n_518 GND efet
M495 Vdd n_1596 dpc27_SBADH GND efet
M496 n_1271 n_1596 GND GND efet
M497 n_182 cclk n_265 GND efet
M498 GND notalucin n_1354 GND efet
M499 n_368 op_T5_rti_rts GND GND efet
M500 n_1635 n_966 GND GND efet
M501 GND n_1214 fetch GND efet
M502 n_770 n_559 GND GND efet
M503 Vdd n_966 dpc29_0ADH17 GND efet
M504 GND n_783 n_1158 GND efet
M505 n_835 n_311 GND GND efet
M506 n_856 n_311 GND GND efet
M507 n_490 cclk notidl4 GND efet
M508 n_1673 cclk op_T__bit GND efet
M509 n_513 cclk pipeUNK06 GND efet
M510 idb2 H1x1 Pout2 GND efet
M511 GND n_610 n_582 GND efet
M512 GND dor4 n_1463 GND efet
M513 GND dor4 n_147 GND efet
M514 op_T0_tsx ir2 GND GND efet
M515 op_T__iny_dey ir2 GND GND efet
M516 op_T__dex ir2 GND GND efet
M517 op_T__inx ir2 GND GND efet
M518 op_T0_dex ir2 GND GND efet
M519 op_T0_txs ir2 GND GND efet
M520 op_T2_ind_x ir2 GND GND efet
M521 x_op_T0_txa ir2 GND GND efet
M522 op_T0_iny_dey ir2 GND GND efet
M523 x_op_T0_tya ir2 GND GND efet
M524 n_1251 dpc0_YSB sb7 GND efet
M525 n_1290 n_1126 GND GND efet
M526 n_1556 nDA_ADD2 n_986 GND efet
M527 n_867 nDA_ADD2 GND GND efet
M528 n_1649 op_T2_abs GND GND efet
M529 GND n_43 n_1541 GND efet
M530 GND n_1529 n_91 GND efet
M531 GND op_T0_tax n_11 GND efet
M532 n_854 cp1 n_1395 GND efet
M533 GND n_1070 n_1538 GND efet
M534 dpc35_PCHC n_1070 GND GND efet
M535 n_1681 n_440 n_905 GND efet
M536 idb6 cclk Vdd GND efet
M537 n_1412 n_1455 GND GND efet
M538 n_726 op_T5_rts GND GND efet
M539 n_468 cp1 n_18 GND efet
M540 n_1039 cp1 n_24 GND efet
M541 n_1649 n_389 GND GND efet
M542 n_A_B_4 dpc13_ORS naluresult4 GND efet
M543 n_993 cclk n_20 GND efet
M544 notalucout DC78_phi2 GND GND efet
M545 n_1480 n_1570 dpc36_nIPC GND efet
M546 GND op_rti_rts n_1377 GND efet
M547 GND n_1316 n_20 GND efet
M548 GND n_AxB_6 _AxB_6_nC56 GND efet
M549 GND n_AxB_6 n_1390 GND efet
M550 nnT2BR cclk n_1269 GND efet
M551 GND n_781 n_1550 GND efet
M552 n_761 alu5 GND GND efet
M553 n_659 n_1153 Vdd GND efet
M554 GND n_1153 n_1639 GND efet
M555 GND pipeT4out n_395 GND efet
M556 AxB1 n_A_B_1 GND GND efet
M557 A_B1 n_A_B_1 GND GND efet
M558 n_1686 n_432 GND GND efet
M559 GND n_440 n_1555 GND efet
M560 GND n_635 ab14 GND efet
M561 n_1097 n_432 GND GND efet
M562 GND n_635 ab14 GND efet
M563 GND op_T0_shift_a n_11 GND efet
M564 n_191 n_790 GND GND efet
M565 GND pipephi2Reset0 n_819 GND efet
M566 op_T0_shift_a notir1 GND GND efet
M567 op_T0_tax notir1 GND GND efet
M568 op_T0_shift_right_a notir1 GND GND efet
M569 op_shift_right notir1 GND GND efet
M570 GND notir1 op_rol_ror GND efet
M571 op_shift notir1 GND GND efet
M572 op_T__shift_a notir1 GND GND efet
M573 op_T0_txa notir1 GND GND efet
M574 op_lsr_ror_dec_inc notir1 GND GND efet
M575 op_asl_rol notir1 GND GND efet
M576 y3 dpc1_SBY sb3 GND efet
M577 pcl7 dpc40_ADLPCL adl7 GND efet
M578 GND noty2 n_1491 GND efet
M579 GND op_T4_rti n_604 GND efet
M580 Vdd n_866 n_9 GND efet
M581 n_161 n_1113 GND GND efet
M582 brk_done n_861 GND GND efet
M583 GND n_1247 dpc8_nDBADD GND efet
M584 db6 n_471 db6 GND efet
M585 GND n_471 db6 GND efet
M586 GND n_471 db6 GND efet
M587 GND n_471 db6 GND efet
M588 GND n_471 db6 GND efet
M589 GND n_471 db6 GND efet
M590 GND n_471 db6 GND efet
M591 n_467 n_470 GND GND efet
M592 op_T2_abs notir2 GND GND efet
M593 n_246 ADL_ABL nABL0 GND efet
M594 GND op_ORS op_SUMS GND efet
M595 GND n_1488 n_545 GND efet
M596 n_570 n_122 GND GND efet
M597 A_B3 n_A_B_3 GND GND efet
M598 dpc0_YSB n_1247 GND GND efet
M599 GND n_572 n_1407 GND efet
M600 n_1501 dor7 GND GND efet
M601 n_23 dor7 GND GND efet
M602 n_1440 notRdy0 GND GND efet
M603 GND nA_B1 n_936 GND efet
M604 GND abh7 n_1153 GND efet
M605 n_659 abh7 GND GND efet
M606 pch1 dpc30_ADHPCH adh1 GND efet
M607 n_590 cp1 n_1178 GND efet
M608 GND nABH5 abh5 GND efet
M609 pch0 dpc30_ADHPCH adh0 GND efet
M610 n_617 abh1 GND GND efet
M611 n_676 abh1 GND GND efet
M612 npchp6 cclk n_1192 GND efet
M613 Vdd abh7 n_1639 GND efet
M614 n_1479 abl1 Vdd GND efet
M615 n_632 cclk n_339 GND efet
M616 D1x1 C1x5Reset GND GND efet
M617 GND n_753 n_1629 GND efet
M618 dasb5 n_753 n_1203 GND efet
M619 cclk n_1467 GND GND efet
M620 dpc35_PCHC n_923 GND GND efet
M621 Vdd n_1364 dpc16_EORS GND efet
M622 GND n_1364 n_108 GND efet
M623 n_1130 n_1258 GND GND efet
M624 idb4 cclk Vdd GND efet
M625 n_356 n_923 GND GND efet
M626 GND n_1619 n_586 GND efet
M627 n_642 n_951 Vdd GND efet
M628 n_1152 n_951 GND GND efet
M629 n_1190 cclk nots2 GND efet
M630 sb2 cclk Vdd GND efet
M631 n_1408 n_1044 n_1000 GND efet
M632 n_1379 cclk pipeUNK07 GND efet
M633 GND n_1643 n_410 GND efet
M634 GND pipeUNK03 n_1614 GND efet
M635 n_1723 pipeUNK03 GND GND efet
M636 PD_xxx010x1 n_1083 GND GND efet
M637 nC78 C67 n_1617 GND efet
M638 GND C67 nC67 GND efet
M639 Vdd n_102 rw GND efet
M640 n_1277 n_1020 GND GND efet
M641 n_548 s7 GND GND efet
M642 GND DBNeg n_648 GND efet
M643 PD_xxxx10x0 n_1083 GND GND efet
M644 npclp1 cclk n_1099 GND efet
M645 n_1130 cclk n_512 GND efet
M646 n_674 cclk n_745 GND efet
M647 GND C34 n_1179 GND efet
M648 n_695 C34 n_619 GND efet
M649 n_882 n_597 GND GND efet
M650 idb2 cclk Vdd GND efet
M651 GND RnWstretched n_298 GND efet
M652 n_269 AxB7 GND GND efet
M653 x_op_T3_ind_y ir2 GND GND efet
M654 op_rti_rts ir2 GND GND efet
M655 op_T2_jsr ir2 GND GND efet
M656 op_T5_jsr ir2 GND GND efet
M657 op_T4_ind_y ir2 GND GND efet
M658 op_T2_ind_y ir2 GND GND efet
M659 op_plp_pla ir2 GND GND efet
M660 op_T4_ind_x ir2 GND GND efet
M661 op_T2_stack_access ir2 GND GND efet
M662 op_T0_tya ir2 GND GND efet
M663 GND op_SRS n_160 GND efet
M664 op_EORS n_837 GND GND efet
M665 GND notidl1 idl1 GND efet
M666 GND n_1253 n_515 GND efet
M667 GND idb7 n_423 GND efet
M668 pipeUNK02 cclk n_774 GND efet
M669 GND n_590 alucin GND efet
M670 n_332 dpc4_SSB sb0 GND efet
M671 op_SRS cclk n_968 GND efet
M672 op_SUMS cclk n_415 GND efet
M673 ab0 n_855 Vdd GND efet
M674 ab0 n_855 Vdd GND efet
M675 ab0 n_855 Vdd GND efet
M676 ab0 n_855 Vdd GND efet
M677 n_202 n_646 GND GND efet
M678 GND notRdy0 n_1343 GND efet
M679 n_1080 n_1056 n_739 GND efet
M680 GND cclk n_881 GND efet
M681 n_631 n_878 GND GND efet
M682 adh7 cclk Vdd GND efet
M683 op_T2_abs ir4 GND GND efet
M684 op_T2_stack ir4 GND GND efet
M685 adl3 dpc21_ADDADL alu3 GND efet
M686 op_T2_jsr ir6 GND GND efet
M687 GND ir6 op_T4_brk_jsr GND efet
M688 op_T5_jsr ir6 GND GND efet
M689 op_shift ir6 GND GND efet
M690 GND ir6 op_T0_jsr GND efet
M691 GND ir6 op_T0_tay_ldy_not_idx GND efet
M692 GND ir6 op_T0_ora GND efet
M693 GND ir6 op_T5_brk GND efet
M694 GND ir6 op_T0_txa GND efet
M695 GND ir6 op_T0_tya GND efet
M696 n_87 cp1 idl1 GND efet
M697 GND ir5 op_T5_brk GND efet
M698 ir6 n_1675 GND GND efet
M699 n_363 n_16 n_1091 GND efet
M700 n_21 n_43 GND GND efet
M701 GND n_1449 n_944 GND efet
M702 n_550 n_384 GND GND efet
M703 n_176 cclk n_598 GND efet
M704 GND op_T0_cpy_iny n_1717 GND efet
M705 n_885 n_384 GND GND efet
M706 n_1592 cclk a7 GND efet
M707 GND cclk n_891 GND efet
M708 n_844 op_T__inx GND GND efet
M709 y2 dpc1_SBY sb2 GND efet
M710 nA_B1 dpc14_SRS naluresult0 GND efet
M711 naluresult1 dpc14_SRS nA_B2 GND efet
M712 nA_B3 dpc14_SRS naluresult2 GND efet
M713 naluresult3 dpc14_SRS nA_B4 GND efet
M714 naluresult4 dpc14_SRS nA_B5 GND efet
M715 naluresult5 dpc14_SRS nA_B6 GND efet
M716 naluresult6 dpc14_SRS nA_B7 GND efet
M717 n_469 cclk n_875 GND efet
M718 n_212 adh4 GND GND efet
M719 pd5_clearIR pd5 GND GND efet
M720 idb3 dpc43_DL_DB n_1661 GND efet
M721 n_830 n_1505 GND GND efet
M722 notx1 x1 GND GND efet
M723 idb0 dpc43_DL_DB n_719 GND efet
M724 GND pipenWR_phi2 notRnWprepad GND efet
M725 op_T__iny_dey ir4 GND GND efet
M726 GND nop_branch_bit6 n_846 GND efet
M727 idl4 notidl4 GND GND efet
M728 idb1 dpc43_DL_DB n_87 GND efet
M729 GND nA_B4 n_1310 GND efet
M730 n_1231 cclk pipeUNK21 GND efet
M731 nC78 n_748 GND GND efet
M732 GND ir7 op_T__asl_rol_a GND efet
M733 op_T__dex ir4 GND GND efet
M734 GND notx3 n_242 GND efet
M735 op_T0_cpx_inx ir4 GND GND efet
M736 y1 dpc1_SBY sb1 GND efet
M737 n_137 n_440 n_504 GND efet
M738 n_1649 brk_done GND GND efet
M739 n_300 brk_done GND GND efet
M740 n_1433 n_90 GND GND efet
M741 GND op_T3 n_256 GND efet
M742 nA_B4 alub4 n_185 GND efet
M743 GND nC12 n_433 GND efet
M744 GND nC12 C12 GND efet
M745 n_913 cp1 n_1274 GND efet
M746 db4 n_147 GND GND efet
M747 db4 n_147 GND GND efet
M748 n_1454 n_852 GND GND efet
M749 GND n_90 p6 GND efet
M750 n_1107 op_inc_nop n_1555 GND efet
M751 n_260 n_852 GND GND efet
M752 Vdd n_769 n_1072 GND efet
M753 GND n_769 n_1325 GND efet
M754 db4 n_147 db4 GND efet
M755 GND pcl4 n_1643 GND efet
M756 adl0 dpc5_SADL n_332 GND efet
M757 GND pcl6 n_232 GND efet
M758 GND s2 n_1190 GND efet
M759 pd0_clearIR pd0 GND GND efet
M760 n_922 n_270 BRtaken GND efet
M761 n_1300 cclk notir2 GND efet
M762 GND n_A_B_2 A_B2 GND efet
M763 n_1115 n_270 GND GND efet
M764 pclp3 npclp3 GND GND efet
M765 GND n_A_B_2 C23 GND efet
M766 GND nABH1 abh1 GND efet
M767 pcl1 dpc40_ADLPCL adl1 GND efet
M768 n_238 pipeUNK35 GND GND efet
M769 op_T5_ind_x _t5 GND GND efet
M770 op_T5_mem_ind_idx _t5 GND GND efet
M771 op_T5_brk _t5 GND GND efet
M772 DA_C01 nA_B0 n_1354 GND efet
M773 n_772 n_1674 GND GND efet
M774 op_T5_rti_rts _t5 GND GND efet
M775 xx_op_T5_jsr _t5 GND GND efet
M776 op_T5_rts _t5 GND GND efet
M777 op_T5_jsr _t5 GND GND efet
M778 op_T5_ind_y _t5 GND GND efet
M779 pcl3 dpc40_ADLPCL adl3 GND efet
M780 n_20 n_344 n_585 GND efet
M781 GND db4 n_490 GND efet
M782 pd3_clearIR pd3 GND GND efet
M783 Vdd n_826 ab8 GND efet
M784 n_1073 n_344 n_557 GND efet
M785 y7 dpc1_SBY sb7 GND efet
M786 alua4 dpc11_SBADD sb4 GND efet
M787 alua3 dpc11_SBADD sb3 GND efet
M788 n_25 n_192 GND GND efet
M789 GND pd0_clearIR n_409 GND efet
M790 n_307 nop_branch_bit7 GND GND efet
M791 n_1456 pipeT3out GND GND efet
M792 sb2 dpc11_SBADD alua2 GND efet
M793 sb1 dpc11_SBADD alua1 GND efet
M794 y1 cclk n_767 GND efet
M795 GND notalu4 alu4 GND efet
M796 GND op_T0_bit n_669 GND efet
M797 adl6 dpc10_ADLADD alub6 GND efet
M798 n_680 cclk n_1688 GND efet
M799 n_106 n_1528 GND GND efet
M800 adl1 dpc10_ADLADD alub1 GND efet
M801 adl4 dpc10_ADLADD alub4 GND efet
M802 adl7 dpc10_ADLADD alub7 GND efet
M803 ab13 n_1608 Vdd GND efet
M804 alub5 dpc10_ADLADD adl5 GND efet
M805 n_1126 cclk VEC0 GND efet
M806 GND n_1262 n_1151 GND efet
M807 n_618 dpc7_SS s6 GND efet
M808 GND n_101 n_1364 GND efet
M809 GND op_T0_ldx_tax_tsx n_844 GND efet
M810 n_998 dpc7_SS s3 GND efet
M811 n_1389 dpc7_SS s2 GND efet
M812 n_280 dpc7_SS s5 GND efet
M813 n_3 dpc7_SS s4 GND efet
M814 n_694 dpc7_SS s1 GND efet
M815 GND adh3 n_883 GND efet
M816 op_T0_bit ir4 GND GND efet
M817 op_T2_pha ir4 GND GND efet
M818 GND n_1642 nWR GND efet
M819 n_1129 cp1 GND GND efet
M820 n_541 cclk notir7 GND efet
M821 ADH_ABH n_1067 GND GND efet
M822 AxB5 n_647 GND GND efet
M823 n_867 nDA_ADD1 GND GND efet
M824 n_1556 nDA_ADD1 GND GND efet
M825 Vdd n_1633 ab5 GND efet
M826 adh3 dpc32_PCHADH pchp3 GND efet
M827 Vdd n_1633 ab5 GND efet
M828 adh1 dpc32_PCHADH pchp1 GND efet
M829 adh2 dpc32_PCHADH pchp2 GND efet
M830 op_T5_rti _t5 GND GND efet
M831 GND clock1 op_T0_clc_sec GND efet
M832 GND clock1 op_T0_cli_sei GND efet
M833 GND clock1 op_T0_jmp GND efet
M834 GND clock1 op_T0_brk_rti GND efet
M835 y2 cclk n_1491 GND efet
M836 op_T0_cld_sed clock1 GND GND efet
M837 op_T0_plp clock1 GND GND efet
M838 GND clock1 x_op_T0_bit GND efet
M839 GND n_587 n_299 GND efet
M840 GND n_236 n_272 GND efet
M841 alu6 dpc20_ADDSB06 sb6 GND efet
M842 alu5 dpc20_ADDSB06 sb5 GND efet
M843 n_388 DA_AxB2 GND GND efet
M844 n_1566 n_1221 GND GND efet
M845 GND n_812 n_1044 GND efet
M846 nWR cclk pipenWR_phi2 GND efet
M847 GND op_T0_cmp n_1560 GND efet
M848 n_1375 cp1 n_95 GND efet
M849 n_1089 cp1 n_1529 GND efet
M850 n_454 n_844 n_946 GND efet
M851 GND n_659 ab15 GND efet
M852 Vdd n_298 db7 GND efet
M853 Vdd n_298 db7 GND efet
M854 Vdd n_298 db7 GND efet
M855 Vdd n_298 db7 GND efet
M856 GND op_T5_rts n_272 GND efet
M857 npclp3 cclk n_1631 GND efet
M858 GND n_344 n_1316 GND efet
M859 GND n_739 n_479 GND efet
M860 GND n_1043 dpc40_ADLPCL GND efet
M861 GND pipeUNK15 H1x1 GND efet
M862 n_1257 n_1218 GND GND efet
M863 GND pd7 pd7_clearIR GND efet
M864 n_994 n_1034 Vdd GND efet
M865 GND n_1034 n_1545 GND efet
M866 GND n_717 n_1087 GND efet
M867 GND n_717 C1x5Reset GND efet
M868 n_1291 cp1 brk_done GND efet
M869 nC34 n_988 GND GND efet
M870 n_854 n_312 n_742 GND efet
M871 n_1558 pipeT2out GND GND efet
M872 GND idb3 DBZ GND efet
M873 GND n_94 n_1024 GND efet
M874 n_1211 n_862 GND GND efet
M875 GND n_849 dpc33_PCHDB GND efet
M876 npclp2 n_1411 GND GND efet
M877 noty3 y3 GND GND efet
M878 GND op_T5_jsr n_1219 GND efet
M879 n_1089 n_1574 GND GND efet
M880 GND clk0 n_519 GND efet
M881 n_644 cp1 n_428 GND efet
M882 ab10 n_1545 Vdd GND efet
M883 nA_B4 dpc15_ANDS naluresult4 GND efet
M884 nA_B2 dpc15_ANDS naluresult2 GND efet
M885 n_676 n_617 Vdd GND efet
M886 n_1474 cp1 notdor1 GND efet
M887 n_666 cp1 n_1380 GND efet
M888 n_334 brk_done GND GND efet
M889 n_1661 cp1 idl3 GND efet
M890 GND irline3 op_sty_cpy_mem GND efet
M891 n_1705 n_630 GND GND efet
M892 dpc39_PCLPCL n_1518 GND GND efet
M893 GND irline3 op_T0_iny_dey GND efet
M894 GND irline3 x_op_T0_tya GND efet
M895 n_171 n_1026 Vdd GND efet
M896 n_455 pipeUNK16 n_1082 GND efet
M897 op_T3_ind_y notir0 GND GND efet
M898 GND RnWstretched n_224 GND efet
M899 nA_B3 dpc15_ANDS naluresult3 GND efet
M900 GND op_rti_rts n_300 GND efet
M901 GND n_1177 n_1614 GND efet
M902 GND RnWstretched n_520 GND efet
M903 GND RnWstretched n_520 GND efet
M904 n_384 op_ANDS GND GND efet
M905 Vdd n_321 dpc33_PCHDB GND efet
M906 n_385 n_1377 GND GND efet
M907 nA_B0 dpc15_ANDS naluresult0 GND efet
M908 nC45 C45 GND GND efet
M909 nC56 C45 n_165 GND efet
M910 idl2 notidl2 GND GND efet
M911 GND notidl2 idl2 GND efet
M912 db2 GND GND GND efet
M913 GND notalu6 alu6 GND efet
M914 idl2 notidl2 GND GND efet
M915 n_1644 n_1457 n_1495 GND efet
M916 n_AxBxC_3 nC23 n_136 GND efet
M917 GND pch3 n_923 GND efet
M918 n_1347 cclk n_1527 GND efet
M919 n_AxB3__C23 nC23 GND GND efet
M920 NMIL cclk n_1252 GND efet
M921 n_1483 alua6 GND GND efet
M922 n_1211 n_1002 GND GND efet
M923 n_1470 n_1416 n_299 GND efet
M924 n_152 n_952 GND GND efet
M925 GND n_862 n_272 GND efet
M926 n_1717 op_T2_idx_x_xy n_1351 GND efet
M927 n_1709 dpc2_XSB sb1 GND efet
M928 op_ANDS n_669 GND GND efet
M929 db4 GND GND GND efet
M930 n_941 pipeUNK07 n_1111 GND efet
M931 n_A_B_1 dpc13_ORS naluresult1 GND efet
M932 GND n_218 n_1716 GND efet
M933 n_1594 cclk n_688 GND efet
M934 GND n_1395 Reset0 GND efet
M935 Reset0 n_1395 GND GND efet
M936 GND n_1072 db0 GND efet
M937 n_AxBxC_5 nC45 n_547 GND efet
M938 n_AxB5__C45 nC45 GND GND efet
M939 ab8 n_826 Vdd GND efet
M940 xx_op_T5_jsr ir4 GND GND efet
M941 op_T2_jmp_abs ir4 GND GND efet
M942 op_T4_jmp ir4 GND GND efet
M943 op_T5_rti_rts ir4 GND GND efet
M944 op_T2_php ir4 GND GND efet
M945 op_T2_php_pha ir4 GND GND efet
M946 op_push_pull ir4 GND GND efet
M947 op_T4_brk ir4 GND GND efet
M948 x_op_T3_plp_pla ir4 GND GND efet
M949 op_T__bit ir4 GND GND efet
M950 n_557 n_410 GND GND efet
M951 n_344 n_410 n_814 GND efet
M952 ab12 n_475 Vdd GND efet
M953 Vdd n_1639 ab15 GND efet
M954 GND cclk n_431 GND efet
M955 dpc10_ADLADD n_1541 Vdd GND efet
M956 GND pipeUNK29 n_1511 GND efet
M957 n_1189 pipeUNK29 GND GND efet
M958 GND RnWstretched n_1072 GND efet
M959 GND RnWstretched n_1072 GND efet
M960 op_T0_txa clock1 GND GND efet
M961 GND clock1 op_T0_tya GND efet
M962 alub7 dpc9_DBADD idb7 GND efet
M963 GND idb1 n_243 GND efet
M964 op_T3_ind_y ir3 GND GND efet
M965 alub6 dpc9_DBADD idb6 GND efet
M966 op_T0_jsr ir3 GND GND efet
M967 op_T2_ind_x ir3 GND GND efet
M968 op_T0_eor clock1 GND GND efet
M969 op_T5_brk ir3 GND GND efet
M970 op_T0 clock1 GND GND efet
M971 op_T0_ora clock1 GND GND efet
M972 GND clock1 op_T0_cmp GND efet
M973 GND clock1 op_T0_cpx_cpy_inx_iny GND efet
M974 GND clock1 op_T0_adc_sbc GND efet
M975 GND clock1 op_T0_sbc GND efet
M976 GND n_643 db3 GND efet
M977 GND n_643 db3 GND efet
M978 n_1181 cp1 n_69 GND efet
M979 nABL7 cclk n_171 GND efet
M980 Vdd n_1295 dpc25_SBDB GND efet
M981 n_1209 cclk n_663 GND efet
M982 n_1339 n_799 GND GND efet
M983 GND n_643 db3 GND efet
M984 dpc10_ADLADD n_1247 GND GND efet
M985 nop_set_C op_T__cpx_cpy_imm_zp GND GND efet
M986 n_388 DA_C01 GND GND efet
M987 n_662 n_625 GND GND efet
M988 GND pipeUNK09 n_781 GND efet
M989 GND pipeUNK09 n_1422 GND efet
M990 GND n_334 n_118 GND efet
M991 GND dpc12_0ADD alua6 GND efet
M992 GND dpc12_0ADD alua5 GND efet
M993 GND dpc12_0ADD alua1 GND efet
M994 GND dpc12_0ADD alua4 GND efet
M995 n_105 notalucin GND GND efet
M996 GND notalucin n_942 GND efet
M997 GND x_op_jmp n_510 GND efet
M998 GND x_op_jmp n_134 GND efet
M999 GND n_23 n_298 GND efet
M1000 db2 n_37 db2 GND efet
M1001 db2 n_37 GND GND efet
M1002 Vdd n_23 n_1501 GND efet
M1003 n_1093 n_968 GND GND efet
M1004 n_1705 cclk n_1020 GND efet
M1005 GND RnWstretched n_37 GND efet
M1006 n_1251 cclk y7 GND efet
M1007 GND n_236 n_1427 GND efet
M1008 GND n_288 n_798 GND efet
M1009 n_367 n_954 GND GND efet
M1010 GND adh1 n_1267 GND efet
M1011 n_494 cp1 n_514 GND efet
M1012 GND db5 n_1588 GND efet
M1013 nABL3 ADL_ABL n_864 GND efet
M1014 n_1347 n_550 GND GND efet
M1015 pipeUNK26 cclk n_132 GND efet
M1016 GND pd6_clearIR n_1309 GND efet
M1017 n_201 nop_branch_bit7 GND GND efet
M1018 aluvout n_408 GND GND efet
M1019 GND n_1699 n_913 GND efet
M1020 n_1141 cp1 n_101 GND efet
M1021 n_779 cclk n_805 GND efet
M1022 n_1480 n_1581 dpc36_nIPC GND efet
M1023 n_408 cclk notaluvout GND efet
M1024 idl6 notidl6 GND GND efet
M1025 GND n_347 n_191 GND efet
M1026 idl6 notidl6 GND GND efet
M1027 GND notidl6 idl6 GND efet
M1028 op_rti_rts irline3 GND GND efet
M1029 op_T2_jsr irline3 GND GND efet
M1030 GND n_698 VEC1 GND efet
M1031 n_1371 n_846 GND GND efet
M1032 nA_B6 dpc15_ANDS naluresult6 GND efet
M1033 naluresult7 dpc15_ANDS nA_B7 GND efet
M1034 op_T3_plp_pla irline3 GND GND efet
M1035 op_T5_rti irline3 GND GND efet
M1036 op_jmp irline3 GND GND efet
M1037 idb7 dpc37_PCLDB pclp7 GND efet
M1038 GND alub7 n_A_B_7 GND efet
M1039 GND irline3 op_T4_brk_jsr GND efet
M1040 GND n_853 n_387 GND efet
M1041 n_670 n_519 GND GND efet
M1042 op_T2_ind notir0 GND GND efet
M1043 op_sta_cmp notir0 GND GND efet
M1044 op_T__adc_sbc notir0 GND GND efet
M1045 op_T__ora_and_eor_adc notir0 GND GND efet
M1046 GND notir0 op_T0_adc_sbc GND efet
M1047 GND notir0 op_T0_sbc GND efet
M1048 op_T5_ind_y notir0 GND GND efet
M1049 GND notir0 op_T0_and GND efet
M1050 GND notir0 op_T0_acc GND efet
M1051 op_T0_lda notir0 GND GND efet
M1052 n_807 n_330 GND GND efet
M1053 GND n_1258 n_1716 GND efet
M1054 GND db3 n_1281 GND efet
M1055 GND nC56 C56 GND efet
M1056 n_112 nC56 C67 GND efet
M1057 n_878 cclk n_462 GND efet
M1058 GND RnWstretched n_1076 GND efet
M1059 GND RnWstretched n_1463 GND efet
M1060 p2 cp1 n_845 GND efet
M1061 n_1358 n_1109 GND GND efet
M1062 op_T4_brk_jsr ir4 GND GND efet
M1063 GND idb3 n_1621 GND efet
M1064 GND n_646 n_182 GND efet
M1065 GND ir7 op_T0_php_pha GND efet
M1066 pipeUNK14 cclk n_318 GND efet
M1067 GND ir7 op_rol_ror GND efet
M1068 op_T0_jsr ir7 GND GND efet
M1069 op_T5_brk ir7 GND GND efet
M1070 n_416 cp1 n_1016 GND efet
M1071 n_586 BRtaken n_1330 GND efet
M1072 n_586 BRtaken n_1330 GND efet
M1073 n_AxB3__C23 AxB3 GND GND efet
M1074 n_136 AxB3 GND GND efet
M1075 n_AxBxC_5 n_AxB5__C45 GND GND efet
M1076 pipeT4out cclk n_188 GND efet
M1077 n_1180 notRdy0 GND GND efet
M1078 n_1132 cp1 n_1087 GND efet
M1079 dpc9_DBADD n_225 GND GND efet
M1080 n_635 abh6 GND GND efet
M1081 n_1523 abh6 GND GND efet
M1082 Vdd abh6 n_963 GND efet
M1083 GND n_171 ab7 GND efet
M1084 GND n_334 Pout2 GND efet
M1085 n_643 RnWstretched GND GND efet
M1086 C78_phi2 cclk C78 GND efet
M1087 n_1517 n_572 GND GND efet
M1088 n_1348 A_B0 n_AxB_0 GND efet
M1089 n_169 n_139 GND GND efet
M1090 GND n_613 n_1159 GND efet
M1091 n_605 n_1440 n_779 GND efet
M1092 GND n_1673 n_754 GND efet
M1093 adh0 dpc32_PCHADH pchp0 GND efet
M1094 n_1636 ADL_ABL nABL2 GND efet
M1095 nABH0 cclk n_381 GND efet
M1096 GND dpc18_nDAA n_700 GND efet
M1097 adh4 dpc32_PCHADH pchp4 GND efet
M1098 Vdd n_1633 ab5 GND efet
M1099 Vdd n_1633 ab5 GND efet
M1100 n_1110 n_756 GND GND efet
M1101 n_146 dpc26_ACDB idb0 GND efet
M1102 n_929 dpc26_ACDB idb1 GND efet
M1103 n_1618 dpc26_ACDB idb2 GND efet
M1104 dpc39_PCLPCL cclk GND GND efet
M1105 GND n_31 n_132 GND efet
M1106 n_1583 A_B4 GND GND efet
M1107 GND nA_B6 n_112 GND efet
M1108 n_1654 dpc26_ACDB idb3 GND efet
M1109 idb4 dpc26_ACDB n_1344 GND efet
M1110 alub5 dpc9_DBADD idb5 GND efet
M1111 alub4 dpc9_DBADD idb4 GND efet
M1112 op_T2_mem_zp ir3 GND GND efet
M1113 op_T5_mem_ind_idx ir3 GND GND efet
M1114 x_op_T4_rti ir3 GND GND efet
M1115 op_T__cpx_cpy_imm_zp ir3 GND GND efet
M1116 alub3 dpc9_DBADD idb3 GND efet
M1117 idb2 dpc9_DBADD alub2 GND efet
M1118 n_1147 cp1 idl7 GND efet
M1119 alub1 dpc9_DBADD idb1 GND efet
M1120 op_T0_ldy_mem notir2 GND GND efet
M1121 GND n_732 clock1 GND efet
M1122 n_366 n_440 n_1012 GND efet
M1123 abh4 nABH4 GND GND efet
M1124 clk2out n_135 GND GND efet
M1125 clk2out n_135 GND GND efet
M1126 n_1090 cclk n_1683 GND efet
M1127 GND n_762 n_1018 GND efet
M1128 adh4 cclk Vdd GND efet
M1129 adl5 cclk Vdd GND efet
M1130 GND n_135 clk2out GND efet
M1131 clk2out n_135 GND GND efet
M1132 n_612 RnWstretched GND GND efet
M1133 n_586 cclk pipeBRtaken GND efet
M1134 GND _t3 op_T3_plp_pla GND efet
M1135 GND _t3 op_T3_stack_bit_jmp GND efet
M1136 op_sty_cpy_mem notir2 GND GND efet
M1137 GND n_621 n_355 GND efet
M1138 GND nDBE n_251 GND efet
M1139 GND D1x1 n_380 GND efet
M1140 GND n_1061 npchp3 GND efet
M1141 n_332 dpc7_SS s0 GND efet
M1142 idb0 cclk Vdd GND efet
M1143 GND n_201 n_1371 GND efet
M1144 GND op_T2_abs_access n_272 GND efet
M1145 n_307 n_846 GND GND efet
M1146 n_1183 fetch n_541 GND efet
M1147 n_1616 pipeUNK05 GND GND efet
M1148 GND idb5 DBZ GND efet
M1149 n_983 cclk nots0 GND efet
M1150 n_1162 cclk n_272 GND efet
M1151 n_472 notRdy0 n_395 GND efet
M1152 n_1615 notRdy0 n_468 GND efet
M1153 n_1100 abl0 GND GND efet
M1154 n_1495 cp1 p3 GND efet
M1155 n_855 abl0 Vdd GND efet
M1156 GND abl0 n_1660 GND efet
M1157 GND idb6 n_1416 GND efet
M1158 GND n_0_ADL2 adl2 GND efet
M1159 GND n_1404 n_133 GND efet
M1160 n_635 cclk nABH6 GND efet
M1161 GND n_1345 n_1500 GND efet
M1162 n_975 n_854 GND GND efet
M1163 pclp3 dpc38_PCLADL adl3 GND efet
M1164 adl2 dpc38_PCLADL pclp2 GND efet
M1165 pclp1 dpc38_PCLADL adl1 GND efet
M1166 GND cclk dpc26_ACDB GND efet
M1167 op_T0_cpy_iny irline3 GND GND efet
M1168 GND n_842 n_1479 GND efet
M1169 GND cclk dpc24_ACSB GND efet
M1170 pipeUNK40 cclk n_191 GND efet
M1171 n_626 DBNeg n_1249 GND efet
M1172 A_B4 n_A_B_4 GND GND efet
M1173 GND op_T__adc_sbc n_1455 GND efet
M1174 n_794 RnWstretched GND GND efet
M1175 op_T__shift_a notir3 GND GND efet
M1176 op_T0_tya notir3 GND GND efet
M1177 op_T3_jmp notir3 GND GND efet
M1178 op_plp_pla notir3 GND GND efet
M1179 op_T0_shift_a notir3 GND GND efet
M1180 op_T0_tay notir3 GND GND efet
M1181 GND notir3 op_T0_pla GND efet
M1182 op_T0_txa notir3 GND GND efet
M1183 op_T4_abs_idx notir3 GND GND efet
M1184 op_T0_tax notir3 GND GND efet
M1185 dasb7 dpc23_SBAC a7 GND efet
M1186 GND n_251 n_1028 GND efet
M1187 dasb5 dpc23_SBAC a5 GND efet
M1188 dasb6 dpc23_SBAC a6 GND efet
M1189 dasb3 dpc23_SBAC a3 GND efet
M1190 sb4 dpc23_SBAC a4 GND efet
M1191 dasb1 dpc23_SBAC a1 GND efet
M1192 a2 dpc23_SBAC dasb2 GND efet
M1193 n_A_B_2 alub2 GND GND efet
M1194 sb0 dpc23_SBAC a0 GND efet
M1195 GND op_T3_ind_x n_1107 GND efet
M1196 GND op_T3_ind_x n_604 GND efet
M1197 n_620 n_1371 GND GND efet
M1198 n_51 Pout3 GND GND efet
M1199 n_476 n_43 GND GND efet
M1200 GND n_453 n_1213 GND efet
M1201 GND n_1002 n_605 GND efet
M1202 n_1541 n_1477 GND GND efet
M1203 GND p2 n_334 GND efet
M1204 GND n_1002 n_605 GND efet
M1205 dpc14_SRS n_1593 Vdd GND efet
M1206 nWR n_335 GND GND efet
M1207 GND n_1696 rw GND efet
M1208 GND n_AxB_2 n_1572 GND efet
M1209 GND n_AxB_2 _AxB_2_nC12 GND efet
M1210 dpc40_ADLPCL n_1247 GND GND efet
M1211 n_440 n_24 GND GND efet
M1212 GND alua5 n_A_B_5 GND efet
M1213 GND op_rmw n_510 GND efet
M1214 GND abh2 n_994 GND efet
M1215 op_T5_jsr ir3 GND GND efet
M1216 op_T5_ind_y ir3 GND GND efet
M1217 op_branch_done ir3 GND GND efet
M1218 op_T2_brk ir3 GND GND efet
M1219 op_T3_jsr ir3 GND GND efet
M1220 op_T2_branch ir3 GND GND efet
M1221 op_T2_zp_zp_idx ir3 GND GND efet
M1222 op_T2_ind ir3 GND GND efet
M1223 op_T5_rts ir3 GND GND efet
M1224 n_937 pcl0 GND GND efet
M1225 n_1500 cclk n_526 GND efet
M1226 GND n_400 n_102 GND efet
M1227 Vdd n_400 n_1696 GND efet
M1228 GND n_834 n_1696 GND efet
M1229 GND n_834 n_400 GND efet
M1230 notx7 x7 GND GND efet
M1231 n_656 n_604 GND GND efet
M1232 ab10 n_1545 Vdd GND efet
M1233 GND op_shift_right n_1012 GND efet
M1234 GND dpc35_PCHC n_949 GND efet
M1235 GND dpc35_PCHC n_1406 GND efet
M1236 n_570 AxB5 GND GND efet
M1237 n_799 cclk nNMIG GND efet
M1238 n_949 n_83 n_523 GND efet
M1239 GND n_83 n_1406 GND efet
M1240 n_1433 nop_branch_bit6 GND GND efet
M1241 Vdd n_1315 n_381 GND efet
M1242 GND op_jsr n_134 GND efet
M1243 dor3 notdor3 GND GND efet
M1244 n_1693 cclk nNMIG GND efet
M1245 n_46 n_992 GND GND efet
M1246 GND op_T0_clc_sec n_889 GND efet
M1247 GND n_17 n_646 GND efet
M1248 Vdd n_17 clock1 GND efet
M1249 GND n_1247 dpc9_DBADD GND efet
M1250 n_992 n_595 GND GND efet
M1251 GND n_91 n_1256 GND efet
M1252 GND n_999 ab12 GND efet
M1253 ab12 n_999 GND GND efet
M1254 GND n_1258 n_813 GND efet
M1255 GND notRdy0 n_720 GND efet
M1256 GND n_1135 n_1203 GND efet
M1257 GND n_1135 n_1629 GND efet
M1258 ab12 n_999 GND GND efet
M1259 GND n_999 ab12 GND efet
M1260 GND n_1045 n_1371 GND efet
M1261 GND n_999 ab12 GND efet
M1262 pipeUNK17 cclk n_334 GND efet
M1263 ab1 n_1479 Vdd GND efet
M1264 AxB3 n_A_B_3 GND GND efet
M1265 n_452 alua2 GND GND efet
M1266 ab2 n_642 GND GND efet
M1267 ab2 n_642 GND GND efet
M1268 n_152 n_1002 GND GND efet
M1269 n_1230 n_43 GND GND efet
M1270 ab12 n_475 Vdd GND efet
M1271 s7 dpc6_SBS sb7 GND efet
M1272 ab2 n_642 GND GND efet
M1273 ab2 n_642 GND GND efet
M1274 DA_C45 nC45 GND GND efet
M1275 GND n_1194 Pout3 GND efet
M1276 GND pipeUNK33 n_1178 GND efet
M1277 n_824 cclk n_398 GND efet
M1278 idb5 dpc25_SBDB sb5 GND efet
M1279 idb6 dpc25_SBDB sb6 GND efet
M1280 sb7 dpc25_SBDB idb7 GND efet
M1281 n_1065 cclk n_1124 GND efet
M1282 n_728 VEC0 GND GND efet
M1283 n_972 n_388 DC34 GND efet
M1284 GND a0 n_5 GND efet
M1285 GND op_T2_abs_y n_1717 GND efet
M1286 ab11 n_359 GND GND efet
M1287 n_636 op_T2_branch GND GND efet
M1288 n_111 cclk pd2 GND efet
M1289 n_62 cclk pd7 GND efet
M1290 GND dor6 n_466 GND efet
M1291 n_1290 cp1 n_698 GND efet
M1292 nIRQP IRQP GND GND efet
M1293 GND notalu1 alu1 GND efet
M1294 n_374 cclk pd6 GND efet
M1295 nIRQP IRQP GND GND efet
M1296 n_1718 cp1 n_671 GND efet
M1297 n_1030 n_757 GND GND efet
M1298 GND n_1024 n_1069 GND efet
M1299 n_1130 n_192 GND GND efet
M1300 idb4 dpc43_DL_DB n_1095 GND efet
M1301 GND op_T0_cli_sei n_1065 GND efet
M1302 n_1610 DA_AB2 GND GND efet
M1303 DA_AxB2 DA_AB2 GND GND efet
M1304 n_566 n_243 n_802 GND efet
M1305 GND pipeUNK17 n_511 GND efet
M1306 idb2 dpc43_DL_DB n_1424 GND efet
M1307 ab14 n_963 Vdd GND efet
M1308 notRdy0 cp1 n_1679 GND efet
M1309 x_op_push_pull ir7 GND GND efet
M1310 n_223 cp1 n_1215 GND efet
M1311 GND notir7 op_T0_txs GND efet
M1312 GND notir7 op_T0_ldx_tax_tsx GND efet
M1313 GND notir7 op_T0_cpx_inx GND efet
M1314 GND notir7 op_from_x GND efet
M1315 GND notir7 x_op_T0_txa GND efet
M1316 GND notir7 op_T0_dex GND efet
M1317 GND notir7 op_T0_cpy_iny GND efet
M1318 op_xy notir7 GND GND efet
M1319 n_A_B_4 alub4 GND GND efet
M1320 GND n_1258 nWR GND efet
M1321 GND notir7 op_T__dex GND efet
M1322 op_T__inx notir7 GND GND efet
M1323 GND notir5 x_op_T0_bit GND efet
M1324 GND notir5 x_op_T__adc_sbc GND efet
M1325 GND notir5 op_T__bit GND efet
M1326 GND notir5 x_op_T3_plp_pla GND efet
M1327 GND notir5 xx_op_T5_jsr GND efet
M1328 GND notir5 op_jsr GND efet
M1329 GND notir5 op_T5_rts GND efet
M1330 GND notir5 op_T3_jsr GND efet
M1331 GND notir5 op_T0_and GND efet
M1332 GND notir5 op_T0_bit GND efet
M1333 n_927 cclk notir4 GND efet
M1334 n_1335 n_628 GND GND efet
M1335 idb5 cclk Vdd GND efet
M1336 GND n_50 n_629 GND efet
M1337 n_440 cclk pipeUNK39 GND efet
M1338 n_1716 op_T3_branch GND GND efet
M1339 n_1708 op_T3_branch GND GND efet
M1340 GND op_T0_jmp n_256 GND efet
M1341 GND npclp4 pclp4 GND efet
M1342 GND GND db7 GND efet
M1343 GND pipenT0 n_964 GND efet
M1344 n_1304 op_T0_sbc GND GND efet
M1345 dpc7_SS n_35 Vdd GND efet
M1346 n_1180 pipenT0 GND GND efet
M1347 _t5 n_378 GND GND efet
M1348 n_71 n_35 GND GND efet
M1349 GND n_1655 n_182 GND efet
M1350 n_1356 a6 GND GND efet
M1351 n_1041 abl3 Vdd GND efet
M1352 GND pipeUNK11 n_1214 GND efet
M1353 GND ir5 op_T2_jmp_abs GND efet
M1354 GND ir5 x_op_T4_rti GND efet
M1355 GND ir5 op_store GND efet
M1356 GND ir5 op_T4_brk GND efet
M1357 GND ir5 op_T2_php GND efet
M1358 GND ir5 op_T2_php_pha GND efet
M1359 GND ir5 op_T2_brk GND efet
M1360 GND ir5 op_sta_cmp GND efet
M1361 GND ir5 op_T0_brk_rti GND efet
M1362 op_brk_rti ir5 GND GND efet
M1363 n_1560 n_1055 GND GND efet
M1364 n_931 cp1 n_1674 GND efet
M1365 n_1526 cp1 n_1450 GND efet
M1366 n_638 op_T0 GND GND efet
M1367 GND n_512 n_154 GND efet
M1368 dpc6_SBS n_1247 GND GND efet
M1369 GND n_1427 n_1448 GND efet
M1370 GND n_223 n_1357 GND efet
M1371 GND n_1219 n_1002 GND efet
M1372 idb0 H1x1 Pout0 GND efet
M1373 n_604 cclk n_1477 GND efet
M1374 GND ir1 n_1133 GND efet
M1375 nABH5 ADH_ABH n_1353 GND efet
M1376 GND ir1 notir1 GND efet
M1377 ab12 n_475 Vdd GND efet
M1378 GND n_1708 n_236 GND efet
M1379 GND n_1399 n_1105 GND efet
M1380 GND x3 notx3 GND efet
M1381 n_14 n_323 GND GND efet
M1382 GND n_355 n_593 GND efet
M1383 Vdd n_355 dpc4_SSB GND efet
M1384 ab1 n_1479 Vdd GND efet
M1385 ab1 n_1479 Vdd GND efet
M1386 Vdd n_1479 ab1 GND efet
M1387 ab1 n_1479 Vdd GND efet
M1388 n_814 n_392 GND GND efet
M1389 n_557 n_392 GND GND efet
M1390 noty4 y4 GND GND efet
M1391 pipeUNK35 cclk n_501 GND efet
M1392 op_T2_abs_y _t2 GND GND efet
M1393 GND n_1565 n_1218 GND efet
M1394 notRdy0 cp1 n_1276 GND efet
M1395 op_T2 _t2 GND GND efet
M1396 op_T2_abs _t2 GND GND efet
M1397 op_T2_idx_x_xy _t2 GND GND efet
M1398 op_T2_ind_x _t2 GND GND efet
M1399 op_T2_ADL_ADD _t2 GND GND efet
M1400 op_T2_stack _t2 GND GND efet
M1401 n_163 n_249 GND GND efet
M1402 dpc22_nDSA n_599 GND GND efet
M1403 GND n_462 n_1278 GND efet
M1404 dpc1_SBY n_692 Vdd GND efet
M1405 n_441 n_692 GND GND efet
M1406 n_1225 op_T2_ind GND GND efet
M1407 Vdd n_291 dpc41_DL_ADL GND efet
M1408 GND n_278 n_1488 GND efet
M1409 GND op_branch_done n_10 GND efet
M1410 INTG n_760 GND GND efet
M1411 GND op_T4_ind_x n_300 GND efet
M1412 n_961 cp1 notdor5 GND efet
M1413 n_186 n_507 n_1082 GND efet
M1414 n_279 n_507 GND GND efet
M1415 p6 H1x1 idb6 GND efet
M1416 n_1501 RnWstretched GND GND efet
M1417 GND n_200 n_57 GND efet
M1418 n_293 n_200 n_1367 GND efet
M1419 GND n_200 n_1486 GND efet
M1420 n_952 cclk n_1509 GND efet
M1421 n_1501 RnWstretched GND GND efet
M1422 Vdd cclk sb3 GND efet
M1423 GND pipeUNK39 n_2 GND efet
M1424 n_1376 cp1 notdor2 GND efet
M1425 GND x_op_T4_rti n_327 GND efet
M1426 AxB3 n_988 GND GND efet
M1427 n_34 cclk nots3 GND efet
M1428 n_AxBxC_4 dpc17_SUMS naluresult4 GND efet
M1429 n_AxBxC_5 dpc17_SUMS naluresult5 GND efet
M1430 naluresult6 dpc17_SUMS n_AxBxC_6 GND efet
M1431 naluresult7 dpc17_SUMS n_AxBxC_7 GND efet
M1432 n_1409 cp1 n_916 GND efet
M1433 GND n_666 n_862 GND efet
M1434 dpc37_PCLDB n_1323 GND GND efet
M1435 GND npchp7 pchp7 GND efet
M1436 n_611 n_1509 GND GND efet
M1437 n_1433 n_201 GND GND efet
M1438 DBNeg idb7 GND GND efet
M1439 GND idb7 DBZ GND efet
M1440 n_146 cclk a0 GND efet
M1441 GND ir7 nop_branch_bit7 GND efet
M1442 n_1244 op_xy GND GND efet
M1443 n_1491 dpc0_YSB sb2 GND efet
M1444 GND n_647 n_570 GND efet
M1445 GND pipeVectorA2 n_815 GND efet
M1446 GND n_1488 n_1547 GND efet
M1447 cp1 n_1105 GND GND efet
M1448 n_494 adh7 GND GND efet
M1449 GND ir5 op_T__dex GND efet
M1450 GND ir5 op_T__iny_dey GND efet
M1451 GND ir5 x_op_T0_tya GND efet
M1452 GND ir5 op_T0_cpy_iny GND efet
M1453 GND ir5 op_sty_cpy_mem GND efet
M1454 GND ir5 op_T0_iny_dey GND efet
M1455 GND ir5 op_from_x GND efet
M1456 op_T0_txs ir5 GND GND efet
M1457 GND ir5 x_op_T0_txa GND efet
M1458 GND ir5 op_T0_dex GND efet
M1459 n_959 pipeUNK20 GND GND efet
M1460 GND n_210 ab5 GND efet
M1461 GND RnWstretched n_42 GND efet
M1462 GND n_128 n_1592 GND efet
M1463 GND n_210 ab5 GND efet
M1464 n_482 A_B6 GND GND efet
M1465 GND n_210 ab5 GND efet
M1466 GND n_210 ab5 GND efet
M1467 GND RnWstretched n_1613 GND efet
M1468 GND RnWstretched n_42 GND efet
M1469 s5 dpc6_SBS sb5 GND efet
M1470 s6 dpc6_SBS sb6 GND efet
M1471 nA_B0 alub0 n_316 GND efet
M1472 GND alub0 n_A_B_0 GND efet
M1473 GND brk_done n_1087 GND efet
M1474 n_1178 pipeUNK32 GND GND efet
M1475 n_1117 cclk pipeVectorA1 GND efet
M1476 n_797 cp1 notdor4 GND efet
M1477 GND n_805 n_1534 GND efet
M1478 n_326 cclk a6 GND efet
M1479 GND n_954 n_513 GND efet
M1480 GND n_1026 n_322 GND efet
M1481 dpc31_PCHPCH n_611 Vdd GND efet
M1482 n_917 notRdy0 GND GND efet
M1483 op_T__cpx_cpy_imm_zp irline3 GND GND efet
M1484 n_255 n_611 GND GND efet
M1485 n_227 pd4_clearIR GND GND efet
M1486 dpc2_XSB n_602 GND GND efet
M1487 ab4 n_634 Vdd GND efet
M1488 n_1099 n_1542 n_1568 GND efet
M1489 Vdd n_634 ab4 GND efet
M1490 Vdd n_634 ab4 GND efet
M1491 GND D1x1 n_1471 GND efet
M1492 n_392 n_386 GND GND efet
M1493 n_1184 n_1253 n_1498 GND efet
M1494 n_903 n_1253 GND GND efet
M1495 dpc34_PCLC n_386 GND GND efet
M1496 n_700 cclk n_1565 GND efet
M1497 GND y7 noty7 GND efet
M1498 n_119 cclk notir1 GND efet
M1499 op_T2_php_pha _t2 GND GND efet
M1500 op_T2_jmp_abs _t2 GND GND efet
M1501 op_T2_mem_zp _t2 GND GND efet
M1502 n_1360 cp1 n_1091 GND efet
M1503 GND op_T2_ind_x n_1106 GND efet
M1504 GND n_1679 n_1262 GND efet
M1505 pipeUNK41 cclk n_504 GND efet
M1506 op_ANDS cclk n_1574 GND efet
M1507 n_384 op_ANDS GND GND efet
M1508 n_515 cclk n_1411 GND efet
M1509 pch1 dpc31_PCHPCH pchp1 GND efet
M1510 pch0 dpc31_PCHPCH pchp0 GND efet
M1511 pch3 dpc31_PCHPCH pchp3 GND efet
M1512 GND dpc29_0ADH17 adh5 GND efet
M1513 n_161 cclk GND GND efet
M1514 GND dpc29_0ADH17 adh3 GND efet
M1515 n_616 op_T0_ldy_mem GND GND efet
M1516 n_1130 n_862 GND GND efet
M1517 idb4 dpc37_PCLDB pclp4 GND efet
M1518 n_133 cclk GND GND efet
M1519 GND dpc29_0ADH17 adh4 GND efet
M1520 n_838 n_581 GND GND efet
M1521 n_835 dpc34_PCLC GND GND efet
M1522 n_134 op_brk_rti GND GND efet
M1523 n_11 n_397 n_1563 GND efet
M1524 GND GND db5 GND efet
M1525 n_1030 n_269 DC78 GND efet
M1526 GND op_sty_cpy_mem n_1397 GND efet
M1527 GND n_1247 dpc24_ACSB GND efet
M1528 n_1312 n_1693 GND GND efet
M1529 GND nnT2BR n_405 GND efet
M1530 nABL0 cclk n_1100 GND efet
M1531 n_793 pipeUNK13 GND GND efet
M1532 GND ir7 op_T3_jmp GND efet
M1533 op_T2_jsr ir7 GND GND efet
M1534 GND ir7 op_rti_rts GND efet
M1535 GND ir7 op_plp_pla GND efet
M1536 GND ir7 op_T__ora_and_eor_adc GND efet
M1537 GND ir7 op_T2_stack_access GND efet
M1538 GND ir7 op_T5_jsr GND efet
M1539 GND ir7 op_shift GND efet
M1540 op_T0_pla ir7 GND GND efet
M1541 GND ir7 op_T__shift_a GND efet
M1542 sync n_417 Vdd GND efet
M1543 sync n_417 Vdd GND efet
M1544 GND NMIP nNMIP GND efet
M1545 GND Reset0 n_14 GND efet
M1546 dpc8_nDBADD n_1534 Vdd GND efet
M1547 GND n_1534 n_763 GND efet
M1548 dasb1 n_36 n_1322 GND efet
M1549 n_1045 n_69 GND GND efet
M1550 Vdd n_417 sync GND efet
M1551 GND n_36 n_735 GND efet
M1552 GND a7 n_128 GND efet
M1553 n_275 n_773 GND GND efet
M1554 n_1348 nA_B0 GND GND efet
M1555 n_1703 n_16 n_468 GND efet
M1556 n_1575 n_1360 GND GND efet
M1557 GND x_op_T__adc_sbc nop_set_C GND efet
M1558 GND nABL5 abl5 GND efet
M1559 GND n_946 n_384 GND efet
M1560 n_366 op_T0_shift_right_a GND GND efet
M1561 n_AxB_4 nA_B4 n_1583 GND efet
M1562 op_T3_ind_x ir4 GND GND efet
M1563 n_577 cp1 n_1046 GND efet
M1564 GND n_476 n_956 GND efet
M1565 dpc12_0ADD n_476 Vdd GND efet
M1566 Vdd n_42 db3 GND efet
M1567 GND s4 n_973 GND efet
M1568 GND n_1471 p4 GND efet
M1569 n_1351 op_xy GND GND efet
M1570 n_961 idb5 GND GND efet
M1571 op_T4_rti ir4 GND GND efet
M1572 op_T2_php notir3 GND GND efet
M1573 op_T3_stack_bit_jmp ir4 GND GND efet
M1574 op_T2_jsr ir4 GND GND efet
M1575 op_rti_rts ir4 GND GND efet
M1576 op_T4_ind_x ir4 GND GND efet
M1577 n_897 cclk n_1211 GND efet
M1578 n_12 notRdy0 n_1091 GND efet
M1579 n_1456 notRdy0 n_428 GND efet
M1580 Vdd n_1076 db4 GND efet
M1581 Vdd n_1076 db4 GND efet
M1582 ab13 n_869 GND GND efet
M1583 ab13 n_869 GND GND efet
M1584 n_757 DA_C45 n_939 GND efet
M1585 GND op_ror n_544 GND efet
M1586 n_280 dpc4_SSB sb5 GND efet
M1587 op_plp_pla ir4 GND GND efet
M1588 dpc3_SBX n_662 GND GND efet
M1589 GND alub1 n_A_B_1 GND efet
M1590 n_86 abl4 GND GND efet
M1591 GND n_469 npchp5 GND efet
M1592 GND op_T2_jsr n_1649 GND efet
M1593 GND op_T4_rts n_1464 GND efet
M1594 nA_B1 alub1 n_189 GND efet
M1595 n_767 dpc0_YSB sb1 GND efet
M1596 n_634 abl4 Vdd GND efet
M1597 GND abl4 n_1676 GND efet
M1598 GND clearIR pd7_clearIR GND efet
M1599 n_705 cp1 n_1668 GND efet
M1600 n_1211 op_T2_abs_access GND GND efet
M1601 GND n_1492 n_1445 GND efet
M1602 GND n_1492 n_1457 GND efet
M1603 GND n_266 n_525 GND efet
M1604 GND n_1357 n_188 GND efet
M1605 n_246 cp1 n_123 GND efet
M1606 n_7 dor6 Vdd GND efet
M1607 GND n_0_ADL0 adl0 GND efet
M1608 GND n_A_B_6 A_B6 GND efet
M1609 n_854 n_975 GND GND efet
M1610 n_678 n_644 GND GND efet
M1611 n_797 idb4 GND GND efet
M1612 n_260 n_1205 GND GND efet
M1613 n_1454 n_1205 dasb7 GND efet
M1614 C67 n_A_B_6 GND GND efet
M1615 op_ORS cclk n_88 GND efet
M1616 sb7 cclk Vdd GND efet
M1617 dpc12_0ADD n_956 GND GND efet
M1618 n_852 sb7 GND GND efet
M1619 n_852 sb7 GND GND efet
M1620 GND n_1464 n_1109 GND efet
M1621 n_227 cp1 n_703 GND efet
M1622 n_62 db7 GND GND efet
M1623 n_1338 cp1 n_720 GND efet
M1624 n_1209 n_609 n_1264 GND efet
M1625 GND n_1412 n_384 GND efet
M1626 Vdd n_7 db6 GND efet
M1627 n_1192 n_609 n_1547 GND efet
M1628 n_629 cclk n_760 GND efet
M1629 GND nnT2BR n_1427 GND efet
M1630 GND db6 n_1638 GND efet
M1631 ab11 n_359 GND GND efet
M1632 GND n_206 n_465 GND efet
M1633 nABH2 ADH_ABH n_836 GND efet
M1634 GND nA_B2 n_716 GND efet
M1635 op_T0_cld_sed notir6 GND GND efet
M1636 op_lsr_ror_dec_inc notir6 GND GND efet
M1637 op_T2_jmp_abs notir6 GND GND efet
M1638 GND notir6 op_T__cpx_cpy_imm_zp GND efet
M1639 GND notir6 op_T__cmp GND efet
M1640 x_op_T4_rti _t4 GND GND efet
M1641 GND _t4 op_T4_jmp GND efet
M1642 GND _t4 op_T4_brk GND efet
M1643 GND _t4 x_op_T4_ind_y GND efet
M1644 GND _t4 op_T4 GND efet
M1645 GND _t4 op_T4_abs_idx GND efet
M1646 op_T4_ind_x _t4 GND GND efet
M1647 op_T4_ind_y _t4 GND GND efet
M1648 GND ir7 op_brk_rti GND efet
M1649 GND ir7 op_T0_jmp GND efet
M1650 n_916 n_1517 GND GND efet
M1651 GND ir7 op_jsr GND efet
M1652 op_T4_brk ir7 GND GND efet
M1653 GND ir7 op_push_pull GND efet
M1654 GND ir7 op_T2_php_pha GND efet
M1655 op_T2_php ir7 GND GND efet
M1656 GND n_1109 n_1649 GND efet
M1657 GND p1 n_318 GND efet
M1658 GND n_43 n_1223 GND efet
M1659 GND notidl0 idl0 GND efet
M1660 idl0 notidl0 GND GND efet
M1661 GND n_1683 n_966 GND efet
M1662 dpc1_SBY n_441 GND GND efet
M1663 dpc6_SBS n_282 GND GND efet
M1664 GND npchp5 pchp5 GND efet
M1665 GND notir7 op_T0_lda GND efet
M1666 GND notir7 op_T0_tay GND efet
M1667 GND notir7 op_T0_tax GND efet
M1668 GND notir7 op_sta_cmp GND efet
M1669 GND notir7 op_store GND efet
M1670 GND notir7 op_T__cmp GND efet
M1671 GND notir7 op_T__cpx_cpy_abs GND efet
M1672 op_T__cpx_cpy_imm_zp notir7 GND GND efet
M1673 op_T0_cld_sed notir7 GND GND efet
M1674 GND notir7 op_clv GND efet
M1675 GND notalu0 alu0 GND efet
M1676 GND n_982 n_1141 GND efet
M1677 n_453 pch7 GND GND efet
M1678 GND op_T2_jmp_abs n_368 GND efet
M1679 GND n_637 notaluvout GND efet
M1680 ab13 n_1608 Vdd GND efet
M1681 n_1231 n_1409 GND GND efet
M1682 n_11 op_ANDS GND GND efet
M1683 n_1135 sb5 GND GND efet
M1684 n_1695 alua7 GND GND efet
M1685 GND alua7 n_A_B_7 GND efet
M1686 nABL4 cclk n_86 GND efet
M1687 n_1117 n_70 GND GND efet
M1688 n_10 n_1211 GND GND efet
M1689 GND n_617 n_1140 GND efet
M1690 GND n_A_B_7 AxB7 GND efet
M1691 A_B7 n_A_B_7 GND GND efet
M1692 GND x_op_T3_ind_y n_300 GND efet
M1693 n_1379 x_op_T0_bit GND GND efet
M1694 GND n_1625 n_90 GND efet
M1695 n_1515 PD_n_0xx0xx0x GND GND efet
M1696 n_1295 n_1527 GND GND efet
M1697 GND op_T5_ind_y n_595 GND efet
M1698 n_275 n_1697 GND GND efet
M1699 n_673 op_T0_adc_sbc n_1053 GND efet
M1700 n_703 fetch n_927 GND efet
M1701 n_340 op_clv GND GND efet
M1702 GND notRdy0 brk_done GND efet
M1703 n_869 abh5 GND GND efet
M1704 idb2 dpc37_PCLDB pclp2 GND efet
M1705 Vdd abh5 n_1608 GND efet
M1706 n_1423 abh5 GND GND efet
M1707 n_931 n_415 GND GND efet
M1708 n_1375 n_88 GND GND efet
M1709 x5 dpc3_SBX sb5 GND efet
M1710 sb6 dpc3_SBX x6 GND efet
M1711 Vdd n_1677 n_999 GND efet
M1712 GND n_1677 n_475 GND efet
M1713 n_865 cclk n_958 GND efet
M1714 x2 dpc3_SBX sb2 GND efet
M1715 x3 dpc3_SBX sb3 GND efet
M1716 ADH_ABH n_582 Vdd GND efet
M1717 GND n_582 n_1067 GND efet
M1718 n_50 cp1 INTG GND efet
M1719 GND n_43 n_611 GND efet
M1720 GND op_T0_txs n_1106 GND efet
M1721 db0 n_1325 Vdd GND efet
M1722 n_396 cclk n_796 GND efet
M1723 n_1105 n_1715 Vdd GND efet
M1724 GND dpc12_0ADD alua7 GND efet
M1725 n_149 alu6 GND GND efet
M1726 GND s1 n_1711 GND efet
M1727 GND op_T0_tya n_1455 GND efet
M1728 y0 cclk n_564 GND efet
M1729 n_659 cclk nABH7 GND efet
M1730 n_726 op_T5_ind_x GND GND efet
M1731 GND op_T5_ind_x n_256 GND efet
M1732 GND n_1463 n_1076 GND efet
M1733 Vdd n_1463 n_147 GND efet
M1734 n_1209 n_1213 GND GND efet
M1735 GND n_228 dpc30_ADHPCH GND efet
M1736 GND op_T0_tay n_11 GND efet
M1737 n_1380 n_819 GND GND efet
M1738 dpc19_ADDSB7 n_714 Vdd GND efet
M1739 n_818 n_43 GND GND efet
M1740 nABL5 cclk n_210 GND efet
M1741 n_1500 dpc36_nIPC n_1706 GND efet
M1742 GND dpc36_nIPC n_1345 GND efet
M1743 n_1101 n_813 n_1508 GND efet
M1744 GND op_plp_pla n_1107 GND efet
M1745 GND n_1002 n_1130 GND efet
M1746 GND ir7 op_T0_eor GND efet
M1747 adl1 dpc5_SADL n_694 GND efet
M1748 n_1592 dpc24_ACSB sb7 GND efet
M1749 pchp0 npchp0 GND GND efet
M1750 nABL2 cclk n_642 GND efet
M1751 op_T2_abs_y notir3 GND GND efet
M1752 GND dpc36_nIPC dpc34_PCLC GND efet
M1753 x_op_T0_tya notir3 GND GND efet
M1754 GND notir3 op_T0_iny_dey GND efet
M1755 op_T0_dex notir3 GND GND efet
M1756 x_op_T0_txa notir3 GND GND efet
M1757 GND pipeUNK21 n_572 GND efet
M1758 n_1092 n_118 GND GND efet
M1759 ab0 n_1100 GND GND efet
M1760 n_61 sb6 GND GND efet
M1761 GND n_1676 n_634 GND efet
M1762 n_1347 op_T0_shift_a GND GND efet
M1763 notir0 cclk n_310 GND efet
M1764 n_86 n_1676 Vdd GND efet
M1765 ab0 n_1100 GND GND efet
M1766 ab0 n_1100 GND GND efet
M1767 adh2 dpc27_SBADH sb2 GND efet
M1768 adh3 dpc27_SBADH sb3 GND efet
M1769 GND cp1 n_1247 GND efet
M1770 n_38 cp1 GND GND efet
M1771 n_882 n_1252 GND GND efet
M1772 sb6 dpc27_SBADH adh6 GND efet
M1773 adh7 dpc27_SBADH sb7 GND efet
M1774 adh0 dpc27_SBADH sb0 GND efet
M1775 y0 dpc1_SBY sb0 GND efet
M1776 GND irline3 op_T5_rti_rts GND efet
M1777 op_T4_jmp irline3 GND GND efet
M1778 GND irline3 op_T2_jmp_abs GND efet
M1779 GND irline3 xx_op_T5_jsr GND efet
M1780 op_T4_brk irline3 GND GND efet
M1781 op_push_pull irline3 GND GND efet
M1782 op_T2_php_pha irline3 GND GND efet
M1783 op_T2_php irline3 GND GND efet
M1784 op_T0_cli_sei irline3 GND GND efet
M1785 x_op_T3_plp_pla irline3 GND GND efet
M1786 dpc26_ACDB n_1247 GND GND efet
M1787 n_1039 pipeUNK40 GND GND efet
M1788 n_1474 idb1 GND GND efet
M1789 dpc30_ADHPCH n_1247 GND GND efet
M1790 GND so n_1650 GND efet
M1791 n_939 n_647 GND GND efet
M1792 nABL3 cclk n_138 GND efet
M1793 n_1270 n_509 GND GND efet
M1794 GND n_653 n_390 GND efet
M1795 GND n_236 n_79 GND efet
M1796 n_14 n_671 GND GND efet
M1797 nC34 C23 n_924 GND efet
M1798 nC23 C23 GND GND efet
M1799 alub2 dpc8_nDBADD n_458 GND efet
M1800 alub4 dpc8_nDBADD n_478 GND efet
M1801 GND n_1269 n_1249 GND efet
M1802 n_753 n_811 GND GND efet
M1803 GND ir0 notir0 GND efet
M1804 n_1133 ir0 GND GND efet
M1805 GND op_T3_jmp n_980 GND efet
M1806 n_80 n_1130 GND GND efet
M1807 dpc26_ACDB n_525 Vdd GND efet
M1808 n_800 n_525 GND GND efet
M1809 GND n_1305 dpc17_SUMS GND efet
M1810 GND n_1708 n_1055 GND efet
M1811 GND op_T0_adc_sbc n_1000 GND efet
M1812 n_861 n_1452 GND GND efet
M1813 GND a3 n_947 GND efet
M1814 n_1247 cp1 GND GND efet
M1815 op_T4_rts ir3 GND GND efet
M1816 GND clock1 op_T0_php_pha GND efet
M1817 PD_1xx000x0 pd4_clearIR GND GND efet
M1818 GND pd4_clearIR PD_0xx0xx0x GND efet
M1819 GND notir5 op_clv GND efet
M1820 GND notir5 op_T0_plp GND efet
M1821 ab6 n_1254 GND GND efet
M1822 n_1497 pipeUNK41 GND GND efet
M1823 GND n_1254 ab6 GND efet
M1824 GND n_1254 ab6 GND efet
M1825 PD_xxx010x1 pd4_clearIR GND GND efet
M1826 GND n_1254 ab6 GND efet
M1827 GND n_1585 n_962 GND efet
M1828 n_1489 n_A_B_7 GND GND efet
M1829 GND nABL0 abl0 GND efet
M1830 nWR n_440 GND GND efet
M1831 n_104 n_440 GND GND efet
M1832 n_812 n_440 GND GND efet
M1833 n_1368 n_1578 GND GND efet
M1834 GND n_1027 n_476 GND efet
M1835 n_368 op_T4_jmp GND GND efet
M1836 n_104 op_T4_jmp GND GND efet
M1837 op_T2_idx_x_xy notir2 GND GND efet
M1838 op_jmp notir2 GND GND efet
M1839 GND op_asl_rol n_790 GND efet
M1840 op_T0_bit notir2 GND GND efet
M1841 op_T3_jmp notir2 GND GND efet
M1842 n_513 n_885 GND GND efet
M1843 sb3 dpc0_YSB n_1531 GND efet
M1844 n_1178 pipeUNK30 GND GND efet
M1845 GND irline3 op_T2_pha GND efet
M1846 op_branch_done irline3 GND GND efet
M1847 op_T0_bit irline3 GND GND efet
M1848 adl2 dpc40_ADLPCL pcl2 GND efet
M1849 pcl5 dpc40_ADLPCL adl5 GND efet
M1850 adl0 dpc40_ADLPCL pcl0 GND efet
M1851 noty6 y6 GND GND efet
M1852 adl4 dpc40_ADLPCL pcl4 GND efet
M1853 adl6 dpc40_ADLPCL pcl6 GND efet
M1854 n_783 pcl2 GND GND efet
M1855 dpc11_SBADD n_1247 GND GND efet
M1856 GND irline3 op_T2_stack_access GND efet
M1857 n_233 n_761 n_970 GND efet
M1858 GND irline3 op_T3_jmp GND efet
M1859 n_604 op_T2_stack GND GND efet
M1860 n_1010 pch0 GND GND efet
M1861 GND op_T0_sbc n_605 GND efet
M1862 GND n_1247 dpc1_SBY GND efet
M1863 n_1264 n_453 GND GND efet
M1864 abl7 nABL7 GND GND efet
M1865 db1 n_798 Vdd GND efet
M1866 db1 n_798 Vdd GND efet
M1867 GND adl6 n_1548 GND efet
M1868 n_1225 op_T2_zp_zp_idx GND GND efet
M1869 n_604 notRdy0 GND GND efet
M1870 GND nots3 n_998 GND efet
M1871 GND db0 n_93 GND efet
M1872 n_419 a2 GND GND efet
M1873 GND alua5 n_1559 GND efet
M1874 n_1508 n_46 GND GND efet
M1875 ab15 n_659 GND GND efet
M1876 ab15 n_659 GND GND efet
M1877 n_1546 n_781 GND GND efet
M1878 dpc13_ORS n_1255 GND GND efet
M1879 GND n_897 n_1369 GND efet
M1880 GND n_781 n_1457 GND efet
M1881 op_T3_mem_abs notir3 GND GND efet
M1882 op_T__asl_rol_a notir3 GND GND efet
M1883 x_op_push_pull notir3 GND GND efet
M1884 op_T0_cld_sed notir3 GND GND efet
M1885 n_299 n_1614 n_1616 GND efet
M1886 n_628 n_55 GND GND efet
M1887 n_176 n_10 GND GND efet
M1888 GND dor2 n_224 GND efet
M1889 n_122 n_AxB_6 GND GND efet
M1890 GND VEC0 nVEC GND efet
M1891 GND n_664 n_1697 GND efet
M1892 GND nop_store n_335 GND efet
M1893 GND n_772 n_1305 GND efet
M1894 n_1030 n_AxB_6 GND GND efet
M1895 x1 dpc3_SBX sb1 GND efet
M1896 GND n_1533 n_964 GND efet
M1897 GND op_T2_stack_access n_1090 GND efet
M1898 GND n_1129 n_1467 GND efet
M1899 n_1619 n_1448 GND GND efet
M1900 n_831 cclk a5 GND efet
M1901 n_1598 n_1511 n_262 GND efet
M1902 Pout1 H1x1 idb1 GND efet
M1903 n_1633 n_172 GND GND efet
M1904 n_210 n_172 Vdd GND efet
M1905 n_678 n_1357 GND GND efet
M1906 GND idb3 n_1600 GND efet
M1907 abh3 nABH3 GND GND efet
M1908 GND idb1 DBZ GND efet
M1909 nTWOCYCLE PD_1xx000x0 GND GND efet
M1910 pipeUNK37 cclk n_944 GND efet
M1911 GND op_T0_php_pha n_1464 GND efet
M1912 GND nC34 C34 GND efet
M1913 n_1310 nC34 C45 GND efet
M1914 GND A_B7 n_1617 GND efet
M1915 GND op_T0_cpx_inx n_1106 GND efet
M1916 n_1684 cp1 notdor6 GND efet
M1917 GND n_1081 n_605 GND efet
M1918 db1 GND GND GND efet
M1919 Vdd n_424 notRdy0 GND efet
M1920 GND pipeUNK01 n_1198 GND efet
M1921 n_1692 n_253 GND GND efet
M1922 n_279 n_253 GND GND efet
M1923 n_906 n_1333 GND GND efet
M1924 Vdd n_1129 cclk GND efet
M1925 notRdy0 n_198 GND GND efet
M1926 GND pipeUNK31 n_1178 GND efet
M1927 op_T0_clc_sec ir2 GND GND efet
M1928 op_T0_cli_sei ir2 GND GND efet
M1929 op_push_pull ir2 GND GND efet
M1930 op_jsr ir2 GND GND efet
M1931 op_T2_php ir2 GND GND efet
M1932 op_T4_brk ir2 GND GND efet
M1933 op_T5_rti_rts ir2 GND GND efet
M1934 op_T2_php_pha ir2 GND GND efet
M1935 x_op_T3_plp_pla ir2 GND GND efet
M1936 xx_op_T5_jsr ir2 GND GND efet
M1937 GND n_1599 n_538 GND efet
M1938 GND notRdy0 fetch GND efet
M1939 notir5 ir5 GND GND efet
M1940 GND DA_C45 n_570 GND efet
M1941 GND n_1719 n_831 GND efet
M1942 Vdd n_224 n_37 GND efet
M1943 GND n_224 n_520 GND efet
M1944 n_436 dpc2_XSB sb4 GND efet
M1945 GND irq n_1599 GND efet
M1946 Vdd n_1296 ab11 GND efet
M1947 op_T2_branch notir4 GND GND efet
M1948 op_branch_done notir4 GND GND efet
M1949 op_T5_ind_y notir4 GND GND efet
M1950 op_T4_abs_idx notir4 GND GND efet
M1951 op_T0_tya notir4 GND GND efet
M1952 x_op_T3_ind_y notir4 GND GND efet
M1953 GND notir4 op_T3_abs_idx GND efet
M1954 op_T2_ind_y notir4 GND GND efet
M1955 x_op_T3_abs_idx notir4 GND GND efet
M1956 GND notir4 x_op_T4_ind_y GND efet
M1957 pipenT0 cclk n_17 GND efet
M1958 GND pipeT5out n_1615 GND efet
M1959 GND clock2 op_T__cpx_cpy_abs GND efet
M1960 GND clock2 op_T__asl_rol_a GND efet
M1961 GND n_604 n_385 GND efet
M1962 op_ORS n_1145 GND GND efet
M1963 GND n_609 n_1213 GND efet
M1964 n_1325 dor0 Vdd GND efet
M1965 GND clock2 op_T__ora_and_eor_adc GND efet
M1966 GND clock2 op_T__adc_sbc GND efet
M1967 GND clock2 op_T__inx GND efet
M1968 GND clock2 op_T__iny_dey GND efet
M1969 x_op_T__adc_sbc clock2 GND GND efet
M1970 GND clock2 op_T__cmp GND efet
M1971 op_T__shift_a clock2 GND GND efet
M1972 GND clock2 op_T__bit GND efet
M1973 GND cclk dpc10_ADLADD GND efet
M1974 GND cclk dpc11_SBADD GND efet
M1975 GND cclk dpc12_0ADD GND efet
M1976 op_T2_mem_zp notir2 GND GND efet
M1977 dpc6_SBS cclk GND GND efet
M1978 GND cclk dpc7_SS GND efet
M1979 GND cclk dpc8_nDBADD GND efet
M1980 GND cclk dpc9_DBADD GND efet
M1981 nTWOCYCLE cp1 nTWOCYCLE_phi1 GND efet
M1982 GND dpc12_0ADD alua0 GND efet
M1983 GND n_747 n_1417 GND efet
M1984 naluresult1 cclk notalu1 GND efet
M1985 n_1137 n_790 n_816 GND efet
M1986 n_1254 cclk nABL6 GND efet
M1987 n_180 notRdy0 GND GND efet
M1988 GND n_1202 n_1367 GND efet
M1989 pipeUNK32 cclk n_1081 GND efet
M1990 n_1199 cclk notidl2 GND efet
M1991 n_824 cclk pipeUNK34 GND efet
M1992 n_1154 notRdy0 GND GND efet
M1993 GND n_310 ir0 GND efet
M1994 pipeUNK31 cclk n_389 GND efet
M1995 adh6 cclk Vdd GND efet
M1996 Vdd cclk adl7 GND efet
M1997 n_501 n_180 GND GND efet
M1998 pclp1 npclp1 GND GND efet
M1999 n_239 nop_branch_done n_192 GND efet
M2000 GND noty3 n_1531 GND efet
M2001 op_clv ir6 GND GND efet
M2002 n_473 cclk pipeUNK33 GND efet
M2003 nA_B5 alub5 n_1559 GND efet
M2004 GND alub5 n_A_B_5 GND efet
M2005 Vdd n_1369 dpc38_PCLADL GND efet
M2006 GND nop_store n_816 GND efet
M2007 n_721 dpc4_SSB sb7 GND efet
M2008 n_618 dpc4_SSB sb6 GND efet
M2009 n_1043 n_818 GND GND efet
M2010 Vdd n_818 dpc40_ADLPCL GND efet
M2011 n_3 dpc4_SSB sb4 GND efet
M2012 n_1426 n_270 GND GND efet
M2013 n_210 abl5 GND GND efet
M2014 notRnWprepad cp1 n_759 GND efet
M2015 n_1633 abl5 Vdd GND efet
M2016 op_T2_php_pha notir3 GND GND efet
M2017 GND cclk nDBE GND efet
M2018 op_T0_jmp notir3 GND GND efet
M2019 GND notir3 op_T2_abs_access GND efet
M2020 op_T0_shift_right_a notir3 GND GND efet
M2021 op_T2_pha notir3 GND GND efet
M2022 GND notir3 op_push_pull GND efet
M2023 x_op_jmp notir3 GND GND efet
M2024 x_op_T3_abs_idx notir3 GND GND efet
M2025 op_T3_abs_idx_ind notir3 GND GND efet
M2026 GND alua0 n_A_B_0 GND efet
M2027 n_696 n_0_ADL0 GND GND efet
M2028 naluresult3 cclk notalu3 GND efet
M2029 GND C12 _AxB_2_nC12 GND efet
M2030 n_1641 cp1 n_237 GND efet
M2031 GND n_1635 dpc29_0ADH17 GND efet
M2032 n_1426 n_1662 n_845 GND efet
M2033 n_724 cp1 n_409 GND efet
M2034 n_387 n_206 n_916 GND efet
M2035 GND n_267 n_80 GND efet
M2036 n_AxBxC_2 C12 n_1572 GND efet
M2037 n_A_B_3 dpc13_ORS naluresult3 GND efet
M2038 n_169 n_1624 GND GND efet
M2039 n_36 n_600 GND GND efet
M2040 Vdd n_1325 db0 GND efet
M2041 GND n_319 n_972 GND efet
M2042 GND n_936 AxB1 GND efet
M2043 GND op_branch_done nop_branch_done GND efet
M2044 n_1636 cp1 n_935 GND efet
M2045 GND n_612 db5 GND efet
M2046 GND n_612 db5 GND efet
M2047 GND n_612 db5 GND efet
M2048 n_1724 notx6 GND GND efet
M2049 GND n_612 db5 GND efet
M2050 db5 n_612 GND GND efet
M2051 db5 n_612 GND GND efet
M2052 GND n_612 db5 GND efet
M2053 GND n_445 n_417 GND efet
M2054 GND n_445 n_317 GND efet
M2055 GND noty5 n_733 GND efet
M2056 nABL1 cclk n_66 GND efet
M2057 n_475 abh4 Vdd GND efet
M2058 GND abh4 n_1677 GND efet
M2059 GND abh4 n_999 GND efet
M2060 naluresult0 cclk notalu0 GND efet
M2061 nC01 C01 GND GND efet
M2062 n_1510 C01 nC12 GND efet
M2063 GND n_1447 n_1175 GND efet
M2064 C78 nC78 GND GND efet
M2065 naluresult4 cclk notalu4 GND efet
M2066 n_1407 n_1262 n_933 GND efet
M2067 dpc35_PCHC n_1010 GND GND efet
M2068 n_311 n_1010 GND GND efet
M2069 n_35 n_796 GND GND efet
M2070 GND n_1047 dpc23_SBAC GND efet
M2071 n_340 cclk pipeUNK12 GND efet
M2072 n_254 cp1 n_1353 GND efet
M2073 short_circuit_branch_add n_1446 n_206 GND efet
M2074 n_433 nA_B2 C23 GND efet
M2075 GND n_383 n_1040 GND efet
M2076 n_1040 n_383 GND GND efet
M2077 GND alu2 nDA_ADD2 GND efet
M2078 n_1445 n_270 n_1495 GND efet
M2079 GND n_1593 n_1552 GND efet
M2080 GND pcl3 n_249 GND efet
M2081 n_AxB_0 dpc16_EORS naluresult0 GND efet
M2082 naluresult1 dpc16_EORS n_AxB_1 GND efet
M2083 n_AxB_2 dpc16_EORS naluresult2 GND efet
M2084 n_AxB_3 dpc16_EORS naluresult3 GND efet
M2085 GND n_1202 n_57 GND efet
M2086 GND n_307 n_620 GND efet
M2087 GND n_902 n_1109 GND efet
M2088 GND n_902 n_1109 GND efet
M2089 n_43 cp1 GND GND efet
M2090 GND cp1 n_1247 GND efet
M2091 GND npchp1 pchp1 GND efet
M2092 n_172 abl5 GND GND efet
M2093 n_1687 idb0 GND GND efet
M2094 n_1618 n_419 GND GND efet
M2095 GND n_541 ir7 GND efet
M2096 alu1 dpc20_ADDSB06 sb1 GND efet
M2097 n_587 pipeUNK12 GND GND efet
M2098 alu0 dpc20_ADDSB06 sb0 GND efet
M2099 n_1716 n_510 GND GND efet
M2100 n_AxB_2 A_B2 n_716 GND efet
M2101 n_674 n_25 GND GND efet
M2102 n_1675 cclk notir6 GND efet
M2103 pd3 cclk n_1281 GND efet
M2104 n_1588 cclk pd5 GND efet
M2105 n_929 cclk a1 GND efet
M2106 pd4 cclk n_1075 GND efet
M2107 n_1638 cclk notidl6 GND efet
M2108 GND n_688 n_1223 GND efet
M2109 GND nots0 n_332 GND efet
M2110 GND dpc29_0ADH17 adh2 GND efet
M2111 n_550 op_ANDS GND GND efet
M2112 Vdd cclk adh3 GND efet
M2113 n_1004 n_1408 GND GND efet
M2114 n_1347 n_862 GND GND efet
M2115 n_1604 op_sty_cpy_mem GND GND efet
M2116 GND n_1380 n_109 GND efet
M2117 n_972 n_1610 DC34 GND efet
M2118 n_653 cp1 n_1497 GND efet
M2119 GND op_T0_ora n_1145 GND efet
M2120 dor1 notdor1 GND GND efet
M2121 alua3 dpc12_0ADD GND GND efet
M2122 GND pd7_clearIR PD_0xx0xx0x GND efet
M2123 n_1346 abh3 GND GND efet
M2124 n_359 abh3 GND GND efet
M2125 abh7 nABH7 GND GND efet
M2126 GND n_467 n_10 GND efet
M2127 n_AxB_5 AxB5 GND GND efet
M2128 GND n_1018 n_100 GND efet
M2129 GND x_op_T3_plp_pla n_368 GND efet
M2130 GND n_231 ONEBYTE GND efet
M2131 n_911 n_877 GND GND efet
M2132 n_911 n_877 GND GND efet
M2133 GND n_133 n_602 GND efet
M2134 GND n_300 n_847 GND efet
M2135 dpc18_nDAA n_709 GND GND efet
M2136 Vdd n_133 dpc2_XSB GND efet
M2137 n_1254 abl6 GND GND efet
M2138 n_1195 abl6 GND GND efet
M2139 Vdd abl6 n_1191 GND efet
M2140 ab3 n_1041 Vdd GND efet
M2141 Vdd n_1041 ab3 GND efet
M2142 Vdd n_1041 ab3 GND efet
M2143 Vdd n_1041 ab3 GND efet
M2144 GND notir6 op_T__dex GND efet
M2145 op_T0_cpx_inx notir6 GND GND efet
M2146 GND notir6 op_T4_rts GND efet
M2147 GND notir6 op_T__inx GND efet
M2148 n_616 cclk n_460 GND efet
M2149 Vdd n_628 dpc24_ACSB GND efet
M2150 GND notir6 op_T0_dex GND efet
M2151 GND notir6 op_T0_cpy_iny GND efet
M2152 op_ror notir6 GND GND efet
M2153 GND notir6 op_T5_rti GND efet
M2154 GND n_1602 n_1596 GND efet
M2155 n_735 n_320 GND GND efet
M2156 adl2 dpc41_DL_ADL n_1424 GND efet
M2157 adl4 dpc41_DL_ADL n_1095 GND efet
M2158 GND RnWstretched n_471 GND efet
M2159 GND n_770 n_19 GND efet
M2160 sb1 cclk Vdd GND efet
M2161 GND notidl7 idl7 GND efet
M2162 GND notidl7 idl7 GND efet
M2163 n_182 n_236 n_1151 GND efet
M2164 n_1161 cp1 n_109 GND efet
M2165 n_564 dpc0_YSB sb0 GND efet
M2166 n_388 AxB1 GND GND efet
M2167 alu2 dpc21_ADDADL adl2 GND efet
M2168 adl0 dpc21_ADDADL alu0 GND efet
M2169 adl1 dpc21_ADDADL alu1 GND efet
M2170 GND Reset0 n_501 GND efet
M2171 GND op_T5_rti n_1464 GND efet
M2172 n_261 x_op_T3_abs_idx GND GND efet
M2173 op_T3_ind_x ir2 GND GND efet
M2174 op_T4_rti ir2 GND GND efet
M2175 op_T5_rti ir2 GND GND efet
M2176 op_T3_plp_pla ir2 GND GND efet
M2177 op_T4_brk_jsr ir2 GND GND efet
M2178 op_T5_brk ir2 GND GND efet
M2179 op_T0_jsr ir2 GND GND efet
M2180 op_T4_rts ir2 GND GND efet
M2181 op_T0_php_pha ir2 GND GND efet
M2182 GND VEC1 nVEC GND efet
M2183 n_728 cclk pipeVectorA0 GND efet
M2184 n_381 abh0 GND GND efet
M2185 pipeUNK13 cclk n_1045 GND efet
M2186 n_1177 cclk n_1069 GND efet
M2187 n_1315 abh0 GND GND efet
M2188 dpc34_PCLC n_232 GND GND efet
M2189 GND n_232 n_1316 GND efet
M2190 dpc0_YSB n_969 GND GND efet
M2191 GND n_232 n_585 GND efet
M2192 AxB5 n_A_B_5 GND GND efet
M2193 A_B5 n_A_B_5 GND GND efet
M2194 Pout0 n_31 GND GND efet
M2195 GND ONEBYTE n_1275 GND efet
M2196 GND notRdy0 n_191 GND efet
M2197 op_T__asl_rol_a notir1 GND GND efet
M2198 Reset0 cclk pipephi2Reset0x GND efet
M2199 ab9 n_1140 Vdd GND efet
M2200 op_SUMS op_ANDS GND GND efet
M2201 Vdd dor3 n_42 GND efet
M2202 GND ir6 op_jsr GND efet
M2203 GND ir6 op_store GND efet
M2204 n_1254 n_1195 Vdd GND efet
M2205 n_1055 n_771 GND GND efet
M2206 GND n_726 n_630 GND efet
M2207 GND n_1195 n_1191 GND efet
M2208 n_721 nots7 GND GND efet
M2209 n_1225 cclk pipedpc28 GND efet
M2210 GND n_43 n_1534 GND efet
M2211 n_1330 nnT2BR GND GND efet
M2212 ab14 n_635 GND GND efet
M2213 ab14 n_635 GND GND efet
M2214 dor7 notdor7 GND GND efet
M2215 GND pipeT4out n_1703 GND efet
M2216 GND op_EORS op_SUMS GND efet
M2217 GND n_1315 n_826 GND efet
M2218 GND nNMIP NMIP GND efet
M2219 GND n_556 n_1344 GND efet
M2220 n_733 cclk y5 GND efet
M2221 Vdd n_1639 ab15 GND efet
M2222 n_1202 n_1265 GND GND efet
M2223 dpc35_PCHC n_1265 GND GND efet
M2224 n_1590 fetch n_1620 GND efet
M2225 n_463 cp1 n_1094 GND efet
M2226 n_1467 n_358 Vdd GND efet
M2227 GND RnWstretched n_769 GND efet
M2228 GND RnWstretched n_1325 GND efet
M2229 GND RnWstretched n_1325 GND efet
M2230 db6 n_471 GND GND efet
M2231 GND n_471 db6 GND efet
M2232 GND notRdy0 n_1275 GND efet
M2233 GND n_645 n_1368 GND efet
M2234 n_1586 cclk n_621 GND efet
M2235 GND xx_op_T5_jsr n_368 GND efet
M2236 n_316 alua0 GND GND efet
M2237 GND n_519 n_670 GND efet
M2238 pclp3 dpc37_PCLDB idb3 GND efet
M2239 pclp1 dpc37_PCLDB idb1 GND efet
M2240 GND irline3 op_T2_stack GND efet
M2241 GND irline3 op_T3_stack_bit_jmp GND efet
M2242 nA_B1 dpc15_ANDS naluresult1 GND efet
M2243 op_T4_rti irline3 GND GND efet
M2244 op_plp_pla irline3 GND GND efet
M2245 GND nABL4 abl4 GND efet
M2246 n_1595 n_754 GND GND efet
M2247 n_648 n_754 n_1181 GND efet
M2248 Vdd n_1545 ab10 GND efet
M2249 nots1 cclk n_1711 GND efet
M2250 n_139 op_SRS GND GND efet
M2251 nop_store op_store GND GND efet
M2252 n_506 n_192 GND GND efet
M2253 adh0 dpc28_0ADH0 GND GND efet
M2254 rw n_1696 GND GND efet
M2255 GND n_1696 rw GND efet
M2256 dpc38_PCLADL n_1462 GND GND efet
M2257 BRtaken n_1115 GND GND efet
M2258 n_935 adl2 GND GND efet
M2259 GND n_5 n_146 GND efet
M2260 GND n_260 dasb7 GND efet
M2261 dasb1 n_735 GND GND efet
M2262 GND n_1467 cclk GND efet
M2263 GND pipeUNK34 n_720 GND efet
M2264 GND notir5 op_T0_cpx_inx GND efet
M2265 GND notir5 op_T0_ldx_tax_tsx GND efet
M2266 nABH5 cclk n_869 GND efet
M2267 idb7 dpc33_PCHDB pchp7 GND efet
M2268 pchp4 dpc33_PCHDB idb4 GND efet
M2269 pchp3 dpc33_PCHDB idb3 GND efet
M2270 idb6 dpc33_PCHDB pchp6 GND efet
M2271 pchp5 dpc33_PCHDB idb5 GND efet
M2272 pchp0 dpc33_PCHDB idb0 GND efet
M2273 n_1279 n_986 n_345 GND efet
M2274 idb2 dpc33_PCHDB pchp2 GND efet
M2275 idb1 dpc33_PCHDB pchp1 GND efet
M2276 n_1358 cclk n_521 GND efet
M2277 GND n_318 Pout1 GND efet
M2278 n_AxBxC_2 _AxB_2_nC12 GND GND efet
M2279 abh6 nABH6 GND GND efet
M2280 Vdd n_466 n_471 GND efet
M2281 n_384 n_1258 GND GND efet
M2282 npclp5 cclk n_1073 GND efet
M2283 GND n_466 n_7 GND efet
M2284 GND C1x5Reset n_1712 GND efet
M2285 n_661 n_1170 n_566 GND efet
M2286 Vdd n_1633 ab5 GND efet
M2287 GND n_506 n_877 GND efet
M2288 C01 nA_B0 n_942 GND efet
M2289 GND pd3_clearIR n_1083 GND efet
M2290 PD_1xx000x0 pd3_clearIR GND GND efet
M2291 n_1480 n_1472 GND GND efet
M2292 n_747 n_670 GND GND efet
M2293 GND adh6 n_880 GND efet
M2294 s7 dpc7_SS n_721 GND efet
M2295 naluresult6 dpc13_ORS n_A_B_6 GND efet
M2296 n_1278 n_824 n_1642 GND efet
M2297 Vdd n_373 db5 GND efet
M2298 GND n_1175 n_267 GND efet
M2299 n_1014 cp1 idl6 GND efet
M2300 n_1546 n_1600 n_1495 GND efet
M2301 Vdd cclk adl2 GND efet
M2302 n_1402 cclk npchp2 GND efet
M2303 clock2 n_1533 GND GND efet
M2304 Vdd n_373 db5 GND efet
M2305 n_1044 n_31 GND GND efet
M2306 GND n_905 n_979 GND efet
M2307 naluresult5 dpc15_ANDS nA_B5 GND efet
M2308 n_1121 cclk n_1225 GND efet
M2309 ab8 n_381 GND GND efet
M2310 GND n_152 n_1343 GND efet
M2311 ab8 n_381 GND GND efet
M2312 GND n_381 ab8 GND efet
M2313 ab8 n_381 GND GND efet
M2314 GND n_381 ab8 GND efet
M2315 GND n_783 dpc34_PCLC GND efet
M2316 GND n_783 n_1253 GND efet
M2317 ab8 n_381 GND GND efet
M2318 ab8 n_381 GND GND efet
M2319 op_T0_shift_right_a ir2 GND GND efet
M2320 op_T2_pha ir2 GND GND efet
M2321 op_T0_tay ir2 GND GND efet
M2322 op_T0_pla ir2 GND GND efet
M2323 op_T0_txa ir2 GND GND efet
M2324 op_T__shift_a ir2 GND GND efet
M2325 op_branch_done ir2 GND GND efet
M2326 op_T5_ind_y ir2 GND GND efet
M2327 op_T0_tax ir2 GND GND efet
M2328 op_T0_shift_a ir2 GND GND efet
M2329 adh5 dpc27_SBADH sb5 GND efet
M2330 pcl2 dpc39_PCLPCL pclp2 GND efet
M2331 GND adh5 n_254 GND efet
M2332 n_618 dpc5_SADL adl6 GND efet
M2333 n_515 n_1542 n_1158 GND efet
M2334 GND nA_B6 n_1038 GND efet
M2335 dpc12_0ADD n_1247 GND GND efet
M2336 GND notidl1 idl1 GND efet
M2337 GND notidl1 idl1 GND efet
M2338 GND n_847 n_104 GND efet
M2339 n_1257 notalucout GND GND efet
M2340 naluresult5 cclk notalu5 GND efet
M2341 n_911 n_79 n_696 GND efet
M2342 DBZ idb4 GND GND efet
M2343 n_1152 abl2 Vdd GND efet
M2344 n_951 abl2 GND GND efet
M2345 n_642 abl2 GND GND efet
M2346 GND n_676 ab9 GND efet
M2347 ab9 n_676 GND GND efet
M2348 GND idb6 n_351 GND efet
M2349 n_AxB_7 AxB7 GND GND efet
M2350 n_1392 nmi GND GND efet
M2351 n_1699 cclk n_1024 GND efet
M2352 pipeT3out cclk n_678 GND efet
M2353 GND pipeUNK22 n_533 GND efet
M2354 GND n_AxB_4 n_375 GND efet
M2355 GND n_AxB_4 _AxB_4_nC34 GND efet
M2356 n_869 n_1423 Vdd GND efet
M2357 n_168 cp1 n_836 GND efet
M2358 GND n_410 n_474 GND efet
M2359 GND n_1423 n_1608 GND efet
M2360 nop_set_C cclk pipeUNK08 GND efet
M2361 notRnWprepad cp1 n_1579 GND efet
M2362 p1 cp1 n_566 GND efet
M2363 dpc3_SBX n_1247 GND GND efet
M2364 n_306 cclk n_581 GND efet
M2365 dpc41_DL_ADL n_1157 GND GND efet
M2366 GND n_562 NMIL GND efet
M2367 dor5 notdor5 GND GND efet
M2368 ab15 n_1639 Vdd GND efet
M2369 DBZ idb2 GND GND efet
M2370 op_rol_ror ir6 GND GND efet
M2371 op_sty_cpy_mem ir6 GND GND efet
M2372 GND ir6 op_T0_txs GND efet
M2373 op_T0_ldx_tax_tsx ir6 GND GND efet
M2374 GND ir6 x_op_T0_txa GND efet
M2375 GND ir6 op_from_x GND efet
M2376 x_op_T0_txa notir1 GND GND efet
M2377 GND notir1 op_xy GND efet
M2378 op_from_x notir1 GND GND efet
M2379 op_T0_dex notir1 GND GND efet
M2380 op_T0_ldx_tax_tsx notir1 GND GND efet
M2381 op_T0_txs notir1 GND GND efet
M2382 op_T0_tsx notir1 GND GND efet
M2383 GND ir7 op_T2_stack GND efet
M2384 op_inc_nop notir1 GND GND efet
M2385 op_ror notir1 GND GND efet
M2386 n_436 cclk x4 GND efet
M2387 GND pcl7 n_641 GND efet
M2388 GND n_1045 p7 GND efet
M2389 n_588 db7 GND GND efet
M2390 GND n_409 PD_xxx010x1 GND efet
M2391 naluresult6 cclk notalu6 GND efet
M2392 sb0 cclk Vdd GND efet
M2393 GND RnWstretched n_1720 GND efet
M2394 GND RnWstretched n_373 GND efet
M2395 GND RnWstretched n_373 GND efet
M2396 n_559 cclk n_608 GND efet
M2397 GND op_T3_mem_zp_idx n_347 GND efet
M2398 n_1380 n_1154 GND GND efet
M2399 GND pipedpc28 dpc28_0ADH0 GND efet
M2400 n_1365 notRdy0 n_1085 GND efet
M2401 GND op_T5_rti n_256 GND efet
M2402 n_1026 abl7 GND GND efet
M2403 n_251 n_221 GND GND efet
M2404 GND n_255 dpc31_PCHPCH GND efet
M2405 n_457 cp1 notdor3 GND efet
M2406 n_626 cp1 n_756 GND efet
M2407 n_359 cclk nABH3 GND efet
M2408 ab11 n_359 GND GND efet
M2409 n_619 n_700 GND GND efet
M2410 GND notRdy0 n_781 GND efet
M2411 n_1118 n_638 n_604 GND efet
M2412 n_467 n_134 GND GND efet
M2413 n_930 n_134 GND GND efet
M2414 GND notalu3 alu3 GND efet
M2415 GND n_1224 n_186 GND efet
M2416 Vdd n_1277 dpc42_DL_ADH GND efet
M2417 ab3 n_138 GND GND efet
M2418 n_363 pipeT_SYNC GND GND efet
M2419 npclp6 n_993 GND GND efet
M2420 GND n_147 db4 GND efet
M2421 GND n_147 db4 GND efet
M2422 n_1376 idb2 GND GND efet
M2423 GND PD_0xx0xx0x PD_n_0xx0xx0x GND efet
M2424 GND n_147 db4 GND efet
M2425 GND n_147 db4 GND efet
M2426 GND n_147 db4 GND efet
M2427 GND n_147 db4 GND efet
M2428 n_717 n_1132 GND GND efet
M2429 GND n_937 n_1345 GND efet
M2430 GND cclk dpc1_SBY GND efet
M2431 dpc2_XSB cclk GND GND efet
M2432 GND cclk dpc3_SBX GND efet
M2433 n_104 cclk n_1221 GND efet
M2434 GND n_937 dpc34_PCLC GND efet
M2435 GND n_937 n_1706 GND efet
M2436 n_47 cp1 n_420 GND efet
M2437 GND cclk dpc0_YSB GND efet
M2438 GND op_T2_abs_access n_773 GND efet
M2439 GND n_964 n_17 GND efet
M2440 GND n_964 clock1 GND efet
M2441 GND n_663 npchp7 GND efet
M2442 adh2 cclk Vdd GND efet
M2443 n_1085 n_372 n_1172 GND efet
M2444 n_912 notRdy0 n_1290 GND efet
M2445 GND RnWstretched n_466 GND efet
M2446 n_1286 n_470 GND GND efet
M2447 n_135 n_127 GND GND efet
M2448 abh0 nABH0 GND GND efet
M2449 GND ir6 op_T0_plp GND efet
M2450 GND ir6 x_op_T0_bit GND efet
M2451 GND RnWstretched n_298 GND efet
M2452 GND RnWstretched n_23 GND efet
M2453 n_1279 n_600 GND GND efet
M2454 GND n_161 n_969 GND efet
M2455 Vdd n_161 dpc0_YSB GND efet
M2456 n_715 n_641 GND GND efet
M2457 dpc34_PCLC n_641 GND GND efet
M2458 GND n_1247 dpc7_SS GND efet
M2459 GND op_T4_brk_jsr n_604 GND efet
M2460 y5 dpc1_SBY sb5 GND efet
M2461 op_T2_php ir6 GND GND efet
M2462 op_T4_brk ir6 GND GND efet
M2463 n_19 cclk pipeUNK18 GND efet
M2464 adl3 dpc10_ADLADD alub3 GND efet
M2465 n_1286 n_930 GND GND efet
M2466 GND dpc22_nDSA n_1179 GND efet
M2467 db6 GND GND GND efet
M2468 GND db0 n_718 GND efet
M2469 GND db2 n_111 GND efet
M2470 n_1618 cclk a2 GND efet
M2471 n_896 db3 GND GND efet
M2472 naluresult7 cclk notalu7 GND efet
M2473 n_1322 n_320 GND GND efet
M2474 adl0 dpc41_DL_ADL n_719 GND efet
M2475 adl1 dpc41_DL_ADL n_87 GND efet
M2476 n_327 op_T0_plp GND GND efet
M2477 adl3 dpc41_DL_ADL n_1661 GND efet
M2478 GND RnWstretched n_471 GND efet
M2479 n_80 cclk n_1333 GND efet
M2480 n_571 pd2_clearIR GND GND efet
M2481 GND n_916 short_circuit_idx_add GND efet
M2482 GND nnT2BR n_272 GND efet
M2483 GND pd2_clearIR PD_1xx000x0 GND efet
M2484 op_T__inx ir4 GND GND efet
M2485 GND pd2_clearIR PD_xxx010x1 GND efet
M2486 PD_xxxx10x0 pd2_clearIR GND GND efet
M2487 op_T0_dex ir4 GND GND efet
M2488 x_op_T0_txa ir4 GND GND efet
M2489 GND notidl4 idl4 GND efet
M2490 idl4 notidl4 GND GND efet
M2491 op_T0_iny_dey ir4 GND GND efet
M2492 GND n_1070 n_200 GND efet
M2493 op_T2_ind_x ir4 GND GND efet
M2494 op_T0_cpy_iny ir4 GND GND efet
M2495 op_T0_pla clock1 GND GND efet
M2496 op_T0_lda clock1 GND GND efet
M2497 GND clock1 op_T0_acc GND efet
M2498 GND clock1 op_T0_tay GND efet
M2499 GND clock1 op_T0_shift_a GND efet
M2500 GND clock1 op_T0_bit GND efet
M2501 op_T0_and clock1 GND GND efet
M2502 op_branch_done clock1 GND GND efet
M2503 op_T0_shift_right_a clock1 GND GND efet
M2504 GND alua4 n_A_B_4 GND efet
M2505 GND alua4 n_185 GND efet
M2506 GND adl0 n_123 GND efet
M2507 GND n_1272 n_608 GND efet
M2508 n_511 n_553 n_845 GND efet
M2509 npchp4 cclk n_1657 GND efet
M2510 nWR op_T4_brk GND GND efet
M2511 n_1391 op_T4_brk GND GND efet
M2512 alu3 dpc20_ADDSB06 sb3 GND efet
M2513 sb4 dpc20_ADDSB06 alu4 GND efet
M2514 Vdd n_1566 dpc43_DL_DB GND efet
M2515 n_1507 cp1 n_864 GND efet
M2516 n_1455 cclk n_1505 GND efet
M2517 n_1240 n_1566 GND GND efet
M2518 C01 n_A_B_0 GND GND efet
M2519 GND dpc29_0ADH17 adh6 GND efet
M2520 pclp5 dpc37_PCLDB idb5 GND efet
M2521 n_1118 op_T2_ADL_ADD GND GND efet
M2522 n_626 n_1401 n_1198 GND efet
M2523 GND notidl7 idl7 GND efet
M2524 GND npchp3 pchp3 GND efet
M2525 n_1528 cp1 n_1215 GND efet
M2526 n_AxBxC_1 n_AxB1__C01 GND GND efet
M2527 n_51 op_T0_sbc n_29 GND efet
M2528 n_732 n_1161 GND GND efet
M2529 GND op_T3_mem_abs n_347 GND efet
M2530 GND ir7 op_T2_brk GND efet
M2531 op_T3_jsr ir7 GND GND efet
M2532 GND n_1613 n_42 GND efet
M2533 GND ir7 op_T0_shift_right_a GND efet
M2534 n_1267 cp1 n_1298 GND efet
M2535 GND n_1097 dasb3 GND efet
M2536 GND nDA_ADD1 n_1682 GND efet
M2537 GND ir7 op_T0_and GND efet
M2538 Vdd n_1613 n_643 GND efet
M2539 GND ir7 op_T2_pha GND efet
M2540 pipeT5out cclk n_378 GND efet
M2541 op_T0_shift_a ir7 GND GND efet
M2542 GND nDA_ADD1 n_1362 GND efet
M2543 GND ir7 op_T0_bit GND efet
M2544 GND notalu2 alu2 GND efet
M2545 n_1510 A_B1 GND GND efet
M2546 PD_0xx0xx0x pd1_clearIR GND GND efet
M2547 n_AxB5__C45 AxB5 GND GND efet
M2548 n_551 n_393 GND GND efet
M2549 pipeUNK23 cclk n_1085 GND efet
M2550 GND pipeT2out n_12 GND efet
M2551 GND adl1 n_1016 GND efet
M2552 n_1013 nC67 n_AxBxC_7 GND efet
M2553 GND nC67 n_AxB7__C67 GND efet
M2554 n_1175 cclk pipeUNK28 GND efet
M2555 n_1312 n_1291 GND GND efet
M2556 n_1681 op_shift GND GND efet
M2557 n_1270 n_43 GND GND efet
M2558 n_794 dor1 GND GND efet
M2559 n_288 dor1 GND GND efet
M2560 n_1390 C56 n_AxBxC_6 GND efet
M2561 GND C56 _AxB_6_nC56 GND efet
M2562 dpc39_PCLPCL n_1247 GND GND efet
M2563 GND n_119 ir1 GND efet
M2564 _t4 n_188 GND GND efet
M2565 n_782 n_1303 n_1040 GND efet
M2566 op_T0_cpx_inx irline3 GND GND efet
M2567 C45 n_A_B_4 GND GND efet
M2568 op_T__iny_dey irline3 GND GND efet
M2569 op_T__inx irline3 GND GND efet
M2570 GND irline3 op_T0_tay_ldy_not_idx GND efet
M2571 op_T0_ldy_mem irline3 GND GND efet
M2572 GND irline3 op_T5_brk GND efet
M2573 GND irline3 op_T0_jsr GND efet
M2574 op_T4_rts irline3 GND GND efet
M2575 op_T0_php_pha irline3 GND GND efet
M2576 Vdd abh1 n_1140 GND efet
M2577 Vdd n_842 n_66 GND efet
M2578 GND n_1149 nNMIG GND efet
M2579 GND n_1565 n_1218 GND efet
M2580 n_1049 cclk n_160 GND efet
M2581 n_647 nA_B5 GND GND efet
M2582 GND n_1501 db7 GND efet
M2583 db7 n_1501 GND GND efet
M2584 db7 n_1501 GND GND efet
M2585 db7 n_1501 GND GND efet
M2586 pipeUNK27 cclk op_SRS GND efet
M2587 GND RnWstretched n_7 GND efet
M2588 n_1092 nNMIG n_480 GND efet
M2589 n_632 op_T2_stack GND GND efet
M2590 n_794 RnWstretched GND GND efet
M2591 GND n_593 dpc4_SSB GND efet
M2592 alua0 dpc11_SBADD sb0 GND efet
M2593 n_613 n_600 n_1362 GND efet
M2594 alua5 dpc11_SBADD sb5 GND efet
M2595 alua6 dpc11_SBADD sb6 GND efet
M2596 GND pch4 n_1400 GND efet
M2597 op_T2_abs_y ir2 GND GND efet
M2598 op_T3_ind_y ir2 GND GND efet
M2599 n_645 NMIP GND GND efet
M2600 GND n_865 n_420 GND efet
M2601 GND noty7 n_1251 GND efet
M2602 GND pch2 n_1265 GND efet
M2603 a4 cclk n_1344 GND efet
M2604 n_388 n_936 GND GND efet
M2605 n_1707 n_936 GND GND efet
M2606 GND alua6 n_A_B_6 GND efet
M2607 adh0 cclk Vdd GND efet
M2608 n_455 n_279 GND GND efet
M2609 GND s6 n_1187 GND efet
M2610 GND op_jmp n_1649 GND efet
M2611 GND pd7_clearIR n_1605 GND efet
M2612 n_719 cp1 idl0 GND efet
M2613 GND op_T4_mem_abs_idx n_347 GND efet
M2614 GND nABL6 abl6 GND efet
M2615 GND n_1413 dpc32_PCHADH GND efet
M2616 n_553 n_781 GND GND efet
M2617 n_1280 op_sta_cmp n_1037 GND efet
M2618 dpc6_SBS n_6 Vdd GND efet
M2619 GND n_6 n_282 GND efet
M2620 GND op_T0_and n_669 GND efet
M2621 GND n_678 _t3 GND efet
M2622 notx6 x6 GND GND efet
M2623 GND idb1 n_583 GND efet
M2624 n_35 n_43 GND GND efet
M2625 pd0 cclk n_93 GND efet
M2626 pd1 cclk n_1319 GND efet
M2627 GND n_636 nnT2BR GND efet
M2628 ab0 n_855 Vdd GND efet
M2629 op_T3_jmp ir4 GND GND efet
M2630 op_T0_cpx_cpy_inx_iny ir4 GND GND efet
M2631 adh6 dpc32_PCHADH pchp6 GND efet
M2632 adh5 dpc32_PCHADH pchp5 GND efet
M2633 n_6 n_43 GND GND efet
M2634 adh7 dpc32_PCHADH pchp7 GND efet
M2635 n_43 n_839 Vdd GND efet
M2636 n_484 cclk npclp7 GND efet
M2637 n_1215 short_circuit_idx_add GND GND efet
M2638 GND adl3 n_1507 GND efet
M2639 n_930 n_1276 GND GND efet
M2640 GND n_1400 n_83 GND efet
M2641 op_EORS cclk n_982 GND efet
M2642 GND clock1 op_T0_ldy_mem GND efet
M2643 GND clock1 op_T0_jsr GND efet
M2644 op_T0_ldx_tax_tsx clock1 GND GND efet
M2645 GND clock1 op_T0_tsx GND efet
M2646 op_T0_cpx_inx clock1 GND GND efet
M2647 op_T0_txs clock1 GND GND efet
M2648 GND clock1 x_op_T0_txa GND efet
M2649 GND clock1 op_T0_dex GND efet
M2650 GND clock1 op_T0_iny_dey GND efet
M2651 GND clock1 x_op_T0_tya GND efet
M2652 GND op_rti_rts n_1649 GND efet
M2653 Vdd n_102 rw GND efet
M2654 Vdd n_102 rw GND efet
M2655 db3 n_643 GND GND efet
M2656 db3 n_643 GND GND efet
M2657 GND n_643 db3 GND efet
M2658 GND n_643 db3 GND efet
M2659 Vdd n_102 rw GND efet
M2660 Vdd n_102 rw GND efet
M2661 Vdd n_102 rw GND efet
M2662 Vdd n_102 rw GND efet
M2663 db2 n_37 GND GND efet
M2664 db2 n_37 GND GND efet
M2665 GND n_37 db2 GND efet
M2666 db2 n_37 GND GND efet
M2667 db2 n_37 GND GND efet
M2668 db2 n_37 GND GND efet
M2669 n_36 n_8 GND GND efet
M2670 GND n_37 db2 GND efet
M2671 n_1030 n_570 DC78 GND efet
M2672 n_150 n_8 GND GND efet
M2673 GND notir7 op_T__iny_dey GND efet
M2674 GND notir7 op_T0_tsx GND efet
M2675 n_1101 cclk n_190 GND efet
M2676 noty1 y1 GND GND efet
M2677 n_501 n_819 GND GND efet
M2678 n_972 n_A_B_2 GND GND efet
M2679 n_1470 n_1111 GND GND efet
M2680 GND cclk n_628 GND efet
M2681 n_313 alua3 GND GND efet
M2682 GND n_1111 n_1614 GND efet
M2683 GND RnWstretched n_798 GND efet
M2684 GND RnWstretched n_798 GND efet
M2685 GND cclk n_525 GND efet
M2686 GND RnWstretched n_288 GND efet
M2687 n_A_B_3 alua3 GND GND efet
M2688 Vdd n_1191 ab6 GND efet
M2689 n_806 GND GND GND efet
M2690 nABH2 cclk n_994 GND efet
M2691 n_1205 n_233 n_569 GND efet
M2692 Vdd n_1499 dpc18_nDAA GND efet
M2693 n_1386 n_1316 n_426 GND efet
M2694 n_1229 cclk npchp0 GND efet
M2695 Vdd n_1191 ab6 GND efet
M2696 op_T2_stack ir2 GND GND efet
M2697 GND n_646 n_773 GND efet
M2698 Vdd n_1720 n_612 GND efet
M2699 n_1076 dor4 Vdd GND efet
M2700 n_405 BRtaken n_1172 GND efet
M2701 GND n_1720 n_373 GND efet
M2702 notir3 ir3 GND GND efet
M2703 n_1609 cclk notir5 GND efet
M2704 op_T__bit irline3 GND GND efet
M2705 op_T0_clc_sec irline3 GND GND efet
M2706 x_op_T0_bit irline3 GND GND efet
M2707 GND irline3 op_T0_plp GND efet
M2708 GND irline3 x_op_T4_rti GND efet
M2709 GND irline3 op_T__cpx_cpy_abs GND efet
M2710 x_op_push_pull irline3 GND GND efet
M2711 op_T0_cld_sed irline3 GND GND efet
M2712 op_clv irline3 GND GND efet
M2713 n_995 n_312 GND GND efet
M2714 n_A_B_0 dpc13_ORS naluresult0 GND efet
M2715 GND n_947 n_1654 GND efet
M2716 GND n_933 n_877 GND efet
M2717 n_1657 n_523 n_1406 GND efet
M2718 n_875 n_523 n_1659 GND efet
M2719 GND n_523 n_743 GND efet
M2720 GND op_T__bit n_513 GND efet
M2721 n_708 n_1230 GND GND efet
M2722 Vdd n_1230 dpc11_SBADD GND efet
M2723 naluresult7 dpc13_ORS n_A_B_7 GND efet
M2724 pipeUNK01 cclk n_1110 GND efet
M2725 Vdd n_21 dpc30_ADHPCH GND efet
M2726 n_228 n_21 GND GND efet
M2727 DC78 dpc18_nDAA GND GND efet
M2728 dpc20_ADDSB06 n_75 GND GND efet
M2729 Vdd n_834 n_102 GND efet
M2730 n_661 pipeUNK14 GND GND efet
M2731 alu7 notalu7 GND GND efet
M2732 GND dor0 n_1072 GND efet
M2733 op_T0_tay irline3 GND GND efet
M2734 GND n_755 n_1170 GND efet
M2735 GND dor0 n_769 GND efet
M2736 GND n_761 n_762 GND efet
M2737 GND irline3 op_T5_jsr GND efet
M2738 GND nop_branch_bit6 n_1293 GND efet
M2739 op_T0_cpx_cpy_inx_iny irline3 GND GND efet
M2740 GND nots1 n_694 GND efet
M2741 GND n_321 n_849 GND efet
M2742 n_533 cp1 n_599 GND efet
M2743 n_1145 notRdy0 GND GND efet
M2744 GND ir7 notir7 GND efet
M2745 GND n_1304 n_1688 GND efet
M2746 GND dpc18_nDAA DC34 GND efet
M2747 GND notir0 op_T3_ind_x GND efet
M2748 y6 dpc1_SBY sb6 GND efet
M2749 n_920 cp1 n_785 GND efet
M2750 GND clearIR pd0_clearIR GND efet
M2751 pd5_clearIR clearIR GND GND efet
M2752 clk2out n_127 Vdd GND efet
M2753 y4 dpc1_SBY sb4 GND efet
M2754 n_748 nA_B7 GND GND efet
M2755 naluresult7 dpc14_SRS Vdd GND efet
M2756 GND op_lsr_ror_dec_inc n_790 GND efet
M2757 GND n_763 dpc8_nDBADD GND efet
M2758 op_T2_brk ir4 GND GND efet
M2759 op_T0_shift_right_a ir4 GND GND efet
M2760 op_T5_rts ir4 GND GND efet
M2761 op_T3_jsr ir4 GND GND efet
M2762 op_T0_jmp ir4 GND GND efet
M2763 op_T0_brk_rti ir4 GND GND efet
M2764 op_brk_rti ir4 GND GND efet
M2765 op_T5_ind_x ir4 GND GND efet
M2766 x_op_jmp ir4 GND GND efet
M2767 op_jsr ir4 GND GND efet
M2768 n_300 n_389 GND GND efet
M2769 GND n_1541 n_491 GND efet
M2770 GND notir0 op_T0_cmp GND efet
M2771 op_T4_brk_jsr ir3 GND GND efet
M2772 op_T4_rti ir3 GND GND efet
M2773 op_T5_rti ir3 GND GND efet
M2774 op_T2_ADL_ADD ir3 GND GND efet
M2775 op_T2_ind_y ir3 GND GND efet
M2776 op_T4_ind_x ir3 GND GND efet
M2777 op_T3_ind_x ir3 GND GND efet
M2778 op_T4_ind_y ir3 GND GND efet
M2779 x_op_T3_ind_y ir3 GND GND efet
M2780 op_rti_rts ir3 GND GND efet
M2781 GND notir5 op_T4_rts GND efet
M2782 GND RnWstretched n_147 GND efet
M2783 GND op_T5_mem_ind_idx n_347 GND efet
M2784 GND idb2 n_458 GND efet
M2785 pchp4 npchp4 GND GND efet
M2786 n_917 n_383 GND GND efet
M2787 GND pcl5 n_386 GND efet
M2788 n_1649 notRdy0 GND GND efet
M2789 n_472 n_16 n_1366 GND efet
M2790 GND pipeUNK18 n_850 GND efet
M2791 GND RnWstretched n_147 GND efet
M2792 n_1656 n_613 dasb2 GND efet
M2793 Vdd cclk idb7 GND efet
M2794 VEC1 cclk n_1452 GND efet
M2795 GND C78_phi2 notalucout GND efet
M2796 GND n_1137 short_circuit_idx_add GND efet
M2797 n_46 notRdy0 GND GND efet
M2798 n_643 RnWstretched GND GND efet
M2799 GND n_1716 n_180 GND efet
M2800 n_896 cclk notidl3 GND efet
M2801 n_AxBxC_3 n_AxB3__C23 GND GND efet
M2802 op_T0_and ir6 GND GND efet
M2803 op_T2_brk ir6 GND GND efet
M2804 GND ir6 op_T3_jsr GND efet
M2805 GND ir6 op_sta_cmp GND efet
M2806 GND ir6 op_T0_lda GND efet
M2807 GND ir6 op_T0_tay GND efet
M2808 op_T0_tax ir6 GND GND efet
M2809 op_T0_bit ir6 GND GND efet
M2810 n_462 n_1338 GND GND efet
M2811 INTG brk_done GND GND efet
M2812 Vdd n_7 db6 GND efet
M2813 Vdd n_7 db6 GND efet
M2814 GND pd1_clearIR n_1641 GND efet
M2815 GND n_680 n_1526 GND efet
M2816 n_1205 n_811 n_100 GND efet
M2817 idb1 cclk Vdd GND efet
M2818 nA_B7 alub7 n_1695 GND efet
M2819 dpc42_DL_ADH n_1441 GND GND efet
M2820 dpc40_ADLPCL cclk GND GND efet
M2821 n_929 n_1549 GND GND efet
M2822 x5 cclk n_578 GND efet
M2823 Vdd n_1191 ab6 GND efet
M2824 adl1 cclk Vdd GND efet
M2825 n_1586 op_T0_tsx GND GND efet
M2826 n_914 n_1316 GND GND efet
M2827 GND n_1499 n_709 GND efet
M2828 Vdd n_1191 ab6 GND efet
M2829 Vdd cclk adl0 GND efet
M2830 GND ir7 op_shift_right GND efet
M2831 n_1667 ADH_ABH nABH3 GND efet
M2832 GND idb5 n_1383 GND efet
M2833 n_1187 cclk nots6 GND efet
M2834 sb6 cclk Vdd GND efet
M2835 pch6 dpc30_ADHPCH adh6 GND efet
M2836 pch7 dpc30_ADHPCH adh7 GND efet
M2837 pch4 dpc30_ADHPCH adh4 GND efet
M2838 pch5 dpc30_ADHPCH adh5 GND efet
M2839 pch2 dpc30_ADHPCH adh2 GND efet
M2840 pch3 dpc30_ADHPCH adh3 GND efet
M2841 GND notir0 op_T4_ind_y GND efet
M2842 GND notir0 op_T2_ind_y GND efet
M2843 op_T4_ind_x notir0 GND GND efet
M2844 op_T2_abs_y notir0 GND GND efet
M2845 op_T2_ind_x notir0 GND GND efet
M2846 GND notir0 op_T0_eor GND efet
M2847 GND notir0 op_T0_ora GND efet
M2848 GND notir0 x_op_T3_ind_y GND efet
M2849 GND cclk n_346 GND efet
M2850 ab9 n_1140 Vdd GND efet
M2851 n_508 op_from_x GND GND efet
M2852 p0 cp1 n_1082 GND efet
M2853 GND n_190 n_220 GND efet
M2854 n_1247 n_38 Vdd GND efet
M2855 n_189 alua1 GND GND efet
M2856 GND alua1 n_A_B_1 GND efet
M2857 n_1451 cp1 n_212 GND efet
M2858 GND n_1247 dpc23_SBAC GND efet
M2859 n_1692 n_270 n_1082 GND efet
M2860 n_126 cclk n_1486 GND efet
M2861 ir2 n_1300 GND GND efet
M2862 op_T3_mem_abs ir4 GND GND efet
M2863 x_op_push_pull ir4 GND GND efet
M2864 op_T__cpx_cpy_imm_zp ir4 GND GND efet
M2865 op_T__asl_rol_a ir4 GND GND efet
M2866 op_T__cpx_cpy_abs ir4 GND GND efet
M2867 x_op_T4_rti ir4 GND GND efet
M2868 op_T0_plp ir4 GND GND efet
M2869 idb4 dpc25_SBDB sb4 GND efet
M2870 sb3 dpc25_SBDB idb3 GND efet
M2871 sb0 dpc25_SBDB idb0 GND efet
M2872 n_19 n_1708 GND GND efet
M2873 idb2 dpc25_SBDB sb2 GND efet
M2874 sb1 dpc25_SBDB idb1 GND efet
M2875 RnWstretched n_251 GND GND efet
M2876 RnWstretched n_251 GND GND efet
M2877 GND n_251 RnWstretched GND efet
M2878 GND n_251 RnWstretched GND efet
M2879 GND notir6 x_op_T__adc_sbc GND efet
M2880 op_T0_cli_sei notir6 GND GND efet
M2881 GND notir6 op_T__cpx_cpy_abs GND efet
M2882 GND notir6 x_op_T4_rti GND efet
M2883 GND n_646 n_272 GND efet
M2884 GND GND rdy GND efet
M2885 GND op_T0_pla n_1455 GND efet
M2886 GND nop_branch_bit7 n_1293 GND efet
M2887 adl5 dpc41_DL_ADL n_1387 GND efet
M2888 GND ir7 op_T5_rti_rts GND efet
M2889 GND ir7 op_T4_jmp GND efet
M2890 GND op_T2_brk n_824 GND efet
M2891 n_1402 n_293 n_57 GND efet
M2892 alub1 dpc8_nDBADD n_583 GND efet
M2893 adl6 dpc21_ADDADL alu6 GND efet
M2894 adl5 dpc21_ADDADL alu5 GND efet
M2895 n_1668 adh0 GND GND efet
M2896 alu7 dpc21_ADDADL adl7 GND efet
M2897 GND ir7 x_op_jmp GND efet
M2898 n_152 op_T2 GND GND efet
M2899 n_568 db5 GND GND efet
M2900 alub3 dpc8_nDBADD n_1621 GND efet
M2901 n_844 cclk n_459 GND efet
M2902 op_T2_mem_zp ir4 GND GND efet
M2903 adl4 dpc21_ADDADL alu4 GND efet
M2904 Vdd n_1399 cp1 GND efet
M2905 op_T4_mem_abs_idx _t4 GND GND efet
M2906 GND pipeUNK02 n_1492 GND efet
M2907 n_378 n_1357 GND GND efet
M2908 x_op_T0_bit ir4 GND GND efet
M2909 op_T5_rti_rts ir3 GND GND efet
M2910 n_831 dpc26_ACDB idb5 GND efet
M2911 op_jsr ir3 GND GND efet
M2912 op_brk_rti ir3 GND GND efet
M2913 op_T3_branch ir3 GND GND efet
M2914 n_1542 n_1345 n_1685 GND efet
M2915 op_T5_ind_x ir3 GND GND efet
M2916 op_T0_brk_rti ir3 GND GND efet
M2917 GND nDBZ n_580 GND efet
M2918 GND s0 n_983 GND efet
M2919 op_T3_mem_zp_idx ir3 GND GND efet
M2920 xx_op_T5_jsr ir3 GND GND efet
M2921 n_635 n_1523 Vdd GND efet
M2922 n_963 n_1523 GND GND efet
M2923 Vdd n_1260 dpc32_PCHADH GND efet
M2924 n_1413 n_1260 GND GND efet
M2925 n_474 cclk n_15 GND efet
M2926 n_21 n_1162 GND GND efet
M2927 GND n_962 nDBE GND efet
M2928 n_1169 dpc2_XSB sb0 GND efet
M2929 ADL_ABL n_220 Vdd GND efet
M2930 GND n_220 n_130 GND efet
M2931 n_1554 n_61 GND GND efet
M2932 n_1575 cclk pipeT2out GND efet
M2933 notx4 x4 GND GND efet
M2934 GND n_61 n_479 GND efet
M2935 GND pipeUNK09 n_941 GND efet
M2936 GND ir5 op_T__cmp GND efet
M2937 n_633 cclk n_1059 GND efet
M2938 n_25 n_256 GND GND efet
M2939 dor4 notdor4 GND GND efet
M2940 dasb6 n_479 GND GND efet
M2941 GND notir0 x_op_T__adc_sbc GND efet
M2942 GND notir0 op_T__cmp GND efet
M2943 op_T5_ind_x notir0 GND GND efet
M2944 x_op_T4_ind_y notir0 GND GND efet
M2945 GND notir0 op_T5_mem_ind_idx GND efet
M2946 GND GND db3 GND efet
M2947 n_330 n_538 n_881 GND efet
M2948 GND op_T5_brk n_689 GND efet
M2949 adh7 dpc42_DL_ADH n_1147 GND efet
M2950 adh6 dpc42_DL_ADH n_1014 GND efet
M2951 adh5 dpc42_DL_ADH n_1387 GND efet
M2952 adh4 dpc42_DL_ADH n_1095 GND efet
M2953 adh3 dpc42_DL_ADH n_1661 GND efet
M2954 adh2 dpc42_DL_ADH n_1424 GND efet
M2955 adh1 dpc42_DL_ADH n_87 GND efet
M2956 adh0 dpc42_DL_ADH n_719 GND efet
M2957 n_188 n_1606 GND GND efet
M2958 n_510 n_347 GND GND efet
M2959 n_1667 cp1 n_883 GND efet
M2960 sb4 cclk Vdd GND efet
M2961 n_973 cclk nots4 GND efet
M2962 n_518 cclk y6 GND efet
M2963 GND p0 n_31 GND efet
M2964 n_928 cp1 n_1378 GND efet
M2965 n_1309 cp1 n_74 GND efet
M2966 n_AxBxC_4 C34 n_375 GND efet
M2967 GND C34 _AxB_4_nC34 GND efet
M2968 pclp7 dpc38_PCLADL adl7 GND efet
M2969 adl0 dpc38_PCLADL pclp0 GND efet
M2970 GND notRdy0 n_1718 GND efet
M2971 clk1out n_747 Vdd GND efet
M2972 GND n_358 n_1715 GND efet
M2973 adl4 dpc38_PCLADL pclp4 GND efet
M2974 GND n_86 ab4 GND efet
M2975 GND n_86 ab4 GND efet
M2976 VEC0 notRdy0 GND GND efet
M2977 GND res n_312 GND efet
M2978 dpc27_SBADH n_1271 GND GND efet
M2979 GND idb0 DBZ GND efet
M2980 GND notRdy0 short_circuit_idx_add GND efet
M2981 nop_set_C op_T__cpx_cpy_abs GND GND efet
M2982 GND n_499 n_743 GND efet
M2983 GND n_499 n_1659 GND efet
M2984 alu2 dpc20_ADDSB06 sb2 GND efet
M2985 n_432 sb3 GND GND efet
M2986 dpc39_PCLPCL n_1270 Vdd GND efet
M2987 GND n_906 n_714 GND efet
M2988 n_432 sb3 GND GND efet
M2989 op_SUMS op_SRS GND GND efet
M2990 n_A_B_2 alua2 GND GND efet
M2991 GND n_1270 n_1518 GND efet
M2992 GND cclk n_1585 GND efet
M2993 op_T2_abs notir3 GND GND efet
M2994 op_T3_abs_idx notir3 GND GND efet
M2995 op_T__iny_dey notir3 GND GND efet
M2996 op_T0_php_pha notir3 GND GND efet
M2997 op_T3_plp_pla notir3 GND GND efet
M2998 op_jmp notir3 GND GND efet
M2999 op_T0_txs notir3 GND GND efet
M3000 op_T__dex notir3 GND GND efet
M3001 op_T__inx notir3 GND GND efet
M3002 op_T0_tsx notir3 GND GND efet
M3003 GND n_1295 n_1238 GND efet
M3004 n_1115 n_620 GND GND efet
M3005 GND op_T0_cld_sed n_774 GND efet
M3006 GND n_616 n_454 GND efet
M3007 GND cclk n_742 GND efet
M3008 GND nABL3 abl3 GND efet
M3009 GND n_620 n_922 GND efet
M3010 n_1147 dpc41_DL_ADL adl7 GND efet
M3011 dor6 notdor6 GND GND efet
M3012 n_1258 n_390 GND GND efet
M3013 GND dor6 n_471 GND efet
M3014 n_AxB1__C01 AxB1 GND GND efet
M3015 n_326 n_1356 GND GND efet
M3016 pclp6 dpc37_PCLDB idb6 GND efet
M3017 DA_AxB2 n_A_B_2 GND GND efet
M3018 n_637 nA_B7 GND GND efet
M3019 idb7 dpc43_DL_DB n_1147 GND efet
M3020 n_1368 NMIL GND GND efet
M3021 idb5 dpc43_DL_DB n_1387 GND efet
M3022 idb6 dpc43_DL_DB n_1014 GND efet
M3023 GND ir7 op_T0_plp GND efet
M3024 GND ir7 x_op_T4_rti GND efet
M3025 Vdd n_322 ab7 GND efet
M3026 ab7 n_322 Vdd GND efet
M3027 op_T0_cli_sei ir7 GND GND efet
M3028 GND ir7 op_T__bit GND efet
M3029 GND clock1 op_T0_cpy_iny GND efet
M3030 GND clock1 op_T0_tay_ldy_not_idx GND efet
M3031 GND ir7 xx_op_T5_jsr GND efet
M3032 GND ir7 op_T2_jmp_abs GND efet
M3033 GND ir7 x_op_T3_plp_pla GND efet
M3034 op_asl_rol ir7 GND GND efet
M3035 pd1_clearIR pd1 GND GND efet
M3036 n_1720 dor5 GND GND efet
M3037 n_612 dor5 GND GND efet
M3038 n_1339 cp1 n_597 GND efet
M3039 pclp5 npclp5 GND GND efet
M3040 n_436 notx4 GND GND efet
M3041 GND notx0 n_1169 GND efet
M3042 GND notir7 x_op_T0_tya GND efet
M3043 GND notir7 op_T0_iny_dey GND efet
M3044 GND n_AxB7__C67 n_AxBxC_7 GND efet
M3045 GND AxB3 n_1610 GND efet
M3046 p7 H1x1 idb7 GND efet
M3047 op_T0_pla irline3 GND GND efet
M3048 op_T0_tya irline3 GND GND efet
M3049 GND op_from_x n_734 GND efet
M3050 n_738 cp1 n_1519 GND efet
M3051 GND pipeUNK36 short_circuit_idx_add GND efet
M3052 GND n_862 n_445 GND efet
M3053 GND op_T3_jsr n_824 GND efet
M3054 n_499 pch5 GND GND efet
M3055 n_733 dpc0_YSB sb5 GND efet
M3056 n_518 dpc0_YSB sb6 GND efet
M3057 n_603 n_47 GND GND efet
M3058 n_658 dpc0_YSB sb4 GND efet
M3059 GND n_358 n_1129 GND efet
M3060 GND n_358 n_1129 GND efet
M3061 n_402 cp1 notRnWprepad GND efet
M3062 alub0 dpc9_DBADD idb0 GND efet
M3063 n_568 cclk notidl5 GND efet
M3064 Vdd cclk adh1 GND efet
M3065 n_871 dpc2_XSB sb7 GND efet
M3066 n_1717 cclk n_1113 GND efet
M3067 n_990 abl3 GND GND efet
M3068 n_138 abl3 GND GND efet
M3069 GND ir5 op_T0_eor GND efet
M3070 GND ir5 op_T5_rti GND efet
M3071 GND ir5 op_T0_php_pha GND efet
M3072 GND ir5 op_T0_tya GND efet
M3073 GND ir5 op_T0_cmp GND efet
M3074 op_T4_rti ir5 GND GND efet
M3075 GND ir5 op_T0_ora GND efet
M3076 GND ir5 op_T2_pha GND efet
M3077 GND ir5 op_T0_txa GND efet
M3078 GND ir7 op_T4_rts GND efet
M3079 GND _t3 op_T3_mem_abs GND efet
M3080 n_613 n_1682 n_150 GND efet
M3081 op_T3_jmp _t3 GND GND efet
M3082 GND _t3 op_T3_jsr GND efet
M3083 GND _t3 op_T3 GND efet
M3084 GND _t3 op_T3_abs_idx_ind GND efet
M3085 GND _t3 x_op_T3_abs_idx GND efet
M3086 GND _t3 op_T3_branch GND efet
M3087 GND _t3 x_op_T3_plp_pla GND efet
M3088 op_T3_mem_zp_idx _t3 GND GND efet
M3089 n_206 alucout GND GND efet
M3090 GND x_op_T0_tya n_1717 GND efet
M3091 GND n_241 n_1033 GND efet
M3092 GND op_T0_dex n_1106 GND efet
M3093 ab12 n_999 GND GND efet
M3094 GND n_999 ab12 GND efet
M3095 GND n_867 n_876 GND efet
M3096 pipeUNK22 cclk n_29 GND efet
M3097 n_975 n_995 n_886 GND efet
M3098 Vdd n_241 dpc21_ADDADL GND efet
M3099 n_612 RnWstretched GND GND efet
M3100 n_14 cclk pipeUNK20 GND efet
M3101 GND _t3 op_T3_ind_y GND efet
M3102 op_T3_ind_x _t3 GND GND efet
M3103 GND _t3 x_op_T3_ind_y GND efet
M3104 GND _t3 op_T3_abs_idx GND efet
M3105 GND n_291 n_1157 GND efet
M3106 n_811 alucout GND GND efet
M3107 n_696 cclk n_610 GND efet
M3108 GND n_794 db1 GND efet
M3109 GND n_794 db1 GND efet
M3110 db1 n_794 GND GND efet
M3111 db1 n_794 GND GND efet
M3112 x_op_T__adc_sbc cclk pipeUNK03 GND efet
M3113 db1 n_794 GND GND efet
M3114 db1 n_794 GND GND efet
M3115 db1 n_794 GND GND efet
M3116 op_T2_jsr _t2 GND GND efet
M3117 op_T2_ind_y _t2 GND GND efet
M3118 op_T2_pha _t2 GND GND efet
M3119 op_T2_stack_access _t2 GND GND efet
M3120 op_T2_branch _t2 GND GND efet
M3121 op_T2_brk _t2 GND GND efet
M3122 op_T2_ind _t2 GND GND efet
M3123 op_T2_zp_zp_idx _t2 GND GND efet
M3124 op_T2_php _t2 GND GND efet
M3125 op_T2_abs_access _t2 GND GND efet
M3126 GND op_T0_jsr n_1058 GND efet
M3127 Vdd n_42 db3 GND efet
M3128 GND n_196 dpc5_SADL GND efet
M3129 n_A_B_5 dpc13_ORS naluresult5 GND efet
M3130 GND op_T3_plp_pla n_1464 GND efet
M3131 GND n_18 n_378 GND efet
M3132 GND n_1247 dpc31_PCHPCH GND efet
M3133 dpc26_ACDB n_800 GND GND efet
M3134 adl6 dpc41_DL_ADL n_1014 GND efet
M3135 GND n_345 n_1097 GND efet
M3136 GND noty1 n_767 GND efet
M3137 GND AxB7 n_AxB7__C67 GND efet
M3138 dasb3 n_345 n_1686 GND efet
M3139 GND n_171 ab7 GND efet
M3140 GND n_171 ab7 GND efet
M3141 n_1154 n_959 GND GND efet
M3142 GND n_171 ab7 GND efet
M3143 n_416 ADL_ABL nABL1 GND efet
M3144 GND n_1007 dpc35_PCHC GND efet
M3145 GND adl7 n_1046 GND efet
M3146 n_389 n_1107 GND GND efet
M3147 noty2 y2 GND GND efet
M3148 GND AxB7 n_1013 GND efet
M3149 n_1387 cp1 idl5 GND efet
M3150 GND n_815 n_0_ADL2 GND efet
M3151 n_1724 cclk x6 GND efet
M3152 GND op_T4_ind_x n_1649 GND efet
M3153 adl3 cclk Vdd GND efet
M3154 n_591 n_1258 GND GND efet
M3155 n_AxBxC_1 dpc17_SUMS naluresult1 GND efet
M3156 n_AxBxC_0 dpc17_SUMS naluresult0 GND efet
M3157 GND n_1238 dpc25_SBDB GND efet
M3158 GND pipeUNK28 n_1598 GND efet
M3159 n_AxBxC_3 dpc17_SUMS naluresult3 GND efet
M3160 n_AxBxC_2 dpc17_SUMS naluresult2 GND efet
M3161 GND n_635 ab14 GND efet
M3162 ab14 n_635 GND GND efet
M3163 nop_branch_bit6 ir6 GND GND efet
M3164 op_T__asl_rol_a ir6 GND GND efet
M3165 GND ir6 op_T0_clc_sec GND efet
M3166 GND ir6 op_T__bit GND efet
M3167 op_asl_rol ir6 GND GND efet
M3168 n_A_B_3 alub3 GND GND efet
M3169 xx_op_T5_jsr ir6 GND GND efet
M3170 pipeUNK09 cclk n_327 GND efet
M3171 ab14 n_635 GND GND efet
M3172 x_op_push_pull ir2 GND GND efet
M3173 op_implied ir2 GND GND efet
M3174 op_clv ir2 GND GND efet
M3175 GND notir5 op_T0_tay GND efet
M3176 GND notir5 op_T0_tax GND efet
M3177 op_T5_mem_ind_idx ir2 GND GND efet
M3178 GND notir5 op_T2_jsr GND efet
M3179 GND notir5 op_T0_sbc GND efet
M3180 GND notir5 op_T0_adc_sbc GND efet
M3181 GND notir5 op_rol_ror GND efet
M3182 GND notir5 op_T5_jsr GND efet
M3183 GND notir5 op_T__adc_sbc GND efet
M3184 GND notir5 op_T0_pla GND efet
M3185 GND notir5 op_T0_lda GND efet
M3186 n_1391 op_T2_php GND GND efet
M3187 GND _AxB_6_nC56 n_AxBxC_6 GND efet
M3188 DC78_phi2 cclk DC78 GND efet
M3189 GND nnT2BR n_104 GND efet
M3190 n_1347 nnT2BR GND GND efet
M3191 n_207 cclk n_1061 GND efet
M3192 n_571 cp1 n_343 GND efet
M3193 GND rdy n_958 GND efet
M3194 n_473 n_980 n_1004 GND efet
M3195 dpc43_DL_DB n_1240 GND GND efet
M3196 Vdd n_963 ab14 GND efet
M3197 n_31 cclk pipeUNK16 GND efet
M3198 notx2 x2 GND GND efet
M3199 dpc34_PCLC n_249 GND GND efet
M3200 GND n_335 n_1280 GND efet
M3201 GND n_440 n_813 GND efet
M3202 nTWOCYCLE PD_xxx010x1 GND GND efet
M3203 n_1549 a1 GND GND efet
M3204 n_1602 cclk n_506 GND efet
M3205 n_1650 cp1 n_94 GND efet
M3206 GND n_95 n_531 GND efet
M3207 GND n_770 n_853 GND efet
M3208 GND op_T0_eor n_837 GND efet
M3209 n_AxBxC_0 n_105 n_406 GND efet
M3210 GND n_1575 _t2 GND efet
M3211 n_818 n_265 GND GND efet
M3212 n_367 n_206 n_1082 GND efet
M3213 n_267 n_544 GND GND efet
M3214 Vdd n_631 dpc37_PCLDB GND efet
M3215 GND n_631 n_1323 GND efet
M3216 GND n_105 _AxB_0_nC0in GND efet
M3217 Vdd cclk adl4 GND efet
M3218 n_616 op_T__iny_dey GND GND efet
M3219 dpc34_PCLC n_329 GND GND efet
M3220 n_1166 n_329 GND GND efet
M3221 db0 n_1072 GND GND efet
M3222 n_1107 op_T4_ind_y GND GND efet
M3223 db0 n_1072 GND GND efet
M3224 GND n_1072 db0 GND efet
M3225 db0 n_1072 GND GND efet
M3226 GND n_1072 db0 GND efet
M3227 db0 n_1072 GND GND efet
M3228 GND n_1072 db0 GND efet
M3229 nA_B2 alub2 n_452 GND efet
M3230 pd6_clearIR pd6 GND GND efet
M3231 n_508 n_335 n_1303 GND efet
M3232 GND op_T5_rts n_256 GND efet
M3233 n_1684 idb6 GND GND efet
M3234 GND n_503 n_270 GND efet
M3235 notRdy0 cp1 n_1272 GND efet
M3236 n_724 fetch n_310 GND efet
M3237 n_237 fetch n_119 GND efet
M3238 op_implied ir0 GND GND efet
M3239 GND n_689 VEC0 GND efet
M3240 n_726 op_T3_abs_idx_ind GND GND efet
M3241 GND pcl1 n_329 GND efet
M3242 GND n_1715 n_1399 GND efet
M3243 GND n_1715 n_1399 GND efet
M3244 GND ir7 op_T3_plp_pla GND efet
M3245 GND ir7 op_T5_rti GND efet
M3246 GND ir7 op_ror GND efet
M3247 op_jmp ir7 GND GND efet
M3248 op_T0_ora ir7 GND GND efet
M3249 GND ir7 op_T3_stack_bit_jmp GND efet
M3250 GND ir7 op_T4_brk_jsr GND efet
M3251 GND ir7 op_T4_rti GND efet
M3252 n_374 db6 GND GND efet
M3253 Pout3 H1x1 idb3 GND efet
M3254 n_AxB_6 nA_B6 n_482 GND efet
M3255 res GND GND GND efet
M3256 GND n_1579 n_221 GND efet
M3257 p4 H1x1 idb4 GND efet
M3258 GND clk0 n_358 GND efet
M3259 GND n_1222 n_1090 GND efet
M3260 GND op_T0_iny_dey n_1717 GND efet
M3261 x0 dpc3_SBX sb0 GND efet
M3262 n_135 n_519 Vdd GND efet
M3263 GND n_519 n_127 GND efet
M3264 Vdd n_543 dpc5_SADL GND efet
M3265 n_196 n_543 GND GND efet
M3266 GND n_1124 n_1662 GND efet
M3267 alub0 dpc8_nDBADD n_624 GND efet
M3268 n_1358 op_T0_txs GND GND efet
M3269 n_1093 cp1 n_226 GND efet
M3270 n_1593 n_226 GND GND efet
M3271 nABH4 ADH_ABH n_1451 GND efet
M3272 n_753 n_811 GND GND efet
M3273 GND n_1269 n_1401 GND efet
M3274 GND ir7 op_T0_clc_sec GND efet
M3275 GND ir7 x_op_T0_bit GND efet
M3276 notir6 ir6 GND GND efet
M3277 GND n_1225 n_1222 GND efet
M3278 GND nots4 n_3 GND efet
M3279 n_1422 pipeUNK06 n_754 GND efet
M3280 n_930 n_1276 GND GND efet
M3281 GND dpc29_0ADH17 adh1 GND efet
M3282 GND RnWstretched n_1076 GND efet
M3283 GND notRdy0 n_16 GND efet
M3284 n_213 db1 GND GND efet
M3285 GND pipeVectorA1 n_0_ADL1 GND efet
M3286 GND nots5 n_280 GND efet
M3287 n_1654 cclk a3 GND efet
M3288 n_705 ADH_ABH nABH0 GND efet
M3289 n_6 n_521 GND GND efet
M3290 Vdd n_317 n_417 GND efet
M3291 GND n_919 n_200 GND efet
M3292 n_1486 n_919 n_1538 GND efet
M3293 n_1229 n_919 n_835 GND efet
M3294 n_871 cclk x7 GND efet
M3295 n_1449 n_958 GND GND efet
M3296 ir4 n_927 GND GND efet
M3297 PD_1xx000x0 n_1605 GND GND efet
M3298 alub7 dpc8_nDBADD n_423 GND efet
M3299 GND clearIR pd1_clearIR GND efet
M3300 n_1655 n_1211 GND GND efet
M3301 y3 cclk n_1531 GND efet
M3302 n_202 n_480 n_629 GND efet
M3303 n_1514 cp1 n_880 GND efet
M3304 dpc11_SBADD n_708 GND GND efet
M3305 n_1304 n_673 GND GND efet
M3306 npclp4 n_15 GND GND efet
M3307 GND alucin notalucin GND efet
M3308 n_472 cp1 n_1606 GND efet
M3309 pipeUNK05 cclk n_90 GND efet
M3310 op_T0_cli_sei notir4 GND GND efet
M3311 op_T4_mem_abs_idx notir4 GND GND efet
M3312 n_889 cclk pipeUNK42 GND efet
M3313 n_1619 n_182 GND GND efet
M3314 n_242 cclk x3 GND efet
M3315 nC34 DC34 GND GND efet
M3316 sb4 dpc6_SBS s4 GND efet
M3317 s3 dpc6_SBS sb3 GND efet
M3318 s2 dpc6_SBS sb2 GND efet
M3319 s1 dpc6_SBS sb1 GND efet
M3320 GND n_AxB_0 n_406 GND efet
M3321 n_802 n_781 GND GND efet
M3322 nC56 n_647 GND GND efet
M3323 GND n_AxB_0 _AxB_0_nC0in GND efet
M3324 sb4 dpc3_SBX x4 GND efet
M3325 n_1080 n_811 GND GND efet
M3326 pipephi2Reset0 cclk Reset0 GND efet
M3327 Vdd n_634 ab4 GND efet
M3328 Vdd n_634 ab4 GND efet
M3329 n_396 n_1358 GND GND efet
M3330 GND notRdy0 n_781 GND efet
M3331 GND C1x5Reset notRnWprepad GND efet
M3332 n_1649 cclk n_1027 GND efet
M3333 ab3 n_138 GND GND efet
M3334 ab3 n_138 GND GND efet
M3335 ab3 n_138 GND GND efet
M3336 GND n_1277 n_1441 GND efet
M3337 n_1037 cclk n_266 GND efet
M3338 n_1675 fetch n_74 GND efet
M3339 n_1609 fetch n_1378 GND efet
M3340 irline3 n_1133 GND GND efet
M3341 n_856 dpc34_PCLC n_919 GND efet
M3342 n_632 n_1289 n_1058 GND efet
M3343 GND pipeUNK37 n_198 GND efet
M3344 GND pipeUNK37 n_198 GND efet
M3345 GND nIRQP n_1092 GND efet
M3346 GND dpc29_0ADH17 adh7 GND efet
M3347 GND op_T3_stack_bit_jmp n_604 GND efet
M3348 n_1230 n_360 GND GND efet
M3349 A_B0 n_A_B_0 GND GND efet
M3350 n_326 dpc26_ACDB idb6 GND efet
M3351 idl0 notidl0 GND GND efet
M3352 op_T3_abs_idx_ind op_push_pull GND GND efet
M3353 op_T4_brk ir3 GND GND efet
M3354 n_970 n_149 GND GND efet
M3355 GND alub6 n_A_B_6 GND efet
M3356 n_1483 alub6 nA_B6 GND efet
M3357 op_branch_done n_603 GND GND efet
M3358 op_T2_abs_access op_push_pull GND GND efet
M3359 pd4_clearIR pd4 GND GND efet
M3360 GND idb4 n_478 GND efet
M3361 GND n_149 n_762 GND efet
M3362 n_1592 dpc26_ACDB idb7 GND efet
M3363 n_1568 n_1345 GND GND efet
M3364 x_op_T4_ind_y ir3 GND GND efet
M3365 naluresult2 dpc13_ORS n_A_B_2 GND efet
M3366 n_1180 cp1 n_1533 GND efet
M3367 op_T5_rts ir7 GND GND efet
M3368 GND ir7 op_T0_brk_rti GND efet
M3369 n_1041 n_990 GND GND efet
M3370 n_138 n_990 Vdd GND efet
M3371 GND n_1357 n_1575 GND efet
M3372 n_795 n_1649 GND GND efet
M3373 n_207 n_293 n_356 GND efet
M3374 n_810 n_293 GND GND efet
M3375 n_734 n_335 n_1106 GND efet
M3376 n_330 n_807 GND GND efet
M3377 adh5 cclk Vdd GND efet
M3378 adl6 cclk Vdd GND efet
M3379 GND pipeUNK04 n_1644 GND efet
M3380 dpc16_EORS n_108 GND GND efet
M3381 dor0 notdor0 GND GND efet
M3382 n_1245 aluvout GND GND efet
M3383 n_1169 cclk x0 GND efet
M3384 n_588 cclk notidl7 GND efet
M3385 n_1446 n_850 GND GND efet
M3386 short_circuit_branch_add n_850 GND GND efet
M3387 GND notir7 op_T0_sbc GND efet
M3388 GND notir7 op_T0_cmp GND efet
M3389 GND notir7 op_T0_cpx_cpy_inx_iny GND efet
M3390 GND notir7 op_inc_nop GND efet
M3391 GND notir7 op_T0_tay_ldy_not_idx GND efet
M3392 GND notir7 op_T0_ldy_mem GND efet
M3393 GND notir7 op_T0_txa GND efet
M3394 GND notir7 op_T0_tya GND efet
M3395 op_T5_jsr ir4 GND GND efet
M3396 op_T2_stack_access ir4 GND GND efet
M3397 n_732 nTWOCYCLE_phi1 n_106 GND efet
M3398 op_T__shift_a ir4 GND GND efet
M3399 op_T0_txa ir4 GND GND efet
M3400 op_T0_pla ir4 GND GND efet
M3401 op_T0_tay ir4 GND GND efet
M3402 op_T0_shift_a ir4 GND GND efet
M3403 op_T0_tax ir4 GND GND efet
M3404 GND n_1542 n_1253 GND efet
M3405 alub6 dpc8_nDBADD n_351 GND efet
M3406 alub5 dpc8_nDBADD n_1383 GND efet
M3407 GND noty4 n_658 GND efet
M3408 GND pipeUNK23 n_819 GND efet
M3409 n_637 C67 GND GND efet
M3410 notaluvout C67 n_1489 GND efet
M3411 GND n_1247 dpc2_XSB GND efet
M3412 nop_set_C op_T__asl_rol_a GND GND efet
M3413 GND n_1335 dpc24_ACSB GND efet
M3414 n_807 n_1599 n_431 GND efet
M3415 n_231 PD_xxxx10x0 GND GND efet
M3416 pclp6 npclp6 GND GND efet
M3417 n_104 n_275 GND GND efet
M3418 n_1515 PD_xxxx10x0 nTWOCYCLE GND efet
M3419 GND nA_B2 DA_AB2 GND efet
M3420 ADL_ABL n_130 GND GND efet
M3421 GND notx1 n_1709 GND efet
M3422 GND nots2 n_1389 GND efet
M3423 GND notRdy0 n_1120 GND efet
M3424 n_1039 notRdy0 n_2 GND efet
M3425 ab3 n_1041 Vdd GND efet
M3426 n_1624 cp1 notRdy0 GND efet
M3427 n_616 op_T0_tay_ldy_not_idx GND GND efet
M3428 ab4 n_86 GND GND efet
M3429 GND n_86 ab4 GND efet
M3430 n_484 n_1386 n_914 GND efet
M3431 n_307 n_31 GND GND efet
M3432 n_1580 sb2 GND GND efet
M3433 n_1580 sb2 GND GND efet
M3434 GND n_759 n_944 GND efet
M3435 n_1300 fetch n_343 GND efet
M3436 n_1189 n_1714 n_262 GND efet
M3437 GND op_T__ora_and_eor_adc n_1455 GND efet
M3438 GND n_676 ab9 GND efet
M3439 ab9 n_676 GND GND efet
M3440 GND n_1346 n_1296 GND efet
M3441 GND op_implied n_664 GND efet
M3442 n_359 n_1346 Vdd GND efet
M3443 IRQP cp1 n_330 GND efet
M3444 GND op_T__shift_a n_1455 GND efet
M3445 alu7 dpc19_ADDSB7 sb7 GND efet
M3446 GND notx7 n_871 GND efet
M3447 n_1712 cclk pipeVectorA2 GND efet
M3448 op_T__asl_rol_a ir2 GND GND efet
M3449 x_op_T4_rti ir2 GND GND efet
M3450 op_T0_plp ir2 GND GND efet
M3451 op_T0_cld_sed ir2 GND GND efet
M3452 n_810 n_923 GND GND efet
M3453 GND AxB1 n_AxB_1 GND efet
M3454 cclk n_1467 GND GND efet
M3455 cclk n_1467 GND GND efet
M3456 GND notir6 op_shift_right GND efet
M3457 op_T5_rts notir6 GND GND efet
M3458 GND notir6 op_T0_jmp GND efet
M3459 GND notir6 x_op_jmp GND efet
M3460 op_T__adc_sbc notir6 GND GND efet
M3461 op_T0_pla notir6 GND GND efet
M3462 GND notir6 op_T2_pha GND efet
M3463 GND notir6 op_T0_shift_right_a GND efet
M3464 GND notir6 op_T4_jmp GND efet
M3465 GND notir6 op_T5_rti_rts GND efet
M3466 GND clearIR pd3_clearIR GND efet
M3467 GND clearIR pd4_clearIR GND efet
M3468 dpc34_PCLC n_1643 GND GND efet
M3469 dpc23_SBAC n_830 Vdd GND efet
M3470 GND n_1643 n_766 GND efet
M3471 GND n_902 n_1289 GND efet
M3472 n_1047 n_830 GND GND efet
M3473 Vdd n_417 sync GND efet
M3474 Vdd n_417 sync GND efet
M3475 Vdd n_417 sync GND efet
M3476 sync n_417 Vdd GND efet
M3477 n_1211 nnT2BR GND GND efet
M3478 n_1211 nnT2BR GND GND efet
M3479 n_1211 n_1286 GND GND efet
M3480 GND _t4 op_T4_rts GND efet
M3481 GND _t4 op_T4_brk_jsr GND efet
M3482 op_T4_rti _t4 GND GND efet
M3483 GND op_T2_jsr n_383 GND efet
M3484 n_1560 op_T0_cpx_cpy_inx_iny GND GND efet
M3485 n_225 n_1223 GND GND efet
M3486 Vdd n_1223 dpc9_DBADD GND efet
M3487 GND pipeUNK06 n_755 GND efet
M3488 n_496 cclk nots5 GND efet
M3489 op_T3_branch notir4 GND GND efet
M3490 op_T3_mem_zp_idx notir4 GND GND efet
M3491 op_T0_clc_sec notir4 GND GND efet
M3492 GND notir4 op_T0_cld_sed GND efet
M3493 GND adh2 n_168 GND efet
M3494 op_clv notir4 GND GND efet
M3495 adl2 dpc10_ADLADD alub2 GND efet
M3496 op_T0_tsx ir6 GND GND efet
M3497 op_T0_ldy_mem ir6 GND GND efet
M3498 GND ir6 x_op_T0_tya GND efet
M3499 GND ir6 op_xy GND efet
M3500 GND idb0 n_1224 GND efet
M3501 n_1303 n_335 n_1397 GND efet
M3502 GND cclk dpc30_ADHPCH GND efet
M3503 GND cclk dpc31_PCHPCH GND efet
M3504 n_600 n_1341 GND GND efet
M3505 GND op_T2_jsr n_300 GND efet
M3506 ab1 n_66 GND GND efet
M3507 ab1 n_66 GND GND efet
M3508 ab1 n_66 GND GND efet
M3509 ab1 n_66 GND GND efet
M3510 n_973 n_973 Vdd GND efet
M3511 n_975 n_975 Vdd GND efet
M3512 n_964 n_964 Vdd GND efet
M3513 n_AxBxC_1 n_AxBxC_1 Vdd GND efet
M3514 n_961 n_961 Vdd GND efet
M3515 n_962 n_962 Vdd GND efet
M3516 n_969 n_969 Vdd GND efet
M3517 _t2 _t2 Vdd GND efet
M3518 n_966 n_966 Vdd GND efet
M3519 nnT2BR nnT2BR Vdd GND efet
M3520 n_200 n_200 Vdd GND efet
M3521 n_201 n_201 Vdd GND efet
M3522 notir0 notir0 Vdd GND efet
M3523 n_191 n_191 Vdd GND efet
M3524 n_A_B_7 n_A_B_7 Vdd GND efet
M3525 op_T0_shift_a op_T0_shift_a Vdd GND efet
M3526 n_1391 n_1391 Vdd GND efet
M3527 n_1389 n_1389 Vdd GND efet
M3528 notir5 notir5 Vdd GND efet
M3529 n_1392 n_1392 Vdd GND efet
M3530 n_1383 n_1383 Vdd GND efet
M3531 n_1386 n_1386 Vdd GND efet
M3532 op_T5_mem_ind_idx op_T5_mem_ind_idx Vdd GND efet
M3533 n_1433 n_1433 Vdd GND efet
M3534 n_428 n_428 Vdd GND efet
M3535 Pout3 Pout3 Vdd GND efet
M3536 n_1368 n_1368 Vdd GND efet
M3537 n_1364 n_1364 Vdd GND efet
M3538 n_1358 n_1358 Vdd GND efet
M3539 n_1357 n_1357 Vdd GND efet
M3540 n_1356 n_1356 Vdd GND efet
M3541 op_T0_cmp op_T0_cmp Vdd GND efet
M3542 nWR nWR Vdd GND efet
M3543 INTG INTG Vdd GND efet
M3544 p7 p7 Vdd GND efet
M3545 n_1369 n_1369 Vdd GND efet
M3546 n_774 n_774 Vdd GND efet
M3547 abh5 abh5 Vdd GND efet
M3548 op_jmp op_jmp Vdd GND efet
M3549 alu7 alu7 Vdd GND efet
M3550 n_767 n_767 Vdd GND efet
M3551 n_769 n_769 Vdd GND efet
M3552 n_770 n_770 Vdd GND efet
M3553 n_771 n_771 Vdd GND efet
M3554 n_772 n_772 Vdd GND efet
M3555 n_773 n_773 Vdd GND efet
M3556 n_1214 n_1214 Vdd GND efet
M3557 n_1213 n_1213 Vdd GND efet
M3558 n_AxB7__C67 n_AxB7__C67 Vdd GND efet
M3559 notx4 notx4 Vdd GND efet
M3560 n_484 n_484 Vdd GND efet
M3561 nA_B5 nA_B5 Vdd GND efet
M3562 n_476 n_476 Vdd GND efet
M3563 n_474 n_474 Vdd GND efet
M3564 n_473 n_473 Vdd GND efet
M3565 pclp2 pclp2 Vdd GND efet
M3566 n_480 n_480 Vdd GND efet
M3567 n_479 n_479 Vdd GND efet
M3568 n_478 n_478 Vdd GND efet
M3569 n_1714 n_1714 Vdd GND efet
M3570 n_1715 n_1715 Vdd GND efet
M3571 n_638 n_638 Vdd GND efet
M3572 n_637 n_637 Vdd GND efet
M3573 n_636 n_636 Vdd GND efet
M3574 n_632 n_632 Vdd GND efet
M3575 n_631 n_631 Vdd GND efet
M3576 n_630 n_630 Vdd GND efet
M3577 n_629 n_629 Vdd GND efet
M3578 n_628 n_628 Vdd GND efet
M3579 n_626 n_626 Vdd GND efet
M3580 n_625 n_625 Vdd GND efet
M3581 ir5 ir5 Vdd GND efet
M3582 ir7 ir7 Vdd GND efet
M3583 n_1316 n_1316 Vdd GND efet
M3584 n_1315 n_1315 Vdd GND efet
M3585 n_1319 n_1319 Vdd GND efet
M3586 nA_B7 nA_B7 Vdd GND efet
M3587 n_1323 n_1323 Vdd GND efet
M3588 notir7 notir7 Vdd GND efet
M3589 nC78 nC78 Vdd GND efet
M3590 op_T__shift_a op_T__shift_a Vdd GND efet
M3591 npclp6 npclp6 Vdd GND efet
M3592 n_732 n_732 Vdd GND efet
M3593 n_728 n_728 Vdd GND efet
M3594 notx6 notx6 Vdd GND efet
M3595 n_739 n_739 Vdd GND efet
M3596 n_743 n_743 Vdd GND efet
M3597 n_733 n_733 Vdd GND efet
M3598 n_735 n_735 Vdd GND efet
M3599 DBZ DBZ Vdd GND efet
M3600 dor1 dor1 Vdd GND efet
M3601 op_T0_cli_sei op_T0_cli_sei Vdd GND efet
M3602 pd2_clearIR pd2_clearIR Vdd GND efet
M3603 n_1668 n_1668 Vdd GND efet
M3604 n_1655 n_1655 Vdd GND efet
M3605 op_T0_cpx_inx op_T0_cpx_inx Vdd GND efet
M3606 n_1657 n_1657 Vdd GND efet
M3607 n_1662 n_1662 Vdd GND efet
M3608 n_1660 n_1660 Vdd GND efet
M3609 op_T__asl_rol_a op_T__asl_rol_a Vdd GND efet
M3610 op_T__inx op_T__inx Vdd GND efet
M3611 n_700 n_700 Vdd GND efet
M3612 n_AxB_2 n_AxB_2 Vdd GND efet
M3613 notir1 notir1 Vdd GND efet
M3614 n_708 n_708 Vdd GND efet
M3615 n_694 n_694 Vdd GND efet
M3616 n_695 n_695 Vdd GND efet
M3617 n_696 n_696 Vdd GND efet
M3618 nDA_ADD2 nDA_ADD2 Vdd GND efet
M3619 n_709 n_709 Vdd GND efet
M3620 op_T2_jsr op_T2_jsr Vdd GND efet
M3621 n_196 n_196 Vdd GND efet
M3622 n_198 n_198 Vdd GND efet
M3623 _AxB_2_nC12 _AxB_2_nC12 Vdd GND efet
M3624 n_192 n_192 Vdd GND efet
M3625 notRnWprepad notRnWprepad Vdd GND efet
M3626 n_188 n_188 Vdd GND efet
M3627 ir2 ir2 Vdd GND efet
M3628 noty0 noty0 Vdd GND efet
M3629 n_1026 n_1026 Vdd GND efet
M3630 n_1010 n_1010 Vdd GND efet
M3631 n_1016 n_1016 Vdd GND efet
M3632 notx5 notx5 Vdd GND efet
M3633 PD_xxxx10x0 PD_xxxx10x0 Vdd GND efet
M3634 A_B1 A_B1 Vdd GND efet
M3635 C23 C23 Vdd GND efet
M3636 n_1024 n_1024 Vdd GND efet
M3637 n_311 n_311 Vdd GND efet
M3638 n_312 n_312 Vdd GND efet
M3639 n_AxB_4 n_AxB_4 Vdd GND efet
M3640 op_T2_jmp_abs op_T2_jmp_abs Vdd GND efet
M3641 n_306 n_306 Vdd GND efet
M3642 n_307 n_307 Vdd GND efet
M3643 PD_xxx010x1 PD_xxx010x1 Vdd GND efet
M3644 op_T0_bit op_T0_bit Vdd GND efet
M3645 alu5 alu5 Vdd GND efet
M3646 n_317 n_317 Vdd GND efet
M3647 ir1 ir1 Vdd GND efet
M3648 op_T0_eor op_T0_eor Vdd GND efet
M3649 pd0_clearIR pd0_clearIR Vdd GND efet
M3650 n_1621 n_1621 Vdd GND efet
M3651 n_A_B_5 n_A_B_5 Vdd GND efet
M3652 n_1631 n_1631 Vdd GND efet
M3653 n_1629 n_1629 Vdd GND efet
M3654 nA_B0 nA_B0 Vdd GND efet
M3655 n_1635 n_1635 Vdd GND efet
M3656 dor2 dor2 Vdd GND efet
M3657 op_T3_abs_idx_ind op_T3_abs_idx_ind Vdd GND efet
M3658 n_678 n_678 Vdd GND efet
M3659 n_673 n_673 Vdd GND efet
M3660 n_674 n_674 Vdd GND efet
M3661 n_669 n_669 Vdd GND efet
M3662 n_670 n_670 Vdd GND efet
M3663 op_T0_ldy_mem op_T0_ldy_mem Vdd GND efet
M3664 pd5_clearIR pd5_clearIR Vdd GND efet
M3665 n_662 n_662 Vdd GND efet
M3666 n_664 n_664 Vdd GND efet
M3667 op_T2_ind_y op_T2_ind_y Vdd GND efet
M3668 n_1295 n_1295 Vdd GND efet
M3669 pchp5 pchp5 Vdd GND efet
M3670 n_1281 n_1281 Vdd GND efet
M3671 C01 C01 Vdd GND efet
M3672 n_1286 n_1286 Vdd GND efet
M3673 n_1289 n_1289 Vdd GND efet
M3674 n_1290 n_1290 Vdd GND efet
M3675 n_1293 n_1293 Vdd GND efet
M3676 PD_1xx000x0 PD_1xx000x0 Vdd GND efet
M3677 n_1045 n_1045 Vdd GND efet
M3678 n_1046 n_1046 Vdd GND efet
M3679 n_1043 n_1043 Vdd GND efet
M3680 n_1044 n_1044 Vdd GND efet
M3681 x_op_push_pull x_op_push_pull Vdd GND efet
M3682 x_op_jmp x_op_jmp Vdd GND efet
M3683 n_1047 n_1047 Vdd GND efet
M3684 nop_branch_done nop_branch_done Vdd GND efet
M3685 n_1054 n_1054 Vdd GND efet
M3686 n_1055 n_1055 Vdd GND efet
M3687 n_1593 n_1593 Vdd GND efet
M3688 n_1592 n_1592 Vdd GND efet
M3689 n_1595 n_1595 Vdd GND efet
M3690 n_1594 n_1594 Vdd GND efet
M3691 pd3_clearIR pd3_clearIR Vdd GND efet
M3692 n_1586 n_1586 Vdd GND efet
M3693 op_T4_jmp op_T4_jmp Vdd GND efet
M3694 n_1588 n_1588 Vdd GND efet
M3695 idl0 idl0 Vdd GND efet
M3696 n_1596 n_1596 Vdd GND efet
M3697 n_334 n_334 Vdd GND efet
M3698 DC78 DC78 Vdd GND efet
M3699 n_332 n_332 Vdd GND efet
M3700 alu6 alu6 Vdd GND efet
M3701 n_340 n_340 Vdd GND efet
M3702 ir6 ir6 Vdd GND efet
M3703 nA_B6 nA_B6 Vdd GND efet
M3704 n_335 n_335 Vdd GND efet
M3705 x_op_T3_ind_y x_op_T3_ind_y Vdd GND efet
M3706 op_T4 op_T4 Vdd GND efet
M3707 n_1082 n_1082 Vdd GND efet
M3708 n_1083 n_1083 Vdd GND efet
M3709 n_A_B_6 n_A_B_6 Vdd GND efet
M3710 n_1085 n_1085 Vdd GND efet
M3711 n_1075 n_1075 Vdd GND efet
M3712 clearIR clearIR Vdd GND efet
M3713 npclp2 npclp2 Vdd GND efet
M3714 n_1081 n_1081 Vdd GND efet
M3715 op_T2_pha op_T2_pha Vdd GND efet
M3716 n_1087 n_1087 Vdd GND efet
M3717 n_1566 n_1566 Vdd GND efet
M3718 notx7 notx7 Vdd GND efet
M3719 n_1560 n_1560 Vdd GND efet
M3720 op_brk_rti op_brk_rti Vdd GND efet
M3721 n_1552 n_1552 Vdd GND efet
M3722 n_1549 n_1549 Vdd GND efet
M3723 BRtaken BRtaken Vdd GND efet
M3724 x_op_T0_txa x_op_T0_txa Vdd GND efet
M3725 pchp4 pchp4 Vdd GND efet
M3726 n_29 n_29 Vdd GND efet
M3727 n_17 n_17 Vdd GND efet
M3728 n_19 n_19 Vdd GND efet
M3729 n_20 n_20 Vdd GND efet
M3730 n_21 n_21 Vdd GND efet
M3731 n_AxBxC_2 n_AxBxC_2 Vdd GND efet
M3732 n_23 n_23 Vdd GND efet
M3733 n_25 n_25 Vdd GND efet
M3734 notir4 notir4 Vdd GND efet
M3735 n_1457 n_1457 Vdd GND efet
M3736 n_1455 n_1455 Vdd GND efet
M3737 n_AxB_6 n_AxB_6 Vdd GND efet
M3738 pclp6 pclp6 Vdd GND efet
M3739 n_1462 n_1462 Vdd GND efet
M3740 pd6_clearIR pd6_clearIR Vdd GND efet
M3741 n_1464 n_1464 Vdd GND efet
M3742 n_1463 n_1463 Vdd GND efet
M3743 op_rol_ror op_rol_ror Vdd GND efet
M3744 n_374 n_374 Vdd GND efet
M3745 n_372 n_372 Vdd GND efet
M3746 n_378 n_378 Vdd GND efet
M3747 abl1 abl1 Vdd GND efet
M3748 n_368 n_368 Vdd GND efet
M3749 n_366 n_366 Vdd GND efet
M3750 n_AxBxC_0 n_AxBxC_0 Vdd GND efet
M3751 op_T5_brk op_T5_brk Vdd GND efet
M3752 op_T0_iny_dey op_T0_iny_dey Vdd GND efet
M3753 dpc36_nIPC dpc36_nIPC Vdd GND efet
M3754 idl6 idl6 Vdd GND efet
M3755 op_T0_clc_sec op_T0_clc_sec Vdd GND efet
M3756 n_1115 n_1115 Vdd GND efet
M3757 n_1111 n_1111 Vdd GND efet
M3758 ir4 ir4 Vdd GND efet
M3759 n_1109 n_1109 Vdd GND efet
M3760 n_1110 n_1110 Vdd GND efet
M3761 n_1106 n_1106 Vdd GND efet
M3762 n_1107 n_1107 Vdd GND efet
M3763 op_T0_and op_T0_and Vdd GND efet
M3764 abl2 abl2 Vdd GND efet
M3765 n_1507 n_1507 Vdd GND efet
M3766 nC01 nC01 Vdd GND efet
M3767 op_T2_abs_y op_T2_abs_y Vdd GND efet
M3768 n_1511 n_1511 Vdd GND efet
M3769 n_1518 n_1518 Vdd GND efet
M3770 n_1517 n_1517 Vdd GND efet
M3771 op_plp_pla op_plp_pla Vdd GND efet
M3772 n_1519 n_1519 Vdd GND efet
M3773 n_1240 n_1240 Vdd GND efet
M3774 n_1231 n_1231 Vdd GND efet
M3775 notalucout notalucout Vdd GND efet
M3776 n_410 n_410 Vdd GND efet
M3777 n_409 n_409 Vdd GND efet
M3778 n_A_B_4 n_A_B_4 Vdd GND efet
M3779 op_T0_ora op_T0_ora Vdd GND efet
M3780 alu0 alu0 Vdd GND efet
M3781 n_400 n_400 Vdd GND efet
M3782 n_397 n_397 Vdd GND efet
M3783 noty1 noty1 Vdd GND efet
M3784 n_1141 n_1141 Vdd GND efet
M3785 n_1145 n_1145 Vdd GND efet
M3786 alucout alucout Vdd GND efet
M3787 n_1153 n_1153 Vdd GND efet
M3788 n_1154 n_1154 Vdd GND efet
M3789 x_op_T__adc_sbc x_op_T__adc_sbc Vdd GND efet
M3790 n_1157 n_1157 Vdd GND efet
M3791 n_108 n_108 Vdd GND efet
M3792 n_109 n_109 Vdd GND efet
M3793 A_B2 A_B2 Vdd GND efet
M3794 n_111 n_111 Vdd GND efet
M3795 n_93 n_93 Vdd GND efet
M3796 dor0 dor0 Vdd GND efet
M3797 n_104 n_104 Vdd GND efet
M3798 n_105 n_105 Vdd GND efet
M3799 npchp1 npchp1 Vdd GND efet
M3800 A_B7 A_B7 Vdd GND efet
M3801 n_889 n_889 Vdd GND efet
M3802 nIRQP nIRQP Vdd GND efet
M3803 n_880 n_880 Vdd GND efet
M3804 fetch fetch Vdd GND efet
M3805 n_877 n_877 Vdd GND efet
M3806 n_876 n_876 Vdd GND efet
M3807 n_885 n_885 Vdd GND efet
M3808 n_AxB_3 n_AxB_3 Vdd GND efet
M3809 n_883 n_883 Vdd GND efet
M3810 n_882 n_882 Vdd GND efet
M3811 A_B6 A_B6 Vdd GND efet
M3812 op_T4_brk_jsr op_T4_brk_jsr Vdd GND efet
M3813 n_797 n_797 Vdd GND efet
M3814 n_800 n_800 Vdd GND efet
M3815 op_push_pull op_push_pull Vdd GND efet
M3816 n_795 n_795 Vdd GND efet
M3817 n_789 n_789 Vdd GND efet
M3818 n_790 n_790 Vdd GND efet
M3819 n_807 n_807 Vdd GND efet
M3820 C78 C78 Vdd GND efet
M3821 n_441 n_441 Vdd GND efet
M3822 n_440 n_440 Vdd GND efet
M3823 dor3 dor3 Vdd GND efet
M3824 n_442 n_442 Vdd GND efet
M3825 op_T5_rti_rts op_T5_rti_rts Vdd GND efet
M3826 n_445 n_445 Vdd GND efet
M3827 dasb2 dasb2 Vdd GND efet
M3828 x_op_T3_abs_idx x_op_T3_abs_idx Vdd GND efet
M3829 n_457 n_457 Vdd GND efet
M3830 n_453 n_453 Vdd GND efet
M3831 n_1159 n_1159 Vdd GND efet
M3832 op_clv op_clv Vdd GND efet
M3833 notalucin notalucin Vdd GND efet
M3834 n_1166 n_1166 Vdd GND efet
M3835 op_T5_ind_y op_T5_ind_y Vdd GND efet
M3836 n_1169 n_1169 Vdd GND efet
M3837 x_op_T0_tya x_op_T0_tya Vdd GND efet
M3838 n_588 n_588 Vdd GND efet
M3839 n_582 n_582 Vdd GND efet
M3840 pclp5 pclp5 Vdd GND efet
M3841 n_75 n_75 Vdd GND efet
M3842 n_70 n_70 Vdd GND efet
M3843 n_71 n_71 Vdd GND efet
M3844 _AxB_4_nC34 _AxB_4_nC34 Vdd GND efet
M3845 Reset0 Reset0 Vdd GND efet
M3846 n_62 n_62 Vdd GND efet
M3847 dor7 dor7 Vdd GND efet
M3848 op_T3_ind_y op_T3_ind_y Vdd GND efet
M3849 n_61 n_61 Vdd GND efet
M3850 n_853 n_853 Vdd GND efet
M3851 n_852 n_852 Vdd GND efet
M3852 n_849 n_849 Vdd GND efet
M3853 n_847 n_847 Vdd GND efet
M3854 nTWOCYCLE nTWOCYCLE Vdd GND efet
M3855 n_850 n_850 Vdd GND efet
M3856 n_844 n_844 Vdd GND efet
M3857 n_842 n_842 Vdd GND efet
M3858 n_846 n_846 Vdd GND efet
M3859 n_845 n_845 Vdd GND efet
M3860 n_1205 n_1205 Vdd GND efet
M3861 n_1195 n_1195 Vdd GND efet
M3862 op_SUMS op_SUMS Vdd GND efet
M3863 n_0_ADL2 n_0_ADL2 Vdd GND efet
M3864 n_1194 n_1194 Vdd GND efet
M3865 DBNeg DBNeg Vdd GND efet
M3866 n_1202 n_1202 Vdd GND efet
M3867 n_AxBxC_6 n_AxBxC_6 Vdd GND efet
M3868 n_1199 n_1199 Vdd GND efet
M3869 n_956 n_956 Vdd GND efet
M3870 n_954 n_954 Vdd GND efet
M3871 n_AxB_1 n_AxB_1 Vdd GND efet
M3872 n_952 n_952 Vdd GND efet
M3873 n_951 n_951 Vdd GND efet
M3874 op_T__cpx_cpy_abs op_T__cpx_cpy_abs Vdd GND efet
M3875 n_947 n_947 Vdd GND efet
M3876 n_946 n_946 Vdd GND efet
M3877 n_959 n_959 Vdd GND efet
M3878 n_958 n_958 Vdd GND efet
M3879 n_587 n_587 Vdd GND efet
M3880 n_571 n_571 Vdd GND efet
M3881 n_572 n_572 Vdd GND efet
M3882 op_T0_adc_sbc op_T0_adc_sbc Vdd GND efet
M3883 n_578 n_578 Vdd GND efet
M3884 op_T3_jsr op_T3_jsr Vdd GND efet
M3885 n_583 n_583 Vdd GND efet
M3886 n_586 n_586 Vdd GND efet
M3887 n_272 n_272 Vdd GND efet
M3888 op_T0_jsr op_T0_jsr Vdd GND efet
M3889 dasb5 dasb5 Vdd GND efet
M3890 n_262 n_262 Vdd GND efet
M3891 n_261 n_261 Vdd GND efet
M3892 n_260 n_260 Vdd GND efet
M3893 n_270 n_270 Vdd GND efet
M3894 n_269 n_269 Vdd GND efet
M3895 n_267 n_267 Vdd GND efet
M3896 nNMIG nNMIG Vdd GND efet
M3897 n_1229 n_1229 Vdd GND efet
M3898 n_1230 n_1230 Vdd GND efet
M3899 n_1225 n_1225 Vdd GND efet
M3900 op_T0_plp op_T0_plp Vdd GND efet
M3901 npclp0 npclp0 Vdd GND efet
M3902 op_ANDS op_ANDS Vdd GND efet
M3903 AxB5 AxB5 Vdd GND efet
M3904 n_1222 n_1222 Vdd GND efet
M3905 n_1223 n_1223 Vdd GND efet
M3906 n_1224 n_1224 Vdd GND efet
M3907 op_xy op_xy Vdd GND efet
M3908 n_1548 n_1548 Vdd GND efet
M3909 n_146 n_146 Vdd GND efet
M3910 n_149 n_149 Vdd GND efet
M3911 n_134 n_134 Vdd GND efet
M3912 n_139 n_139 Vdd GND efet
M3913 n_132 n_132 Vdd GND efet
M3914 n_133 n_133 Vdd GND efet
M3915 n_A_B_0 n_A_B_0 Vdd GND efet
M3916 op_sta_cmp op_sta_cmp Vdd GND efet
M3917 pchp3 pchp3 Vdd GND efet
M3918 C45 C45 Vdd GND efet
M3919 n_929 n_929 Vdd GND efet
M3920 n_928 n_928 Vdd GND efet
M3921 n_917 n_917 Vdd GND efet
M3922 n_916 n_916 Vdd GND efet
M3923 n_919 n_919 Vdd GND efet
M3924 A_B4 A_B4 Vdd GND efet
M3925 n_923 n_923 Vdd GND efet
M3926 n_920 n_920 Vdd GND efet
M3927 C1x5Reset C1x5Reset Vdd GND efet
M3928 nop_store nop_store Vdd GND efet
M3929 n_611 n_611 Vdd GND efet
M3930 n_613 n_613 Vdd GND efet
M3931 n_608 n_608 Vdd GND efet
M3932 n_609 n_609 Vdd GND efet
M3933 n_618 n_618 Vdd GND efet
M3934 n_620 n_620 Vdd GND efet
M3935 n_616 n_616 Vdd GND efet
M3936 n_617 n_617 Vdd GND efet
M3937 DA_C01 DA_C01 Vdd GND efet
M3938 n_624 n_624 Vdd GND efet
M3939 VEC0 VEC0 Vdd GND efet
M3940 op_T0_txs op_T0_txs Vdd GND efet
M3941 op_ror op_ror Vdd GND efet
M3942 n_241 n_241 Vdd GND efet
M3943 idl5 idl5 Vdd GND efet
M3944 n_243 n_243 Vdd GND efet
M3945 n_242 n_242 Vdd GND efet
M3946 abl5 abl5 Vdd GND efet
M3947 n_233 n_233 Vdd GND efet
M3948 n_238 n_238 Vdd GND efet
M3949 n_236 n_236 Vdd GND efet
M3950 n_1256 n_1256 Vdd GND efet
M3951 n_1257 n_1257 Vdd GND efet
M3952 n_1253 n_1253 Vdd GND efet
M3953 n_1255 n_1255 Vdd GND efet
M3954 abl3 abl3 Vdd GND efet
M3955 n_1251 n_1251 Vdd GND efet
M3956 n_1245 n_1245 Vdd GND efet
M3957 op_shift_right op_shift_right Vdd GND efet
M3958 n_1258 n_1258 Vdd GND efet
M3959 op_T4_ind_x op_T4_ind_x Vdd GND efet
M3960 op_SRS op_SRS Vdd GND efet
M3961 dor4 dor4 Vdd GND efet
M3962 n_1709 n_1709 Vdd GND efet
M3963 op_T__cpx_cpy_imm_zp op_T__cpx_cpy_imm_zp Vdd GND efet
M3964 abl0 abl0 Vdd GND efet
M3965 n_1711 n_1711 Vdd GND efet
M3966 n_1712 n_1712 Vdd GND efet
M3967 n_1697 n_1697 Vdd GND efet
M3968 dpc34_PCLC dpc34_PCLC Vdd GND efet
M3969 n_1705 n_1705 Vdd GND efet
M3970 n_1708 n_1708 Vdd GND efet
M3971 C12 C12 Vdd GND efet
M3972 n_506 n_506 Vdd GND efet
M3973 n_507 n_507 Vdd GND efet
M3974 n_510 n_510 Vdd GND efet
M3975 C56 C56 Vdd GND efet
M3976 n_501 n_501 Vdd GND efet
M3977 n_503 n_503 Vdd GND efet
M3978 n_504 n_504 Vdd GND efet
M3979 n_513 n_513 Vdd GND efet
M3980 n_515 n_515 Vdd GND efet
M3981 DA_AB2 DA_AB2 Vdd GND efet
M3982 n_213 n_213 Vdd GND efet
M3983 n_212 n_212 Vdd GND efet
M3984 pchp1 pchp1 Vdd GND efet
M3985 pclp4 pclp4 Vdd GND efet
M3986 n_207 n_207 Vdd GND efet
M3987 n_206 n_206 Vdd GND efet
M3988 op_T2_ADL_ADD op_T2_ADL_ADD Vdd GND efet
M3989 n_218 n_218 Vdd GND efet
M3990 n_0_ADL0 n_0_ADL0 Vdd GND efet
M3991 n_990 n_990 Vdd GND efet
M3992 n_988 n_988 Vdd GND efet
M3993 n_550 n_550 Vdd GND efet
M3994 n_551 n_551 Vdd GND efet
M3995 op_shift op_shift Vdd GND efet
M3996 n_548 n_548 Vdd GND efet
M3997 n_543 n_543 Vdd GND efet
M3998 n_544 n_544 Vdd GND efet
M3999 n_538 n_538 Vdd GND efet
M4000 pd4_clearIR pd4_clearIR Vdd GND efet
M4001 n_533 n_533 Vdd GND efet
M4002 npchp7 npchp7 Vdd GND efet
M4003 noty3 noty3 Vdd GND efet
M4004 n_182 n_182 Vdd GND efet
M4005 n_172 n_172 Vdd GND efet
M4006 n_169 n_169 Vdd GND efet
M4007 n_176 n_176 Vdd GND efet
M4008 _AxB_6_nC56 _AxB_6_nC56 Vdd GND efet
M4009 abl6 abl6 Vdd GND efet
M4010 n_AxB_7 n_AxB_7 Vdd GND efet
M4011 n_180 n_180 Vdd GND efet
M4012 op_T0_txa op_T0_txa Vdd GND efet
M4013 n_1449 n_1449 Vdd GND efet
M4014 dor5 dor5 Vdd GND efet
M4015 notx1 notx1 Vdd GND efet
M4016 noty6 noty6 Vdd GND efet
M4017 n_1440 n_1440 Vdd GND efet
M4018 n_1441 n_1441 Vdd GND efet
M4019 Pout1 Pout1 Vdd GND efet
M4020 n_1446 n_1446 Vdd GND efet
M4021 n_1448 n_1448 Vdd GND efet
M4022 n_1401 n_1401 Vdd GND efet
M4023 n_1402 n_1402 Vdd GND efet
M4024 n_1399 n_1399 Vdd GND efet
M4025 n_1400 n_1400 Vdd GND efet
M4026 n_1412 n_1412 Vdd GND efet
M4027 n_1413 n_1413 Vdd GND efet
M4028 n_1408 n_1408 Vdd GND efet
M4029 pd7_clearIR pd7_clearIR Vdd GND efet
M4030 alu3 alu3 Vdd GND efet
M4031 dor6 dor6 Vdd GND efet
M4032 op_T2 op_T2 Vdd GND efet
M4033 op_T0_sbc op_T0_sbc Vdd GND efet
M4034 n_781 n_781 Vdd GND efet
M4035 n_779 n_779 Vdd GND efet
M4036 ONEBYTE ONEBYTE Vdd GND efet
M4037 op_T5_jsr op_T5_jsr Vdd GND efet
M4038 op_T__dex op_T__dex Vdd GND efet
M4039 op_T5_rti op_T5_rti Vdd GND efet
M4040 n_783 n_783 Vdd GND efet
M4041 n_782 n_782 Vdd GND efet
M4042 n_1117 n_1117 Vdd GND efet
M4043 n_1694 n_1694 Vdd GND efet
M4044 n_A_B_2 n_A_B_2 Vdd GND efet
M4045 op_EORS op_EORS Vdd GND efet
M4046 n_1688 n_1688 Vdd GND efet
M4047 n_1687 n_1687 Vdd GND efet
M4048 n_1684 n_1684 Vdd GND efet
M4049 n_1682 n_1682 Vdd GND efet
M4050 n_1677 n_1677 Vdd GND efet
M4051 n_1676 n_1676 Vdd GND efet
M4052 so so Vdd GND efet
M4053 n_1376 n_1376 Vdd GND efet
M4054 n_1377 n_1377 Vdd GND efet
M4055 n_1379 n_1379 Vdd GND efet
M4056 n_1380 n_1380 Vdd GND efet
M4057 n_1371 n_1371 Vdd GND efet
M4058 DC34 DC34 Vdd GND efet
M4059 NMIL NMIL Vdd GND efet
M4060 n_1375 n_1375 Vdd GND efet
M4061 op_T3_jmp op_T3_jmp Vdd GND efet
M4062 brk_done brk_done Vdd GND efet
M4063 n_763 n_763 Vdd GND efet
M4064 n_762 n_762 Vdd GND efet
M4065 n_755 n_755 Vdd GND efet
M4066 n_754 n_754 Vdd GND efet
M4067 n_761 n_761 Vdd GND efet
M4068 n_757 n_757 Vdd GND efet
M4069 n_748 n_748 Vdd GND efet
M4070 n_747 n_747 Vdd GND efet
M4071 n_753 n_753 Vdd GND efet
M4072 op_T2_php op_T2_php Vdd GND efet
M4073 n_470 n_470 Vdd GND efet
M4074 n_472 n_472 Vdd GND efet
M4075 n_458 n_458 Vdd GND efet
M4076 x_op_T4_ind_y x_op_T4_ind_y Vdd GND efet
M4077 n_462 n_462 Vdd GND efet
M4078 idl3 idl3 Vdd GND efet
M4079 n_465 n_465 Vdd GND efet
M4080 n_466 n_466 Vdd GND efet
M4081 n_467 n_467 Vdd GND efet
M4082 n_468 n_468 Vdd GND efet
M4083 n_1717 n_1717 Vdd GND efet
M4084 n_1716 n_1716 Vdd GND efet
M4085 n_1719 n_1719 Vdd GND efet
M4086 n_1718 n_1718 Vdd GND efet
M4087 op_branch_done op_branch_done Vdd GND efet
M4088 n_1720 n_1720 Vdd GND efet
M4089 n_1724 n_1724 Vdd GND efet
M4090 pchp0 pchp0 Vdd GND efet
M4091 n_658 n_658 Vdd GND efet
M4092 op_T3_branch op_T3_branch Vdd GND efet
M4093 n_647 n_647 Vdd GND efet
M4094 n_A_B_3 n_A_B_3 Vdd GND efet
M4095 n_AxBxC_4 n_AxBxC_4 Vdd GND efet
M4096 pchp6 pchp6 Vdd GND efet
M4097 AxB3 AxB3 Vdd GND efet
M4098 n_641 n_641 Vdd GND efet
M4099 n_645 n_645 Vdd GND efet
M4100 n_646 n_646 Vdd GND efet
M4101 n_1346 n_1346 Vdd GND efet
M4102 n_1347 n_1347 Vdd GND efet
M4103 n_1344 n_1344 Vdd GND efet
M4104 n_1345 n_1345 Vdd GND efet
M4105 op_T0_acc op_T0_acc Vdd GND efet
M4106 n_1343 n_1343 Vdd GND efet
M4107 op_T0_cpx_cpy_inx_iny op_T0_cpx_cpy_inx_iny Vdd GND efet
M4108 n_1339 n_1339 Vdd GND efet
M4109 dpc35_PCHC dpc35_PCHC Vdd GND efet
M4110 n_1335 n_1335 Vdd GND efet
M4111 pclp3 pclp3 Vdd GND efet
M4112 n_721 n_721 Vdd GND efet
M4113 n_720 n_720 Vdd GND efet
M4114 n_718 n_718 Vdd GND efet
M4115 n_717 n_717 Vdd GND efet
M4116 n_715 n_715 Vdd GND efet
M4117 n_714 n_714 Vdd GND efet
M4118 n_726 n_726 Vdd GND efet
M4119 dpc22_nDSA dpc22_nDSA Vdd GND efet
M4120 n_355 n_355 Vdd GND efet
M4121 dasb1 dasb1 Vdd GND efet
M4122 n_1007 n_1007 Vdd GND efet
M4123 abh6 abh6 Vdd GND efet
M4124 irline3 irline3 Vdd GND efet
M4125 n_995 n_995 Vdd GND efet
M4126 n_992 n_992 Vdd GND efet
M4127 op_implied op_implied Vdd GND efet
M4128 nC23 nC23 Vdd GND efet
M4129 n_1002 n_1002 Vdd GND efet
M4130 n_998 n_998 Vdd GND efet
M4131 abh2 abh2 Vdd GND efet
M4132 op_T0_tay_ldy_not_idx op_T0_tay_ldy_not_idx Vdd GND efet
M4133 n_291 n_291 Vdd GND efet
M4134 n_288 n_288 Vdd GND efet
M4135 n_AxB1__C01 n_AxB1__C01 Vdd GND efet
M4136 n_293 n_293 Vdd GND efet
M4137 n_299 n_299 Vdd GND efet
M4138 nNMIP nNMIP Vdd GND efet
M4139 op_T__cmp op_T__cmp Vdd GND efet
M4140 n_300 n_300 Vdd GND efet
M4141 n_1649 n_1649 Vdd GND efet
M4142 n_1650 n_1650 Vdd GND efet
M4143 op_T__bit op_T__bit Vdd GND efet
M4144 pclp7 pclp7 Vdd GND efet
M4145 n_1642 n_1642 Vdd GND efet
M4146 n_1643 n_1643 Vdd GND efet
M4147 noty7 noty7 Vdd GND efet
M4148 n_1641 n_1641 Vdd GND efet
M4149 alu2 alu2 Vdd GND efet
M4150 n_1638 n_1638 Vdd GND efet
M4151 A_B0 A_B0 Vdd GND efet
M4152 n_692 n_692 Vdd GND efet
M4153 nA_B2 nA_B2 Vdd GND efet
M4154 dasb6 dasb6 Vdd GND efet
M4155 n_0_ADL1 n_0_ADL1 Vdd GND efet
M4156 op_T0_tsx op_T0_tsx Vdd GND efet
M4157 n_689 n_689 Vdd GND efet
M4158 Pout0 Pout0 Vdd GND efet
M4159 op_asl_rol op_asl_rol Vdd GND efet
M4160 _t4 _t4 Vdd GND efet
M4161 C67 C67 Vdd GND efet
M4162 A_B3 A_B3 Vdd GND efet
M4163 idl4 idl4 Vdd GND efet
M4164 n_1305 n_1305 Vdd GND efet
M4165 n_1304 n_1304 Vdd GND efet
M4166 n_1303 n_1303 Vdd GND efet
M4167 n_1312 n_1312 Vdd GND efet
M4168 op_T4_rti op_T4_rti Vdd GND efet
M4169 n_1309 n_1309 Vdd GND efet
M4170 notaluvout notaluvout Vdd GND efet
M4171 H1x1 H1x1 Vdd GND efet
M4172 nDBE nDBE Vdd GND efet
M4173 n_1034 n_1034 Vdd GND efet
M4174 n_1038 n_1038 Vdd GND efet
M4175 n_1037 n_1037 Vdd GND efet
M4176 op_T3_stack_bit_jmp op_T3_stack_bit_jmp Vdd GND efet
M4177 n_1028 n_1028 Vdd GND efet
M4178 n_1033 n_1033 Vdd GND efet
M4179 NMIP NMIP Vdd GND efet
M4180 n_1599 n_1599 Vdd GND efet
M4181 n_1600 n_1600 Vdd GND efet
M4182 op_sty_cpy_mem op_sty_cpy_mem Vdd GND efet
M4183 n_1605 n_1605 Vdd GND efet
M4184 n_1610 n_1610 Vdd GND efet
M4185 op_T4_rts op_T4_rts Vdd GND efet
M4186 n_1613 n_1613 Vdd GND efet
M4187 n_1614 n_1614 Vdd GND efet
M4188 n_1618 n_1618 Vdd GND efet
M4189 n_1619 n_1619 Vdd GND efet
M4190 n_1070 n_1070 Vdd GND efet
M4191 n_1069 n_1069 Vdd GND efet
M4192 n_1067 n_1067 Vdd GND efet
M4193 idl2 idl2 Vdd GND efet
M4194 n_1065 n_1065 Vdd GND efet
M4195 nA_B4 nA_B4 Vdd GND efet
M4196 op_T2_abs op_T2_abs Vdd GND efet
M4197 n_1056 n_1056 Vdd GND efet
M4198 op_T0_shift_right_a op_T0_shift_right_a Vdd GND efet
M4199 n_1073 n_1073 Vdd GND efet
M4200 op_T2_stack op_T2_stack Vdd GND efet
M4201 n_1585 n_1585 Vdd GND efet
M4202 nC45 nC45 Vdd GND efet
M4203 n_1573 n_1573 Vdd GND efet
M4204 _t3 _t3 Vdd GND efet
M4205 x_op_T4_rti x_op_T4_rti Vdd GND efet
M4206 n_1578 n_1578 Vdd GND efet
M4207 n_1580 n_1580 Vdd GND efet
M4208 n_1575 n_1575 Vdd GND efet
M4209 ir3 ir3 Vdd GND efet
M4210 op_T3_abs_idx op_T3_abs_idx Vdd GND efet
M4211 op_lsr_ror_dec_inc op_lsr_ror_dec_inc Vdd GND efet
M4212 n_35 n_35 Vdd GND efet
M4213 n_34 n_34 Vdd GND efet
M4214 npchp5 npchp5 Vdd GND efet
M4215 n_31 n_31 Vdd GND efet
M4216 n_46 n_46 Vdd GND efet
M4217 npclp4 npclp4 Vdd GND efet
M4218 n_38 n_38 Vdd GND efet
M4219 n_36 n_36 Vdd GND efet
M4220 abh1 abh1 Vdd GND efet
M4221 n_420 n_420 Vdd GND efet
M4222 n_419 n_419 Vdd GND efet
M4223 n_318 n_318 Vdd GND efet
M4224 n_319 n_319 Vdd GND efet
M4225 n_320 n_320 Vdd GND efet
M4226 n_321 n_321 Vdd GND efet
M4227 op_inc_nop op_inc_nop Vdd GND efet
M4228 n_326 n_326 Vdd GND efet
M4229 n_327 n_327 Vdd GND efet
M4230 ir0 ir0 Vdd GND efet
M4231 n_329 n_329 Vdd GND efet
M4232 n_330 n_330 Vdd GND efet
M4233 n_1101 n_1101 Vdd GND efet
M4234 n_1099 n_1099 Vdd GND efet
M4235 n_1089 n_1089 Vdd GND efet
M4236 n_1091 n_1091 Vdd GND efet
M4237 n_1090 n_1090 Vdd GND efet
M4238 n_1094 n_1094 Vdd GND efet
M4239 n_1093 n_1093 Vdd GND efet
M4240 n_1097 n_1097 Vdd GND efet
M4241 n_1541 n_1541 Vdd GND efet
M4242 n_1542 n_1542 Vdd GND efet
M4243 n_1526 n_1526 Vdd GND efet
M4244 n_1531 n_1531 Vdd GND efet
M4245 n_1534 n_1534 Vdd GND efet
M4246 op_from_x op_from_x Vdd GND efet
M4247 notx3 notx3 Vdd GND efet
M4248 n_1523 n_1523 Vdd GND efet
M4249 op_T2_ind op_T2_ind Vdd GND efet
M4250 n_AxB_0 n_AxB_0 Vdd GND efet
M4251 n_16 n_16 Vdd GND efet
M4252 n_14 n_14 Vdd GND efet
M4253 n_8 n_8 Vdd GND efet
M4254 n_6 n_6 Vdd GND efet
M4255 n_11 n_11 Vdd GND efet
M4256 n_10 n_10 Vdd GND efet
M4257 n_3 n_3 Vdd GND efet
M4258 op_T5_rts op_T5_rts Vdd GND efet
M4259 n_5 n_5 Vdd GND efet
M4260 op_T0_tay op_T0_tay Vdd GND efet
M4261 VEC1 VEC1 Vdd GND efet
M4262 op_T__iny_dey op_T__iny_dey Vdd GND efet
M4263 x_op_T0_bit x_op_T0_bit Vdd GND efet
M4264 op_T0_brk_rti op_T0_brk_rti Vdd GND efet
M4265 n_1474 n_1474 Vdd GND efet
M4266 dasb3 dasb3 Vdd GND efet
M4267 n_AxB_5 n_AxB_5 Vdd GND efet
M4268 n_1471 n_1471 Vdd GND efet
M4269 noty2 noty2 Vdd GND efet
M4270 n_1486 n_1486 Vdd GND efet
M4271 abh4 abh4 Vdd GND efet
M4272 n_358 n_358 Vdd GND efet
M4273 PD_0xx0xx0x PD_0xx0xx0x Vdd GND efet
M4274 n_347 n_347 Vdd GND efet
M4275 nA_B3 nA_B3 Vdd GND efet
M4276 n_344 n_344 Vdd GND efet
M4277 n_345 n_345 Vdd GND efet
M4278 op_T4_abs_idx op_T4_abs_idx Vdd GND efet
M4279 n_351 n_351 Vdd GND efet
M4280 op_T4_brk op_T4_brk Vdd GND efet
M4281 notir3 notir3 Vdd GND efet
M4282 nC12 nC12 Vdd GND efet
M4283 n_1120 n_1120 Vdd GND efet
M4284 p4 p4 Vdd GND efet
M4285 nVEC nVEC Vdd GND efet
M4286 n_1133 n_1133 Vdd GND efet
M4287 n_1130 n_1130 Vdd GND efet
M4288 n_1129 n_1129 Vdd GND efet
M4289 n_1137 n_1137 Vdd GND efet
M4290 n_1135 n_1135 Vdd GND efet
M4291 n_1654 n_1654 Vdd GND efet
M4292 pchp2 pchp2 Vdd GND efet
M4293 n_1497 n_1497 Vdd GND efet
M4294 dasb7 dasb7 Vdd GND efet
M4295 n_1495 n_1495 Vdd GND efet
M4296 n_1491 n_1491 Vdd GND efet
M4297 n_1492 n_1492 Vdd GND efet
M4298 op_T3_plp_pla op_T3_plp_pla Vdd GND efet
M4299 n_1488 n_1488 Vdd GND efet
M4300 n_1499 n_1499 Vdd GND efet
M4301 n_1500 n_1500 Vdd GND efet
M4302 n_128 n_128 Vdd GND efet
M4303 n_127 n_127 Vdd GND efet
M4304 PD_n_0xx0xx0x PD_n_0xx0xx0x Vdd GND efet
M4305 npchp3 npchp3 Vdd GND efet
M4306 n_123 n_123 Vdd GND efet
M4307 n_122 n_122 Vdd GND efet
M4308 op_T3 op_T3 Vdd GND efet
M4309 n_118 n_118 Vdd GND efet
M4310 op_T0_pla op_T0_pla Vdd GND efet
M4311 n_130 n_130 Vdd GND efet
M4312 n_810 n_810 Vdd GND efet
M4313 pd1_clearIR pd1_clearIR Vdd GND efet
M4314 n_812 n_812 Vdd GND efet
M4315 n_811 n_811 Vdd GND efet
M4316 n_815 n_815 Vdd GND efet
M4317 n_813 n_813 Vdd GND efet
M4318 n_818 n_818 Vdd GND efet
M4319 n_AxB5__C45 n_AxB5__C45 Vdd GND efet
M4320 op_T__adc_sbc op_T__adc_sbc Vdd GND efet
M4321 n_819 n_819 Vdd GND efet
M4322 n_392 n_392 Vdd GND efet
M4323 n_396 n_396 Vdd GND efet
M4324 n_388 n_388 Vdd GND efet
M4325 n_389 n_389 Vdd GND efet
M4326 n_390 n_390 Vdd GND efet
M4327 idl7 idl7 Vdd GND efet
M4328 n_383 n_383 Vdd GND efet
M4329 n_384 n_384 Vdd GND efet
M4330 n_385 n_385 Vdd GND efet
M4331 n_386 n_386 Vdd GND efet
M4332 n_1181 n_1181 Vdd GND efet
M4333 n_1180 n_1180 Vdd GND efet
M4334 n_1179 n_1179 Vdd GND efet
M4335 n_1178 n_1178 Vdd GND efet
M4336 n_1184 n_1184 Vdd GND efet
M4337 notir2 notir2 Vdd GND efet
M4338 n_91 n_91 Vdd GND efet
M4339 n_90 n_90 Vdd GND efet
M4340 p6 p6 Vdd GND efet
M4341 op_T0_dex op_T0_dex Vdd GND efet
M4342 n_79 n_79 Vdd GND efet
M4343 C34 C34 Vdd GND efet
M4344 n_83 n_83 Vdd GND efet
M4345 n_80 n_80 Vdd GND efet
M4346 rdy rdy Vdd GND efet
M4347 op_T2_ind_x op_T2_ind_x Vdd GND efet
M4348 alu1 alu1 Vdd GND efet
M4349 n_875 n_875 Vdd GND efet
M4350 n_854 n_854 Vdd GND efet
M4351 op_rti_rts op_rti_rts Vdd GND efet
M4352 n_AxB3__C23 n_AxB3__C23 Vdd GND efet
M4353 n_861 n_861 Vdd GND efet
M4354 n_862 n_862 Vdd GND efet
M4355 n_867 n_867 Vdd GND efet
M4356 idl1 idl1 Vdd GND efet
M4357 n_871 n_871 Vdd GND efet
M4358 n_432 n_432 Vdd GND efet
M4359 op_rmw op_rmw Vdd GND efet
M4360 nC56 nC56 Vdd GND efet
M4361 n_424 n_424 Vdd GND efet
M4362 AxB1 AxB1 Vdd GND efet
M4363 abh3 abh3 Vdd GND efet
M4364 n_423 n_423 Vdd GND efet
M4365 n_436 n_436 Vdd GND efet
M4366 n_1211 n_1211 Vdd GND efet
M4367 op_T5_ind_x op_T5_ind_x Vdd GND efet
M4368 n_1219 n_1219 Vdd GND efet
M4369 n_1218 n_1218 Vdd GND efet
M4370 n_1187 n_1187 Vdd GND efet
M4371 short_circuit_idx_add short_circuit_idx_add Vdd GND efet
M4372 n_1192 n_1192 Vdd GND efet
M4373 n_1190 n_1190 Vdd GND efet
M4374 n_830 n_830 Vdd GND efet
M4375 n_831 n_831 Vdd GND efet
M4376 n_824 n_824 Vdd GND efet
M4377 D1x1 D1x1 Vdd GND efet
M4378 n_838 n_838 Vdd GND efet
M4379 n_839 n_839 Vdd GND efet
M4380 n_834 n_834 Vdd GND efet
M4381 n_837 n_837 Vdd GND efet
M4382 nop_branch_bit6 nop_branch_bit6 Vdd GND efet
M4383 nA_B1 nA_B1 Vdd GND efet
M4384 n_570 n_570 Vdd GND efet
M4385 n_568 n_568 Vdd GND efet
M4386 n_556 n_556 Vdd GND efet
M4387 _AxB_0_nC0in _AxB_0_nC0in Vdd GND efet
M4388 n_553 n_553 Vdd GND efet
M4389 op_T0_php_pha op_T0_php_pha Vdd GND efet
M4390 abl7 abl7 Vdd GND efet
M4391 n_566 n_566 Vdd GND efet
M4392 noty4 noty4 Vdd GND efet
M4393 n_564 n_564 Vdd GND efet
M4394 n_1244 n_1244 Vdd GND efet
M4395 op_T__ora_and_eor_adc op_T__ora_and_eor_adc Vdd GND efet
M4396 AxB7 AxB7 Vdd GND efet
M4397 op_T2_branch op_T2_branch Vdd GND efet
M4398 n_1238 n_1238 Vdd GND efet
M4399 A_B5 A_B5 Vdd GND efet
M4400 op_T0_cpy_iny op_T0_cpy_iny Vdd GND efet
M4401 abl4 abl4 Vdd GND efet
M4402 n_160 n_160 Vdd GND efet
M4403 op_T2_stack_access op_T2_stack_access Vdd GND efet
M4404 n_163 n_163 Vdd GND efet
M4405 n_161 n_161 Vdd GND efet
M4406 n_154 n_154 Vdd GND efet
M4407 n_152 n_152 Vdd GND efet
M4408 clock2 clock2 Vdd GND efet
M4409 n_A_B_1 n_A_B_1 Vdd GND efet
M4410 n_168 n_168 Vdd GND efet
M4411 op_T0_tax op_T0_tax Vdd GND efet
M4412 n_935 n_935 Vdd GND efet
M4413 n_936 n_936 Vdd GND efet
M4414 n_937 n_937 Vdd GND efet
M4415 n_930 n_930 Vdd GND efet
M4416 n_931 n_931 Vdd GND efet
M4417 op_T2_php_pha op_T2_php_pha Vdd GND efet
M4418 n_933 n_933 Vdd GND efet
M4419 aluvout aluvout Vdd GND efet
M4420 n_944 n_944 Vdd GND efet
M4421 n_1039 n_1039 Vdd GND efet
M4422 n_1018 n_1018 Vdd GND efet
M4423 op_T3_mem_abs op_T3_mem_abs Vdd GND efet
M4424 alu4 alu4 Vdd GND efet
M4425 n_602 n_602 Vdd GND efet
M4426 n_600 n_600 Vdd GND efet
M4427 n_604 n_604 Vdd GND efet
M4428 n_603 n_603 Vdd GND efet
M4429 n_593 n_593 Vdd GND efet
M4430 nC67 nC67 Vdd GND efet
M4431 n_595 n_595 Vdd GND efet
M4432 op_T0_jmp op_T0_jmp Vdd GND efet
M4433 n_284 n_284 Vdd GND efet
M4434 op_T2_zp_zp_idx op_T2_zp_zp_idx Vdd GND efet
M4435 op_T2_abs_access op_T2_abs_access Vdd GND efet
M4436 n_AxBxC_3 n_AxBxC_3 Vdd GND efet
M4437 n_275 n_275 Vdd GND efet
M4438 n_278 n_278 Vdd GND efet
M4439 n_279 n_279 Vdd GND efet
M4440 n_280 n_280 Vdd GND efet
M4441 op_T4_mem_abs_idx op_T4_mem_abs_idx Vdd GND efet
M4442 n_282 n_282 Vdd GND efet
M4443 n_1262 n_1262 Vdd GND efet
M4444 n_1260 n_1260 Vdd GND efet
M4445 n_1267 n_1267 Vdd GND efet
M4446 n_1265 n_1265 Vdd GND efet
M4447 n_1270 n_1270 Vdd GND efet
M4448 nDBZ nDBZ Vdd GND efet
M4449 op_T0 op_T0 Vdd GND efet
M4450 n_1271 n_1271 Vdd GND efet
M4451 n_1277 n_1277 Vdd GND efet
M4452 n_1275 n_1275 Vdd GND efet
M4453 alucin alucin Vdd GND efet
M4454 n_913 n_913 Vdd GND efet
M4455 n_906 n_906 Vdd GND efet
M4456 _t5 _t5 Vdd GND efet
M4457 op_T3_mem_zp_idx op_T3_mem_zp_idx Vdd GND efet
M4458 n_905 n_905 Vdd GND efet
M4459 n_896 n_896 Vdd GND efet
M4460 nDA_ADD1 nDA_ADD1 Vdd GND efet
M4461 notx2 notx2 Vdd GND efet
M4462 notir6 notir6 Vdd GND efet
M4463 notx0 notx0 Vdd GND efet
M4464 n_986 n_986 Vdd GND efet
M4465 pclp1 pclp1 Vdd GND efet
M4466 n_980 n_980 Vdd GND efet
M4467 n_494 n_494 Vdd GND efet
M4468 op_T4_ind_y op_T4_ind_y Vdd GND efet
M4469 n_491 n_491 Vdd GND efet
M4470 n_490 n_490 Vdd GND efet
M4471 abh7 abh7 Vdd GND efet
M4472 pclp0 pclp0 Vdd GND efet
M4473 op_T2_brk op_T2_brk Vdd GND efet
M4474 n_AxBxC_5 n_AxBxC_5 Vdd GND efet
M4475 n_499 n_499 Vdd GND efet
M4476 n_496 n_496 Vdd GND efet
M4477 nop_set_C nop_set_C Vdd GND efet
M4478 n_253 n_253 Vdd GND efet
M4479 n_249 n_249 Vdd GND efet
M4480 n_251 n_251 Vdd GND efet
M4481 n_256 n_256 Vdd GND efet
M4482 op_T0_tya op_T0_tya Vdd GND efet
M4483 n_254 n_254 Vdd GND efet
M4484 n_255 n_255 Vdd GND efet
M4485 op_T2_idx_x_xy op_T2_idx_x_xy Vdd GND efet
M4486 op_jsr op_jsr Vdd GND efet
M4487 op_T0_ldx_tax_tsx op_T0_ldx_tax_tsx Vdd GND efet
M4488 n_983 n_983 Vdd GND efet
M4489 n_979 n_979 Vdd GND efet
M4490 noty5 noty5 Vdd GND efet
M4491 n_1170 n_1170 Vdd GND efet
M4492 nop_branch_bit7 nop_branch_bit7 Vdd GND efet
M4493 n_1175 n_1175 Vdd GND efet
M4494 DA_C45 DA_C45 Vdd GND efet
M4495 n_AxBxC_7 n_AxBxC_7 Vdd GND efet
M4496 n_531 n_531 Vdd GND efet
M4497 op_store op_store Vdd GND efet
M4498 DA_AxB2 DA_AxB2 Vdd GND efet
M4499 n_519 n_519 Vdd GND efet
M4500 n_518 n_518 Vdd GND efet
M4501 n_523 n_523 Vdd GND efet
M4502 op_ORS op_ORS Vdd GND efet
M4503 xx_op_T5_jsr xx_op_T5_jsr Vdd GND efet
M4504 n_525 n_525 Vdd GND efet
M4505 n_1215 n_1215 Vdd GND efet
M4506 n_1209 n_1209 Vdd GND efet
M4507 pchp7 pchp7 Vdd GND efet
M4508 n_225 n_225 Vdd GND efet
M4509 n_227 n_227 Vdd GND efet
M4510 n_228 n_228 Vdd GND efet
M4511 dpc28_0ADH0 dpc28_0ADH0 Vdd GND efet
M4512 op_T2_mem_zp op_T2_mem_zp Vdd GND efet
M4513 n_220 n_220 Vdd GND efet
M4514 n_221 n_221 Vdd GND efet
M4515 n_224 n_224 Vdd GND efet
M4516 n_231 n_231 Vdd GND efet
M4517 n_232 n_232 Vdd GND efet
M4518 x_op_T3_plp_pla x_op_T3_plp_pla Vdd GND efet
M4519 abh0 abh0 Vdd GND efet
M4520 Pout2 Pout2 Vdd GND efet
M4521 op_T0_lda op_T0_lda Vdd GND efet
M4522 op_T0_cld_sed op_T0_cld_sed Vdd GND efet
M4523 n_1416 n_1416 Vdd GND efet
M4524 op_T3_ind_x op_T3_ind_x Vdd GND efet
M4525 n_1427 n_1427 Vdd GND efet
M4526 nC34 nC34 Vdd GND efet
M4527 n_1423 n_1423 Vdd GND efet
