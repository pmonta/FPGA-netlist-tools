`include "common.h"

module chip_4004(
  input eclk, ereset,
  input clk1,
  input clk2,
  output sync,
  input reset,
  input test,
  input d0_i,
  output d0_o,
  output d0_t,
  input d1_i,
  output d1_o,
  output d1_t,
  input d2_i,
  output d2_o,
  output d2_t,
  input d3_i,
  output d3_o,
  output d3_t,
  output cm_rom,
  output cm_ram3,
  output cm_ram2,
  output cm_ram1,
  output cm_ram0
);

  function v;   // convert an analog node value to 2-level
  input [`W-1:0] x;
  begin
    v = ~x[`W-1];
  end
  endfunction

  function [`W-1:0] a;   // convert a 2-level node value to analog
  input x;
  begin
    a = x ? `HI2 : `LO2;
  end
  endfunction

  wire signed [`W-1:0] N0556_port_2, N0556_port_1, N0556_v;
  wire signed [`W-1:0] S00819_port_0, S00819_v;
  wire signed [`W-1:0] CY_ADA_port_2, CY_ADA_port_3, CY_ADA_port_0, CY_ADA_v;
  wire signed [`W-1:0] N0449_port_3, N0449_port_1, N0449_port_6, N0449_port_4, N0449_port_5, N0449_v;
  wire signed [`W-1:0] N0448_port_2, N0448_port_3, N0448_port_0, N0448_port_1, N0448_v;
  wire signed [`W-1:0] N0443_port_2, N0443_port_1, N0443_v;
  wire signed [`W-1:0] N0442_port_0, N0442_port_1, N0442_v;
  wire signed [`W-1:0] N0441_port_0, N0441_port_1, N0441_v;
  wire signed [`W-1:0] N0440_port_3, N0440_port_4, N0440_port_5, N0440_v;
  wire signed [`W-1:0] N0447_port_2, N0447_port_3, N0447_port_1, N0447_v;
  wire signed [`W-1:0] N0446_port_2, N0446_port_3, N0446_v;
  wire signed [`W-1:0] N0445_port_2, N0445_port_1, N0445_v;
  wire signed [`W-1:0] N0444_port_12, N0444_port_13, N0444_v;
  wire signed [`W-1:0] N0991_port_0, N0991_port_1, N0991_v;
  wire signed [`W-1:0] N0990_port_0, N0990_port_1, N0990_v;
  wire signed [`W-1:0] N0993_port_2, N0993_port_3, N0993_v;
  wire signed [`W-1:0] N0992_port_2, N0992_port_3, N0992_v;
  wire signed [`W-1:0] N0995_port_2, N0995_port_3, N0995_v;
  wire signed [`W-1:0] N0994_port_2, N0994_port_3, N0994_v;
  wire signed [`W-1:0] N0997_port_3, N0997_port_1, N0997_v;
  wire signed [`W-1:0] N0999_port_2, N0999_port_3, N0999_v;
  wire signed [`W-1:0] N0998_port_0, N0998_port_1, N0998_v;
  wire signed [`W-1:0] N0883_port_8, N0883_port_9, N0883_port_2, N0883_port_3, N0883_port_0, N0883_port_6, N0883_port_7, N0883_port_4, N0883_port_5, N0883_port_10, N0883_v;
  wire signed [`W-1:0] N0880_port_8, N0880_port_9, N0880_port_2, N0880_port_3, N0880_port_0, N0880_port_6, N0880_port_7, N0880_port_4, N0880_port_5, N0880_port_10, N0880_v;
  wire signed [`W-1:0] N0887_port_3, N0887_port_5, N0887_v;
  wire signed [`W-1:0] N0886_port_0, N0886_port_1, N0886_v;
  wire signed [`W-1:0] N0530_port_3, N0530_port_4, N0530_v;
  wire signed [`W-1:0] N0536_port_8, N0536_port_9, N0536_port_2, N0536_port_3, N0536_port_0, N0536_port_1, N0536_port_6, N0536_port_7, N0536_port_4, N0536_port_5, N0536_port_10, N0536_v;
  wire signed [`W-1:0] N0535_port_8, N0535_port_9, N0535_port_2, N0535_port_3, N0535_port_0, N0535_port_1, N0535_port_6, N0535_port_7, N0535_port_4, N0535_port_5, N0535_port_10, N0535_v;
  wire signed [`W-1:0] N0534_port_8, N0534_port_9, N0534_port_2, N0534_port_3, N0534_port_0, N0534_port_1, N0534_port_6, N0534_port_7, N0534_port_4, N0534_port_5, N0534_port_10, N0534_v;
  wire signed [`W-1:0] N0539_port_2, N0539_port_3, N0539_port_0, N0539_port_1, N0539_v;
  wire signed [`W-1:0] N0538_port_8, N0538_port_9, N0538_port_2, N0538_port_3, N0538_port_0, N0538_port_1, N0538_port_6, N0538_port_7, N0538_port_4, N0538_port_5, N0538_port_10, N0538_v;
  wire signed [`W-1:0] S00579_port_1, S00579_v;
  wire signed [`W-1:0] S00578_port_1, S00578_v;
  wire signed [`W-1:0] N0939_port_3, N0939_port_4, N0939_v;
  wire signed [`W-1:0] N0418_port_0, N0418_port_1, N0418_v;
  wire signed [`W-1:0] S00757_port_1, S00757_v;
  wire signed [`W-1:0] N0528_port_0, N0528_port_1, N0528_v;
  wire signed [`W-1:0] INC_ISZ_port_2, INC_ISZ_port_3, INC_ISZ_port_0, INC_ISZ_port_1, INC_ISZ_port_4, INC_ISZ_v;
  wire signed [`W-1:0] LD_port_2, LD_port_3, LD_port_0, LD_port_1, LD_port_4, LD_v;
  wire signed [`W-1:0] N0331_port_2, N0331_port_0, N0331_port_1, N0331_v;
  wire signed [`W-1:0] S00817_port_0, S00817_v;
  wire signed [`W-1:0] N0330_port_0, N0330_port_1, N0330_v;
  wire signed [`W-1:0] SUB_GROUP_6__port_2, SUB_GROUP_6__port_3, SUB_GROUP_6__port_0, SUB_GROUP_6__port_1, SUB_GROUP_6__port_6, SUB_GROUP_6__v;
  wire signed [`W-1:0] N0525_port_0, N0525_port_1, N0525_v;
  wire signed [`W-1:0] INC_ISZ_XCH_port_2, INC_ISZ_XCH_port_3, INC_ISZ_XCH_port_1, INC_ISZ_XCH_port_4, INC_ISZ_XCH_port_5, INC_ISZ_XCH_v;
  wire signed [`W-1:0] R8_3_port_1, R8_3_v;
  wire signed [`W-1:0] R8_2_port_0, R8_2_v;
  wire signed [`W-1:0] R8_1_port_1, R8_1_v;
  wire signed [`W-1:0] R8_0_port_0, R8_0_v;
  wire signed [`W-1:0] N0668_port_3, N0668_port_0, N0668_port_4, N0668_v;
  wire signed [`W-1:0] N0332_port_2, N0332_port_0, N0332_port_1, N0332_port_5, N0332_v;
  wire signed [`W-1:0] N0527_port_0, N0527_port_1, N0527_v;
  wire signed [`W-1:0] N0335_port_0, N0335_port_1, N0335_v;
  wire signed [`W-1:0] _TMP_1_port_2, _TMP_1_port_0, _TMP_1_port_1, _TMP_1_v;
  wire signed [`W-1:0] _TMP_0_port_2, _TMP_0_port_0, _TMP_0_port_1, _TMP_0_v;
  wire signed [`W-1:0] _TMP_3_port_2, _TMP_3_port_0, _TMP_3_port_1, _TMP_3_v;
  wire signed [`W-1:0] _TMP_2_port_2, _TMP_2_port_0, _TMP_2_port_1, _TMP_2_v;
  wire signed [`W-1:0] N0337_port_2, N0337_port_0, N0337_port_1, N0337_v;
  wire signed [`W-1:0] TMP_3_port_2, TMP_3_port_0, TMP_3_port_1, TMP_3_v;
  wire signed [`W-1:0] TMP_2_port_2, TMP_2_port_0, TMP_2_port_1, TMP_2_v;
  wire signed [`W-1:0] TMP_1_port_2, TMP_1_port_0, TMP_1_port_1, TMP_1_v;
  wire signed [`W-1:0] TMP_0_port_2, TMP_0_port_0, TMP_0_port_1, TMP_0_v;
  wire signed [`W-1:0] JIN_FIN_port_8, JIN_FIN_port_6, JIN_FIN_port_7, JIN_FIN_port_4, JIN_FIN_port_5, JIN_FIN_v;
  wire signed [`W-1:0] N0336_port_0, N0336_port_1, N0336_v;
  wire signed [`W-1:0] N0523_port_2, N0523_port_3, N0523_port_0, N0523_port_1, N0523_v;
  wire signed [`W-1:0] N0454_port_0, N0454_v;
  wire signed [`W-1:0] N0455_port_3, N0455_port_6, N0455_port_4, N0455_v;
  wire signed [`W-1:0] N0456_port_0, N0456_port_1, N0456_v;
  wire signed [`W-1:0] N0457_port_2, N0457_port_0, N0457_port_1, N0457_v;
  wire signed [`W-1:0] N0450_port_2, N0450_port_0, N0450_v;
  wire signed [`W-1:0] N0451_port_2, N0451_port_0, N0451_v;
  wire signed [`W-1:0] N0452_port_1, N0452_v;
  wire signed [`W-1:0] N0453_port_2, N0453_port_0, N0453_port_1, N0453_v;
  wire signed [`W-1:0] N0458_port_0, N0458_v;
  wire signed [`W-1:0] N0459_port_6, N0459_port_4, N0459_port_5, N0459_v;
  wire signed [`W-1:0] JCN_ISZ_port_8, JCN_ISZ_port_3, JCN_ISZ_port_6, JCN_ISZ_port_7, JCN_ISZ_port_5, JCN_ISZ_v;
  wire signed [`W-1:0] R3_0_port_1, R3_0_v;
  wire signed [`W-1:0] R3_1_port_0, R3_1_v;
  wire signed [`W-1:0] R3_3_port_0, R3_3_v;
  wire signed [`W-1:0] LDM_BBL_port_2, LDM_BBL_port_3, LDM_BBL_port_0, LDM_BBL_port_1, LDM_BBL_v;
  wire signed [`W-1:0] N0982_port_0, N0982_port_1, N0982_v;
  wire signed [`W-1:0] N0983_port_2, N0983_port_3, N0983_v;
  wire signed [`W-1:0] N0980_port_0, N0980_port_1, N0980_v;
  wire signed [`W-1:0] N0981_port_0, N0981_port_1, N0981_v;
  wire signed [`W-1:0] N0986_port_0, N0986_port_1, N0986_v;
  wire signed [`W-1:0] N0987_port_0, N0987_port_1, N0987_v;
  wire signed [`W-1:0] N0984_port_0, N0984_port_1, N0984_v;
  wire signed [`W-1:0] N0985_port_0, N0985_port_1, N0985_v;
  wire signed [`W-1:0] R1_2_port_1, R1_2_v;
  wire signed [`W-1:0] R1_3_port_0, R1_3_v;
  wire signed [`W-1:0] N0988_port_0, N0988_port_1, N0988_v;
  wire signed [`W-1:0] N0989_port_0, N0989_port_1, N0989_v;
  wire signed [`W-1:0] N0366_port_2, N0366_port_3, N0366_port_0, N0366_port_1, N0366_port_6, N0366_port_4, N0366_port_5, N0366_v;
  wire signed [`W-1:0] RRAB0_port_6, RRAB0_port_7, RRAB0_port_4, RRAB0_port_5, RRAB0_v;
  wire signed [`W-1:0] RRAB1_port_6, RRAB1_port_7, RRAB1_port_4, RRAB1_port_5, RRAB1_v;
  wire signed [`W-1:0] N0872_port_3, N0872_port_0, N0872_port_5, N0872_v;
  wire signed [`W-1:0] R7_0_port_1, R7_0_v;
  wire signed [`W-1:0] R7_1_port_0, R7_1_v;
  wire signed [`W-1:0] R7_2_port_1, R7_2_v;
  wire signed [`W-1:0] R7_3_port_0, R7_3_v;
  wire signed [`W-1:0] S00699_port_1, S00699_v;
  wire signed [`W-1:0] N0902_port_2, N0902_port_3, N0902_v;
  wire signed [`W-1:0] R5_2_port_1, R5_2_v;
  wire signed [`W-1:0] R5_0_port_1, R5_0_v;
  wire signed [`W-1:0] N0524_port_2, N0524_port_3, N0524_port_1, N0524_port_4, N0524_v;
  wire signed [`W-1:0] N0526_port_2, N0526_port_0, N0526_port_1, N0526_v;
  wire signed [`W-1:0] N0522_port_2, N0522_port_1, N0522_v;
  wire signed [`W-1:0] BBL_port_2, BBL_port_3, BBL_port_1, BBL_port_4, BBL_port_5, BBL_v;
  wire signed [`W-1:0] N0906_port_0, N0906_port_1, N0906_v;
  wire signed [`W-1:0] _OPR_1_port_15, _OPR_1_port_16, _OPR_1_v;
  wire signed [`W-1:0] N0964_port_2, N0964_port_1, N0964_v;
  wire signed [`W-1:0] _OPR_0_port_10, _OPR_0_port_11, _OPR_0_v;
  wire signed [`W-1:0] POC_port_3, POC_port_4, POC_v;
  wire signed [`W-1:0] N0650_port_0, N0650_port_1, N0650_v;
  wire signed [`W-1:0] N0357_port_2, N0357_port_3, N0357_port_0, N0357_port_1, N0357_port_4, N0357_port_5, N0357_v;
  wire signed [`W-1:0] N0996_port_2, N0996_port_0, N0996_v;
  wire signed [`W-1:0] cm_rom_port_0, cm_rom_port_1, cm_rom_v;
  wire signed [`W-1:0] N0585_port_0, N0585_port_1, N0585_v;
  wire signed [`W-1:0] cm_ram0_port_0, cm_ram0_port_1, cm_ram0_v;
  wire signed [`W-1:0] N0344_port_2, N0344_port_0, N0344_v;
  wire signed [`W-1:0] d2_port_2, d2_port_0, d2_port_1, d2_port_4, d2_port_5, d2_v;
  wire signed [`W-1:0] d3_port_2, d3_port_0, d3_port_1, d3_port_4, d3_port_5, d3_v;
  wire signed [`W-1:0] WRAB1_port_4, WRAB1_port_5, WRAB1_v;
  wire signed [`W-1:0] WRAB0_port_4, WRAB0_port_5, WRAB0_v;
  wire signed [`W-1:0] DCL_port_2, DCL_port_3, DCL_port_0, DCL_port_1, DCL_port_4, DCL_port_5, DCL_v;
  wire signed [`W-1:0] N0348_port_2, N0348_port_1, N0348_port_5, N0348_v;
  wire signed [`W-1:0] N0349_port_2, N0349_port_0, N0349_v;
  wire signed [`W-1:0] N0617_port_2, N0617_port_1, N0617_v;
  wire signed [`W-1:0] KBP_port_2, KBP_port_3, KBP_port_0, KBP_port_1, KBP_port_4, KBP_port_5, KBP_v;
  wire signed [`W-1:0] N0615_port_1, N0615_v;
  wire signed [`W-1:0] N0612_port_0, N0612_port_1, N0612_v;
  wire signed [`W-1:0] N0610_port_3, N0610_port_0, N0610_port_4, N0610_v;
  wire signed [`W-1:0] N0611_port_0, N0611_port_1, N0611_v;
  wire signed [`W-1:0] N0834_port_0, N0834_port_1, N0834_v;
  wire signed [`W-1:0] ACC_ADA_port_0, ACC_ADA_port_1, ACC_ADA_port_5, ACC_ADA_v;
  wire signed [`W-1:0] __POC__CLK2_SC_A32_X12__port_8, __POC__CLK2_SC_A32_X12__port_9, __POC__CLK2_SC_A32_X12__port_2, __POC__CLK2_SC_A32_X12__port_3, __POC__CLK2_SC_A32_X12__port_0, __POC__CLK2_SC_A32_X12__port_1, __POC__CLK2_SC_A32_X12__port_6, __POC__CLK2_SC_A32_X12__port_7, __POC__CLK2_SC_A32_X12__port_4, __POC__CLK2_SC_A32_X12__port_5, __POC__CLK2_SC_A32_X12__v;
  wire signed [`W-1:0] N0341_port_0, N0341_port_1, N0341_v;
  wire signed [`W-1:0] N0342_port_0, N0342_port_1, N0342_v;
  wire signed [`W-1:0] PC0_9_port_1, PC0_9_v;
  wire signed [`W-1:0] PC0_8_port_0, PC0_8_v;
  wire signed [`W-1:0] RADB2_port_6, RADB2_port_4, RADB2_port_5, RADB2_v;
  wire signed [`W-1:0] RADB0_port_6, RADB0_port_4, RADB0_port_5, RADB0_v;
  wire signed [`W-1:0] RADB1_port_6, RADB1_port_4, RADB1_port_5, RADB1_v;
  wire signed [`W-1:0] PC0_1_port_1, PC0_1_v;
  wire signed [`W-1:0] PC0_0_port_0, PC0_0_v;
  wire signed [`W-1:0] PC0_3_port_1, PC0_3_v;
  wire signed [`W-1:0] PC0_2_port_0, PC0_2_v;
  wire signed [`W-1:0] PC0_5_port_0, PC0_5_v;
  wire signed [`W-1:0] PC0_4_port_1, PC0_4_v;
  wire signed [`W-1:0] PC0_7_port_0, PC0_7_v;
  wire signed [`W-1:0] PC0_6_port_1, PC0_6_v;
  wire signed [`W-1:0] N0421_port_2, N0421_port_0, N0421_port_1, N0421_v;
  wire signed [`W-1:0] N0420_port_3, N0420_port_4, N0420_v;
  wire signed [`W-1:0] N0423_port_0, N0423_port_1, N0423_v;
  wire signed [`W-1:0] N0422_port_0, N0422_v;
  wire signed [`W-1:0] N0425_port_0, N0425_v;
  wire signed [`W-1:0] N0424_port_12, N0424_port_13, N0424_v;
  wire signed [`W-1:0] N0427_port_3, N0427_port_4, N0427_port_5, N0427_v;
  wire signed [`W-1:0] N0426_port_12, N0426_port_13, N0426_v;
  wire signed [`W-1:0] N0429_port_0, N0429_port_1, N0429_v;
  wire signed [`W-1:0] N0428_port_2, N0428_port_3, N0428_port_0, N0428_port_1, N0428_v;
  wire signed [`W-1:0] N0343_port_2, N0343_v;
  wire signed [`W-1:0] S00582_port_1, S00582_v;
  wire signed [`W-1:0] S00583_port_1, S00583_v;
  wire signed [`W-1:0] O_IB_port_2, O_IB_port_0, O_IB_port_1, O_IB_v;
  wire signed [`W-1:0] WRITE_CARRY_2__port_8, WRITE_CARRY_2__port_9, WRITE_CARRY_2__port_2, WRITE_CARRY_2__port_3, WRITE_CARRY_2__port_0, WRITE_CARRY_2__port_1, WRITE_CARRY_2__port_6, WRITE_CARRY_2__port_7, WRITE_CARRY_2__port_4, WRITE_CARRY_2__port_5, WRITE_CARRY_2__port_10, WRITE_CARRY_2__port_11, WRITE_CARRY_2__port_12, WRITE_CARRY_2__port_13, WRITE_CARRY_2__v;
  wire signed [`W-1:0] N0739_port_0, N0739_v;
  wire signed [`W-1:0] N0738_port_3, N0738_port_0, N0738_v;
  wire signed [`W-1:0] N0735_port_0, N0735_port_1, N0735_v;
  wire signed [`W-1:0] N0734_port_0, N0734_port_1, N0734_v;
  wire signed [`W-1:0] N0737_port_2, N0737_port_1, N0737_v;
  wire signed [`W-1:0] N0736_port_0, N0736_port_1, N0736_v;
  wire signed [`W-1:0] N0731_port_2, N0731_v;
  wire signed [`W-1:0] N0730_port_2, N0730_port_0, N0730_port_1, N0730_v;
  wire signed [`W-1:0] N0733_port_0, N0733_port_1, N0733_v;
  wire signed [`W-1:0] N0732_port_2, N0732_port_1, N0732_v;
  wire signed [`W-1:0] N0956_port_0, N0956_port_1, N0956_v;
  wire signed [`W-1:0] N0951_port_0, N0951_port_1, N0951_v;
  wire signed [`W-1:0] N0950_port_0, N0950_port_1, N0950_v;
  wire signed [`W-1:0] N0953_port_0, N0953_port_1, N0953_v;
  wire signed [`W-1:0] N0952_port_0, N0952_port_1, N0952_v;
  wire signed [`W-1:0] N0959_port_0, N0959_port_1, N0959_v;
  wire signed [`W-1:0] N0958_port_0, N0958_port_1, N0958_v;
  wire signed [`W-1:0] CY_port_2, CY_port_3, CY_port_0, CY_port_1, CY_port_5, CY_v;
  wire signed [`W-1:0] S00685_port_0, S00685_v;
  wire signed [`W-1:0] S00687_port_0, S00687_v;
  wire signed [`W-1:0] S00689_port_0, S00689_v;
  wire signed [`W-1:0] N0559_port_2, N0559_port_1, N0559_v;
  wire signed [`W-1:0] N0558_port_2, N0558_port_0, N0558_port_1, N0558_v;
  wire signed [`W-1:0] N0882_port_8, N0882_port_9, N0882_port_2, N0882_port_3, N0882_port_1, N0882_port_6, N0882_port_7, N0882_port_4, N0882_port_5, N0882_port_10, N0882_v;
  wire signed [`W-1:0] N0881_port_8, N0881_port_9, N0881_port_2, N0881_port_3, N0881_port_0, N0881_port_6, N0881_port_7, N0881_port_4, N0881_port_5, N0881_port_10, N0881_v;
  wire signed [`W-1:0] S00731_port_1, S00731_v;
  wire signed [`W-1:0] N0397_port_2, N0397_v;
  wire signed [`W-1:0] N0533_port_8, N0533_port_9, N0533_port_2, N0533_port_3, N0533_port_0, N0533_port_1, N0533_port_6, N0533_port_7, N0533_port_4, N0533_port_5, N0533_port_10, N0533_v;
  wire signed [`W-1:0] N0383_port_2, N0383_port_0, N0383_port_1, N0383_v;
  wire signed [`W-1:0] N0532_port_8, N0532_port_9, N0532_port_2, N0532_port_3, N0532_port_0, N0532_port_1, N0532_port_6, N0532_port_7, N0532_port_4, N0532_port_5, N0532_port_10, N0532_v;
  wire signed [`W-1:0] N0531_port_8, N0531_port_9, N0531_port_2, N0531_port_3, N0531_port_0, N0531_port_1, N0531_port_6, N0531_port_7, N0531_port_4, N0531_port_5, N0531_port_10, N0531_v;
  wire signed [`W-1:0] N0537_port_8, N0537_port_9, N0537_port_2, N0537_port_3, N0537_port_0, N0537_port_1, N0537_port_6, N0537_port_7, N0537_port_4, N0537_port_5, N0537_port_10, N0537_v;
  wire signed [`W-1:0] S00836_port_0, S00836_v;
  wire signed [`W-1:0] N0641_port_2, N0641_port_0, N0641_port_1, N0641_v;
  wire signed [`W-1:0] S00724_port_1, S00724_v;
  wire signed [`W-1:0] IOW_port_2, IOW_port_0, IOW_port_1, IOW_v;
  wire signed [`W-1:0] IOR_port_3, IOR_port_1, IOR_port_5, IOR_v;
  wire signed [`W-1:0] N0356_port_8, N0356_port_9, N0356_port_6, N0356_v;
  wire signed [`W-1:0] N0643_port_2, N0643_port_1, N0643_v;
  wire signed [`W-1:0] N0642_port_3, N0642_port_0, N0642_port_4, N0642_v;
  wire signed [`W-1:0] S00833_port_0, S00833_v;
  wire signed [`W-1:0] PC2_11_port_1, PC2_11_v;
  wire signed [`W-1:0] PC2_10_port_0, PC2_10_v;
  wire signed [`W-1:0] N0890_port_0, N0890_port_1, N0890_v;
  wire signed [`W-1:0] N0644_port_0, N0644_port_1, N0644_v;
  wire signed [`W-1:0] N0891_port_4, N0891_port_5, N0891_v;
  wire signed [`W-1:0] JMS_port_2, JMS_port_3, JMS_port_1, JMS_port_4, JMS_port_5, JMS_v;
  wire signed [`W-1:0] N0892_port_0, N0892_port_1, N0892_v;
  wire signed [`W-1:0] CY_IB_port_2, CY_IB_port_0, CY_IB_port_1, CY_IB_v;
  wire signed [`W-1:0] N0358_port_2, N0358_port_3, N0358_port_0, N0358_port_1, N0358_port_6, N0358_port_7, N0358_port_4, N0358_port_5, N0358_v;
  wire signed [`W-1:0] SUB_port_2, SUB_port_3, SUB_port_0, SUB_port_1, SUB_port_4, SUB_v;
  wire signed [`W-1:0] N0432_port_0, N0432_port_1, N0432_v;
  wire signed [`W-1:0] N0433_port_0, N0433_v;
  wire signed [`W-1:0] N0430_port_2, N0430_port_0, N0430_port_1, N0430_v;
  wire signed [`W-1:0] N0431_port_0, N0431_v;
  wire signed [`W-1:0] N0436_port_3, N0436_port_0, N0436_port_4, N0436_port_5, N0436_v;
  wire signed [`W-1:0] N0437_port_2, N0437_port_0, N0437_v;
  wire signed [`W-1:0] N0434_port_12, N0434_port_13, N0434_v;
  wire signed [`W-1:0] N0435_port_2, N0435_port_1, N0435_v;
  wire signed [`W-1:0] N0438_port_1, N0438_v;
  wire signed [`W-1:0] N0439_port_12, N0439_port_13, N0439_v;
  wire signed [`W-1:0] ADD_port_2, ADD_port_3, ADD_port_0, ADD_port_1, ADD_port_4, ADD_v;
  wire signed [`W-1:0] ADM_port_2, ADM_port_3, ADM_port_0, ADM_port_1, ADM_port_4, ADM_port_5, ADM_v;
  wire signed [`W-1:0] reset_port_2, reset_port_0, reset_v;
  wire signed [`W-1:0] N0728_port_2, N0728_port_0, N0728_port_1, N0728_v;
  wire signed [`W-1:0] N0729_port_2, N0729_v;
  wire signed [`W-1:0] N0726_port_2, N0726_port_0, N0726_port_1, N0726_v;
  wire signed [`W-1:0] N0727_port_2, N0727_v;
  wire signed [`W-1:0] N0724_port_2, N0724_port_0, N0724_port_1, N0724_v;
  wire signed [`W-1:0] N0725_port_2, N0725_v;
  wire signed [`W-1:0] N0722_port_2, N0722_port_0, N0722_port_1, N0722_v;
  wire signed [`W-1:0] N0723_port_2, N0723_v;
  wire signed [`W-1:0] N0720_port_2, N0720_port_0, N0720_port_1, N0720_v;
  wire signed [`W-1:0] N0721_port_2, N0721_v;
  wire signed [`W-1:0] N0946_port_2, N0946_port_1, N0946_v;
  wire signed [`W-1:0] N0944_port_2, N0944_port_1, N0944_v;
  wire signed [`W-1:0] N0942_port_2, N0942_port_1, N0942_v;
  wire signed [`W-1:0] N0943_port_3, N0943_port_4, N0943_v;
  wire signed [`W-1:0] N0940_port_2, N0940_port_1, N0940_v;
  wire signed [`W-1:0] N0948_port_0, N0948_port_1, N0948_v;
  wire signed [`W-1:0] N0949_port_0, N0949_port_1, N0949_v;
  wire signed [`W-1:0] N0894_port_0, N0894_port_1, N0894_v;
  wire signed [`W-1:0] N0895_port_0, N0895_port_1, N0895_v;
  wire signed [`W-1:0] N0897_port_0, N0897_port_1, N0897_v;
  wire signed [`W-1:0] N0893_port_4, N0893_port_5, N0893_v;
  wire signed [`W-1:0] N0898_port_2, N0898_port_3, N0898_port_0, N0898_port_1, N0898_v;
  wire signed [`W-1:0] N0899_port_2, N0899_port_3, N0899_port_0, N0899_port_1, N0899_v;
  wire signed [`W-1:0] N0548_port_2, N0548_port_0, N0548_port_1, N0548_v;
  wire signed [`W-1:0] N0549_port_2, N0549_port_0, N0549_port_1, N0549_v;
  wire signed [`W-1:0] S00839_port_1, S00839_v;
  wire signed [`W-1:0] N0542_port_4, N0542_port_5, N0542_v;
  wire signed [`W-1:0] N0543_port_8, N0543_port_9, N0543_v;
  wire signed [`W-1:0] N0540_port_1, N0540_port_5, N0540_v;
  wire signed [`W-1:0] N0541_port_4, N0541_port_5, N0541_v;
  wire signed [`W-1:0] N0546_port_2, N0546_port_0, N0546_port_1, N0546_v;
  wire signed [`W-1:0] N0547_port_2, N0547_port_0, N0547_v;
  wire signed [`W-1:0] N0544_port_8, N0544_port_9, N0544_v;
  wire signed [`W-1:0] N0545_port_3, N0545_port_6, N0545_port_7, N0545_port_4, N0545_port_5, N0545_v;
  wire signed [`W-1:0] N0467_port_2, N0467_port_3, N0467_port_1, N0467_port_4, N0467_port_5, N0467_v;
  wire signed [`W-1:0] N0466_port_2, N0466_port_3, N0466_port_6, N0466_v;
  wire signed [`W-1:0] INC_GROUP_5__port_2, INC_GROUP_5__port_3, INC_GROUP_5__port_0, INC_GROUP_5__port_1, INC_GROUP_5__v;
  wire signed [`W-1:0] N0502_port_2, N0502_port_0, N0502_v;
  wire signed [`W-1:0] N0682_port_2, N0682_port_3, N0682_port_0, N0682_port_1, N0682_port_4, N0682_v;
  wire signed [`W-1:0] _OPR_3_port_10, _OPR_3_port_11, _OPR_3_v;
  wire signed [`W-1:0] _OPR_2_port_12, _OPR_2_port_13, _OPR_2_v;
  wire signed [`W-1:0] N0966_port_0, N0966_port_1, N0966_v;
  wire signed [`W-1:0] N0517_port_1, N0517_v;
  wire signed [`W-1:0] N0516_port_0, N0516_port_1, N0516_v;
  wire signed [`W-1:0] XCH_port_2, XCH_port_3, XCH_port_0, XCH_port_1, XCH_port_4, XCH_v;
  wire signed [`W-1:0] CMC_port_2, CMC_port_3, CMC_port_0, CMC_port_1, CMC_port_4, CMC_port_5, CMC_v;
  wire signed [`W-1:0] CMA_port_2, CMA_port_3, CMA_port_0, CMA_port_1, CMA_port_4, CMA_port_5, CMA_v;
  wire signed [`W-1:0] N0510_port_0, N0510_port_1, N0510_v;
  wire signed [`W-1:0] N0513_port_2, N0513_port_3, N0513_port_0, N0513_port_1, N0513_v;
  wire signed [`W-1:0] M22_port_8, M22_port_10, M22_port_11, M22_v;
  wire signed [`W-1:0] JUN2_JMS2_port_2, JUN2_JMS2_port_3, JUN2_JMS2_port_0, JUN2_JMS2_port_1, JUN2_JMS2_v;
  wire signed [`W-1:0] N0361_port_2, N0361_port_0, N0361_port_1, N0361_v;
  wire signed [`W-1:0] N0512_port_0, N0512_port_1, N0512_v;
  wire signed [`W-1:0] N0345_port_2, N0345_port_3, N0345_port_0, N0345_port_1, N0345_port_4, N0345_port_5, N0345_v;
  wire signed [`W-1:0] SC_A22_M22_CLK2_port_8, SC_A22_M22_CLK2_port_9, SC_A22_M22_CLK2_v;
  wire signed [`W-1:0] OPA_IB_port_6, OPA_IB_port_4, OPA_IB_port_5, OPA_IB_v;
  wire signed [`W-1:0] S00654_port_1, S00654_v;
  wire signed [`W-1:0] S00818_port_0, S00818_v;
  wire signed [`W-1:0] N0367_port_0, N0367_port_1, N0367_v;
  wire signed [`W-1:0] N0364_port_3, N0364_port_0, N0364_port_1, N0364_v;
  wire signed [`W-1:0] N0362_port_1, N0362_v;
  wire signed [`W-1:0] N0363_port_2, N0363_port_3, N0363_port_0, N0363_port_1, N0363_port_4, N0363_port_5, N0363_v;
  wire signed [`W-1:0] N0360_port_1, N0360_v;
  wire signed [`W-1:0] S00729_port_1, S00729_v;
  wire signed [`W-1:0] N0399_port_2, N0399_port_0, N0399_v;
  wire signed [`W-1:0] N0396_port_2, N0396_port_3, N0396_port_0, N0396_port_1, N0396_port_6, N0396_port_4, N0396_port_5, N0396_v;
  wire signed [`W-1:0] N0395_port_2, N0395_port_3, N0395_port_0, N0395_port_1, N0395_port_6, N0395_port_4, N0395_port_5, N0395_v;
  wire signed [`W-1:0] N0394_port_2, N0394_port_3, N0394_port_0, N0394_port_1, N0394_port_6, N0394_port_4, N0394_port_5, N0394_v;
  wire signed [`W-1:0] N0393_port_2, N0393_port_3, N0393_port_0, N0393_port_1, N0393_port_6, N0393_port_4, N0393_port_5, N0393_v;
  wire signed [`W-1:0] N0392_port_2, N0392_port_3, N0392_port_0, N0392_port_1, N0392_port_6, N0392_port_4, N0392_port_5, N0392_v;
  wire signed [`W-1:0] N0391_port_2, N0391_port_3, N0391_port_0, N0391_port_1, N0391_port_6, N0391_port_4, N0391_port_5, N0391_v;
  wire signed [`W-1:0] N0390_port_2, N0390_port_3, N0390_port_0, N0390_port_1, N0390_port_6, N0390_port_4, N0390_port_5, N0390_v;
  wire signed [`W-1:0] N0409_port_3, N0409_port_4, N0409_v;
  wire signed [`W-1:0] N0408_port_0, N0408_v;
  wire signed [`W-1:0] N0407_port_2, N0407_port_0, N0407_port_1, N0407_v;
  wire signed [`W-1:0] N0406_port_12, N0406_port_13, N0406_v;
  wire signed [`W-1:0] N0405_port_1, N0405_v;
  wire signed [`W-1:0] N0404_port_2, N0404_port_0, N0404_port_1, N0404_v;
  wire signed [`W-1:0] N0403_port_3, N0403_port_0, N0403_port_1, N0403_v;
  wire signed [`W-1:0] N0402_port_2, N0402_port_0, N0402_port_1, N0402_v;
  wire signed [`W-1:0] N0401_port_2, N0401_port_3, N0401_v;
  wire signed [`W-1:0] N0400_port_0, N0400_port_1, N0400_v;
  wire signed [`W-1:0] SBM_port_2, SBM_port_3, SBM_port_0, SBM_port_1, SBM_port_4, SBM_port_5, SBM_v;
  wire signed [`W-1:0] _CN_port_2, _CN_port_3, _CN_v;
  wire signed [`W-1:0] S00678_port_1, S00678_v;
  wire signed [`W-1:0] N0719_port_2, N0719_v;
  wire signed [`W-1:0] N0718_port_2, N0718_port_0, N0718_port_1, N0718_v;
  wire signed [`W-1:0] N0713_port_2, N0713_port_0, N0713_port_1, N0713_v;
  wire signed [`W-1:0] N0712_port_2, N0712_port_0, N0712_port_1, N0712_v;
  wire signed [`W-1:0] N0711_port_2, N0711_port_0, N0711_port_1, N0711_v;
  wire signed [`W-1:0] N0710_port_2, N0710_port_1, N0710_v;
  wire signed [`W-1:0] N0717_port_2, N0717_port_3, N0717_port_4, N0717_v;
  wire signed [`W-1:0] N0715_port_0, N0715_port_1, N0715_port_4, N0715_v;
  wire signed [`W-1:0] N0714_port_2, N0714_port_0, N0714_port_1, N0714_v;
  wire signed [`W-1:0] N0973_port_0, N0973_port_1, N0973_v;
  wire signed [`W-1:0] N0972_port_0, N0972_port_1, N0972_v;
  wire signed [`W-1:0] N0971_port_0, N0971_port_1, N0971_v;
  wire signed [`W-1:0] N0970_port_0, N0970_port_1, N0970_v;
  wire signed [`W-1:0] N0977_port_0, N0977_port_1, N0977_v;
  wire signed [`W-1:0] N0976_port_0, N0976_port_1, N0976_v;
  wire signed [`W-1:0] N0975_port_0, N0975_port_1, N0975_v;
  wire signed [`W-1:0] N0974_port_2, N0974_port_3, N0974_v;
  wire signed [`W-1:0] N0979_port_0, N0979_port_1, N0979_v;
  wire signed [`W-1:0] N0978_port_0, N0978_port_1, N0978_v;
  wire signed [`W-1:0] SC_M12_CLK2_port_0, SC_M12_CLK2_port_1, SC_M12_CLK2_v;
  wire signed [`W-1:0] N0577_port_6, N0577_port_5, N0577_v;
  wire signed [`W-1:0] N0576_port_0, N0576_port_1, N0576_v;
  wire signed [`W-1:0] N0575_port_2, N0575_port_0, N0575_port_1, N0575_v;
  wire signed [`W-1:0] N0574_port_3, N0574_port_0, N0574_port_4, N0574_v;
  wire signed [`W-1:0] N0573_port_2, N0573_port_0, N0573_port_1, N0573_v;
  wire signed [`W-1:0] N0572_port_0, N0572_port_1, N0572_v;
  wire signed [`W-1:0] N0571_port_2, N0571_port_0, N0571_port_1, N0571_v;
  wire signed [`W-1:0] N0570_port_3, N0570_port_6, N0570_port_7, N0570_port_4, N0570_port_5, N0570_v;
  wire signed [`W-1:0] N0579_port_0, N0579_port_1, N0579_v;
  wire signed [`W-1:0] N0578_port_2, N0578_port_1, N0578_v;
  wire signed [`W-1:0] S00825_port_0, S00825_v;
  wire signed [`W-1:0] S00531_port_0, S00531_v;
  wire signed [`W-1:0] N0379_port_2, N0379_port_0, N0379_port_1, N0379_v;
  wire signed [`W-1:0] S00536_port_1, S00536_v;
  wire signed [`W-1:0] PC1_0_port_0, PC1_0_v;
  wire signed [`W-1:0] R14_1_port_1, R14_1_v;
  wire signed [`W-1:0] R14_0_port_0, R14_0_v;
  wire signed [`W-1:0] R14_3_port_1, R14_3_v;
  wire signed [`W-1:0] R14_2_port_0, R14_2_v;
  wire signed [`W-1:0] R10_1_port_1, R10_1_v;
  wire signed [`W-1:0] R10_0_port_0, R10_0_v;
  wire signed [`W-1:0] R10_3_port_1, R10_3_v;
  wire signed [`W-1:0] R10_2_port_0, R10_2_v;
  wire signed [`W-1:0] N0889_port_4, N0889_port_5, N0889_v;
  wire signed [`W-1:0] N0515_port_2, N0515_port_0, N0515_v;
  wire signed [`W-1:0] N0514_port_2, N0514_port_3, N0514_port_0, N0514_port_6, N0514_port_4, N0514_port_5, N0514_v;
  wire signed [`W-1:0] N0888_port_0, N0888_port_1, N0888_v;
  wire signed [`W-1:0] N0845_port_0, N0845_port_1, N0845_v;
  wire signed [`W-1:0] N0844_port_0, N0844_port_1, N0844_v;
  wire signed [`W-1:0] N0511_port_2, N0511_port_3, N0511_port_0, N0511_port_1, N0511_v;
  wire signed [`W-1:0] N0842_port_0, N0842_port_1, N0842_v;
  wire signed [`W-1:0] N0371_port_2, N0371_port_3, N0371_port_0, N0371_v;
  wire signed [`W-1:0] N0849_port_1, N0849_v;
  wire signed [`W-1:0] N0848_port_2, N0848_port_0, N0848_port_1, N0848_port_6, N0848_port_4, N0848_port_5, N0848_v;
  wire signed [`W-1:0] ISZ_port_2, ISZ_port_3, ISZ_port_0, ISZ_port_1, ISZ_port_4, ISZ_v;
  wire signed [`W-1:0] N0370_port_2, N0370_port_3, N0370_port_0, N0370_port_1, N0370_port_4, N0370_port_5, N0370_v;
  wire signed [`W-1:0] N0875_port_3, N0875_port_1, N0875_port_4, N0875_v;
  wire signed [`W-1:0] R12_3_port_1, R12_3_v;
  wire signed [`W-1:0] CLB_port_2, CLB_port_3, CLB_port_0, CLB_port_1, CLB_port_4, CLB_port_5, CLB_v;
  wire signed [`W-1:0] CLC_port_2, CLC_port_3, CLC_port_0, CLC_port_1, CLC_port_4, CLC_port_5, CLC_v;
  wire signed [`W-1:0] M12_port_10, M12_port_11, M12_port_8, M12_port_7, M12_v;
  wire signed [`W-1:0] __X21__CLK2__port_2, __X21__CLK2__port_3, __X21__CLK2__v;
  wire signed [`W-1:0] DC_port_4, DC_port_5, DC_v;
  wire signed [`W-1:0] N0388_port_2, N0388_port_3, N0388_port_0, N0388_port_1, N0388_port_6, N0388_port_4, N0388_port_5, N0388_v;
  wire signed [`W-1:0] N0389_port_2, N0389_port_3, N0389_port_0, N0389_port_1, N0389_port_6, N0389_port_4, N0389_port_5, N0389_v;
  wire signed [`W-1:0] N0380_port_0, N0380_v;
  wire signed [`W-1:0] N0381_port_12, N0381_port_13, N0381_v;
  wire signed [`W-1:0] N0382_port_3, N0382_port_4, N0382_port_5, N0382_v;
  wire signed [`W-1:0] N0384_port_1, N0384_v;
  wire signed [`W-1:0] N0385_port_2, N0385_port_3, N0385_port_0, N0385_port_1, N0385_port_6, N0385_port_4, N0385_port_5, N0385_v;
  wire signed [`W-1:0] N0386_port_2, N0386_port_3, N0386_port_0, N0386_port_1, N0386_port_6, N0386_port_4, N0386_port_5, N0386_v;
  wire signed [`W-1:0] N0387_port_2, N0387_port_3, N0387_port_0, N0387_port_1, N0387_port_6, N0387_port_4, N0387_port_5, N0387_v;
  wire signed [`W-1:0] R12_0_port_0, R12_0_v;
  wire signed [`W-1:0] N0419_port_2, N0419_port_3, N0419_port_1, N0419_v;
  wire signed [`W-1:0] N0410_port_12, N0410_port_13, N0410_v;
  wire signed [`W-1:0] N0411_port_3, N0411_port_4, N0411_port_5, N0411_v;
  wire signed [`W-1:0] N0412_port_0, N0412_port_1, N0412_v;
  wire signed [`W-1:0] N0413_port_2, N0413_port_3, N0413_port_0, N0413_port_1, N0413_v;
  wire signed [`W-1:0] N0414_port_0, N0414_v;
  wire signed [`W-1:0] N0415_port_2, N0415_port_0, N0415_port_1, N0415_v;
  wire signed [`W-1:0] N0416_port_1, N0416_v;
  wire signed [`W-1:0] N0417_port_0, N0417_port_1, N0417_v;
  wire signed [`W-1:0] _COM_port_0, _COM_port_1, _COM_v;
  wire signed [`W-1:0] N0901_port_2, N0901_port_3, N0901_port_0, N0901_port_1, N0901_v;
  wire signed [`W-1:0] N0704_port_0, N0704_port_1, N0704_v;
  wire signed [`W-1:0] N0705_port_2, N0705_port_3, N0705_port_0, N0705_port_1, N0705_v;
  wire signed [`W-1:0] N0706_port_0, N0706_port_1, N0706_v;
  wire signed [`W-1:0] N0707_port_0, N0707_v;
  wire signed [`W-1:0] N0700_port_2, N0700_port_3, N0700_v;
  wire signed [`W-1:0] N0701_port_2, N0701_port_3, N0701_port_0, N0701_port_1, N0701_v;
  wire signed [`W-1:0] N0702_port_0, N0702_port_1, N0702_v;
  wire signed [`W-1:0] N0703_port_0, N0703_v;
  wire signed [`W-1:0] N0708_port_2, N0708_port_3, N0708_port_4, N0708_port_5, N0708_v;
  wire signed [`W-1:0] N0709_port_0, N0709_port_1, N0709_v;
  wire signed [`W-1:0] N0885_port_2, N0885_port_1, N0885_v;
  wire signed [`W-1:0] N0378_port_2, N0378_port_0, N0378_port_1, N0378_v;
  wire signed [`W-1:0] D2_port_8, D2_port_9, D2_port_2, D2_port_3, D2_port_0, D2_port_1, D2_port_6, D2_port_7, D2_port_4, D2_port_5, D2_port_10, D2_port_11, D2_port_13, D2_port_14, D2_port_15, D2_port_16, D2_port_17, D2_port_18, D2_v;
  wire signed [`W-1:0] D3_port_8, D3_port_9, D3_port_2, D3_port_3, D3_port_0, D3_port_1, D3_port_6, D3_port_7, D3_port_4, D3_port_5, D3_port_11, D3_port_12, D3_port_13, D3_port_14, D3_port_15, D3_port_16, D3_port_17, D3_port_18, D3_v;
  wire signed [`W-1:0] D0_port_8, D0_port_9, D0_port_2, D0_port_3, D0_port_0, D0_port_1, D0_port_6, D0_port_7, D0_port_4, D0_port_5, D0_port_10, D0_port_11, D0_port_12, D0_port_13, D0_port_14, D0_port_15, D0_port_16, D0_port_17, D0_v;
  wire signed [`W-1:0] D1_port_8, D1_port_9, D1_port_2, D1_port_3, D1_port_0, D1_port_1, D1_port_6, D1_port_7, D1_port_4, D1_port_5, D1_port_10, D1_port_11, D1_port_12, D1_port_13, D1_port_14, D1_port_15, D1_port_16, D1_port_17, D1_v;
  wire signed [`W-1:0] N0968_port_0, N0968_port_1, N0968_v;
  wire signed [`W-1:0] N0969_port_0, N0969_port_1, N0969_v;
  wire signed [`W-1:0] N0965_port_2, N0965_port_3, N0965_v;
  wire signed [`W-1:0] N0967_port_0, N0967_port_1, N0967_v;
  wire signed [`W-1:0] N0960_port_0, N0960_port_1, N0960_v;
  wire signed [`W-1:0] N0961_port_0, N0961_port_1, N0961_v;
  wire signed [`W-1:0] N0962_port_0, N0962_port_1, N0962_v;
  wire signed [`W-1:0] N0963_port_0, N0963_port_1, N0963_v;
  wire signed [`W-1:0] N0907_port_0, N0907_port_1, N0907_v;
  wire signed [`W-1:0] N0884_port_2, N0884_port_1, N0884_v;
  wire signed [`W-1:0] N0560_port_6, N0560_port_5, N0560_v;
  wire signed [`W-1:0] N0561_port_0, N0561_port_1, N0561_v;
  wire signed [`W-1:0] N0562_port_2, N0562_port_0, N0562_port_1, N0562_v;
  wire signed [`W-1:0] N0563_port_0, N0563_port_1, N0563_v;
  wire signed [`W-1:0] N0564_port_3, N0564_port_0, N0564_v;
  wire signed [`W-1:0] N0565_port_8, N0565_port_9, N0565_v;
  wire signed [`W-1:0] N0566_port_0, N0566_v;
  wire signed [`W-1:0] N0567_port_0, N0567_port_1, N0567_v;
  wire signed [`W-1:0] N0568_port_0, N0568_port_1, N0568_v;
  wire signed [`W-1:0] N0569_port_8, N0569_port_9, N0569_v;
  wire signed [`W-1:0] N0365_port_2, N0365_port_0, N0365_port_1, N0365_v;
  wire signed [`W-1:0] S00814_port_0, S00814_v;
  wire signed [`W-1:0] N0368_port_2, N0368_port_3, N0368_port_0, N0368_port_1, N0368_v;
  wire signed [`W-1:0] N0369_port_2, N0369_port_0, N0369_port_1, N0369_v;
  wire signed [`W-1:0] S00676_port_0, S00676_v;
  wire signed [`W-1:0] N0640_port_0, N0640_port_1, N0640_v;
  wire signed [`W-1:0] N0314_port_2, N0314_port_0, N0314_port_1, N0314_v;
  wire signed [`W-1:0] _OPA_0_port_13, _OPA_0_port_14, _OPA_0_v;
  wire signed [`W-1:0] N0311_port_0, N0311_port_1, N0311_v;
  wire signed [`W-1:0] _OPA_2_port_6, _OPA_2_port_7, _OPA_2_v;
  wire signed [`W-1:0] _OPA_3_port_10, _OPA_3_port_11, _OPA_3_v;
  wire signed [`W-1:0] N0646_port_2, N0646_port_1, N0646_v;
  wire signed [`W-1:0] ADD_GROUP_4__port_2, ADD_GROUP_4__port_3, ADD_GROUP_4__port_0, ADD_GROUP_4__port_1, ADD_GROUP_4__port_4, ADD_GROUP_4__v;
  wire signed [`W-1:0] ___SC__JIN_FIN__CLK1_M11_X21_INH__port_2, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_3, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_0, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_1, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_4, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_5, ___SC__JIN_FIN__CLK1_M11_X21_INH__v;
  wire signed [`W-1:0] N0486_port_2, N0486_port_3, N0486_port_4, N0486_port_5, N0486_v;
  wire signed [`W-1:0] N0860_port_0, N0860_port_1, N0860_v;
  wire signed [`W-1:0] N0947_port_0, N0947_port_1, N0947_v;
  wire signed [`W-1:0] N0941_port_3, N0941_port_4, N0941_v;
  wire signed [`W-1:0] N0861_port_2, N0861_port_3, N0861_port_0, N0861_v;
  wire signed [`W-1:0] N0863_port_2, N0863_port_3, N0863_port_0, N0863_port_1, N0863_v;
  wire signed [`W-1:0] N0862_port_2, N0862_port_3, N0862_port_0, N0862_port_1, N0862_v;
  wire signed [`W-1:0] N0865_port_2, N0865_port_3, N0865_port_0, N0865_port_1, N0865_v;
  wire signed [`W-1:0] N0864_port_2, N0864_port_3, N0864_port_0, N0864_port_1, N0864_v;
  wire signed [`W-1:0] WRITE_ACC_1__port_8, WRITE_ACC_1__port_9, WRITE_ACC_1__port_2, WRITE_ACC_1__port_3, WRITE_ACC_1__port_0, WRITE_ACC_1__port_1, WRITE_ACC_1__port_6, WRITE_ACC_1__port_7, WRITE_ACC_1__port_4, WRITE_ACC_1__port_5, WRITE_ACC_1__port_10, WRITE_ACC_1__port_11, WRITE_ACC_1__port_12, WRITE_ACC_1__port_13, WRITE_ACC_1__port_14, WRITE_ACC_1__port_15, WRITE_ACC_1__v;
  wire signed [`W-1:0] N0866_port_8, N0866_port_9, N0866_port_2, N0866_port_3, N0866_port_0, N0866_port_6, N0866_port_7, N0866_port_4, N0866_port_5, N0866_port_10, N0866_v;
  wire signed [`W-1:0] N0855_port_2, N0855_port_3, N0855_port_1, N0855_port_4, N0855_v;
  wire signed [`W-1:0] N0896_port_0, N0896_port_1, N0896_v;
  wire signed [`W-1:0] IO_port_2, IO_port_3, IO_port_0, IO_port_1, IO_port_4, IO_v;
  wire signed [`W-1:0] N0911_port_2, N0911_port_0, N0911_port_1, N0911_v;
  wire signed [`W-1:0] N0621_port_0, N0621_port_1, N0621_v;
  wire signed [`W-1:0] N0910_port_0, N0910_port_1, N0910_v;
  wire signed [`W-1:0] N0280_port_0, N0280_v;
  wire signed [`W-1:0] N0284_port_1, N0284_v;
  wire signed [`W-1:0] N0286_port_1, N0286_v;
  wire signed [`W-1:0] N0289_port_3, N0289_v;
  wire signed [`W-1:0] N0288_port_8, N0288_port_2, N0288_port_3, N0288_port_0, N0288_port_1, N0288_port_6, N0288_port_7, N0288_port_4, N0288_port_5, N0288_v;
  wire signed [`W-1:0] N0771_port_2, N0771_port_3, N0771_port_1, N0771_port_6, N0771_port_4, N0771_port_5, N0771_v;
  wire signed [`W-1:0] N0770_port_2, N0770_port_3, N0770_port_1, N0770_port_6, N0770_port_4, N0770_port_5, N0770_v;
  wire signed [`W-1:0] N0773_port_2, N0773_port_3, N0773_port_1, N0773_port_6, N0773_port_4, N0773_port_5, N0773_v;
  wire signed [`W-1:0] N0772_port_2, N0772_port_3, N0772_port_1, N0772_port_6, N0772_port_4, N0772_port_5, N0772_v;
  wire signed [`W-1:0] N0775_port_2, N0775_port_3, N0775_port_0, N0775_port_6, N0775_port_4, N0775_port_5, N0775_v;
  wire signed [`W-1:0] N0774_port_2, N0774_port_3, N0774_port_0, N0774_port_6, N0774_port_4, N0774_port_5, N0774_v;
  wire signed [`W-1:0] N0777_port_2, N0777_port_3, N0777_port_1, N0777_port_6, N0777_port_4, N0777_port_5, N0777_v;
  wire signed [`W-1:0] N0776_port_2, N0776_port_3, N0776_port_0, N0776_port_6, N0776_port_4, N0776_port_5, N0776_v;
  wire signed [`W-1:0] N0779_port_2, N0779_port_3, N0779_port_0, N0779_port_6, N0779_port_4, N0779_port_5, N0779_v;
  wire signed [`W-1:0] N0778_port_2, N0778_port_3, N0778_port_0, N0778_port_6, N0778_port_4, N0778_port_5, N0778_v;
  wire signed [`W-1:0] N0919_port_2, N0919_port_3, N0919_v;
  wire signed [`W-1:0] N0918_port_0, N0918_port_1, N0918_v;
  wire signed [`W-1:0] N0626_port_3, N0626_port_1, N0626_port_4, N0626_v;
  wire signed [`W-1:0] N0914_port_2, N0914_port_0, N0914_port_1, N0914_v;
  wire signed [`W-1:0] test_port_2, test_port_0, test_v;
  wire signed [`W-1:0] S00834_port_0, S00834_v;
  wire signed [`W-1:0] N0915_port_0, N0915_port_1, N0915_v;
  wire signed [`W-1:0] S00804_port_0, S00804_v;
  wire signed [`W-1:0] N0599_port_3, N0599_port_6, N0599_port_7, N0599_port_4, N0599_port_5, N0599_v;
  wire signed [`W-1:0] N0598_port_8, N0598_port_9, N0598_v;
  wire signed [`W-1:0] S00801_port_1, S00801_v;
  wire signed [`W-1:0] S00800_port_0, S00800_v;
  wire signed [`W-1:0] N0595_port_0, N0595_port_1, N0595_v;
  wire signed [`W-1:0] N0594_port_0, N0594_port_1, N0594_v;
  wire signed [`W-1:0] N0597_port_0, N0597_port_1, N0597_v;
  wire signed [`W-1:0] N0596_port_0, N0596_port_1, N0596_v;
  wire signed [`W-1:0] N0591_port_8, N0591_port_9, N0591_v;
  wire signed [`W-1:0] N0590_port_2, N0590_port_1, N0590_v;
  wire signed [`W-1:0] N0593_port_0, N0593_v;
  wire signed [`W-1:0] N0592_port_1, N0592_v;
  wire signed [`W-1:0] N0609_port_2, N0609_port_0, N0609_port_1, N0609_v;
  wire signed [`W-1:0] N0359_port_2, N0359_port_3, N0359_port_0, N0359_port_1, N0359_port_4, N0359_port_5, N0359_v;
  wire signed [`W-1:0] N0606_port_0, N0606_port_1, N0606_v;
  wire signed [`W-1:0] N0601_port_0, N0601_port_1, N0601_v;
  wire signed [`W-1:0] N0600_port_2, N0600_port_3, N0600_port_0, N0600_v;
  wire signed [`W-1:0] N0603_port_2, N0603_port_1, N0603_v;
  wire signed [`W-1:0] N0602_port_2, N0602_port_0, N0602_port_1, N0602_v;
  wire signed [`W-1:0] N0825_port_0, N0825_port_1, N0825_v;
  wire signed [`W-1:0] N0827_port_0, N0827_port_1, N0827_v;
  wire signed [`W-1:0] N0826_port_0, N0826_port_1, N0826_v;
  wire signed [`W-1:0] N0821_port_0, N0821_port_1, N0821_v;
  wire signed [`W-1:0] N0917_port_0, N0917_port_1, N0917_v;
  wire signed [`W-1:0] __INH__X11_X31_CLK1_port_12, __INH__X11_X31_CLK1_port_13, __INH__X11_X31_CLK1_port_14, __INH__X11_X31_CLK1_port_15, __INH__X11_X31_CLK1_v;
  wire signed [`W-1:0] S00761_port_0, S00761_v;
  wire signed [`W-1:0] N0817_port_0, N0817_port_1, N0817_v;
  wire signed [`W-1:0] N0811_port_0, N0811_port_1, N0811_v;
  wire signed [`W-1:0] S00781_port_1, S00781_v;
  wire signed [`W-1:0] CY_ADAC_port_2, CY_ADAC_port_0, CY_ADAC_port_1, CY_ADAC_v;
  wire signed [`W-1:0] N0652_port_0, N0652_port_1, N0652_v;
  wire signed [`W-1:0] CLK2_SC_A12_M12__port_8, CLK2_SC_A12_M12__port_9, CLK2_SC_A12_M12__port_2, CLK2_SC_A12_M12__port_3, CLK2_SC_A12_M12__port_0, CLK2_SC_A12_M12__port_1, CLK2_SC_A12_M12__port_6, CLK2_SC_A12_M12__port_7, CLK2_SC_A12_M12__port_4, CLK2_SC_A12_M12__port_5, CLK2_SC_A12_M12__v;
  wire signed [`W-1:0] N0292_port_4, N0292_v;
  wire signed [`W-1:0] N0293_port_2, N0293_port_3, N0293_v;
  wire signed [`W-1:0] N0290_port_0, N0290_v;
  wire signed [`W-1:0] N0291_port_5, N0291_v;
  wire signed [`W-1:0] N0296_port_2, N0296_port_3, N0296_port_0, N0296_port_1, N0296_v;
  wire signed [`W-1:0] N0297_port_0, N0297_port_1, N0297_v;
  wire signed [`W-1:0] N0294_port_2, N0294_port_3, N0294_port_0, N0294_port_1, N0294_v;
  wire signed [`W-1:0] N0295_port_1, N0295_v;
  wire signed [`W-1:0] N0298_port_3, N0298_port_0, N0298_v;
  wire signed [`W-1:0] N0299_port_0, N0299_port_1, N0299_v;
  wire signed [`W-1:0] N0762_port_2, N0762_port_3, N0762_port_0, N0762_port_1, N0762_port_4, N0762_port_5, N0762_v;
  wire signed [`W-1:0] N0763_port_2, N0763_port_3, N0763_port_0, N0763_port_1, N0763_port_4, N0763_port_5, N0763_v;
  wire signed [`W-1:0] N0760_port_2, N0760_port_0, N0760_port_1, N0760_v;
  wire signed [`W-1:0] N0761_port_2, N0761_port_3, N0761_port_0, N0761_port_1, N0761_port_4, N0761_port_5, N0761_v;
  wire signed [`W-1:0] N0766_port_0, N0766_port_1, N0766_v;
  wire signed [`W-1:0] N0767_port_2, N0767_port_0, N0767_v;
  wire signed [`W-1:0] N0764_port_2, N0764_port_3, N0764_port_0, N0764_port_1, N0764_port_4, N0764_port_5, N0764_v;
  wire signed [`W-1:0] N0765_port_2, N0765_port_1, N0765_v;
  wire signed [`W-1:0] N0768_port_2, N0768_port_0, N0768_v;
  wire signed [`W-1:0] N0769_port_2, N0769_port_0, N0769_port_1, N0769_v;
  wire signed [`W-1:0] N0908_port_0, N0908_port_1, N0908_v;
  wire signed [`W-1:0] N0909_port_0, N0909_port_1, N0909_v;
  wire signed [`W-1:0] N0903_port_0, N0903_port_1, N0903_v;
  wire signed [`W-1:0] sync_port_0, sync_port_1, sync_v;
  wire signed [`W-1:0] N0904_port_0, N0904_port_1, N0904_v;
  wire signed [`W-1:0] N0905_port_0, N0905_port_1, N0905_v;
  wire signed [`W-1:0] SC_A12_CLK2_port_2, SC_A12_CLK2_port_3, SC_A12_CLK2_v;
  wire signed [`W-1:0] R3_2_port_1, R3_2_v;
  wire signed [`W-1:0] N0588_port_2, N0588_port_3, N0588_port_0, N0588_port_1, N0588_v;
  wire signed [`W-1:0] N0589_port_0, N0589_port_1, N0589_v;
  wire signed [`W-1:0] N0586_port_0, N0586_v;
  wire signed [`W-1:0] N0587_port_2, N0587_port_3, N0587_port_0, N0587_port_1, N0587_port_6, N0587_port_4, N0587_port_5, N0587_v;
  wire signed [`W-1:0] N0584_port_3, N0584_port_6, N0584_port_7, N0584_port_4, N0584_port_5, N0584_v;
  wire signed [`W-1:0] N0582_port_2, N0582_port_1, N0582_v;
  wire signed [`W-1:0] N0583_port_8, N0583_port_9, N0583_v;
  wire signed [`W-1:0] N0580_port_2, N0580_port_1, N0580_v;
  wire signed [`W-1:0] N0581_port_8, N0581_port_9, N0581_v;
  wire signed [`W-1:0] N0618_port_2, N0618_port_0, N0618_port_1, N0618_v;
  wire signed [`W-1:0] N0619_port_8, N0619_port_9, N0619_v;
  wire signed [`W-1:0] N0616_port_8, N0616_port_9, N0616_v;
  wire signed [`W-1:0] N0614_port_0, N0614_port_1, N0614_v;
  wire signed [`W-1:0] N0613_port_0, N0613_port_6, N0613_v;
  wire signed [`W-1:0] N0836_port_0, N0836_port_1, N0836_v;
  wire signed [`W-1:0] N0837_port_0, N0837_port_1, N0837_v;
  wire signed [`W-1:0] N0835_port_0, N0835_port_1, N0835_v;
  wire signed [`W-1:0] N0832_port_0, N0832_port_1, N0832_v;
  wire signed [`W-1:0] N0833_port_2, N0833_port_3, N0833_v;
  wire signed [`W-1:0] N0830_port_0, N0830_port_1, N0830_v;
  wire signed [`W-1:0] N0831_port_0, N0831_port_1, N0831_v;
  wire signed [`W-1:0] S00612_port_1, S00612_v;
  wire signed [`W-1:0] S00613_port_0, S00613_v;
  wire signed [`W-1:0] N0838_port_0, N0838_port_1, N0838_v;
  wire signed [`W-1:0] N0839_port_0, N0839_port_1, N0839_v;
  wire signed [`W-1:0] S00580_port_1, S00580_v;
  wire signed [`W-1:0] S00581_port_1, S00581_v;
  wire signed [`W-1:0] S00584_port_1, S00584_v;
  wire signed [`W-1:0] S00585_port_1, S00585_v;
  wire signed [`W-1:0] cm_ram2_port_0, cm_ram2_port_1, cm_ram2_v;
  wire signed [`W-1:0] S00725_port_0, S00725_v;
  wire signed [`W-1:0] R2_1_port_1, R2_1_v;
  wire signed [`W-1:0] R2_0_port_0, R2_0_v;
  wire signed [`W-1:0] R2_3_port_1, R2_3_v;
  wire signed [`W-1:0] R2_2_port_0, R2_2_v;
  wire signed [`W-1:0] R0_3_port_1, R0_3_v;
  wire signed [`W-1:0] R0_2_port_0, R0_2_v;
  wire signed [`W-1:0] R0_1_port_1, R0_1_v;
  wire signed [`W-1:0] R0_0_port_0, R0_0_v;
  wire signed [`W-1:0] SC_port_4, SC_port_13, SC_v;
  wire signed [`W-1:0] R1_0_port_1, R1_0_v;
  wire signed [`W-1:0] R1_1_port_0, R1_1_v;
  wire signed [`W-1:0] R6_1_port_1, R6_1_v;
  wire signed [`W-1:0] R6_0_port_0, R6_0_v;
  wire signed [`W-1:0] R6_3_port_1, R6_3_v;
  wire signed [`W-1:0] R6_2_port_0, R6_2_v;
  wire signed [`W-1:0] N0629_port_2, N0629_port_0, N0629_port_1, N0629_v;
  wire signed [`W-1:0] N0628_port_2, N0628_port_3, N0628_port_0, N0628_port_1, N0628_port_4, N0628_v;
  wire signed [`W-1:0] N0851_port_1, N0851_v;
  wire signed [`W-1:0] R4_3_port_1, R4_3_v;
  wire signed [`W-1:0] R4_2_port_0, R4_2_v;
  wire signed [`W-1:0] R4_1_port_1, R4_1_v;
  wire signed [`W-1:0] R4_0_port_0, R4_0_v;
  wire signed [`W-1:0] N0623_port_0, N0623_port_1, N0623_v;
  wire signed [`W-1:0] N0622_port_2, N0622_port_3, N0622_v;
  wire signed [`W-1:0] N0333_port_0, N0333_port_1, N0333_v;
  wire signed [`W-1:0] N0620_port_3, N0620_port_6, N0620_port_7, N0620_port_4, N0620_port_5, N0620_v;
  wire signed [`W-1:0] N0627_port_2, N0627_port_0, N0627_v;
  wire signed [`W-1:0] N0334_port_0, N0334_port_1, N0334_v;
  wire signed [`W-1:0] N0625_port_0, N0625_v;
  wire signed [`W-1:0] N0624_port_0, N0624_port_1, N0624_v;
  wire signed [`W-1:0] N0803_port_3, N0803_port_1, N0803_port_4, N0803_v;
  wire signed [`W-1:0] N0854_port_0, N0854_port_6, N0854_v;
  wire signed [`W-1:0] ADSR_port_2, ADSR_port_0, ADSR_port_1, ADSR_v;
  wire signed [`W-1:0] ADDR_PTR_1_port_2, ADDR_PTR_1_port_3, ADDR_PTR_1_port_0, ADDR_PTR_1_port_1, ADDR_PTR_1_v;
  wire signed [`W-1:0] ADDR_PTR_0_port_2, ADDR_PTR_0_port_3, ADDR_PTR_0_port_0, ADDR_PTR_0_port_1, ADDR_PTR_0_v;
  wire signed [`W-1:0] READ_ACC_3__port_8, READ_ACC_3__port_9, READ_ACC_3__port_2, READ_ACC_3__port_3, READ_ACC_3__port_0, READ_ACC_3__port_1, READ_ACC_3__port_6, READ_ACC_3__port_7, READ_ACC_3__port_4, READ_ACC_3__port_5, READ_ACC_3__v;
  wire signed [`W-1:0] L_port_2, L_port_0, L_port_1, L_port_5, L_v;
  wire signed [`W-1:0] N0856_port_2, N0856_port_3, N0856_port_0, N0856_port_1, N0856_v;
  wire signed [`W-1:0] N0857_port_2, N0857_port_3, N0857_port_1, N0857_port_4, N0857_v;
  wire signed [`W-1:0] _OPE_port_0, _OPE_port_1, _OPE_v;
  wire signed [`W-1:0] N0858_port_2, N0858_port_3, N0858_port_0, N0858_port_1, N0858_v;
  wire signed [`W-1:0] N0759_port_0, N0759_port_1, N0759_v;
  wire signed [`W-1:0] N0758_port_2, N0758_port_3, N0758_port_1, N0758_v;
  wire signed [`W-1:0] N0757_port_0, N0757_port_1, N0757_v;
  wire signed [`W-1:0] N0756_port_2, N0756_port_0, N0756_port_1, N0756_v;
  wire signed [`W-1:0] N0755_port_0, N0755_port_1, N0755_v;
  wire signed [`W-1:0] N0754_port_2, N0754_port_3, N0754_port_1, N0754_v;
  wire signed [`W-1:0] N0753_port_0, N0753_port_1, N0753_v;
  wire signed [`W-1:0] N0752_port_3, N0752_port_0, N0752_v;
  wire signed [`W-1:0] N0751_port_2, N0751_port_0, N0751_port_1, N0751_v;
  wire signed [`W-1:0] N0750_port_2, N0750_port_0, N0750_port_1, N0750_v;
  wire signed [`W-1:0] S00690_port_1, S00690_v;
  wire signed [`W-1:0] N0920_port_0, N0920_port_1, N0920_v;
  wire signed [`W-1:0] N0339_port_2, N0339_port_0, N0339_port_1, N0339_v;
  wire signed [`W-1:0] N0338_port_0, N0338_port_1, N0338_v;
  wire signed [`W-1:0] S00609_port_0, S00609_v;
  wire signed [`W-1:0] N0802_port_2, N0802_port_1, N0802_v;
  wire signed [`W-1:0] N0801_port_2, N0801_port_1, N0801_v;
  wire signed [`W-1:0] N0800_port_0, N0800_port_1, N0800_v;
  wire signed [`W-1:0] N0807_port_0, N0807_port_1, N0807_v;
  wire signed [`W-1:0] N0806_port_0, N0806_port_1, N0806_v;
  wire signed [`W-1:0] N0805_port_2, N0805_port_1, N0805_v;
  wire signed [`W-1:0] N0804_port_2, N0804_port_3, N0804_v;
  wire signed [`W-1:0] S00601_port_1, S00601_v;
  wire signed [`W-1:0] S00600_port_1, S00600_v;
  wire signed [`W-1:0] N0809_port_0, N0809_port_1, N0809_v;
  wire signed [`W-1:0] N0808_port_0, N0808_port_1, N0808_v;
  wire signed [`W-1:0] S00599_port_1, S00599_v;
  wire signed [`W-1:0] S00598_port_1, S00598_v;
  wire signed [`W-1:0] ADSL_port_2, ADSL_port_0, ADSL_port_1, ADSL_v;
  wire signed [`W-1:0] A32_port_8, A32_port_9, A32_port_6, A32_v;
  wire signed [`W-1:0] N0936_port_0, N0936_port_1, N0936_v;
  wire signed [`W-1:0] N0935_port_0, N0935_port_1, N0935_v;
  wire signed [`W-1:0] N0931_port_0, N0931_port_1, N0931_v;
  wire signed [`W-1:0] N0930_port_0, N0930_port_1, N0930_v;
  wire signed [`W-1:0] S00734_port_1, S00734_v;
  wire signed [`W-1:0] R9_2_port_1, R9_2_v;
  wire signed [`W-1:0] R9_3_port_0, R9_3_v;
  wire signed [`W-1:0] R9_0_port_1, R9_0_v;
  wire signed [`W-1:0] R9_1_port_0, R9_1_v;
  wire signed [`W-1:0] N0520_port_0, N0520_port_1, N0520_v;
  wire signed [`W-1:0] N0521_port_0, N0521_v;
  wire signed [`W-1:0] S00732_port_1, S00732_v;
  wire signed [`W-1:0] FIN_FIM_port_2, FIN_FIM_port_3, FIN_FIM_port_0, FIN_FIM_port_4, FIN_FIM_port_5, FIN_FIM_v;
  wire signed [`W-1:0] __POC_CLK2_X12_X32__INH_port_2, __POC_CLK2_X12_X32__INH_port_3, __POC_CLK2_X12_X32__INH_port_0, __POC_CLK2_X12_X32__INH_port_1, __POC_CLK2_X12_X32__INH_port_4, __POC_CLK2_X12_X32__INH_port_5, __POC_CLK2_X12_X32__INH_v;
  wire signed [`W-1:0] INC_ISZ_ADD_SUB_XCH_LD_port_2, INC_ISZ_ADD_SUB_XCH_LD_port_3, INC_ISZ_ADD_SUB_XCH_LD_port_4, INC_ISZ_ADD_SUB_XCH_LD_port_5, INC_ISZ_ADD_SUB_XCH_LD_v;
  wire signed [`W-1:0] M12_M22_CLK1__M11_M12__port_8, M12_M22_CLK1__M11_M12__port_9, M12_M22_CLK1__M11_M12__v;
  wire signed [`W-1:0] S00828_port_1, S00828_v;
  wire signed [`W-1:0] N0847_port_3, N0847_port_0, N0847_port_1, N0847_port_6, N0847_port_4, N0847_port_5, N0847_v;
  wire signed [`W-1:0] ACC_ADAC_port_3, ACC_ADAC_port_0, ACC_ADAC_port_1, ACC_ADAC_v;
  wire signed [`W-1:0] _OPA_1_port_8, _OPA_1_port_7, _OPA_1_v;
  wire signed [`W-1:0] IAC_port_2, IAC_port_3, IAC_port_0, IAC_port_1, IAC_port_4, IAC_port_5, IAC_v;
  wire signed [`W-1:0] ADD_ACC_port_2, ADD_ACC_port_0, ADD_ACC_port_1, ADD_ACC_v;
  wire signed [`W-1:0] N0281_port_1, N0281_v;
  wire signed [`W-1:0] N0283_port_1, N0283_v;
  wire signed [`W-1:0] N0282_port_1, N0282_v;
  wire signed [`W-1:0] ACC_3_port_3, ACC_3_port_0, ACC_3_port_1, ACC_3_port_4, ACC_3_v;
  wire signed [`W-1:0] ACC_2_port_2, ACC_2_port_3, ACC_2_port_0, ACC_2_port_4, ACC_2_v;
  wire signed [`W-1:0] ACC_1_port_3, ACC_1_port_0, ACC_1_port_1, ACC_1_port_4, ACC_1_v;
  wire signed [`W-1:0] ACC_0_port_8, ACC_0_port_9, ACC_0_port_2, ACC_0_port_1, ACC_0_port_6, ACC_0_port_7, ACC_0_port_4, ACC_0_port_5, ACC_0_port_10, ACC_0_v;
  wire signed [`W-1:0] N0285_port_1, N0285_v;
  wire signed [`W-1:0] N0287_port_1, N0287_v;
  wire signed [`W-1:0] N0945_port_3, N0945_port_4, N0945_v;
  wire signed [`W-1:0] cm_ram1_port_0, cm_ram1_port_1, cm_ram1_v;
  wire signed [`W-1:0] TCS_port_2, TCS_port_3, TCS_port_0, TCS_port_1, TCS_port_4, TCS_port_5, TCS_v;
  wire signed [`W-1:0] cm_ram3_port_0, cm_ram3_port_1, cm_ram3_v;
  wire signed [`W-1:0] SC_A22_port_3, SC_A22_port_4, SC_A22_v;
  wire signed [`W-1:0] TCC_port_2, TCC_port_3, TCC_port_0, TCC_port_1, TCC_port_4, TCC_port_5, TCC_v;
  wire signed [`W-1:0] REG_RFSH_2_port_2, REG_RFSH_2_port_3, REG_RFSH_2_port_0, REG_RFSH_2_port_1, REG_RFSH_2_v;
  wire signed [`W-1:0] REG_RFSH_1_port_2, REG_RFSH_1_port_3, REG_RFSH_1_port_0, REG_RFSH_1_port_1, REG_RFSH_1_v;
  wire signed [`W-1:0] REG_RFSH_0_port_2, REG_RFSH_0_port_3, REG_RFSH_0_port_0, REG_RFSH_0_port_1, REG_RFSH_0_v;
  wire signed [`W-1:0] N0748_port_2, N0748_port_1, N0748_v;
  wire signed [`W-1:0] N0749_port_2, N0749_port_0, N0749_port_1, N0749_v;
  wire signed [`W-1:0] N0740_port_2, N0740_port_1, N0740_v;
  wire signed [`W-1:0] N0741_port_0, N0741_port_1, N0741_v;
  wire signed [`W-1:0] N0742_port_2, N0742_port_1, N0742_v;
  wire signed [`W-1:0] N0743_port_2, N0743_port_1, N0743_v;
  wire signed [`W-1:0] N0744_port_2, N0744_port_1, N0744_v;
  wire signed [`W-1:0] N0745_port_2, N0745_port_1, N0745_v;
  wire signed [`W-1:0] N0746_port_2, N0746_port_1, N0746_v;
  wire signed [`W-1:0] N0747_port_2, N0747_port_1, N0747_v;
  wire signed [`W-1:0] N0670_port_3, N0670_port_0, N0670_port_4, N0670_v;
  wire signed [`W-1:0] CY_1_port_2, CY_1_port_3, CY_1_port_1, CY_1_port_6, CY_1_port_4, CY_1_v;
  wire signed [`W-1:0] N0674_port_2, N0674_port_0, N0674_port_1, N0674_v;
  wire signed [`W-1:0] N0676_port_0, N0676_port_1, N0676_v;
  wire signed [`W-1:0] N0677_port_0, N0677_port_1, N0677_v;
  wire signed [`W-1:0] N0634_port_8, N0634_port_9, N0634_v;
  wire signed [`W-1:0] N0635_port_3, N0635_port_6, N0635_port_7, N0635_port_4, N0635_port_5, N0635_v;
  wire signed [`W-1:0] N0636_port_2, N0636_port_3, N0636_port_1, N0636_port_4, N0636_port_5, N0636_v;
  wire signed [`W-1:0] N0637_port_2, N0637_port_0, N0637_port_1, N0637_v;
  wire signed [`W-1:0] N0630_port_2, N0630_port_1, N0630_v;
  wire signed [`W-1:0] N0631_port_0, N0631_port_1, N0631_v;
  wire signed [`W-1:0] N0632_port_8, N0632_port_9, N0632_v;
  wire signed [`W-1:0] N0633_port_0, N0633_v;
  wire signed [`W-1:0] N0638_port_0, N0638_port_1, N0638_v;
  wire signed [`W-1:0] N0639_port_0, N0639_port_1, N0639_v;
  wire signed [`W-1:0] N0329_port_0, N0329_port_1, N0329_v;
  wire signed [`W-1:0] N0322_port_2, N0322_port_1, N0322_port_4, N0322_v;
  wire signed [`W-1:0] N0323_port_2, N0323_port_0, N0323_port_1, N0323_v;
  wire signed [`W-1:0] N0320_port_0, N0320_port_1, N0320_v;
  wire signed [`W-1:0] N0321_port_0, N0321_port_1, N0321_v;
  wire signed [`W-1:0] N0326_port_2, N0326_port_3, N0326_port_1, N0326_port_4, N0326_port_5, N0326_v;
  wire signed [`W-1:0] N0324_port_0, N0324_port_1, N0324_v;
  wire signed [`W-1:0] N0325_port_6, N0325_v;
  wire signed [`W-1:0] ACB_IB_port_2, ACB_IB_port_0, ACB_IB_port_1, ACB_IB_v;
  wire signed [`W-1:0] N0818_port_0, N0818_port_1, N0818_v;
  wire signed [`W-1:0] N0814_port_0, N0814_port_1, N0814_v;
  wire signed [`W-1:0] R5_3_port_0, R5_3_v;
  wire signed [`W-1:0] A22_port_8, A22_port_9, A22_port_6, A22_port_5, A22_v;
  wire signed [`W-1:0] N0473_port_2, N0473_port_3, N0473_port_0, N0473_port_1, N0473_v;
  wire signed [`W-1:0] N0921_port_0, N0921_port_1, N0921_v;
  wire signed [`W-1:0] N0922_port_0, N0922_port_1, N0922_v;
  wire signed [`W-1:0] N0923_port_0, N0923_port_1, N0923_v;
  wire signed [`W-1:0] N0924_port_0, N0924_port_1, N0924_v;
  wire signed [`W-1:0] N0925_port_0, N0925_port_1, N0925_v;
  wire signed [`W-1:0] N0926_port_0, N0926_port_1, N0926_v;
  wire signed [`W-1:0] N0927_port_0, N0927_port_1, N0927_v;
  wire signed [`W-1:0] N0928_port_2, N0928_port_3, N0928_v;
  wire signed [`W-1:0] N0929_port_0, N0929_port_1, N0929_v;
  wire signed [`W-1:0] N0697_port_0, N0697_v;
  wire signed [`W-1:0] S00709_port_1, S00709_v;
  wire signed [`W-1:0] R5_1_port_0, R5_1_v;
  wire signed [`W-1:0] N0690_port_2, N0690_port_0, N0690_port_1, N0690_v;
  wire signed [`W-1:0] N0691_port_0, N0691_v;
  wire signed [`W-1:0] N0694_port_0, N0694_v;
  wire signed [`W-1:0] N0933_port_0, N0933_port_1, N0933_v;
  wire signed [`W-1:0] INH_port_2, INH_port_4, INH_v;
  wire signed [`W-1:0] N0913_port_2, N0913_port_0, N0913_port_1, N0913_v;
  wire signed [`W-1:0] N0912_port_2, N0912_port_0, N0912_port_1, N0912_v;
  wire signed [`W-1:0] S00564_port_0, S00564_v;
  wire signed [`W-1:0] N0932_port_0, N0932_port_1, N0932_v;
  wire signed [`W-1:0] N0916_port_0, N0916_port_1, N0916_v;
  wire signed [`W-1:0] N0693_port_2, N0693_port_3, N0693_port_1, N0693_v;
  wire signed [`W-1:0] N0820_port_2, N0820_port_3, N0820_v;
  wire signed [`W-1:0] PC1_1_port_1, PC1_1_v;
  wire signed [`W-1:0] PC1_2_port_0, PC1_2_v;
  wire signed [`W-1:0] PC1_3_port_1, PC1_3_v;
  wire signed [`W-1:0] PC1_4_port_1, PC1_4_v;
  wire signed [`W-1:0] PC1_5_port_0, PC1_5_v;
  wire signed [`W-1:0] PC1_6_port_1, PC1_6_v;
  wire signed [`W-1:0] PC1_7_port_0, PC1_7_v;
  wire signed [`W-1:0] PC1_8_port_0, PC1_8_v;
  wire signed [`W-1:0] PC1_9_port_1, PC1_9_v;
  wire signed [`W-1:0] N0822_port_0, N0822_port_1, N0822_v;
  wire signed [`W-1:0] PC3_6_port_1, PC3_6_v;
  wire signed [`W-1:0] PC3_7_port_0, PC3_7_v;
  wire signed [`W-1:0] PC3_4_port_1, PC3_4_v;
  wire signed [`W-1:0] PC3_5_port_0, PC3_5_v;
  wire signed [`W-1:0] PC3_2_port_0, PC3_2_v;
  wire signed [`W-1:0] PC3_3_port_1, PC3_3_v;
  wire signed [`W-1:0] PC3_0_port_0, PC3_0_v;
  wire signed [`W-1:0] PC3_1_port_1, PC3_1_v;
  wire signed [`W-1:0] S00803_port_1, S00803_v;
  wire signed [`W-1:0] PC3_8_port_0, PC3_8_v;
  wire signed [`W-1:0] PC3_9_port_1, PC3_9_v;
  wire signed [`W-1:0] N0900_port_2, N0900_port_3, N0900_port_0, N0900_port_1, N0900_v;
  wire signed [`W-1:0] N0353_port_2, N0353_port_1, N0353_v;
  wire signed [`W-1:0] N0352_port_0, N0352_port_1, N0352_v;
  wire signed [`W-1:0] N0351_port_2, N0351_port_0, N0351_port_1, N0351_v;
  wire signed [`W-1:0] N0350_port_0, N0350_port_1, N0350_v;
  wire signed [`W-1:0] N0608_port_2, N0608_port_0, N0608_port_1, N0608_v;
  wire signed [`W-1:0] N0355_port_3, N0355_port_0, N0355_port_1, N0355_v;
  wire signed [`W-1:0] N0354_port_2, N0354_port_3, N0354_port_0, N0354_port_1, N0354_port_4, N0354_port_5, N0354_v;
  wire signed [`W-1:0] N0605_port_0, N0605_port_1, N0605_v;
  wire signed [`W-1:0] N0604_port_0, N0604_port_1, N0604_v;
  wire signed [`W-1:0] N0607_port_0, N0607_port_1, N0607_v;
  wire signed [`W-1:0] ADC_CY_port_2, ADC_CY_port_3, ADC_CY_port_1, ADC_CY_v;
  wire signed [`W-1:0] OPR_3_port_14, OPR_3_port_15, OPR_3_v;
  wire signed [`W-1:0] N0852_port_1, N0852_v;
  wire signed [`W-1:0] N0938_port_2, N0938_port_3, N0938_v;
  wire signed [`W-1:0] N0824_port_0, N0824_port_1, N0824_v;
  wire signed [`W-1:0] ADD_IB_port_2, ADD_IB_port_0, ADD_IB_port_1, ADD_IB_v;
  wire signed [`W-1:0] N0823_port_0, N0823_port_1, N0823_v;
  wire signed [`W-1:0] PC2_9_port_1, PC2_9_v;
  wire signed [`W-1:0] PC2_8_port_0, PC2_8_v;
  wire signed [`W-1:0] PC2_7_port_0, PC2_7_v;
  wire signed [`W-1:0] PC2_6_port_1, PC2_6_v;
  wire signed [`W-1:0] PC2_5_port_0, PC2_5_v;
  wire signed [`W-1:0] PC2_4_port_1, PC2_4_v;
  wire signed [`W-1:0] PC2_3_port_1, PC2_3_v;
  wire signed [`W-1:0] PC2_2_port_0, PC2_2_v;
  wire signed [`W-1:0] PC2_1_port_1, PC2_1_v;
  wire signed [`W-1:0] PC2_0_port_0, PC2_0_v;
  wire signed [`W-1:0] N0793_port_0, N0793_port_1, N0793_v;
  wire signed [`W-1:0] N0792_port_0, N0792_port_1, N0792_v;
  wire signed [`W-1:0] N0791_port_0, N0791_port_1, N0791_v;
  wire signed [`W-1:0] N0790_port_0, N0790_port_1, N0790_v;
  wire signed [`W-1:0] N0797_port_2, N0797_port_1, N0797_v;
  wire signed [`W-1:0] N0796_port_0, N0796_port_1, N0796_v;
  wire signed [`W-1:0] N0795_port_0, N0795_port_1, N0795_v;
  wire signed [`W-1:0] N0794_port_0, N0794_port_1, N0794_v;
  wire signed [`W-1:0] N0829_port_0, N0829_port_1, N0829_v;
  wire signed [`W-1:0] N0799_port_0, N0799_port_1, N0799_v;
  wire signed [`W-1:0] N0798_port_0, N0798_port_1, N0798_v;
  wire signed [`W-1:0] N0828_port_0, N0828_port_1, N0828_v;
  wire signed [`W-1:0] __X31__CLK2__port_2, __X31__CLK2__port_1, __X31__CLK2__v;
  wire signed [`W-1:0] clk1_port_0, clk1_port_1, clk1_port_28, clk1_v;
  wire signed [`W-1:0] clk2_port_51, clk2_port_0, clk2_v;
  wire signed [`W-1:0] N0317_port_0, N0317_v;
  wire signed [`W-1:0] N0316_port_2, N0316_port_0, N0316_port_1, N0316_v;
  wire signed [`W-1:0] N0315_port_0, N0315_v;
  wire signed [`W-1:0] N0645_port_8, N0645_port_9, N0645_v;
  wire signed [`W-1:0] N0312_port_0, N0312_port_1, N0312_v;
  wire signed [`W-1:0] N0647_port_8, N0647_port_9, N0647_v;
  wire signed [`W-1:0] N0310_port_3, N0310_port_4, N0310_v;
  wire signed [`W-1:0] N0649_port_2, N0649_port_1, N0649_v;
  wire signed [`W-1:0] N0648_port_3, N0648_port_6, N0648_port_7, N0648_port_4, N0648_port_5, N0648_v;
  wire signed [`W-1:0] S00840_port_1, S00840_v;
  wire signed [`W-1:0] N0319_port_0, N0319_port_1, N0319_v;
  wire signed [`W-1:0] N0318_port_2, N0318_port_3, N0318_port_1, N0318_port_4, N0318_port_5, N0318_v;
  wire signed [`W-1:0] N0487_port_2, N0487_port_1, N0487_v;
  wire signed [`W-1:0] N0485_port_0, N0485_port_1, N0485_v;
  wire signed [`W-1:0] N0484_port_0, N0484_port_1, N0484_v;
  wire signed [`W-1:0] N0483_port_0, N0483_port_1, N0483_v;
  wire signed [`W-1:0] N0482_port_0, N0482_port_1, N0482_v;
  wire signed [`W-1:0] N0481_port_2, N0481_port_3, N0481_port_0, N0481_port_1, N0481_v;
  wire signed [`W-1:0] N0480_port_0, N0480_port_1, N0480_v;
  wire signed [`W-1:0] WADB2_port_6, WADB2_port_4, WADB2_port_5, WADB2_v;
  wire signed [`W-1:0] WADB1_port_6, WADB1_port_4, WADB1_port_5, WADB1_v;
  wire signed [`W-1:0] WADB0_port_6, WADB0_port_4, WADB0_port_5, WADB0_v;
  wire signed [`W-1:0] N0489_port_0, N0489_v;
  wire signed [`W-1:0] N0488_port_0, N0488_port_1, N0488_v;
  wire signed [`W-1:0] N0869_port_8, N0869_port_9, N0869_port_2, N0869_port_3, N0869_port_0, N0869_port_6, N0869_port_7, N0869_port_4, N0869_port_5, N0869_port_10, N0869_v;
  wire signed [`W-1:0] N0868_port_8, N0868_port_9, N0868_port_2, N0868_port_3, N0868_port_0, N0868_port_6, N0868_port_7, N0868_port_4, N0868_port_5, N0868_port_10, N0868_v;
  wire signed [`W-1:0] N0867_port_8, N0867_port_9, N0867_port_2, N0867_port_3, N0867_port_0, N0867_port_6, N0867_port_7, N0867_port_4, N0867_port_5, N0867_port_10, N0867_v;
  wire signed [`W-1:0] N0853_port_0, N0853_port_1, N0853_v;
  wire signed [`W-1:0] A12_port_9, A12_port_7, A12_port_10, A12_v;
  wire signed [`W-1:0] S00716_port_1, S00716_v;
  wire signed [`W-1:0] S00710_port_0, S00710_v;
  wire signed [`W-1:0] __INH__X32_CLK2_port_2, __INH__X32_CLK2_port_3, __INH__X32_CLK2_v;
  wire signed [`W-1:0] S00620_port_1, S00620_v;
  wire signed [`W-1:0] S00627_port_1, S00627_v;
  wire signed [`W-1:0] S00624_port_1, S00624_v;
  wire signed [`W-1:0] S00628_port_0, S00628_v;
  wire signed [`W-1:0] N0684_port_0, N0684_port_1, N0684_v;
  wire signed [`W-1:0] N0850_port_1, N0850_v;
  wire signed [`W-1:0] N0507_port_0, N0507_port_1, N0507_v;
  wire signed [`W-1:0] N0346_port_3, N0346_port_0, N0346_port_1, N0346_v;
  wire signed [`W-1:0] N0504_port_0, N0504_v;
  wire signed [`W-1:0] N0505_port_2, N0505_port_0, N0505_port_1, N0505_v;
  wire signed [`W-1:0] SC_M22_CLK2_port_3, SC_M22_CLK2_port_4, SC_M22_CLK2_v;
  wire signed [`W-1:0] N0503_port_2, N0503_port_0, N0503_port_1, N0503_v;
  wire signed [`W-1:0] N0500_port_1, N0500_v;
  wire signed [`W-1:0] N0501_port_0, N0501_port_1, N0501_v;
  wire signed [`W-1:0] ADD_0_port_2, ADD_0_port_3, ADD_0_port_1, ADD_0_port_4, ADD_0_port_5, ADD_0_v;
  wire signed [`W-1:0] _I_O_port_0, _I_O_port_1, _I_O_v;
  wire signed [`W-1:0] d0_port_2, d0_port_3, d0_port_0, d0_port_4, d0_port_5, d0_v;
  wire signed [`W-1:0] d1_port_2, d1_port_3, d1_port_0, d1_port_4, d1_port_5, d1_v;
  wire signed [`W-1:0] N0347_port_3, N0347_port_1, N0347_port_4, N0347_v;
  wire signed [`W-1:0] N1013_port_1, N1013_v;
  wire signed [`W-1:0] N1012_port_1, N1012_v;
  wire signed [`W-1:0] N1011_port_0, N1011_v;
  wire signed [`W-1:0] N1010_port_0, N1010_v;
  wire signed [`W-1:0] N1015_port_1, N1015_v;
  wire signed [`W-1:0] N1014_port_1, N1014_v;
  wire signed [`W-1:0] R15_0_port_1, R15_0_v;
  wire signed [`W-1:0] R15_1_port_0, R15_1_v;
  wire signed [`W-1:0] R15_2_port_1, R15_2_v;
  wire signed [`W-1:0] R15_3_port_0, R15_3_v;
  wire signed [`W-1:0] N0937_port_0, N0937_port_1, N0937_port_6, N0937_v;
  wire signed [`W-1:0] R11_0_port_1, R11_0_v;
  wire signed [`W-1:0] R11_1_port_0, R11_1_v;
  wire signed [`W-1:0] R11_2_port_1, R11_2_v;
  wire signed [`W-1:0] R11_3_port_0, R11_3_v;
  wire signed [`W-1:0] R13_2_port_1, R13_2_v;
  wire signed [`W-1:0] R13_3_port_0, R13_3_v;
  wire signed [`W-1:0] R13_0_port_1, R13_0_v;
  wire signed [`W-1:0] R13_1_port_0, R13_1_v;
  wire signed [`W-1:0] OPR_1_port_9, OPR_1_port_10, OPR_1_v;
  wire signed [`W-1:0] OPR_0_port_3, OPR_0_port_6, OPR_0_v;
  wire signed [`W-1:0] OPR_2_port_8, OPR_2_port_14, OPR_2_v;
  wire signed [`W-1:0] N0340_port_2, N0340_port_0, N0340_v;
  wire signed [`W-1:0] N0859_port_2, N0859_port_3, N0859_port_1, N0859_port_4, N0859_v;
  wire signed [`W-1:0] N0688_port_0, N0688_v;
  wire signed [`W-1:0] N0788_port_0, N0788_port_1, N0788_v;
  wire signed [`W-1:0] N0789_port_0, N0789_port_1, N0789_v;
  wire signed [`W-1:0] N0784_port_0, N0784_port_1, N0784_v;
  wire signed [`W-1:0] N0785_port_0, N0785_port_1, N0785_v;
  wire signed [`W-1:0] N0786_port_0, N0786_port_1, N0786_v;
  wire signed [`W-1:0] N0787_port_0, N0787_port_1, N0787_v;
  wire signed [`W-1:0] N0780_port_2, N0780_port_3, N0780_port_0, N0780_port_6, N0780_port_4, N0780_port_5, N0780_v;
  wire signed [`W-1:0] N0781_port_2, N0781_port_3, N0781_port_0, N0781_port_6, N0781_port_4, N0781_port_5, N0781_v;
  wire signed [`W-1:0] N0782_port_2, N0782_port_3, N0782_port_4, N0782_port_5, N0782_v;
  wire signed [`W-1:0] N0783_port_2, N0783_port_3, N0783_v;
  wire signed [`W-1:0] N0300_port_3, N0300_port_4, N0300_v;
  wire signed [`W-1:0] N0301_port_2, N0301_port_3, N0301_v;
  wire signed [`W-1:0] N0302_port_0, N0302_port_1, N0302_v;
  wire signed [`W-1:0] N0303_port_0, N0303_port_1, N0303_v;
  wire signed [`W-1:0] N0304_port_2, N0304_port_3, N0304_port_1, N0304_v;
  wire signed [`W-1:0] N0305_port_2, N0305_port_0, N0305_port_1, N0305_v;
  wire signed [`W-1:0] N0306_port_0, N0306_port_1, N0306_v;
  wire signed [`W-1:0] N0307_port_3, N0307_port_4, N0307_port_5, N0307_v;
  wire signed [`W-1:0] N0308_port_0, N0308_port_1, N0308_v;
  wire signed [`W-1:0] N0309_port_0, N0309_port_1, N0309_v;
  wire signed [`W-1:0] N0658_port_3, N0658_port_0, N0658_port_1, N0658_v;
  wire signed [`W-1:0] N0659_port_4, N0659_port_5, N0659_v;
  wire signed [`W-1:0] N0490_port_2, N0490_port_0, N0490_v;
  wire signed [`W-1:0] N0491_port_0, N0491_port_1, N0491_v;
  wire signed [`W-1:0] N0492_port_0, N0492_v;
  wire signed [`W-1:0] N0493_port_0, N0493_port_1, N0493_v;
  wire signed [`W-1:0] N0494_port_2, N0494_port_0, N0494_v;
  wire signed [`W-1:0] N0495_port_0, N0495_port_1, N0495_v;
  wire signed [`W-1:0] N0496_port_0, N0496_port_1, N0496_v;
  wire signed [`W-1:0] N0497_port_0, N0497_v;
  wire signed [`W-1:0] N0498_port_1, N0498_v;
  wire signed [`W-1:0] N0499_port_0, N0499_v;
  wire signed [`W-1:0] N0878_port_2, N0878_port_3, N0878_port_4, N0878_v;
  wire signed [`W-1:0] N0879_port_3, N0879_port_1, N0879_port_4, N0879_v;
  wire signed [`W-1:0] N0653_port_0, N0653_v;
  wire signed [`W-1:0] N0651_port_0, N0651_port_1, N0651_v;
  wire signed [`W-1:0] N0656_port_0, N0656_port_1, N0656_v;
  wire signed [`W-1:0] X12_port_10, X12_port_12, X12_port_13, X12_port_15, X12_v;
  wire signed [`W-1:0] N0657_port_8, N0657_port_9, N0657_v;
  wire signed [`W-1:0] N0654_port_2, N0654_port_0, N0654_port_1, N0654_v;
  wire signed [`W-1:0] N0655_port_2, N0655_port_1, N0655_v;
  wire signed [`W-1:0] S00762_port_1, S00762_v;
  wire signed [`W-1:0] RAL_port_2, RAL_port_3, RAL_port_0, RAL_port_1, RAL_port_4, RAL_port_5, RAL_v;
  wire signed [`W-1:0] RAR_port_2, RAR_port_3, RAR_port_0, RAR_port_1, RAR_port_4, RAR_port_5, RAR_v;
  wire signed [`W-1:0] N0716_port_2, N0716_port_3, N0716_port_0, N0716_port_1, N0716_port_4, N0716_v;
  wire signed [`W-1:0] N0313_port_0, N0313_port_1, N0313_v;
  wire signed [`W-1:0] OPA_2_port_0, OPA_2_port_4, OPA_2_port_13, OPA_2_v;
  wire signed [`W-1:0] OPA_3_port_2, OPA_3_port_0, OPA_3_port_13, OPA_3_v;
  wire signed [`W-1:0] OPA_0_port_11, OPA_0_port_12, OPA_0_port_13, OPA_0_v;
  wire signed [`W-1:0] _INH_port_0, _INH_port_1, _INH_v;
  wire signed [`W-1:0] N0934_port_0, N0934_port_1, N0934_v;
  wire signed [`W-1:0] STC_port_2, STC_port_3, STC_port_0, STC_port_1, STC_port_4, STC_port_5, STC_v;
  wire signed [`W-1:0] N0873_port_0, N0873_port_4, N0873_port_5, N0873_v;
  wire signed [`W-1:0] N0870_port_2, N0870_port_0, N0870_port_6, N0870_v;
  wire signed [`W-1:0] FIN_FIM_SRC_JIN_port_3, FIN_FIM_SRC_JIN_port_6, FIN_FIM_SRC_JIN_port_4, FIN_FIM_SRC_JIN_port_5, FIN_FIM_SRC_JIN_v;
  wire signed [`W-1:0] N0871_port_0, N0871_port_6, N0871_port_5, N0871_v;
  wire signed [`W-1:0] N0876_port_2, N0876_port_1, N0876_v;
  wire signed [`W-1:0] N0877_port_2, N0877_port_3, N0877_port_4, N0877_v;
  wire signed [`W-1:0] N0874_port_2, N0874_port_1, N0874_v;
  wire signed [`W-1:0] N1008_port_1, N1008_v;
  wire signed [`W-1:0] N1009_port_0, N1009_v;
  wire signed [`W-1:0] N1004_port_3, N1004_port_4, N1004_v;
  wire signed [`W-1:0] N1005_port_2, N1005_port_3, N1005_v;
  wire signed [`W-1:0] N1006_port_3, N1006_port_4, N1006_v;
  wire signed [`W-1:0] N1007_port_2, N1007_port_3, N1007_v;
  wire signed [`W-1:0] N1000_port_3, N1000_port_4, N1000_v;
  wire signed [`W-1:0] N1001_port_2, N1001_port_3, N1001_v;
  wire signed [`W-1:0] N1002_port_3, N1002_port_4, N1002_v;
  wire signed [`W-1:0] N1003_port_2, N1003_port_3, N1003_v;
  wire signed [`W-1:0] OPA_1_port_10, OPA_1_port_11, OPA_1_port_12, OPA_1_v;
  wire signed [`W-1:0] PC3_10_port_0, PC3_10_v;
  wire signed [`W-1:0] PC3_11_port_1, PC3_11_v;
  wire signed [`W-1:0] FIM_SRC_port_2, FIM_SRC_port_3, FIM_SRC_port_0, FIM_SRC_port_1, FIM_SRC_port_4, FIM_SRC_v;
  wire signed [`W-1:0] ADDR_RFSH_1_port_2, ADDR_RFSH_1_port_3, ADDR_RFSH_1_port_0, ADDR_RFSH_1_port_1, ADDR_RFSH_1_v;
  wire signed [`W-1:0] ADDR_RFSH_0_port_2, ADDR_RFSH_0_port_3, ADDR_RFSH_0_port_0, ADDR_RFSH_0_port_1, ADDR_RFSH_0_v;
  wire signed [`W-1:0] S00778_port_0, S00778_v;
  wire signed [`W-1:0] N0375_port_3, N0375_port_0, N0375_port_1, N0375_v;
  wire signed [`W-1:0] N0374_port_1, N0374_v;
  wire signed [`W-1:0] N0696_port_2, N0696_port_3, N0696_port_0, N0696_v;
  wire signed [`W-1:0] N0377_port_0, N0377_port_1, N0377_v;
  wire signed [`W-1:0] N0376_port_2, N0376_port_3, N0376_port_0, N0376_port_1, N0376_port_4, N0376_port_5, N0376_v;
  wire signed [`W-1:0] N0278_port_1, N0278_v;
  wire signed [`W-1:0] N0279_port_2, N0279_port_3, N0279_port_0, N0279_port_1, N0279_v;
  wire signed [`W-1:0] DCL_1_port_2, DCL_1_port_3, DCL_1_port_1, DCL_1_v;
  wire signed [`W-1:0] DCL_0_port_3, DCL_0_port_0, DCL_0_port_4, DCL_0_v;
  wire signed [`W-1:0] DCL_2_port_2, DCL_2_port_3, DCL_2_port_1, DCL_2_v;
  wire signed [`W-1:0] N0373_port_2, N0373_port_3, N0373_port_0, N0373_port_1, N0373_v;
  wire signed [`W-1:0] N0372_port_2, N0372_port_3, N0372_port_0, N0372_port_1, N0372_v;
  wire signed [`W-1:0] N0669_port_3, N0669_port_0, N0669_port_1, N0669_v;
  wire signed [`W-1:0] N0667_port_2, N0667_port_0, N0667_port_1, N0667_v;
  wire signed [`W-1:0] N0666_port_2, N0666_port_3, N0666_port_4, N0666_v;
  wire signed [`W-1:0] N0665_port_2, N0665_port_0, N0665_port_1, N0665_v;
  wire signed [`W-1:0] N0664_port_2, N0664_port_1, N0664_port_4, N0664_v;
  wire signed [`W-1:0] N0663_port_2, N0663_port_3, N0663_port_1, N0663_v;
  wire signed [`W-1:0] N0662_port_0, N0662_port_1, N0662_v;
  wire signed [`W-1:0] N0661_port_0, N0661_port_1, N0661_v;
  wire signed [`W-1:0] N0660_port_0, N0660_port_1, N0660_v;
  wire signed [`W-1:0] N0469_port_0, N0469_port_1, N0469_port_4, N0469_v;
  wire signed [`W-1:0] N0468_port_2, N0468_port_3, N0468_port_0, N0468_port_1, N0468_v;
  wire signed [`W-1:0] N0465_port_0, N0465_port_1, N0465_v;
  wire signed [`W-1:0] N0464_port_2, N0464_port_3, N0464_port_4, N0464_v;
  wire signed [`W-1:0] PC1_10_port_0, PC1_10_v;
  wire signed [`W-1:0] PC1_11_port_1, PC1_11_v;
  wire signed [`W-1:0] N0461_port_2, N0461_port_1, N0461_port_4, N0461_v;
  wire signed [`W-1:0] N0460_port_0, N0460_port_1, N0460_v;
  wire signed [`W-1:0] N0463_port_2, N0463_port_3, N0463_port_6, N0463_v;
  wire signed [`W-1:0] N0462_port_0, N0462_port_1, N0462_v;
  wire signed [`W-1:0] N0685_port_0, N0685_v;
  wire signed [`W-1:0] N0687_port_2, N0687_port_0, N0687_port_1, N0687_v;
  wire signed [`W-1:0] N0681_port_0, N0681_port_1, N0681_v;
  wire signed [`W-1:0] N0680_port_0, N0680_port_1, N0680_v;
  wire signed [`W-1:0] N0683_port_2, N0683_port_0, N0683_port_1, N0683_v;
  wire signed [`W-1:0] S00557_port_1, S00557_v;
  wire signed [`W-1:0] N0689_port_2, N0689_port_0, N0689_port_1, N0689_v;
  wire signed [`W-1:0] X22_port_6, X22_port_7, X22_port_5, X22_v;
  wire signed [`W-1:0] N0398_port_0, N0398_port_1, N0398_v;
  wire signed [`W-1:0] R12_2_port_0, R12_2_v;
  wire signed [`W-1:0] R12_1_port_1, R12_1_v;
  wire signed [`W-1:0] N0846_port_2, N0846_port_0, N0846_port_1, N0846_port_6, N0846_port_4, N0846_port_5, N0846_v;
  wire signed [`W-1:0] N0843_port_0, N0843_port_1, N0843_v;
  wire signed [`W-1:0] N0841_port_0, N0841_port_1, N0841_v;
  wire signed [`W-1:0] N0840_port_0, N0840_port_1, N0840_v;
  wire signed [`W-1:0] N0519_port_0, N0519_v;
  wire signed [`W-1:0] N0518_port_0, N0518_port_1, N0518_v;
  wire signed [`W-1:0] N0692_port_2, N0692_port_0, N0692_port_1, N0692_v;
  wire signed [`W-1:0] OPE_port_2, OPE_port_3, OPE_port_0, OPE_port_1, OPE_port_4, OPE_v;
  wire signed [`W-1:0] N0695_port_2, N0695_port_3, N0695_port_1, N0695_v;
  wire signed [`W-1:0] N0686_port_0, N0686_port_1, N0686_v;
  wire signed [`W-1:0] JCN_port_2, JCN_port_3, JCN_port_0, JCN_port_1, JCN_port_4, JCN_v;
  wire signed [`W-1:0] N0678_port_3, N0678_port_0, N0678_port_1, N0678_port_4, N0678_v;
  wire signed [`W-1:0] N0679_port_2, N0679_port_0, N0679_v;
  wire signed [`W-1:0] N0671_port_2, N0671_port_0, N0671_port_1, N0671_v;
  wire signed [`W-1:0] N0672_port_2, N0672_port_0, N0672_port_1, N0672_v;
  wire signed [`W-1:0] N0673_port_2, N0673_port_0, N0673_port_1, N0673_v;
  wire signed [`W-1:0] N0675_port_2, N0675_port_3, N0675_port_0, N0675_v;
  wire signed [`W-1:0] N0478_port_2, N0478_port_3, N0478_port_0, N0478_port_1, N0478_port_4, N0478_v;
  wire signed [`W-1:0] N0479_port_2, N0479_port_0, N0479_v;
  wire signed [`W-1:0] N0476_port_2, N0476_port_0, N0476_v;
  wire signed [`W-1:0] N0477_port_2, N0477_port_0, N0477_port_1, N0477_v;
  wire signed [`W-1:0] N0474_port_2, N0474_port_3, N0474_port_0, N0474_port_1, N0474_v;
  wire signed [`W-1:0] N0475_port_0, N0475_port_1, N0475_port_4, N0475_v;
  wire signed [`W-1:0] N0472_port_2, N0472_port_3, N0472_port_0, N0472_port_1, N0472_v;
  wire signed [`W-1:0] N0470_port_2, N0470_port_3, N0470_port_0, N0470_port_1, N0470_v;
  wire signed [`W-1:0] N0471_port_2, N0471_port_3, N0471_port_0, N0471_port_1, N0471_v;
  wire signed [`W-1:0] X32_port_11, X32_port_12, X32_v;
  wire signed [`W-1:0] N0698_port_2, N0698_port_3, N0698_port_1, N0698_v;
  wire signed [`W-1:0] N0699_port_1, N0699_v;
  wire signed [`W-1:0] CLK2_JMS_DC_M22_BBL_M22_X12_X22___port_2, CLK2_JMS_DC_M22_BBL_M22_X12_X22___port_3, CLK2_JMS_DC_M22_BBL_M22_X12_X22___port_4, CLK2_JMS_DC_M22_BBL_M22_X12_X22___v;
  wire signed [`W-1:0] N0506_port_0, N0506_v;
  wire signed [`W-1:0] N0508_port_0, N0508_port_1, N0508_v;
  wire signed [`W-1:0] N0509_port_0, N0509_port_1, N0509_v;
  wire signed [`W-1:0] S00740_port_0, S00740_v;
  wire signed [`W-1:0] N0328_port_2, N0328_port_0, N0328_port_1, N0328_v;
  wire signed [`W-1:0] S00766_port_0, S00766_v;
  wire signed [`W-1:0] N0551_port_2, N0551_port_0, N0551_port_1, N0551_v;
  wire signed [`W-1:0] S00767_port_0, S00767_v;
  wire signed [`W-1:0] N0550_port_2, N0550_port_3, N0550_port_0, N0550_port_1, N0550_v;
  wire signed [`W-1:0] N0327_port_3, N0327_port_0, N0327_port_4, N0327_v;
  wire signed [`W-1:0] S00764_port_1, S00764_v;
  wire signed [`W-1:0] N0553_port_2, N0553_port_1, N0553_v;
  wire signed [`W-1:0] N0955_port_2, N0955_port_3, N0955_v;
  wire signed [`W-1:0] N0954_port_0, N0954_port_1, N0954_v;
  wire signed [`W-1:0] N0957_port_0, N0957_port_1, N0957_v;
  wire signed [`W-1:0] S00765_port_0, S00765_v;
  wire signed [`W-1:0] N0552_port_2, N0552_port_0, N0552_port_1, N0552_v;
  wire signed [`W-1:0] N0819_port_2, N0819_port_0, N0819_port_1, N0819_v;
  wire signed [`W-1:0] DAA_port_2, DAA_port_3, DAA_port_0, DAA_port_1, DAA_port_4, DAA_port_5, DAA_v;
  wire signed [`W-1:0] DAC_port_2, DAC_port_3, DAC_port_0, DAC_port_1, DAC_port_4, DAC_port_5, DAC_v;
  wire signed [`W-1:0] _SRC_port_0, _SRC_port_1, _SRC_v;
  wire signed [`W-1:0] N0529_port_8, N0529_port_9, N0529_v;
  wire signed [`W-1:0] N0815_port_0, N0815_port_1, N0815_v;
  wire signed [`W-1:0] N0555_port_2, N0555_port_0, N0555_port_1, N0555_v;
  wire signed [`W-1:0] N0816_port_0, N0816_port_1, N0816_v;
  wire signed [`W-1:0] __FIN_X12__port_2, __FIN_X12__port_3, __FIN_X12__v;
  wire signed [`W-1:0] JUN_JMS_port_8, JUN_JMS_port_7, JUN_JMS_port_4, JUN_JMS_port_5, JUN_JMS_v;
  wire signed [`W-1:0] N0810_port_0, N0810_port_1, N0810_v;
  wire signed [`W-1:0] S00835_port_0, S00835_v;
  wire signed [`W-1:0] N0812_port_0, N0812_port_1, N0812_v;
  wire signed [`W-1:0] N0554_port_2, N0554_port_0, N0554_port_1, N0554_v;
  wire signed [`W-1:0] N0813_port_0, N0813_port_1, N0813_v;
  wire signed [`W-1:0] PC0_11_port_1, PC0_11_v;
  wire signed [`W-1:0] PC0_10_port_0, PC0_10_v;
  wire signed [`W-1:0] N0557_port_2, N0557_port_0, N0557_port_1, N0557_v;


  spice_pin_input pin_2245(reset, reset_v, reset_port_2);
  spice_pin_input pin_2242(clk1, clk1_v, clk1_port_28);
  spice_pin_input pin_2246(test, test_v, test_port_2);
  spice_pin_input pin_2243(clk2, clk2_v, clk2_port_51);

  spice_pin_output pin_2253(cm_ram2, cm_ram2_v);
  spice_pin_output pin_2252(cm_ram3, cm_ram3_v);
  spice_pin_output pin_2251(cm_rom, cm_rom_v);
  spice_pin_output pin_2244(sync, sync_v);
  spice_pin_output pin_2255(cm_ram0, cm_ram0_v);
  spice_pin_output pin_2254(cm_ram1, cm_ram1_v);

  spice_pin_bidirectional pin_2247(d0_i, d0_o, d0_t, d0_v, d0_port_5);
  spice_pin_bidirectional pin_2248(d1_i, d1_o, d1_t, d1_v, d1_port_5);
  spice_pin_bidirectional pin_2249(d2_i, d2_o, d2_t, d2_v, d2_port_5);
  spice_pin_bidirectional pin_2250(d3_i, d3_o, d3_t, d3_v, d3_port_5);

  spice_transistor_nmos_vdd tM3268(v(S00839_v), N0698_v, N0698_port_3);
  spice_transistor_nmos_gnd tM2689(v(N1014_v), N1004_v, N1004_port_3);
  spice_transistor_nmos_gnd tM2688(v(N1012_v), N1000_v, N1000_port_3);
  spice_transistor_nmos tM1190(v(N0426_v), N0390_v, PC2_10_v, N0390_port_4, PC2_10_port_0);
  spice_transistor_nmos_gnd tM1935(v(X22_v), N0511_v, N0511_port_3);
  spice_transistor_nmos_gnd tM2926(v(N0875_v), N0884_v, N0884_port_1);
  spice_transistor_nmos_gnd tM1949(v(N0600_v), N0610_v, N0610_port_3);
  spice_transistor_nmos_gnd tM1948(v(clk2_v), N0460_v, N0460_port_1);
  spice_transistor_nmos tM1944(v(DC_v), N0467_v, N0484_v, N0467_port_2, N0484_port_1);
  spice_transistor_nmos tM1947(v(clk2_v), N0592_v, N0588_v, N0592_port_1, N0588_port_1);
  spice_transistor_nmos tM1940(v(N0528_v), N0526_v, N0527_v, N0526_port_1, N0527_port_0);
  spice_transistor_nmos_gnd tM1936(v(DC_v), N0526_v, N0526_port_0);
  spice_transistor_nmos_gnd tM1942(v(JMS_v), N0485_v, N0485_port_0);
  spice_transistor_nmos tM1383(v(N0434_v), N0830_v, N0781_v, N0830_port_0, N0781_port_4);
  spice_transistor_nmos tM1382(v(N0424_v), N0781_v, N0815_v, N0781_port_3, N0815_port_1);
  spice_transistor_nmos tM1381(v(N0406_v), N0795_v, N0777_v, N0795_port_1, N0777_port_2);
  spice_transistor_nmos_gnd tM1380(v(N0306_v), N0314_v, N0314_port_0);
  spice_transistor_nmos_gnd tM1387(v(PC1_4_v), N0816_v, N0816_port_0);
  spice_transistor_nmos_gnd tM1386(v(PC3_0_v), N0843_v, N0843_port_0);
  spice_transistor_nmos tM1385(v(N0439_v), PC3_0_v, N0394_v, PC3_0_port_0, N0394_port_5);
  spice_transistor_nmos_gnd tM1384(v(PC2_0_v), N0830_v, N0830_port_1);
  spice_transistor_nmos_gnd tM1389(v(N0773_v), N0396_v, N0396_port_1);
  spice_transistor_nmos tM1388(v(N0424_v), N0777_v, N0816_v, N0777_port_3, N0816_port_1);
  spice_transistor_nmos_gnd tM3157(v(N0735_v), cm_ram2_v, cm_ram2_port_1);
  spice_transistor_nmos tM1203(v(WADB0_v), N0780_v, N0763_v, N0780_port_0, N0763_port_5);
  spice_transistor_nmos_gnd tM1200(v(PC2_10_v), N0826_v, N0826_port_1);
  spice_transistor_nmos_gnd tM3095(v(POC_v), DCL_2_v, DCL_2_port_3);
  spice_transistor_nmos_vdd tM1201(v(__INH__X11_X31_CLK1_v), N0775_v, N0775_port_6);
  spice_transistor_nmos tM1206(v(N0381_v), N0391_v, PC0_9_v, N0391_port_2, PC0_9_port_1);
  spice_transistor_nmos_gnd tM1207(v(PC1_9_v), N0812_v, N0812_port_0);
  spice_transistor_nmos_gnd tM3096(v(DCL_2_v), N0749_v, N0749_port_1);
  spice_transistor_nmos tM1204(v(WADB0_v), N0781_v, N0764_v, N0781_port_0, N0764_port_3);
  spice_transistor_nmos_gnd tM1169(v(R11_0_v), N0966_v, N0966_port_0);
  spice_transistor_nmos_gnd tM1168(v(R9_0_v), N0956_v, N0956_port_1);
  spice_transistor_nmos tM1167(v(N0616_v), N0956_v, N0866_v, N0956_port_0, N0866_port_6);
  spice_transistor_nmos tM1166(v(N0591_v), N0866_v, N0947_v, N0866_port_5, N0947_port_1);
  spice_transistor_nmos_gnd tM1165(v(R7_0_v), N0947_v, N0947_port_0);
  spice_transistor_nmos_gnd tM1164(v(R5_0_v), N0929_v, N0929_port_1);
  spice_transistor_nmos tM1163(v(N0581_v), N0929_v, N0866_v, N0929_port_0, N0866_port_4);
  spice_transistor_nmos tM1162(v(N0565_v), N0866_v, N0920_v, N0866_port_3, N0920_port_1);
  spice_transistor_nmos_gnd tM1161(v(R3_0_v), N0920_v, N0920_port_0);
  spice_transistor_nmos_gnd tM1160(v(R1_0_v), N0903_v, N0903_port_1);
  spice_transistor_nmos_gnd tM1562(v(N0530_v), N0902_v, N0902_port_3);
  spice_transistor_nmos tM1561(v(N0584_v), N0591_v, __POC__CLK2_SC_A32_X12__v, N0591_port_9, __POC__CLK2_SC_A32_X12__port_3);
  spice_transistor_nmos tM1541(v(N0434_v), N0832_v, N0773_v, N0832_port_0, N0773_port_4);
  spice_transistor_nmos tM1540(v(N0424_v), N0773_v, N0817_v, N0773_port_3, N0817_port_1);
  spice_transistor_nmos_gnd tM1543(v(PC2_8_v), N0832_v, N0832_port_1);
  spice_transistor_nmos tM1545(v(N0444_v), N0773_v, N0845_v, N0773_port_5, N0845_port_1);
  spice_transistor_nmos_gnd tM1549(v(N0489_v), N0488_v, N0488_port_1);
  spice_transistor_nmos_gnd tM2945(v(N0871_v), N0899_v, N0899_port_0);
  spice_transistor_nmos_gnd tM1742(v(N0401_v), N0382_v, N0382_port_4);
  spice_transistor_nmos_gnd tM2016(v(DC_v), N0597_v, N0597_port_0);
  spice_transistor_nmos tM2017(v(FIN_FIM_SRC_JIN_v), N0597_v, N0596_v, N0597_port_1, N0596_port_0);
  spice_transistor_nmos_gnd tM2014(v(FIN_FIM_SRC_JIN_v), N0602_v, N0602_port_2);
  spice_transistor_nmos_gnd tM2015(v(_OPA_0_v), N0580_v, N0580_port_1);
  spice_transistor_nmos_gnd tM2012(v(SC_v), N0612_v, N0612_port_0);
  spice_transistor_nmos_gnd tM1037(v(N0298_v), N0756_v, N0756_port_2);
  spice_transistor_nmos_gnd tM2010(v(N0636_v), N0640_v, N0640_port_1);
  spice_transistor_nmos_gnd tM2011(v(INC_ISZ_ADD_SUB_XCH_LD_v), N0614_v, N0614_port_1);
  spice_transistor_nmos_vdd tM1769(v(S00581_v), N0584_v, N0584_port_7);
  spice_transistor_nmos_vdd tM1761(v(S00578_v), N0530_v, N0530_port_4);
  spice_transistor_nmos tM1760(v(N0466_v), N0464_v, N0465_v, N0464_port_4, N0465_port_1);
  spice_transistor_nmos_vdd tM1763(v(S00579_v), N0545_v, N0545_port_7);
  spice_transistor_nmos_vdd tM1764(v(S00580_v), N0570_v, N0570_port_7);
  spice_transistor_nmos_gnd tM2492(v(OPA_0_v), DAC_v, DAC_port_5);
  spice_transistor_nmos_vdd tM2493(v(N1002_v), _OPA_2_v, _OPA_2_port_7);
  spice_transistor_nmos_gnd tM2490(v(OPA_0_v), KBP_v, KBP_port_5);
  spice_transistor_nmos_gnd tM2496(v(OPA_0_v), STC_v, STC_port_5);
  spice_transistor_nmos_gnd tM1745(v(N0420_v), N0440_v, N0440_port_4);
  spice_transistor_nmos_gnd tM2494(v(N1004_v), OPA_1_v, OPA_1_port_10);
  spice_transistor_nmos_gnd tM2495(v(OPA_0_v), CMA_v, CMA_port_5);
  spice_transistor_nmos_gnd tM2498(v(OPA_0_v), CLB_v, CLB_port_5);
  spice_transistor_nmos_vdd tM1032(v(N0325_v), N0298_v, N0298_port_0);
  spice_transistor_nmos_vdd tM3252(v(N0696_v), d0_v, d0_port_2);
  spice_transistor_nmos_vdd tM2702(v(N0659_v), D0_v, D0_port_9);
  spice_transistor_nmos_gnd tM2703(v(N0700_v), N0687_v, N0687_port_1);
  spice_transistor_nmos_vdd tM2700(v(S00689_v), N0689_v, N0689_port_0);
  spice_transistor_nmos tM2707(v(SC_M22_CLK2_v), D0_v, N1015_v, D0_port_10, N1015_port_1);
  spice_transistor_nmos_gnd tM2704(v(N0700_v), N0689_v, N0689_port_1);
  spice_transistor_nmos_vdd tM2708(v(N0659_v), D2_v, D2_port_10);
  spice_transistor_nmos tM2032(v(_OPA_0_v), N0596_v, N0590_v, N0596_port_1, N0590_port_1);
  spice_transistor_nmos tM2034(v(N0564_v), N0563_v, N0562_v, N0563_port_0, N0562_port_0);
  spice_transistor_nmos_gnd tM2035(v(M12_v), N0563_v, N0563_port_1);
  spice_transistor_nmos_gnd tM1615(v(N0783_v), N0381_v, N0381_port_12);
  spice_transistor_nmos_gnd tM1614(v(N0783_v), N0406_v, N0406_port_12);
  spice_transistor_nmos_gnd tM1617(v(N0804_v), N0424_v, N0424_port_12);
  spice_transistor_nmos_gnd tM1616(v(N0804_v), N0410_v, N0410_port_12);
  spice_transistor_nmos_gnd tM1611(v(N0304_v), WADB2_v, WADB2_port_5);
  spice_transistor_nmos_gnd tM1610(v(N0318_v), WADB1_v, WADB1_port_5);
  spice_transistor_nmos_gnd tM1613(v(N0300_v), WADB2_v, WADB2_port_6);
  spice_transistor_nmos_gnd tM1612(v(N0300_v), WADB1_v, WADB1_port_6);
  spice_transistor_nmos tM2122(v(JCN_ISZ_v), N0373_v, N0372_v, N0373_port_0, N0372_port_0);
  spice_transistor_nmos tM2123(v(FIN_FIM_v), N0372_v, N0373_v, N0372_port_1, N0373_port_1);
  spice_transistor_nmos_gnd tM2120(v(_OPR_2_v), INC_ISZ_v, INC_ISZ_port_2);
  spice_transistor_nmos_gnd tM2121(v(_OPR_2_v), BBL_v, BBL_port_2);
  spice_transistor_nmos tM1619(v(N0382_v), N0381_v, ___SC__JIN_FIN__CLK1_M11_X21_INH__v, N0381_port_13, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_0);
  spice_transistor_nmos tM1618(v(N0382_v), N0406_v, __POC_CLK2_X12_X32__INH_v, N0406_port_13, __POC_CLK2_X12_X32__INH_port_0);
  spice_transistor_nmos_gnd tM2124(v(_OPR_2_v), JMS_v, JMS_port_2);
  spice_transistor_nmos_gnd tM2125(v(OPR_3_v), FIN_FIM_SRC_JIN_v, FIN_FIM_SRC_JIN_port_3);
  spice_transistor_nmos_gnd tM2830(v(N0727_v), A32_v, A32_port_9);
  spice_transistor_nmos_gnd tM2832(v(N0727_v), N0746_v, N0746_port_1);
  spice_transistor_nmos_vdd tM2834(v(S00778_v), N0746_v, N0746_port_2);
  spice_transistor_nmos_gnd tM2774(v(N0477_v), ADC_CY_v, ADC_CY_port_2);
  spice_transistor_nmos_gnd tM2838(v(N0348_v), N0819_v, N0819_port_1);
  spice_transistor_nmos_gnd tM2839(v(N0347_v), N0819_v, N0819_port_2);
  spice_transistor_nmos_gnd tM1079(v(N0295_v), N0738_v, N0738_port_3);
  spice_transistor_nmos_gnd tM1583(v(N0620_v), N0965_v, N0965_port_2);
  spice_transistor_nmos_gnd tM2237(v(OPA_0_v), N0516_v, N0516_port_0);
  spice_transistor_nmos_gnd tM2773(v(N0678_v), N0676_v, N0676_port_1);
  spice_transistor_nmos tM2934(v(clk2_v), N0285_v, A22_v, N0285_port_1, A22_port_6);
  spice_transistor_nmos_gnd tM3277(v(N0676_v), N0668_v, N0668_port_3);
  spice_transistor_nmos tM2238(v(FIM_SRC_v), N0516_v, _SRC_v, N0516_port_1, _SRC_port_0);
  spice_transistor_nmos_gnd tM2239(v(SC_v), N0417_v, N0417_port_0);
  spice_transistor_nmos tM1588(v(N0635_v), N0645_v, __POC__CLK2_SC_A32_X12__v, N0645_port_9, __POC__CLK2_SC_A32_X12__port_6);
  spice_transistor_nmos_gnd tM3154(v(N0345_v), N0359_v, N0359_port_1);
  spice_transistor_nmos_gnd tM3059(v(N0556_v), N0900_v, N0900_port_2);
  spice_transistor_nmos_gnd tM3058(v(N0872_v), N0900_v, N0900_port_1);
  spice_transistor_nmos tM3051(v(clk2_v), N0286_v, A12_v, N0286_port_1, A12_port_7);
  spice_transistor_nmos tM3050(v(clk1_v), N0729_v, N0728_v, N0729_port_2, N0728_port_1);
  spice_transistor_nmos_gnd tM3053(v(N0348_v), N0345_v, N0345_port_4);
  spice_transistor_nmos_gnd tM3052(v(N0768_v), DCL_2_v, DCL_2_port_1);
  spice_transistor_nmos_gnd tM3054(v(N0348_v), N0363_v, N0363_port_4);
  spice_transistor_nmos tM3057(v(N0559_v), N0900_v, N0879_v, N0900_port_0, N0879_port_4);
  spice_transistor_nmos tM1862(v(JCN_ISZ_v), N0338_v, N0326_v, N0338_port_0, N0326_port_5);
  spice_transistor_nmos tM1863(v(N0322_v), N0339_v, N0338_v, N0339_port_1, N0338_port_1);
  spice_transistor_nmos tM1860(v(N0310_v), N0341_v, N0339_v, N0341_port_0, N0339_port_0);
  spice_transistor_nmos tM1861(v(JUN_JMS_v), N0326_v, N0341_v, N0326_port_4, N0341_port_1);
  spice_transistor_nmos_gnd tM2139(v(OPR_2_v), N0636_v, N0636_port_2);
  spice_transistor_nmos_gnd tM1864(v(M22_v), N0339_v, N0339_port_2);
  spice_transistor_nmos_gnd tM1865(v(SC_v), N0310_v, N0310_port_3);
  spice_transistor_nmos_vdd tM1868(v(S00654_v), N0344_v, N0344_port_0);
  spice_transistor_nmos_gnd tM2138(v(OPR_2_v), XCH_v, XCH_port_1);
  spice_transistor_nmos_vdd tM1869(v(N0344_v), SC_v, SC_port_4);
  spice_transistor_nmos_gnd tM2693(v(N1006_v), N1007_v, N1007_port_3);
  spice_transistor_nmos_vdd tM2725(v(N0659_v), D1_v, D1_port_11);
  spice_transistor_nmos tM2723(v(SC_M22_CLK2_v), D3_v, N1012_v, D3_port_11, N1012_port_1);
  spice_transistor_nmos tM2457(v(clk1_v), N0719_v, N0718_v, N0719_port_2, N0718_port_1);
  spice_transistor_nmos_vdd tM2454(v(S00710_v), N0742_v, N0742_port_2);
  spice_transistor_nmos_gnd tM2455(v(N0281_v), N0718_v, N0718_port_0);
  spice_transistor_nmos tM1943(v(M22_v), N0484_v, N0485_v, N0484_port_0, N0485_port_1);
  spice_transistor_nmos_gnd tM2101(v(_OPR_3_v), LDM_BBL_v, LDM_BBL_port_0);
  spice_transistor_nmos_gnd tM1970(v(DC_v), RRAB0_v, RRAB0_port_5);
  spice_transistor_nmos_gnd tM1972(v(N0615_v), RRAB0_v, RRAB0_port_6);
  spice_transistor_nmos_gnd tM1973(v(N0460_v), CLK2_JMS_DC_M22_BBL_M22_X12_X22___v, CLK2_JMS_DC_M22_BBL_M22_X12_X22___port_4);
  spice_transistor_nmos tM1976(v(N0580_v), N0594_v, N0588_v, N0594_port_0, N0588_port_2);
  spice_transistor_nmos tM1977(v(FIN_FIM_SRC_JIN_v), N0588_v, N0589_v, N0588_port_3, N0589_port_1);
  spice_transistor_nmos_gnd tM1908(v(N0467_v), CLK2_JMS_DC_M22_BBL_M22_X12_X22___v, CLK2_JMS_DC_M22_BBL_M22_X12_X22___port_2);
  spice_transistor_nmos tM1378(v(RADB2_v), N0396_v, D0_v, N0396_port_0, D0_port_6);
  spice_transistor_nmos tM1376(v(WADB1_v), N0764_v, N0777_v, N0764_port_4, N0777_port_1);
  spice_transistor_nmos tM1377(v(RADB1_v), D0_v, N0395_v, D0_port_5, N0395_port_1);
  spice_transistor_nmos_gnd tM1374(v(N0777_v), N0395_v, N0395_port_0);
  spice_transistor_nmos_gnd tM1375(v(PC0_4_v), N0795_v, N0795_port_0);
  spice_transistor_nmos_gnd tM1372(v(PC1_0_v), N0815_v, N0815_port_0);
  spice_transistor_nmos tM1373(v(N0426_v), N0394_v, PC2_0_v, N0394_port_4, PC2_0_port_0);
  spice_transistor_nmos_gnd tM1370(v(PC0_0_v), N0794_v, N0794_port_1);
  spice_transistor_nmos tM1371(v(N0410_v), PC1_0_v, N0394_v, PC1_0_port_0, N0394_port_3);
  spice_transistor_nmos_gnd tM2131(v(OPR_2_v), FIN_FIM_v, FIN_FIM_port_2);
  spice_transistor_nmos tM1118(v(N0444_v), N0774_v, N0835_v, N0774_port_5, N0835_port_1);
  spice_transistor_nmos_vdd tM1119(v(__INH__X11_X31_CLK1_v), N0774_v, N0774_port_6);
  spice_transistor_nmos_gnd tM1112(v(N0497_v), N0862_v, N0862_port_1);
  spice_transistor_nmos_gnd tM1117(v(PC3_7_v), N0835_v, N0835_port_0);
  spice_transistor_nmos tM1115(v(N0424_v), N0778_v, N0808_v, N0778_port_3, N0808_port_1);
  spice_transistor_nmos tM1288(v(N0543_v), N0906_v, N0867_v, N0906_port_0, N0867_port_2);
  spice_transistor_nmos_gnd tM1289(v(R1_1_v), N0906_v, N0906_port_1);
  spice_transistor_nmos tM1282(v(N0634_v), N0532_v, R12_0_v, N0532_port_8, R12_0_port_0);
  spice_transistor_nmos_gnd tM1283(v(R6_1_v), N0949_v, N0949_port_0);
  spice_transistor_nmos tM1280(v(N0634_v), N0531_v, R13_0_v, N0531_port_8, R13_0_port_1);
  spice_transistor_nmos tM1281(v(N0647_v), R15_0_v, N0531_v, R15_0_port_1, N0531_port_9);
  spice_transistor_nmos tM1286(v(N0529_v), N0534_v, R1_1_v, N0534_port_2, R1_1_port_0);
  spice_transistor_nmos tM1287(v(N0544_v), R3_1_v, N0534_v, R3_1_port_0, N0534_port_3);
  spice_transistor_nmos tM1284(v(N0591_v), N0881_v, N0949_v, N0881_port_5, N0949_port_1);
  spice_transistor_nmos tM1285(v(N0544_v), R2_1_v, N0533_v, R2_1_port_1, N0533_port_3);
  spice_transistor_nmos tM2953(v(N0854_v), N0857_v, N0850_v, N0857_port_3, N0850_port_1);
  spice_transistor_nmos_gnd tM2952(v(N0850_v), N0347_v, N0347_port_4);
  spice_transistor_nmos tM2950(v(ADSR_v), N0848_v, ACC_1_v, N0848_port_0, ACC_1_port_4);
  spice_transistor_nmos tM2959(v(ACC_ADA_v), N0871_v, N0857_v, N0871_port_6, N0857_port_4);
  spice_transistor_nmos_gnd tM2958(v(N0889_v), N0899_v, N0899_port_3);
  spice_transistor_nmos_gnd tM1579(v(N0455_v), N0463_v, N0463_port_3);
  spice_transistor_nmos_gnd tM1261(v(R2_1_v), N0922_v, N0922_port_0);
  spice_transistor_nmos_vdd tM1575(v(S00557_v), RRAB1_v, RRAB1_port_4);
  spice_transistor_nmos_vdd tM1577(v(__INH__X11_X31_CLK1_v), N0773_v, N0773_port_6);
  spice_transistor_nmos tM1570(v(N0599_v), CLK2_SC_A12_M12__v, N0598_v, CLK2_SC_A12_M12__port_4, N0598_port_9);
  spice_transistor_nmos tM1571(v(N0620_v), N0619_v, CLK2_SC_A12_M12__v, N0619_port_9, CLK2_SC_A12_M12__port_5);
  spice_transistor_nmos_gnd tM1573(v(N0599_v), N0955_v, N0955_port_2);
  spice_transistor_nmos_vdd tM1754(v(S00599_v), N0411_v, N0411_port_5);
  spice_transistor_nmos_vdd tM1755(v(S00600_v), N0427_v, N0427_port_5);
  spice_transistor_nmos_gnd tM1756(v(N0420_v), N0401_v, N0401_port_2);
  spice_transistor_nmos_gnd tM1023(v(N0740_v), sync_v, sync_port_0);
  spice_transistor_nmos tM1020(v(N0290_v), N0311_v, N0312_v, N0311_port_1, N0312_port_0);
  spice_transistor_nmos tM1021(v(N0290_v), N0301_v, N0302_v, N0301_port_3, N0302_port_0);
  spice_transistor_nmos_gnd tM2005(v(N0627_v), __POC__CLK2_SC_A32_X12__v, __POC__CLK2_SC_A32_X12__port_8);
  spice_transistor_nmos_gnd tM2007(v(N0547_v), WRAB0_v, WRAB0_port_5);
  spice_transistor_nmos tM1758(v(N0466_v), N0491_v, N0475_v, N0491_port_1, N0475_port_4);
  spice_transistor_nmos_gnd tM1759(v(N0458_v), N0465_v, N0465_port_0);
  spice_transistor_nmos_vdd tM1028(v(S00536_v), N0738_v, N0738_port_0);
  spice_transistor_nmos tM1265(v(N0632_v), N0866_v, N0966_v, N0866_port_7, N0966_port_1);
  spice_transistor_nmos_gnd tM1594(v(N0635_v), N0974_v, N0974_port_2);
  spice_transistor_nmos_gnd tM1595(v(N0648_v), N0983_v, N0983_port_2);
  spice_transistor_nmos tM1266(v(N0645_v), N0975_v, N0866_v, N0975_port_0, N0866_port_8);
  spice_transistor_nmos tM1591(v(N0648_v), N0657_v, __POC__CLK2_SC_A32_X12__v, N0657_port_9, __POC__CLK2_SC_A32_X12__port_7);
  spice_transistor_nmos_gnd tM1267(v(R13_0_v), N0975_v, N0975_port_1);
  spice_transistor_nmos_gnd tM2481(v(OPA_0_v), N0512_v, N0512_port_1);
  spice_transistor_nmos tM2480(v(N0432_v), N0512_v, N0486_v, N0512_port_0, N0486_port_5);
  spice_transistor_nmos_gnd tM2483(v(_OPA_0_v), TCS_v, TCS_port_5);
  spice_transistor_nmos_gnd tM2482(v(_OPA_0_v), DCL_v, DCL_port_5);
  spice_transistor_nmos_gnd tM2485(v(_OPA_0_v), RAL_v, RAL_port_5);
  spice_transistor_nmos_gnd tM2484(v(_OPA_0_v), DAA_v, DAA_port_5);
  spice_transistor_nmos_gnd tM2487(v(_OPA_0_v), CMC_v, CMC_port_5);
  spice_transistor_nmos_gnd tM2486(v(_OPA_0_v), TCC_v, TCC_port_5);
  spice_transistor_nmos_gnd tM2489(v(_OPA_0_v), ADM_v, ADM_port_5);
  spice_transistor_nmos_gnd tM2488(v(_OPA_0_v), CLC_v, CLC_port_5);
  spice_transistor_nmos_gnd tM2710(v(LDM_BBL_v), N0658_v, N0658_port_1);
  spice_transistor_nmos tM2715(v(SC_M22_CLK2_v), D2_v, N1013_v, D2_port_11, N1013_port_1);
  spice_transistor_nmos_gnd tM2717(v(N0658_v), OPA_IB_v, OPA_IB_port_4);
  spice_transistor_nmos_gnd tM2716(v(N0689_v), d3_v, d3_port_0);
  spice_transistor_nmos_gnd tM2719(v(__X21__CLK2__v), OPA_IB_v, OPA_IB_port_5);
  spice_transistor_nmos tM1620(v(N0411_v), N0410_v, ___SC__JIN_FIN__CLK1_M11_X21_INH__v, N0410_port_13, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_1);
  spice_transistor_nmos tM1621(v(N0411_v), N0424_v, __POC_CLK2_X12_X32__INH_v, N0424_port_13, __POC_CLK2_X12_X32__INH_port_1);
  spice_transistor_nmos tM1623(v(N0732_v), N0711_v, N0712_v, N0711_port_2, N0712_port_2);
  spice_transistor_nmos_gnd tM1624(v(N0820_v), N0434_v, N0434_port_12);
  spice_transistor_nmos_gnd tM1625(v(N0820_v), N0426_v, N0426_port_12);
  spice_transistor_nmos_gnd tM1626(v(N0833_v), N0439_v, N0439_port_12);
  spice_transistor_nmos_gnd tM1627(v(N0833_v), N0444_v, N0444_port_12);
  spice_transistor_nmos tM1628(v(clk1_v), ADDR_RFSH_0_v, N0519_v, ADDR_RFSH_0_port_2, N0519_port_0);
  spice_transistor_nmos_gnd tM1629(v(N0540_v), N0545_v, N0545_port_3);
  spice_transistor_nmos_gnd tM2133(v(OPR_2_v), FIM_SRC_v, FIM_SRC_port_1);
  spice_transistor_nmos_gnd tM2132(v(OPR_2_v), JCN_v, JCN_port_1);
  spice_transistor_nmos_gnd tM2135(v(OPR_2_v), JIN_FIN_v, JIN_FIN_port_5);
  spice_transistor_nmos_gnd tM2134(v(_OPR_2_v), JUN2_JMS2_v, JUN2_JMS2_port_1);
  spice_transistor_nmos_gnd tM2137(v(_OPR_1_v), ISZ_v, ISZ_port_2);
  spice_transistor_nmos_gnd tM2136(v(_OPR_1_v), FIN_FIM_v, FIN_FIM_port_3);
  spice_transistor_nmos_vdd tM2829(v(N0746_v), A32_v, A32_port_8);
  spice_transistor_nmos tM2828(v(N0356_v), N0803_v, N0819_v, N0803_port_3, N0819_port_0);
  spice_transistor_nmos_gnd tM2826(v(KBP_v), N0350_v, N0350_port_1);
  spice_transistor_nmos_gnd tM2825(v(O_IB_v), N0378_v, N0378_port_1);
  spice_transistor_nmos tM2824(v(DAA_v), N0378_v, N0818_v, N0378_port_0, N0818_port_1);
  spice_transistor_nmos_gnd tM2823(v(N0803_v), N0818_v, N0818_port_0);
  spice_transistor_nmos_gnd tM2821(v(A32_v), N0288_v, N0288_port_4);
  spice_transistor_nmos tM3198(v(N0861_v), N0901_v, N0877_v, N0901_port_1, N0877_port_3);
  spice_transistor_nmos tM3191(v(ADSL_v), N0514_v, N0513_v, N0514_port_6, N0513_port_2);
  spice_transistor_nmos tM3192(v(N0854_v), N0859_v, N0852_v, N0859_port_3, N0852_port_1);
  spice_transistor_nmos tM3193(v(ADSR_v), N0513_v, ACC_3_v, N0513_port_3, ACC_3_port_4);
  spice_transistor_nmos tM3194(v(N0893_v), N0914_v, N0557_v, N0914_port_0, N0557_port_1);
  spice_transistor_nmos_gnd tM3195(v(N0873_v), N0901_v, N0901_port_0);
  spice_transistor_nmos_gnd tM2224(v(OPR_0_v), ADD_v, ADD_port_3);
  spice_transistor_nmos_gnd tM2221(v(OPR_0_v), BBL_v, BBL_port_4);
  spice_transistor_nmos_gnd tM2223(v(OPR_0_v), LD_v, LD_port_3);
  spice_transistor_nmos_vdd tM2222(v(N0999_v), OPR_0_v, OPR_0_port_3);
  spice_transistor_nmos_gnd tM2851(v(ACC_0_v), N0856_v, N0856_port_3);
  spice_transistor_nmos_gnd tM2856(v(N0846_v), ADD_0_v, ADD_0_port_1);
  spice_transistor_nmos_gnd tM3288(v(POC_v), d0_v, d0_port_4);
  spice_transistor_nmos tM2854(v(ACB_IB_v), N0346_v, D0_v, N0346_port_3, D0_port_12);
  spice_transistor_nmos_gnd tM3284(v(N0664_v), D3_v, D3_port_17);
  spice_transistor_nmos_vdd tM3285(v(N0663_v), D3_v, D3_port_18);
  spice_transistor_nmos_gnd tM3286(v(POC_v), d3_v, d3_port_2);
  spice_transistor_nmos_vdd tM3287(v(N0693_v), d1_v, d1_port_2);
  spice_transistor_nmos_gnd tM3281(v(D1_v), N0673_v, N0673_port_0);
  spice_transistor_nmos tM3282(v(N0702_v), N0673_v, N0694_v, N0673_port_1, N0694_port_0);
  spice_transistor_nmos tM3064(v(N0964_v), D2_v, N0606_v, D2_port_15, N0606_port_0);
  spice_transistor_nmos_gnd tM3060(v(N0891_v), N0900_v, N0900_port_3);
  spice_transistor_nmos tM3062(v(N0556_v), N0554_v, N0555_v, N0554_port_2, N0555_port_2);
  spice_transistor_nmos_gnd tM3063(v(N0691_v), N0690_v, N0690_port_2);
  spice_transistor_nmos_gnd tM3068(v(N0944_v), _TMP_2_v, _TMP_2_port_0);
  spice_transistor_nmos tM3069(v(N0937_v), _TMP_2_v, N0891_v, _TMP_2_port_1, N0891_port_4);
  spice_transistor_nmos_gnd tM3266(v(N0696_v), N0698_v, N0698_port_1);
  spice_transistor_nmos_gnd tM3267(v(N0700_v), N0698_v, N0698_port_2);
  spice_transistor_nmos_gnd tM3262(v(N0700_v), N0696_v, N0696_port_2);
  spice_transistor_nmos_gnd tM3260(v(N0736_v), cm_ram0_v, cm_ram0_port_1);
  spice_transistor_nmos_gnd tM3261(v(N0698_v), d0_v, d0_port_3);
  spice_transistor_nmos_gnd tM1105(v(PC1_3_v), N0808_v, N0808_port_0);
  spice_transistor_nmos_gnd tM2924(v(N0857_v), N0472_v, N0472_port_3);
  spice_transistor_nmos_gnd tM1314(v(R12_1_v), N0977_v, N0977_port_1);
  spice_transistor_nmos_gnd tM2359(v(OPA_3_v), N0481_v, N0481_port_3);
  spice_transistor_nmos_vdd tM2799(v(N0704_v), N0700_v, N0700_port_2);
  spice_transistor_nmos_gnd tM1311(v(R5_1_v), N0932_v, N0932_port_1);
  spice_transistor_nmos_gnd tM2751(v(N0855_v), N0470_v, N0470_port_3);
  spice_transistor_nmos_gnd tM2664(v(SUB_v), READ_ACC_3__v, READ_ACC_3__port_8);
  spice_transistor_nmos_gnd tM2129(v(_OPR_2_v), LDM_BBL_v, LDM_BBL_port_1);
  spice_transistor_nmos_gnd tM1965(v(N0637_v), N0642_v, N0642_port_3);
  spice_transistor_nmos_gnd tM1964(v(N0637_v), N0641_v, N0641_port_2);
  spice_transistor_nmos tM1369(v(N0406_v), N0794_v, N0781_v, N0794_port_0, N0781_port_2);
  spice_transistor_nmos tM1368(v(N0381_v), N0394_v, PC0_0_v, N0394_port_2, PC0_0_port_0);
  spice_transistor_nmos tM1365(v(N0444_v), N0780_v, N0842_v, N0780_port_5, N0842_port_1);
  spice_transistor_nmos tM1364(v(N0410_v), PC1_1_v, N0393_v, PC1_1_port_1, N0393_port_3);
  spice_transistor_nmos tM1367(v(N0439_v), PC3_1_v, N0393_v, PC3_1_port_1, N0393_port_5);
  spice_transistor_nmos tM1366(v(N0426_v), N0393_v, PC2_1_v, N0393_port_4, PC2_1_port_1);
  spice_transistor_nmos tM1361(v(RRAB1_v), D3_v, N0538_v, D3_port_5, N0538_port_0);
  spice_transistor_nmos tM1360(v(M12_M22_CLK1__M11_M12__v), N0500_v, D3_v, N0500_port_1, D3_port_4);
  spice_transistor_nmos_gnd tM1363(v(PC3_1_v), N0842_v, N0842_port_0);
  spice_transistor_nmos tM1362(v(RRAB0_v), N0537_v, D3_v, N0537_port_0, D3_port_6);
  spice_transistor_nmos tM1109(v(WRAB1_v), N0862_v, N0866_v, N0862_port_0, N0866_port_0);
  spice_transistor_nmos tM1108(v(M12_M22_CLK1__M11_M12__v), D0_v, N0497_v, D0_port_2, N0497_port_0);
  spice_transistor_nmos tM1101(v(N0434_v), N0822_v, N0774_v, N0822_port_0, N0774_port_4);
  spice_transistor_nmos tM1100(v(N0424_v), N0774_v, N0807_v, N0774_port_3, N0807_port_1);
  spice_transistor_nmos_gnd tM1103(v(N0779_v), N0388_v, N0388_port_1);
  spice_transistor_nmos_gnd tM1102(v(PC2_7_v), N0822_v, N0822_port_1);
  spice_transistor_nmos_vdd tM1107(v(__INH__X11_X31_CLK1_v), N0770_v, N0770_port_6);
  spice_transistor_nmos tM1106(v(N0439_v), PC3_7_v, N0386_v, PC3_7_port_0, N0386_port_5);
  spice_transistor_nmos tM1299(v(N0632_v), N0881_v, N0968_v, N0881_port_7, N0968_port_1);
  spice_transistor_nmos_gnd tM1298(v(R10_1_v), N0968_v, N0968_port_0);
  spice_transistor_nmos tM1291(v(N0616_v), N0958_v, N0881_v, N0958_port_0, N0881_port_6);
  spice_transistor_nmos tM1290(v(N0569_v), N0533_v, R4_1_v, N0533_port_4, R4_1_port_1);
  spice_transistor_nmos_gnd tM1293(v(R10_0_v), N0967_v, N0967_port_0);
  spice_transistor_nmos_gnd tM1292(v(R8_1_v), N0958_v, N0958_port_1);
  spice_transistor_nmos tM1295(v(N0645_v), N0976_v, N0880_v, N0976_port_0, N0880_port_8);
  spice_transistor_nmos tM1294(v(N0632_v), N0880_v, N0967_v, N0880_port_7, N0967_port_1);
  spice_transistor_nmos tM1297(v(N0647_v), R14_0_v, N0532_v, R14_0_port_0, N0532_port_9);
  spice_transistor_nmos_gnd tM1296(v(R12_0_v), N0976_v, N0976_port_1);
  spice_transistor_nmos tM2923(v(M12_v), N0472_v, ACC_1_v, N0472_port_2, ACC_1_port_0);
  spice_transistor_nmos tM2920(v(N0889_v), N0875_v, N0888_v, N0875_port_1, N0888_port_1);
  spice_transistor_nmos_gnd tM2921(v(N0347_v), ACC_0_v, ACC_0_port_8);
  spice_transistor_nmos tM2927(v(N0553_v), N0551_v, N0552_v, N0551_port_0, N0552_port_0);
  spice_transistor_nmos tM2925(v(ADSL_v), N0846_v, ACC_1_v, N0846_port_6, ACC_1_port_1);
  spice_transistor_nmos_gnd tM2928(v(N0871_v), N0551_v, N0551_port_1);
  spice_transistor_nmos_gnd tM2929(v(N0889_v), N0552_v, N0552_port_1);
  spice_transistor_nmos tM1569(v(N0599_v), N0616_v, __POC__CLK2_SC_A32_X12__v, N0616_port_9, __POC__CLK2_SC_A32_X12__port_4);
  spice_transistor_nmos_gnd tM1568(v(N0965_v), N0632_v, N0632_port_8);
  spice_transistor_nmos_gnd tM1563(v(N0545_v), N0919_v, N0919_port_2);
  spice_transistor_nmos tM1560(v(N0584_v), N0583_v, CLK2_SC_A12_M12__v, N0583_port_9, CLK2_SC_A12_M12__port_3);
  spice_transistor_nmos_gnd tM1567(v(N0965_v), N0619_v, N0619_port_8);
  spice_transistor_nmos_gnd tM1566(v(N0955_v), N0598_v, N0598_port_8);
  spice_transistor_nmos_gnd tM1565(v(N0584_v), N0938_v, N0938_port_2);
  spice_transistor_nmos_gnd tM1564(v(N0570_v), N0928_v, N0928_port_2);
  spice_transistor_nmos_gnd tM1743(v(N0401_v), N0411_v, N0411_port_4);
  spice_transistor_nmos_gnd tM1034(v(N0290_v), N0756_v, N0756_port_0);
  spice_transistor_nmos_gnd tM1741(v(N0409_v), N0411_v, N0411_port_3);
  spice_transistor_nmos_gnd tM1740(v(N0400_v), N0382_v, N0382_port_3);
  spice_transistor_nmos tM1031(v(RADB0_v), N0388_v, D2_v, N0388_port_0, D2_port_1);
  spice_transistor_nmos_vdd tM1030(v(N0738_v), sync_v, sync_port_1);
  spice_transistor_nmos tM1033(v(N0298_v), N0762_v, N0755_v, N0762_port_0, N0755_port_1);
  spice_transistor_nmos_gnd tM1744(v(N0420_v), N0427_v, N0427_port_4);
  spice_transistor_nmos_gnd tM2031(v(N0603_v), N0568_v, N0568_port_0);
  spice_transistor_nmos_vdd tM1749(v(S00598_v), N0382_v, N0382_port_5);
  spice_transistor_nmos_gnd tM1039(v(N0758_v), N0763_v, N0763_port_0);
  spice_transistor_nmos_gnd tM1038(v(N0756_v), N0762_v, N0762_port_2);
  spice_transistor_nmos_gnd tM2036(v(M22_v), N0576_v, N0576_port_0);
  spice_transistor_nmos tM2037(v(N0564_v), N0575_v, N0576_v, N0575_port_0, N0576_port_1);
  spice_transistor_nmos_gnd tM1585(v(N0974_v), N0634_v, N0634_port_8);
  spice_transistor_nmos_gnd tM1584(v(N0974_v), N0645_v, N0645_port_8);
  spice_transistor_nmos_gnd tM1587(v(N0983_v), N0657_v, N0657_port_8);
  spice_transistor_nmos_gnd tM1586(v(N0983_v), N0647_v, N0647_port_8);
  spice_transistor_nmos_gnd tM1580(v(N0463_v), N0455_v, N0455_port_3);
  spice_transistor_nmos tM1589(v(N0635_v), N0634_v, CLK2_SC_A12_M12__v, N0634_port_9, CLK2_SC_A12_M12__port_6);
  spice_transistor_nmos_gnd tM1930(v(SC_v), N0435_v, N0435_port_1);
  spice_transistor_nmos_vdd tM2724(v(S00716_v), OPA_IB_v, OPA_IB_port_6);
  spice_transistor_nmos_vdd tM2726(v(N0659_v), D3_v, D3_port_12);
  spice_transistor_nmos_gnd tM1933(v(A32_v), N0428_v, N0428_port_3);
  spice_transistor_nmos tM2720(v(SC_M22_CLK2_v), D1_v, N1014_v, D1_port_10, N1014_port_1);
  spice_transistor_nmos_vdd tM2721(v(N0687_v), d3_v, d3_port_1);
  spice_transistor_nmos_gnd tM1544(v(PC3_8_v), N0845_v, N0845_port_0);
  spice_transistor_nmos_gnd tM2104(v(IOR_v), N0683_v, N0683_port_2);
  spice_transistor_nmos_gnd tM2105(v(A32_v), N0682_v, N0682_port_2);
  spice_transistor_nmos_gnd tM2106(v(M12_v), N0682_v, N0682_port_3);
  spice_transistor_nmos_gnd tM2107(v(N0703_v), L_v, L_port_0);
  spice_transistor_nmos_gnd tM2100(v(OPR_3_v), N0636_v, N0636_port_1);
  spice_transistor_nmos tM1547(v(N0463_v), N0488_v, N0469_v, N0488_port_0, N0469_port_4);
  spice_transistor_nmos_gnd tM2102(v(A32_v), N0629_v, N0629_port_1);
  spice_transistor_nmos tM2103(v(SC_v), N0629_v, N0631_v, N0629_port_2, N0631_port_0);
  spice_transistor_nmos tM2753(v(CY_IB_v), D0_v, CY_1_v, D0_port_11, CY_1_port_2);
  spice_transistor_nmos_vdd tM1546(v(__INH__X11_X31_CLK1_v), N0777_v, N0777_port_6);
  spice_transistor_nmos_gnd tM2108(v(N0703_v), L_v, L_port_1);
  spice_transistor_nmos tM2109(v(clk2_v), N0631_v, N0630_v, N0631_port_1, N0630_port_1);
  spice_transistor_nmos_gnd tM2459(v(X22_v), N0383_v, N0383_port_0);
  spice_transistor_nmos_gnd tM3231(v(vss_v), d0_v, d0_port_0);
  spice_transistor_nmos_gnd tM1639(v(N0541_v), N0545_v, N0545_port_4);
  spice_transistor_nmos_gnd tM1638(v(N0541_v), N0539_v, N0539_port_1);
  spice_transistor_nmos_gnd tM1637(v(N0646_v), N0613_v, N0613_port_6);
  spice_transistor_nmos_gnd tM1636(v(N0613_v), N0648_v, N0648_port_3);
  spice_transistor_nmos_gnd tM1635(v(N0613_v), N0635_v, N0635_port_3);
  spice_transistor_nmos_gnd tM1634(v(N0613_v), N0620_v, N0620_port_3);
  spice_transistor_nmos_gnd tM1633(v(N0613_v), N0540_v, N0540_port_5);
  spice_transistor_nmos_gnd tM1632(v(N0613_v), N0599_v, N0599_port_3);
  spice_transistor_nmos_gnd tM1631(v(N0540_v), N0584_v, N0584_port_3);
  spice_transistor_nmos_gnd tM1630(v(N0540_v), N0570_v, N0570_port_3);
  spice_transistor_nmos_gnd tM2943(v(N0342_v), N0964_v, N0964_port_1);
  spice_transistor_nmos_gnd tM3178(v(N0859_v), N0474_v, N0474_port_3);
  spice_transistor_nmos_gnd tM2588(v(XCH_v), WRITE_ACC_1__v, WRITE_ACC_1__port_3);
  spice_transistor_nmos_gnd tM2589(v(POC_v), WRITE_ACC_1__v, WRITE_ACC_1__port_4);
  spice_transistor_nmos tM2858(v(ADD_ACC_v), N0846_v, ACC_0_v, N0846_port_4, ACC_0_port_6);
  spice_transistor_nmos_gnd tM2859(v(N0878_v), N0874_v, N0874_port_1);
  spice_transistor_nmos_gnd tM2946(v(ACC_1_v), N0857_v, N0857_port_1);
  spice_transistor_nmos_gnd tM2580(v(N0803_v), N0403_v, N0403_port_0);
  spice_transistor_nmos_gnd tM2581(v(N0725_v), M12_v, M12_port_11);
  spice_transistor_nmos tM2850(v(ADSL_v), CY_1_v, ACC_0_v, CY_1_port_6, ACC_0_port_2);
  spice_transistor_nmos_gnd tM2583(v(POC_v), N0717_v, N0717_port_2);
  spice_transistor_nmos_vdd tM2584(v(S00757_v), N0717_v, N0717_port_3);
  spice_transistor_nmos tM2857(v(M12_v), ACC_0_v, N0471_v, ACC_0_port_5, N0471_port_1);
  spice_transistor_nmos_gnd tM2586(v(N0802_v), N0403_v, N0403_port_1);
  spice_transistor_nmos_gnd tM2587(v(__X21__CLK2__v), N0448_v, N0448_port_1);
  spice_transistor_nmos_vdd tM3272(v(S00819_v), N0937_v, N0937_port_6);
  spice_transistor_nmos_gnd tM2210(v(_OPR_0_v), N0636_v, N0636_port_4);
  spice_transistor_nmos_gnd tM2211(v(_OPR_0_v), SUB_v, SUB_port_3);
  spice_transistor_nmos_vdd tM2212(v(N0998_v), _OPR_0_v, _OPR_0_port_10);
  spice_transistor_nmos_gnd tM2213(v(OPA_0_v), FIN_FIM_v, FIN_FIM_port_4);
  spice_transistor_nmos_gnd tM2214(v(OPR_0_v), FIM_SRC_v, FIM_SRC_port_3);
  spice_transistor_nmos_gnd tM2215(v(OPR_0_v), IO_v, IO_port_3);
  spice_transistor_nmos_gnd tM3173(v(N0363_v), N0357_v, N0357_port_2);
  spice_transistor_nmos_gnd tM2219(v(A12_v), N0769_v, N0769_port_1);
  spice_transistor_nmos_gnd tM2401(v(OPA_2_v), DAA_v, DAA_port_3);
  spice_transistor_nmos_gnd tM3299(v(N0700_v), N0695_v, N0695_port_2);
  spice_transistor_nmos_gnd tM3298(v(N0693_v), N0695_v, N0695_port_1);
  spice_transistor_nmos_gnd tM3174(v(N0377_v), N0357_v, N0357_port_3);
  spice_transistor_nmos_gnd tM3293(v(N0695_v), d1_v, d1_port_3);
  spice_transistor_nmos_vdd tM3292(v(S00836_v), N0693_v, N0693_port_3);
  spice_transistor_nmos tM3175(v(N0415_v), D1_v, N0359_v, D1_port_15, N0359_port_5);
  spice_transistor_nmos_gnd tM3297(v(N0676_v), N0664_v, N0664_port_2);
  spice_transistor_nmos_gnd tM3073(v(N0676_v), N0665_v, N0665_port_0);
  spice_transistor_nmos_vdd tM3072(v(M12_v), N0606_v, N0606_port_1);
  spice_transistor_nmos_gnd tM3071(v(N0692_v), d2_v, d2_port_1);
  spice_transistor_nmos_vdd tM3070(v(N0943_v), _TMP_2_v, _TMP_2_port_2);
  spice_transistor_nmos_vdd tM3077(v(N0913_v), N0559_v, N0559_port_2);
  spice_transistor_nmos_gnd tM3076(v(N0917_v), N0559_v, N0559_port_1);
  spice_transistor_nmos_gnd tM3074(v(N0913_v), N0917_v, N0917_port_0);
  spice_transistor_nmos_gnd tM2013(v(SC_v), DC_v, DC_port_5);
  spice_transistor_nmos_gnd tM3275(v(N0668_v), N0667_v, N0667_port_0);
  spice_transistor_nmos_gnd tM3274(v(N0668_v), D1_v, D1_port_16);
  spice_transistor_nmos_gnd tM3276(v(N0676_v), N0667_v, N0667_port_1);
  spice_transistor_nmos_gnd tM3271(v(d1_v), N0668_v, N0668_port_0);
  spice_transistor_nmos_gnd tM2407(v(OPA_2_v), CMC_v, CMC_port_3);
  spice_transistor_nmos_gnd tM3273(v(vss_v), d2_v, d2_port_4);
  spice_transistor_nmos_vdd tM2870(v(N0939_v), _TMP_0_v, _TMP_0_port_2);
  spice_transistor_nmos_vdd tM3279(v(N0667_v), D1_v, D1_port_17);
  spice_transistor_nmos tM1440(v(N0543_v), N0910_v, N0869_v, N0910_port_0, N0869_port_2);
  spice_transistor_nmos_gnd tM1441(v(R1_3_v), N0910_v, N0910_port_1);
  spice_transistor_nmos_gnd tM3187(v(N0893_v), N0558_v, N0558_port_0);
  spice_transistor_nmos_gnd tM3186(v(N0873_v), N0557_v, N0557_port_0);
  spice_transistor_nmos tM3179(v(ADSL_v), N0848_v, ACC_3_v, N0848_port_6, ACC_3_port_1);
  spice_transistor_nmos tM3184(v(N0559_v), N0892_v, N0897_v, N0892_port_0, N0897_port_1);
  spice_transistor_nmos_gnd tM3183(v(N0877_v), N0885_v, N0885_port_1);
  spice_transistor_nmos_gnd tM3182(v(N0873_v), N0897_v, N0897_port_0);
  spice_transistor_nmos tM3189(v(ADD_ACC_v), N0514_v, ACC_3_v, N0514_port_5, ACC_3_port_3);
  spice_transistor_nmos_gnd tM3188(v(ACC_3_v), N0859_v, N0859_port_1);
  spice_transistor_nmos_gnd tM2792(v(N0452_v), CY_1_v, CY_1_port_3);
  spice_transistor_nmos tM3185(v(N0893_v), N0877_v, N0892_v, N0877_port_2, N0892_port_1);
  spice_transistor_nmos_gnd tM2971(v(POC_v), d2_v, d2_port_0);
  spice_transistor_nmos_gnd tM2403(v(N1002_v), OPA_2_v, OPA_2_port_4);
  spice_transistor_nmos_gnd tM2796(v(SUB_GROUP_6__v), N0937_v, N0937_port_0);
  spice_transistor_nmos_gnd tM3181(v(N0606_v), N0943_v, N0943_port_4);
  spice_transistor_nmos_gnd tM2491(v(OPA_0_v), RAR_v, RAR_port_5);
  spice_transistor_nmos_gnd tM2497(v(OPA_0_v), IAC_v, IAC_port_5);
  spice_transistor_nmos tM2884(v(SUB_GROUP_6__v), TMP_0_v, N0887_v, TMP_0_port_0, N0887_port_5);
  spice_transistor_nmos_gnd tM2499(v(OPA_0_v), SBM_v, SBM_port_5);
  spice_transistor_nmos tM2881(v(ACC_ADA_v), N0870_v, N0471_v, N0870_port_6, N0471_port_3);
  spice_transistor_nmos_gnd tM1912(v(N0600_v), N0609_v, N0609_port_2);
  spice_transistor_nmos tM1913(v(N0574_v), N0600_v, N0601_v, N0600_port_2, N0601_port_0);
  spice_transistor_nmos tM1910(v(SC_A12_CLK2_v), N0574_v, N0585_v, N0574_port_4, N0585_port_0);
  spice_transistor_nmos tM1911(v(N0571_v), N0625_v, N0609_v, N0625_port_0, N0609_port_1);
  spice_transistor_nmos_gnd tM1916(v(N0586_v), N0585_v, N0585_port_1);
  spice_transistor_nmos_gnd tM1917(v(N0593_v), N0601_v, N0601_port_1);
  spice_transistor_nmos_gnd tM1914(v(N0610_v), REG_RFSH_1_v, REG_RFSH_1_port_3);
  spice_transistor_nmos_gnd tM1915(v(N0610_v), N0600_v, N0600_port_3);
  spice_transistor_nmos_gnd tM1918(v(clk2_v), RRAB1_v, RRAB1_port_7);
  spice_transistor_nmos_gnd tM2069(v(POC_v), N0626_v, N0626_port_4);
  spice_transistor_nmos_gnd tM2068(v(N0630_v), N0626_v, N0626_port_3);
  spice_transistor_nmos_gnd tM2789(v(N0705_v), N0704_v, N0704_port_0);
  spice_transistor_nmos_gnd tM2706(v(N0687_v), N0689_v, N0689_port_2);
  spice_transistor_nmos_vdd tM1359(v(__INH__X11_X31_CLK1_v), N0776_v, N0776_port_6);
  spice_transistor_nmos_gnd tM1350(v(R9_2_v), N0960_v, N0960_port_1);
  spice_transistor_nmos tM1351(v(N0647_v), R15_1_v, N0534_v, R15_1_port_0, N0534_port_9);
  spice_transistor_nmos_gnd tM1352(v(R15_1_v), N0987_v, N0987_port_0);
  spice_transistor_nmos_gnd tM1353(v(R11_2_v), N0970_v, N0970_port_0);
  spice_transistor_nmos tM1354(v(N0569_v), N0535_v, R5_2_v, N0535_port_4, R5_2_port_1);
  spice_transistor_nmos tM1355(v(N0583_v), R7_2_v, N0535_v, R7_2_port_1, N0535_port_5);
  spice_transistor_nmos tM1356(v(N0569_v), N0536_v, R4_2_v, N0536_port_4, R4_2_port_0);
  spice_transistor_nmos_gnd tM1357(v(R0_3_v), N0909_v, N0909_port_0);
  spice_transistor_nmos_gnd tM2406(v(OPA_2_v), STC_v, STC_port_3);
  spice_transistor_nmos tM2869(v(N0937_v), _TMP_0_v, N0887_v, _TMP_0_port_1, N0887_port_3);
  spice_transistor_nmos_gnd tM1828(v(N0449_v), N0450_v, N0450_port_2);
  spice_transistor_nmos tM1826(v(JCN_ISZ_v), N0321_v, N0323_v, N0321_port_0, N0323_port_2);
  spice_transistor_nmos tM1827(v(N0322_v), N0318_v, N0321_v, N0318_port_4, N0321_port_1);
  spice_transistor_nmos tM1824(v(X22_v), N0318_v, N0319_v, N0318_port_2, N0319_port_1);
  spice_transistor_nmos tM1825(v(N0310_v), N0324_v, N0318_v, N0324_port_1, N0318_port_3);
  spice_transistor_nmos_gnd tM1822(v(SC_v), N0320_v, N0320_port_0);
  spice_transistor_nmos tM1823(v(JIN_FIN_v), N0319_v, N0320_v, N0319_port_0, N0320_port_1);
  spice_transistor_nmos_gnd tM1820(v(A32_v), N0304_v, N0304_port_3);
  spice_transistor_nmos tM1821(v(JUN_JMS_v), N0323_v, N0324_v, N0323_port_1, N0324_port_0);
  spice_transistor_nmos tM2534(v(N0328_v), N0332_v, N0336_v, N0332_port_0, N0336_port_1);
  spice_transistor_nmos tM1804(v(X32_v), ADDR_PTR_0_v, N0420_v, ADDR_PTR_0_port_0, N0420_port_4);
  spice_transistor_nmos tM3228(v(N0964_v), D3_v, N0607_v, D3_port_16, N0607_port_1);
  spice_transistor_nmos tM2537(v(POC_v), N0332_v, N0331_v, N0332_port_2, N0331_port_2);
  spice_transistor_nmos_gnd tM2536(v(clk2_v), N0423_v, N0423_port_0);
  spice_transistor_nmos tM2531(v(clk2_v), N0360_v, N0369_v, N0360_port_1, N0369_port_2);
  spice_transistor_nmos_gnd tM2530(v(X12_v), N0369_v, N0369_port_1);
  spice_transistor_nmos_gnd tM2933(v(N0285_v), N0726_v, N0726_port_0);
  spice_transistor_nmos tM2935(v(clk1_v), N0727_v, N0726_v, N0727_port_2, N0726_port_1);
  spice_transistor_nmos tM2533(v(N0337_v), N0336_v, N0335_v, N0336_port_0, N0335_port_1);
  spice_transistor_nmos_gnd tM2937(v(DCL_1_v), N0716_v, N0716_port_1);
  spice_transistor_nmos tM2939(v(N0889_v), N0912_v, N0551_v, N0912_port_0, N0551_port_2);
  spice_transistor_nmos tM2938(v(N0351_v), N0371_v, N0767_v, N0371_port_3, N0767_port_2);
  spice_transistor_nmos_gnd tM2532(v(clk1_v), N0335_v, N0335_port_0);
  spice_transistor_nmos_gnd tM1000(v(N0770_v), N0385_v, N0385_port_0);
  spice_transistor_nmos_gnd tM1001(v(vss_v), test_v, test_port_0);
  spice_transistor_nmos_gnd tM1002(v(vss_v), reset_v, reset_port_0);
  spice_transistor_nmos_gnd tM1003(v(N0754_v), N0761_v, N0761_port_0);
  spice_transistor_nmos_gnd tM1004(v(PC0_11_v), N0785_v, N0785_port_0);
  spice_transistor_nmos tM1005(v(N0406_v), N0785_v, N0770_v, N0785_port_1, N0770_port_1);
  spice_transistor_nmos_gnd tM1006(v(N0301_v), N0754_v, N0754_port_1);
  spice_transistor_nmos tM1007(v(N0301_v), N0761_v, N0753_v, N0761_port_1, N0753_port_0);
  spice_transistor_nmos_gnd tM1009(v(N0289_v), N0754_v, N0754_port_3);
  spice_transistor_nmos_gnd tM2085(v(OPR_3_v), FIN_FIM_v, FIN_FIM_port_0);
  spice_transistor_nmos_gnd tM2084(v(OPR_3_v), JCN_v, JCN_port_0);
  spice_transistor_nmos_gnd tM2128(v(_OPR_2_v), N0587_v, N0587_port_2);
  spice_transistor_nmos tM1134(v(N0426_v), N0388_v, PC2_2_v, N0388_port_4, PC2_2_port_0);
  spice_transistor_nmos tM1135(v(N0439_v), PC3_2_v, N0388_v, PC3_2_port_0, N0388_port_5);
  spice_transistor_nmos_gnd tM1136(v(N0775_v), N0389_v, N0389_port_1);
  spice_transistor_nmos_gnd tM1137(v(N0771_v), N0390_v, N0390_port_1);
  spice_transistor_nmos tM1130(v(N0426_v), N0387_v, PC2_3_v, N0387_port_4, PC2_3_port_1);
  spice_transistor_nmos_vdd tM1131(v(__INH__X11_X31_CLK1_v), N0778_v, N0778_port_6);
  spice_transistor_nmos tM1133(v(N0439_v), PC3_3_v, N0387_v, PC3_3_port_1, N0387_port_5);
  spice_transistor_nmos_gnd tM2732(v(INC_GROUP_5__v), N0546_v, N0546_port_0);
  spice_transistor_nmos_gnd tM2730(v(N0675_v), N0659_v, N0659_port_5);
  spice_transistor_nmos tM1138(v(WADB2_v), N0771_v, N0762_v, N0771_port_1, N0762_port_5);
  spice_transistor_nmos tM1139(v(N0406_v), N0789_v, N0775_v, N0789_port_0, N0775_port_2);
  spice_transistor_nmos_gnd tM2735(v(L_v), N0701_v, N0701_port_1);
  spice_transistor_nmos_gnd tM2734(v(L_v), N0686_v, N0686_port_0);
  spice_transistor_nmos_gnd tM2113(v(SC_v), N0644_v, N0644_port_1);
  spice_transistor_nmos tM2112(v(A22_v), N0644_v, N0643_v, N0644_port_0, N0643_port_1);
  spice_transistor_nmos tM2111(v(SC_v), N0662_v, N0661_v, N0662_port_1, N0661_port_0);
  spice_transistor_nmos_gnd tM2110(v(M12_v), N0662_v, N0662_port_0);
  spice_transistor_nmos tM2117(v(OPR_3_v), INC_ISZ_ADD_SUB_XCH_LD_v, N0628_v, INC_ISZ_ADD_SUB_XCH_LD_port_2, N0628_port_1);
  spice_transistor_nmos tM2440(v(N0801_v), N0800_v, N0782_v, N0800_port_0, N0782_port_2);
  spice_transistor_nmos tM2443(v(N0799_v), N0782_v, N0798_v, N0782_port_3, N0798_port_1);
  spice_transistor_nmos tM2114(v(clk2_v), N0661_v, N0660_v, N0661_port_1, N0660_port_0);
  spice_transistor_nmos_gnd tM2119(v(_OPR_2_v), N0523_v, N0523_port_0);
  spice_transistor_nmos_gnd tM2118(v(OPR_3_v), N0587_v, N0587_port_1);
  spice_transistor_nmos_gnd tM2449(v(N0719_v), X22_v, X22_port_7);
  spice_transistor_nmos_vdd tM2448(v(N0742_v), X22_v, X22_port_6);
  spice_transistor_nmos_gnd tM2561(v(N0340_v), N0342_v, N0342_port_1);
  spice_transistor_nmos_gnd tM1649(v(N0542_v), N0570_v, N0570_port_5);
  spice_transistor_nmos_gnd tM1642(v(N0577_v), N0570_v, N0570_port_4);
  spice_transistor_nmos_gnd tM1643(v(N0542_v), N0539_v, N0539_port_2);
  spice_transistor_nmos_gnd tM1640(v(N0541_v), N0599_v, N0599_port_4);
  spice_transistor_nmos_gnd tM1641(v(N0541_v), N0620_v, N0620_port_4);
  spice_transistor_nmos_gnd tM1646(v(N0577_v), N0635_v, N0635_port_4);
  spice_transistor_nmos_gnd tM1647(v(N0577_v), N0648_v, N0648_port_4);
  spice_transistor_nmos_gnd tM1644(v(N0577_v), N0584_v, N0584_port_4);
  spice_transistor_nmos_gnd tM2597(v(CLB_v), WRITE_ACC_1__v, WRITE_ACC_1__port_9);
  spice_transistor_nmos_gnd tM2596(v(N1005_v), _OPA_1_v, _OPA_1_port_7);
  spice_transistor_nmos_gnd tM2595(v(IAC_v), WRITE_ACC_1__v, WRITE_ACC_1__port_8);
  spice_transistor_nmos_gnd tM2593(v(TCC_v), WRITE_ACC_1__v, WRITE_ACC_1__port_6);
  spice_transistor_nmos_gnd tM2592(v(CMA_v), WRITE_ACC_1__v, WRITE_ACC_1__port_5);
  spice_transistor_nmos_gnd tM2591(v(POC_v), WRITE_CARRY_2__v, WRITE_CARRY_2__port_1);
  spice_transistor_nmos_gnd tM2590(v(INC_ISZ_v), INC_GROUP_5__v, INC_GROUP_5__port_0);
  spice_transistor_nmos_gnd tM2126(v(OPR_3_v), JUN2_JMS2_v, JUN2_JMS2_port_0);
  spice_transistor_nmos_vdd tM2599(v(N1005_v), OPA_1_v, OPA_1_port_11);
  spice_transistor_nmos tM2127(v(_OPR_2_v), N0628_v, INC_ISZ_ADD_SUB_XCH_LD_v, N0628_port_2, INC_ISZ_ADD_SUB_XCH_LD_port_3);
  spice_transistor_nmos_gnd tM2027(v(_OPR_3_v), IO_v, IO_port_0);
  spice_transistor_nmos_gnd tM2025(v(N0590_v), N0564_v, N0564_port_0);
  spice_transistor_nmos tM2024(v(X32_v), N0612_v, N0611_v, N0612_port_1, N0611_port_0);
  spice_transistor_nmos_vdd tM2023(v(S00627_v), N0626_v, N0626_port_1);
  spice_transistor_nmos tM2022(v(clk2_v), N0649_v, N0650_v, N0649_port_2, N0650_port_0);
  spice_transistor_nmos tM2021(v(clk2_v), N0655_v, N0656_v, N0655_port_2, N0656_port_0);
  spice_transistor_nmos_gnd tM2029(v(DC_v), INC_ISZ_v, INC_ISZ_port_0);
  spice_transistor_nmos_gnd tM2028(v(_OPR_3_v), OPE_v, OPE_port_0);
  spice_transistor_nmos tM1245(v(N0424_v), N0780_v, N0814_v, N0780_port_3, N0814_port_1);
  spice_transistor_nmos tM1242(v(N0381_v), N0393_v, PC0_1_v, N0393_port_2, PC0_1_port_1);
  spice_transistor_nmos_gnd tM1243(v(PC1_1_v), N0814_v, N0814_port_0);
  spice_transistor_nmos tM1240(v(N0444_v), N0776_v, N0841_v, N0776_port_5, N0841_port_1);
  spice_transistor_nmos_gnd tM2206(v(_OPR_0_v), JCN_ISZ_v, JCN_ISZ_port_7);
  spice_transistor_nmos_gnd tM2205(v(_OPR_0_v), XCH_v, XCH_port_3);
  spice_transistor_nmos_gnd tM1241(v(N0781_v), N0394_v, N0394_port_1);
  spice_transistor_nmos tM2203(v(clk2_v), N0362_v, N0368_v, N0362_port_1, N0368_port_2);
  spice_transistor_nmos tM2202(v(N0343_v), N0368_v, N0367_v, N0368_port_1, N0367_port_1);
  spice_transistor_nmos_gnd tM2201(v(N0352_v), N0367_v, N0367_port_0);
  spice_transistor_nmos_gnd tM2200(v(X32_v), N0352_v, N0352_port_1);
  spice_transistor_nmos_vdd tM3089(v(S00803_v), ACC_ADA_v, ACC_ADA_port_5);
  spice_transistor_nmos_gnd tM3086(v(N0666_v), N0665_v, N0665_port_2);
  spice_transistor_nmos_vdd tM3084(v(N0690_v), d2_v, d2_port_2);
  spice_transistor_nmos tM3083(v(SUB_GROUP_6__v), TMP_2_v, N0891_v, TMP_2_port_2, N0891_port_5);
  spice_transistor_nmos_vdd tM3081(v(N0944_v), TMP_2_v, TMP_2_port_0);
  spice_transistor_nmos_gnd tM3240(v(vss_v), d1_v, d1_port_0);
  spice_transistor_nmos_gnd tM2997(v(N0851_v), N0348_v, N0348_port_1);
  spice_transistor_nmos_gnd tM3243(v(N0676_v), N0670_v, N0670_port_3);
  spice_transistor_nmos_gnd tM3244(v(N0676_v), N0669_v, N0669_port_1);
  spice_transistor_nmos_vdd tM3245(v(N0669_v), D0_v, D0_port_17);
  spice_transistor_nmos_gnd tM2150(v(_OPR_1_v), N0523_v, N0523_port_2);
  spice_transistor_nmos_gnd tM2919(v(N0871_v), N0895_v, N0895_port_1);
  spice_transistor_nmos tM2912(v(ADD_IB_v), N0847_v, D1_v, N0847_port_3, D1_port_12);
  spice_transistor_nmos_gnd tM1331(v(R9_1_v), N0959_v, N0959_port_1);
  spice_transistor_nmos tM1898(v(N0571_v), REG_RFSH_1_v, N0593_v, REG_RFSH_1_port_2, N0593_port_0);
  spice_transistor_nmos_gnd tM1897(v(N0571_v), N0574_v, N0574_port_3);
  spice_transistor_nmos_gnd tM1903(v(N0506_v), N0509_v, N0509_port_0);
  spice_transistor_nmos tM1902(v(CLK2_JMS_DC_M22_BBL_M22_X12_X22___v), N0520_v, N0466_v, N0520_port_1, N0466_port_6);
  spice_transistor_nmos_gnd tM1905(v(N0592_v), RRAB1_v, RRAB1_port_5);
  spice_transistor_nmos tM1904(v(CLK2_JMS_DC_M22_BBL_M22_X12_X22___v), N0459_v, N0509_v, N0459_port_6, N0509_port_1);
  spice_transistor_nmos_gnd tM1896(v(N0571_v), N0573_v, N0573_port_2);
  spice_transistor_nmos_gnd tM1909(v(DC_v), RRAB1_v, RRAB1_port_6);
  spice_transistor_nmos_gnd tM1894(v(N0574_v), N0571_v, N0571_port_2);
  spice_transistor_nmos tM1891(v(SC_A12_CLK2_v), N0571_v, N0572_v, N0571_port_1, N0572_port_0);
  spice_transistor_nmos tM1890(v(clk1_v), REG_RFSH_0_v, N0566_v, REG_RFSH_0_port_2, N0566_port_0);
  spice_transistor_nmos_gnd tM2768(v(N0678_v), N0677_v, N0677_port_1);
  spice_transistor_nmos_gnd tM1144(v(PC2_2_v), N0824_v, N0824_port_1);
  spice_transistor_nmos_vdd tM2681(v(S00676_v), N0702_v, N0702_port_1);
  spice_transistor_nmos_gnd tM2680(v(N1006_v), OPA_0_v, OPA_0_port_12);
  spice_transistor_nmos_gnd tM1141(v(PC1_2_v), N0809_v, N0809_port_0);
  spice_transistor_nmos_gnd tM1140(v(PC0_6_v), N0789_v, N0789_port_1);
  spice_transistor_nmos_gnd tM1839(v(N0517_v), __INH__X11_X31_CLK1_v, __INH__X11_X31_CLK1_port_13);
  spice_transistor_nmos tM1143(v(N0434_v), N0824_v, N0779_v, N0824_port_0, N0779_port_4);
  spice_transistor_nmos_vdd tM1834(v(S00628_v), __INH__X11_X31_CLK1_v, __INH__X11_X31_CLK1_port_12);
  spice_transistor_nmos_gnd tM1837(v(N0436_v), N0437_v, N0437_port_2);
  spice_transistor_nmos_vdd tM1836(v(N0436_v), ___SC__JIN_FIN__CLK1_M11_X21_INH__v, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_5);
  spice_transistor_nmos_vdd tM1831(v(S00612_v), N0436_v, N0436_port_0);
  spice_transistor_nmos_gnd tM1830(v(N0437_v), ___SC__JIN_FIN__CLK1_M11_X21_INH__v, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_4);
  spice_transistor_nmos_gnd tM2761(v(N0342_v), CY_ADA_v, CY_ADA_port_2);
  spice_transistor_nmos tM1060(v(N0292_v), N0313_v, N0305_v, N0313_port_1, N0305_port_0);
  spice_transistor_nmos_vdd tM1066(v(N0325_v), N0305_v, N0305_port_1);
  spice_transistor_nmos_gnd tM2765(v(WRITE_ACC_1__v), ADD_ACC_v, ADD_ACC_port_0);
  spice_transistor_nmos_gnd tM2904(v(N0350_v), N0376_v, N0376_port_1);
  spice_transistor_nmos_gnd tM2905(v(N0767_v), DCL_0_v, DCL_0_port_4);
  spice_transistor_nmos_gnd tM2906(v(N0350_v), N0345_v, N0345_port_1);
  spice_transistor_nmos_gnd tM2907(v(N0350_v), N0354_v, N0354_port_1);
  spice_transistor_nmos_gnd tM2900(v(N0351_v), N0766_v, N0766_port_1);
  spice_transistor_nmos_gnd tM2901(v(DCL_0_v), N0716_v, N0716_port_0);
  spice_transistor_nmos_gnd tM1347(v(R0_2_v), N0908_v, N0908_port_1);
  spice_transistor_nmos tM1346(v(N0543_v), N0908_v, N0882_v, N0908_port_0, N0882_port_2);
  spice_transistor_nmos tM1345(v(N0544_v), R2_2_v, N0536_v, R2_2_port_0, N0536_port_3);
  spice_transistor_nmos tM1344(v(N0529_v), N0536_v, R0_2_v, N0536_port_2, R0_2_port_0);
  spice_transistor_nmos tM1343(v(N0544_v), R3_2_v, N0535_v, R3_2_port_1, N0535_port_3);
  spice_transistor_nmos tM1342(v(N0529_v), N0535_v, R1_2_v, N0535_port_2, R1_2_port_1);
  spice_transistor_nmos_gnd tM1341(v(R7_2_v), N0951_v, N0951_port_0);
  spice_transistor_nmos_gnd tM1340(v(R13_1_v), N0978_v, N0978_port_1);
  spice_transistor_nmos tM1349(v(N0616_v), N0960_v, N0868_v, N0960_port_0, N0868_port_6);
  spice_transistor_nmos tM1348(v(N0591_v), N0868_v, N0951_v, N0868_port_5, N0951_port_1);
  spice_transistor_nmos_gnd tM2694(v(N1013_v), N1002_v, N1002_port_3);
  spice_transistor_nmos_gnd tM2695(v(N1015_v), N1006_v, N1006_port_3);
  spice_transistor_nmos_gnd tM2690(v(JUN2_JMS2_v), N0658_v, N0658_port_0);
  spice_transistor_nmos_gnd tM2691(v(N1002_v), N1003_v, N1003_port_3);
  spice_transistor_nmos tM1019(v(M12_M22_CLK1__M11_M12__v), N0290_v, D2_v, N0290_port_0, D2_port_0);
  spice_transistor_nmos tM1018(v(RADB0_v), N0387_v, D3_v, N0387_port_0, D3_port_3);
  spice_transistor_nmos tM1017(v(M12_M22_CLK1__M11_M12__v), N0289_v, D3_v, N0289_port_3, D3_port_2);
  spice_transistor_nmos_vdd tM1016(v(N0325_v), N0301_v, N0301_port_2);
  spice_transistor_nmos_gnd tM1015(v(N0289_v), N0311_v, N0311_port_0);
  spice_transistor_nmos tM1014(v(WADB2_v), N0770_v, N0761_v, N0770_port_2, N0761_port_3);
  spice_transistor_nmos tM1012(v(RADB1_v), D3_v, N0386_v, D3_port_0, N0386_port_0);
  spice_transistor_nmos_gnd tM1011(v(N0289_v), N0753_v, N0753_port_1);
  spice_transistor_nmos_gnd tM1123(v(PC3_3_v), N0836_v, N0836_port_0);
  spice_transistor_nmos tM1121(v(RRAB0_v), N0532_v, D0_v, N0532_port_0, D0_port_4);
  spice_transistor_nmos tM1120(v(RRAB1_v), D0_v, N0531_v, D0_port_3, N0531_port_1);
  spice_transistor_nmos tM1127(v(N0410_v), PC1_2_v, N0388_v, PC1_2_port_0, N0388_port_3);
  spice_transistor_nmos tM1126(v(N0381_v), N0388_v, PC0_2_v, N0388_port_2, PC0_2_port_0);
  spice_transistor_nmos tM1125(v(N0410_v), PC1_3_v, N0387_v, PC1_3_port_1, N0387_port_3);
  spice_transistor_nmos tM1124(v(N0444_v), N0778_v, N0836_v, N0778_port_5, N0836_port_1);
  spice_transistor_nmos_gnd tM1129(v(PC0_2_v), N0788_v, N0788_port_1);
  spice_transistor_nmos tM1128(v(N0406_v), N0788_v, N0779_v, N0788_port_0, N0779_port_2);
  spice_transistor_nmos_gnd tM2474(v(OPA_1_v), RAL_v, RAL_port_4);
  spice_transistor_nmos_gnd tM2475(v(OPA_1_v), CMA_v, CMA_port_4);
  spice_transistor_nmos_gnd tM2476(v(OPA_1_v), DAC_v, DAC_port_4);
  spice_transistor_nmos_gnd tM2477(v(OPA_1_v), CLC_v, CLC_port_4);
  spice_transistor_nmos_gnd tM2478(v(OPA_1_v), CLB_v, CLB_port_4);
  spice_transistor_nmos_gnd tM2479(v(OPA_1_v), SBM_v, SBM_port_4);
  spice_transistor_nmos_gnd tM1659(v(N0542_v), N0599_v, N0599_port_5);
  spice_transistor_nmos_gnd tM1658(v(N0504_v), N0508_v, N0508_port_0);
  spice_transistor_nmos tM1173(v(N0529_v), N0532_v, R0_0_v, N0532_port_2, R0_0_port_0);
  spice_transistor_nmos tM1651(v(N0427_v), N0426_v, ___SC__JIN_FIN__CLK1_M11_X21_INH__v, N0426_port_13, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_2);
  spice_transistor_nmos tM1650(v(N0427_v), N0434_v, __POC_CLK2_X12_X32__INH_v, N0434_port_13, __POC_CLK2_X12_X32__INH_port_2);
  spice_transistor_nmos tM1653(v(N0440_v), N0444_v, __POC_CLK2_X12_X32__INH_v, N0444_port_13, __POC_CLK2_X12_X32__INH_port_3);
  spice_transistor_nmos tM1652(v(N0440_v), N0439_v, ___SC__JIN_FIN__CLK1_M11_X21_INH__v, N0439_port_13, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_3);
  spice_transistor_nmos_gnd tM1655(v(N0382_v), N0783_v, N0783_port_2);
  spice_transistor_nmos_gnd tM1654(v(N0519_v), N0518_v, N0518_port_0);
  spice_transistor_nmos tM1657(v(__INH__X32_CLK2_v), N0518_v, N0463_v, N0518_port_1, N0463_port_6);
  spice_transistor_nmos_gnd tM1656(v(N0411_v), N0804_v, N0804_port_2);
  spice_transistor_nmos tM2874(v(N0553_v), N0898_v, N0878_v, N0898_port_0, N0878_port_4);
  spice_transistor_nmos_gnd tM2876(v(N0550_v), N0898_v, N0898_port_2);
  spice_transistor_nmos tM2053(v(clk2_v), N0622_v, N0623_v, N0622_port_3, N0623_port_0);
  spice_transistor_nmos_gnd tM2056(v(A12_v), N0618_v, N0618_port_1);
  spice_transistor_nmos_gnd tM2057(v(A22_v), N0654_v, N0654_port_2);
  spice_transistor_nmos_gnd tM2054(v(M12_v), N0618_v, N0618_port_0);
  spice_transistor_nmos tM2055(v(X12_v), N0682_v, N0683_v, N0682_port_0, N0683_port_0);
  spice_transistor_nmos_vdd tM2791(v(N0546_v), N0550_v, N0550_port_2);
  spice_transistor_nmos tM2058(v(clk2_v), N0578_v, N0575_v, N0578_port_1, N0575_port_2);
  spice_transistor_nmos_gnd tM3258(v(N0716_v), N0736_v, N0736_port_1);
  spice_transistor_nmos_gnd tM2273(v(_I_O_v), IOW_v, IOW_port_1);
  spice_transistor_nmos_gnd tM3099(v(N0731_v), N0748_v, N0748_port_1);
  spice_transistor_nmos_gnd tM1521(v(A22_v), N0712_v, N0712_port_1);
  spice_transistor_nmos_vdd tM3094(v(N0748_v), A12_v, A12_port_9);
  spice_transistor_nmos_gnd tM3097(v(N0731_v), A12_v, A12_port_10);
  spice_transistor_nmos_gnd tM1520(v(N0737_v), cm_rom_v, cm_rom_port_1);
  spice_transistor_nmos_gnd tM3091(v(A12_v), N0288_v, N0288_port_6);
  spice_transistor_nmos_gnd tM2306(v(__X31__CLK2__v), N0480_v, N0480_port_0);
  spice_transistor_nmos_gnd tM2966(v(N0879_v), N0848_v, N0848_port_1);
  spice_transistor_nmos_gnd tM2304(v(_I_O_v), ADM_v, ADM_port_1);
  spice_transistor_nmos_gnd tM2303(v(_I_O_v), SBM_v, SBM_port_1);
  spice_transistor_nmos_gnd tM3259(v(N0733_v), cm_ram1_v, cm_ram1_port_1);
  spice_transistor_nmos tM2301(v(OPA_IB_v), D3_v, OPA_3_v, D3_port_9, OPA_3_port_0);
  spice_transistor_nmos_vdd tM3255(v(N0716_v), cm_ram0_v, cm_ram0_port_0);
  spice_transistor_nmos_vdd tM3254(v(N0713_v), cm_ram1_v, cm_ram1_port_0);
  spice_transistor_nmos_gnd tM3253(v(N0713_v), N0733_v, N0733_port_0);
  spice_transistor_nmos tM2308(v(N0480_v), N0482_v, N0477_v, N0482_port_0, N0477_port_1);
  spice_transistor_nmos tM3250(v(N0702_v), N0674_v, N0697_v, N0674_port_2, N0697_port_0);
  spice_transistor_nmos_gnd tM2965(v(N0346_v), N0376_v, N0376_port_2);
  spice_transistor_nmos_gnd tM2610(v(CLC_v), WRITE_CARRY_2__v, WRITE_CARRY_2__port_8);
  spice_transistor_nmos_gnd tM2611(v(CLB_v), WRITE_CARRY_2__v, WRITE_CARRY_2__port_9);
  spice_transistor_nmos tM2940(v(N0871_v), N0552_v, N0912_v, N0552_port_2, N0912_port_1);
  spice_transistor_nmos tM2469(v(clk2_v), N0380_v, N0383_v, N0380_port_0, N0383_port_1);
  spice_transistor_nmos_gnd tM3055(v(N0348_v), N0370_v, N0370_port_4);
  spice_transistor_nmos_vdd tM2468(v(S00699_v), N0782_v, N0782_port_5);
  spice_transistor_nmos_gnd tM3056(v(N0348_v), N0376_v, N0376_port_4);
  spice_transistor_nmos_gnd tM2463(v(N0721_v), X12_v, X12_port_13);
  spice_transistor_nmos_gnd tM3251(v(N0697_v), N0696_v, N0696_port_0);
  spice_transistor_nmos_gnd tM1938(v(SC_v), N0525_v, N0525_port_0);
  spice_transistor_nmos tM1939(v(JIN_FIN_v), N0525_v, N0524_v, N0525_port_1, N0524_port_1);
  spice_transistor_nmos_gnd tM1937(v(_CN_v), N0528_v, N0528_port_1);
  spice_transistor_nmos_gnd tM2863(v(N0856_v), N0471_v, N0471_port_2);
  spice_transistor_nmos_gnd tM3117(v(N0354_v), N0358_v, N0358_port_2);
  spice_transistor_nmos_gnd tM2862(v(N0887_v), N0549_v, N0549_port_1);
  spice_transistor_nmos tM2860(v(N0887_v), N0878_v, N0886_v, N0878_port_2, N0886_port_1);
  spice_transistor_nmos_vdd tM1800(v(S00601_v), N0440_v, N0440_port_5);
  spice_transistor_nmos tM1801(v(X12_v), N0409_v, ADDR_RFSH_1_v, N0409_port_3, ADDR_RFSH_1_port_3);
  spice_transistor_nmos tM1802(v(X32_v), ADDR_PTR_1_v, N0409_v, ADDR_PTR_1_port_3, N0409_port_4);
  spice_transistor_nmos tM1803(v(X12_v), N0420_v, ADDR_RFSH_0_v, N0420_port_3, ADDR_RFSH_0_port_3);
  spice_transistor_nmos tM2947(v(ADD_ACC_v), N0847_v, ACC_1_v, N0847_port_5, ACC_1_port_3);
  spice_transistor_nmos_vdd tM2462(v(N0743_v), X12_v, X12_port_12);
  spice_transistor_nmos_gnd tM2868(v(N0705_v), N0700_v, N0700_port_3);
  spice_transistor_nmos_vdd tM1248(v(__INH__X11_X31_CLK1_v), N0772_v, N0772_port_6);
  spice_transistor_nmos tM1246(v(N0434_v), N0829_v, N0780_v, N0829_port_1, N0780_port_4);
  spice_transistor_nmos_gnd tM1244(v(PC2_1_v), N0829_v, N0829_port_0);
  spice_transistor_nmos_gnd tM2911(v(N0847_v), ADD_0_v, ADD_0_port_3);
  spice_transistor_nmos tM2917(v(ACC_ADAC_v), N0871_v, N0472_v, N0871_port_0, N0472_port_0);
  spice_transistor_nmos tM2916(v(ACB_IB_v), D1_v, N0347_v, D1_port_13, N0347_port_1);
  spice_transistor_nmos_vdd tM2914(v(N0875_v), N0847_v, N0847_port_4);
  spice_transistor_nmos tM1332(v(N0619_v), R11_1_v, N0534_v, R11_1_port_0, N0534_port_7);
  spice_transistor_nmos tM1333(v(N0634_v), N0533_v, R12_1_v, N0533_port_8, R12_1_port_1);
  spice_transistor_nmos tM1330(v(N0616_v), N0959_v, N0867_v, N0959_port_0, N0867_port_6);
  spice_transistor_nmos tM1336(v(N0634_v), N0534_v, R13_1_v, N0534_port_8, R13_1_port_0);
  spice_transistor_nmos_gnd tM1337(v(R11_1_v), N0969_v, N0969_port_0);
  spice_transistor_nmos tM1334(v(N0657_v), N0881_v, N0986_v, N0881_port_9, N0986_port_1);
  spice_transistor_nmos tM1335(v(N0647_v), R14_1_v, N0533_v, R14_1_port_1, N0533_port_9);
  spice_transistor_nmos tM1338(v(N0632_v), N0867_v, N0969_v, N0867_port_7, N0969_port_1);
  spice_transistor_nmos tM1339(v(N0645_v), N0978_v, N0867_v, N0978_port_0, N0867_port_8);
  spice_transistor_nmos_gnd tM2683(v(D3_v), N0671_v, N0671_port_2);
  spice_transistor_nmos tM1799(v(SC_A22_v), N0617_v, REG_RFSH_1_v, N0617_port_2, REG_RFSH_1_port_1);
  spice_transistor_nmos_vdd tM1068(v(N0325_v), N0752_v, N0752_port_0);
  spice_transistor_nmos tM1069(v(N0752_v), N0764_v, N0759_v, N0764_port_0, N0759_port_1);
  spice_transistor_nmos_gnd tM2687(v(N1004_v), N1005_v, N1005_port_3);
  spice_transistor_nmos tM1062(v(N0292_v), N0299_v, N0294_v, N0299_port_1, N0294_port_1);
  spice_transistor_nmos tM1063(v(N0292_v), N0293_v, N0294_v, N0293_port_3, N0294_port_2);
  spice_transistor_nmos tM1061(v(N0292_v), N0303_v, N0294_v, N0303_port_1, N0294_port_0);
  spice_transistor_nmos tM1794(v(SC_A22_v), N0582_v, REG_RFSH_0_v, N0582_port_2, REG_RFSH_0_port_0);
  spice_transistor_nmos tM1067(v(RADB0_v), N0394_v, D0_v, N0394_port_0, D0_port_1);
  spice_transistor_nmos tM1064(v(M12_M22_CLK1__M11_M12__v), N0292_v, D0_v, N0292_port_4, D0_port_0);
  spice_transistor_nmos_gnd tM1065(v(N0292_v), N0759_v, N0759_port_0);
  spice_transistor_nmos_gnd tM1488(v(vss_v), clk2_v, clk2_port_0);
  spice_transistor_nmos_gnd tM1489(v(vss_v), clk1_v, clk1_port_0);
  spice_transistor_nmos tM1484(v(N0632_v), N0869_v, N0973_v, N0869_port_7, N0973_port_1);
  spice_transistor_nmos tM1485(v(N0645_v), N0982_v, N0869_v, N0982_port_0, N0869_port_8);
  spice_transistor_nmos_gnd tM1486(v(R13_3_v), N0982_v, N0982_port_1);
  spice_transistor_nmos_vdd tM1480(v(SC_A22_M22_CLK2_v), N0883_v, N0883_port_10);
  spice_transistor_nmos tM1481(v(N0647_v), R14_3_v, N0537_v, R14_3_port_1, N0537_port_9);
  spice_transistor_nmos tM1482(v(N0634_v), N0538_v, R13_3_v, N0538_port_8, R13_3_port_0);
  spice_transistor_nmos tM1483(v(N0647_v), R15_3_v, N0538_v, R15_3_port_0, N0538_port_9);
  spice_transistor_nmos tM1664(v(__FIN_X12__v), N0539_v, N0530_v, N0539_port_3, N0530_port_3);
  spice_transistor_nmos_gnd tM1666(v(__FIN_X12__v), N0561_v, N0561_port_1);
  spice_transistor_nmos_gnd tM1660(v(N0542_v), N0635_v, N0635_port_5);
  spice_transistor_nmos_gnd tM1661(v(N0577_v), N0541_v, N0541_port_5);
  spice_transistor_nmos_gnd tM1662(v(N0617_v), N0577_v, N0577_port_5);
  spice_transistor_nmos tM1663(v(__INH__X32_CLK2_v), N0455_v, N0508_v, N0455_port_6, N0508_port_1);
  spice_transistor_nmos_vdd tM2467(v(S00725_v), N0743_v, N0743_port_2);
  spice_transistor_nmos_gnd tM2465(v(N0721_v), N0743_v, N0743_port_1);
  spice_transistor_nmos_gnd tM1668(v(N0427_v), N0820_v, N0820_port_2);
  spice_transistor_nmos_gnd tM1669(v(N0440_v), N0833_v, N0833_port_3);
  spice_transistor_nmos_gnd tM2461(v(X12_v), N0288_v, N0288_port_1);
  spice_transistor_nmos_vdd tM1467(v(SC_A22_M22_CLK2_v), N0882_v, N0882_port_10);
  spice_transistor_nmos_vdd tM1464(v(SC_A22_M22_CLK2_v), N0868_v, N0868_port_10);
  spice_transistor_nmos_gnd tM1462(v(R14_2_v), N0989_v, N0989_port_0);
  spice_transistor_nmos tM1463(v(N0657_v), N0882_v, N0989_v, N0882_port_9, N0989_port_1);
  spice_transistor_nmos tM1460(v(N0645_v), N0981_v, N0883_v, N0981_port_0, N0883_port_8);
  spice_transistor_nmos_gnd tM1461(v(R12_3_v), N0981_v, N0981_port_1);
  spice_transistor_nmos_gnd tM1468(v(R14_3_v), N0990_v, N0990_port_0);
  spice_transistor_nmos tM1469(v(N0657_v), N0883_v, N0990_v, N0883_port_9, N0990_port_1);
  spice_transistor_nmos_gnd tM2861(v(N0870_v), N0548_v, N0548_port_1);
  spice_transistor_nmos_gnd tM2867(v(N0940_v), _TMP_0_v, _TMP_0_port_0);
  spice_transistor_nmos tM2866(v(N0887_v), N0911_v, N0548_v, N0911_port_1, N0548_port_2);
  spice_transistor_nmos tM2865(v(N0870_v), N0549_v, N0911_v, N0549_port_2, N0911_port_0);
  spice_transistor_nmos tM2040(v(INC_ISZ_XCH_v), N0603_v, N0611_v, N0603_port_1, N0611_port_1);
  spice_transistor_nmos_gnd tM2043(v(N0568_v), N0579_v, N0579_port_0);
  spice_transistor_nmos tM2045(v(N0580_v), N0575_v, N0579_v, N0575_port_1, N0579_port_1);
  spice_transistor_nmos_gnd tM2044(v(N0568_v), N0567_v, N0567_port_1);
  spice_transistor_nmos tM2047(v(A12_v), N0651_v, N0650_v, N0651_port_0, N0650_port_1);
  spice_transistor_nmos tM2046(v(SC_v), N0654_v, N0656_v, N0654_port_0, N0656_port_1);
  spice_transistor_nmos_gnd tM2049(v(M22_v), N0654_v, N0654_port_1);
  spice_transistor_nmos_gnd tM2048(v(SC_v), N0651_v, N0651_port_1);
  spice_transistor_nmos tM1980(v(JCN_ISZ_v), N0527_v, N0524_v, N0527_port_1, N0524_port_2);
  spice_transistor_nmos tM1983(v(X22_v), N0467_v, N0468_v, N0467_port_4, N0468_port_2);
  spice_transistor_nmos tM1982(v(M22_v), N0468_v, N0467_v, N0468_port_1, N0467_port_3);
  spice_transistor_nmos tM1987(v(X12_v), N0608_v, N0602_v, N0608_port_2, N0602_port_0);
  spice_transistor_nmos_gnd tM1986(v(clk2_v), RRAB0_v, RRAB0_port_7);
  spice_transistor_nmos_gnd tM2315(v(clk2_v), N0297_v, N0297_port_0);
  spice_transistor_nmos_gnd tM2314(v(N0769_v), N0327_v, N0327_port_3);
  spice_transistor_nmos tM2317(v(clk2_v), X22_v, N0280_v, X22_port_5, N0280_port_0);
  spice_transistor_nmos tM2979(v(N0702_v), N0691_v, N0672_v, N0691_port_0, N0672_port_2);
  spice_transistor_nmos_gnd tM2311(v(IOR_v), N0479_v, N0479_port_2);
  spice_transistor_nmos_gnd tM2310(v(N0479_v), N0482_v, N0482_port_1);
  spice_transistor_nmos tM2313(v(N0419_v), N0418_v, N0413_v, N0418_port_1, N0413_port_1);
  spice_transistor_nmos tM2312(v(N0399_v), N0412_v, N0413_v, N0412_port_1, N0413_port_0);
  spice_transistor_nmos_vdd tM3222(v(M12_v), N0607_v, N0607_port_0);
  spice_transistor_nmos tM3223(v(N0937_v), TMP_3_v, N0893_v, TMP_3_port_0, N0893_port_5);
  spice_transistor_nmos_gnd tM3221(v(N0945_v), N0946_v, N0946_port_2);
  spice_transistor_nmos_vdd tM2318(v(S00678_v), N0297_v, N0297_port_1);
  spice_transistor_nmos_vdd tM3224(v(N0946_v), TMP_3_v, TMP_3_port_1);
  spice_transistor_nmos_vdd tM3225(v(N0914_v), N0861_v, N0861_port_3);
  spice_transistor_nmos_vdd tM1504(v(__INH__X11_X31_CLK1_v), N0781_v, N0781_port_6);
  spice_transistor_nmos_gnd tM3136(v(_COM_v), N0715_v, N0715_port_1);
  spice_transistor_nmos_gnd tM3137(v(N0354_v), N0366_v, N0366_port_1);
  spice_transistor_nmos_vdd tM3134(v(N0714_v), cm_ram3_v, cm_ram3_port_0);
  spice_transistor_nmos_gnd tM3135(v(N0714_v), N0734_v, N0734_port_0);
  spice_transistor_nmos_gnd tM3133(v(N0750_v), N0715_v, N0715_port_0);
  spice_transistor_nmos_gnd tM1502(v(N0919_v), N0565_v, N0565_port_8);
  spice_transistor_nmos_gnd tM3138(v(N0363_v), N0366_v, N0366_port_2);
  spice_transistor_nmos_gnd tM3139(v(N0370_v), N0366_v, N0366_port_3);
  spice_transistor_nmos_gnd tM2790(v(M12_v), N0550_v, N0550_port_1);
  spice_transistor_nmos_vdd tM2816(v(S00761_v), N0745_v, N0745_port_2);
  spice_transistor_nmos_vdd tM2545(v(N0332_v), N0342_v, N0342_port_0);
  spice_transistor_nmos_gnd tM2815(v(_COM_v), N0717_v, N0717_port_4);
  spice_transistor_nmos_gnd tM2931(v(N0346_v), N0371_v, N0371_port_2);
  spice_transistor_nmos_gnd tM2810(v(N0870_v), N0894_v, N0894_port_1);
  spice_transistor_nmos_gnd tM2930(v(N0371_v), N0370_v, N0370_port_2);
  spice_transistor_nmos_gnd tM2811(v(CY_1_v), N0803_v, N0803_port_1);
  spice_transistor_nmos tM1929(v(_INH_v), N0428_v, N0429_v, N0428_port_1, N0429_port_1);
  spice_transistor_nmos tM1928(v(clk2_v), N0438_v, N0428_v, N0438_port_1, N0428_port_0);
  spice_transistor_nmos_gnd tM1923(v(N0524_v), INH_v, INH_port_4);
  spice_transistor_nmos_gnd tM1922(v(INH_v), _INH_v, _INH_port_1);
  spice_transistor_nmos tM1921(v(X32_v), N0496_v, N0495_v, N0496_port_1, N0495_port_0);
  spice_transistor_nmos_gnd tM1920(v(clk2_v), N0496_v, N0496_port_0);
  spice_transistor_nmos_gnd tM1927(v(X12_v), N0429_v, N0429_port_0);
  spice_transistor_nmos tM1926(v(_INH_v), N0495_v, N0494_v, N0495_port_1, N0494_port_2);
  spice_transistor_nmos_gnd tM1925(v(clk1_v), N0522_v, N0522_port_2);
  spice_transistor_nmos_gnd tM1924(v(M22_v), N0511_v, N0511_port_2);
  spice_transistor_nmos_vdd tM2976(v(S00766_v), N0692_v, N0692_port_0);
  spice_transistor_nmos tM1186(v(N0406_v), N0790_v, N0771_v, N0790_port_0, N0771_port_2);
  spice_transistor_nmos tM2819(v(clk2_v), N0284_v, A32_v, N0284_port_1, A32_port_6);
  spice_transistor_nmos tM1817(v(X22_v), N0308_v, N0304_v, N0308_port_0, N0304_port_2);
  spice_transistor_nmos_gnd tM1815(v(N0450_v), __POC_CLK2_X12_X32__INH_v, __POC_CLK2_X12_X32__INH_port_5);
  spice_transistor_nmos_vdd tM1814(v(S00613_v), N0449_v, N0449_port_1);
  spice_transistor_nmos_gnd tM1813(v(JUN_JMS_v), N0309_v, N0309_port_0);
  spice_transistor_nmos_vdd tM1811(v(N0449_v), __POC_CLK2_X12_X32__INH_v, __POC_CLK2_X12_X32__INH_port_4);
  spice_transistor_nmos_gnd tM1819(v(M12_v), N0323_v, N0323_port_0);
  spice_transistor_nmos tM1818(v(N0310_v), N0309_v, N0308_v, N0309_port_1, N0308_port_1);
  spice_transistor_nmos tM1259(v(N0569_v), N0532_v, R4_0_v, N0532_port_4, R4_0_port_0);
  spice_transistor_nmos tM1258(v(N0581_v), N0930_v, N0880_v, N0930_port_0, N0880_port_4);
  spice_transistor_nmos tM1255(v(N0543_v), N0905_v, N0881_v, N0905_port_1, N0881_port_2);
  spice_transistor_nmos_gnd tM1254(v(N0867_v), N0534_v, N0534_port_1);
  spice_transistor_nmos tM1257(v(N0565_v), N0880_v, N0921_v, N0880_port_3, N0921_port_1);
  spice_transistor_nmos_gnd tM1256(v(R2_0_v), N0921_v, N0921_port_0);
  spice_transistor_nmos_gnd tM1251(v(N0500_v), N0865_v, N0865_port_1);
  spice_transistor_nmos_gnd tM1253(v(N0881_v), N0533_v, N0533_port_1);
  spice_transistor_nmos tM1252(v(RRAB0_v), N0536_v, D2_v, N0536_port_0, D2_port_6);
  spice_transistor_nmos tM1321(v(N0598_v), N0534_v, R9_1_v, N0534_port_6, R9_1_port_0);
  spice_transistor_nmos tM1320(v(N0619_v), R10_1_v, N0533_v, R10_1_port_1, N0533_port_7);
  spice_transistor_nmos tM1323(v(WRAB0_v), N0882_v, N0864_v, N0882_port_1, N0864_port_3);
  spice_transistor_nmos_gnd tM1322(v(N0882_v), N0536_v, N0536_port_1);
  spice_transistor_nmos_gnd tM1324(v(R3_2_v), N0924_v, N0924_port_0);
  spice_transistor_nmos_gnd tM1327(v(R5_2_v), N0933_v, N0933_port_1);
  spice_transistor_nmos tM1326(v(N0581_v), N0933_v, N0868_v, N0933_port_0, N0868_port_4);
  spice_transistor_nmos tM1329(v(N0591_v), N0867_v, N0950_v, N0867_port_5, N0950_port_1);
  spice_transistor_nmos_gnd tM1328(v(R7_1_v), N0950_v, N0950_port_0);
  spice_transistor_nmos tM1078(v(N0307_v), N0305_v, N0306_v, N0305_port_2, N0306_port_0);
  spice_transistor_nmos_gnd tM1073(v(N0307_v), N0294_v, N0294_port_3);
  spice_transistor_nmos_gnd tM1075(v(N0307_v), N0752_v, N0752_port_3);
  spice_transistor_nmos_gnd tM1074(v(N0752_v), N0760_v, N0760_port_2);
  spice_transistor_nmos_gnd tM1077(v(N0738_v), N0740_v, N0740_port_2);
  spice_transistor_nmos_gnd tM1076(v(N0760_v), N0764_v, N0764_port_2);
  spice_transistor_nmos_gnd tM3227(v(N0945_v), TMP_3_v, TMP_3_port_2);
  spice_transistor_nmos_gnd tM1499(v(N0902_v), N0543_v, N0543_port_8);
  spice_transistor_nmos_gnd tM1498(v(N0469_v), N0453_v, N0453_port_0);
  spice_transistor_nmos_vdd tM1493(v(SC_A22_M22_CLK2_v), N0869_v, N0869_port_10);
  spice_transistor_nmos tM1492(v(N0657_v), N0869_v, N0991_v, N0869_port_9, N0991_port_1);
  spice_transistor_nmos_gnd tM1491(v(R15_3_v), N0991_v, N0991_port_0);
  spice_transistor_nmos_gnd tM1497(v(N0461_v), ADDR_RFSH_1_v, ADDR_RFSH_1_port_1);
  spice_transistor_nmos_gnd tM1673(v(N0416_v), RADB0_v, RADB0_port_4);
  spice_transistor_nmos_gnd tM1672(v(N0711_v), N0307_v, N0307_port_3);
  spice_transistor_nmos_gnd tM2418(v(N0739_v), X32_v, X32_port_11);
  spice_transistor_nmos_gnd tM1670(v(N0317_v), N0732_v, N0732_port_1);
  spice_transistor_nmos_gnd tM1677(v(clk1_v), N0307_v, N0307_port_5);
  spice_transistor_nmos_gnd tM1675(v(clk2_v), N0300_v, N0300_port_3);
  spice_transistor_nmos_gnd tM2412(v(_OPA_1_v), DAA_v, DAA_port_4);
  spice_transistor_nmos_gnd tM2413(v(clk2_v), N0398_v, N0398_port_1);
  spice_transistor_nmos_gnd tM1679(v(N0717_v), N0737_v, N0737_port_2);
  spice_transistor_nmos_gnd tM2411(v(OPA_2_v), CLB_v, CLB_port_3);
  spice_transistor_nmos_vdd tM2416(v(S00690_v), N0741_v, N0741_port_1);
  spice_transistor_nmos tM1475(v(N0616_v), N0963_v, N0869_v, N0963_port_0, N0869_port_6);
  spice_transistor_nmos tM1474(v(N0591_v), N0869_v, N0954_v, N0869_port_5, N0954_port_1);
  spice_transistor_nmos tM1477(v(N0619_v), R11_3_v, N0538_v, R11_3_port_0, N0538_port_7);
  spice_transistor_nmos_gnd tM1476(v(R9_3_v), N0963_v, N0963_port_1);
  spice_transistor_nmos tM1471(v(N0619_v), R10_3_v, N0537_v, R10_3_port_1, N0537_port_7);
  spice_transistor_nmos tM1470(v(N0598_v), N0537_v, R8_3_v, N0537_port_6, R8_3_port_1);
  spice_transistor_nmos_gnd tM1473(v(R7_3_v), N0954_v, N0954_port_0);
  spice_transistor_nmos tM1472(v(N0598_v), N0538_v, R9_3_v, N0538_port_6, R9_3_port_0);
  spice_transistor_nmos tM2782(v(clk2_v), N0675_v, N0684_v, N0675_port_3, N0684_port_0);
  spice_transistor_nmos_gnd tM2783(v(N0685_v), N0684_v, N0684_port_1);
  spice_transistor_nmos tM2741(v(clk1_v), N0685_v, N0701_v, N0685_port_0, N0701_port_2);
  spice_transistor_nmos tM1479(v(N0634_v), N0537_v, R12_3_v, N0537_port_8, R12_3_port_1);
  spice_transistor_nmos_gnd tM1478(v(R11_3_v), N0973_v, N0973_port_0);
  spice_transistor_nmos_gnd tM2784(v(N0707_v), N0705_v, N0705_port_0);
  spice_transistor_nmos tM2785(v(L_v), N0705_v, N0706_v, N0705_port_1, N0706_port_0);
  spice_transistor_nmos_gnd tM2899(v(DCL_0_v), N0751_v, N0751_port_1);
  spice_transistor_nmos_vdd tM2893(v(N0911_v), N0553_v, N0553_port_2);
  spice_transistor_nmos_gnd tM2890(v(N0604_v), N0939_v, N0939_port_3);
  spice_transistor_nmos_gnd tM2078(v(_OPR_3_v), N0628_v, N0628_port_0);
  spice_transistor_nmos tM2079(v(_OPR_3_v), INC_ISZ_XCH_v, N0587_v, INC_ISZ_XCH_port_1, N0587_port_0);
  spice_transistor_nmos tM1781(v(SC_M22_CLK2_v), D2_v, N0617_v, D2_port_7, N0617_port_1);
  spice_transistor_nmos tM1780(v(SC_M22_CLK2_v), D1_v, N0582_v, D1_port_7, N0582_port_1);
  spice_transistor_nmos_gnd tM2074(v(SC_v), N0681_v, N0681_port_1);
  spice_transistor_nmos_gnd tM2075(v(X12_v), N0629_v, N0629_port_0);
  spice_transistor_nmos_gnd tM2076(v(_OPR_3_v), XCH_v, XCH_port_0);
  spice_transistor_nmos_gnd tM2077(v(_OPR_3_v), BBL_v, BBL_port_1);
  spice_transistor_nmos tM2070(v(M22_v), N0679_v, N0680_v, N0679_port_2, N0680_port_0);
  spice_transistor_nmos_gnd tM2071(v(N0643_v), SC_A22_v, SC_A22_port_4);
  spice_transistor_nmos tM2072(v(clk2_v), N0703_v, N0682_v, N0703_port_0, N0682_port_1);
  spice_transistor_nmos tM2073(v(clk2_v), N0681_v, N0680_v, N0681_port_0, N0680_port_1);
  spice_transistor_nmos_gnd tM2254(v(OPE_v), _OPE_v, _OPE_port_1);
  spice_transistor_nmos_gnd tM2527(v(POC_v), N0328_v, N0328_port_2);
  spice_transistor_nmos_gnd tM2524(v(clk2_v), N0337_v, N0337_port_2);
  spice_transistor_nmos_gnd tM2525(v(N0337_v), __X21__CLK2__v, __X21__CLK2__port_3);
  spice_transistor_nmos_gnd tM2250(v(IO_v), _I_O_v, _I_O_port_0);
  spice_transistor_nmos_vdd tM2251(v(N0493_v), _I_O_v, _I_O_port_1);
  spice_transistor_nmos_gnd tM2252(v(ISZ_v), N0456_v, N0456_port_0);
  spice_transistor_nmos_gnd tM2253(v(JCN_v), N0476_v, N0476_port_0);
  spice_transistor_nmos_gnd tM3305(v(d3_v), N0664_v, N0664_port_4);
  spice_transistor_nmos_gnd tM3304(v(N0676_v), N0663_v, N0663_port_3);
  spice_transistor_nmos_gnd tM3307(v(POC_v), d1_v, d1_port_4);
  spice_transistor_nmos_gnd tM3306(v(vss_v), d3_v, d3_port_4);
  spice_transistor_nmos_vdd tM3300(v(S00840_v), N0695_v, N0695_port_3);
  spice_transistor_nmos tM2528(v(X22_v), N0330_v, N0331_v, N0330_port_0, N0331_port_0);
  spice_transistor_nmos_gnd tM2529(v(clk2_v), N0330_v, N0330_port_1);
  spice_transistor_nmos_gnd tM2096(v(_OPR_2_v), IO_v, IO_port_1);
  spice_transistor_nmos_gnd tM2097(v(_OPR_2_v), OPE_v, OPE_port_1);
  spice_transistor_nmos_gnd tM2094(v(OPR_3_v), INC_ISZ_v, INC_ISZ_port_1);
  spice_transistor_nmos_gnd tM2095(v(_OPR_2_v), ISZ_v, ISZ_port_1);
  spice_transistor_nmos_gnd tM2092(v(OPR_3_v), JIN_FIN_v, JIN_FIN_port_4);
  spice_transistor_nmos_gnd tM2093(v(OPR_3_v), JUN_JMS_v, JUN_JMS_port_4);
  spice_transistor_nmos_gnd tM2091(v(OPR_3_v), FIM_SRC_v, FIM_SRC_port_0);
  spice_transistor_nmos_vdd tM2892(v(S00762_v), N0939_v, N0939_port_4);
  spice_transistor_nmos tM2320(v(N0297_v), N0295_v, N0296_v, N0295_port_1, N0296_port_0);
  spice_transistor_nmos_gnd tM2321(v(N0280_v), N0296_v, N0296_port_1);
  spice_transistor_nmos tM2323(v(clk1_v), N0739_v, N0296_v, N0739_port_0, N0296_port_3);
  spice_transistor_nmos tM2324(v(clk1_v), N0404_v, N0397_v, N0404_port_0, N0397_port_2);
  spice_transistor_nmos_gnd tM2325(v(N0405_v), N0404_v, N0404_port_1);
  spice_transistor_nmos tM2326(v(clk2_v), N0413_v, N0405_v, N0413_port_2, N0405_port_1);
  spice_transistor_nmos_gnd tM3230(v(N0607_v), N0945_v, N0945_port_3);
  spice_transistor_nmos_gnd tM3233(v(N0403_v), N0357_v, N0357_port_5);
  spice_transistor_nmos_gnd tM2539(v(INC_ISZ_v), N0442_v, N0442_port_0);
  spice_transistor_nmos_gnd tM3124(v(N0287_v), N0730_v, N0730_port_1);
  spice_transistor_nmos_gnd tM3127(v(_COM_v), N0714_v, N0714_port_1);
  spice_transistor_nmos tM3126(v(clk2_v), N0287_v, N0288_v, N0287_port_1, N0288_port_7);
  spice_transistor_nmos tM3123(v(clk1_v), N0731_v, N0730_v, N0731_port_2, N0730_port_0);
  spice_transistor_nmos_gnd tM3122(v(N0749_v), N0714_v, N0714_port_0);
  spice_transistor_nmos_gnd tM2963(v(A22_v), N0288_v, N0288_port_5);
  spice_transistor_nmos_vdd tM3129(v(S00818_v), N0714_v, N0714_port_2);
  spice_transistor_nmos_gnd tM2739(v(ADD_GROUP_4__v), CY_ADA_v, CY_ADA_port_0);
  spice_transistor_nmos_vdd tM2631(v(S00709_v), SUB_GROUP_6__v, SUB_GROUP_6__port_1);
  spice_transistor_nmos_gnd tM2636(v(__X31__CLK2__v), ADSL_v, ADSL_port_0);
  spice_transistor_nmos tM2968(v(N0937_v), TMP_1_v, N0889_v, TMP_1_port_0, N0889_port_4);
  spice_transistor_nmos_gnd tM2981(v(N0912_v), N0916_v, N0916_port_0);
  spice_transistor_nmos tM1978(v(X12_v), N0595_v, N0594_v, N0595_port_0, N0594_port_1);
  spice_transistor_nmos_gnd tM1979(v(BBL_v), N0468_v, N0468_port_0);
  spice_transistor_nmos_gnd tM2635(v(RAR_v), N0490_v, N0490_port_0);
  spice_transistor_nmos_gnd tM2969(v(N0942_v), _TMP_1_v, _TMP_1_port_0);
  spice_transistor_nmos_vdd tM2639(v(S00729_v), ADD_IB_v, ADD_IB_port_2);
  spice_transistor_nmos_gnd tM2737(v(N0342_v), N0546_v, N0546_port_2);
  spice_transistor_nmos_gnd tM2445(v(clk2_v), N0375_v, N0375_port_0);
  spice_transistor_nmos_gnd tM2444(v(N0797_v), N0782_v, N0782_port_4);
  spice_transistor_nmos tM1974(v(clk2_v), N0608_v, N0615_v, N0608_port_1, N0615_port_1);
  spice_transistor_nmos_gnd tM3038(v(N0879_v), N0876_v, N0876_port_1);
  spice_transistor_nmos_gnd tM1975(v(X22_v), N0589_v, N0589_port_0);
  spice_transistor_nmos_gnd tM2446(v(N0408_v), N0797_v, N0797_port_1);
  spice_transistor_nmos_vdd tM2967(v(S00767_v), N0912_v, N0912_port_2);
  spice_transistor_nmos_gnd tM2441(v(N0329_v), N0800_v, N0800_port_1);
  spice_transistor_nmos_gnd tM2442(v(N0805_v), N0798_v, N0798_port_0);
  spice_transistor_nmos_gnd tM2562(v(N0332_v), N0340_v, N0340_port_2);
  spice_transistor_nmos_gnd tM2964(v(N0765_v), DCL_1_v, DCL_1_port_1);
  spice_transistor_nmos_vdd tM2563(v(S00731_v), N0332_v, N0332_port_5);
  spice_transistor_nmos tM2560(v(clk2_v), M12_v, N0433_v, M12_port_8, N0433_port_0);
  spice_transistor_nmos tM2293(v(SC_M12_CLK2_v), D3_v, N1008_v, D3_port_8, N1008_port_1);
  spice_transistor_nmos_gnd tM2962(v(N0346_v), N0363_v, N0363_port_2);
  spice_transistor_nmos_gnd tM2526(v(N0329_v), N0328_v, N0328_port_1);
  spice_transistor_nmos_gnd tM1268(v(R15_0_v), N0984_v, N0984_port_0);
  spice_transistor_nmos tM1269(v(N0657_v), N0866_v, N0984_v, N0866_port_9, N0984_port_1);
  spice_transistor_nmos tM1723(v(clk2_v), N0402_v, N0416_v, N0402_port_2, N0416_port_1);
  spice_transistor_nmos_gnd tM1260(v(R4_0_v), N0930_v, N0930_port_1);
  spice_transistor_nmos tM1262(v(N0529_v), N0533_v, R0_1_v, N0533_port_2, R0_1_port_1);
  spice_transistor_nmos tM1263(v(N0583_v), R6_0_v, N0532_v, R6_0_port_0, N0532_port_5);
  spice_transistor_nmos_gnd tM1264(v(R6_0_v), N0948_v, N0948_port_0);
  spice_transistor_nmos_vdd tM1379(v(N0325_v), N0306_v, N0306_port_1);
  spice_transistor_nmos_vdd tM1318(v(SC_A22_M22_CLK2_v), N0880_v, N0880_port_10);
  spice_transistor_nmos_gnd tM1319(v(R14_1_v), N0986_v, N0986_port_0);
  spice_transistor_nmos_vdd tM1315(v(SC_A22_M22_CLK2_v), N0866_v, N0866_port_10);
  spice_transistor_nmos tM1645(v(clk1_v), N0503_v, N0504_v, N0503_port_2, N0504_port_0);
  spice_transistor_nmos tM1310(v(N0581_v), N0932_v, N0867_v, N0932_port_0, N0867_port_4);
  spice_transistor_nmos tM1312(v(N0598_v), N0533_v, R8_1_v, N0533_port_6, R8_1_port_1);
  spice_transistor_nmos tM1313(v(N0645_v), N0977_v, N0881_v, N0977_port_0, N0881_port_8);
  spice_transistor_nmos_gnd tM2667(v(ADD_v), ADD_GROUP_4__v, ADD_GROUP_4__port_4);
  spice_transistor_nmos_gnd tM2666(v(ADD_v), READ_ACC_3__v, READ_ACC_3__port_9);
  spice_transistor_nmos_gnd tM2661(v(SBM_v), SUB_GROUP_6__v, SUB_GROUP_6__port_2);
  spice_transistor_nmos_gnd tM2660(v(ADM_v), ADD_GROUP_4__v, ADD_GROUP_4__port_2);
  spice_transistor_nmos_gnd tM2594(v(DAC_v), WRITE_ACC_1__v, WRITE_ACC_1__port_7);
  spice_transistor_nmos_gnd tM2450(v(X22_v), N0288_v, N0288_port_0);
  spice_transistor_nmos_gnd tM2409(v(OPA_2_v), IAC_v, IAC_port_3);
  spice_transistor_nmos_gnd tM2408(v(OPA_2_v), DAC_v, DAC_port_3);
  spice_transistor_nmos_gnd tM2098(v(_OPR_2_v), JUN_JMS_v, JUN_JMS_port_5);
  spice_transistor_nmos_gnd tM1689(v(clk2_v), RADB1_v, RADB1_port_5);
  spice_transistor_nmos_gnd tM1686(v(X32_v), N0402_v, N0402_port_1);
  spice_transistor_nmos_gnd tM2400(v(OPA_2_v), TCS_v, TCS_port_3);
  spice_transistor_nmos_gnd tM1684(v(N0708_v), N0710_v, N0710_port_1);
  spice_transistor_nmos_gnd tM2402(v(N1003_v), _OPA_2_v, _OPA_2_port_6);
  spice_transistor_nmos_vdd tM2405(v(N1001_v), OPA_3_v, OPA_3_port_13);
  spice_transistor_nmos_vdd tM2404(v(N1000_v), _OPA_3_v, _OPA_3_port_11);
  spice_transistor_nmos_vdd tM1680(v(N0710_v), M12_M22_CLK1__M11_M12__v, M12_M22_CLK1__M11_M12__port_8);
  spice_transistor_nmos_gnd tM1681(v(N0708_v), M12_M22_CLK1__M11_M12__v, M12_M22_CLK1__M11_M12__port_9);
  spice_transistor_nmos tM1442(v(N0569_v), N0537_v, R4_3_v, N0537_port_4, R4_3_port_1);
  spice_transistor_nmos tM1443(v(N0591_v), N0883_v, N0953_v, N0883_port_5, N0953_port_1);
  spice_transistor_nmos tM1444(v(N0616_v), N0962_v, N0883_v, N0962_port_0, N0883_port_6);
  spice_transistor_nmos_gnd tM1445(v(R8_3_v), N0962_v, N0962_port_1);
  spice_transistor_nmos_gnd tM1446(v(R12_2_v), N0980_v, N0980_port_1);
  spice_transistor_nmos_gnd tM1447(v(R10_3_v), N0972_v, N0972_port_0);
  spice_transistor_nmos tM1448(v(N0583_v), R6_3_v, N0537_v, R6_3_port_1, N0537_port_5);
  spice_transistor_nmos tM1449(v(N0569_v), N0538_v, R5_3_v, N0538_port_4, R5_3_port_0);
  spice_transistor_nmos_vdd tM2598(v(N1004_v), _OPA_1_v, _OPA_1_port_8);
  spice_transistor_nmos tM2794(v(N0854_v), N0855_v, N0452_v, N0855_port_3, N0452_port_1);
  spice_transistor_nmos_gnd tM2797(v(M12_v), N0937_v, N0937_port_1);
  spice_transistor_nmos_gnd tM2849(v(N0346_v), ACC_0_v, ACC_0_port_1);
  spice_transistor_nmos tM2889(v(N0964_v), D0_v, N0604_v, D0_port_14, N0604_port_1);
  spice_transistor_nmos_gnd tM2888(v(N0915_v), N0553_v, N0553_port_1);
  spice_transistor_nmos tM2848(v(N0378_v), N0377_v, N0376_v, N0377_port_0, N0376_port_0);
  spice_transistor_nmos_vdd tM2885(v(N0940_v), TMP_0_v, TMP_0_port_1);
  spice_transistor_nmos_vdd tM2887(v(M12_v), N0604_v, N0604_port_0);
  spice_transistor_nmos_gnd tM2886(v(N0939_v), TMP_0_v, TMP_0_port_2);
  spice_transistor_nmos tM2880(v(ADD_IB_v), D0_v, N0846_v, D0_port_13, N0846_port_5);
  spice_transistor_nmos_gnd tM2883(v(N0939_v), N0940_v, N0940_port_2);
  spice_transistor_nmos_gnd tM1045(v(N0291_v), N0757_v, N0757_port_1);
  spice_transistor_nmos tM1046(v(N0291_v), N0298_v, N0299_v, N0298_port_3, N0299_port_0);
  spice_transistor_nmos tM1047(v(N0291_v), N0312_v, N0313_v, N0312_port_1, N0313_port_0);
  spice_transistor_nmos_gnd tM1040(v(N0293_v), N0758_v, N0758_port_1);
  spice_transistor_nmos tM1041(v(N0293_v), N0763_v, N0757_v, N0763_port_1, N0757_port_0);
  spice_transistor_nmos_gnd tM1043(v(N0291_v), N0758_v, N0758_port_3);
  spice_transistor_nmos_gnd tM2062(v(POC_v), N0683_v, N0683_port_1);
  spice_transistor_nmos tM2061(v(SC_v), N0618_v, N0623_v, N0618_port_2, N0623_port_1);
  spice_transistor_nmos tM1048(v(N0291_v), N0302_v, N0303_v, N0302_port_1, N0303_port_0);
  spice_transistor_nmos_vdd tM1049(v(N0325_v), N0293_v, N0293_port_2);
  spice_transistor_nmos_vdd tM2064(v(N0626_v), __POC__CLK2_SC_A32_X12__v, __POC__CLK2_SC_A32_X12__port_9);
  spice_transistor_nmos_gnd tM2243(v(N0327_v), POC_v, POC_port_4);
  spice_transistor_nmos_gnd tM2242(v(N0327_v), N0769_v, N0769_port_2);
  spice_transistor_nmos_gnd tM2241(v(N0397_v), _CN_v, _CN_port_3);
  spice_transistor_nmos_gnd tM2240(v(reset_v), N0327_v, N0327_port_0);
  spice_transistor_nmos_gnd tM2247(v(IO_v), N0493_v, N0493_port_1);
  spice_transistor_nmos tM2246(v(X32_v), N0417_v, N0418_v, N0417_port_1, N0418_port_0);
  spice_transistor_nmos_gnd tM2245(v(X32_v), N0399_v, N0399_port_0);
  spice_transistor_nmos_gnd tM2244(v(N0397_v), N0412_v, N0412_port_0);
  spice_transistor_nmos_vdd tM2249(v(N0510_v), _OPE_v, _OPE_port_0);
  spice_transistor_nmos_gnd tM2248(v(OPE_v), N0510_v, N0510_port_1);
  spice_transistor_nmos_gnd tM2081(v(_OPR_3_v), SUB_v, SUB_port_0);
  spice_transistor_nmos_gnd tM2080(v(_OPR_3_v), LD_v, LD_port_0);
  spice_transistor_nmos_gnd tM2083(v(OPR_3_v), JCN_ISZ_v, JCN_ISZ_port_3);
  spice_transistor_nmos_gnd tM2082(v(_OPR_3_v), ADD_v, ADD_port_0);
  spice_transistor_nmos_gnd tM2089(v(N0343_v), N0344_v, N0344_port_2);
  spice_transistor_nmos_gnd tM2088(v(N0343_v), SC_v, SC_port_13);
  spice_transistor_nmos_gnd tM2993(v(N0605_v), N0941_v, N0941_port_3);
  spice_transistor_nmos_gnd tM2183(v(N0992_v), OPR_3_v, OPR_3_port_15);
  spice_transistor_nmos tM3204(v(N0559_v), N0557_v, N0558_v, N0557_port_2, N0558_port_2);
  spice_transistor_nmos tM3200(v(ACC_ADA_v), N0873_v, N0859_v, N0873_port_5, N0859_port_4);
  spice_transistor_nmos tM3201(v(N0873_v), N0558_v, N0914_v, N0558_port_1, N0914_port_1);
  spice_transistor_nmos_gnd tM3202(v(N0559_v), N0901_v, N0901_port_2);
  spice_transistor_nmos_gnd tM3203(v(N0893_v), N0901_v, N0901_port_3);
  spice_transistor_nmos_gnd tM3208(v(N0666_v), D2_v, D2_port_17);
  spice_transistor_nmos_vdd tM3209(v(N0665_v), D2_v, D2_port_18);
  spice_transistor_nmos_gnd tM2992(v(N0700_v), N0692_v, N0692_port_1);
  spice_transistor_nmos_gnd tM2339(v(_OPE_v), O_IB_v, O_IB_port_1);
  spice_transistor_nmos_gnd tM2338(v(_OPE_v), DCL_v, DCL_port_1);
  spice_transistor_nmos_gnd tM2337(v(N0476_v), N0478_v, N0478_port_0);
  spice_transistor_nmos_gnd tM2333(v(N0739_v), N0741_v, N0741_port_0);
  spice_transistor_nmos_gnd tM2361(v(_OPE_v), STC_v, STC_port_1);
  spice_transistor_nmos tM2456(v(clk2_v), N0281_v, X12_v, N0281_port_1, X12_port_10);
  spice_transistor_nmos tM3110(v(ADD_IB_v), N0514_v, D3_v, N0514_port_2, D3_port_13);
  spice_transistor_nmos_vdd tM3112(v(N0877_v), N0514_v, N0514_port_3);
  spice_transistor_nmos tM3113(v(ACB_IB_v), D3_v, N0356_v, D3_port_14, N0356_port_6);
  spice_transistor_nmos tM3114(v(ACC_ADAC_v), N0873_v, N0474_v, N0873_port_0, N0474_port_0);
  spice_transistor_nmos_gnd tM3115(v(N0377_v), N0358_v, N0358_port_0);
  spice_transistor_nmos_gnd tM3116(v(N0345_v), N0358_v, N0358_port_1);
  spice_transistor_nmos_gnd tM3118(v(N0363_v), N0358_v, N0358_port_3);
  spice_transistor_nmos_gnd tM3119(v(N0370_v), N0358_v, N0358_port_4);
  spice_transistor_nmos tM2209(v(_OPR_0_v), INC_ISZ_XCH_v, N0587_v, INC_ISZ_XCH_port_4, N0587_port_6);
  spice_transistor_nmos_gnd tM2659(v(ADM_v), READ_ACC_3__v, READ_ACC_3__port_7);
  spice_transistor_nmos_gnd tM2208(v(OPR_1_v), JUN2_JMS2_v, JUN2_JMS2_port_2);
  spice_transistor_nmos_gnd tM2207(v(_OPR_0_v), JMS_v, JMS_port_4);
  spice_transistor_nmos_gnd tM1110(v(N0866_v), N0531_v, N0531_port_0);
  spice_transistor_nmos tM1116(v(N0434_v), N0823_v, N0778_v, N0823_port_1, N0778_port_4);
  spice_transistor_nmos_gnd tM1114(v(PC2_3_v), N0823_v, N0823_port_0);
  spice_transistor_nmos_gnd tM2451(v(N0719_v), N0742_v, N0742_port_1);
  spice_transistor_nmos_gnd tM1871(v(X12_v), N0447_v, N0447_port_1);
  spice_transistor_nmos_gnd tM1872(v(X32_v), N0447_v, N0447_port_2);
  spice_transistor_nmos_gnd tM1875(v(clk1_v), N0443_v, N0443_port_2);
  spice_transistor_nmos tM1879(v(clk2_v), N0517_v, N0511_v, N0517_port_1, N0511_port_1);
  spice_transistor_nmos_gnd tM2875(v(N0870_v), N0898_v, N0898_port_1);
  spice_transistor_nmos_gnd tM2957(v(N0553_v), N0899_v, N0899_port_2);
  spice_transistor_nmos tM2956(v(N0556_v), N0899_v, N0875_v, N0899_port_1, N0875_port_4);
  spice_transistor_nmos_vdd tM2954(v(M12_v), N0871_v, N0871_port_5);
  spice_transistor_nmos_gnd tM2960(v(N0346_v), N0345_v, N0345_port_2);
  spice_transistor_nmos tM1309(v(N0565_v), N0867_v, N0923_v, N0867_port_3, N0923_port_1);
  spice_transistor_nmos tM1308(v(N0543_v), N0907_v, N0868_v, N0907_port_1, N0868_port_2);
  spice_transistor_nmos tM1303(v(N0569_v), N0534_v, R5_1_v, N0534_port_4, R5_1_port_0);
  spice_transistor_nmos tM1302(v(N0583_v), R6_1_v, N0533_v, R6_1_port_1, N0533_port_5);
  spice_transistor_nmos tM1301(v(N0657_v), N0880_v, N0985_v, N0880_port_9, N0985_port_1);
  spice_transistor_nmos_gnd tM1300(v(R14_0_v), N0985_v, N0985_port_0);
  spice_transistor_nmos_gnd tM1307(v(N0868_v), N0535_v, N0535_port_1);
  spice_transistor_nmos_gnd tM1306(v(R1_2_v), N0907_v, N0907_port_0);
  spice_transistor_nmos_gnd tM1305(v(R3_1_v), N0923_v, N0923_port_0);
  spice_transistor_nmos tM1304(v(N0583_v), R7_1_v, N0534_v, R7_1_port_0, N0534_port_5);
  spice_transistor_nmos_gnd tM2654(v(N0515_v), ACC_ADAC_v, ACC_ADAC_port_0);
  spice_transistor_nmos_gnd tM2655(v(N0342_v), ACC_ADAC_v, ACC_ADAC_port_1);
  spice_transistor_nmos tM1276(v(N0616_v), N0957_v, N0880_v, N0957_port_1, N0880_port_6);
  spice_transistor_nmos tM1275(v(N0619_v), R10_0_v, N0532_v, R10_0_port_0, N0532_port_7);
  spice_transistor_nmos_gnd tM1277(v(R4_1_v), N0931_v, N0931_port_0);
  spice_transistor_nmos_gnd tM1274(v(R8_0_v), N0957_v, N0957_port_0);
  spice_transistor_nmos tM1273(v(N0598_v), N0532_v, R8_0_v, N0532_port_6, R8_0_port_0);
  spice_transistor_nmos tM1279(v(N0581_v), N0931_v, N0881_v, N0931_port_1, N0881_port_4);
  spice_transistor_nmos tM1278(v(N0565_v), N0881_v, N0922_v, N0881_port_3, N0922_port_1);
  spice_transistor_nmos_gnd tM1699(v(N0560_v), N0620_v, N0620_port_5);
  spice_transistor_nmos_gnd tM1698(v(N0560_v), N0584_v, N0584_port_5);
  spice_transistor_nmos_gnd tM3082(v(N0943_v), TMP_2_v, TMP_2_port_1);
  spice_transistor_nmos_gnd tM1697(v(N0560_v), N0545_v, N0545_port_5);
  spice_transistor_nmos tM1270(v(N0591_v), N0880_v, N0948_v, N0880_port_5, N0948_port_1);
  spice_transistor_nmos_gnd tM1691(v(clk2_v), RADB2_v, RADB2_port_5);
  spice_transistor_nmos_gnd tM1690(v(N0384_v), RADB1_v, RADB1_port_6);
  spice_transistor_nmos_gnd tM1692(v(N0374_v), RADB2_v, RADB2_port_6);
  spice_transistor_nmos tM1459(v(N0632_v), N0883_v, N0972_v, N0883_port_7, N0972_port_1);
  spice_transistor_nmos tM1458(v(N0583_v), R7_3_v, N0538_v, R7_3_port_0, N0538_port_5);
  spice_transistor_nmos_gnd tM1457(v(R5_3_v), N0936_v, N0936_port_1);
  spice_transistor_nmos tM1456(v(N0581_v), N0936_v, N0869_v, N0936_port_0, N0869_port_4);
  spice_transistor_nmos tM1455(v(N0565_v), N0869_v, N0927_v, N0869_port_3, N0927_port_1);
  spice_transistor_nmos_gnd tM1454(v(R3_3_v), N0927_v, N0927_port_0);
  spice_transistor_nmos_gnd tM1453(v(N0469_v), N0461_v, N0461_port_1);
  spice_transistor_nmos_gnd tM1451(v(N0461_v), N0469_v, N0469_port_0);
  spice_transistor_nmos_vdd tM3241(v(S00828_v), N0854_v, N0854_port_6);
  spice_transistor_nmos tM1053(v(WADB0_v), N0779_v, N0762_v, N0779_port_0, N0762_port_3);
  spice_transistor_nmos tM1052(v(WADB0_v), N0778_v, N0761_v, N0778_port_0, N0761_port_5);
  spice_transistor_nmos tM1051(v(WADB1_v), N0761_v, N0774_v, N0761_port_4, N0774_port_0);
  spice_transistor_nmos tM1050(v(M12_M22_CLK1__M11_M12__v), N0291_v, D1_v, N0291_port_5, D1_port_0);
  spice_transistor_nmos tM1057(v(RADB1_v), D1_v, N0392_v, D1_port_1, N0392_port_0);
  spice_transistor_nmos tM1056(v(RADB2_v), N0390_v, D2_v, N0390_port_0, D2_port_3);
  spice_transistor_nmos tM1055(v(RADB1_v), D2_v, N0389_v, D2_port_2, N0389_port_0);
  spice_transistor_nmos tM1054(v(WADB1_v), N0762_v, N0775_v, N0762_port_4, N0775_port_0);
  spice_transistor_nmos tM1059(v(RADB0_v), N0393_v, D1_v, N0393_port_0, D1_port_3);
  spice_transistor_nmos tM1058(v(RADB2_v), N0391_v, D1_v, N0391_port_0, D1_port_2);
  spice_transistor_nmos_gnd tM2500(v(_OPE_v), N0415_v, N0415_port_1);
  spice_transistor_nmos_vdd tM1026(v(S00531_v), N0740_v, N0740_port_1);
  spice_transistor_nmos_gnd tM2502(v(__X21__CLK2__v), N0351_v, N0351_port_1);
  spice_transistor_nmos_gnd tM2503(v(DCL_v), N0353_v, N0353_port_1);
  spice_transistor_nmos_gnd tM2504(v(KBP_v), WRITE_ACC_1__v, WRITE_ACC_1__port_0);
  spice_transistor_nmos_gnd tM2505(v(__X21__CLK2__v), N0415_v, N0415_port_2);
  spice_transistor_nmos_gnd tM2507(v(N0380_v), N0375_v, N0375_port_1);
  spice_transistor_nmos_gnd tM3248(v(D0_v), N0674_v, N0674_port_0);
  spice_transistor_nmos_gnd tM3160(v(_COM_v), N0716_v, N0716_port_3);
  spice_transistor_nmos_gnd tM1022(v(N0290_v), N0755_v, N0755_port_0);
  spice_transistor_nmos tM2008(v(_OPA_0_v), N0602_v, N0614_v, N0602_port_1, N0614_port_0);
  spice_transistor_nmos_gnd tM1752(v(N0492_v), N0491_v, N0491_port_0);
  spice_transistor_nmos_gnd tM3165(v(N0377_v), N0359_v, N0359_port_3);
  spice_transistor_nmos_gnd tM3164(v(N0370_v), N0359_v, N0359_port_2);
  spice_transistor_nmos_gnd tM2435(v(OPA_2_v), SBM_v, SBM_port_3);
  spice_transistor_nmos_gnd tM2436(v(OPA_2_v), ADM_v, ADM_port_3);
  spice_transistor_nmos_gnd tM2437(v(_OPA_1_v), ADM_v, ADM_port_4);
  spice_transistor_nmos_gnd tM2430(v(_OPA_1_v), TCC_v, TCC_port_4);
  spice_transistor_nmos_gnd tM2431(v(OPA_1_v), N0507_v, N0507_port_1);
  spice_transistor_nmos_gnd tM2432(v(_OPA_1_v), STC_v, STC_port_4);
  spice_transistor_nmos tM3166(v(N0415_v), D2_v, N0366_v, D2_port_16, N0366_port_6);
  spice_transistor_nmos_vdd tM2438(v(N0782_v), _COM_v, _COM_port_0);
  spice_transistor_nmos_gnd tM2439(v(N0784_v), _COM_v, _COM_port_1);
  spice_transistor_nmos_gnd tM3213(v(d2_v), N0666_v, N0666_port_3);
  spice_transistor_nmos_gnd tM3212(v(N0946_v), _TMP_3_v, _TMP_3_port_0);
  spice_transistor_nmos_gnd tM1696(v(N0409_v), N0400_v, N0400_port_0);
  spice_transistor_nmos_gnd tM3217(v(N0914_v), N0918_v, N0918_port_0);
  spice_transistor_nmos_vdd tM3216(v(N0945_v), _TMP_3_v, _TMP_3_port_2);
  spice_transistor_nmos_gnd tM3215(v(N0676_v), N0666_v, N0666_port_4);
  spice_transistor_nmos tM3214(v(SUB_GROUP_6__v), _TMP_3_v, N0893_v, _TMP_3_port_1, N0893_port_4);
  spice_transistor_nmos_gnd tM2001(v(N0622_v), CLK2_SC_A12_M12__v, CLK2_SC_A12_M12__port_8);
  spice_transistor_nmos_gnd tM3219(v(N0918_v), N0861_v, N0861_port_2);
  spice_transistor_nmos tM2348(v(N0456_v), N0478_v, N0419_v, N0478_port_3, N0419_port_1);
  spice_transistor_nmos_gnd tM2342(v(_OPE_v), DAA_v, DAA_port_1);
  spice_transistor_nmos_gnd tM2343(v(_OPE_v), RAR_v, RAR_port_1);
  spice_transistor_nmos_gnd tM2340(v(_OPE_v), KBP_v, KBP_port_1);
  spice_transistor_nmos_gnd tM2002(v(N0626_v), N0627_v, N0627_port_0);
  spice_transistor_nmos tM2346(v(N0487_v), N0478_v, N0481_v, N0478_port_1, N0481_port_0);
  spice_transistor_nmos tM2347(v(_OPA_3_v), N0478_v, N0481_v, N0478_port_2, N0481_port_1);
  spice_transistor_nmos_gnd tM2344(v(_OPE_v), RAL_v, RAL_port_1);
  spice_transistor_nmos_gnd tM2345(v(_OPE_v), CMA_v, CMA_port_1);
  spice_transistor_nmos_gnd tM2878(v(N0911_v), N0915_v, N0915_port_0);
  spice_transistor_nmos tM1590(v(N0648_v), N0647_v, CLK2_SC_A12_M12__v, N0647_port_9, CLK2_SC_A12_M12__port_7);
  spice_transistor_nmos_vdd tM3109(v(S00814_v), N0748_v, N0748_port_2);
  spice_transistor_nmos_gnd tM3108(v(N0356_v), N0376_v, N0376_port_5);
  spice_transistor_nmos_gnd tM3107(v(N0356_v), N0370_v, N0370_port_5);
  spice_transistor_nmos_gnd tM3106(v(N0356_v), N0363_v, N0363_port_5);
  spice_transistor_nmos_gnd tM3105(v(N0514_v), ADD_0_v, ADD_0_port_5);
  spice_transistor_nmos_gnd tM3104(v(N0356_v), N0349_v, N0349_port_2);
  spice_transistor_nmos_gnd tM3103(v(N0356_v), N0354_v, N0354_port_5);
  spice_transistor_nmos_gnd tM3102(v(N0349_v), N0345_v, N0345_port_5);
  spice_transistor_nmos tM3101(v(N0766_v), N0768_v, N0749_v, N0768_port_2, N0749_port_2);
  spice_transistor_nmos_gnd tM2983(v(N0941_v), N0942_v, N0942_port_2);
  spice_transistor_nmos_gnd tM1848(v(N0451_v), N0449_v, N0449_port_6);
  spice_transistor_nmos_gnd tM1849(v(JIN_FIN_v), N0441_v, N0441_port_1);
  spice_transistor_nmos_gnd tM1844(v(N0443_v), N0436_v, N0436_port_3);
  spice_transistor_nmos tM1845(v(N0435_v), N0436_v, N0441_v, N0436_port_4, N0441_port_0);
  spice_transistor_nmos_gnd tM1846(v(POC_v), N0449_v, N0449_port_4);
  spice_transistor_nmos_gnd tM1847(v(N0447_v), N0449_v, N0449_port_5);
  spice_transistor_nmos_gnd tM1840(v(INH_v), __INH__X11_X31_CLK1_v, __INH__X11_X31_CLK1_port_14);
  spice_transistor_nmos_gnd tM1841(v(N0522_v), __INH__X11_X31_CLK1_v, __INH__X11_X31_CLK1_port_15);
  spice_transistor_nmos_gnd tM1843(v(INH_v), N0449_v, N0449_port_3);
  spice_transistor_nmos_gnd tM2501(v(N0353_v), N0351_v, N0351_port_0);
  spice_transistor_nmos_gnd tM3012(v(N0347_v), N0370_v, N0370_port_3);
  spice_transistor_nmos_gnd tM1998(v(N0622_v), N0621_v, N0621_port_0);
  spice_transistor_nmos_gnd tM1997(v(N0653_v), N0652_v, N0652_port_1);
  spice_transistor_nmos tM1518(v(clk2_v), N0314_v, N0315_v, N0314_port_2, N0315_port_0);
  spice_transistor_nmos_vdd tM1519(v(N0717_v), cm_rom_v, cm_rom_port_0);
  spice_transistor_nmos_gnd tM1517(v(A32_v), N0712_v, N0712_port_0);
  spice_transistor_nmos tM1514(v(N0381_v), N0396_v, PC0_8_v, N0396_port_2, PC0_8_port_0);
  spice_transistor_nmos tM1515(v(N0406_v), N0796_v, N0773_v, N0796_port_0, N0773_port_2);
  spice_transistor_nmos tM1512(v(N0455_v), N0453_v, N0454_v, N0453_port_2, N0454_port_0);
  spice_transistor_nmos tM1513(v(N0410_v), PC1_4_v, N0395_v, PC1_4_port_1, N0395_port_3);
  spice_transistor_nmos_gnd tM1510(v(PC3_4_v), N0844_v, N0844_port_0);
  spice_transistor_nmos tM1511(v(N0455_v), ADDR_RFSH_1_v, N0489_v, ADDR_RFSH_1_port_2, N0489_port_0);
  spice_transistor_nmos tM2039(v(_OPA_0_v), N0567_v, N0562_v, N0567_port_0, N0562_port_2);
  spice_transistor_nmos_gnd tM1192(v(N0772_v), N0391_v, N0391_port_1);
  spice_transistor_nmos tM1193(v(WADB2_v), N0772_v, N0763_v, N0772_port_1, N0763_port_3);
  spice_transistor_nmos tM1191(v(N0439_v), PC3_10_v, N0390_v, PC3_10_port_0, N0390_port_5);
  spice_transistor_nmos_gnd tM1196(v(PC0_9_v), N0791_v, N0791_port_1);
  spice_transistor_nmos_gnd tM1197(v(PC1_10_v), N0811_v, N0811_port_0);
  spice_transistor_nmos tM1194(v(WADB1_v), N0763_v, N0776_v, N0763_port_4, N0776_port_0);
  spice_transistor_nmos tM1195(v(N0406_v), N0791_v, N0772_v, N0791_port_0, N0772_port_2);
  spice_transistor_nmos tM1198(v(N0424_v), N0771_v, N0811_v, N0771_port_3, N0811_port_1);
  spice_transistor_nmos tM1199(v(N0434_v), N0826_v, N0771_v, N0826_port_0, N0771_port_4);
  spice_transistor_nmos tM1202(v(M12_M22_CLK1__M11_M12__v), N0499_v, D2_v, N0499_port_0, D2_port_4);
  spice_transistor_nmos_gnd tM1208(v(PC2_9_v), N0827_v, N0827_port_0);
  spice_transistor_nmos tM1209(v(N0424_v), N0772_v, N0812_v, N0772_port_3, N0812_port_1);
  spice_transistor_nmos tM1394(v(N0444_v), N0781_v, N0843_v, N0781_port_5, N0843_port_1);
  spice_transistor_nmos tM1428(v(N0634_v), N0535_v, R13_2_v, N0535_port_8, R13_2_port_1);
  spice_transistor_nmos tM1429(v(N0647_v), R15_2_v, N0535_v, R15_2_port_1, N0535_port_9);
  spice_transistor_nmos tM2535(v(N0329_v), N0331_v, N0332_v, N0331_port_1, N0332_port_1);
  spice_transistor_nmos tM2130(v(OPR_2_v), N0523_v, JCN_ISZ_v, N0523_port_1, JCN_ISZ_port_5);
  spice_transistor_nmos_gnd tM1422(v(R4_3_v), N0935_v, N0935_port_1);
  spice_transistor_nmos_gnd tM1423(v(R6_2_v), N0952_v, N0952_port_0);
  spice_transistor_nmos tM1420(v(N0565_v), N0883_v, N0926_v, N0883_port_3, N0926_port_1);
  spice_transistor_nmos tM1421(v(N0581_v), N0935_v, N0883_v, N0935_port_0, N0883_port_4);
  spice_transistor_nmos_gnd tM1426(v(R8_2_v), N0961_v, N0961_port_1);
  spice_transistor_nmos tM1427(v(N0619_v), R10_2_v, N0536_v, R10_2_port_0, N0536_port_7);
  spice_transistor_nmos tM1424(v(N0591_v), N0882_v, N0952_v, N0882_port_5, N0952_port_1);
  spice_transistor_nmos tM1425(v(N0616_v), N0961_v, N0882_v, N0961_port_0, N0882_port_6);
  spice_transistor_nmos_gnd tM2647(v(CMA_v), N0515_v, N0515_port_0);
  spice_transistor_nmos_gnd tM2646(v(N0490_v), ADSR_v, ADSR_port_1);
  spice_transistor_nmos_gnd tM2645(v(__X31__CLK2__v), ADSR_v, ADSR_port_0);
  spice_transistor_nmos_gnd tM2642(v(N0502_v), ADSL_v, ADSL_port_1);
  spice_transistor_nmos_vdd tM2649(v(S00724_v), ACB_IB_v, ACB_IB_port_2);
  spice_transistor_nmos_gnd tM2519(v(N0282_v), N0720_v, N0720_port_0);
  spice_transistor_nmos_gnd tM2961(v(N0346_v), N0354_v, N0354_port_2);
  spice_transistor_nmos_gnd tM2514(v(N0375_v), __X31__CLK2__v, __X31__CLK2__port_2);
  spice_transistor_nmos_gnd tM2511(v(DAA_v), WRITE_ACC_1__v, WRITE_ACC_1__port_2);
  spice_transistor_nmos_gnd tM2510(v(TCS_v), WRITE_ACC_1__v, WRITE_ACC_1__port_1);
  spice_transistor_nmos tM1737(v(clk2_v), N0278_v, N0279_v, N0278_port_1, N0279_port_1);
  spice_transistor_nmos_gnd tM1734(v(M12_v), N0708_v, N0708_port_4);
  spice_transistor_nmos_gnd tM1735(v(M22_v), N0708_v, N0708_port_5);
  spice_transistor_nmos_gnd tM1732(v(N0278_v), N0709_v, N0709_port_1);
  spice_transistor_nmos tM1731(v(clk1_v), N0708_v, N0709_v, N0708_port_3, N0709_port_0);
  spice_transistor_nmos_gnd tM1738(v(M12_v), N0279_v, N0279_port_2);
  spice_transistor_nmos_gnd tM1739(v(clk2_v), RADB0_v, RADB0_port_6);
  spice_transistor_nmos_gnd tM2423(v(N0414_v), N0407_v, N0407_port_0);
  spice_transistor_nmos_gnd tM2422(v(_SRC_v), N0799_v, N0799_port_1);
  spice_transistor_nmos tM2421(v(clk2_v), N0414_v, A22_v, N0414_port_0, A22_port_5);
  spice_transistor_nmos_vdd tM2420(v(N0741_v), X32_v, X32_port_12);
  spice_transistor_nmos_vdd tM2426(v(S00685_v), N0415_v, N0415_port_0);
  spice_transistor_nmos tM2424(v(N0398_v), N0407_v, N0408_v, N0407_port_1, N0408_port_0);
  spice_transistor_nmos_gnd tM2429(v(_OPA_1_v), RAR_v, RAR_port_4);
  spice_transistor_nmos tM2428(v(CY_1_v), N0507_v, N0486_v, N0507_port_0, N0486_port_4);
  spice_transistor_nmos tM1236(v(N0434_v), N0828_v, N0776_v, N0828_port_0, N0776_port_4);
  spice_transistor_nmos_gnd tM2358(v(N0486_v), N0481_v, N0481_port_2);
  spice_transistor_nmos tM2351(v(ADD_0_v), N0478_v, N0419_v, N0478_port_4, N0419_port_2);
  spice_transistor_nmos_gnd tM2355(v(_OPA_3_v), KBP_v, KBP_port_2);
  spice_transistor_nmos_gnd tM2354(v(_OPA_3_v), DCL_v, DCL_port_2);
  spice_transistor_nmos_gnd tM2357(v(_OPA_3_v), DAA_v, DAA_port_2);
  spice_transistor_nmos_gnd tM2356(v(_OPA_3_v), TCS_v, TCS_port_2);
  spice_transistor_nmos_gnd tM2434(v(_OPA_1_v), IAC_v, IAC_port_4);
  spice_transistor_nmos tM2795(v(CY_ADAC_v), N0550_v, N0855_v, N0550_port_3, N0855_port_4);
  spice_transistor_nmos_gnd tM2433(v(_OPA_1_v), CMC_v, CMC_port_4);
  spice_transistor_nmos_gnd tM3172(v(N0345_v), N0357_v, N0357_port_1);
  spice_transistor_nmos_vdd tM3170(v(S00833_v), N0716_v, N0716_port_4);
  spice_transistor_nmos_vdd tM3171(v(S00834_v), N0713_v, N0713_port_2);
  spice_transistor_nmos tM3176(v(N0415_v), D0_v, N0357_v, D0_port_15, N0357_port_4);
  spice_transistor_nmos tM3177(v(M12_v), N0474_v, ACC_3_v, N0474_port_2, ACC_3_port_0);
  spice_transistor_nmos_gnd tM2822(v(DAA_v), N0802_v, N0802_port_1);
  spice_transistor_nmos_gnd tM2769(v(N0699_v), N0678_v, N0678_port_3);
  spice_transistor_nmos_gnd tM3006(v(N0347_v), N0345_v, N0345_port_3);
  spice_transistor_nmos_gnd tM3007(v(N0347_v), N0354_v, N0354_port_3);
  spice_transistor_nmos tM3004(v(N0351_v), N0364_v, N0765_v, N0364_port_1, N0765_port_1);
  spice_transistor_nmos_gnd tM3005(v(N0364_v), N0363_v, N0363_port_3);
  spice_transistor_nmos_gnd tM3002(v(POC_v), DCL_1_v, DCL_1_port_2);
  spice_transistor_nmos_vdd tM3000(v(N0747_v), A22_v, A22_port_8);
  spice_transistor_nmos_gnd tM3001(v(N0729_v), A22_v, A22_port_9);
  spice_transistor_nmos_gnd tM3008(v(N0347_v), N0364_v, N0364_port_3);
  spice_transistor_nmos tM3009(v(ACC_ADAC_v), N0872_v, N0858_v, N0872_port_0, N0858_port_1);
  spice_transistor_nmos tM1325(v(N0565_v), N0868_v, N0924_v, N0868_port_3, N0924_port_1);
  spice_transistor_nmos tM2998(v(N0854_v), N0858_v, N0851_v, N0858_port_0, N0851_port_1);
  spice_transistor_nmos_vdd tM3197(v(M12_v), N0873_v, N0873_port_4);
  spice_transistor_nmos tM2817(v(clk1_v), N0725_v, N0724_v, N0725_port_2, N0724_port_0);
  spice_transistor_nmos_gnd tM2349(v(_I_O_v), N0329_v, N0329_port_1);
  spice_transistor_nmos tM2781(v(clk1_v), L_v, N0707_v, L_port_5, N0707_port_0);
  spice_transistor_nmos_gnd tM1858(v(X32_v), N0334_v, N0334_port_1);
  spice_transistor_nmos_gnd tM1853(v(_CN_v), N0322_v, N0322_port_1);
  spice_transistor_nmos_gnd tM1852(v(clk2_v), N0451_v, N0451_port_2);
  spice_transistor_nmos_gnd tM1851(v(A22_v), N0318_v, N0318_port_5);
  spice_transistor_nmos_gnd tM1850(v(N0438_v), N0436_v, N0436_port_5);
  spice_transistor_nmos tM1857(v(JIN_FIN_v), N0334_v, N0333_v, N0334_port_0, N0333_port_1);
  spice_transistor_nmos_gnd tM1856(v(A12_v), N0326_v, N0326_port_2);
  spice_transistor_nmos tM1855(v(SC_v), N0333_v, N0326_v, N0333_port_0, N0326_port_1);
  spice_transistor_nmos_gnd tM1854(v(SC_v), N0322_v, N0322_port_2);
  spice_transistor_nmos_gnd tM2341(v(_OPE_v), TCS_v, TCS_port_1);
  spice_transistor_nmos_gnd tM1070(v(N0292_v), N0760_v, N0760_port_0);
  spice_transistor_nmos_gnd tM2674(v(clk2_v), N0702_v, N0702_port_0);
  spice_transistor_nmos_gnd tM2671(v(N1000_v), N1001_v, N1001_port_3);
  spice_transistor_nmos tM1572(v(N0620_v), N0632_v, __POC__CLK2_SC_A32_X12__v, N0632_port_9, __POC__CLK2_SC_A32_X12__port_5);
  spice_transistor_nmos tM1988(v(X12_v), __FIN_X12__v, N0639_v, __FIN_X12__port_3, N0639_port_0);
  spice_transistor_nmos tM1981(v(JUN_JMS_v), N0524_v, N0526_v, N0524_port_3, N0526_port_2);
  spice_transistor_nmos_gnd tM1985(v(INC_ISZ_ADD_SUB_XCH_LD_v), N0595_v, N0595_port_1);
  spice_transistor_nmos tM1984(v(X12_v), N0467_v, N0468_v, N0467_port_5, N0468_port_3);
  spice_transistor_nmos tM1509(v(N0545_v), N0565_v, __POC__CLK2_SC_A32_X12__v, N0565_port_9, __POC__CLK2_SC_A32_X12__port_1);
  spice_transistor_nmos tM1508(v(N0545_v), N0544_v, CLK2_SC_A12_M12__v, N0544_port_9, CLK2_SC_A12_M12__port_1);
  spice_transistor_nmos tM1507(v(N0530_v), N0529_v, CLK2_SC_A12_M12__v, N0529_port_9, CLK2_SC_A12_M12__port_0);
  spice_transistor_nmos tM1506(v(N0530_v), N0543_v, __POC__CLK2_SC_A32_X12__v, N0543_port_9, __POC__CLK2_SC_A32_X12__port_0);
  spice_transistor_nmos_gnd tM1501(v(N0919_v), N0544_v, N0544_port_8);
  spice_transistor_nmos_gnd tM1500(v(N0902_v), N0529_v, N0529_port_8);
  spice_transistor_nmos_gnd tM2764(v(WRITE_CARRY_2__v), ADC_CY_v, ADC_CY_port_1);
  spice_transistor_nmos_gnd tM2762(v(READ_ACC_3__v), ACC_ADA_v, ACC_ADA_port_0);
  spice_transistor_nmos_gnd tM2067(v(N0679_v), SC_M22_CLK2_v, SC_M22_CLK2_port_4);
  spice_transistor_nmos_gnd tM2658(v(N0853_v), N0854_v, N0854_port_0);
  spice_transistor_nmos tM1181(v(N0444_v), N0775_v, N0838_v, N0775_port_5, N0838_port_1);
  spice_transistor_nmos_gnd tM1180(v(PC3_6_v), N0838_v, N0838_port_0);
  spice_transistor_nmos tM1183(v(N0410_v), PC1_6_v, N0389_v, PC1_6_port_1, N0389_port_3);
  spice_transistor_nmos tM1182(v(N0381_v), N0389_v, PC0_6_v, N0389_port_2, PC0_6_port_1);
  spice_transistor_nmos tM1185(v(N0410_v), PC1_10_v, N0390_v, PC1_10_port_0, N0390_port_3);
  spice_transistor_nmos tM1184(v(N0381_v), N0390_v, PC0_10_v, N0390_port_2, PC0_10_port_0);
  spice_transistor_nmos_gnd tM1187(v(PC0_10_v), N0790_v, N0790_port_1);
  spice_transistor_nmos tM1189(v(N0439_v), PC3_6_v, N0389_v, PC3_6_port_1, N0389_port_5);
  spice_transistor_nmos tM1188(v(N0426_v), N0389_v, PC2_6_v, N0389_port_4, PC2_6_port_1);
  spice_transistor_nmos_gnd tM1747(v(A32_v), N0279_v, N0279_port_3);
  spice_transistor_nmos_gnd tM1211(v(PC3_10_v), N0839_v, N0839_port_0);
  spice_transistor_nmos tM1210(v(N0434_v), N0827_v, N0772_v, N0827_port_1, N0772_port_4);
  spice_transistor_nmos_gnd tM2763(v(N0342_v), ACC_ADA_v, ACC_ADA_port_1);
  spice_transistor_nmos tM1212(v(N0444_v), N0771_v, N0839_v, N0771_port_5, N0839_port_1);
  spice_transistor_nmos_gnd tM1215(v(N0499_v), N0864_v, N0864_port_0);
  spice_transistor_nmos tM1214(v(RRAB1_v), D2_v, N0535_v, D2_port_5, N0535_port_0);
  spice_transistor_nmos_vdd tM1217(v(__INH__X11_X31_CLK1_v), N0771_v, N0771_port_6);
  spice_transistor_nmos_vdd tM2978(v(N0941_v), _TMP_1_v, _TMP_1_port_1);
  spice_transistor_nmos tM1219(v(WRAB1_v), N0863_v, N0867_v, N0863_port_3, N0867_port_0);
  spice_transistor_nmos tM1218(v(WRAB0_v), N0881_v, N0863_v, N0881_port_0, N0863_port_2);
  spice_transistor_nmos_gnd tM2738(v(SUB_GROUP_6__v), CY_ADAC_v, CY_ADAC_port_0);
  spice_transistor_nmos tM2748(v(M12_v), CY_v, N0470_v, CY_port_1, N0470_port_0);
  spice_transistor_nmos tM2749(v(CY_ADA_v), N0550_v, N0470_v, N0550_port_0, N0470_port_1);
  spice_transistor_nmos_vdd tM2746(v(N0403_v), N0860_v, N0860_port_1);
  spice_transistor_nmos tM2745(v(N0415_v), CY_v, N0860_v, CY_port_0, N0860_port_0);
  spice_transistor_nmos tM2742(v(ADSR_v), CY_1_v, N0513_v, CY_1_port_1, N0513_port_0);
  spice_transistor_nmos tM1439(v(N0544_v), R3_3_v, N0538_v, R3_3_port_0, N0538_port_3);
  spice_transistor_nmos tM1438(v(N0529_v), N0538_v, R1_3_v, N0538_port_2, R1_3_port_0);
  spice_transistor_nmos tM1431(v(N0647_v), R14_2_v, N0536_v, R14_2_port_0, N0536_port_9);
  spice_transistor_nmos tM1430(v(N0634_v), N0536_v, R12_2_v, N0536_port_8, R12_2_port_0);
  spice_transistor_nmos tM1433(v(N0632_v), N0882_v, N0971_v, N0882_port_7, N0971_port_1);
  spice_transistor_nmos_gnd tM1432(v(R10_2_v), N0971_v, N0971_port_0);
  spice_transistor_nmos_gnd tM1435(v(R6_3_v), N0953_v, N0953_port_0);
  spice_transistor_nmos tM1434(v(N0645_v), N0980_v, N0882_v, N0980_port_0, N0882_port_8);
  spice_transistor_nmos tM1437(v(N0544_v), R2_3_v, N0537_v, R2_3_port_1, N0537_port_3);
  spice_transistor_nmos tM1436(v(N0529_v), N0537_v, R0_3_v, N0537_port_2, R0_3_port_1);
  spice_transistor_nmos_gnd tM2632(v(IAC_v), INC_GROUP_5__v, INC_GROUP_5__port_2);
  spice_transistor_nmos_vdd tM2985(v(M12_v), N0605_v, N0605_port_0);
  spice_transistor_nmos_gnd tM2630(v(CMC_v), SUB_GROUP_6__v, SUB_GROUP_6__port_0);
  spice_transistor_nmos_gnd tM2637(v(__X31__CLK2__v), ADD_IB_v, ADD_IB_port_1);
  spice_transistor_nmos_gnd tM2988(v(N0941_v), TMP_1_v, TMP_1_port_2);
  spice_transistor_nmos_gnd tM2989(v(N0700_v), N0690_v, N0690_port_1);
  spice_transistor_nmos tM2568(v(clk2_v), X12_v, N0425_v, X12_port_15, N0425_port_0);
  spice_transistor_nmos_gnd tM3065(v(N0690_v), N0692_v, N0692_port_2);
  spice_transistor_nmos_gnd tM2290(v(N1010_v), N0996_v, N0996_port_2);
  spice_transistor_nmos_gnd tM2291(v(N0994_v), N0995_v, N0995_port_2);
  spice_transistor_nmos_gnd tM2292(v(N0996_v), N0997_v, N0997_port_1);
  spice_transistor_nmos_gnd tM1906(v(N0494_v), __INH__X32_CLK2_v, __INH__X32_CLK2_port_3);
  spice_transistor_nmos_gnd tM2294(v(N0992_v), N0993_v, N0993_port_2);
  spice_transistor_nmos_gnd tM2296(v(N0997_v), _OPR_1_v, _OPR_1_port_16);
  spice_transistor_nmos_gnd tM2297(v(N0996_v), OPR_1_v, OPR_1_port_10);
  spice_transistor_nmos tM1725(v(clk2_v), N0374_v, N0365_v, N0374_port_1, N0365_port_0);
  spice_transistor_nmos tM1724(v(clk2_v), N0384_v, N0379_v, N0384_port_1, N0379_port_0);
  spice_transistor_nmos_gnd tM1727(v(A12_v), N0379_v, N0379_port_1);
  spice_transistor_nmos_vdd tM1726(v(S00609_v), N0710_v, N0710_port_2);
  spice_transistor_nmos tM1721(v(N0459_v), ADDR_PTR_1_v, N0492_v, ADDR_PTR_1_port_2, N0492_port_0);
  spice_transistor_nmos_gnd tM1720(v(N0409_v), N0440_v, N0440_port_3);
  spice_transistor_nmos tM1722(v(N0459_v), N0457_v, N0458_v, N0457_port_2, N0458_port_0);
  spice_transistor_nmos tM2009(v(_OPA_0_v), N0640_v, N0639_v, N0640_port_0, N0639_port_1);
  spice_transistor_nmos_gnd tM1728(v(A22_v), N0365_v, N0365_port_1);
  spice_transistor_nmos tM2767(v(clk1_v), N0686_v, N0675_v, N0686_port_1, N0675_port_2);
  spice_transistor_nmos_gnd tM2188(v(N1008_v), N0992_v, N0992_port_2);
  spice_transistor_nmos tM2189(v(SC_M12_CLK2_v), D1_v, N1010_v, D1_port_8, N1010_port_0);
  spice_transistor_nmos_gnd tM2184(v(N0993_v), _OPR_3_v, _OPR_3_port_11);
  spice_transistor_nmos_gnd tM2187(v(N1011_v), N0998_v, N0998_port_1);
  spice_transistor_nmos tM2181(v(SC_M12_CLK2_v), D0_v, N1011_v, D0_port_7, N1011_port_0);
  spice_transistor_nmos tM2182(v(SC_M12_CLK2_v), D2_v, N1009_v, D2_port_8, N1009_port_0);
  spice_transistor_nmos_gnd tM2364(v(_OPE_v), IAC_v, IAC_port_1);
  spice_transistor_nmos_gnd tM2365(v(_I_O_v), IOR_v, IOR_port_3);
  spice_transistor_nmos tM2366(v(A12_v), N0477_v, N0483_v, N0477_port_2, N0483_port_0);
  spice_transistor_nmos tM2367(v(OPA_IB_v), D2_v, OPA_2_v, D2_port_9, OPA_2_port_0);
  spice_transistor_nmos_gnd tM2360(v(_OPE_v), TCC_v, TCC_port_1);
  spice_transistor_nmos_gnd tM2362(v(_OPE_v), CMC_v, CMC_port_1);
  spice_transistor_nmos_gnd tM2363(v(_OPE_v), DAC_v, DAC_port_1);
  spice_transistor_nmos_gnd tM2368(v(IOR_v), N0483_v, N0483_port_1);
  spice_transistor_nmos_gnd tM2369(v(_OPE_v), CLC_v, CLC_port_1);
  spice_transistor_nmos tM2166(v(OPR_1_v), N0523_v, JCN_ISZ_v, N0523_port_3, JCN_ISZ_port_6);
  spice_transistor_nmos_gnd tM2167(v(OPR_1_v), BBL_v, BBL_port_3);
  spice_transistor_nmos_gnd tM2164(v(OPR_1_v), JUN_JMS_v, JUN_JMS_port_7);
  spice_transistor_nmos_gnd tM2165(v(_OPR_1_v), N0636_v, N0636_port_3);
  spice_transistor_nmos tM2162(v(SC_v), N0368_v, N0373_v, N0368_port_0, N0373_port_3);
  spice_transistor_nmos_gnd tM2163(v(OPR_1_v), JCN_v, JCN_port_2);
  spice_transistor_nmos_gnd tM2160(v(N0362_v), N0361_v, N0361_port_2);
  spice_transistor_nmos tM2161(v(JUN_JMS_v), N0373_v, N0372_v, N0373_port_2, N0372_port_3);
  spice_transistor_nmos_gnd tM2601(v(SUB_v), WRITE_ACC_1__v, WRITE_ACC_1__port_11);
  spice_transistor_nmos_gnd tM2168(v(OPR_1_v), JMS_v, JMS_port_3);
  spice_transistor_nmos tM2169(v(_OPR_1_v), INC_ISZ_XCH_v, N0587_v, INC_ISZ_XCH_port_3, N0587_port_5);
  spice_transistor_nmos_gnd tM2600(v(LD_v), WRITE_ACC_1__v, WRITE_ACC_1__port_10);
  spice_transistor_nmos_gnd tM2970(v(D2_v), N0672_v, N0672_port_0);
  spice_transistor_nmos_gnd tM2605(v(TCC_v), WRITE_CARRY_2__v, WRITE_CARRY_2__port_3);
  spice_transistor_nmos_gnd tM2604(v(SUB_v), WRITE_CARRY_2__v, WRITE_CARRY_2__port_2);
  spice_transistor_nmos_gnd tM3168(v(TCS_v), N0359_v, N0359_port_4);
  spice_transistor_nmos_gnd tM3163(v(N0751_v), N0713_v, N0713_port_1);
  spice_transistor_nmos_vdd tM2004(v(N0621_v), CLK2_SC_A12_M12__v, CLK2_SC_A12_M12__port_9);
  spice_transistor_nmos_gnd tM2410(v(OPA_2_v), CLC_v, CLC_port_3);
  spice_transistor_nmos_gnd tM3014(v(DCL_1_v), N0750_v, N0750_port_0);
  spice_transistor_nmos_gnd tM3017(v(N0729_v), N0747_v, N0747_port_1);
  spice_transistor_nmos_vdd tM3010(v(N0876_v), N0848_v, N0848_port_2);
  spice_transistor_nmos_gnd tM3013(v(N0347_v), N0376_v, N0376_port_3);
  spice_transistor_nmos_gnd tM2609(v(IAC_v), WRITE_CARRY_2__v, WRITE_CARRY_2__port_7);
  spice_transistor_nmos_vdd tM3019(v(S00800_v), N0747_v, N0747_port_2);
  spice_transistor_nmos_gnd tM2608(v(DAC_v), WRITE_CARRY_2__v, WRITE_CARRY_2__port_6);
  spice_transistor_nmos_vdd tM3264(v(S00835_v), N0696_v, N0696_port_3);
  spice_transistor_nmos_gnd tM2419(v(N0782_v), N0784_v, N0784_port_1);
  spice_transistor_nmos_gnd tM3290(v(N0700_v), N0693_v, N0693_port_2);
  spice_transistor_nmos_vdd tM2000(v(S00620_v), N0621_v, N0621_port_1);
  spice_transistor_nmos_gnd tM2786(v(POC_v), N0705_v, N0705_port_2);
  spice_transistor_nmos_gnd tM2787(v(N0702_v), N0706_v, N0706_port_1);
  spice_transistor_nmos tM2759(v(ADSR_v), N0846_v, CY_v, N0846_port_0, CY_port_5);
  spice_transistor_nmos_gnd tM2376(v(N1001_v), _OPA_3_v, _OPA_3_port_10);
  spice_transistor_nmos_gnd tM2894(v(N0884_v), N0847_v, N0847_port_1);
  spice_transistor_nmos_vdd tM2895(v(S00764_v), ACC_ADAC_v, ACC_ADAC_port_3);
  spice_transistor_nmos tM1538(v(N0439_v), PC3_8_v, N0396_v, PC3_8_port_0, N0396_port_5);
  spice_transistor_nmos_gnd tM1539(v(PC1_8_v), N0817_v, N0817_port_0);
  spice_transistor_nmos tM1530(v(clk1_v), N0317_v, N0316_v, N0317_port_0, N0316_port_2);
  spice_transistor_nmos_gnd tM1531(v(N0326_v), WADB0_v, WADB0_port_6);
  spice_transistor_nmos_gnd tM1532(v(PC0_8_v), N0796_v, N0796_port_1);
  spice_transistor_nmos tM1533(v(N0410_v), PC1_8_v, N0396_v, PC1_8_port_0, N0396_port_3);
  spice_transistor_nmos tM1534(v(N0444_v), N0777_v, N0844_v, N0777_port_5, N0844_port_1);
  spice_transistor_nmos tM1535(v(N0426_v), N0395_v, PC2_4_v, N0395_port_4, PC2_4_port_1);
  spice_transistor_nmos tM1536(v(N0439_v), PC3_4_v, N0395_v, PC3_4_port_1, N0395_port_5);
  spice_transistor_nmos tM1537(v(N0426_v), N0396_v, PC2_8_v, N0396_port_4, PC2_8_port_0);
  spice_transistor_nmos_gnd tM1881(v(N0459_v), N0466_v, N0466_port_3);
  spice_transistor_nmos_gnd tM1882(v(N0459_v), ADDR_PTR_0_v, ADDR_PTR_0_port_1);
  spice_transistor_nmos tM1228(v(N0444_v), N0772_v, N0840_v, N0772_port_5, N0840_port_1);
  spice_transistor_nmos tM1229(v(N0439_v), PC3_9_v, N0391_v, PC3_9_port_1, N0391_port_5);
  spice_transistor_nmos_gnd tM1886(v(N0466_v), N0505_v, N0505_port_0);
  spice_transistor_nmos tM1224(v(N0381_v), N0392_v, PC0_5_v, N0392_port_3, PC0_5_port_0);
  spice_transistor_nmos tM1225(v(N0406_v), N0792_v, N0776_v, N0792_port_0, N0776_port_2);
  spice_transistor_nmos_gnd tM1226(v(PC0_5_v), N0792_v, N0792_port_1);
  spice_transistor_nmos tM1227(v(N0426_v), N0391_v, PC2_9_v, N0391_port_4, PC2_9_port_1);
  spice_transistor_nmos tM1220(v(WRAB1_v), N0864_v, N0868_v, N0864_port_1, N0868_port_0);
  spice_transistor_nmos_gnd tM1221(v(PC3_9_v), N0840_v, N0840_port_0);
  spice_transistor_nmos tM1222(v(N0410_v), PC1_9_v, N0391_v, PC1_9_port_1, N0391_port_3);
  spice_transistor_nmos tM1223(v(N0410_v), PC1_5_v, N0392_v, PC1_5_port_0, N0392_port_2);
  spice_transistor_nmos tM1156(v(RRAB0_v), N0533_v, D1_v, N0533_port_0, D1_port_5);
  spice_transistor_nmos tM1157(v(WRAB0_v), N0880_v, N0862_v, N0880_port_0, N0862_port_3);
  spice_transistor_nmos_vdd tM1154(v(__INH__X11_X31_CLK1_v), N0779_v, N0779_port_6);
  spice_transistor_nmos tM1155(v(RRAB1_v), D1_v, N0534_v, D1_port_4, N0534_port_0);
  spice_transistor_nmos tM1152(v(N0434_v), N0825_v, N0775_v, N0825_port_1, N0775_port_4);
  spice_transistor_nmos tM1153(v(N0444_v), N0779_v, N0837_v, N0779_port_5, N0837_port_1);
  spice_transistor_nmos tM1402(v(N0581_v), N0934_v, N0882_v, N0934_port_0, N0882_port_4);
  spice_transistor_nmos tM1151(v(N0424_v), N0775_v, N0810_v, N0775_port_3, N0810_port_1);
  spice_transistor_nmos_gnd tM2754(v(N0342_v), CY_ADAC_v, CY_ADAC_port_1);
  spice_transistor_nmos_gnd tM2757(v(CY_v), N0855_v, N0855_port_1);
  spice_transistor_nmos tM2756(v(ADC_CY_v), N0861_v, CY_v, N0861_port_0, CY_port_3);
  spice_transistor_nmos_gnd tM1408(v(R13_2_v), N0979_v, N0979_port_1);
  spice_transistor_nmos tM1409(v(N0598_v), N0535_v, R9_2_v, N0535_port_6, R9_2_port_1);
  spice_transistor_nmos_gnd tM1158(v(N0880_v), N0532_v, N0532_port_1);
  spice_transistor_nmos tM1159(v(N0543_v), N0903_v, N0866_v, N0903_port_0, N0866_port_2);
  spice_transistor_nmos_gnd tM2523(v(N0360_v), N0337_v, N0337_port_1);
  spice_transistor_nmos tM2520(v(clk2_v), N0282_v, M22_v, N0282_port_1, M22_port_8);
  spice_transistor_nmos tM2521(v(clk1_v), N0721_v, N0720_v, N0721_port_2, N0720_port_1);
  spice_transistor_nmos tM1088(v(N0410_v), PC1_11_v, N0385_v, PC1_11_port_1, N0385_port_3);
  spice_transistor_nmos tM1089(v(N0381_v), N0386_v, PC0_7_v, N0386_port_2, PC0_7_port_0);
  spice_transistor_nmos_gnd tM2623(v(IAC_v), READ_ACC_3__v, READ_ACC_3__port_3);
  spice_transistor_nmos_gnd tM2622(v(TCC_v), ADD_GROUP_4__v, ADD_GROUP_4__port_1);
  spice_transistor_nmos_gnd tM2624(v(DAC_v), READ_ACC_3__v, READ_ACC_3__port_4);
  spice_transistor_nmos_gnd tM2627(v(STC_v), INC_GROUP_5__v, INC_GROUP_5__port_1);
  spice_transistor_nmos_vdd tM2994(v(N0912_v), N0556_v, N0556_port_2);
  spice_transistor_nmos_gnd tM1080(v(PC2_11_v), N0821_v, N0821_port_0);
  spice_transistor_nmos_gnd tM1081(v(PC1_11_v), N0806_v, N0806_port_0);
  spice_transistor_nmos tM1082(v(N0424_v), N0770_v, N0806_v, N0770_port_3, N0806_port_1);
  spice_transistor_nmos tM1083(v(N0434_v), N0821_v, N0770_v, N0821_port_1, N0770_port_4);
  spice_transistor_nmos tM1084(v(N0444_v), N0770_v, N0834_v, N0770_port_5, N0834_port_0);
  spice_transistor_nmos_gnd tM1085(v(PC3_11_v), N0834_v, N0834_port_1);
  spice_transistor_nmos_gnd tM1086(v(N0774_v), N0386_v, N0386_port_1);
  spice_transistor_nmos tM1087(v(N0381_v), N0385_v, PC0_11_v, N0385_port_2, PC0_11_port_1);
  spice_transistor_nmos_vdd tM2579(v(N0745_v), M12_v, M12_port_10);
  spice_transistor_nmos_gnd tM2578(v(M12_v), N0288_v, N0288_port_3);
  spice_transistor_nmos_gnd tM2852(v(M12_v), N0870_v, N0870_port_2);
  spice_transistor_nmos_gnd tM2571(v(N0422_v), N0805_v, N0805_port_2);
  spice_transistor_nmos tM2570(v(N0423_v), N0421_v, N0422_v, N0421_port_1, N0422_port_0);
  spice_transistor_nmos_gnd tM2573(v(N0433_v), N0430_v, N0430_port_2);
  spice_transistor_nmos_gnd tM2572(v(X12_v), N0853_v, N0853_port_1);
  spice_transistor_nmos_gnd tM1711(v(N0400_v), N0427_v, N0427_port_3);
  spice_transistor_nmos_gnd tM1713(v(N0464_v), N0475_v, N0475_port_1);
  spice_transistor_nmos_gnd tM1715(v(N0464_v), ADDR_PTR_1_v, ADDR_PTR_1_port_1);
  spice_transistor_nmos_gnd tM1716(v(N0475_v), N0464_v, N0464_port_2);
  spice_transistor_nmos_gnd tM1718(v(N0475_v), N0457_v, N0457_port_0);
  spice_transistor_nmos tM2987(v(SUB_GROUP_6__v), _TMP_1_v, N0889_v, _TMP_1_port_2, N0889_port_5);
  spice_transistor_nmos_gnd tM2199(v(_OPR_0_v), JIN_FIN_v, JIN_FIN_port_7);
  spice_transistor_nmos_gnd tM2198(v(_OPR_0_v), OPE_v, OPE_port_3);
  spice_transistor_nmos_gnd tM2193(v(OPR_1_v), SUB_v, SUB_port_2);
  spice_transistor_nmos_gnd tM2191(v(N1009_v), N0994_v, N0994_port_3);
  spice_transistor_nmos tM2038(v(clk2_v), N0562_v, N0547_v, N0562_port_1, N0547_port_2);
  spice_transistor_nmos_gnd tM2196(v(_OPR_0_v), ISZ_v, ISZ_port_3);
  spice_transistor_nmos_gnd tM2195(v(OPR_1_v), LDM_BBL_v, LDM_BBL_port_2);
  spice_transistor_nmos_gnd tM2194(v(OPR_1_v), ADD_v, ADD_port_2);
  spice_transistor_nmos_gnd tM2373(v(_OPA_3_v), SBM_v, SBM_port_2);
  spice_transistor_nmos_gnd tM2371(v(_OPA_3_v), STC_v, STC_port_2);
  spice_transistor_nmos_gnd tM2370(v(_OPE_v), CLB_v, CLB_port_1);
  spice_transistor_nmos_gnd tM2377(v(N1000_v), OPA_3_v, OPA_3_port_2);
  spice_transistor_nmos_gnd tM2090(v(OPR_3_v), ISZ_v, ISZ_port_0);
  spice_transistor_nmos_gnd tM2375(v(_OPA_3_v), IOR_v, IOR_port_5);
  spice_transistor_nmos_gnd tM2379(v(OPA_3_v), IOW_v, IOW_port_2);
  spice_transistor_nmos_gnd tM2378(v(OPA_3_v), O_IB_v, O_IB_port_2);
  spice_transistor_nmos_vdd tM2175(v(N0993_v), OPR_3_v, OPR_3_port_14);
  spice_transistor_nmos_vdd tM2176(v(N0992_v), _OPR_3_v, _OPR_3_port_10);
  spice_transistor_nmos_gnd tM2171(v(_OPR_1_v), LD_v, LD_port_2);
  spice_transistor_nmos_gnd tM2170(v(_OPR_1_v), FIN_FIM_SRC_JIN_v, FIN_FIM_SRC_JIN_port_5);
  spice_transistor_nmos_gnd tM2173(v(N0994_v), OPR_2_v, OPR_2_port_14);
  spice_transistor_nmos_gnd tM2172(v(N0995_v), _OPR_2_v, _OPR_2_port_13);
  spice_transistor_nmos_gnd tM2179(v(N0660_v), SC_M12_CLK2_v, SC_M12_CLK2_port_0);
  spice_transistor_nmos_gnd tM2668(v(SUB_v), SUB_GROUP_6__v, SUB_GROUP_6__port_3);
  spice_transistor_nmos_vdd tM2287(v(N0996_v), _OPR_1_v, _OPR_1_port_15);
  spice_transistor_nmos_gnd tM2286(v(N0999_v), _OPR_0_v, _OPR_0_port_11);
  spice_transistor_nmos_gnd tM2285(v(N0998_v), OPR_0_v, OPR_0_port_6);
  spice_transistor_nmos_gnd tM2099(v(OPR_3_v), JMS_v, JMS_port_1);
  spice_transistor_nmos_gnd tM2289(v(N0998_v), N0999_v, N0999_port_2);
  spice_transistor_nmos_vdd tM2288(v(N0997_v), OPR_1_v, OPR_1_port_9);
  spice_transistor_nmos_gnd tM3151(v(N0715_v), N0735_v, N0735_port_1);
  spice_transistor_nmos_vdd tM3152(v(S00825_v), N0715_v, N0715_port_4);
  spice_transistor_nmos_gnd tM3158(v(N0734_v), cm_ram3_v, cm_ram3_port_1);
  spice_transistor_nmos_gnd tM3159(v(_COM_v), N0713_v, N0713_port_0);
  spice_transistor_nmos_gnd tM1404(v(R2_3_v), N0926_v, N0926_port_0);
  spice_transistor_nmos_gnd tM3080(v(N0943_v), N0944_v, N0944_port_2);
  spice_transistor_nmos_vdd tM2986(v(N0942_v), TMP_1_v, TMP_1_port_1);
  spice_transistor_nmos_gnd tM2665(v(IOR_v), WRITE_ACC_1__v, WRITE_ACC_1__port_14);
  spice_transistor_nmos tM3020(v(N0766_v), N0750_v, N0765_v, N0750_port_2, N0765_port_2);
  spice_transistor_nmos tM3022(v(N0351_v), N0355_v, N0768_v, N0355_port_1, N0768_port_0);
  spice_transistor_nmos_gnd tM3023(v(N0355_v), N0354_v, N0354_port_4);
  spice_transistor_nmos_gnd tM3024(v(N0348_v), N0355_v, N0355_port_3);
  spice_transistor_nmos_gnd tM3025(v(N0348_v), ACC_0_v, ACC_0_port_9);
  spice_transistor_nmos tM3026(v(ADSL_v), N0847_v, ACC_2_v, N0847_port_6, ACC_2_port_0);
  spice_transistor_nmos_gnd tM3027(v(ACC_2_v), N0858_v, N0858_port_3);
  spice_transistor_nmos_gnd tM3029(v(N0848_v), ADD_0_v, ADD_0_port_4);
  spice_transistor_nmos_gnd tM2805(v(N0849_v), N0346_v, N0346_port_0);
  spice_transistor_nmos tM2801(v(N0550_v), N0886_v, N0894_v, N0886_port_0, N0894_port_0);
  spice_transistor_nmos_gnd tM2800(v(M12_v), SUB_GROUP_6__v, SUB_GROUP_6__port_6);
  spice_transistor_nmos_gnd tM2908(v(N0350_v), N0363_v, N0363_port_1);
  spice_transistor_nmos_gnd tM2909(v(N0350_v), N0370_v, N0370_port_1);
  spice_transistor_nmos tM1401(v(N0565_v), N0882_v, N0925_v, N0882_port_3, N0925_port_1);
  spice_transistor_nmos_gnd tM2618(v(N0442_v), ADD_IB_v, ADD_IB_port_0);
  spice_transistor_nmos_vdd tM3087(v(S00801_v), N0943_v, N0943_port_3);
  spice_transistor_nmos tM2902(v(N0766_v), N0751_v, N0767_v, N0751_port_2, N0767_port_0);
  spice_transistor_nmos_gnd tM2903(v(POC_v), DCL_0_v, DCL_0_port_3);
  spice_transistor_nmos tM3167(v(N0415_v), D3_v, N0358_v, D3_port_15, N0358_port_7);
  spice_transistor_nmos_gnd tM2619(v(XCH_v), N0445_v, N0445_port_1);
  spice_transistor_nmos_gnd tM2663(v(ADD_v), WRITE_CARRY_2__v, WRITE_CARRY_2__port_13);
  spice_transistor_nmos tM1888(v(clk1_v), N0521_v, ADDR_PTR_0_v, N0521_port_0, ADDR_PTR_0_port_3);
  spice_transistor_nmos tM1889(v(clk1_v), N0505_v, N0506_v, N0505_port_2, N0506_port_0);
  spice_transistor_nmos_gnd tM3239(v(N0670_v), N0669_v, N0669_port_0);
  spice_transistor_nmos_gnd tM3238(v(N0670_v), D0_v, D0_port_16);
  spice_transistor_nmos tM1405(v(N0583_v), R6_2_v, N0536_v, R6_2_port_0, N0536_port_5);
  spice_transistor_nmos tM1406(v(N0632_v), N0868_v, N0970_v, N0868_port_7, N0970_port_1);
  spice_transistor_nmos_gnd tM2328(v(test_v), N0432_v, N0432_port_0);
  spice_transistor_nmos tM1407(v(N0645_v), N0979_v, N0868_v, N0979_port_0, N0868_port_8);
  spice_transistor_nmos_gnd tM1400(v(R2_2_v), N0925_v, N0925_port_0);
  spice_transistor_nmos_gnd tM3303(v(N0664_v), N0663_v, N0663_port_2);
  spice_transistor_nmos_gnd tM1150(v(PC2_6_v), N0825_v, N0825_port_0);
  spice_transistor_nmos_vdd tM3235(v(S00817_v), N0945_v, N0945_port_4);
  spice_transistor_nmos_gnd tM1403(v(R4_2_v), N0934_v, N0934_port_1);
  spice_transistor_nmos_gnd tM1239(v(PC3_5_v), N0841_v, N0841_port_0);
  spice_transistor_nmos tM1238(v(N0439_v), PC3_5_v, N0392_v, PC3_5_port_0, N0392_port_5);
  spice_transistor_nmos_gnd tM3237(v(d0_v), N0670_v, N0670_port_0);
  spice_transistor_nmos_gnd tM1899(v(N0521_v), N0520_v, N0520_port_0);
  spice_transistor_nmos_gnd tM1233(v(N0780_v), N0393_v, N0393_port_1);
  spice_transistor_nmos_gnd tM1232(v(PC0_1_v), N0793_v, N0793_port_0);
  spice_transistor_nmos_gnd tM1231(v(PC1_5_v), N0813_v, N0813_port_0);
  spice_transistor_nmos tM1230(v(N0426_v), N0392_v, PC2_5_v, N0392_port_4, PC2_5_port_0);
  spice_transistor_nmos_gnd tM1237(v(PC2_5_v), N0828_v, N0828_port_1);
  spice_transistor_nmos tM1235(v(N0424_v), N0776_v, N0813_v, N0776_port_3, N0813_port_1);
  spice_transistor_nmos tM1234(v(N0406_v), N0793_v, N0780_v, N0793_port_1, N0780_port_2);
  spice_transistor_nmos_gnd tM1145(v(N0498_v), N0863_v, N0863_port_1);
  spice_transistor_nmos_vdd tM1412(v(SC_A22_M22_CLK2_v), N0881_v, N0881_port_10);
  spice_transistor_nmos tM1411(v(N0657_v), N0867_v, N0987_v, N0867_port_9, N0987_port_1);
  spice_transistor_nmos tM1410(v(N0619_v), R11_2_v, N0535_v, R11_2_port_1, N0535_port_7);
  spice_transistor_nmos tM1417(v(N0657_v), N0868_v, N0988_v, N0868_port_9, N0988_port_1);
  spice_transistor_nmos_gnd tM1416(v(R15_2_v), N0988_v, N0988_port_0);
  spice_transistor_nmos_vdd tM1415(v(SC_A22_M22_CLK2_v), N0867_v, N0867_port_10);
  spice_transistor_nmos tM1142(v(N0424_v), N0779_v, N0809_v, N0779_port_3, N0809_port_1);
  spice_transistor_nmos_vdd tM2760(v(S00732_v), CY_ADAC_v, CY_ADAC_port_2);
  spice_transistor_nmos tM1013(v(RADB2_v), N0385_v, D3_v, N0385_port_1, D3_port_1);
  spice_transistor_nmos_gnd tM1419(v(N0869_v), N0538_v, N0538_port_1);
  spice_transistor_nmos tM1418(v(N0598_v), N0536_v, R8_2_v, N0536_port_6, R8_2_port_0);
  spice_transistor_nmos_gnd tM1149(v(PC1_6_v), N0810_v, N0810_port_0);
  spice_transistor_nmos_gnd tM1148(v(PC3_2_v), N0837_v, N0837_port_0);
  spice_transistor_nmos_gnd tM2766(v(clk1_v), N0678_v, N0678_port_1);
  spice_transistor_nmos_vdd tM2699(v(S00687_v), N0687_v, N0687_port_0);
  spice_transistor_nmos tM2752(v(ADSL_v), N0513_v, CY_v, N0513_port_1, CY_port_2);
  spice_transistor_nmos tM1097(v(N0406_v), N0787_v, N0778_v, N0787_port_0, N0778_port_2);
  spice_transistor_nmos_gnd tM1096(v(N0778_v), N0387_v, N0387_port_1);
  spice_transistor_nmos tM1095(v(N0426_v), N0386_v, PC2_7_v, N0386_port_4, PC2_7_port_0);
  spice_transistor_nmos tM1094(v(N0439_v), PC3_11_v, N0385_v, PC3_11_port_1, N0385_port_5);
  spice_transistor_nmos tM1093(v(N0426_v), N0385_v, PC2_11_v, N0385_port_4, PC2_11_port_1);
  spice_transistor_nmos_gnd tM1092(v(PC0_7_v), N0786_v, N0786_port_1);
  spice_transistor_nmos tM1091(v(N0406_v), N0786_v, N0774_v, N0786_port_0, N0774_port_2);
  spice_transistor_nmos tM1090(v(N0410_v), PC1_7_v, N0386_v, PC1_7_port_0, N0386_port_3);
  spice_transistor_nmos_gnd tM1099(v(PC1_7_v), N0807_v, N0807_port_0);
  spice_transistor_nmos_gnd tM1098(v(PC0_3_v), N0787_v, N0787_port_1);
  spice_transistor_nmos_gnd tM1527(v(N0300_v), WADB0_v, WADB0_port_5);
  spice_transistor_nmos_gnd tM1525(v(N0315_v), N0316_v, N0316_port_0);
  spice_transistor_nmos_gnd tM1524(v(A12_v), N0711_v, N0711_port_0);
  spice_transistor_nmos tM1522(v(vcc_v), N0325_v, clk1_v, N0325_port_6, clk1_port_1);
  spice_transistor_nmos_gnd tM2614(v(RAR_v), READ_ACC_3__v, READ_ACC_3__port_1);
  spice_transistor_nmos_gnd tM2615(v(RAL_v), READ_ACC_3__v, READ_ACC_3__port_2);
  spice_transistor_nmos tM2616(v(N0445_v), N0448_v, ACB_IB_v, N0448_port_2, ACB_IB_port_0);
  spice_transistor_nmos tM2617(v(__X31__CLK2__v), ACB_IB_v, N0448_v, ACB_IB_port_1, N0448_port_3);
  spice_transistor_nmos_gnd tM2612(v(SBM_v), WRITE_CARRY_2__v, WRITE_CARRY_2__port_10);
  spice_transistor_nmos_gnd tM2613(v(ADM_v), WRITE_CARRY_2__v, WRITE_CARRY_2__port_11);
  spice_transistor_nmos tM2918(v(N0553_v), N0888_v, N0895_v, N0888_port_0, N0895_port_0);
  spice_transistor_nmos_gnd tM1707(v(N0561_v), N0648_v, N0648_port_6);
  spice_transistor_nmos_gnd tM1706(v(N0561_v), N0635_v, N0635_port_6);
  spice_transistor_nmos_gnd tM1705(v(N0561_v), N0620_v, N0620_port_6);
  spice_transistor_nmos_gnd tM1704(v(N0561_v), N0599_v, N0599_port_6);
  spice_transistor_nmos_gnd tM1703(v(N0561_v), N0584_v, N0584_port_6);
  spice_transistor_nmos_gnd tM1702(v(N0561_v), N0570_v, N0570_port_6);
  spice_transistor_nmos_gnd tM1701(v(N0561_v), N0545_v, N0545_port_6);
  spice_transistor_nmos_gnd tM1700(v(N0560_v), N0648_v, N0648_port_5);
  spice_transistor_nmos_gnd tM1205(v(N0776_v), N0392_v, N0392_port_1);
  spice_transistor_nmos_gnd tM2388(v(OPA_2_v), N0501_v, N0501_port_0);
  spice_transistor_nmos tM2389(v(ACC_0_v), N0501_v, N0486_v, N0501_port_1, N0486_port_2);
  spice_transistor_nmos_gnd tM2386(v(N0486_v), N0487_v, N0487_port_1);
  spice_transistor_nmos_gnd tM2387(v(_OPA_2_v), DCL_v, DCL_port_3);
  spice_transistor_nmos_gnd tM2384(v(OPA_3_v), CMC_v, CMC_port_2);
  spice_transistor_nmos_gnd tM2385(v(OPA_3_v), IAC_v, IAC_port_2);
  spice_transistor_nmos_gnd tM2382(v(OPA_3_v), CMA_v, CMA_port_2);
  spice_transistor_nmos_gnd tM2383(v(OPA_3_v), TCC_v, TCC_port_2);
  spice_transistor_nmos_gnd tM2380(v(OPA_3_v), RAR_v, RAR_port_2);
  spice_transistor_nmos_gnd tM2381(v(OPA_3_v), RAL_v, RAL_port_2);
  spice_transistor_nmos_gnd tM2140(v(OPR_2_v), N0628_v, N0628_port_3);
  spice_transistor_nmos_vdd tM2141(v(N0995_v), OPR_2_v, OPR_2_port_8);
  spice_transistor_nmos_vdd tM2142(v(N0994_v), _OPR_2_v, _OPR_2_port_12);
  spice_transistor_nmos tM2143(v(OPR_2_v), N0587_v, INC_ISZ_XCH_v, N0587_port_3, INC_ISZ_XCH_port_2);
  spice_transistor_nmos_gnd tM2144(v(OPR_2_v), FIN_FIM_SRC_JIN_v, FIN_FIM_SRC_JIN_port_4);
  spice_transistor_nmos_gnd tM2145(v(_OPR_1_v), FIM_SRC_v, FIM_SRC_port_2);
  spice_transistor_nmos_gnd tM2146(v(_OPR_1_v), IO_v, IO_port_2);
  spice_transistor_nmos_gnd tM2147(v(_OPR_1_v), OPE_v, OPE_port_2);
  spice_transistor_nmos_gnd tM2148(v(_OPR_1_v), JIN_FIN_v, JIN_FIN_port_6);
  spice_transistor_nmos_gnd tM2149(v(_OPR_1_v), INC_ISZ_v, INC_ISZ_port_3);
  spice_transistor_nmos_gnd tM1967(v(N0578_v), WRAB1_v, WRAB1_port_4);
  spice_transistor_nmos_gnd tM2544(v(N0446_v), N0448_v, N0448_port_0);
  spice_transistor_nmos_gnd tM2547(v(M22_v), N0288_v, N0288_port_2);
  spice_transistor_nmos_gnd tM2812(v(N0725_v), N0745_v, N0745_port_1);
  spice_transistor_nmos_gnd tM2541(v(TCS_v), WRITE_CARRY_2__v, WRITE_CARRY_2__port_0);
  spice_transistor_nmos_gnd tM2542(v(TCS_v), ADD_GROUP_4__v, ADD_GROUP_4__port_0);
  spice_transistor_nmos_gnd tM2543(v(DAA_v), READ_ACC_3__v, READ_ACC_3__port_0);
  spice_transistor_nmos tM1963(v(N0600_v), N0653_v, N0641_v, N0653_port_0, N0641_port_1);
  spice_transistor_nmos_vdd tM2548(v(N0744_v), M22_v, M22_port_10);
  spice_transistor_nmos_gnd tM2549(v(N0723_v), M22_v, M22_port_11);
  spice_transistor_nmos_gnd tM2818(v(N0284_v), N0724_v, N0724_port_1);
  spice_transistor_nmos_gnd tM1962(v(N0633_v), N0638_v, N0638_port_1);
  spice_transistor_nmos_gnd tM3142(v(N0356_v), ACC_0_v, ACC_0_port_10);
  spice_transistor_nmos_gnd tM3141(v(N0403_v), N0358_v, N0358_port_6);
  spice_transistor_nmos_gnd tM3140(v(N0377_v), N0366_v, N0366_port_4);
  spice_transistor_nmos_gnd tM1961(v(N0642_v), N0637_v, N0637_port_2);
  spice_transistor_nmos_gnd tM3144(v(N0852_v), N0356_v, N0356_port_8);
  spice_transistor_nmos_gnd tM1960(v(N0642_v), REG_RFSH_2_v, REG_RFSH_2_port_3);
  spice_transistor_nmos_gnd tM2621(v(IOW_v), N0446_v, N0446_port_2);
  spice_transistor_nmos_gnd tM2620(v(N0446_v), CY_IB_v, CY_IB_port_0);
  spice_transistor_nmos_gnd tM2991(v(N0916_v), N0556_v, N0556_port_1);
  spice_transistor_nmos tM2678(v(OPA_IB_v), D0_v, OPA_0_v, D0_port_8, OPA_0_port_11);
  spice_transistor_nmos tM2990(v(N0964_v), D1_v, N0605_v, D1_port_14, N0605_port_1);
  spice_transistor_nmos_gnd tM2625(v(SBM_v), READ_ACC_3__v, READ_ACC_3__port_5);
  spice_transistor_nmos_gnd tM1968(v(N0649_v), SC_A12_CLK2_v, SC_A12_CLK2_port_2);
  spice_transistor_nmos_vdd tM2996(v(S00781_v), N0941_v, N0941_port_4);
  spice_transistor_nmos_gnd tM2679(v(N1007_v), _OPA_0_v, _OPA_0_port_13);
  spice_transistor_nmos_gnd tM2629(v(__X31__CLK2__v), CY_IB_v, CY_IB_port_1);
  spice_transistor_nmos_gnd tM3039(v(M12_v), N0872_v, N0872_port_3);
  spice_transistor_nmos_gnd tM2628(v(RAL_v), N0502_v, N0502_port_0);
  spice_transistor_nmos_gnd tM3037(v(N0872_v), N0554_v, N0554_port_0);
  spice_transistor_nmos tM3036(v(N0891_v), N0879_v, N0890_v, N0879_port_1, N0890_port_1);
  spice_transistor_nmos_gnd tM3035(v(N0872_v), N0896_v, N0896_port_1);
  spice_transistor_nmos tM3034(v(N0556_v), N0890_v, N0896_v, N0890_port_0, N0896_port_0);
  spice_transistor_nmos_gnd tM3033(v(N0858_v), N0473_v, N0473_port_2);
  spice_transistor_nmos tM3032(v(M12_v), ACC_2_v, N0473_v, ACC_2_port_3, N0473_port_1);
  spice_transistor_nmos tM3031(v(ADD_ACC_v), N0848_v, ACC_2_v, N0848_port_4, ACC_2_port_2);
  spice_transistor_nmos tM3030(v(ACB_IB_v), N0348_v, D2_v, N0348_port_5, D2_port_13);
  spice_transistor_nmos_gnd tM3146(v(TCS_v), N0366_v, N0366_port_5);
  spice_transistor_nmos_gnd tM2471(v(OPA_1_v), DCL_v, DCL_port_4);
  spice_transistor_nmos_gnd tM2472(v(OPA_1_v), KBP_v, KBP_port_4);
  spice_transistor_nmos tM3042(v(N0872_v), N0555_v, N0913_v, N0555_port_1, N0913_port_0);
  spice_transistor_nmos_gnd tM2473(v(OPA_1_v), TCS_v, TCS_port_4);
  spice_transistor_nmos_vdd tM2977(v(S00765_v), N0690_v, N0690_port_0);
  spice_transistor_nmos_gnd tM3041(v(N0891_v), N0555_v, N0555_port_0);
  spice_transistor_nmos tM3046(v(ACC_ADA_v), N0872_v, N0473_v, N0872_port_5, N0473_port_3);
  spice_transistor_nmos tM1895(v(clk1_v), N0586_v, N0573_v, N0586_port_0, N0573_port_1);
  spice_transistor_nmos tM3045(v(ADD_IB_v), D2_v, N0848_v, D2_port_14, N0848_port_5);
  spice_transistor_nmos_gnd tM2574(v(N0425_v), N0421_v, N0421_port_2);
  spice_transistor_nmos_gnd tM3180(v(N0885_v), N0514_v, N0514_port_4);
  spice_transistor_nmos_gnd tM2577(v(N0431_v), N0801_v, N0801_port_2);
  spice_transistor_nmos_gnd tM1893(v(N0574_v), REG_RFSH_0_v, REG_RFSH_0_port_3);
  spice_transistor_nmos tM2673(v(OPA_IB_v), D1_v, OPA_1_v, D1_port_9, OPA_1_port_12);
  spice_transistor_nmos_gnd tM1892(v(N0566_v), N0572_v, N0572_port_1);
  spice_transistor_nmos_vdd tM2670(v(N1003_v), OPA_2_v, OPA_2_port_13);
  spice_transistor_nmos tM1958(v(N0600_v), REG_RFSH_2_v, N0633_v, REG_RFSH_2_port_2, N0633_port_0);
  spice_transistor_nmos tM1959(v(N0610_v), N0637_v, N0638_v, N0637_port_1, N0638_port_0);
  spice_transistor_nmos tM1956(v(SC_A22_v), N0646_v, REG_RFSH_2_v, N0646_port_2, REG_RFSH_2_port_0);
  spice_transistor_nmos tM1952(v(SC_M22_CLK2_v), D3_v, N0646_v, D3_port_7, N0646_port_1);
  spice_transistor_nmos tM1950(v(N0574_v), N0610_v, N0624_v, N0610_port_4, N0624_port_0);
  spice_transistor_nmos_gnd tM1951(v(N0625_v), N0624_v, N0624_port_1);
  spice_transistor_nmos_gnd tM2705(v(N0688_v), N0687_v, N0687_port_2);
  spice_transistor_nmos_vdd tM1395(v(__INH__X11_X31_CLK1_v), N0780_v, N0780_port_6);
  spice_transistor_nmos tM1396(v(WRAB0_v), N0883_v, N0865_v, N0883_port_0, N0865_port_2);
  spice_transistor_nmos tM1397(v(WRAB1_v), N0865_v, N0869_v, N0865_port_3, N0869_port_0);
  spice_transistor_nmos tM1390(v(WADB2_v), N0773_v, N0764_v, N0773_port_1, N0764_port_5);
  spice_transistor_nmos tM1391(v(N0381_v), N0395_v, PC0_4_v, N0395_port_2, PC0_4_port_1);
  spice_transistor_nmos tM1392(v(N0434_v), N0831_v, N0777_v, N0831_port_0, N0777_port_4);
  spice_transistor_nmos_gnd tM1393(v(PC2_4_v), N0831_v, N0831_port_1);
  spice_transistor_nmos_gnd tM1398(v(N0883_v), N0537_v, N0537_port_1);
  spice_transistor_nmos tM1399(v(N0543_v), N0909_v, N0883_v, N0909_port_1, N0883_port_2);
  spice_transistor_nmos_gnd tM2877(v(N0887_v), N0898_v, N0898_port_3);
  spice_transistor_nmos tM2872(v(ADSR_v), N0847_v, ACC_0_v, N0847_port_0, ACC_0_port_7);
  spice_transistor_nmos_gnd tM3289(v(N0694_v), N0693_v, N0693_port_1);
  spice_transistor_nmos_vdd tM3210(v(S00804_v), N0914_v, N0914_port_2);
  spice_transistor_nmos tM1170(v(N0529_v), N0531_v, R1_0_v, N0531_port_2, R1_0_port_1);
  spice_transistor_nmos tM1171(v(N0544_v), R3_0_v, N0531_v, R3_0_port_1, N0531_port_3);
  spice_transistor_nmos tM1172(v(N0569_v), N0531_v, R5_0_v, N0531_port_4, R5_0_port_1);
  spice_transistor_nmos tM1174(v(N0544_v), R2_0_v, N0532_v, R2_0_port_0, N0532_port_3);
  spice_transistor_nmos tM1175(v(N0543_v), N0904_v, N0880_v, N0904_port_0, N0880_port_2);
  spice_transistor_nmos_gnd tM1176(v(R0_0_v), N0904_v, N0904_port_1);
  spice_transistor_nmos tM1177(v(N0583_v), R7_0_v, N0531_v, R7_0_port_1, N0531_port_5);
  spice_transistor_nmos_gnd tM1178(v(R0_1_v), N0905_v, N0905_port_0);
  spice_transistor_nmos tM1179(v(M12_M22_CLK1__M11_M12__v), N0498_v, D1_v, N0498_port_1, D1_port_6);
  spice_transistor_nmos_gnd tM1553(v(N0928_v), N0581_v, N0581_port_8);
  spice_transistor_nmos_gnd tM1550(v(N0454_v), N0462_v, N0462_port_0);
  spice_transistor_nmos tM1551(v(N0463_v), N0461_v, N0462_v, N0461_port_4, N0462_port_1);
  spice_transistor_nmos_gnd tM1556(v(N0938_v), N0591_v, N0591_port_8);
  spice_transistor_nmos_gnd tM1557(v(N0955_v), N0616_v, N0616_port_8);
  spice_transistor_nmos_gnd tM1554(v(N0928_v), N0569_v, N0569_port_8);
  spice_transistor_nmos_gnd tM1555(v(N0938_v), N0583_v, N0583_port_8);
  spice_transistor_nmos_gnd tM2603(v(LDM_BBL_v), WRITE_ACC_1__v, WRITE_ACC_1__port_13);
  spice_transistor_nmos_gnd tM2602(v(ADD_v), WRITE_ACC_1__v, WRITE_ACC_1__port_12);
  spice_transistor_nmos tM1558(v(N0570_v), N0581_v, __POC__CLK2_SC_A32_X12__v, N0581_port_9, __POC__CLK2_SC_A32_X12__port_2);
  spice_transistor_nmos tM1559(v(N0570_v), N0569_v, CLK2_SC_A12_M12__v, N0569_port_9, CLK2_SC_A12_M12__port_2);
  spice_transistor_nmos_gnd tM2607(v(CMC_v), WRITE_CARRY_2__v, WRITE_CARRY_2__port_5);
  spice_transistor_nmos_gnd tM2606(v(STC_v), WRITE_CARRY_2__v, WRITE_CARRY_2__port_4);
  spice_transistor_nmos_vdd tM1779(v(S00585_v), N0648_v, N0648_port_7);
  spice_transistor_nmos tM1272(v(N0619_v), R11_0_v, N0531_v, R11_0_port_1, N0531_port_7);
  spice_transistor_nmos_vdd tM1772(v(S00584_v), N0635_v, N0635_port_7);
  spice_transistor_nmos_vdd tM1770(v(S00582_v), N0599_v, N0599_port_7);
  spice_transistor_nmos_vdd tM1771(v(S00583_v), N0620_v, N0620_port_7);
  spice_transistor_nmos_gnd tM1776(v(N0560_v), N0542_v, N0542_port_5);
  spice_transistor_nmos_gnd tM1777(v(N0582_v), N0560_v, N0560_port_5);
  spice_transistor_nmos_gnd tM2197(v(_OPR_0_v), JCN_v, JCN_port_3);
  spice_transistor_nmos_vdd tM2777(v(S00734_v), CY_ADA_v, CY_ADA_port_3);
  spice_transistor_nmos_gnd tM2775(v(N0477_v), ADD_ACC_v, ADD_ACC_port_1);
  spice_transistor_nmos tM1271(v(N0598_v), N0531_v, R9_0_v, N0531_port_6, R9_0_port_1);
  spice_transistor_nmos_gnd tM2772(v(N0685_v), N0678_v, N0678_port_4);
  spice_transistor_nmos_vdd tM2771(v(N0677_v), N0676_v, N0676_port_0);
  spice_transistor_nmos tM2770(v(N0702_v), N0701_v, N0699_v, N0701_port_3, N0699_port_1);
  spice_transistor_nmos_gnd tM2398(v(_OPA_2_v), TCC_v, TCC_port_3);
  spice_transistor_nmos tM2682(v(N0702_v), N0671_v, N0688_v, N0671_port_1, N0688_port_0);
  spice_transistor_nmos_gnd tM2372(v(_OPA_3_v), DAC_v, DAC_port_2);
  spice_transistor_nmos_gnd tM2395(v(OPA_3_v), CLC_v, CLC_port_2);
  spice_transistor_nmos_gnd tM2394(v(_OPA_2_v), RAL_v, RAL_port_3);
  spice_transistor_nmos_gnd tM2397(v(_OPA_2_v), CMA_v, CMA_port_3);
  spice_transistor_nmos_gnd tM2396(v(OPA_3_v), CLB_v, CLB_port_2);
  spice_transistor_nmos_gnd tM2393(v(_OPA_2_v), RAR_v, RAR_port_3);
  spice_transistor_nmos_gnd tM2392(v(_OPA_2_v), KBP_v, KBP_port_3);
  spice_transistor_nmos_gnd tM1604(v(N0455_v), ADDR_RFSH_0_v, ADDR_RFSH_0_port_1);
  spice_transistor_nmos_gnd tM1605(v(N0463_v), N0503_v, N0503_port_0);
  spice_transistor_nmos_gnd tM1600(v(N0540_v), N0539_v, N0539_port_0);
  spice_transistor_nmos_gnd tM2158(v(X32_v), N0372_v, N0372_port_2);
  spice_transistor_nmos tM2157(v(clk1_v), N0361_v, N0343_v, N0361_port_1, N0343_port_2);
  spice_transistor_nmos_gnd tM2156(v(_OPR_1_v), N0587_v, N0587_port_4);
  spice_transistor_nmos tM2155(v(_OPR_1_v), N0628_v, INC_ISZ_ADD_SUB_XCH_LD_v, N0628_port_4, INC_ISZ_ADD_SUB_XCH_LD_port_4);
  spice_transistor_nmos_gnd tM2154(v(OPR_2_v), ADD_v, ADD_port_1);
  spice_transistor_nmos_gnd tM2153(v(OPR_2_v), SUB_v, SUB_port_1);
  spice_transistor_nmos_gnd tM2152(v(OPR_2_v), LD_v, LD_port_1);
  spice_transistor_nmos_gnd tM2151(v(_OPR_1_v), XCH_v, XCH_port_2);
  spice_transistor_nmos_vdd tM1609(v(S00564_v), RRAB0_v, RRAB0_port_4);
  spice_transistor_nmos_gnd tM2374(v(_OPA_3_v), ADM_v, ADM_port_2);
  spice_transistor_nmos_vdd tM2553(v(S00740_v), N0744_v, N0744_port_2);
  spice_transistor_nmos_gnd tM2551(v(N0723_v), N0744_v, N0744_port_1);
  spice_transistor_nmos tM2806(v(N0854_v), N0856_v, N0849_v, N0856_port_0, N0849_port_1);
  spice_transistor_nmos_gnd tM2557(v(N0283_v), N0722_v, N0722_port_0);
  spice_transistor_nmos tM2556(v(N0423_v), N0430_v, N0431_v, N0430_port_1, N0431_port_0);
  spice_transistor_nmos_gnd tM2803(v(N0878_v), N0846_v, N0846_port_1);
  spice_transistor_nmos tM2802(v(N0550_v), N0548_v, N0549_v, N0548_port_0, N0549_port_0);
  spice_transistor_nmos tM2559(v(clk1_v), N0723_v, N0722_v, N0723_port_2, N0722_port_1);
  spice_transistor_nmos tM2558(v(clk2_v), N0283_v, M12_v, N0283_port_1, M12_port_7);
  spice_transistor_nmos_vdd tM2809(v(N0874_v), N0846_v, N0846_port_2);
  spice_transistor_nmos tM2808(v(ACC_ADAC_v), N0870_v, N0856_v, N0870_port_0, N0856_port_1);
  spice_transistor_nmos tM1996(v(N0610_v), N0642_v, N0652_v, N0642_port_4, N0652_port_0);
  spice_transistor_nmos_gnd tM1884(v(N0466_v), N0459_v, N0459_port_4);
  spice_transistor_nmos_vdd tM1994(v(S00624_v), SC_A22_M22_CLK2_v, SC_A22_M22_CLK2_port_8);
  spice_transistor_nmos_gnd tM1995(v(N0655_v), SC_A22_M22_CLK2_v, SC_A22_M22_CLK2_port_9);
  spice_transistor_nmos_gnd tM3048(v(DCL_2_v), N0716_v, N0716_port_2);
  spice_transistor_nmos_gnd tM3049(v(N0286_v), N0728_v, N0728_port_0);
  spice_transistor_nmos tM3043(v(N0891_v), N0913_v, N0554_v, N0913_port_1, N0554_port_1);
  spice_transistor_nmos tM3040(v(ADSR_v), N0514_v, ACC_2_v, N0514_port_0, ACC_2_port_4);
  spice_transistor_nmos_vdd tM2685(v(N1007_v), OPA_0_v, OPA_0_port_13);
  spice_transistor_nmos_vdd tM2684(v(N1006_v), _OPA_0_v, _OPA_0_port_14);
  spice_transistor_nmos tM1104(v(N0381_v), N0387_v, PC0_3_v, N0387_port_2, PC0_3_port_1);
  spice_transistor_nmos_vdd tM3148(v(N0715_v), cm_ram2_v, cm_ram2_port_0);

  spice_pullup pullup_1153(N0643_v, N0643_port_2);
  spice_pullup pullup_2139(N0885_v, N0885_port_2);
  spice_pullup pullup_492(N0394_v, N0394_port_6);
  spice_pullup pullup_493(N0461_v, N0461_port_2);
  spice_pullup pullup_494(ADDR_RFSH_1_v, ADDR_RFSH_1_port_0);
  spice_pullup pullup_703(N0400_v, N0400_port_1);
  spice_pullup pullup_707(ADDR_PTR_1_v, ADDR_PTR_1_port_0);
  spice_pullup pullup_705(N0475_v, N0475_port_0);
  spice_pullup pullup_1604(N0445_v, N0445_port_2);
  spice_pullup pullup_814(S00612_v, S00612_port_1);
  spice_pullup pullup_815(S00628_v, S00628_port_0);
  spice_pullup pullup_811(N0437_v, N0437_port_0);
  spice_pullup pullup_726(N0279_v, N0279_port_0);
  spice_pullup pullup_1276(N0993_v, N0993_port_3);
  spice_pullup pullup_1274(N0995_v, N0995_port_3);
  spice_pullup pullup_1275(N0997_v, N0997_port_3);
  spice_pullup pullup_1271(N0999_v, N0999_port_3);
  spice_pullup pullup_1625(ADD_GROUP_4__v, ADD_GROUP_4__port_3);
  spice_pullup pullup_921(N0467_v, N0467_port_1);
  spice_pullup pullup_926(N0588_v, N0588_port_0);
  spice_pullup pullup_8(N0754_v, N0754_port_2);
  spice_pullup pullup_1852(N0377_v, N0377_port_1);
  spice_pullup pullup_1851(ADD_0_v, ADD_0_port_2);
  spice_pullup pullup_1294(S00678_v, S00678_port_1);
  spice_pullup pullup_1297(N0296_v, N0296_port_2);
  spice_pullup pullup_2148(S00801_v, S00801_port_1);
  spice_pullup pullup_2033(N0665_v, N0665_port_1);
  spice_pullup pullup_2036(N0349_v, N0349_port_0);
  spice_pullup pullup_2105(S00834_v, S00834_port_0);
  spice_pullup pullup_2100(N0357_v, N0357_port_0);
  spice_pullup pullup_667(N0732_v, N0732_port_2);
  spice_pullup pullup_661(N0561_v, N0561_port_0);
  spice_pullup pullup_663(N0833_v, N0833_port_2);
  spice_pullup pullup_485(N0537_v, N0537_port_10);
  spice_pullup pullup_710(N0464_v, N0464_port_3);
  spice_pullup pullup_247(N0391_v, N0391_port_6);
  spice_pullup pullup_245(N0864_v, N0864_port_2);
  spice_pullup pullup_1619(WRITE_CARRY_2__v, WRITE_CARRY_2__port_12);
  spice_pullup pullup_1784(N0856_v, N0856_port_2);
  spice_pullup pullup_1040(SC_A22_v, SC_A22_port_3);
  spice_pullup pullup_1043(SC_M22_CLK2_v, SC_M22_CLK2_port_3);
  spice_pullup pullup_1042(N0679_v, N0679_port_0);
  spice_pullup pullup_933(N0637_v, N0637_port_0);
  spice_pullup pullup_935(N0641_v, N0641_port_0);
  spice_pullup pullup_934(N0642_v, N0642_port_0);
  spice_pullup pullup_937(REG_RFSH_2_v, REG_RFSH_2_port_1);
  spice_pullup pullup_1827(N0911_v, N0911_port_2);
  spice_pullup pullup_1820(N0874_v, N0874_port_2);
  spice_pullup pullup_1829(N0878_v, N0878_port_3);
  spice_pullup pullup_1695(N0546_v, N0546_port_1);
  spice_pullup pullup_776(N0600_v, N0600_port_0);
  spice_pullup pullup_774(N0574_v, N0574_port_0);
  spice_pullup pullup_773(N0571_v, N0571_port_0);
  spice_pullup pullup_772(S00585_v, S00585_port_1);
  spice_pullup pullup_771(S00584_v, S00584_port_1);
  spice_pullup pullup_2026(S00804_v, S00804_port_0);
  spice_pullup pullup_2027(N0944_v, N0944_port_1);
  spice_pullup pullup_770(S00583_v, S00583_port_1);
  spice_pullup pullup_2023(N0917_v, N0917_port_1);
  spice_pullup pullup_674(N0300_v, N0300_port_4);
  spice_pullup pullup_672(N0307_v, N0307_port_4);
  spice_pullup pullup_779(N0610_v, N0610_port_0);
  spice_pullup pullup_2112(S00833_v, S00833_port_0);
  spice_pullup pullup_1440(N0407_v, N0407_port_2);
  spice_pullup pullup_120(N0862_v, N0862_port_2);
  spice_pullup pullup_1599(READ_ACC_3__v, READ_ACC_3__port_6);
  spice_pullup pullup_1598(INC_GROUP_5__v, INC_GROUP_5__port_3);
  spice_pullup pullup_722(N0365_v, N0365_port_2);
  spice_pullup pullup_723(N0708_v, N0708_port_2);
  spice_pullup pullup_1620(N0515_v, N0515_port_2);
  spice_pullup pullup_729(N0379_v, N0379_port_2);
  spice_pullup pullup_839(N0326_v, N0326_port_3);
  spice_pullup pullup_1135(N0352_v, N0352_port_0);
  spice_pullup pullup_2142(N0877_v, N0877_port_4);
  spice_pullup pullup_1792(N0751_v, N0751_port_0);
  spice_pullup pullup_1835(N0915_v, N0915_port_1);
  spice_pullup pullup_1168(N0992_v, N0992_port_3);
  spice_pullup pullup_1838(N0940_v, N0940_port_1);
  spice_pullup pullup_1166(N0996_v, N0996_port_0);
  spice_pullup pullup_1534(N0805_v, N0805_port_1);
  spice_pullup pullup_2231(N0664_v, N0664_port_1);
  spice_pullup pullup_1901(N0884_v, N0884_port_2);
  spice_pullup pullup_1902(N0857_v, N0857_port_2);
  spice_pullup pullup_1904(N0347_v, N0347_port_3);
  spice_pullup pullup_1908(N0875_v, N0875_port_3);
  spice_pullup pullup_1607(N0446_v, N0446_port_3);
  spice_pullup pullup_1606(CY_IB_v, CY_IB_port_2);
  spice_pullup pullup_1799(N0354_v, N0354_port_0);
  spice_pullup pullup_1798(N0802_v, N0802_port_2);
  spice_pullup pullup_2167(S00817_v, S00817_port_0);
  spice_pullup pullup_130(N0863_v, N0863_port_0);
  spice_pullup pullup_644(N0541_v, N0541_port_4);
  spice_pullup pullup_2230(N0663_v, N0663_port_1);
  spice_pullup pullup_1638(S00676_v, S00676_port_0);
  spice_pullup pullup_1639(N0671_v, N0671_port_0);
  spice_pullup pullup_1635(N1005_v, N1005_port_2);
  spice_pullup pullup_1632(N1001_v, N1001_port_2);
  spice_pullup pullup_356(N0392_v, N0392_port_6);
  spice_pullup pullup_1029(N0627_v, N0627_port_2);
  spice_pullup pullup_1028(S00627_v, S00627_port_1);
  spice_pullup pullup_1027(N0622_v, N0622_port_2);
  spice_pullup pullup_912(N0428_v, N0428_port_2);
  spice_pullup pullup_911(N0528_v, N0528_port_0);
  spice_pullup pullup_914(N0435_v, N0435_port_2);
  spice_pullup pullup_1690(N0678_v, N0678_port_0);
  spice_pullup pullup_1692(N0701_v, N0701_port_0);
  spice_pullup pullup_2227(S00836_v, S00836_port_0);
  spice_pullup pullup_1934(N0916_v, N0916_port_1);
  spice_pullup pullup_1809(N0471_v, N0471_port_0);
  spice_pullup pullup_1801(N0370_v, N0370_port_0);
  spice_pullup pullup_1803(N0378_v, N0378_port_2);
  spice_pullup pullup_1802(N0345_v, N0345_port_0);
  spice_pullup pullup_211(N0389_v, N0389_port_6);
  spice_pullup pullup_2173(S00819_v, S00819_port_0);
  spice_pullup pullup_2236(S00840_v, S00840_port_1);
  spice_pullup pullup_1278(IOR_v, IOR_port_1);
  spice_pullup pullup_109(N0385_v, N0385_port_6);
  spice_pullup pullup_214(N0390_v, N0390_port_6);
  spice_pullup pullup_589(N0938_v, N0938_port_3);
  spice_pullup pullup_925(N0460_v, N0460_port_0);
  spice_pullup pullup_1488(N0328_v, N0328_port_0);
  spice_pullup pullup_1485(N0375_v, N0375_port_3);
  spice_pullup pullup_1715(N0855_v, N0855_port_2);
  spice_pullup pullup_1487(N0337_v, N0337_port_0);
  spice_pullup pullup_1486(N0369_v, N0369_port_0);
  spice_pullup pullup_1483(__X21__CLK2__v, __X21__CLK2__port_2);
  spice_pullup pullup_1482(S00699_v, S00699_port_1);
  spice_pullup pullup_1156(SC_M12_CLK2_v, SC_M12_CLK2_port_1);
  spice_pullup pullup_1154(N0660_v, N0660_port_1);
  spice_pullup pullup_690(N0820_v, N0820_port_3);
  spice_pullup pullup_1036(N0578_v, N0578_port_2);
  spice_pullup pullup_1037(N0590_v, N0590_port_2);
  spice_pullup pullup_968(DC_v, DC_port_4);
  spice_pullup pullup_969(WRAB1_v, WRAB1_port_5);
  spice_pullup pullup_1476(N0383_v, N0383_port_2);
  spice_pullup pullup_111(N0386_v, N0386_port_6);
  spice_pullup pullup_1325(N0476_v, N0476_port_2);
  spice_pullup pullup_1327(N0419_v, N0419_port_3);
  spice_pullup pullup_1328(_SRC_v, _SRC_port_1);
  spice_pullup pullup_2216(N0668_v, N0668_port_4);
  spice_pullup pullup_2219(N0673_v, N0673_port_2);
  spice_pullup pullup_1926(S00765_v, S00765_port_0);
  spice_pullup pullup_1927(S00766_v, S00766_port_0);
  spice_pullup pullup_1925(N0672_v, N0672_port_1);
  spice_pullup pullup_2161(N0946_v, N0946_port_1);
  spice_pullup pullup_1970(N0355_v, N0355_port_0);
  spice_pullup pullup_1977(N0473_v, N0473_port_0);
  spice_pullup pullup_1811(ACC_0_v, ACC_0_port_4);
  spice_pullup pullup_70(N0764_v, N0764_port_1);
  spice_pullup pullup_1516(N0423_v, N0423_port_1);
  spice_pullup pullup_1510(N0442_v, N0442_port_1);
  spice_pullup pullup_758(N0542_v, N0542_port_4);
  spice_pullup pullup_757(N0577_v, N0577_port_6);
  spice_pullup pullup_599(N0455_v, N0455_port_4);
  spice_pullup pullup_598(N0540_v, N0540_port_1);
  spice_pullup pullup_596(N0983_v, N0983_port_3);
  spice_pullup pullup_595(N0974_v, N0974_port_3);
  spice_pullup pullup_594(N0965_v, N0965_port_3);
  spice_pullup pullup_593(N0613_v, N0613_port_0);
  spice_pullup pullup_590(N0955_v, N0955_port_3);
  spice_pullup pullup_1492(N0720_v, N0720_port_2);
  spice_pullup pullup_683(RADB0_v, RADB0_port_5);
  spice_pullup pullup_682(RADB1_v, RADB1_port_4);
  spice_pullup pullup_680(N0402_v, N0402_port_0);
  spice_pullup pullup_689(N0804_v, N0804_port_3);
  spice_pullup pullup_688(N0783_v, N0783_port_3);
  spice_pullup pullup_1003(N0524_v, N0524_port_4);
  spice_pullup pullup_1007(N0580_v, N0580_port_2);
  spice_pullup pullup_971(WRAB0_v, WRAB0_port_4);
  spice_pullup pullup_970(N0547_v, N0547_port_0);
  spice_pullup pullup_972(SC_A12_CLK2_v, SC_A12_CLK2_port_3);
  spice_pullup pullup_1311(N0456_v, N0456_port_1);
  spice_pullup pullup_1310(N0413_v, N0413_port_3);
  spice_pullup pullup_2206(S00839_v, S00839_port_1);
  spice_pullup pullup_2201(S00835_v, S00835_port_0);
  spice_pullup pullup_1953(DCL_1_v, DCL_1_port_3);
  spice_pullup pullup_2159(N0918_v, N0918_port_1);
  spice_pullup pullup_2152(N0666_v, N0666_port_2);
  spice_pullup pullup_69(N0760_v, N0760_port_1);
  spice_pullup pullup_1793(DCL_0_v, DCL_0_port_0);
  spice_pullup pullup_1797(N0403_v, N0403_port_3);
  spice_pullup pullup_1796(N0803_v, N0803_port_4);
  spice_pullup pullup_765(S00578_v, S00578_port_1);
  spice_pullup pullup_766(S00579_v, S00579_port_1);
  spice_pullup pullup_767(S00580_v, S00580_port_1);
  spice_pullup pullup_768(S00581_v, S00581_port_1);
  spice_pullup pullup_769(S00582_v, S00582_port_1);
  spice_pullup pullup_2214(N0667_v, N0667_port_2);
  spice_pullup pullup_778(REG_RFSH_0_v, REG_RFSH_0_port_1);
  spice_pullup pullup_1771(S00757_v, S00757_port_1);
  spice_pullup pullup_1770(S00761_v, S00761_port_0);
  spice_pullup pullup_1777(N0724_v, N0724_port_2);
  spice_pullup pullup_1010(N0568_v, N0568_port_1);
  spice_pullup pullup_412(N0534_v, N0534_port_10);
  spice_pullup pullup_411(N0533_v, N0533_port_10);
  spice_pullup pullup_946(__FIN_X12__v, __FIN_X12__port_2);
  spice_pullup pullup_1019(N0564_v, N0564_port_3);
  spice_pullup pullup_788(N0450_v, N0450_port_0);
  spice_pullup pullup_789(S00598_v, S00598_port_1);
  spice_pullup pullup_780(N0609_v, N0609_port_0);
  spice_pullup pullup_781(REG_RFSH_1_v, REG_RFSH_1_port_0);
  spice_pullup pullup_1737(S00732_v, S00732_port_1);
  spice_pullup pullup_1302(N0399_v, N0399_port_2);
  spice_pullup pullup_1306(N0404_v, N0404_port_2);
  spice_pullup pullup_1307(N0784_v, N0784_port_0);
  spice_pullup pullup_1304(N0432_v, N0432_port_1);
  spice_pullup pullup_1305(N0327_v, N0327_port_4);
  spice_pullup pullup_761(N0560_v, N0560_port_6);
  spice_pullup pullup_1949(N0348_v, N0348_port_2);
  spice_pullup pullup_514(N0314_v, N0314_port_1);
  spice_pullup pullup_2095(N0735_v, N0735_port_0);
  spice_pullup pullup_2092(S00825_v, S00825_port_0);
  spice_pullup pullup_2090(N0356_v, N0356_port_9);
  spice_pullup pullup_1543(N0801_v, N0801_port_1);
  spice_pullup pullup_1544(N0722_v, N0722_port_2);
  spice_pullup pullup_1478(__X31__CLK2__v, __X31__CLK2__port_1);
  spice_pullup pullup_1479(N0353_v, N0353_port_2);
  spice_pullup pullup_775(N0573_v, N0573_port_0);
  spice_pullup pullup_573(S00557_v, S00557_port_1);
  spice_pullup pullup_575(N0463_v, N0463_port_2);
  spice_pullup pullup_579(N0928_v, N0928_port_3);
  spice_pullup pullup_578(N0919_v, N0919_port_3);
  spice_pullup pullup_315(N0532_v, N0532_port_10);
  spice_pullup pullup_314(N0531_v, N0531_port_10);
  spice_pullup pullup_1162(N0994_v, N0994_port_2);
  spice_pullup pullup_1161(N0998_v, N0998_port_0);
  spice_pullup pullup_1761(N0350_v, N0350_port_0);
  spice_pullup pullup_1764(N0346_v, N0346_port_1);
  spice_pullup pullup_1366(N0398_v, N0398_port_0);
  spice_pullup pullup_950(N0608_v, N0608_port_0);
  spice_pullup pullup_798(N0318_v, N0318_port_1);
  spice_pullup pullup_791(S00600_v, S00600_port_1);
  spice_pullup pullup_790(S00599_v, S00599_port_1);
  spice_pullup pullup_792(S00601_v, S00601_port_1);
  spice_pullup pullup_794(S00613_v, S00613_port_0);
  spice_pullup pullup_2133(N0859_v, N0859_port_2);
  spice_pullup pullup_1932(N0942_v, N0942_port_1);
  spice_pullup pullup_1374(N0486_v, N0486_port_3);
  spice_pullup pullup_1791(N0766_v, N0766_port_0);
  spice_pullup pullup_1203(FIM_SRC_v, FIM_SRC_port_4);
  spice_pullup pullup_1202(JCN_v, JCN_port_4);
  spice_pullup pullup_1201(ISZ_v, ISZ_port_4);
  spice_pullup pullup_1207(JIN_FIN_v, JIN_FIN_port_8);
  spice_pullup pullup_1206(OPE_v, OPE_port_4);
  spice_pullup pullup_1205(N0493_v, N0493_port_0);
  spice_pullup pullup_1204(IO_v, IO_port_4);
  spice_pullup pullup_1209(JUN_JMS_v, JUN_JMS_port_8);
  spice_pullup pullup_1208(N0510_v, N0510_port_0);
  spice_pullup pullup_1993(N0876_v, N0876_port_2);
  spice_pullup pullup_1996(N0879_v, N0879_port_3);
  spice_pullup pullup_2088(N0474_v, N0474_port_1);
  spice_pullup pullup_1789(S00778_v, S00778_port_0);
  spice_pullup pullup_1688(N0659_v, N0659_port_4);
  spice_pullup pullup_1687(N0675_v, N0675_port_0);
  spice_pullup pullup_1686(S00716_v, S00716_port_1);
  spice_pullup pullup_40(N0758_v, N0758_port_2);
  spice_pullup pullup_42(N0763_v, N0763_port_2);
  spice_pullup pullup_546(N0395_v, N0395_port_6);
  spice_pullup pullup_540(WADB2_v, WADB2_port_4);
  spice_pullup pullup_144(N0387_v, N0387_port_6);
  spice_pullup pullup_145(N0388_v, N0388_port_6);
  spice_pullup pullup_899(CLK2_JMS_DC_M22_BBL_M22_X12_X22___v, CLK2_JMS_DC_M22_BBL_M22_X12_X22___port_3);
  spice_pullup pullup_1193(POC_v, POC_port_3);
  spice_pullup pullup_1192(N0769_v, N0769_port_0);
  spice_pullup pullup_1196(FIN_FIM_v, FIN_FIM_port_5);
  spice_pullup pullup_1755(N0704_v, N0704_port_1);
  spice_pullup pullup_1750(CY_1_v, CY_1_port_4);
  spice_pullup pullup_712(N0457_v, N0457_port_1);
  spice_pullup pullup_1194(_CN_v, _CN_port_2);
  spice_pullup pullup_1210(JCN_ISZ_v, JCN_ISZ_port_8);
  spice_pullup pullup_1211(INC_ISZ_v, INC_ISZ_port_4);
  spice_pullup pullup_1212(DCL_v, DCL_port_0);
  spice_pullup pullup_248(N0865_v, N0865_port_0);
  spice_pullup pullup_1961(N0858_v, N0858_port_2);
  spice_pullup pullup_2094(N0734_v, N0734_port_1);
  spice_pullup pullup_1614(N0502_v, N0502_port_2);
  spice_pullup pullup_1615(N0490_v, N0490_port_2);
  spice_pullup pullup_1616(ADSR_v, ADSR_port_2);
  spice_pullup pullup_2098(N0359_v, N0359_port_0);
  spice_pullup pullup_1611(S00709_v, S00709_port_1);
  spice_pullup pullup_1613(ADSL_v, ADSL_port_2);
  spice_pullup pullup_2185(N0669_v, N0669_port_3);
  spice_pullup pullup_2184(N0670_v, N0670_port_4);
  spice_pullup pullup_2187(N0674_v, N0674_port_1);
  spice_pullup pullup_2180(S00828_v, S00828_port_1);
  spice_pullup pullup_34(N0762_v, N0762_port_1);
  spice_pullup pullup_33(N0756_v, N0756_port_1);
  spice_pullup pullup_2058(S00803_v, S00803_port_1);
  spice_pullup pullup_1699(N0677_v, N0677_port_0);
  spice_pullup pullup_887(N0522_v, N0522_port_1);
  spice_pullup pullup_881(__INH__X32_CLK2_v, __INH__X32_CLK2_port_2);
  spice_pullup pullup_880(N0494_v, N0494_port_0);
  spice_pullup pullup_1180(N0368_v, N0368_port_3);
  spice_pullup pullup_1745(N0705_v, N0705_port_3);
  spice_pullup pullup_678(S00609_v, S00609_port_0);
  spice_pullup pullup_2194(N0733_v, N0733_port_1);
  spice_pullup pullup_2195(N0736_v, N0736_port_0);
  spice_pullup pullup_27(S00536_v, S00536_port_1);
  spice_pullup pullup_24(S00531_v, S00531_port_0);
  spice_pullup pullup_2038(N0728_v, N0728_port_2);
  spice_pullup pullup_1365(N0487_v, N0487_port_2);
  spice_pullup pullup_670(RADB2_v, RADB2_port_4);
  spice_pullup pullup_603(N0503_v, N0503_port_1);
  spice_pullup pullup_2040(DCL_2_v, DCL_2_port_2);
  spice_pullup pullup_2041(N0749_v, N0749_port_0);
  spice_pullup pullup_2047(S00814_v, S00814_port_0);
  spice_pullup pullup_1800(N0363_v, N0363_port_0);
  spice_pullup pullup_526(N0316_v, N0316_port_1);
  spice_pullup pullup_527(N0711_v, N0711_port_1);
  spice_pullup pullup_521(WADB1_v, WADB1_port_4);
  spice_pullup pullup_1420(N0797_v, N0797_port_2);
  spice_pullup pullup_1425(S00710_v, S00710_port_0);
  spice_pullup pullup_822(N0451_v, N0451_port_0);
  spice_pullup pullup_1736(S00734_v, S00734_port_1);
  spice_pullup pullup_1735(ADC_CY_v, ADC_CY_port_3);
  spice_pullup pullup_1733(ADD_ACC_v, ADD_ACC_port_2);
  spice_pullup pullup_524(WADB0_v, WADB0_port_4);
  spice_pullup pullup_450(N0469_v, N0469_port_1);
  spice_pullup pullup_1648(N1003_v, N1003_port_2);
  spice_pullup pullup_858(N0511_v, N0511_port_0);
  spice_pullup pullup_853(N0443_v, N0443_port_1);
  spice_pullup pullup_850(S00654_v, S00654_port_1);
  spice_pullup pullup_856(_INH_v, _INH_port_0);
  spice_pullup pullup_857(INH_v, INH_port_2);
  spice_pullup pullup_854(N0447_v, N0447_port_3);
  spice_pullup pullup_1238(N0636_v, N0636_port_5);
  spice_pullup pullup_1239(INC_ISZ_ADD_SUB_XCH_LD_v, INC_ISZ_ADD_SUB_XCH_LD_port_5);
  spice_pullup pullup_1232(KBP_v, KBP_port_0);
  spice_pullup pullup_1233(TCS_v, TCS_port_0);
  spice_pullup pullup_1231(O_IB_v, O_IB_port_0);
  spice_pullup pullup_1236(BBL_v, BBL_port_5);
  spice_pullup pullup_1237(JMS_v, JMS_port_5);
  spice_pullup pullup_1234(DAA_v, DAA_port_0);
  spice_pullup pullup_1235(XCH_v, XCH_port_4);
  spice_pullup pullup_1965(N0750_v, N0750_port_1);
  spice_pullup pullup_1508(N0351_v, N0351_port_2);
  spice_pullup pullup_10(N0761_v, N0761_port_2);
  spice_pullup pullup_983(S00624_v, S00624_port_1);
  spice_pullup pullup_2074(S00818_v, S00818_port_0);
  spice_pullup pullup_2077(N0288_v, N0288_port_8);
  spice_pullup pullup_2076(N0366_v, N0366_port_0);
  spice_pullup pullup_2071(N0730_v, N0730_port_2);
  spice_pullup pullup_1430(N0718_v, N0718_port_2);
  spice_pullup pullup_1436(S00725_v, S00725_port_0);
  spice_pullup pullup_997(S00620_v, S00620_port_1);
  spice_pullup pullup_996(N0655_v, N0655_port_1);
  spice_pullup pullup_995(N0649_v, N0649_port_1);
  spice_pullup pullup_448(N0393_v, N0393_port_6);
  spice_pullup pullup_1658(S00689_v, S00689_port_0);
  spice_pullup pullup_1659(S00687_v, S00687_port_0);
  spice_pullup pullup_1654(N1007_v, N1007_port_2);
  spice_pullup pullup_847(N0322_v, N0322_port_4);
  spice_pullup pullup_846(N0310_v, N0310_port_4);
  spice_pullup pullup_1018(N0603_v, N0603_port_2);
  spice_pullup pullup_1248(FIN_FIM_SRC_JIN_v, FIN_FIM_SRC_JIN_port_6);
  spice_pullup pullup_1247(LD_v, LD_port_4);
  spice_pullup pullup_1246(INC_ISZ_XCH_v, INC_ISZ_XCH_port_5);
  spice_pullup pullup_1245(STC_v, STC_port_0);
  spice_pullup pullup_1244(TCC_v, TCC_port_0);
  spice_pullup pullup_1243(CMA_v, CMA_port_0);
  spice_pullup pullup_1242(RAL_v, RAL_port_0);
  spice_pullup pullup_1241(RAR_v, RAR_port_0);
  spice_pullup pullup_1240(IOW_v, IOW_port_0);
  spice_pullup pullup_1967(S00800_v, S00800_port_0);
  spice_pullup pullup_1886(N0364_v, N0364_port_0);
  spice_pullup pullup_1399(S00685_v, S00685_port_0);
  spice_pullup pullup_1391(S00690_v, S00690_port_1);
  spice_pullup pullup_1869(S00767_v, S00767_port_0);
  spice_pullup pullup_1867(S00764_v, S00764_port_1);
  spice_pullup pullup_1864(N0371_v, N0371_port_0);
  spice_pullup pullup_2067(N0358_v, N0358_port_5);
  spice_pullup pullup_1533(S00731_v, S00731_port_1);
  spice_pullup pullup_1535(N0853_v, N0853_port_0);
  spice_pullup pullup_1537(N0421_v, N0421_port_0);
  spice_pullup pullup_1309(N0329_v, N0329_port_0);
  spice_pullup pullup_501(N0453_v, N0453_port_1);
  spice_pullup pullup_503(N0902_v, N0902_port_2);
  spice_pullup pullup_746(N0401_v, N0401_port_3);
  spice_pullup pullup_740(N0304_v, N0304_port_1);
  spice_pullup pullup_618(N0737_v, N0737_port_1);
  spice_pullup pullup_1669(N1000_v, N1000_port_4);
  spice_pullup pullup_1258(CLB_v, CLB_port_0);
  spice_pullup pullup_1259(SBM_v, SBM_port_0);
  spice_pullup pullup_1254(SUB_v, SUB_port_4);
  spice_pullup pullup_1255(ADD_v, ADD_port_4);
  spice_pullup pullup_1256(LDM_BBL_v, LDM_BBL_port_3);
  spice_pullup pullup_1257(JUN2_JMS2_v, JUN2_JMS2_port_3);
  spice_pullup pullup_1250(CMC_v, CMC_port_0);
  spice_pullup pullup_1251(DAC_v, DAC_port_0);
  spice_pullup pullup_1252(IAC_v, IAC_port_0);
  spice_pullup pullup_1253(CLC_v, CLC_port_0);
  spice_pullup pullup_1092(N0630_v, N0630_port_2);
  spice_pullup pullup_1091(N0682_v, N0682_port_4);
  spice_pullup pullup_1897(N0964_v, N0964_port_2);
  spice_pullup pullup_1895(S00762_v, S00762_port_1);
  spice_pullup pullup_1890(N0726_v, N0726_port_2);
  spice_pullup pullup_1389(N0799_v, N0799_port_0);
  spice_pullup pullup_1876(N0472_v, N0472_port_1);
  spice_pullup pullup_2015(N0913_v, N0913_port_2);
  spice_pullup pullup_2014(S00781_v, S00781_port_1);
  spice_pullup pullup_1524(N0340_v, N0340_port_0);
  spice_pullup pullup_1523(N0430_v, N0430_port_0);
  spice_pullup pullup_1521(S00740_v, S00740_port_0);
  spice_pullup pullup_1150(L_v, L_port_2);
  spice_pullup pullup_600(ADDR_RFSH_0_v, ADDR_RFSH_0_port_0);
  spice_pullup pullup_604(S00564_v, S00564_port_0);
  spice_pullup pullup_1708(N0470_v, N0470_port_2);
  spice_pullup pullup_1702(S00729_v, S00729_port_1);
  spice_pullup pullup_1703(S00724_v, S00724_port_1);
  spice_pullup pullup_464(N0536_v, N0536_port_10);
  spice_pullup pullup_463(N0535_v, N0535_port_10);
  spice_pullup pullup_1672(N1004_v, N1004_port_4);
  spice_pullup pullup_1673(N1002_v, N1002_port_4);
  spice_pullup pullup_1671(WRITE_ACC_1__v, WRITE_ACC_1__port_15);
  spice_pullup pullup_1674(N1006_v, N1006_port_4);
  spice_pullup pullup_1678(N0658_v, N0658_port_3);
  spice_pullup pullup_863(ADDR_PTR_0_v, ADDR_PTR_0_port_2);
  spice_pullup pullup_860(N0466_v, N0466_port_2);
  spice_pullup pullup_867(N0505_v, N0505_port_1);
  spice_pullup pullup_865(N0459_v, N0459_port_5);
  spice_pullup pullup_1260(ADM_v, ADM_port_0);
  spice_pullup pullup_1063(N0361_v, N0361_port_0);
  spice_pullup pullup_488(N0538_v, N0538_port_10);
  spice_pullup pullup_550(N0396_v, N0396_port_6);
  spice_pullup pullup_1283(N0480_v, N0480_port_1);
  spice_pullup pullup_1281(N0477_v, N0477_port_0);
  spice_pullup pullup_1285(N0479_v, N0479_port_0);




  spice_node_2 n_N0556(eclk, ereset, N0556_port_2,N0556_port_1, N0556_v);
  spice_node_1 n_S00819(eclk, ereset, S00819_port_0, S00819_v);
  spice_node_3 n_CY_ADA(eclk, ereset, CY_ADA_port_2,CY_ADA_port_3,CY_ADA_port_0, CY_ADA_v);
  spice_node_5 n_N0449(eclk, ereset, N0449_port_3,N0449_port_1,N0449_port_6,N0449_port_4,N0449_port_5, N0449_v);
  spice_node_4 n_N0448(eclk, ereset, N0448_port_2,N0448_port_3,N0448_port_0,N0448_port_1, N0448_v);
  spice_node_2 n_N0443(eclk, ereset, N0443_port_2,N0443_port_1, N0443_v);
  spice_node_2 n_N0442(eclk, ereset, N0442_port_0,N0442_port_1, N0442_v);
  spice_node_2 n_N0441(eclk, ereset, N0441_port_0,N0441_port_1, N0441_v);
  spice_node_3 n_N0440(eclk, ereset, N0440_port_3,N0440_port_4,N0440_port_5, N0440_v);
  spice_node_3 n_N0447(eclk, ereset, N0447_port_2,N0447_port_3,N0447_port_1, N0447_v);
  spice_node_2 n_N0446(eclk, ereset, N0446_port_2,N0446_port_3, N0446_v);
  spice_node_2 n_N0445(eclk, ereset, N0445_port_2,N0445_port_1, N0445_v);
  spice_node_2 n_N0444(eclk, ereset, N0444_port_12,N0444_port_13, N0444_v);
  spice_node_2 n_N0991(eclk, ereset, N0991_port_0,N0991_port_1, N0991_v);
  spice_node_2 n_N0990(eclk, ereset, N0990_port_0,N0990_port_1, N0990_v);
  spice_node_2 n_N0993(eclk, ereset, N0993_port_2,N0993_port_3, N0993_v);
  spice_node_2 n_N0992(eclk, ereset, N0992_port_2,N0992_port_3, N0992_v);
  spice_node_2 n_N0995(eclk, ereset, N0995_port_2,N0995_port_3, N0995_v);
  spice_node_2 n_N0994(eclk, ereset, N0994_port_2,N0994_port_3, N0994_v);
  spice_node_2 n_N0997(eclk, ereset, N0997_port_3,N0997_port_1, N0997_v);
  spice_node_2 n_N0999(eclk, ereset, N0999_port_2,N0999_port_3, N0999_v);
  spice_node_2 n_N0998(eclk, ereset, N0998_port_0,N0998_port_1, N0998_v);
  spice_node_10 n_N0883(eclk, ereset, N0883_port_8,N0883_port_9,N0883_port_2,N0883_port_3,N0883_port_0,N0883_port_6,N0883_port_7,N0883_port_4,N0883_port_5,N0883_port_10, N0883_v);
  spice_node_10 n_N0880(eclk, ereset, N0880_port_8,N0880_port_9,N0880_port_2,N0880_port_3,N0880_port_0,N0880_port_6,N0880_port_7,N0880_port_4,N0880_port_5,N0880_port_10, N0880_v);
  spice_node_2 n_N0887(eclk, ereset, N0887_port_3,N0887_port_5, N0887_v);
  spice_node_2 n_N0886(eclk, ereset, N0886_port_0,N0886_port_1, N0886_v);
  spice_node_2 n_N0530(eclk, ereset, N0530_port_3,N0530_port_4, N0530_v);
  spice_node_11 n_N0536(eclk, ereset, N0536_port_8,N0536_port_9,N0536_port_2,N0536_port_3,N0536_port_0,N0536_port_1,N0536_port_6,N0536_port_7,N0536_port_4,N0536_port_5,N0536_port_10, N0536_v);
  spice_node_11 n_N0535(eclk, ereset, N0535_port_8,N0535_port_9,N0535_port_2,N0535_port_3,N0535_port_0,N0535_port_1,N0535_port_6,N0535_port_7,N0535_port_4,N0535_port_5,N0535_port_10, N0535_v);
  spice_node_11 n_N0534(eclk, ereset, N0534_port_8,N0534_port_9,N0534_port_2,N0534_port_3,N0534_port_0,N0534_port_1,N0534_port_6,N0534_port_7,N0534_port_4,N0534_port_5,N0534_port_10, N0534_v);
  spice_node_4 n_N0539(eclk, ereset, N0539_port_2,N0539_port_3,N0539_port_0,N0539_port_1, N0539_v);
  spice_node_11 n_N0538(eclk, ereset, N0538_port_8,N0538_port_9,N0538_port_2,N0538_port_3,N0538_port_0,N0538_port_1,N0538_port_6,N0538_port_7,N0538_port_4,N0538_port_5,N0538_port_10, N0538_v);
  spice_node_1 n_S00579(eclk, ereset, S00579_port_1, S00579_v);
  spice_node_1 n_S00578(eclk, ereset, S00578_port_1, S00578_v);
  spice_node_2 n_N0939(eclk, ereset, N0939_port_3,N0939_port_4, N0939_v);
  spice_node_2 n_N0418(eclk, ereset, N0418_port_0,N0418_port_1, N0418_v);
  spice_node_1 n_S00757(eclk, ereset, S00757_port_1, S00757_v);
  spice_node_2 n_N0528(eclk, ereset, N0528_port_0,N0528_port_1, N0528_v);
  spice_node_5 n_INC_ISZ(eclk, ereset, INC_ISZ_port_2,INC_ISZ_port_3,INC_ISZ_port_0,INC_ISZ_port_1,INC_ISZ_port_4, INC_ISZ_v);
  spice_node_5 n_LD(eclk, ereset, LD_port_2,LD_port_3,LD_port_0,LD_port_1,LD_port_4, LD_v);
  spice_node_3 n_N0331(eclk, ereset, N0331_port_2,N0331_port_0,N0331_port_1, N0331_v);
  spice_node_1 n_S00817(eclk, ereset, S00817_port_0, S00817_v);
  spice_node_2 n_N0330(eclk, ereset, N0330_port_0,N0330_port_1, N0330_v);
  spice_node_5 n_SUB_GROUP_6_(eclk, ereset, SUB_GROUP_6__port_2,SUB_GROUP_6__port_3,SUB_GROUP_6__port_0,SUB_GROUP_6__port_1,SUB_GROUP_6__port_6, SUB_GROUP_6__v);
  spice_node_2 n_N0525(eclk, ereset, N0525_port_0,N0525_port_1, N0525_v);
  spice_node_5 n_INC_ISZ_XCH(eclk, ereset, INC_ISZ_XCH_port_2,INC_ISZ_XCH_port_3,INC_ISZ_XCH_port_1,INC_ISZ_XCH_port_4,INC_ISZ_XCH_port_5, INC_ISZ_XCH_v);
  spice_node_1 n_R8_3(eclk, ereset, R8_3_port_1, R8_3_v);
  spice_node_1 n_R8_2(eclk, ereset, R8_2_port_0, R8_2_v);
  spice_node_1 n_R8_1(eclk, ereset, R8_1_port_1, R8_1_v);
  spice_node_1 n_R8_0(eclk, ereset, R8_0_port_0, R8_0_v);
  spice_node_3 n_N0668(eclk, ereset, N0668_port_3,N0668_port_0,N0668_port_4, N0668_v);
  spice_node_4 n_N0332(eclk, ereset, N0332_port_2,N0332_port_0,N0332_port_1,N0332_port_5, N0332_v);
  spice_node_2 n_N0527(eclk, ereset, N0527_port_0,N0527_port_1, N0527_v);
  spice_node_2 n_N0335(eclk, ereset, N0335_port_0,N0335_port_1, N0335_v);
  spice_node_3 n__TMP_1(eclk, ereset, _TMP_1_port_2,_TMP_1_port_0,_TMP_1_port_1, _TMP_1_v);
  spice_node_3 n__TMP_0(eclk, ereset, _TMP_0_port_2,_TMP_0_port_0,_TMP_0_port_1, _TMP_0_v);
  spice_node_3 n__TMP_3(eclk, ereset, _TMP_3_port_2,_TMP_3_port_0,_TMP_3_port_1, _TMP_3_v);
  spice_node_3 n__TMP_2(eclk, ereset, _TMP_2_port_2,_TMP_2_port_0,_TMP_2_port_1, _TMP_2_v);
  spice_node_3 n_N0337(eclk, ereset, N0337_port_2,N0337_port_0,N0337_port_1, N0337_v);
  spice_node_3 n_TMP_3(eclk, ereset, TMP_3_port_2,TMP_3_port_0,TMP_3_port_1, TMP_3_v);
  spice_node_3 n_TMP_2(eclk, ereset, TMP_2_port_2,TMP_2_port_0,TMP_2_port_1, TMP_2_v);
  spice_node_3 n_TMP_1(eclk, ereset, TMP_1_port_2,TMP_1_port_0,TMP_1_port_1, TMP_1_v);
  spice_node_3 n_TMP_0(eclk, ereset, TMP_0_port_2,TMP_0_port_0,TMP_0_port_1, TMP_0_v);
  spice_node_5 n_JIN_FIN(eclk, ereset, JIN_FIN_port_8,JIN_FIN_port_6,JIN_FIN_port_7,JIN_FIN_port_4,JIN_FIN_port_5, JIN_FIN_v);
  spice_node_2 n_N0336(eclk, ereset, N0336_port_0,N0336_port_1, N0336_v);
  spice_node_4 n_N0523(eclk, ereset, N0523_port_2,N0523_port_3,N0523_port_0,N0523_port_1, N0523_v);
  spice_node_1 n_N0454(eclk, ereset, N0454_port_0, N0454_v);
  spice_node_3 n_N0455(eclk, ereset, N0455_port_3,N0455_port_6,N0455_port_4, N0455_v);
  spice_node_2 n_N0456(eclk, ereset, N0456_port_0,N0456_port_1, N0456_v);
  spice_node_3 n_N0457(eclk, ereset, N0457_port_2,N0457_port_0,N0457_port_1, N0457_v);
  spice_node_2 n_N0450(eclk, ereset, N0450_port_2,N0450_port_0, N0450_v);
  spice_node_2 n_N0451(eclk, ereset, N0451_port_2,N0451_port_0, N0451_v);
  spice_node_1 n_N0452(eclk, ereset, N0452_port_1, N0452_v);
  spice_node_3 n_N0453(eclk, ereset, N0453_port_2,N0453_port_0,N0453_port_1, N0453_v);
  spice_node_1 n_N0458(eclk, ereset, N0458_port_0, N0458_v);
  spice_node_3 n_N0459(eclk, ereset, N0459_port_6,N0459_port_4,N0459_port_5, N0459_v);
  spice_node_5 n_JCN_ISZ(eclk, ereset, JCN_ISZ_port_8,JCN_ISZ_port_3,JCN_ISZ_port_6,JCN_ISZ_port_7,JCN_ISZ_port_5, JCN_ISZ_v);
  spice_node_1 n_R3_0(eclk, ereset, R3_0_port_1, R3_0_v);
  spice_node_1 n_R3_1(eclk, ereset, R3_1_port_0, R3_1_v);
  spice_node_1 n_R3_3(eclk, ereset, R3_3_port_0, R3_3_v);
  spice_node_4 n_LDM_BBL(eclk, ereset, LDM_BBL_port_2,LDM_BBL_port_3,LDM_BBL_port_0,LDM_BBL_port_1, LDM_BBL_v);
  spice_node_2 n_N0982(eclk, ereset, N0982_port_0,N0982_port_1, N0982_v);
  spice_node_2 n_N0983(eclk, ereset, N0983_port_2,N0983_port_3, N0983_v);
  spice_node_2 n_N0980(eclk, ereset, N0980_port_0,N0980_port_1, N0980_v);
  spice_node_2 n_N0981(eclk, ereset, N0981_port_0,N0981_port_1, N0981_v);
  spice_node_2 n_N0986(eclk, ereset, N0986_port_0,N0986_port_1, N0986_v);
  spice_node_2 n_N0987(eclk, ereset, N0987_port_0,N0987_port_1, N0987_v);
  spice_node_2 n_N0984(eclk, ereset, N0984_port_0,N0984_port_1, N0984_v);
  spice_node_2 n_N0985(eclk, ereset, N0985_port_0,N0985_port_1, N0985_v);
  spice_node_1 n_R1_2(eclk, ereset, R1_2_port_1, R1_2_v);
  spice_node_1 n_R1_3(eclk, ereset, R1_3_port_0, R1_3_v);
  spice_node_2 n_N0988(eclk, ereset, N0988_port_0,N0988_port_1, N0988_v);
  spice_node_2 n_N0989(eclk, ereset, N0989_port_0,N0989_port_1, N0989_v);
  spice_node_7 n_N0366(eclk, ereset, N0366_port_2,N0366_port_3,N0366_port_0,N0366_port_1,N0366_port_6,N0366_port_4,N0366_port_5, N0366_v);
  spice_node_4 n_RRAB0(eclk, ereset, RRAB0_port_6,RRAB0_port_7,RRAB0_port_4,RRAB0_port_5, RRAB0_v);
  spice_node_4 n_RRAB1(eclk, ereset, RRAB1_port_6,RRAB1_port_7,RRAB1_port_4,RRAB1_port_5, RRAB1_v);
  spice_node_3 n_N0872(eclk, ereset, N0872_port_3,N0872_port_0,N0872_port_5, N0872_v);
  spice_node_1 n_R7_0(eclk, ereset, R7_0_port_1, R7_0_v);
  spice_node_1 n_R7_1(eclk, ereset, R7_1_port_0, R7_1_v);
  spice_node_1 n_R7_2(eclk, ereset, R7_2_port_1, R7_2_v);
  spice_node_1 n_R7_3(eclk, ereset, R7_3_port_0, R7_3_v);
  spice_node_1 n_S00699(eclk, ereset, S00699_port_1, S00699_v);
  spice_node_2 n_N0902(eclk, ereset, N0902_port_2,N0902_port_3, N0902_v);
  spice_node_1 n_R5_2(eclk, ereset, R5_2_port_1, R5_2_v);
  spice_node_1 n_R5_0(eclk, ereset, R5_0_port_1, R5_0_v);
  spice_node_4 n_N0524(eclk, ereset, N0524_port_2,N0524_port_3,N0524_port_1,N0524_port_4, N0524_v);
  spice_node_3 n_N0526(eclk, ereset, N0526_port_2,N0526_port_0,N0526_port_1, N0526_v);
  spice_node_2 n_N0522(eclk, ereset, N0522_port_2,N0522_port_1, N0522_v);
  spice_node_5 n_BBL(eclk, ereset, BBL_port_2,BBL_port_3,BBL_port_1,BBL_port_4,BBL_port_5, BBL_v);
  spice_node_2 n_N0906(eclk, ereset, N0906_port_0,N0906_port_1, N0906_v);
  spice_node_2 n__OPR_1(eclk, ereset, _OPR_1_port_15,_OPR_1_port_16, _OPR_1_v);
  spice_node_2 n_N0964(eclk, ereset, N0964_port_2,N0964_port_1, N0964_v);
  spice_node_2 n__OPR_0(eclk, ereset, _OPR_0_port_10,_OPR_0_port_11, _OPR_0_v);
  spice_node_2 n_POC(eclk, ereset, POC_port_3,POC_port_4, POC_v);
  spice_node_2 n_N0650(eclk, ereset, N0650_port_0,N0650_port_1, N0650_v);
  spice_node_6 n_N0357(eclk, ereset, N0357_port_2,N0357_port_3,N0357_port_0,N0357_port_1,N0357_port_4,N0357_port_5, N0357_v);
  spice_node_2 n_N0996(eclk, ereset, N0996_port_2,N0996_port_0, N0996_v);
  spice_node_2 n_cm_rom(eclk, ereset, cm_rom_port_0,cm_rom_port_1, cm_rom_v);
  spice_node_2 n_N0585(eclk, ereset, N0585_port_0,N0585_port_1, N0585_v);
  spice_node_2 n_cm_ram0(eclk, ereset, cm_ram0_port_0,cm_ram0_port_1, cm_ram0_v);
  spice_node_2 n_N0344(eclk, ereset, N0344_port_2,N0344_port_0, N0344_v);
  spice_node_5 n_d2(eclk, ereset, d2_port_2,d2_port_0,d2_port_1,d2_port_4,d2_port_5, d2_v);
  spice_node_5 n_d3(eclk, ereset, d3_port_2,d3_port_0,d3_port_1,d3_port_4,d3_port_5, d3_v);
  spice_node_2 n_WRAB1(eclk, ereset, WRAB1_port_4,WRAB1_port_5, WRAB1_v);
  spice_node_2 n_WRAB0(eclk, ereset, WRAB0_port_4,WRAB0_port_5, WRAB0_v);
  spice_node_6 n_DCL(eclk, ereset, DCL_port_2,DCL_port_3,DCL_port_0,DCL_port_1,DCL_port_4,DCL_port_5, DCL_v);
  spice_node_3 n_N0348(eclk, ereset, N0348_port_2,N0348_port_1,N0348_port_5, N0348_v);
  spice_node_2 n_N0349(eclk, ereset, N0349_port_2,N0349_port_0, N0349_v);
  spice_node_2 n_N0617(eclk, ereset, N0617_port_2,N0617_port_1, N0617_v);
  spice_node_6 n_KBP(eclk, ereset, KBP_port_2,KBP_port_3,KBP_port_0,KBP_port_1,KBP_port_4,KBP_port_5, KBP_v);
  spice_node_1 n_N0615(eclk, ereset, N0615_port_1, N0615_v);
  spice_node_2 n_N0612(eclk, ereset, N0612_port_0,N0612_port_1, N0612_v);
  spice_node_3 n_N0610(eclk, ereset, N0610_port_3,N0610_port_0,N0610_port_4, N0610_v);
  spice_node_2 n_N0611(eclk, ereset, N0611_port_0,N0611_port_1, N0611_v);
  spice_node_2 n_N0834(eclk, ereset, N0834_port_0,N0834_port_1, N0834_v);
  spice_node_3 n_ACC_ADA(eclk, ereset, ACC_ADA_port_0,ACC_ADA_port_1,ACC_ADA_port_5, ACC_ADA_v);
  spice_node_10 n___POC__CLK2_SC_A32_X12_(eclk, ereset, __POC__CLK2_SC_A32_X12__port_8,__POC__CLK2_SC_A32_X12__port_9,__POC__CLK2_SC_A32_X12__port_2,__POC__CLK2_SC_A32_X12__port_3,__POC__CLK2_SC_A32_X12__port_0,__POC__CLK2_SC_A32_X12__port_1,__POC__CLK2_SC_A32_X12__port_6,__POC__CLK2_SC_A32_X12__port_7,__POC__CLK2_SC_A32_X12__port_4,__POC__CLK2_SC_A32_X12__port_5, __POC__CLK2_SC_A32_X12__v);
  spice_node_2 n_N0341(eclk, ereset, N0341_port_0,N0341_port_1, N0341_v);
  spice_node_2 n_N0342(eclk, ereset, N0342_port_0,N0342_port_1, N0342_v);
  spice_node_1 n_PC0_9(eclk, ereset, PC0_9_port_1, PC0_9_v);
  spice_node_1 n_PC0_8(eclk, ereset, PC0_8_port_0, PC0_8_v);
  spice_node_3 n_RADB2(eclk, ereset, RADB2_port_6,RADB2_port_4,RADB2_port_5, RADB2_v);
  spice_node_3 n_RADB0(eclk, ereset, RADB0_port_6,RADB0_port_4,RADB0_port_5, RADB0_v);
  spice_node_3 n_RADB1(eclk, ereset, RADB1_port_6,RADB1_port_4,RADB1_port_5, RADB1_v);
  spice_node_1 n_PC0_1(eclk, ereset, PC0_1_port_1, PC0_1_v);
  spice_node_1 n_PC0_0(eclk, ereset, PC0_0_port_0, PC0_0_v);
  spice_node_1 n_PC0_3(eclk, ereset, PC0_3_port_1, PC0_3_v);
  spice_node_1 n_PC0_2(eclk, ereset, PC0_2_port_0, PC0_2_v);
  spice_node_1 n_PC0_5(eclk, ereset, PC0_5_port_0, PC0_5_v);
  spice_node_1 n_PC0_4(eclk, ereset, PC0_4_port_1, PC0_4_v);
  spice_node_1 n_PC0_7(eclk, ereset, PC0_7_port_0, PC0_7_v);
  spice_node_1 n_PC0_6(eclk, ereset, PC0_6_port_1, PC0_6_v);
  spice_node_3 n_N0421(eclk, ereset, N0421_port_2,N0421_port_0,N0421_port_1, N0421_v);
  spice_node_2 n_N0420(eclk, ereset, N0420_port_3,N0420_port_4, N0420_v);
  spice_node_2 n_N0423(eclk, ereset, N0423_port_0,N0423_port_1, N0423_v);
  spice_node_1 n_N0422(eclk, ereset, N0422_port_0, N0422_v);
  spice_node_1 n_N0425(eclk, ereset, N0425_port_0, N0425_v);
  spice_node_2 n_N0424(eclk, ereset, N0424_port_12,N0424_port_13, N0424_v);
  spice_node_3 n_N0427(eclk, ereset, N0427_port_3,N0427_port_4,N0427_port_5, N0427_v);
  spice_node_2 n_N0426(eclk, ereset, N0426_port_12,N0426_port_13, N0426_v);
  spice_node_2 n_N0429(eclk, ereset, N0429_port_0,N0429_port_1, N0429_v);
  spice_node_4 n_N0428(eclk, ereset, N0428_port_2,N0428_port_3,N0428_port_0,N0428_port_1, N0428_v);
  spice_node_1 n_N0343(eclk, ereset, N0343_port_2, N0343_v);
  spice_node_1 n_S00582(eclk, ereset, S00582_port_1, S00582_v);
  spice_node_1 n_S00583(eclk, ereset, S00583_port_1, S00583_v);
  spice_node_3 n_O_IB(eclk, ereset, O_IB_port_2,O_IB_port_0,O_IB_port_1, O_IB_v);
  spice_node_14 n_WRITE_CARRY_2_(eclk, ereset, WRITE_CARRY_2__port_8,WRITE_CARRY_2__port_9,WRITE_CARRY_2__port_2,WRITE_CARRY_2__port_3,WRITE_CARRY_2__port_0,WRITE_CARRY_2__port_1,WRITE_CARRY_2__port_6,WRITE_CARRY_2__port_7,WRITE_CARRY_2__port_4,WRITE_CARRY_2__port_5,WRITE_CARRY_2__port_10,WRITE_CARRY_2__port_11,WRITE_CARRY_2__port_12,WRITE_CARRY_2__port_13, WRITE_CARRY_2__v);
  spice_node_1 n_N0739(eclk, ereset, N0739_port_0, N0739_v);
  spice_node_2 n_N0738(eclk, ereset, N0738_port_3,N0738_port_0, N0738_v);
  spice_node_2 n_N0735(eclk, ereset, N0735_port_0,N0735_port_1, N0735_v);
  spice_node_2 n_N0734(eclk, ereset, N0734_port_0,N0734_port_1, N0734_v);
  spice_node_2 n_N0737(eclk, ereset, N0737_port_2,N0737_port_1, N0737_v);
  spice_node_2 n_N0736(eclk, ereset, N0736_port_0,N0736_port_1, N0736_v);
  spice_node_1 n_N0731(eclk, ereset, N0731_port_2, N0731_v);
  spice_node_3 n_N0730(eclk, ereset, N0730_port_2,N0730_port_0,N0730_port_1, N0730_v);
  spice_node_2 n_N0733(eclk, ereset, N0733_port_0,N0733_port_1, N0733_v);
  spice_node_2 n_N0732(eclk, ereset, N0732_port_2,N0732_port_1, N0732_v);
  spice_node_2 n_N0956(eclk, ereset, N0956_port_0,N0956_port_1, N0956_v);
  spice_node_2 n_N0951(eclk, ereset, N0951_port_0,N0951_port_1, N0951_v);
  spice_node_2 n_N0950(eclk, ereset, N0950_port_0,N0950_port_1, N0950_v);
  spice_node_2 n_N0953(eclk, ereset, N0953_port_0,N0953_port_1, N0953_v);
  spice_node_2 n_N0952(eclk, ereset, N0952_port_0,N0952_port_1, N0952_v);
  spice_node_2 n_N0959(eclk, ereset, N0959_port_0,N0959_port_1, N0959_v);
  spice_node_2 n_N0958(eclk, ereset, N0958_port_0,N0958_port_1, N0958_v);
  spice_node_5 n_CY(eclk, ereset, CY_port_2,CY_port_3,CY_port_0,CY_port_1,CY_port_5, CY_v);
  spice_node_1 n_S00685(eclk, ereset, S00685_port_0, S00685_v);
  spice_node_1 n_S00687(eclk, ereset, S00687_port_0, S00687_v);
  spice_node_1 n_S00689(eclk, ereset, S00689_port_0, S00689_v);
  spice_node_2 n_N0559(eclk, ereset, N0559_port_2,N0559_port_1, N0559_v);
  spice_node_3 n_N0558(eclk, ereset, N0558_port_2,N0558_port_0,N0558_port_1, N0558_v);
  spice_node_10 n_N0882(eclk, ereset, N0882_port_8,N0882_port_9,N0882_port_2,N0882_port_3,N0882_port_1,N0882_port_6,N0882_port_7,N0882_port_4,N0882_port_5,N0882_port_10, N0882_v);
  spice_node_10 n_N0881(eclk, ereset, N0881_port_8,N0881_port_9,N0881_port_2,N0881_port_3,N0881_port_0,N0881_port_6,N0881_port_7,N0881_port_4,N0881_port_5,N0881_port_10, N0881_v);
  spice_node_1 n_S00731(eclk, ereset, S00731_port_1, S00731_v);
  spice_node_1 n_N0397(eclk, ereset, N0397_port_2, N0397_v);
  spice_node_11 n_N0533(eclk, ereset, N0533_port_8,N0533_port_9,N0533_port_2,N0533_port_3,N0533_port_0,N0533_port_1,N0533_port_6,N0533_port_7,N0533_port_4,N0533_port_5,N0533_port_10, N0533_v);
  spice_node_3 n_N0383(eclk, ereset, N0383_port_2,N0383_port_0,N0383_port_1, N0383_v);
  spice_node_11 n_N0532(eclk, ereset, N0532_port_8,N0532_port_9,N0532_port_2,N0532_port_3,N0532_port_0,N0532_port_1,N0532_port_6,N0532_port_7,N0532_port_4,N0532_port_5,N0532_port_10, N0532_v);
  spice_node_11 n_N0531(eclk, ereset, N0531_port_8,N0531_port_9,N0531_port_2,N0531_port_3,N0531_port_0,N0531_port_1,N0531_port_6,N0531_port_7,N0531_port_4,N0531_port_5,N0531_port_10, N0531_v);
  spice_node_11 n_N0537(eclk, ereset, N0537_port_8,N0537_port_9,N0537_port_2,N0537_port_3,N0537_port_0,N0537_port_1,N0537_port_6,N0537_port_7,N0537_port_4,N0537_port_5,N0537_port_10, N0537_v);
  spice_node_1 n_S00836(eclk, ereset, S00836_port_0, S00836_v);
  spice_node_3 n_N0641(eclk, ereset, N0641_port_2,N0641_port_0,N0641_port_1, N0641_v);
  spice_node_1 n_S00724(eclk, ereset, S00724_port_1, S00724_v);
  spice_node_3 n_IOW(eclk, ereset, IOW_port_2,IOW_port_0,IOW_port_1, IOW_v);
  spice_node_3 n_IOR(eclk, ereset, IOR_port_3,IOR_port_1,IOR_port_5, IOR_v);
  spice_node_3 n_N0356(eclk, ereset, N0356_port_8,N0356_port_9,N0356_port_6, N0356_v);
  spice_node_2 n_N0643(eclk, ereset, N0643_port_2,N0643_port_1, N0643_v);
  spice_node_3 n_N0642(eclk, ereset, N0642_port_3,N0642_port_0,N0642_port_4, N0642_v);
  spice_node_1 n_S00833(eclk, ereset, S00833_port_0, S00833_v);
  spice_node_1 n_PC2_11(eclk, ereset, PC2_11_port_1, PC2_11_v);
  spice_node_1 n_PC2_10(eclk, ereset, PC2_10_port_0, PC2_10_v);
  spice_node_2 n_N0890(eclk, ereset, N0890_port_0,N0890_port_1, N0890_v);
  spice_node_2 n_N0644(eclk, ereset, N0644_port_0,N0644_port_1, N0644_v);
  spice_node_2 n_N0891(eclk, ereset, N0891_port_4,N0891_port_5, N0891_v);
  spice_node_5 n_JMS(eclk, ereset, JMS_port_2,JMS_port_3,JMS_port_1,JMS_port_4,JMS_port_5, JMS_v);
  spice_node_2 n_N0892(eclk, ereset, N0892_port_0,N0892_port_1, N0892_v);
  spice_node_3 n_CY_IB(eclk, ereset, CY_IB_port_2,CY_IB_port_0,CY_IB_port_1, CY_IB_v);
  spice_node_8 n_N0358(eclk, ereset, N0358_port_2,N0358_port_3,N0358_port_0,N0358_port_1,N0358_port_6,N0358_port_7,N0358_port_4,N0358_port_5, N0358_v);
  spice_node_5 n_SUB(eclk, ereset, SUB_port_2,SUB_port_3,SUB_port_0,SUB_port_1,SUB_port_4, SUB_v);
  spice_node_2 n_N0432(eclk, ereset, N0432_port_0,N0432_port_1, N0432_v);
  spice_node_1 n_N0433(eclk, ereset, N0433_port_0, N0433_v);
  spice_node_3 n_N0430(eclk, ereset, N0430_port_2,N0430_port_0,N0430_port_1, N0430_v);
  spice_node_1 n_N0431(eclk, ereset, N0431_port_0, N0431_v);
  spice_node_4 n_N0436(eclk, ereset, N0436_port_3,N0436_port_0,N0436_port_4,N0436_port_5, N0436_v);
  spice_node_2 n_N0437(eclk, ereset, N0437_port_2,N0437_port_0, N0437_v);
  spice_node_2 n_N0434(eclk, ereset, N0434_port_12,N0434_port_13, N0434_v);
  spice_node_2 n_N0435(eclk, ereset, N0435_port_2,N0435_port_1, N0435_v);
  spice_node_1 n_N0438(eclk, ereset, N0438_port_1, N0438_v);
  spice_node_2 n_N0439(eclk, ereset, N0439_port_12,N0439_port_13, N0439_v);
  spice_node_5 n_ADD(eclk, ereset, ADD_port_2,ADD_port_3,ADD_port_0,ADD_port_1,ADD_port_4, ADD_v);
  spice_node_6 n_ADM(eclk, ereset, ADM_port_2,ADM_port_3,ADM_port_0,ADM_port_1,ADM_port_4,ADM_port_5, ADM_v);
  spice_node_2 n_reset(eclk, ereset, reset_port_2,reset_port_0, reset_v);
  spice_node_3 n_N0728(eclk, ereset, N0728_port_2,N0728_port_0,N0728_port_1, N0728_v);
  spice_node_1 n_N0729(eclk, ereset, N0729_port_2, N0729_v);
  spice_node_3 n_N0726(eclk, ereset, N0726_port_2,N0726_port_0,N0726_port_1, N0726_v);
  spice_node_1 n_N0727(eclk, ereset, N0727_port_2, N0727_v);
  spice_node_3 n_N0724(eclk, ereset, N0724_port_2,N0724_port_0,N0724_port_1, N0724_v);
  spice_node_1 n_N0725(eclk, ereset, N0725_port_2, N0725_v);
  spice_node_3 n_N0722(eclk, ereset, N0722_port_2,N0722_port_0,N0722_port_1, N0722_v);
  spice_node_1 n_N0723(eclk, ereset, N0723_port_2, N0723_v);
  spice_node_3 n_N0720(eclk, ereset, N0720_port_2,N0720_port_0,N0720_port_1, N0720_v);
  spice_node_1 n_N0721(eclk, ereset, N0721_port_2, N0721_v);
  spice_node_2 n_N0946(eclk, ereset, N0946_port_2,N0946_port_1, N0946_v);
  spice_node_2 n_N0944(eclk, ereset, N0944_port_2,N0944_port_1, N0944_v);
  spice_node_2 n_N0942(eclk, ereset, N0942_port_2,N0942_port_1, N0942_v);
  spice_node_2 n_N0943(eclk, ereset, N0943_port_3,N0943_port_4, N0943_v);
  spice_node_2 n_N0940(eclk, ereset, N0940_port_2,N0940_port_1, N0940_v);
  spice_node_2 n_N0948(eclk, ereset, N0948_port_0,N0948_port_1, N0948_v);
  spice_node_2 n_N0949(eclk, ereset, N0949_port_0,N0949_port_1, N0949_v);
  spice_node_2 n_N0894(eclk, ereset, N0894_port_0,N0894_port_1, N0894_v);
  spice_node_2 n_N0895(eclk, ereset, N0895_port_0,N0895_port_1, N0895_v);
  spice_node_2 n_N0897(eclk, ereset, N0897_port_0,N0897_port_1, N0897_v);
  spice_node_2 n_N0893(eclk, ereset, N0893_port_4,N0893_port_5, N0893_v);
  spice_node_4 n_N0898(eclk, ereset, N0898_port_2,N0898_port_3,N0898_port_0,N0898_port_1, N0898_v);
  spice_node_4 n_N0899(eclk, ereset, N0899_port_2,N0899_port_3,N0899_port_0,N0899_port_1, N0899_v);
  spice_node_3 n_N0548(eclk, ereset, N0548_port_2,N0548_port_0,N0548_port_1, N0548_v);
  spice_node_3 n_N0549(eclk, ereset, N0549_port_2,N0549_port_0,N0549_port_1, N0549_v);
  spice_node_1 n_S00839(eclk, ereset, S00839_port_1, S00839_v);
  spice_node_2 n_N0542(eclk, ereset, N0542_port_4,N0542_port_5, N0542_v);
  spice_node_2 n_N0543(eclk, ereset, N0543_port_8,N0543_port_9, N0543_v);
  spice_node_2 n_N0540(eclk, ereset, N0540_port_1,N0540_port_5, N0540_v);
  spice_node_2 n_N0541(eclk, ereset, N0541_port_4,N0541_port_5, N0541_v);
  spice_node_3 n_N0546(eclk, ereset, N0546_port_2,N0546_port_0,N0546_port_1, N0546_v);
  spice_node_2 n_N0547(eclk, ereset, N0547_port_2,N0547_port_0, N0547_v);
  spice_node_2 n_N0544(eclk, ereset, N0544_port_8,N0544_port_9, N0544_v);
  spice_node_5 n_N0545(eclk, ereset, N0545_port_3,N0545_port_6,N0545_port_7,N0545_port_4,N0545_port_5, N0545_v);
  spice_node_5 n_N0467(eclk, ereset, N0467_port_2,N0467_port_3,N0467_port_1,N0467_port_4,N0467_port_5, N0467_v);
  spice_node_3 n_N0466(eclk, ereset, N0466_port_2,N0466_port_3,N0466_port_6, N0466_v);
  spice_node_4 n_INC_GROUP_5_(eclk, ereset, INC_GROUP_5__port_2,INC_GROUP_5__port_3,INC_GROUP_5__port_0,INC_GROUP_5__port_1, INC_GROUP_5__v);
  spice_node_2 n_N0502(eclk, ereset, N0502_port_2,N0502_port_0, N0502_v);
  spice_node_5 n_N0682(eclk, ereset, N0682_port_2,N0682_port_3,N0682_port_0,N0682_port_1,N0682_port_4, N0682_v);
  spice_node_2 n__OPR_3(eclk, ereset, _OPR_3_port_10,_OPR_3_port_11, _OPR_3_v);
  spice_node_2 n__OPR_2(eclk, ereset, _OPR_2_port_12,_OPR_2_port_13, _OPR_2_v);
  spice_node_2 n_N0966(eclk, ereset, N0966_port_0,N0966_port_1, N0966_v);
  spice_node_1 n_N0517(eclk, ereset, N0517_port_1, N0517_v);
  spice_node_2 n_N0516(eclk, ereset, N0516_port_0,N0516_port_1, N0516_v);
  spice_node_5 n_XCH(eclk, ereset, XCH_port_2,XCH_port_3,XCH_port_0,XCH_port_1,XCH_port_4, XCH_v);
  spice_node_6 n_CMC(eclk, ereset, CMC_port_2,CMC_port_3,CMC_port_0,CMC_port_1,CMC_port_4,CMC_port_5, CMC_v);
  spice_node_6 n_CMA(eclk, ereset, CMA_port_2,CMA_port_3,CMA_port_0,CMA_port_1,CMA_port_4,CMA_port_5, CMA_v);
  spice_node_2 n_N0510(eclk, ereset, N0510_port_0,N0510_port_1, N0510_v);
  spice_node_4 n_N0513(eclk, ereset, N0513_port_2,N0513_port_3,N0513_port_0,N0513_port_1, N0513_v);
  spice_node_3 n_M22(eclk, ereset, M22_port_8,M22_port_10,M22_port_11, M22_v);
  spice_node_4 n_JUN2_JMS2(eclk, ereset, JUN2_JMS2_port_2,JUN2_JMS2_port_3,JUN2_JMS2_port_0,JUN2_JMS2_port_1, JUN2_JMS2_v);
  spice_node_3 n_N0361(eclk, ereset, N0361_port_2,N0361_port_0,N0361_port_1, N0361_v);
  spice_node_2 n_N0512(eclk, ereset, N0512_port_0,N0512_port_1, N0512_v);
  spice_node_6 n_N0345(eclk, ereset, N0345_port_2,N0345_port_3,N0345_port_0,N0345_port_1,N0345_port_4,N0345_port_5, N0345_v);
  spice_node_2 n_SC_A22_M22_CLK2(eclk, ereset, SC_A22_M22_CLK2_port_8,SC_A22_M22_CLK2_port_9, SC_A22_M22_CLK2_v);
  spice_node_3 n_OPA_IB(eclk, ereset, OPA_IB_port_6,OPA_IB_port_4,OPA_IB_port_5, OPA_IB_v);
  spice_node_1 n_S00654(eclk, ereset, S00654_port_1, S00654_v);
  spice_node_1 n_S00818(eclk, ereset, S00818_port_0, S00818_v);
  spice_node_2 n_N0367(eclk, ereset, N0367_port_0,N0367_port_1, N0367_v);
  spice_node_3 n_N0364(eclk, ereset, N0364_port_3,N0364_port_0,N0364_port_1, N0364_v);
  spice_node_1 n_N0362(eclk, ereset, N0362_port_1, N0362_v);
  spice_node_6 n_N0363(eclk, ereset, N0363_port_2,N0363_port_3,N0363_port_0,N0363_port_1,N0363_port_4,N0363_port_5, N0363_v);
  spice_node_1 n_N0360(eclk, ereset, N0360_port_1, N0360_v);
  spice_node_1 n_S00729(eclk, ereset, S00729_port_1, S00729_v);
  spice_node_2 n_N0399(eclk, ereset, N0399_port_2,N0399_port_0, N0399_v);
  spice_node_7 n_N0396(eclk, ereset, N0396_port_2,N0396_port_3,N0396_port_0,N0396_port_1,N0396_port_6,N0396_port_4,N0396_port_5, N0396_v);
  spice_node_7 n_N0395(eclk, ereset, N0395_port_2,N0395_port_3,N0395_port_0,N0395_port_1,N0395_port_6,N0395_port_4,N0395_port_5, N0395_v);
  spice_node_7 n_N0394(eclk, ereset, N0394_port_2,N0394_port_3,N0394_port_0,N0394_port_1,N0394_port_6,N0394_port_4,N0394_port_5, N0394_v);
  spice_node_7 n_N0393(eclk, ereset, N0393_port_2,N0393_port_3,N0393_port_0,N0393_port_1,N0393_port_6,N0393_port_4,N0393_port_5, N0393_v);
  spice_node_7 n_N0392(eclk, ereset, N0392_port_2,N0392_port_3,N0392_port_0,N0392_port_1,N0392_port_6,N0392_port_4,N0392_port_5, N0392_v);
  spice_node_7 n_N0391(eclk, ereset, N0391_port_2,N0391_port_3,N0391_port_0,N0391_port_1,N0391_port_6,N0391_port_4,N0391_port_5, N0391_v);
  spice_node_7 n_N0390(eclk, ereset, N0390_port_2,N0390_port_3,N0390_port_0,N0390_port_1,N0390_port_6,N0390_port_4,N0390_port_5, N0390_v);
  spice_node_2 n_N0409(eclk, ereset, N0409_port_3,N0409_port_4, N0409_v);
  spice_node_1 n_N0408(eclk, ereset, N0408_port_0, N0408_v);
  spice_node_3 n_N0407(eclk, ereset, N0407_port_2,N0407_port_0,N0407_port_1, N0407_v);
  spice_node_2 n_N0406(eclk, ereset, N0406_port_12,N0406_port_13, N0406_v);
  spice_node_1 n_N0405(eclk, ereset, N0405_port_1, N0405_v);
  spice_node_3 n_N0404(eclk, ereset, N0404_port_2,N0404_port_0,N0404_port_1, N0404_v);
  spice_node_3 n_N0403(eclk, ereset, N0403_port_3,N0403_port_0,N0403_port_1, N0403_v);
  spice_node_3 n_N0402(eclk, ereset, N0402_port_2,N0402_port_0,N0402_port_1, N0402_v);
  spice_node_2 n_N0401(eclk, ereset, N0401_port_2,N0401_port_3, N0401_v);
  spice_node_2 n_N0400(eclk, ereset, N0400_port_0,N0400_port_1, N0400_v);
  spice_node_6 n_SBM(eclk, ereset, SBM_port_2,SBM_port_3,SBM_port_0,SBM_port_1,SBM_port_4,SBM_port_5, SBM_v);
  spice_node_2 n__CN(eclk, ereset, _CN_port_2,_CN_port_3, _CN_v);
  spice_node_1 n_S00678(eclk, ereset, S00678_port_1, S00678_v);
  spice_node_1 n_N0719(eclk, ereset, N0719_port_2, N0719_v);
  spice_node_3 n_N0718(eclk, ereset, N0718_port_2,N0718_port_0,N0718_port_1, N0718_v);
  spice_node_3 n_N0713(eclk, ereset, N0713_port_2,N0713_port_0,N0713_port_1, N0713_v);
  spice_node_3 n_N0712(eclk, ereset, N0712_port_2,N0712_port_0,N0712_port_1, N0712_v);
  spice_node_3 n_N0711(eclk, ereset, N0711_port_2,N0711_port_0,N0711_port_1, N0711_v);
  spice_node_2 n_N0710(eclk, ereset, N0710_port_2,N0710_port_1, N0710_v);
  spice_node_3 n_N0717(eclk, ereset, N0717_port_2,N0717_port_3,N0717_port_4, N0717_v);
  spice_node_3 n_N0715(eclk, ereset, N0715_port_0,N0715_port_1,N0715_port_4, N0715_v);
  spice_node_3 n_N0714(eclk, ereset, N0714_port_2,N0714_port_0,N0714_port_1, N0714_v);
  spice_node_2 n_N0973(eclk, ereset, N0973_port_0,N0973_port_1, N0973_v);
  spice_node_2 n_N0972(eclk, ereset, N0972_port_0,N0972_port_1, N0972_v);
  spice_node_2 n_N0971(eclk, ereset, N0971_port_0,N0971_port_1, N0971_v);
  spice_node_2 n_N0970(eclk, ereset, N0970_port_0,N0970_port_1, N0970_v);
  spice_node_2 n_N0977(eclk, ereset, N0977_port_0,N0977_port_1, N0977_v);
  spice_node_2 n_N0976(eclk, ereset, N0976_port_0,N0976_port_1, N0976_v);
  spice_node_2 n_N0975(eclk, ereset, N0975_port_0,N0975_port_1, N0975_v);
  spice_node_2 n_N0974(eclk, ereset, N0974_port_2,N0974_port_3, N0974_v);
  spice_node_2 n_N0979(eclk, ereset, N0979_port_0,N0979_port_1, N0979_v);
  spice_node_2 n_N0978(eclk, ereset, N0978_port_0,N0978_port_1, N0978_v);
  spice_node_2 n_SC_M12_CLK2(eclk, ereset, SC_M12_CLK2_port_0,SC_M12_CLK2_port_1, SC_M12_CLK2_v);
  spice_node_2 n_N0577(eclk, ereset, N0577_port_6,N0577_port_5, N0577_v);
  spice_node_2 n_N0576(eclk, ereset, N0576_port_0,N0576_port_1, N0576_v);
  spice_node_3 n_N0575(eclk, ereset, N0575_port_2,N0575_port_0,N0575_port_1, N0575_v);
  spice_node_3 n_N0574(eclk, ereset, N0574_port_3,N0574_port_0,N0574_port_4, N0574_v);
  spice_node_3 n_N0573(eclk, ereset, N0573_port_2,N0573_port_0,N0573_port_1, N0573_v);
  spice_node_2 n_N0572(eclk, ereset, N0572_port_0,N0572_port_1, N0572_v);
  spice_node_3 n_N0571(eclk, ereset, N0571_port_2,N0571_port_0,N0571_port_1, N0571_v);
  spice_node_5 n_N0570(eclk, ereset, N0570_port_3,N0570_port_6,N0570_port_7,N0570_port_4,N0570_port_5, N0570_v);
  spice_node_2 n_N0579(eclk, ereset, N0579_port_0,N0579_port_1, N0579_v);
  spice_node_2 n_N0578(eclk, ereset, N0578_port_2,N0578_port_1, N0578_v);
  spice_node_1 n_S00825(eclk, ereset, S00825_port_0, S00825_v);
  spice_node_1 n_S00531(eclk, ereset, S00531_port_0, S00531_v);
  spice_node_3 n_N0379(eclk, ereset, N0379_port_2,N0379_port_0,N0379_port_1, N0379_v);
  spice_node_1 n_S00536(eclk, ereset, S00536_port_1, S00536_v);
  spice_node_1 n_PC1_0(eclk, ereset, PC1_0_port_0, PC1_0_v);
  spice_node_1 n_R14_1(eclk, ereset, R14_1_port_1, R14_1_v);
  spice_node_1 n_R14_0(eclk, ereset, R14_0_port_0, R14_0_v);
  spice_node_1 n_R14_3(eclk, ereset, R14_3_port_1, R14_3_v);
  spice_node_1 n_R14_2(eclk, ereset, R14_2_port_0, R14_2_v);
  spice_node_1 n_R10_1(eclk, ereset, R10_1_port_1, R10_1_v);
  spice_node_1 n_R10_0(eclk, ereset, R10_0_port_0, R10_0_v);
  spice_node_1 n_R10_3(eclk, ereset, R10_3_port_1, R10_3_v);
  spice_node_1 n_R10_2(eclk, ereset, R10_2_port_0, R10_2_v);
  spice_node_2 n_N0889(eclk, ereset, N0889_port_4,N0889_port_5, N0889_v);
  spice_node_2 n_N0515(eclk, ereset, N0515_port_2,N0515_port_0, N0515_v);
  spice_node_6 n_N0514(eclk, ereset, N0514_port_2,N0514_port_3,N0514_port_0,N0514_port_6,N0514_port_4,N0514_port_5, N0514_v);
  spice_node_2 n_N0888(eclk, ereset, N0888_port_0,N0888_port_1, N0888_v);
  spice_node_2 n_N0845(eclk, ereset, N0845_port_0,N0845_port_1, N0845_v);
  spice_node_2 n_N0844(eclk, ereset, N0844_port_0,N0844_port_1, N0844_v);
  spice_node_4 n_N0511(eclk, ereset, N0511_port_2,N0511_port_3,N0511_port_0,N0511_port_1, N0511_v);
  spice_node_2 n_N0842(eclk, ereset, N0842_port_0,N0842_port_1, N0842_v);
  spice_node_3 n_N0371(eclk, ereset, N0371_port_2,N0371_port_3,N0371_port_0, N0371_v);
  spice_node_1 n_N0849(eclk, ereset, N0849_port_1, N0849_v);
  spice_node_6 n_N0848(eclk, ereset, N0848_port_2,N0848_port_0,N0848_port_1,N0848_port_6,N0848_port_4,N0848_port_5, N0848_v);
  spice_node_5 n_ISZ(eclk, ereset, ISZ_port_2,ISZ_port_3,ISZ_port_0,ISZ_port_1,ISZ_port_4, ISZ_v);
  spice_node_6 n_N0370(eclk, ereset, N0370_port_2,N0370_port_3,N0370_port_0,N0370_port_1,N0370_port_4,N0370_port_5, N0370_v);
  spice_node_3 n_N0875(eclk, ereset, N0875_port_3,N0875_port_1,N0875_port_4, N0875_v);
  spice_node_1 n_R12_3(eclk, ereset, R12_3_port_1, R12_3_v);
  spice_node_6 n_CLB(eclk, ereset, CLB_port_2,CLB_port_3,CLB_port_0,CLB_port_1,CLB_port_4,CLB_port_5, CLB_v);
  spice_node_6 n_CLC(eclk, ereset, CLC_port_2,CLC_port_3,CLC_port_0,CLC_port_1,CLC_port_4,CLC_port_5, CLC_v);
  spice_node_4 n_M12(eclk, ereset, M12_port_10,M12_port_11,M12_port_8,M12_port_7, M12_v);
  spice_node_2 n___X21__CLK2_(eclk, ereset, __X21__CLK2__port_2,__X21__CLK2__port_3, __X21__CLK2__v);
  spice_node_2 n_DC(eclk, ereset, DC_port_4,DC_port_5, DC_v);
  spice_node_7 n_N0388(eclk, ereset, N0388_port_2,N0388_port_3,N0388_port_0,N0388_port_1,N0388_port_6,N0388_port_4,N0388_port_5, N0388_v);
  spice_node_7 n_N0389(eclk, ereset, N0389_port_2,N0389_port_3,N0389_port_0,N0389_port_1,N0389_port_6,N0389_port_4,N0389_port_5, N0389_v);
  spice_node_1 n_N0380(eclk, ereset, N0380_port_0, N0380_v);
  spice_node_2 n_N0381(eclk, ereset, N0381_port_12,N0381_port_13, N0381_v);
  spice_node_3 n_N0382(eclk, ereset, N0382_port_3,N0382_port_4,N0382_port_5, N0382_v);
  spice_node_1 n_N0384(eclk, ereset, N0384_port_1, N0384_v);
  spice_node_7 n_N0385(eclk, ereset, N0385_port_2,N0385_port_3,N0385_port_0,N0385_port_1,N0385_port_6,N0385_port_4,N0385_port_5, N0385_v);
  spice_node_7 n_N0386(eclk, ereset, N0386_port_2,N0386_port_3,N0386_port_0,N0386_port_1,N0386_port_6,N0386_port_4,N0386_port_5, N0386_v);
  spice_node_7 n_N0387(eclk, ereset, N0387_port_2,N0387_port_3,N0387_port_0,N0387_port_1,N0387_port_6,N0387_port_4,N0387_port_5, N0387_v);
  spice_node_1 n_R12_0(eclk, ereset, R12_0_port_0, R12_0_v);
  spice_node_3 n_N0419(eclk, ereset, N0419_port_2,N0419_port_3,N0419_port_1, N0419_v);
  spice_node_2 n_N0410(eclk, ereset, N0410_port_12,N0410_port_13, N0410_v);
  spice_node_3 n_N0411(eclk, ereset, N0411_port_3,N0411_port_4,N0411_port_5, N0411_v);
  spice_node_2 n_N0412(eclk, ereset, N0412_port_0,N0412_port_1, N0412_v);
  spice_node_4 n_N0413(eclk, ereset, N0413_port_2,N0413_port_3,N0413_port_0,N0413_port_1, N0413_v);
  spice_node_1 n_N0414(eclk, ereset, N0414_port_0, N0414_v);
  spice_node_3 n_N0415(eclk, ereset, N0415_port_2,N0415_port_0,N0415_port_1, N0415_v);
  spice_node_1 n_N0416(eclk, ereset, N0416_port_1, N0416_v);
  spice_node_2 n_N0417(eclk, ereset, N0417_port_0,N0417_port_1, N0417_v);
  spice_node_2 n__COM(eclk, ereset, _COM_port_0,_COM_port_1, _COM_v);
  spice_node_4 n_N0901(eclk, ereset, N0901_port_2,N0901_port_3,N0901_port_0,N0901_port_1, N0901_v);
  spice_node_2 n_N0704(eclk, ereset, N0704_port_0,N0704_port_1, N0704_v);
  spice_node_4 n_N0705(eclk, ereset, N0705_port_2,N0705_port_3,N0705_port_0,N0705_port_1, N0705_v);
  spice_node_2 n_N0706(eclk, ereset, N0706_port_0,N0706_port_1, N0706_v);
  spice_node_1 n_N0707(eclk, ereset, N0707_port_0, N0707_v);
  spice_node_2 n_N0700(eclk, ereset, N0700_port_2,N0700_port_3, N0700_v);
  spice_node_4 n_N0701(eclk, ereset, N0701_port_2,N0701_port_3,N0701_port_0,N0701_port_1, N0701_v);
  spice_node_2 n_N0702(eclk, ereset, N0702_port_0,N0702_port_1, N0702_v);
  spice_node_1 n_N0703(eclk, ereset, N0703_port_0, N0703_v);
  spice_node_4 n_N0708(eclk, ereset, N0708_port_2,N0708_port_3,N0708_port_4,N0708_port_5, N0708_v);
  spice_node_2 n_N0709(eclk, ereset, N0709_port_0,N0709_port_1, N0709_v);
  spice_node_2 n_N0885(eclk, ereset, N0885_port_2,N0885_port_1, N0885_v);
  spice_node_3 n_N0378(eclk, ereset, N0378_port_2,N0378_port_0,N0378_port_1, N0378_v);
  spice_node_18 n_D2(eclk, ereset, D2_port_8,D2_port_9,D2_port_2,D2_port_3,D2_port_0,D2_port_1,D2_port_6,D2_port_7,D2_port_4,D2_port_5,D2_port_10,D2_port_11,D2_port_13,D2_port_14,D2_port_15,D2_port_16,D2_port_17,D2_port_18, D2_v);
  spice_node_18 n_D3(eclk, ereset, D3_port_8,D3_port_9,D3_port_2,D3_port_3,D3_port_0,D3_port_1,D3_port_6,D3_port_7,D3_port_4,D3_port_5,D3_port_11,D3_port_12,D3_port_13,D3_port_14,D3_port_15,D3_port_16,D3_port_17,D3_port_18, D3_v);
  spice_node_18 n_D0(eclk, ereset, D0_port_8,D0_port_9,D0_port_2,D0_port_3,D0_port_0,D0_port_1,D0_port_6,D0_port_7,D0_port_4,D0_port_5,D0_port_10,D0_port_11,D0_port_12,D0_port_13,D0_port_14,D0_port_15,D0_port_16,D0_port_17, D0_v);
  spice_node_18 n_D1(eclk, ereset, D1_port_8,D1_port_9,D1_port_2,D1_port_3,D1_port_0,D1_port_1,D1_port_6,D1_port_7,D1_port_4,D1_port_5,D1_port_10,D1_port_11,D1_port_12,D1_port_13,D1_port_14,D1_port_15,D1_port_16,D1_port_17, D1_v);
  spice_node_2 n_N0968(eclk, ereset, N0968_port_0,N0968_port_1, N0968_v);
  spice_node_2 n_N0969(eclk, ereset, N0969_port_0,N0969_port_1, N0969_v);
  spice_node_2 n_N0965(eclk, ereset, N0965_port_2,N0965_port_3, N0965_v);
  spice_node_2 n_N0967(eclk, ereset, N0967_port_0,N0967_port_1, N0967_v);
  spice_node_2 n_N0960(eclk, ereset, N0960_port_0,N0960_port_1, N0960_v);
  spice_node_2 n_N0961(eclk, ereset, N0961_port_0,N0961_port_1, N0961_v);
  spice_node_2 n_N0962(eclk, ereset, N0962_port_0,N0962_port_1, N0962_v);
  spice_node_2 n_N0963(eclk, ereset, N0963_port_0,N0963_port_1, N0963_v);
  spice_node_2 n_N0907(eclk, ereset, N0907_port_0,N0907_port_1, N0907_v);
  spice_node_2 n_N0884(eclk, ereset, N0884_port_2,N0884_port_1, N0884_v);
  spice_node_2 n_N0560(eclk, ereset, N0560_port_6,N0560_port_5, N0560_v);
  spice_node_2 n_N0561(eclk, ereset, N0561_port_0,N0561_port_1, N0561_v);
  spice_node_3 n_N0562(eclk, ereset, N0562_port_2,N0562_port_0,N0562_port_1, N0562_v);
  spice_node_2 n_N0563(eclk, ereset, N0563_port_0,N0563_port_1, N0563_v);
  spice_node_2 n_N0564(eclk, ereset, N0564_port_3,N0564_port_0, N0564_v);
  spice_node_2 n_N0565(eclk, ereset, N0565_port_8,N0565_port_9, N0565_v);
  spice_node_1 n_N0566(eclk, ereset, N0566_port_0, N0566_v);
  spice_node_2 n_N0567(eclk, ereset, N0567_port_0,N0567_port_1, N0567_v);
  spice_node_2 n_N0568(eclk, ereset, N0568_port_0,N0568_port_1, N0568_v);
  spice_node_2 n_N0569(eclk, ereset, N0569_port_8,N0569_port_9, N0569_v);
  spice_node_3 n_N0365(eclk, ereset, N0365_port_2,N0365_port_0,N0365_port_1, N0365_v);
  spice_node_1 n_S00814(eclk, ereset, S00814_port_0, S00814_v);
  spice_node_4 n_N0368(eclk, ereset, N0368_port_2,N0368_port_3,N0368_port_0,N0368_port_1, N0368_v);
  spice_node_3 n_N0369(eclk, ereset, N0369_port_2,N0369_port_0,N0369_port_1, N0369_v);
  spice_node_1 n_S00676(eclk, ereset, S00676_port_0, S00676_v);
  spice_node_2 n_N0640(eclk, ereset, N0640_port_0,N0640_port_1, N0640_v);
  spice_node_3 n_N0314(eclk, ereset, N0314_port_2,N0314_port_0,N0314_port_1, N0314_v);
  spice_node_2 n__OPA_0(eclk, ereset, _OPA_0_port_13,_OPA_0_port_14, _OPA_0_v);
  spice_node_2 n_N0311(eclk, ereset, N0311_port_0,N0311_port_1, N0311_v);
  spice_node_2 n__OPA_2(eclk, ereset, _OPA_2_port_6,_OPA_2_port_7, _OPA_2_v);
  spice_node_2 n__OPA_3(eclk, ereset, _OPA_3_port_10,_OPA_3_port_11, _OPA_3_v);
  spice_node_2 n_N0646(eclk, ereset, N0646_port_2,N0646_port_1, N0646_v);
  spice_node_5 n_ADD_GROUP_4_(eclk, ereset, ADD_GROUP_4__port_2,ADD_GROUP_4__port_3,ADD_GROUP_4__port_0,ADD_GROUP_4__port_1,ADD_GROUP_4__port_4, ADD_GROUP_4__v);
  spice_node_6 n____SC__JIN_FIN__CLK1_M11_X21_INH_(eclk, ereset, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_2,___SC__JIN_FIN__CLK1_M11_X21_INH__port_3,___SC__JIN_FIN__CLK1_M11_X21_INH__port_0,___SC__JIN_FIN__CLK1_M11_X21_INH__port_1,___SC__JIN_FIN__CLK1_M11_X21_INH__port_4,___SC__JIN_FIN__CLK1_M11_X21_INH__port_5, ___SC__JIN_FIN__CLK1_M11_X21_INH__v);
  spice_node_4 n_N0486(eclk, ereset, N0486_port_2,N0486_port_3,N0486_port_4,N0486_port_5, N0486_v);
  spice_node_2 n_N0860(eclk, ereset, N0860_port_0,N0860_port_1, N0860_v);
  spice_node_2 n_N0947(eclk, ereset, N0947_port_0,N0947_port_1, N0947_v);
  spice_node_2 n_N0941(eclk, ereset, N0941_port_3,N0941_port_4, N0941_v);
  spice_node_3 n_N0861(eclk, ereset, N0861_port_2,N0861_port_3,N0861_port_0, N0861_v);
  spice_node_4 n_N0863(eclk, ereset, N0863_port_2,N0863_port_3,N0863_port_0,N0863_port_1, N0863_v);
  spice_node_4 n_N0862(eclk, ereset, N0862_port_2,N0862_port_3,N0862_port_0,N0862_port_1, N0862_v);
  spice_node_4 n_N0865(eclk, ereset, N0865_port_2,N0865_port_3,N0865_port_0,N0865_port_1, N0865_v);
  spice_node_4 n_N0864(eclk, ereset, N0864_port_2,N0864_port_3,N0864_port_0,N0864_port_1, N0864_v);
  spice_node_16 n_WRITE_ACC_1_(eclk, ereset, WRITE_ACC_1__port_8,WRITE_ACC_1__port_9,WRITE_ACC_1__port_2,WRITE_ACC_1__port_3,WRITE_ACC_1__port_0,WRITE_ACC_1__port_1,WRITE_ACC_1__port_6,WRITE_ACC_1__port_7,WRITE_ACC_1__port_4,WRITE_ACC_1__port_5,WRITE_ACC_1__port_10,WRITE_ACC_1__port_11,WRITE_ACC_1__port_12,WRITE_ACC_1__port_13,WRITE_ACC_1__port_14,WRITE_ACC_1__port_15, WRITE_ACC_1__v);
  spice_node_10 n_N0866(eclk, ereset, N0866_port_8,N0866_port_9,N0866_port_2,N0866_port_3,N0866_port_0,N0866_port_6,N0866_port_7,N0866_port_4,N0866_port_5,N0866_port_10, N0866_v);
  spice_node_4 n_N0855(eclk, ereset, N0855_port_2,N0855_port_3,N0855_port_1,N0855_port_4, N0855_v);
  spice_node_2 n_N0896(eclk, ereset, N0896_port_0,N0896_port_1, N0896_v);
  spice_node_5 n_IO(eclk, ereset, IO_port_2,IO_port_3,IO_port_0,IO_port_1,IO_port_4, IO_v);
  spice_node_3 n_N0911(eclk, ereset, N0911_port_2,N0911_port_0,N0911_port_1, N0911_v);
  spice_node_2 n_N0621(eclk, ereset, N0621_port_0,N0621_port_1, N0621_v);
  spice_node_2 n_N0910(eclk, ereset, N0910_port_0,N0910_port_1, N0910_v);
  spice_node_1 n_N0280(eclk, ereset, N0280_port_0, N0280_v);
  spice_node_1 n_N0284(eclk, ereset, N0284_port_1, N0284_v);
  spice_node_1 n_N0286(eclk, ereset, N0286_port_1, N0286_v);
  spice_node_1 n_N0289(eclk, ereset, N0289_port_3, N0289_v);
  spice_node_9 n_N0288(eclk, ereset, N0288_port_8,N0288_port_2,N0288_port_3,N0288_port_0,N0288_port_1,N0288_port_6,N0288_port_7,N0288_port_4,N0288_port_5, N0288_v);
  spice_node_6 n_N0771(eclk, ereset, N0771_port_2,N0771_port_3,N0771_port_1,N0771_port_6,N0771_port_4,N0771_port_5, N0771_v);
  spice_node_6 n_N0770(eclk, ereset, N0770_port_2,N0770_port_3,N0770_port_1,N0770_port_6,N0770_port_4,N0770_port_5, N0770_v);
  spice_node_6 n_N0773(eclk, ereset, N0773_port_2,N0773_port_3,N0773_port_1,N0773_port_6,N0773_port_4,N0773_port_5, N0773_v);
  spice_node_6 n_N0772(eclk, ereset, N0772_port_2,N0772_port_3,N0772_port_1,N0772_port_6,N0772_port_4,N0772_port_5, N0772_v);
  spice_node_6 n_N0775(eclk, ereset, N0775_port_2,N0775_port_3,N0775_port_0,N0775_port_6,N0775_port_4,N0775_port_5, N0775_v);
  spice_node_6 n_N0774(eclk, ereset, N0774_port_2,N0774_port_3,N0774_port_0,N0774_port_6,N0774_port_4,N0774_port_5, N0774_v);
  spice_node_6 n_N0777(eclk, ereset, N0777_port_2,N0777_port_3,N0777_port_1,N0777_port_6,N0777_port_4,N0777_port_5, N0777_v);
  spice_node_6 n_N0776(eclk, ereset, N0776_port_2,N0776_port_3,N0776_port_0,N0776_port_6,N0776_port_4,N0776_port_5, N0776_v);
  spice_node_6 n_N0779(eclk, ereset, N0779_port_2,N0779_port_3,N0779_port_0,N0779_port_6,N0779_port_4,N0779_port_5, N0779_v);
  spice_node_6 n_N0778(eclk, ereset, N0778_port_2,N0778_port_3,N0778_port_0,N0778_port_6,N0778_port_4,N0778_port_5, N0778_v);
  spice_node_2 n_N0919(eclk, ereset, N0919_port_2,N0919_port_3, N0919_v);
  spice_node_2 n_N0918(eclk, ereset, N0918_port_0,N0918_port_1, N0918_v);
  spice_node_3 n_N0626(eclk, ereset, N0626_port_3,N0626_port_1,N0626_port_4, N0626_v);
  spice_node_3 n_N0914(eclk, ereset, N0914_port_2,N0914_port_0,N0914_port_1, N0914_v);
  spice_node_2 n_test(eclk, ereset, test_port_2,test_port_0, test_v);
  spice_node_1 n_S00834(eclk, ereset, S00834_port_0, S00834_v);
  spice_node_2 n_N0915(eclk, ereset, N0915_port_0,N0915_port_1, N0915_v);
  spice_node_1 n_S00804(eclk, ereset, S00804_port_0, S00804_v);
  spice_node_5 n_N0599(eclk, ereset, N0599_port_3,N0599_port_6,N0599_port_7,N0599_port_4,N0599_port_5, N0599_v);
  spice_node_2 n_N0598(eclk, ereset, N0598_port_8,N0598_port_9, N0598_v);
  spice_node_1 n_S00801(eclk, ereset, S00801_port_1, S00801_v);
  spice_node_1 n_S00800(eclk, ereset, S00800_port_0, S00800_v);
  spice_node_2 n_N0595(eclk, ereset, N0595_port_0,N0595_port_1, N0595_v);
  spice_node_2 n_N0594(eclk, ereset, N0594_port_0,N0594_port_1, N0594_v);
  spice_node_2 n_N0597(eclk, ereset, N0597_port_0,N0597_port_1, N0597_v);
  spice_node_2 n_N0596(eclk, ereset, N0596_port_0,N0596_port_1, N0596_v);
  spice_node_2 n_N0591(eclk, ereset, N0591_port_8,N0591_port_9, N0591_v);
  spice_node_2 n_N0590(eclk, ereset, N0590_port_2,N0590_port_1, N0590_v);
  spice_node_1 n_N0593(eclk, ereset, N0593_port_0, N0593_v);
  spice_node_1 n_N0592(eclk, ereset, N0592_port_1, N0592_v);
  spice_node_3 n_N0609(eclk, ereset, N0609_port_2,N0609_port_0,N0609_port_1, N0609_v);
  spice_node_6 n_N0359(eclk, ereset, N0359_port_2,N0359_port_3,N0359_port_0,N0359_port_1,N0359_port_4,N0359_port_5, N0359_v);
  spice_node_2 n_N0606(eclk, ereset, N0606_port_0,N0606_port_1, N0606_v);
  spice_node_2 n_N0601(eclk, ereset, N0601_port_0,N0601_port_1, N0601_v);
  spice_node_3 n_N0600(eclk, ereset, N0600_port_2,N0600_port_3,N0600_port_0, N0600_v);
  spice_node_2 n_N0603(eclk, ereset, N0603_port_2,N0603_port_1, N0603_v);
  spice_node_3 n_N0602(eclk, ereset, N0602_port_2,N0602_port_0,N0602_port_1, N0602_v);
  spice_node_2 n_N0825(eclk, ereset, N0825_port_0,N0825_port_1, N0825_v);
  spice_node_2 n_N0827(eclk, ereset, N0827_port_0,N0827_port_1, N0827_v);
  spice_node_2 n_N0826(eclk, ereset, N0826_port_0,N0826_port_1, N0826_v);
  spice_node_2 n_N0821(eclk, ereset, N0821_port_0,N0821_port_1, N0821_v);
  spice_node_2 n_N0917(eclk, ereset, N0917_port_0,N0917_port_1, N0917_v);
  spice_node_4 n___INH__X11_X31_CLK1(eclk, ereset, __INH__X11_X31_CLK1_port_12,__INH__X11_X31_CLK1_port_13,__INH__X11_X31_CLK1_port_14,__INH__X11_X31_CLK1_port_15, __INH__X11_X31_CLK1_v);
  spice_node_1 n_S00761(eclk, ereset, S00761_port_0, S00761_v);
  spice_node_2 n_N0817(eclk, ereset, N0817_port_0,N0817_port_1, N0817_v);
  spice_node_2 n_N0811(eclk, ereset, N0811_port_0,N0811_port_1, N0811_v);
  spice_node_1 n_S00781(eclk, ereset, S00781_port_1, S00781_v);
  spice_node_3 n_CY_ADAC(eclk, ereset, CY_ADAC_port_2,CY_ADAC_port_0,CY_ADAC_port_1, CY_ADAC_v);
  spice_node_2 n_N0652(eclk, ereset, N0652_port_0,N0652_port_1, N0652_v);
  spice_node_10 n_CLK2_SC_A12_M12_(eclk, ereset, CLK2_SC_A12_M12__port_8,CLK2_SC_A12_M12__port_9,CLK2_SC_A12_M12__port_2,CLK2_SC_A12_M12__port_3,CLK2_SC_A12_M12__port_0,CLK2_SC_A12_M12__port_1,CLK2_SC_A12_M12__port_6,CLK2_SC_A12_M12__port_7,CLK2_SC_A12_M12__port_4,CLK2_SC_A12_M12__port_5, CLK2_SC_A12_M12__v);
  spice_node_1 n_N0292(eclk, ereset, N0292_port_4, N0292_v);
  spice_node_2 n_N0293(eclk, ereset, N0293_port_2,N0293_port_3, N0293_v);
  spice_node_1 n_N0290(eclk, ereset, N0290_port_0, N0290_v);
  spice_node_1 n_N0291(eclk, ereset, N0291_port_5, N0291_v);
  spice_node_4 n_N0296(eclk, ereset, N0296_port_2,N0296_port_3,N0296_port_0,N0296_port_1, N0296_v);
  spice_node_2 n_N0297(eclk, ereset, N0297_port_0,N0297_port_1, N0297_v);
  spice_node_4 n_N0294(eclk, ereset, N0294_port_2,N0294_port_3,N0294_port_0,N0294_port_1, N0294_v);
  spice_node_1 n_N0295(eclk, ereset, N0295_port_1, N0295_v);
  spice_node_2 n_N0298(eclk, ereset, N0298_port_3,N0298_port_0, N0298_v);
  spice_node_2 n_N0299(eclk, ereset, N0299_port_0,N0299_port_1, N0299_v);
  spice_node_6 n_N0762(eclk, ereset, N0762_port_2,N0762_port_3,N0762_port_0,N0762_port_1,N0762_port_4,N0762_port_5, N0762_v);
  spice_node_6 n_N0763(eclk, ereset, N0763_port_2,N0763_port_3,N0763_port_0,N0763_port_1,N0763_port_4,N0763_port_5, N0763_v);
  spice_node_3 n_N0760(eclk, ereset, N0760_port_2,N0760_port_0,N0760_port_1, N0760_v);
  spice_node_6 n_N0761(eclk, ereset, N0761_port_2,N0761_port_3,N0761_port_0,N0761_port_1,N0761_port_4,N0761_port_5, N0761_v);
  spice_node_2 n_N0766(eclk, ereset, N0766_port_0,N0766_port_1, N0766_v);
  spice_node_2 n_N0767(eclk, ereset, N0767_port_2,N0767_port_0, N0767_v);
  spice_node_6 n_N0764(eclk, ereset, N0764_port_2,N0764_port_3,N0764_port_0,N0764_port_1,N0764_port_4,N0764_port_5, N0764_v);
  spice_node_2 n_N0765(eclk, ereset, N0765_port_2,N0765_port_1, N0765_v);
  spice_node_2 n_N0768(eclk, ereset, N0768_port_2,N0768_port_0, N0768_v);
  spice_node_3 n_N0769(eclk, ereset, N0769_port_2,N0769_port_0,N0769_port_1, N0769_v);
  spice_node_2 n_N0908(eclk, ereset, N0908_port_0,N0908_port_1, N0908_v);
  spice_node_2 n_N0909(eclk, ereset, N0909_port_0,N0909_port_1, N0909_v);
  spice_node_2 n_N0903(eclk, ereset, N0903_port_0,N0903_port_1, N0903_v);
  spice_node_2 n_sync(eclk, ereset, sync_port_0,sync_port_1, sync_v);
  spice_node_2 n_N0904(eclk, ereset, N0904_port_0,N0904_port_1, N0904_v);
  spice_node_2 n_N0905(eclk, ereset, N0905_port_0,N0905_port_1, N0905_v);
  spice_node_2 n_SC_A12_CLK2(eclk, ereset, SC_A12_CLK2_port_2,SC_A12_CLK2_port_3, SC_A12_CLK2_v);
  spice_node_1 n_R3_2(eclk, ereset, R3_2_port_1, R3_2_v);
  spice_node_4 n_N0588(eclk, ereset, N0588_port_2,N0588_port_3,N0588_port_0,N0588_port_1, N0588_v);
  spice_node_2 n_N0589(eclk, ereset, N0589_port_0,N0589_port_1, N0589_v);
  spice_node_1 n_N0586(eclk, ereset, N0586_port_0, N0586_v);
  spice_node_7 n_N0587(eclk, ereset, N0587_port_2,N0587_port_3,N0587_port_0,N0587_port_1,N0587_port_6,N0587_port_4,N0587_port_5, N0587_v);
  spice_node_5 n_N0584(eclk, ereset, N0584_port_3,N0584_port_6,N0584_port_7,N0584_port_4,N0584_port_5, N0584_v);
  spice_node_2 n_N0582(eclk, ereset, N0582_port_2,N0582_port_1, N0582_v);
  spice_node_2 n_N0583(eclk, ereset, N0583_port_8,N0583_port_9, N0583_v);
  spice_node_2 n_N0580(eclk, ereset, N0580_port_2,N0580_port_1, N0580_v);
  spice_node_2 n_N0581(eclk, ereset, N0581_port_8,N0581_port_9, N0581_v);
  spice_node_3 n_N0618(eclk, ereset, N0618_port_2,N0618_port_0,N0618_port_1, N0618_v);
  spice_node_2 n_N0619(eclk, ereset, N0619_port_8,N0619_port_9, N0619_v);
  spice_node_2 n_N0616(eclk, ereset, N0616_port_8,N0616_port_9, N0616_v);
  spice_node_2 n_N0614(eclk, ereset, N0614_port_0,N0614_port_1, N0614_v);
  spice_node_2 n_N0613(eclk, ereset, N0613_port_0,N0613_port_6, N0613_v);
  spice_node_2 n_N0836(eclk, ereset, N0836_port_0,N0836_port_1, N0836_v);
  spice_node_2 n_N0837(eclk, ereset, N0837_port_0,N0837_port_1, N0837_v);
  spice_node_2 n_N0835(eclk, ereset, N0835_port_0,N0835_port_1, N0835_v);
  spice_node_2 n_N0832(eclk, ereset, N0832_port_0,N0832_port_1, N0832_v);
  spice_node_2 n_N0833(eclk, ereset, N0833_port_2,N0833_port_3, N0833_v);
  spice_node_2 n_N0830(eclk, ereset, N0830_port_0,N0830_port_1, N0830_v);
  spice_node_2 n_N0831(eclk, ereset, N0831_port_0,N0831_port_1, N0831_v);
  spice_node_1 n_S00612(eclk, ereset, S00612_port_1, S00612_v);
  spice_node_1 n_S00613(eclk, ereset, S00613_port_0, S00613_v);
  spice_node_2 n_N0838(eclk, ereset, N0838_port_0,N0838_port_1, N0838_v);
  spice_node_2 n_N0839(eclk, ereset, N0839_port_0,N0839_port_1, N0839_v);
  spice_node_1 n_S00580(eclk, ereset, S00580_port_1, S00580_v);
  spice_node_1 n_S00581(eclk, ereset, S00581_port_1, S00581_v);
  spice_node_1 n_S00584(eclk, ereset, S00584_port_1, S00584_v);
  spice_node_1 n_S00585(eclk, ereset, S00585_port_1, S00585_v);
  spice_node_2 n_cm_ram2(eclk, ereset, cm_ram2_port_0,cm_ram2_port_1, cm_ram2_v);
  spice_node_1 n_S00725(eclk, ereset, S00725_port_0, S00725_v);
  spice_node_1 n_R2_1(eclk, ereset, R2_1_port_1, R2_1_v);
  spice_node_1 n_R2_0(eclk, ereset, R2_0_port_0, R2_0_v);
  spice_node_1 n_R2_3(eclk, ereset, R2_3_port_1, R2_3_v);
  spice_node_1 n_R2_2(eclk, ereset, R2_2_port_0, R2_2_v);
  spice_node_1 n_R0_3(eclk, ereset, R0_3_port_1, R0_3_v);
  spice_node_1 n_R0_2(eclk, ereset, R0_2_port_0, R0_2_v);
  spice_node_1 n_R0_1(eclk, ereset, R0_1_port_1, R0_1_v);
  spice_node_1 n_R0_0(eclk, ereset, R0_0_port_0, R0_0_v);
  spice_node_2 n_SC(eclk, ereset, SC_port_4,SC_port_13, SC_v);
  spice_node_1 n_R1_0(eclk, ereset, R1_0_port_1, R1_0_v);
  spice_node_1 n_R1_1(eclk, ereset, R1_1_port_0, R1_1_v);
  spice_node_1 n_R6_1(eclk, ereset, R6_1_port_1, R6_1_v);
  spice_node_1 n_R6_0(eclk, ereset, R6_0_port_0, R6_0_v);
  spice_node_1 n_R6_3(eclk, ereset, R6_3_port_1, R6_3_v);
  spice_node_1 n_R6_2(eclk, ereset, R6_2_port_0, R6_2_v);
  spice_node_3 n_N0629(eclk, ereset, N0629_port_2,N0629_port_0,N0629_port_1, N0629_v);
  spice_node_5 n_N0628(eclk, ereset, N0628_port_2,N0628_port_3,N0628_port_0,N0628_port_1,N0628_port_4, N0628_v);
  spice_node_1 n_N0851(eclk, ereset, N0851_port_1, N0851_v);
  spice_node_1 n_R4_3(eclk, ereset, R4_3_port_1, R4_3_v);
  spice_node_1 n_R4_2(eclk, ereset, R4_2_port_0, R4_2_v);
  spice_node_1 n_R4_1(eclk, ereset, R4_1_port_1, R4_1_v);
  spice_node_1 n_R4_0(eclk, ereset, R4_0_port_0, R4_0_v);
  spice_node_2 n_N0623(eclk, ereset, N0623_port_0,N0623_port_1, N0623_v);
  spice_node_2 n_N0622(eclk, ereset, N0622_port_2,N0622_port_3, N0622_v);
  spice_node_2 n_N0333(eclk, ereset, N0333_port_0,N0333_port_1, N0333_v);
  spice_node_5 n_N0620(eclk, ereset, N0620_port_3,N0620_port_6,N0620_port_7,N0620_port_4,N0620_port_5, N0620_v);
  spice_node_2 n_N0627(eclk, ereset, N0627_port_2,N0627_port_0, N0627_v);
  spice_node_2 n_N0334(eclk, ereset, N0334_port_0,N0334_port_1, N0334_v);
  spice_node_1 n_N0625(eclk, ereset, N0625_port_0, N0625_v);
  spice_node_2 n_N0624(eclk, ereset, N0624_port_0,N0624_port_1, N0624_v);
  spice_node_3 n_N0803(eclk, ereset, N0803_port_3,N0803_port_1,N0803_port_4, N0803_v);
  spice_node_2 n_N0854(eclk, ereset, N0854_port_0,N0854_port_6, N0854_v);
  spice_node_3 n_ADSR(eclk, ereset, ADSR_port_2,ADSR_port_0,ADSR_port_1, ADSR_v);
  spice_node_4 n_ADDR_PTR_1(eclk, ereset, ADDR_PTR_1_port_2,ADDR_PTR_1_port_3,ADDR_PTR_1_port_0,ADDR_PTR_1_port_1, ADDR_PTR_1_v);
  spice_node_4 n_ADDR_PTR_0(eclk, ereset, ADDR_PTR_0_port_2,ADDR_PTR_0_port_3,ADDR_PTR_0_port_0,ADDR_PTR_0_port_1, ADDR_PTR_0_v);
  spice_node_10 n_READ_ACC_3_(eclk, ereset, READ_ACC_3__port_8,READ_ACC_3__port_9,READ_ACC_3__port_2,READ_ACC_3__port_3,READ_ACC_3__port_0,READ_ACC_3__port_1,READ_ACC_3__port_6,READ_ACC_3__port_7,READ_ACC_3__port_4,READ_ACC_3__port_5, READ_ACC_3__v);
  spice_node_4 n_L(eclk, ereset, L_port_2,L_port_0,L_port_1,L_port_5, L_v);
  spice_node_4 n_N0856(eclk, ereset, N0856_port_2,N0856_port_3,N0856_port_0,N0856_port_1, N0856_v);
  spice_node_4 n_N0857(eclk, ereset, N0857_port_2,N0857_port_3,N0857_port_1,N0857_port_4, N0857_v);
  spice_node_2 n__OPE(eclk, ereset, _OPE_port_0,_OPE_port_1, _OPE_v);
  spice_node_4 n_N0858(eclk, ereset, N0858_port_2,N0858_port_3,N0858_port_0,N0858_port_1, N0858_v);
  spice_node_2 n_N0759(eclk, ereset, N0759_port_0,N0759_port_1, N0759_v);
  spice_node_3 n_N0758(eclk, ereset, N0758_port_2,N0758_port_3,N0758_port_1, N0758_v);
  spice_node_2 n_N0757(eclk, ereset, N0757_port_0,N0757_port_1, N0757_v);
  spice_node_3 n_N0756(eclk, ereset, N0756_port_2,N0756_port_0,N0756_port_1, N0756_v);
  spice_node_2 n_N0755(eclk, ereset, N0755_port_0,N0755_port_1, N0755_v);
  spice_node_3 n_N0754(eclk, ereset, N0754_port_2,N0754_port_3,N0754_port_1, N0754_v);
  spice_node_2 n_N0753(eclk, ereset, N0753_port_0,N0753_port_1, N0753_v);
  spice_node_2 n_N0752(eclk, ereset, N0752_port_3,N0752_port_0, N0752_v);
  spice_node_3 n_N0751(eclk, ereset, N0751_port_2,N0751_port_0,N0751_port_1, N0751_v);
  spice_node_3 n_N0750(eclk, ereset, N0750_port_2,N0750_port_0,N0750_port_1, N0750_v);
  spice_node_1 n_S00690(eclk, ereset, S00690_port_1, S00690_v);
  spice_node_2 n_N0920(eclk, ereset, N0920_port_0,N0920_port_1, N0920_v);
  spice_node_3 n_N0339(eclk, ereset, N0339_port_2,N0339_port_0,N0339_port_1, N0339_v);
  spice_node_2 n_N0338(eclk, ereset, N0338_port_0,N0338_port_1, N0338_v);
  spice_node_1 n_S00609(eclk, ereset, S00609_port_0, S00609_v);
  spice_node_2 n_N0802(eclk, ereset, N0802_port_2,N0802_port_1, N0802_v);
  spice_node_2 n_N0801(eclk, ereset, N0801_port_2,N0801_port_1, N0801_v);
  spice_node_2 n_N0800(eclk, ereset, N0800_port_0,N0800_port_1, N0800_v);
  spice_node_2 n_N0807(eclk, ereset, N0807_port_0,N0807_port_1, N0807_v);
  spice_node_2 n_N0806(eclk, ereset, N0806_port_0,N0806_port_1, N0806_v);
  spice_node_2 n_N0805(eclk, ereset, N0805_port_2,N0805_port_1, N0805_v);
  spice_node_2 n_N0804(eclk, ereset, N0804_port_2,N0804_port_3, N0804_v);
  spice_node_1 n_S00601(eclk, ereset, S00601_port_1, S00601_v);
  spice_node_1 n_S00600(eclk, ereset, S00600_port_1, S00600_v);
  spice_node_2 n_N0809(eclk, ereset, N0809_port_0,N0809_port_1, N0809_v);
  spice_node_2 n_N0808(eclk, ereset, N0808_port_0,N0808_port_1, N0808_v);
  spice_node_1 n_S00599(eclk, ereset, S00599_port_1, S00599_v);
  spice_node_1 n_S00598(eclk, ereset, S00598_port_1, S00598_v);
  spice_node_3 n_ADSL(eclk, ereset, ADSL_port_2,ADSL_port_0,ADSL_port_1, ADSL_v);
  spice_node_3 n_A32(eclk, ereset, A32_port_8,A32_port_9,A32_port_6, A32_v);
  spice_node_2 n_N0936(eclk, ereset, N0936_port_0,N0936_port_1, N0936_v);
  spice_node_2 n_N0935(eclk, ereset, N0935_port_0,N0935_port_1, N0935_v);
  spice_node_2 n_N0931(eclk, ereset, N0931_port_0,N0931_port_1, N0931_v);
  spice_node_2 n_N0930(eclk, ereset, N0930_port_0,N0930_port_1, N0930_v);
  spice_node_1 n_S00734(eclk, ereset, S00734_port_1, S00734_v);
  spice_node_1 n_R9_2(eclk, ereset, R9_2_port_1, R9_2_v);
  spice_node_1 n_R9_3(eclk, ereset, R9_3_port_0, R9_3_v);
  spice_node_1 n_R9_0(eclk, ereset, R9_0_port_1, R9_0_v);
  spice_node_1 n_R9_1(eclk, ereset, R9_1_port_0, R9_1_v);
  spice_node_2 n_N0520(eclk, ereset, N0520_port_0,N0520_port_1, N0520_v);
  spice_node_1 n_N0521(eclk, ereset, N0521_port_0, N0521_v);
  spice_node_1 n_S00732(eclk, ereset, S00732_port_1, S00732_v);
  spice_node_5 n_FIN_FIM(eclk, ereset, FIN_FIM_port_2,FIN_FIM_port_3,FIN_FIM_port_0,FIN_FIM_port_4,FIN_FIM_port_5, FIN_FIM_v);
  spice_node_6 n___POC_CLK2_X12_X32__INH(eclk, ereset, __POC_CLK2_X12_X32__INH_port_2,__POC_CLK2_X12_X32__INH_port_3,__POC_CLK2_X12_X32__INH_port_0,__POC_CLK2_X12_X32__INH_port_1,__POC_CLK2_X12_X32__INH_port_4,__POC_CLK2_X12_X32__INH_port_5, __POC_CLK2_X12_X32__INH_v);
  spice_node_4 n_INC_ISZ_ADD_SUB_XCH_LD(eclk, ereset, INC_ISZ_ADD_SUB_XCH_LD_port_2,INC_ISZ_ADD_SUB_XCH_LD_port_3,INC_ISZ_ADD_SUB_XCH_LD_port_4,INC_ISZ_ADD_SUB_XCH_LD_port_5, INC_ISZ_ADD_SUB_XCH_LD_v);
  spice_node_2 n_M12_M22_CLK1__M11_M12_(eclk, ereset, M12_M22_CLK1__M11_M12__port_8,M12_M22_CLK1__M11_M12__port_9, M12_M22_CLK1__M11_M12__v);
  spice_node_1 n_S00828(eclk, ereset, S00828_port_1, S00828_v);
  spice_node_6 n_N0847(eclk, ereset, N0847_port_3,N0847_port_0,N0847_port_1,N0847_port_6,N0847_port_4,N0847_port_5, N0847_v);
  spice_node_3 n_ACC_ADAC(eclk, ereset, ACC_ADAC_port_3,ACC_ADAC_port_0,ACC_ADAC_port_1, ACC_ADAC_v);
  spice_node_2 n__OPA_1(eclk, ereset, _OPA_1_port_8,_OPA_1_port_7, _OPA_1_v);
  spice_node_6 n_IAC(eclk, ereset, IAC_port_2,IAC_port_3,IAC_port_0,IAC_port_1,IAC_port_4,IAC_port_5, IAC_v);
  spice_node_3 n_ADD_ACC(eclk, ereset, ADD_ACC_port_2,ADD_ACC_port_0,ADD_ACC_port_1, ADD_ACC_v);
  spice_node_1 n_N0281(eclk, ereset, N0281_port_1, N0281_v);
  spice_node_1 n_N0283(eclk, ereset, N0283_port_1, N0283_v);
  spice_node_1 n_N0282(eclk, ereset, N0282_port_1, N0282_v);
  spice_node_4 n_ACC_3(eclk, ereset, ACC_3_port_3,ACC_3_port_0,ACC_3_port_1,ACC_3_port_4, ACC_3_v);
  spice_node_4 n_ACC_2(eclk, ereset, ACC_2_port_2,ACC_2_port_3,ACC_2_port_0,ACC_2_port_4, ACC_2_v);
  spice_node_4 n_ACC_1(eclk, ereset, ACC_1_port_3,ACC_1_port_0,ACC_1_port_1,ACC_1_port_4, ACC_1_v);
  spice_node_9 n_ACC_0(eclk, ereset, ACC_0_port_8,ACC_0_port_9,ACC_0_port_2,ACC_0_port_1,ACC_0_port_6,ACC_0_port_7,ACC_0_port_4,ACC_0_port_5,ACC_0_port_10, ACC_0_v);
  spice_node_1 n_N0285(eclk, ereset, N0285_port_1, N0285_v);
  spice_node_1 n_N0287(eclk, ereset, N0287_port_1, N0287_v);
  spice_node_2 n_N0945(eclk, ereset, N0945_port_3,N0945_port_4, N0945_v);
  spice_node_2 n_cm_ram1(eclk, ereset, cm_ram1_port_0,cm_ram1_port_1, cm_ram1_v);
  spice_node_6 n_TCS(eclk, ereset, TCS_port_2,TCS_port_3,TCS_port_0,TCS_port_1,TCS_port_4,TCS_port_5, TCS_v);
  spice_node_2 n_cm_ram3(eclk, ereset, cm_ram3_port_0,cm_ram3_port_1, cm_ram3_v);
  spice_node_2 n_SC_A22(eclk, ereset, SC_A22_port_3,SC_A22_port_4, SC_A22_v);
  spice_node_6 n_TCC(eclk, ereset, TCC_port_2,TCC_port_3,TCC_port_0,TCC_port_1,TCC_port_4,TCC_port_5, TCC_v);
  spice_node_4 n_REG_RFSH_2(eclk, ereset, REG_RFSH_2_port_2,REG_RFSH_2_port_3,REG_RFSH_2_port_0,REG_RFSH_2_port_1, REG_RFSH_2_v);
  spice_node_4 n_REG_RFSH_1(eclk, ereset, REG_RFSH_1_port_2,REG_RFSH_1_port_3,REG_RFSH_1_port_0,REG_RFSH_1_port_1, REG_RFSH_1_v);
  spice_node_4 n_REG_RFSH_0(eclk, ereset, REG_RFSH_0_port_2,REG_RFSH_0_port_3,REG_RFSH_0_port_0,REG_RFSH_0_port_1, REG_RFSH_0_v);
  spice_node_2 n_N0748(eclk, ereset, N0748_port_2,N0748_port_1, N0748_v);
  spice_node_3 n_N0749(eclk, ereset, N0749_port_2,N0749_port_0,N0749_port_1, N0749_v);
  spice_node_2 n_N0740(eclk, ereset, N0740_port_2,N0740_port_1, N0740_v);
  spice_node_2 n_N0741(eclk, ereset, N0741_port_0,N0741_port_1, N0741_v);
  spice_node_2 n_N0742(eclk, ereset, N0742_port_2,N0742_port_1, N0742_v);
  spice_node_2 n_N0743(eclk, ereset, N0743_port_2,N0743_port_1, N0743_v);
  spice_node_2 n_N0744(eclk, ereset, N0744_port_2,N0744_port_1, N0744_v);
  spice_node_2 n_N0745(eclk, ereset, N0745_port_2,N0745_port_1, N0745_v);
  spice_node_2 n_N0746(eclk, ereset, N0746_port_2,N0746_port_1, N0746_v);
  spice_node_2 n_N0747(eclk, ereset, N0747_port_2,N0747_port_1, N0747_v);
  spice_node_3 n_N0670(eclk, ereset, N0670_port_3,N0670_port_0,N0670_port_4, N0670_v);
  spice_node_5 n_CY_1(eclk, ereset, CY_1_port_2,CY_1_port_3,CY_1_port_1,CY_1_port_6,CY_1_port_4, CY_1_v);
  spice_node_3 n_N0674(eclk, ereset, N0674_port_2,N0674_port_0,N0674_port_1, N0674_v);
  spice_node_2 n_N0676(eclk, ereset, N0676_port_0,N0676_port_1, N0676_v);
  spice_node_2 n_N0677(eclk, ereset, N0677_port_0,N0677_port_1, N0677_v);
  spice_node_2 n_N0634(eclk, ereset, N0634_port_8,N0634_port_9, N0634_v);
  spice_node_5 n_N0635(eclk, ereset, N0635_port_3,N0635_port_6,N0635_port_7,N0635_port_4,N0635_port_5, N0635_v);
  spice_node_5 n_N0636(eclk, ereset, N0636_port_2,N0636_port_3,N0636_port_1,N0636_port_4,N0636_port_5, N0636_v);
  spice_node_3 n_N0637(eclk, ereset, N0637_port_2,N0637_port_0,N0637_port_1, N0637_v);
  spice_node_2 n_N0630(eclk, ereset, N0630_port_2,N0630_port_1, N0630_v);
  spice_node_2 n_N0631(eclk, ereset, N0631_port_0,N0631_port_1, N0631_v);
  spice_node_2 n_N0632(eclk, ereset, N0632_port_8,N0632_port_9, N0632_v);
  spice_node_1 n_N0633(eclk, ereset, N0633_port_0, N0633_v);
  spice_node_2 n_N0638(eclk, ereset, N0638_port_0,N0638_port_1, N0638_v);
  spice_node_2 n_N0639(eclk, ereset, N0639_port_0,N0639_port_1, N0639_v);
  spice_node_2 n_N0329(eclk, ereset, N0329_port_0,N0329_port_1, N0329_v);
  spice_node_3 n_N0322(eclk, ereset, N0322_port_2,N0322_port_1,N0322_port_4, N0322_v);
  spice_node_3 n_N0323(eclk, ereset, N0323_port_2,N0323_port_0,N0323_port_1, N0323_v);
  spice_node_2 n_N0320(eclk, ereset, N0320_port_0,N0320_port_1, N0320_v);
  spice_node_2 n_N0321(eclk, ereset, N0321_port_0,N0321_port_1, N0321_v);
  spice_node_5 n_N0326(eclk, ereset, N0326_port_2,N0326_port_3,N0326_port_1,N0326_port_4,N0326_port_5, N0326_v);
  spice_node_2 n_N0324(eclk, ereset, N0324_port_0,N0324_port_1, N0324_v);
  spice_node_1 n_N0325(eclk, ereset, N0325_port_6, N0325_v);
  spice_node_3 n_ACB_IB(eclk, ereset, ACB_IB_port_2,ACB_IB_port_0,ACB_IB_port_1, ACB_IB_v);
  spice_node_2 n_N0818(eclk, ereset, N0818_port_0,N0818_port_1, N0818_v);
  spice_node_2 n_N0814(eclk, ereset, N0814_port_0,N0814_port_1, N0814_v);
  spice_node_1 n_R5_3(eclk, ereset, R5_3_port_0, R5_3_v);
  spice_node_4 n_A22(eclk, ereset, A22_port_8,A22_port_9,A22_port_6,A22_port_5, A22_v);
  spice_node_4 n_N0473(eclk, ereset, N0473_port_2,N0473_port_3,N0473_port_0,N0473_port_1, N0473_v);
  spice_node_2 n_N0921(eclk, ereset, N0921_port_0,N0921_port_1, N0921_v);
  spice_node_2 n_N0922(eclk, ereset, N0922_port_0,N0922_port_1, N0922_v);
  spice_node_2 n_N0923(eclk, ereset, N0923_port_0,N0923_port_1, N0923_v);
  spice_node_2 n_N0924(eclk, ereset, N0924_port_0,N0924_port_1, N0924_v);
  spice_node_2 n_N0925(eclk, ereset, N0925_port_0,N0925_port_1, N0925_v);
  spice_node_2 n_N0926(eclk, ereset, N0926_port_0,N0926_port_1, N0926_v);
  spice_node_2 n_N0927(eclk, ereset, N0927_port_0,N0927_port_1, N0927_v);
  spice_node_2 n_N0928(eclk, ereset, N0928_port_2,N0928_port_3, N0928_v);
  spice_node_2 n_N0929(eclk, ereset, N0929_port_0,N0929_port_1, N0929_v);
  spice_node_1 n_N0697(eclk, ereset, N0697_port_0, N0697_v);
  spice_node_1 n_S00709(eclk, ereset, S00709_port_1, S00709_v);
  spice_node_1 n_R5_1(eclk, ereset, R5_1_port_0, R5_1_v);
  spice_node_3 n_N0690(eclk, ereset, N0690_port_2,N0690_port_0,N0690_port_1, N0690_v);
  spice_node_1 n_N0691(eclk, ereset, N0691_port_0, N0691_v);
  spice_node_1 n_N0694(eclk, ereset, N0694_port_0, N0694_v);
  spice_node_2 n_N0933(eclk, ereset, N0933_port_0,N0933_port_1, N0933_v);
  spice_node_2 n_INH(eclk, ereset, INH_port_2,INH_port_4, INH_v);
  spice_node_3 n_N0913(eclk, ereset, N0913_port_2,N0913_port_0,N0913_port_1, N0913_v);
  spice_node_3 n_N0912(eclk, ereset, N0912_port_2,N0912_port_0,N0912_port_1, N0912_v);
  spice_node_1 n_S00564(eclk, ereset, S00564_port_0, S00564_v);
  spice_node_2 n_N0932(eclk, ereset, N0932_port_0,N0932_port_1, N0932_v);
  spice_node_2 n_N0916(eclk, ereset, N0916_port_0,N0916_port_1, N0916_v);
  spice_node_3 n_N0693(eclk, ereset, N0693_port_2,N0693_port_3,N0693_port_1, N0693_v);
  spice_node_2 n_N0820(eclk, ereset, N0820_port_2,N0820_port_3, N0820_v);
  spice_node_1 n_PC1_1(eclk, ereset, PC1_1_port_1, PC1_1_v);
  spice_node_1 n_PC1_2(eclk, ereset, PC1_2_port_0, PC1_2_v);
  spice_node_1 n_PC1_3(eclk, ereset, PC1_3_port_1, PC1_3_v);
  spice_node_1 n_PC1_4(eclk, ereset, PC1_4_port_1, PC1_4_v);
  spice_node_1 n_PC1_5(eclk, ereset, PC1_5_port_0, PC1_5_v);
  spice_node_1 n_PC1_6(eclk, ereset, PC1_6_port_1, PC1_6_v);
  spice_node_1 n_PC1_7(eclk, ereset, PC1_7_port_0, PC1_7_v);
  spice_node_1 n_PC1_8(eclk, ereset, PC1_8_port_0, PC1_8_v);
  spice_node_1 n_PC1_9(eclk, ereset, PC1_9_port_1, PC1_9_v);
  spice_node_2 n_N0822(eclk, ereset, N0822_port_0,N0822_port_1, N0822_v);
  spice_node_1 n_PC3_6(eclk, ereset, PC3_6_port_1, PC3_6_v);
  spice_node_1 n_PC3_7(eclk, ereset, PC3_7_port_0, PC3_7_v);
  spice_node_1 n_PC3_4(eclk, ereset, PC3_4_port_1, PC3_4_v);
  spice_node_1 n_PC3_5(eclk, ereset, PC3_5_port_0, PC3_5_v);
  spice_node_1 n_PC3_2(eclk, ereset, PC3_2_port_0, PC3_2_v);
  spice_node_1 n_PC3_3(eclk, ereset, PC3_3_port_1, PC3_3_v);
  spice_node_1 n_PC3_0(eclk, ereset, PC3_0_port_0, PC3_0_v);
  spice_node_1 n_PC3_1(eclk, ereset, PC3_1_port_1, PC3_1_v);
  spice_node_1 n_S00803(eclk, ereset, S00803_port_1, S00803_v);
  spice_node_1 n_PC3_8(eclk, ereset, PC3_8_port_0, PC3_8_v);
  spice_node_1 n_PC3_9(eclk, ereset, PC3_9_port_1, PC3_9_v);
  spice_node_4 n_N0900(eclk, ereset, N0900_port_2,N0900_port_3,N0900_port_0,N0900_port_1, N0900_v);
  spice_node_2 n_N0353(eclk, ereset, N0353_port_2,N0353_port_1, N0353_v);
  spice_node_2 n_N0352(eclk, ereset, N0352_port_0,N0352_port_1, N0352_v);
  spice_node_3 n_N0351(eclk, ereset, N0351_port_2,N0351_port_0,N0351_port_1, N0351_v);
  spice_node_2 n_N0350(eclk, ereset, N0350_port_0,N0350_port_1, N0350_v);
  spice_node_3 n_N0608(eclk, ereset, N0608_port_2,N0608_port_0,N0608_port_1, N0608_v);
  spice_node_3 n_N0355(eclk, ereset, N0355_port_3,N0355_port_0,N0355_port_1, N0355_v);
  spice_node_6 n_N0354(eclk, ereset, N0354_port_2,N0354_port_3,N0354_port_0,N0354_port_1,N0354_port_4,N0354_port_5, N0354_v);
  spice_node_2 n_N0605(eclk, ereset, N0605_port_0,N0605_port_1, N0605_v);
  spice_node_2 n_N0604(eclk, ereset, N0604_port_0,N0604_port_1, N0604_v);
  spice_node_2 n_N0607(eclk, ereset, N0607_port_0,N0607_port_1, N0607_v);
  spice_node_3 n_ADC_CY(eclk, ereset, ADC_CY_port_2,ADC_CY_port_3,ADC_CY_port_1, ADC_CY_v);
  spice_node_2 n_OPR_3(eclk, ereset, OPR_3_port_14,OPR_3_port_15, OPR_3_v);
  spice_node_1 n_N0852(eclk, ereset, N0852_port_1, N0852_v);
  spice_node_2 n_N0938(eclk, ereset, N0938_port_2,N0938_port_3, N0938_v);
  spice_node_2 n_N0824(eclk, ereset, N0824_port_0,N0824_port_1, N0824_v);
  spice_node_3 n_ADD_IB(eclk, ereset, ADD_IB_port_2,ADD_IB_port_0,ADD_IB_port_1, ADD_IB_v);
  spice_node_2 n_N0823(eclk, ereset, N0823_port_0,N0823_port_1, N0823_v);
  spice_node_1 n_PC2_9(eclk, ereset, PC2_9_port_1, PC2_9_v);
  spice_node_1 n_PC2_8(eclk, ereset, PC2_8_port_0, PC2_8_v);
  spice_node_1 n_PC2_7(eclk, ereset, PC2_7_port_0, PC2_7_v);
  spice_node_1 n_PC2_6(eclk, ereset, PC2_6_port_1, PC2_6_v);
  spice_node_1 n_PC2_5(eclk, ereset, PC2_5_port_0, PC2_5_v);
  spice_node_1 n_PC2_4(eclk, ereset, PC2_4_port_1, PC2_4_v);
  spice_node_1 n_PC2_3(eclk, ereset, PC2_3_port_1, PC2_3_v);
  spice_node_1 n_PC2_2(eclk, ereset, PC2_2_port_0, PC2_2_v);
  spice_node_1 n_PC2_1(eclk, ereset, PC2_1_port_1, PC2_1_v);
  spice_node_1 n_PC2_0(eclk, ereset, PC2_0_port_0, PC2_0_v);
  spice_node_2 n_N0793(eclk, ereset, N0793_port_0,N0793_port_1, N0793_v);
  spice_node_2 n_N0792(eclk, ereset, N0792_port_0,N0792_port_1, N0792_v);
  spice_node_2 n_N0791(eclk, ereset, N0791_port_0,N0791_port_1, N0791_v);
  spice_node_2 n_N0790(eclk, ereset, N0790_port_0,N0790_port_1, N0790_v);
  spice_node_2 n_N0797(eclk, ereset, N0797_port_2,N0797_port_1, N0797_v);
  spice_node_2 n_N0796(eclk, ereset, N0796_port_0,N0796_port_1, N0796_v);
  spice_node_2 n_N0795(eclk, ereset, N0795_port_0,N0795_port_1, N0795_v);
  spice_node_2 n_N0794(eclk, ereset, N0794_port_0,N0794_port_1, N0794_v);
  spice_node_2 n_N0829(eclk, ereset, N0829_port_0,N0829_port_1, N0829_v);
  spice_node_2 n_N0799(eclk, ereset, N0799_port_0,N0799_port_1, N0799_v);
  spice_node_2 n_N0798(eclk, ereset, N0798_port_0,N0798_port_1, N0798_v);
  spice_node_2 n_N0828(eclk, ereset, N0828_port_0,N0828_port_1, N0828_v);
  spice_node_2 n___X31__CLK2_(eclk, ereset, __X31__CLK2__port_2,__X31__CLK2__port_1, __X31__CLK2__v);
  spice_node_3 n_clk1(eclk, ereset, clk1_port_0,clk1_port_1,clk1_port_28, clk1_v);
  spice_node_2 n_clk2(eclk, ereset, clk2_port_51,clk2_port_0, clk2_v);
  spice_node_1 n_N0317(eclk, ereset, N0317_port_0, N0317_v);
  spice_node_3 n_N0316(eclk, ereset, N0316_port_2,N0316_port_0,N0316_port_1, N0316_v);
  spice_node_1 n_N0315(eclk, ereset, N0315_port_0, N0315_v);
  spice_node_2 n_N0645(eclk, ereset, N0645_port_8,N0645_port_9, N0645_v);
  spice_node_2 n_N0312(eclk, ereset, N0312_port_0,N0312_port_1, N0312_v);
  spice_node_2 n_N0647(eclk, ereset, N0647_port_8,N0647_port_9, N0647_v);
  spice_node_2 n_N0310(eclk, ereset, N0310_port_3,N0310_port_4, N0310_v);
  spice_node_2 n_N0649(eclk, ereset, N0649_port_2,N0649_port_1, N0649_v);
  spice_node_5 n_N0648(eclk, ereset, N0648_port_3,N0648_port_6,N0648_port_7,N0648_port_4,N0648_port_5, N0648_v);
  spice_node_1 n_S00840(eclk, ereset, S00840_port_1, S00840_v);
  spice_node_2 n_N0319(eclk, ereset, N0319_port_0,N0319_port_1, N0319_v);
  spice_node_5 n_N0318(eclk, ereset, N0318_port_2,N0318_port_3,N0318_port_1,N0318_port_4,N0318_port_5, N0318_v);
  spice_node_2 n_N0487(eclk, ereset, N0487_port_2,N0487_port_1, N0487_v);
  spice_node_2 n_N0485(eclk, ereset, N0485_port_0,N0485_port_1, N0485_v);
  spice_node_2 n_N0484(eclk, ereset, N0484_port_0,N0484_port_1, N0484_v);
  spice_node_2 n_N0483(eclk, ereset, N0483_port_0,N0483_port_1, N0483_v);
  spice_node_2 n_N0482(eclk, ereset, N0482_port_0,N0482_port_1, N0482_v);
  spice_node_4 n_N0481(eclk, ereset, N0481_port_2,N0481_port_3,N0481_port_0,N0481_port_1, N0481_v);
  spice_node_2 n_N0480(eclk, ereset, N0480_port_0,N0480_port_1, N0480_v);
  spice_node_3 n_WADB2(eclk, ereset, WADB2_port_6,WADB2_port_4,WADB2_port_5, WADB2_v);
  spice_node_3 n_WADB1(eclk, ereset, WADB1_port_6,WADB1_port_4,WADB1_port_5, WADB1_v);
  spice_node_3 n_WADB0(eclk, ereset, WADB0_port_6,WADB0_port_4,WADB0_port_5, WADB0_v);
  spice_node_1 n_N0489(eclk, ereset, N0489_port_0, N0489_v);
  spice_node_2 n_N0488(eclk, ereset, N0488_port_0,N0488_port_1, N0488_v);
  spice_node_10 n_N0869(eclk, ereset, N0869_port_8,N0869_port_9,N0869_port_2,N0869_port_3,N0869_port_0,N0869_port_6,N0869_port_7,N0869_port_4,N0869_port_5,N0869_port_10, N0869_v);
  spice_node_10 n_N0868(eclk, ereset, N0868_port_8,N0868_port_9,N0868_port_2,N0868_port_3,N0868_port_0,N0868_port_6,N0868_port_7,N0868_port_4,N0868_port_5,N0868_port_10, N0868_v);
  spice_node_10 n_N0867(eclk, ereset, N0867_port_8,N0867_port_9,N0867_port_2,N0867_port_3,N0867_port_0,N0867_port_6,N0867_port_7,N0867_port_4,N0867_port_5,N0867_port_10, N0867_v);
  spice_node_2 n_N0853(eclk, ereset, N0853_port_0,N0853_port_1, N0853_v);
  spice_node_3 n_A12(eclk, ereset, A12_port_9,A12_port_7,A12_port_10, A12_v);
  spice_node_1 n_S00716(eclk, ereset, S00716_port_1, S00716_v);
  spice_node_1 n_S00710(eclk, ereset, S00710_port_0, S00710_v);
  spice_node_2 n___INH__X32_CLK2(eclk, ereset, __INH__X32_CLK2_port_2,__INH__X32_CLK2_port_3, __INH__X32_CLK2_v);
  spice_node_1 n_S00620(eclk, ereset, S00620_port_1, S00620_v);
  spice_node_1 n_S00627(eclk, ereset, S00627_port_1, S00627_v);
  spice_node_1 n_S00624(eclk, ereset, S00624_port_1, S00624_v);
  spice_node_1 n_S00628(eclk, ereset, S00628_port_0, S00628_v);
  spice_node_2 n_N0684(eclk, ereset, N0684_port_0,N0684_port_1, N0684_v);
  spice_node_1 n_N0850(eclk, ereset, N0850_port_1, N0850_v);
  spice_node_2 n_N0507(eclk, ereset, N0507_port_0,N0507_port_1, N0507_v);
  spice_node_3 n_N0346(eclk, ereset, N0346_port_3,N0346_port_0,N0346_port_1, N0346_v);
  spice_node_1 n_N0504(eclk, ereset, N0504_port_0, N0504_v);
  spice_node_3 n_N0505(eclk, ereset, N0505_port_2,N0505_port_0,N0505_port_1, N0505_v);
  spice_node_2 n_SC_M22_CLK2(eclk, ereset, SC_M22_CLK2_port_3,SC_M22_CLK2_port_4, SC_M22_CLK2_v);
  spice_node_3 n_N0503(eclk, ereset, N0503_port_2,N0503_port_0,N0503_port_1, N0503_v);
  spice_node_1 n_N0500(eclk, ereset, N0500_port_1, N0500_v);
  spice_node_2 n_N0501(eclk, ereset, N0501_port_0,N0501_port_1, N0501_v);
  spice_node_5 n_ADD_0(eclk, ereset, ADD_0_port_2,ADD_0_port_3,ADD_0_port_1,ADD_0_port_4,ADD_0_port_5, ADD_0_v);
  spice_node_2 n__I_O(eclk, ereset, _I_O_port_0,_I_O_port_1, _I_O_v);
  spice_node_5 n_d0(eclk, ereset, d0_port_2,d0_port_3,d0_port_0,d0_port_4,d0_port_5, d0_v);
  spice_node_5 n_d1(eclk, ereset, d1_port_2,d1_port_3,d1_port_0,d1_port_4,d1_port_5, d1_v);
  spice_node_3 n_N0347(eclk, ereset, N0347_port_3,N0347_port_1,N0347_port_4, N0347_v);
  spice_node_1 n_N1013(eclk, ereset, N1013_port_1, N1013_v);
  spice_node_1 n_N1012(eclk, ereset, N1012_port_1, N1012_v);
  spice_node_1 n_N1011(eclk, ereset, N1011_port_0, N1011_v);
  spice_node_1 n_N1010(eclk, ereset, N1010_port_0, N1010_v);
  spice_node_1 n_N1015(eclk, ereset, N1015_port_1, N1015_v);
  spice_node_1 n_N1014(eclk, ereset, N1014_port_1, N1014_v);
  spice_node_1 n_R15_0(eclk, ereset, R15_0_port_1, R15_0_v);
  spice_node_1 n_R15_1(eclk, ereset, R15_1_port_0, R15_1_v);
  spice_node_1 n_R15_2(eclk, ereset, R15_2_port_1, R15_2_v);
  spice_node_1 n_R15_3(eclk, ereset, R15_3_port_0, R15_3_v);
  spice_node_3 n_N0937(eclk, ereset, N0937_port_0,N0937_port_1,N0937_port_6, N0937_v);
  spice_node_1 n_R11_0(eclk, ereset, R11_0_port_1, R11_0_v);
  spice_node_1 n_R11_1(eclk, ereset, R11_1_port_0, R11_1_v);
  spice_node_1 n_R11_2(eclk, ereset, R11_2_port_1, R11_2_v);
  spice_node_1 n_R11_3(eclk, ereset, R11_3_port_0, R11_3_v);
  spice_node_1 n_R13_2(eclk, ereset, R13_2_port_1, R13_2_v);
  spice_node_1 n_R13_3(eclk, ereset, R13_3_port_0, R13_3_v);
  spice_node_1 n_R13_0(eclk, ereset, R13_0_port_1, R13_0_v);
  spice_node_1 n_R13_1(eclk, ereset, R13_1_port_0, R13_1_v);
  spice_node_2 n_OPR_1(eclk, ereset, OPR_1_port_9,OPR_1_port_10, OPR_1_v);
  spice_node_2 n_OPR_0(eclk, ereset, OPR_0_port_3,OPR_0_port_6, OPR_0_v);
  spice_node_2 n_OPR_2(eclk, ereset, OPR_2_port_8,OPR_2_port_14, OPR_2_v);
  spice_node_2 n_N0340(eclk, ereset, N0340_port_2,N0340_port_0, N0340_v);
  spice_node_4 n_N0859(eclk, ereset, N0859_port_2,N0859_port_3,N0859_port_1,N0859_port_4, N0859_v);
  spice_node_1 n_N0688(eclk, ereset, N0688_port_0, N0688_v);
  spice_node_2 n_N0788(eclk, ereset, N0788_port_0,N0788_port_1, N0788_v);
  spice_node_2 n_N0789(eclk, ereset, N0789_port_0,N0789_port_1, N0789_v);
  spice_node_2 n_N0784(eclk, ereset, N0784_port_0,N0784_port_1, N0784_v);
  spice_node_2 n_N0785(eclk, ereset, N0785_port_0,N0785_port_1, N0785_v);
  spice_node_2 n_N0786(eclk, ereset, N0786_port_0,N0786_port_1, N0786_v);
  spice_node_2 n_N0787(eclk, ereset, N0787_port_0,N0787_port_1, N0787_v);
  spice_node_6 n_N0780(eclk, ereset, N0780_port_2,N0780_port_3,N0780_port_0,N0780_port_6,N0780_port_4,N0780_port_5, N0780_v);
  spice_node_6 n_N0781(eclk, ereset, N0781_port_2,N0781_port_3,N0781_port_0,N0781_port_6,N0781_port_4,N0781_port_5, N0781_v);
  spice_node_4 n_N0782(eclk, ereset, N0782_port_2,N0782_port_3,N0782_port_4,N0782_port_5, N0782_v);
  spice_node_2 n_N0783(eclk, ereset, N0783_port_2,N0783_port_3, N0783_v);
  spice_node_2 n_N0300(eclk, ereset, N0300_port_3,N0300_port_4, N0300_v);
  spice_node_2 n_N0301(eclk, ereset, N0301_port_2,N0301_port_3, N0301_v);
  spice_node_2 n_N0302(eclk, ereset, N0302_port_0,N0302_port_1, N0302_v);
  spice_node_2 n_N0303(eclk, ereset, N0303_port_0,N0303_port_1, N0303_v);
  spice_node_3 n_N0304(eclk, ereset, N0304_port_2,N0304_port_3,N0304_port_1, N0304_v);
  spice_node_3 n_N0305(eclk, ereset, N0305_port_2,N0305_port_0,N0305_port_1, N0305_v);
  spice_node_2 n_N0306(eclk, ereset, N0306_port_0,N0306_port_1, N0306_v);
  spice_node_3 n_N0307(eclk, ereset, N0307_port_3,N0307_port_4,N0307_port_5, N0307_v);
  spice_node_2 n_N0308(eclk, ereset, N0308_port_0,N0308_port_1, N0308_v);
  spice_node_2 n_N0309(eclk, ereset, N0309_port_0,N0309_port_1, N0309_v);
  spice_node_3 n_N0658(eclk, ereset, N0658_port_3,N0658_port_0,N0658_port_1, N0658_v);
  spice_node_2 n_N0659(eclk, ereset, N0659_port_4,N0659_port_5, N0659_v);
  spice_node_2 n_N0490(eclk, ereset, N0490_port_2,N0490_port_0, N0490_v);
  spice_node_2 n_N0491(eclk, ereset, N0491_port_0,N0491_port_1, N0491_v);
  spice_node_1 n_N0492(eclk, ereset, N0492_port_0, N0492_v);
  spice_node_2 n_N0493(eclk, ereset, N0493_port_0,N0493_port_1, N0493_v);
  spice_node_2 n_N0494(eclk, ereset, N0494_port_2,N0494_port_0, N0494_v);
  spice_node_2 n_N0495(eclk, ereset, N0495_port_0,N0495_port_1, N0495_v);
  spice_node_2 n_N0496(eclk, ereset, N0496_port_0,N0496_port_1, N0496_v);
  spice_node_1 n_N0497(eclk, ereset, N0497_port_0, N0497_v);
  spice_node_1 n_N0498(eclk, ereset, N0498_port_1, N0498_v);
  spice_node_1 n_N0499(eclk, ereset, N0499_port_0, N0499_v);
  spice_node_3 n_N0878(eclk, ereset, N0878_port_2,N0878_port_3,N0878_port_4, N0878_v);
  spice_node_3 n_N0879(eclk, ereset, N0879_port_3,N0879_port_1,N0879_port_4, N0879_v);
  spice_node_1 n_N0653(eclk, ereset, N0653_port_0, N0653_v);
  spice_node_2 n_N0651(eclk, ereset, N0651_port_0,N0651_port_1, N0651_v);
  spice_node_2 n_N0656(eclk, ereset, N0656_port_0,N0656_port_1, N0656_v);
  spice_node_4 n_X12(eclk, ereset, X12_port_10,X12_port_12,X12_port_13,X12_port_15, X12_v);
  spice_node_2 n_N0657(eclk, ereset, N0657_port_8,N0657_port_9, N0657_v);
  spice_node_3 n_N0654(eclk, ereset, N0654_port_2,N0654_port_0,N0654_port_1, N0654_v);
  spice_node_2 n_N0655(eclk, ereset, N0655_port_2,N0655_port_1, N0655_v);
  spice_node_1 n_S00762(eclk, ereset, S00762_port_1, S00762_v);
  spice_node_6 n_RAL(eclk, ereset, RAL_port_2,RAL_port_3,RAL_port_0,RAL_port_1,RAL_port_4,RAL_port_5, RAL_v);
  spice_node_6 n_RAR(eclk, ereset, RAR_port_2,RAR_port_3,RAR_port_0,RAR_port_1,RAR_port_4,RAR_port_5, RAR_v);
  spice_node_5 n_N0716(eclk, ereset, N0716_port_2,N0716_port_3,N0716_port_0,N0716_port_1,N0716_port_4, N0716_v);
  spice_node_2 n_N0313(eclk, ereset, N0313_port_0,N0313_port_1, N0313_v);
  spice_node_3 n_OPA_2(eclk, ereset, OPA_2_port_0,OPA_2_port_4,OPA_2_port_13, OPA_2_v);
  spice_node_3 n_OPA_3(eclk, ereset, OPA_3_port_2,OPA_3_port_0,OPA_3_port_13, OPA_3_v);
  spice_node_3 n_OPA_0(eclk, ereset, OPA_0_port_11,OPA_0_port_12,OPA_0_port_13, OPA_0_v);
  spice_node_2 n__INH(eclk, ereset, _INH_port_0,_INH_port_1, _INH_v);
  spice_node_2 n_N0934(eclk, ereset, N0934_port_0,N0934_port_1, N0934_v);
  spice_node_6 n_STC(eclk, ereset, STC_port_2,STC_port_3,STC_port_0,STC_port_1,STC_port_4,STC_port_5, STC_v);
  spice_node_3 n_N0873(eclk, ereset, N0873_port_0,N0873_port_4,N0873_port_5, N0873_v);
  spice_node_3 n_N0870(eclk, ereset, N0870_port_2,N0870_port_0,N0870_port_6, N0870_v);
  spice_node_4 n_FIN_FIM_SRC_JIN(eclk, ereset, FIN_FIM_SRC_JIN_port_3,FIN_FIM_SRC_JIN_port_6,FIN_FIM_SRC_JIN_port_4,FIN_FIM_SRC_JIN_port_5, FIN_FIM_SRC_JIN_v);
  spice_node_3 n_N0871(eclk, ereset, N0871_port_0,N0871_port_6,N0871_port_5, N0871_v);
  spice_node_2 n_N0876(eclk, ereset, N0876_port_2,N0876_port_1, N0876_v);
  spice_node_3 n_N0877(eclk, ereset, N0877_port_2,N0877_port_3,N0877_port_4, N0877_v);
  spice_node_2 n_N0874(eclk, ereset, N0874_port_2,N0874_port_1, N0874_v);
  spice_node_1 n_N1008(eclk, ereset, N1008_port_1, N1008_v);
  spice_node_1 n_N1009(eclk, ereset, N1009_port_0, N1009_v);
  spice_node_2 n_N1004(eclk, ereset, N1004_port_3,N1004_port_4, N1004_v);
  spice_node_2 n_N1005(eclk, ereset, N1005_port_2,N1005_port_3, N1005_v);
  spice_node_2 n_N1006(eclk, ereset, N1006_port_3,N1006_port_4, N1006_v);
  spice_node_2 n_N1007(eclk, ereset, N1007_port_2,N1007_port_3, N1007_v);
  spice_node_2 n_N1000(eclk, ereset, N1000_port_3,N1000_port_4, N1000_v);
  spice_node_2 n_N1001(eclk, ereset, N1001_port_2,N1001_port_3, N1001_v);
  spice_node_2 n_N1002(eclk, ereset, N1002_port_3,N1002_port_4, N1002_v);
  spice_node_2 n_N1003(eclk, ereset, N1003_port_2,N1003_port_3, N1003_v);
  spice_node_3 n_OPA_1(eclk, ereset, OPA_1_port_10,OPA_1_port_11,OPA_1_port_12, OPA_1_v);
  spice_node_1 n_PC3_10(eclk, ereset, PC3_10_port_0, PC3_10_v);
  spice_node_1 n_PC3_11(eclk, ereset, PC3_11_port_1, PC3_11_v);
  spice_node_5 n_FIM_SRC(eclk, ereset, FIM_SRC_port_2,FIM_SRC_port_3,FIM_SRC_port_0,FIM_SRC_port_1,FIM_SRC_port_4, FIM_SRC_v);
  spice_node_4 n_ADDR_RFSH_1(eclk, ereset, ADDR_RFSH_1_port_2,ADDR_RFSH_1_port_3,ADDR_RFSH_1_port_0,ADDR_RFSH_1_port_1, ADDR_RFSH_1_v);
  spice_node_4 n_ADDR_RFSH_0(eclk, ereset, ADDR_RFSH_0_port_2,ADDR_RFSH_0_port_3,ADDR_RFSH_0_port_0,ADDR_RFSH_0_port_1, ADDR_RFSH_0_v);
  spice_node_1 n_S00778(eclk, ereset, S00778_port_0, S00778_v);
  spice_node_3 n_N0375(eclk, ereset, N0375_port_3,N0375_port_0,N0375_port_1, N0375_v);
  spice_node_1 n_N0374(eclk, ereset, N0374_port_1, N0374_v);
  spice_node_3 n_N0696(eclk, ereset, N0696_port_2,N0696_port_3,N0696_port_0, N0696_v);
  spice_node_2 n_N0377(eclk, ereset, N0377_port_0,N0377_port_1, N0377_v);
  spice_node_6 n_N0376(eclk, ereset, N0376_port_2,N0376_port_3,N0376_port_0,N0376_port_1,N0376_port_4,N0376_port_5, N0376_v);
  spice_node_1 n_N0278(eclk, ereset, N0278_port_1, N0278_v);
  spice_node_4 n_N0279(eclk, ereset, N0279_port_2,N0279_port_3,N0279_port_0,N0279_port_1, N0279_v);
  spice_node_3 n_DCL_1(eclk, ereset, DCL_1_port_2,DCL_1_port_3,DCL_1_port_1, DCL_1_v);
  spice_node_3 n_DCL_0(eclk, ereset, DCL_0_port_3,DCL_0_port_0,DCL_0_port_4, DCL_0_v);
  spice_node_3 n_DCL_2(eclk, ereset, DCL_2_port_2,DCL_2_port_3,DCL_2_port_1, DCL_2_v);
  spice_node_4 n_N0373(eclk, ereset, N0373_port_2,N0373_port_3,N0373_port_0,N0373_port_1, N0373_v);
  spice_node_4 n_N0372(eclk, ereset, N0372_port_2,N0372_port_3,N0372_port_0,N0372_port_1, N0372_v);
  spice_node_3 n_N0669(eclk, ereset, N0669_port_3,N0669_port_0,N0669_port_1, N0669_v);
  spice_node_3 n_N0667(eclk, ereset, N0667_port_2,N0667_port_0,N0667_port_1, N0667_v);
  spice_node_3 n_N0666(eclk, ereset, N0666_port_2,N0666_port_3,N0666_port_4, N0666_v);
  spice_node_3 n_N0665(eclk, ereset, N0665_port_2,N0665_port_0,N0665_port_1, N0665_v);
  spice_node_3 n_N0664(eclk, ereset, N0664_port_2,N0664_port_1,N0664_port_4, N0664_v);
  spice_node_3 n_N0663(eclk, ereset, N0663_port_2,N0663_port_3,N0663_port_1, N0663_v);
  spice_node_2 n_N0662(eclk, ereset, N0662_port_0,N0662_port_1, N0662_v);
  spice_node_2 n_N0661(eclk, ereset, N0661_port_0,N0661_port_1, N0661_v);
  spice_node_2 n_N0660(eclk, ereset, N0660_port_0,N0660_port_1, N0660_v);
  spice_node_3 n_N0469(eclk, ereset, N0469_port_0,N0469_port_1,N0469_port_4, N0469_v);
  spice_node_4 n_N0468(eclk, ereset, N0468_port_2,N0468_port_3,N0468_port_0,N0468_port_1, N0468_v);
  spice_node_2 n_N0465(eclk, ereset, N0465_port_0,N0465_port_1, N0465_v);
  spice_node_3 n_N0464(eclk, ereset, N0464_port_2,N0464_port_3,N0464_port_4, N0464_v);
  spice_node_1 n_PC1_10(eclk, ereset, PC1_10_port_0, PC1_10_v);
  spice_node_1 n_PC1_11(eclk, ereset, PC1_11_port_1, PC1_11_v);
  spice_node_3 n_N0461(eclk, ereset, N0461_port_2,N0461_port_1,N0461_port_4, N0461_v);
  spice_node_2 n_N0460(eclk, ereset, N0460_port_0,N0460_port_1, N0460_v);
  spice_node_3 n_N0463(eclk, ereset, N0463_port_2,N0463_port_3,N0463_port_6, N0463_v);
  spice_node_2 n_N0462(eclk, ereset, N0462_port_0,N0462_port_1, N0462_v);
  spice_node_1 n_N0685(eclk, ereset, N0685_port_0, N0685_v);
  spice_node_3 n_N0687(eclk, ereset, N0687_port_2,N0687_port_0,N0687_port_1, N0687_v);
  spice_node_2 n_N0681(eclk, ereset, N0681_port_0,N0681_port_1, N0681_v);
  spice_node_2 n_N0680(eclk, ereset, N0680_port_0,N0680_port_1, N0680_v);
  spice_node_3 n_N0683(eclk, ereset, N0683_port_2,N0683_port_0,N0683_port_1, N0683_v);
  spice_node_1 n_S00557(eclk, ereset, S00557_port_1, S00557_v);
  spice_node_3 n_N0689(eclk, ereset, N0689_port_2,N0689_port_0,N0689_port_1, N0689_v);
  spice_node_3 n_X22(eclk, ereset, X22_port_6,X22_port_7,X22_port_5, X22_v);
  spice_node_2 n_N0398(eclk, ereset, N0398_port_0,N0398_port_1, N0398_v);
  spice_node_1 n_R12_2(eclk, ereset, R12_2_port_0, R12_2_v);
  spice_node_1 n_R12_1(eclk, ereset, R12_1_port_1, R12_1_v);
  spice_node_6 n_N0846(eclk, ereset, N0846_port_2,N0846_port_0,N0846_port_1,N0846_port_6,N0846_port_4,N0846_port_5, N0846_v);
  spice_node_2 n_N0843(eclk, ereset, N0843_port_0,N0843_port_1, N0843_v);
  spice_node_2 n_N0841(eclk, ereset, N0841_port_0,N0841_port_1, N0841_v);
  spice_node_2 n_N0840(eclk, ereset, N0840_port_0,N0840_port_1, N0840_v);
  spice_node_1 n_N0519(eclk, ereset, N0519_port_0, N0519_v);
  spice_node_2 n_N0518(eclk, ereset, N0518_port_0,N0518_port_1, N0518_v);
  spice_node_3 n_N0692(eclk, ereset, N0692_port_2,N0692_port_0,N0692_port_1, N0692_v);
  spice_node_5 n_OPE(eclk, ereset, OPE_port_2,OPE_port_3,OPE_port_0,OPE_port_1,OPE_port_4, OPE_v);
  spice_node_3 n_N0695(eclk, ereset, N0695_port_2,N0695_port_3,N0695_port_1, N0695_v);
  spice_node_2 n_N0686(eclk, ereset, N0686_port_0,N0686_port_1, N0686_v);
  spice_node_5 n_JCN(eclk, ereset, JCN_port_2,JCN_port_3,JCN_port_0,JCN_port_1,JCN_port_4, JCN_v);
  spice_node_4 n_N0678(eclk, ereset, N0678_port_3,N0678_port_0,N0678_port_1,N0678_port_4, N0678_v);
  spice_node_2 n_N0679(eclk, ereset, N0679_port_2,N0679_port_0, N0679_v);
  spice_node_3 n_N0671(eclk, ereset, N0671_port_2,N0671_port_0,N0671_port_1, N0671_v);
  spice_node_3 n_N0672(eclk, ereset, N0672_port_2,N0672_port_0,N0672_port_1, N0672_v);
  spice_node_3 n_N0673(eclk, ereset, N0673_port_2,N0673_port_0,N0673_port_1, N0673_v);
  spice_node_3 n_N0675(eclk, ereset, N0675_port_2,N0675_port_3,N0675_port_0, N0675_v);
  spice_node_5 n_N0478(eclk, ereset, N0478_port_2,N0478_port_3,N0478_port_0,N0478_port_1,N0478_port_4, N0478_v);
  spice_node_2 n_N0479(eclk, ereset, N0479_port_2,N0479_port_0, N0479_v);
  spice_node_2 n_N0476(eclk, ereset, N0476_port_2,N0476_port_0, N0476_v);
  spice_node_3 n_N0477(eclk, ereset, N0477_port_2,N0477_port_0,N0477_port_1, N0477_v);
  spice_node_4 n_N0474(eclk, ereset, N0474_port_2,N0474_port_3,N0474_port_0,N0474_port_1, N0474_v);
  spice_node_3 n_N0475(eclk, ereset, N0475_port_0,N0475_port_1,N0475_port_4, N0475_v);
  spice_node_4 n_N0472(eclk, ereset, N0472_port_2,N0472_port_3,N0472_port_0,N0472_port_1, N0472_v);
  spice_node_4 n_N0470(eclk, ereset, N0470_port_2,N0470_port_3,N0470_port_0,N0470_port_1, N0470_v);
  spice_node_4 n_N0471(eclk, ereset, N0471_port_2,N0471_port_3,N0471_port_0,N0471_port_1, N0471_v);
  spice_node_2 n_X32(eclk, ereset, X32_port_11,X32_port_12, X32_v);
  spice_node_3 n_N0698(eclk, ereset, N0698_port_2,N0698_port_3,N0698_port_1, N0698_v);
  spice_node_1 n_N0699(eclk, ereset, N0699_port_1, N0699_v);
  spice_node_3 n_CLK2_JMS_DC_M22_BBL_M22_X12_X22__(eclk, ereset, CLK2_JMS_DC_M22_BBL_M22_X12_X22___port_2,CLK2_JMS_DC_M22_BBL_M22_X12_X22___port_3,CLK2_JMS_DC_M22_BBL_M22_X12_X22___port_4, CLK2_JMS_DC_M22_BBL_M22_X12_X22___v);
  spice_node_1 n_N0506(eclk, ereset, N0506_port_0, N0506_v);
  spice_node_2 n_N0508(eclk, ereset, N0508_port_0,N0508_port_1, N0508_v);
  spice_node_2 n_N0509(eclk, ereset, N0509_port_0,N0509_port_1, N0509_v);
  spice_node_1 n_S00740(eclk, ereset, S00740_port_0, S00740_v);
  spice_node_3 n_N0328(eclk, ereset, N0328_port_2,N0328_port_0,N0328_port_1, N0328_v);
  spice_node_1 n_S00766(eclk, ereset, S00766_port_0, S00766_v);
  spice_node_3 n_N0551(eclk, ereset, N0551_port_2,N0551_port_0,N0551_port_1, N0551_v);
  spice_node_1 n_S00767(eclk, ereset, S00767_port_0, S00767_v);
  spice_node_4 n_N0550(eclk, ereset, N0550_port_2,N0550_port_3,N0550_port_0,N0550_port_1, N0550_v);
  spice_node_3 n_N0327(eclk, ereset, N0327_port_3,N0327_port_0,N0327_port_4, N0327_v);
  spice_node_1 n_S00764(eclk, ereset, S00764_port_1, S00764_v);
  spice_node_2 n_N0553(eclk, ereset, N0553_port_2,N0553_port_1, N0553_v);
  spice_node_2 n_N0955(eclk, ereset, N0955_port_2,N0955_port_3, N0955_v);
  spice_node_2 n_N0954(eclk, ereset, N0954_port_0,N0954_port_1, N0954_v);
  spice_node_2 n_N0957(eclk, ereset, N0957_port_0,N0957_port_1, N0957_v);
  spice_node_1 n_S00765(eclk, ereset, S00765_port_0, S00765_v);
  spice_node_3 n_N0552(eclk, ereset, N0552_port_2,N0552_port_0,N0552_port_1, N0552_v);
  spice_node_3 n_N0819(eclk, ereset, N0819_port_2,N0819_port_0,N0819_port_1, N0819_v);
  spice_node_6 n_DAA(eclk, ereset, DAA_port_2,DAA_port_3,DAA_port_0,DAA_port_1,DAA_port_4,DAA_port_5, DAA_v);
  spice_node_6 n_DAC(eclk, ereset, DAC_port_2,DAC_port_3,DAC_port_0,DAC_port_1,DAC_port_4,DAC_port_5, DAC_v);
  spice_node_2 n__SRC(eclk, ereset, _SRC_port_0,_SRC_port_1, _SRC_v);
  spice_node_2 n_N0529(eclk, ereset, N0529_port_8,N0529_port_9, N0529_v);
  spice_node_2 n_N0815(eclk, ereset, N0815_port_0,N0815_port_1, N0815_v);
  spice_node_3 n_N0555(eclk, ereset, N0555_port_2,N0555_port_0,N0555_port_1, N0555_v);
  spice_node_2 n_N0816(eclk, ereset, N0816_port_0,N0816_port_1, N0816_v);
  spice_node_2 n___FIN_X12_(eclk, ereset, __FIN_X12__port_2,__FIN_X12__port_3, __FIN_X12__v);
  spice_node_4 n_JUN_JMS(eclk, ereset, JUN_JMS_port_8,JUN_JMS_port_7,JUN_JMS_port_4,JUN_JMS_port_5, JUN_JMS_v);
  spice_node_2 n_N0810(eclk, ereset, N0810_port_0,N0810_port_1, N0810_v);
  spice_node_1 n_S00835(eclk, ereset, S00835_port_0, S00835_v);
  spice_node_2 n_N0812(eclk, ereset, N0812_port_0,N0812_port_1, N0812_v);
  spice_node_3 n_N0554(eclk, ereset, N0554_port_2,N0554_port_0,N0554_port_1, N0554_v);
  spice_node_2 n_N0813(eclk, ereset, N0813_port_0,N0813_port_1, N0813_v);
  spice_node_1 n_PC0_11(eclk, ereset, PC0_11_port_1, PC0_11_v);
  spice_node_1 n_PC0_10(eclk, ereset, PC0_10_port_0, PC0_10_v);
  spice_node_3 n_N0557(eclk, ereset, N0557_port_2,N0557_port_0,N0557_port_1, N0557_v);

endmodule

module spice_node_0(input eclk,ereset, output signed [`W-1:0] v);
  assign v = 0;
endmodule

module spice_node_1(input eclk,ereset, input signed [`W-1:0] i0, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_2(input eclk,ereset, input signed [`W-1:0] i0,i1, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_3(input eclk,ereset, input signed [`W-1:0] i0,i1,i2, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_4(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_5(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_6(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_7(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_8(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6,i7, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6+i7;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_9(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6,i7,i8, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6+i7+i8;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_10(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6+i7+i8+i9;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_11(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6+i7+i8+i9+i10;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_14(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6+i7+i8+i9+i10+i11+i12+i13;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_16(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6+i7+i8+i9+i10+i11+i12+i13+i14+i15;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_18(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12,i13,i14,i15,i16,i17, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6+i7+i8+i9+i10+i11+i12+i13+i14+i15+i16+i17;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

