`include "common.h"

module chip_6502(
  input eclk, ereset,
  output ab0,
  output ab1,
  output ab2,
  output ab3,
  output ab4,
  output ab5,
  output ab6,
  output ab7,
  output ab8,
  output ab9,
  output ab10,
  output ab11,
  output ab12,
  output ab13,
  output ab14,
  output ab15,
  input db0_i,
  output db0_o,
  output db0_t,
  input db1_i,
  output db1_o,
  output db1_t,
  input db2_i,
  output db2_o,
  output db2_t,
  input db3_i,
  output db3_o,
  output db3_t,
  input db4_i,
  output db4_o,
  output db4_t,
  input db5_i,
  output db5_o,
  output db5_t,
  input db6_i,
  output db6_o,
  output db6_t,
  input db7_i,
  output db7_o,
  output db7_t,
  input res,
  output rw,
  output sync,
  input so,
  input clk0,
  output clk1out,
  output clk2out,
  input rdy,
  input nmi,
  input irq
);

  function v;   // convert an analog node value to 2-level
  input [`W-1:0] x;
  begin
    v = ~x[`W-1];
  end
  endfunction

  function [`W-1:0] a;   // convert a 2-level node value to analog
  input x;
  begin
    a = x ? `HI2 : `LO2;
  end
  endfunction

  wire signed [`W-1:0] n_1387_port_2, n_1387_port_3, n_1387_port_0, n_1387_port_1, n_1387_v;
  wire signed [`W-1:0] irq_port_2, irq_v;
  wire signed [`W-1:0] so_port_2, so_port_3, so_v;
  wire signed [`W-1:0] n_304_port_2, n_304_port_3, n_304_port_0, n_304_port_1, n_304_port_4, n_304_v;
  wire signed [`W-1:0] n_330_port_7, n_330_port_4, n_330_v;
  wire signed [`W-1:0] rdy_port_2, rdy_port_3, rdy_v;
  wire signed [`W-1:0] db1_port_1, db1_port_4, db1_port_5, db1_v;
  wire signed [`W-1:0] db0_port_1, db0_port_4, db0_port_5, db0_v;
  wire signed [`W-1:0] db3_port_2, db3_port_3, db3_port_5, db3_v;
  wire signed [`W-1:0] db2_port_2, db2_port_3, db2_port_5, db2_v;
  wire signed [`W-1:0] db5_port_0, db5_port_4, db5_port_5, db5_v;
  wire signed [`W-1:0] db4_port_3, db4_port_0, db4_port_5, db4_v;
  wire signed [`W-1:0] db7_port_3, db7_port_1, db7_port_5, db7_v;
  wire signed [`W-1:0] db6_port_0, db6_port_4, db6_port_5, db6_v;
  wire signed [`W-1:0] n_1661_port_2, n_1661_port_3, n_1661_port_0, n_1661_port_1, n_1661_v;
  wire signed [`W-1:0] idb1_port_8, idb1_port_9, idb1_port_3, idb1_port_0, idb1_port_4, idb1_port_5, idb1_port_10, idb1_v;
  wire signed [`W-1:0] idb0_port_8, idb0_port_2, idb0_port_1, idb0_port_6, idb0_port_7, idb0_port_5, idb0_port_10, idb0_v;
  wire signed [`W-1:0] idb3_port_9, idb3_port_3, idb3_port_0, idb3_port_1, idb3_port_6, idb3_port_5, idb3_port_10, idb3_v;
  wire signed [`W-1:0] idb2_port_3, idb2_port_0, idb2_port_1, idb2_port_6, idb2_port_4, idb2_port_5, idb2_port_10, idb2_v;
  wire signed [`W-1:0] idb5_port_9, idb5_port_2, idb5_port_6, idb5_port_7, idb5_port_4, idb5_port_5, idb5_v;
  wire signed [`W-1:0] idb4_port_9, idb4_port_0, idb4_port_6, idb4_port_7, idb4_port_4, idb4_port_5, idb4_port_10, idb4_v;
  wire signed [`W-1:0] idb7_port_9, idb7_port_2, idb7_port_3, idb7_port_0, idb7_port_7, idb7_port_4, idb7_port_10, idb7_v;
  wire signed [`W-1:0] idb6_port_9, idb6_port_3, idb6_port_0, idb6_port_6, idb6_port_7, idb6_port_5, idb6_port_11, idb6_v;
  wire signed [`W-1:0] n_719_port_2, n_719_port_3, n_719_port_0, n_719_port_1, n_719_v;
  wire signed [`W-1:0] nmi_port_2, nmi_v;
  wire signed [`W-1:0] n_633_port_0, n_633_v;
  wire signed [`W-1:0] n_866_v;
  wire signed [`W-1:0] n_806_v;
  wire signed [`W-1:0] n_807_port_3, n_807_port_5, n_807_v;
  wire signed [`W-1:0] n_87_port_2, n_87_port_3, n_87_port_0, n_87_port_1, n_87_v;
  wire signed [`W-1:0] sb2_port_8, sb2_port_9, sb2_port_3, sb2_port_1, sb2_port_7, sb2_port_10, sb2_port_11, sb2_port_12, sb2_v;
  wire signed [`W-1:0] sb3_port_9, sb3_port_3, sb3_port_1, sb3_port_7, sb3_port_4, sb3_port_5, sb3_port_10, sb3_port_11, sb3_v;
  wire signed [`W-1:0] sb0_port_9, sb0_port_2, sb0_port_1, sb0_port_6, sb0_port_4, sb0_port_10, sb0_port_11, sb0_port_12, sb0_v;
  wire signed [`W-1:0] sb1_port_8, sb1_port_9, sb1_port_2, sb1_port_6, sb1_port_7, sb1_port_10, sb1_port_11, sb1_port_12, sb1_v;
  wire signed [`W-1:0] sb6_port_8, sb6_port_9, sb6_port_2, sb6_port_6, sb6_port_4, sb6_port_10, sb6_port_11, sb6_port_12, sb6_v;
  wire signed [`W-1:0] sb7_port_8, sb7_port_9, sb7_port_3, sb7_port_0, sb7_port_1, sb7_port_6, sb7_port_7, sb7_port_5, sb7_v;
  wire signed [`W-1:0] sb4_port_8, sb4_port_9, sb4_port_3, sb4_port_0, sb4_port_5, sb4_port_10, sb4_port_11, sb4_port_12, sb4_v;
  wire signed [`W-1:0] sb5_port_8, sb5_port_2, sb5_port_3, sb5_port_6, sb5_port_7, sb5_port_10, sb5_port_11, sb5_port_12, sb5_v;
  wire signed [`W-1:0] res_port_2, res_v;
  wire signed [`W-1:0] adl7_port_2, adl7_port_3, adl7_port_0, adl7_port_7, adl7_port_5, adl7_v;
  wire signed [`W-1:0] adl6_port_2, adl6_port_3, adl6_port_1, adl6_port_4, adl6_port_5, adl6_v;
  wire signed [`W-1:0] adl5_port_2, adl5_port_3, adl5_port_0, adl5_port_1, adl5_port_4, adl5_v;
  wire signed [`W-1:0] adl4_port_3, adl4_port_0, adl4_port_1, adl4_port_4, adl4_port_5, adl4_v;
  wire signed [`W-1:0] adl3_port_2, adl3_port_3, adl3_port_0, adl3_port_1, adl3_port_4, adl3_v;
  wire signed [`W-1:0] adl2_port_2, adl2_port_3, adl2_port_0, adl2_port_6, adl2_port_4, adl2_port_5, adl2_v;
  wire signed [`W-1:0] adl1_port_2, adl1_port_3, adl1_port_0, adl1_port_1, adl1_port_4, adl1_port_5, adl1_v;
  wire signed [`W-1:0] adl0_port_3, adl0_port_0, adl0_port_6, adl0_port_7, adl0_port_4, adl0_port_5, adl0_v;
  wire signed [`W-1:0] n_1014_port_2, n_1014_port_3, n_1014_port_0, n_1014_port_1, n_1014_v;
  wire signed [`W-1:0] n_1424_port_2, n_1424_port_3, n_1424_port_0, n_1424_port_1, n_1424_v;
  wire signed [`W-1:0] notaluoutmux0_port_2, notaluoutmux0_port_3, notaluoutmux0_port_0, notaluoutmux0_port_1, notaluoutmux0_port_5, notaluoutmux0_v;
  wire signed [`W-1:0] notaluoutmux1_port_2, notaluoutmux1_port_0, notaluoutmux1_port_1, notaluoutmux1_port_4, notaluoutmux1_port_5, notaluoutmux1_v;
  wire signed [`W-1:0] n_277_port_2, n_277_port_3, n_277_port_1, n_277_port_4, n_277_port_5, n_277_v;
  wire signed [`W-1:0] n_1095_port_2, n_1095_port_3, n_1095_port_0, n_1095_port_1, n_1095_v;
  wire signed [`W-1:0] adh3_port_3, adh3_port_0, adh3_port_6, adh3_port_4, adh3_port_5, adh3_v;
  wire signed [`W-1:0] adh2_port_3, adh2_port_0, adh2_port_6, adh2_port_4, adh2_port_5, adh2_v;
  wire signed [`W-1:0] adh1_port_2, adh1_port_0, adh1_port_1, adh1_port_6, adh1_port_4, adh1_v;
  wire signed [`W-1:0] adh0_port_2, adh0_port_3, adh0_port_0, adh0_port_1, adh0_port_6, adh0_v;
  wire signed [`W-1:0] adh7_port_2, adh7_port_3, adh7_port_0, adh7_port_4, adh7_port_5, adh7_v;
  wire signed [`W-1:0] adh6_port_3, adh6_port_0, adh6_port_6, adh6_port_4, adh6_port_5, adh6_v;
  wire signed [`W-1:0] adh5_port_2, adh5_port_3, adh5_port_0, adh5_port_4, adh5_port_5, adh5_v;
  wire signed [`W-1:0] adh4_port_2, adh4_port_0, adh4_port_6, adh4_port_4, adh4_port_5, adh4_v;
  wire signed [`W-1:0] NMIP_port_7, NMIP_port_4, NMIP_v;
  wire signed [`W-1:0] n_1071_port_2, n_1071_port_3, n_1071_port_0, n_1071_port_4, n_1071_port_5, n_1071_v;
  wire signed [`W-1:0] n_1147_port_2, n_1147_port_3, n_1147_port_0, n_1147_port_1, n_1147_v;
  wire signed [`W-1:0] n_722_port_2, n_722_port_0, n_722_port_1, n_722_port_4, n_722_port_5, n_722_v;
  wire signed [`W-1:0] n_1059_port_0, n_1059_v;
  wire signed [`W-1:0] n_740_port_2, n_740_port_3, n_740_port_0, n_740_port_1, n_740_port_4, n_740_v;
  wire signed [`W-1:0] n_975_port_3, n_975_port_6, n_975_v;
  wire signed [`W-1:0] clk0_port_3, clk0_v;
  wire signed [`W-1:0] _ABH3_port_3, _ABH3_v;
  wire signed [`W-1:0] _ABH1_port_3, _ABH1_v;
  wire signed [`W-1:0] _ABH0_port_3, _ABH0_v;
  wire signed [`W-1:0] _ABH7_port_3, _ABH7_v;
  wire signed [`W-1:0] _ABH6_port_3, _ABH6_v;
  wire signed [`W-1:0] _ABH5_port_3, _ABH5_v;
  wire signed [`W-1:0] n_854_port_6, n_854_port_4, n_854_v;
  wire signed [`W-1:0] n_297_port_3, n_297_port_5, n_297_v;
  wire signed [`W-1:0] n_296_port_3, n_296_port_0, n_296_port_1, n_296_port_4, n_296_port_5, n_296_v;

  wire pipedpc28_v;
  wire dor5_v;
  wire dor4_v;
  wire dor7_v;
  wire dor6_v;
  wire dor1_v;
  wire dor0_v;
  wire dor3_v;
  wire dor2_v;
  wire _DBZ_v;
  wire _DBE_v;
  wire n_1714_v;
  wire n_1715_v;
  wire n_1716_v;
  wire n_1717_v;
  wire n_1247_v;
  wire n_1244_v;
  wire n_1245_v;
  wire n_1718_v;
  wire n_1719_v;
  wire _ABL7_v;
  wire _ABL6_v;
  wire _ABL5_v;
  wire _ABL3_v;
  wire _ABL2_v;
  wire _ABL1_v;
  wire _ABL0_v;
  wire dpc5_SADL_v;
  wire n_604_v;
  wire n_600_v;
  wire n_602_v;
  wire n_603_v;
  wire n_608_v;
  wire n_609_v;
  wire pd6_clearIR_v;
  wire n_460_v;
  wire n_462_v;
  wire n_465_v;
  wire n_466_v;
  wire n_467_v;
  wire n_468_v;
  wire n_469_v;
  wire op_T4_brk_v;
  wire n_1162_v;
  wire n_1161_v;
  wire rw_v;
  wire x_op_T3_plp_pla_v;
  wire idl7_v;
  wire idl6_v;
  wire idl5_v;
  wire idl4_v;
  wire idl3_v;
  wire idl2_v;
  wire idl1_v;
  wire idl0_v;
  wire n_1529_v;
  wire n_1528_v;
  wire n_1523_v;
  wire n_1521_v;
  wire n_1527_v;
  wire n_1526_v;
  wire n_733_v;
  wire dpc20_ADDSB06_v;
  wire n_1389_v;
  wire n_1386_v;
  wire n_1383_v;
  wire n_1380_v;
  wire x6_v;
  wire n_819_v;
  wire n_818_v;
  wire n_811_v;
  wire n_810_v;
  wire n_813_v;
  wire n_812_v;
  wire n_815_v;
  wire ir0_v;
  wire ir1_v;
  wire ir2_v;
  wire ir3_v;
  wire ir4_v;
  wire ir5_v;
  wire ir6_v;
  wire ir7_v;
  wire n_599_v;
  wire n_1267_v;
  wire n_1260_v;
  wire op_T__inx_v;
  wire n_9_v;
  wire n_5_v;
  wire n_6_v;
  wire n_7_v;
  wire n_3_v;
  wire aluanandb0_v;
  wire aluanandb1_v;
  wire n_1240_v;
  wire n_1711_v;
  wire n_1712_v;
  wire op_T0_php_pha_v;
  wire dasb6_v;
  wire dasb5_v;
  wire dasb3_v;
  wire dasb2_v;
  wire dasb1_v;
  wire n_662_v;
  wire n_663_v;
  wire n_666_v;
  wire n_664_v;
  wire alu4_v;
  wire alu5_v;
  wire alu6_v;
  wire alu7_v;
  wire alu0_v;
  wire alu1_v;
  wire alu2_v;
  wire alu3_v;
  wire _ABL4_v;
  wire n_488_v;
  wire n_484_v;
  wire n_485_v;
  wire n_480_v;
  wire n_481_v;
  wire PD_xxx010x1_v;
  wire op_shift_v;
  wire op_xy_v;
  wire op_T0_cld_sed_v;
  wire n_327_v;
  wire n_326_v;
  wire _AxB_0__C0in_v;
  wire n_321_v;
  wire n_320_v;
  wire n_1105_v;
  wire n_1107_v;
  wire n_1106_v;
  wire n_1101_v;
  wire n_1100_v;
  wire n_1109_v;
  wire pd4_clearIR_v;
  wire op_ror_v;
  wire dpc6_SBS_v;
  wire n_345_v;
  wire n_347_v;
  wire n_340_v;
  wire n_831_v;
  wire n_830_v;
  wire n_839_v;
  wire n_838_v;
  wire op_T0_ldy_mem_v;
  wire D1x1_v;
  wire s3_v;
  wire s2_v;
  wire s1_v;
  wire s0_v;
  wire s7_v;
  wire s6_v;
  wire s5_v;
  wire s4_v;
  wire dpc15_ANDS_v;
  wire n_1585_v;
  wire n_1586_v;
  wire _TWOCYCLE_v;
  wire dpc27_SBADH_v;
  wire pd3_clearIR_v;
  wire n_1450_v;
  wire n_649_v;
  wire n_138_v;
  wire n_139_v;
  wire n_641_v;
  wire n_642_v;
  wire n_643_v;
  wire n_132_v;
  wire n_645_v;
  wire n_646_v;
  wire n_647_v;
  wire n_1632_v;
  wire n_1635_v;
  wire _AxB_6__C56_v;
  wire pd0_clearIR_v;
  wire op_T0_shift_a_v;
  wire __AxB7__C67_v;
  wire n_1439_v;
  wire _VEC_v;
  wire n_1129_v;
  wire n_1126_v;
  wire n_1124_v;
  wire n_1121_v;
  wire n_1120_v;
  wire n_587_v;
  wire n_586_v;
  wire n_583_v;
  wire n_582_v;
  wire n_588_v;
  wire op_rmw_v;
  wire n_360_v;
  wire n_366_v;
  wire n_368_v;
  wire op_jmp_v;
  wire C12_v;
  wire n_1433_v;
  wire op_shift_right_v;
  wire op_EORS_v;
  wire x_op_T__adc_sbc_v;
  wire n_1631_v;
  wire notir0_v;
  wire notir1_v;
  wire notir2_v;
  wire notir3_v;
  wire notir4_v;
  wire notir5_v;
  wire notir6_v;
  wire notir7_v;
  wire n_94_v;
  wire n_95_v;
  wire n_93_v;
  wire n_90_v;
  wire n_91_v;
  wire op_lsr_ror_dec_inc_v;
  wire n_110_v;
  wire n_111_v;
  wire n_118_v;
  wire n_119_v;
  wire cp1_v;
  wire a3_v;
  wire a6_v;
  wire n_696_v;
  wire n_698_v;
  wire n_1199_v;
  wire n_930_v;
  wire DA_AxB2_v;
  wire n_1479_v;
  wire pipeVectorA2_v;
  wire sync_v;
  wire n_745_v;
  wire n_1499_v;
  wire n_1325_v;
  wire n_1496_v;
  wire n_1495_v;
  wire n_1492_v;
  wire n_1323_v;
  wire n_1141_v;
  wire n_568_v;
  wire n_565_v;
  wire n_564_v;
  wire n_567_v;
  wire n_566_v;
  wire n_562_v;
  wire __AxBxC_6_v;
  wire __AxBxC_7_v;
  wire __AxBxC_4_v;
  wire __AxBxC_5_v;
  wire __AxBxC_2_v;
  wire __AxBxC_3_v;
  wire __AxBxC_0_v;
  wire __AxBxC_1_v;
  wire n_300_v;
  wire n_307_v;
  wire n_306_v;
  wire aluaorb0_v;
  wire x_op_T0_tya_v;
  wire x_op_T4_ind_y_v;
  wire pclp0_v;
  wire pclp1_v;
  wire pclp2_v;
  wire pclp3_v;
  wire pclp4_v;
  wire pclp5_v;
  wire pclp6_v;
  wire pclp7_v;
  wire op_T3_branch_v;
  wire ab12_v;
  wire ab13_v;
  wire ab10_v;
  wire ab11_v;
  wire n_79_v;
  wire ab14_v;
  wire ab15_v;
  wire n_75_v;
  wire n_70_v;
  wire n_71_v;
  wire n_72_v;
  wire n_1252_v;
  wire n_1705_v;
  wire n_1256_v;
  wire op_T0_tya_v;
  wire n_172_v;
  wire n_176_v;
  wire n_177_v;
  wire n_796_v;
  wire n_797_v;
  wire n_794_v;
  wire n_795_v;
  wire n_790_v;
  wire n_798_v;
  wire n_799_v;
  wire pd7_v;
  wire pd6_v;
  wire pd5_v;
  wire pd4_v;
  wire pd3_v;
  wire pd2_v;
  wire pd1_v;
  wire pd0_v;
  wire n_1305_v;
  wire n_1304_v;
  wire n_1303_v;
  wire n_1301_v;
  wire n_1300_v;
  wire n_1309_v;
  wire n_332_v;
  wire n_1166_v;
  wire n_1169_v;
  wire n_339_v;
  wire PD_1xx000x0_v;
  wire n_548_v;
  wire op_T2_brk_v;
  wire n_543_v;
  wire n_541_v;
  wire n_544_v;
  wire C56_v;
  wire n_890_v;
  wire n_323_v;
  wire n_322_v;
  wire n_897_v;
  wire n_896_v;
  wire n_329_v;
  wire pipeUNK31_v;
  wire xx_op_T5_jsr_v;
  wire PD_xxxx10x0_v;
  wire n_1028_v;
  wire dpc24_ACSB_v;
  wire n_50_v;
  wire n_55_v;
  wire n_152_v;
  wire n_154_v;
  wire n_1347_v;
  wire op_ORS_v;
  wire n_1346_v;
  wire _AxB_2__C12_v;
  wire n_1360_v;
  wire n_1364_v;
  wire n_1369_v;
  wire n_1368_v;
  wire clearIR_v;
  wire op_T__cpx_cpy_imm_zp_v;
  wire n_1187_v;
  wire n_1181_v;
  wire n_1180_v;
  wire op_T5_mem_ind_idx_v;
  wire n_521_v;
  wire n_520_v;
  wire n_523_v;
  wire n_525_v;
  wire n_526_v;
  wire C78_v;
  wire dpc21_ADDADL_v;
  wire n_1592_v;
  wire n_31_v;
  wire n_34_v;
  wire n_35_v;
  wire n_36_v;
  wire n_37_v;
  wire pchp4_v;
  wire pchp5_v;
  wire pchp6_v;
  wire pchp7_v;
  wire pchp0_v;
  wire pchp1_v;
  wire pchp2_v;
  wire pchp3_v;
  wire clk1out_v;
  wire _WR_v;
  wire n_1647_v;
  wire n_1642_v;
  wire n_1643_v;
  wire n_1640_v;
  wire n_1641_v;
  wire n_1649_v;
  wire _op_branch_bit6_v;
  wire _op_branch_bit7_v;
  wire n_1184_v;
  wire op_rol_ror_v;
  wire n_1491_v;
  wire n_201_v;
  wire n_206_v;
  wire clock1_v;
  wire clock2_v;
  wire n_1434_v;
  wire n_1341_v;
  wire n_1344_v;
  wire op_asl_rol_v;
  wire short_circuit_idx_add_v;
  wire n_509_v;
  wire n_507_v;
  wire n_506_v;
  wire n_504_v;
  wire n_503_v;
  wire n_501_v;
  wire x_op_T0_bit_v;
  wire n_18_v;
  wire n_16_v;
  wire n_17_v;
  wire n_14_v;
  wire n_15_v;
  wire n_10_v;
  wire n_11_v;
  wire n_1084_v;
  wire n_1085_v;
  wire n_1087_v;
  wire n_1081_v;
  wire n_1082_v;
  wire n_1083_v;
  wire n_1089_v;
  wire n_1269_v;
  wire dpc35_PCHC_v;
  wire n_1265_v;
  wire n_1662_v;
  wire n_1262_v;
  wire n_1668_v;
  wire op_T2_abs_y_v;
  wire n_267_v;
  wire n_264_v;
  wire n_265_v;
  wire n_262_v;
  wire n_260_v;
  wire n_261_v;
  wire n_269_v;
  wire dpc32_PCHADH_v;
  wire n_8_v;
  wire op_T3_mem_abs_v;
  wire op_T2_ADL_ADD_v;
  wire n_1417_v;
  wire n_1416_v;
  wire n_1413_v;
  wire n_1412_v;
  wire n_1411_v;
  wire n_381_v;
  wire n_383_v;
  wire n_385_v;
  wire n_384_v;
  wire n_386_v;
  wire n_389_v;
  wire n_388_v;
  wire op_T__shift_a_v;
  wire n_927_v;
  wire n_920_v;
  wire n_923_v;
  wire n_928_v;
  wire n_1039_v;
  wire alub2_v;
  wire pch7_v;
  wire pch6_v;
  wire pch5_v;
  wire pch4_v;
  wire pch3_v;
  wire pch2_v;
  wire pch1_v;
  wire pch0_v;
  wire op_T3_mem_zp_idx_v;
  wire notalucin_v;
  wire dpc13_ORS_v;
  wire n_1069_v;
  wire n_1067_v;
  wire n_1065_v;
  wire n_1063_v;
  wire n_1061_v;
  wire op_T0_tay_v;
  wire op_T0_tax_v;
  wire n_1608_v;
  wire n_1609_v;
  wire n_1606_v;
  wire n_1605_v;
  wire op_T0_brk_rti_v;
  wire n_249_v;
  wire n_718_v;
  wire n_717_v;
  wire n_715_v;
  wire n_241_v;
  wire n_242_v;
  wire n_243_v;
  wire dasb7_v;
  wire notidl0_v;
  wire op_T5_rti_rts_v;
  wire pipeT3out_v;
  wire n_669_v;
  wire _C23_v;
  wire nnT2BR_v;
  wire n_1472_v;
  wire n_1474_v;
  wire n_1477_v;
  wire op_T4_ind_y_v;
  wire n_1295_v;
  wire n_1296_v;
  wire n_1291_v;
  wire n_1290_v;
  wire n_1293_v;
  wire dpc7_SS_v;
  wire op_T__iny_dey_v;
  wire n_902_v;
  wire n_906_v;
  wire n_905_v;
  wire n_1356_v;
  wire n_1423_v;
  wire pipeUNK18_v;
  wire pipeUNK16_v;
  wire pipeUNK17_v;
  wire pipeUNK14_v;
  wire pipeUNK15_v;
  wire pipeUNK12_v;
  wire pipeUNK13_v;
  wire pipeUNK11_v;
  wire n_38_v;
  wire n_1599_v;
  wire n_1041_v;
  wire n_1043_v;
  wire n_1596_v;
  wire n_1045_v;
  wire n_1046_v;
  wire n_1595_v;
  wire n_1624_v;
  wire n_1625_v;
  wire n_1620_v;
  wire n_1621_v;
  wire n_1629_v;
  wire n_228_v;
  wire n_223_v;
  wire n_220_v;
  wire n_221_v;
  wire n_226_v;
  wire n_227_v;
  wire n_224_v;
  wire n_225_v;
  wire op_T4_abs_idx_v;
  wire op_implied_v;
  wire n_735_v;
  wire n_730_v;
  wire n_732_v;
  wire dpc22__DSA_v;
  wire n_739_v;
  wire x2_v;
  wire x3_v;
  wire x0_v;
  wire x1_v;
  wire op_T__dex_v;
  wire x7_v;
  wire x4_v;
  wire x5_v;
  wire n_415_v;
  wire _C01_v;
  wire op_T0_sbc_v;
  wire n_410_v;
  wire n_1458_v;
  wire n_1452_v;
  wire n_1457_v;
  wire n_1455_v;
  wire DA_AB2_v;
  wire n_692_v;
  wire n_695_v;
  wire n_694_v;
  wire n_969_v;
  wire n_968_v;
  wire n_961_v;
  wire n_963_v;
  wire n_962_v;
  wire n_964_v;
  wire n_966_v;
  wire irline3_v;
  wire pcl3_v;
  wire pcl2_v;
  wire pcl1_v;
  wire pcl0_v;
  wire pcl7_v;
  wire pcl6_v;
  wire pcl5_v;
  wire pcl4_v;
  wire dpc0_YSB_v;
  wire pipeUNK34_v;
  wire pipeUNK35_v;
  wire pipeUNK36_v;
  wire pipeUNK37_v;
  wire pipeUNK30_v;
  wire pipeUNK32_v;
  wire pipeUNK33_v;
  wire pipeUNK39_v;
  wire n_1020_v;
  wire n_1026_v;
  wire n_1027_v;
  wire n_1024_v;
  wire n_1025_v;
  wire alua6_v;
  wire alua7_v;
  wire alua4_v;
  wire alua5_v;
  wire alua2_v;
  wire alua3_v;
  wire alua0_v;
  wire alua1_v;
  wire n_1271_v;
  wire op_T2_branch_v;
  wire dpc41_DL_ADL_v;
  wire n_200_v;
  wire n_753_v;
  wire n_756_v;
  wire n_757_v;
  wire n_754_v;
  wire n_207_v;
  wire n_208_v;
  wire n_209_v;
  wire n_759_v;
  wire _C67_v;
  wire dpc37_PCLDB_v;
  wire __AxB3__C23_v;
  wire pipephi2Reset0_v;
  wire pd5_clearIR_v;
  wire dpc12_0ADD_v;
  wire dpc4_SSB_v;
  wire n_134_v;
  wire n_947_v;
  wire n_946_v;
  wire n_417_v;
  wire n_944_v;
  wire op_T0_cpy_iny_v;
  wire n_419_v;
  wire y1_v;
  wire y0_v;
  wire y3_v;
  wire y2_v;
  wire y5_v;
  wire y4_v;
  wire y7_v;
  wire y6_v;
  wire n_1007_v;
  wire n_1002_v;
  wire abh5_v;
  wire abh4_v;
  wire abh7_v;
  wire abh6_v;
  wire abh1_v;
  wire abh0_v;
  wire abh3_v;
  wire abh2_v;
  wire n_1552_v;
  wire alucin_v;
  wire x_op_push_pull_v;
  wire dpc11_SBADD_v;
  wire dpc10_ADLADD_v;
  wire n_779_v;
  wire n_770_v;
  wire n_771_v;
  wire n_772_v;
  wire n_773_v;
  wire n_774_v;
  wire n_837_v;
  wire op_T0_bit_v;
  wire n_344_v;
  wire n_834_v;
  wire dpc29_0ADH17_v;
  wire dpc26_ACDB_v;
  wire _C45_v;
  wire VEC0_v;
  wire VEC1_v;
  wire op_T4_rts_v;
  wire n_430_v;
  wire n_436_v;
  wire op_T4_rti_v;
  wire op_SRS_v;
  wire n_1343_v;
  wire n_1345_v;
  wire n_1578_v;
  wire n_1579_v;
  wire n_1573_v;
  wire n_1574_v;
  wire DC78_v;
  wire op_sta_cmp_v;
  wire op_SUMS_v;
  wire n_1688_v;
  wire pipeT2out_v;
  wire n_404_v;
  wire n_954_v;
  wire n_400_v;
  wire op_T4_brk_jsr_v;
  wire n_1219_v;
  wire n_1215_v;
  wire n_1214_v;
  wire n_1211_v;
  wire n_1213_v;
  wire n_1655_v;
  wire pd2_clearIR_v;
  wire n_1654_v;
  wire n_1657_v;
  wire n_1650_v;
  wire n_182_v;
  wire n_180_v;
  wire n_184_v;
  wire n_635_v;
  wire n_634_v;
  wire n_637_v;
  wire n_636_v;
  wire n_631_v;
  wire n_630_v;
  wire n_632_v;
  wire n_459_v;
  wire n_458_v;
  wire n_988_v;
  wire n_983_v;
  wire n_982_v;
  wire n_981_v;
  wire n_987_v;
  wire n_986_v;
  wire n_457_v;
  wire op_T0_lda_v;
  wire abl1_v;
  wire abl0_v;
  wire abl4_v;
  wire pipe_WR_phi2_v;
  wire op_T3_plp_pla_v;
  wire n_1517_v;
  wire n_1518_v;
  wire n_1519_v;
  wire DC78_phi2_v;
  wire n_279_v;
  wire n_846_v;
  wire n_847_v;
  wire n_844_v;
  wire n_845_v;
  wire n_842_v;
  wire op_T3_jmp_v;
  wire n_849_v;
  wire __AxB5__C45_v;
  wire dpc16_EORS_v;
  wire n_1231_v;
  wire n_1230_v;
  wire n_1238_v;
  wire n_1722_v;
  wire op_branch_done_v;
  wire aluvout_v;
  wire n_618_v;
  wire n_613_v;
  wire n_612_v;
  wire n_611_v;
  wire n_610_v;
  wire n_617_v;
  wire n_616_v;
  wire n_1137_v;
  wire n_620_v;
  wire n_884_v;
  wire Pout0_v;
  wire n_1545_v;
  wire n_1010_v;
  wire n_1017_v;
  wire n_1542_v;
  wire dpc19_ADDSB7_v;
  wire n_477_v;
  wire n_476_v;
  wire n_475_v;
  wire n_474_v;
  wire n_473_v;
  wire n_472_v;
  wire n_471_v;
  wire n_470_v;
  wire n_479_v;
  wire n_478_v;
  wire brk_done_v;
  wire p2_v;
  wire p3_v;
  wire op_T0_txa_v;
  wire p0_v;
  wire p6_v;
  wire p7_v;
  wire DC34_v;
  wire op_T2_stack_v;
  wire n_1534_v;
  wire n_1531_v;
  wire n_1533_v;
  wire n_1391_v;
  wire n_1392_v;
  wire n_1395_v;
  wire n_1398_v;
  wire n_1399_v;
  wire n_288_v;
  wire n_280_v;
  wire n_282_v;
  wire n_284_v;
  wire n_135_v;
  wire n_644_v;
  wire n_133_v;
  wire n_130_v;
  wire n_869_v;
  wire n_865_v;
  wire n_867_v;
  wire n_861_v;
  wire n_862_v;
  wire pipeT4out_v;
  wire n_350_v;
  wire dpc17_SUMS_v;
  wire pipeT_SYNC_v;
  wire _op_branch_done_v;
  wire op_T0_acc_v;
  wire BRtaken_v;
  wire n_1251_v;
  wire n_1253_v;
  wire n_1257_v;
  wire n_1258_v;
  wire n_1709_v;
  wire n_1708_v;
  wire dpc3_SBX_v;
  wire op_T2_php_v;
  wire op_T2_pha_v;
  wire dpc31_PCHPCH_v;
  wire n_671_v;
  wire n_670_v;
  wire n_673_v;
  wire n_675_v;
  wire n_674_v;
  wire n_676_v;
  wire n_678_v;
  wire Pout1_v;
  wire Pout3_v;
  wire Pout2_v;
  wire n_499_v;
  wire n_494_v;
  wire n_496_v;
  wire n_491_v;
  wire n_490_v;
  wire pd7_clearIR_v;
  wire n_1401_v;
  wire n_1404_v;
  wire op_T4_jmp_v;
  wire n_19_v;
  wire n_1117_v;
  wire n_1115_v;
  wire n_1113_v;
  wire n_1110_v;
  wire n_1111_v;
  wire n_803_v;
  wire n_800_v;
  wire n_805_v;
  wire n_432_v;
  wire n_1272_v;
  wire n_1277_v;
  wire n_1276_v;
  wire n_1275_v;
  wire n_1274_v;
  wire n_1660_v;
  wire op_inc_nop_v;
  wire n_128_v;
  wire n_659_v;
  wire n_658_v;
  wire n_127_v;
  wire n_126_v;
  wire n_653_v;
  wire n_652_v;
  wire n_123_v;
  wire n_122_v;
  wire op_T0_shift_right_a_v;
  wire op_T0_adc_sbc_v;
  wire op_push_pull_v;
  wire pipe_VEC_v;
  wire n_266_v;
  wire n_1130_v;
  wire n_1132_v;
  wire n_1133_v;
  wire n_1135_v;
  wire n_1138_v;
  wire op_T2_mem_zp_v;
  wire n_355_v;
  wire n_824_v;
  wire n_826_v;
  wire n_351_v;
  wire dpc9_DBADD_v;
  wire n_358_v;
  wire n_359_v;
  wire dpc33_PCHDB_v;
  wire INTG_v;
  wire n_755_v;
  wire op_T2_ind_v;
  wire op_rti_rts_v;
  wire dpc8_nDBADD_v;
  wire notdor1_v;
  wire notdor0_v;
  wire notdor3_v;
  wire notdor2_v;
  wire notdor5_v;
  wire notdor4_v;
  wire notdor7_v;
  wire notdor6_v;
  wire n_1570_v;
  wire n_109_v;
  wire n_108_v;
  wire n_102_v;
  wire n_101_v;
  wire n_105_v;
  wire n_104_v;
  wire n_1575_v;
  wire dpc39_PCLPCL_v;
  wire ADH_ABH_v;
  wire n_581_v;
  wire Reset0_v;
  wire dpc25_SBDB_v;
  wire n_1541_v;
  wire dpc23_SBAC_v;
  wire n_1484_v;
  wire x_op_jmp_v;
  wire n_1338_v;
  wire n_1339_v;
  wire n_1488_v;
  wire n_1335_v;
  wire n_1333_v;
  wire n_1159_v;
  wire n_1152_v;
  wire n_1157_v;
  wire n_1154_v;
  wire _t2_v;
  wire _t3_v;
  wire n_595_v;
  wire n_597_v;
  wire _t4_v;
  wire _t5_v;
  wire nots3_v;
  wire nots2_v;
  wire nots1_v;
  wire nots0_v;
  wire nots7_v;
  wire nots6_v;
  wire nots5_v;
  wire nots4_v;
  wire n_1682_v;
  wire n_378_v;
  wire n_1683_v;
  wire n_374_v;
  wire n_372_v;
  wire n_373_v;
  wire x_op_T0_txa_v;
  wire C01_v;
  wire op_store_v;
  wire n_1687_v;
  wire ab0_v;
  wire ab1_v;
  wire ab2_v;
  wire ab3_v;
  wire ab4_v;
  wire ab5_v;
  wire ab6_v;
  wire ab7_v;
  wire ab8_v;
  wire ab9_v;
  wire n_80_v;
  wire n_83_v;
  wire n_86_v;
  wire n_88_v;
  wire n_1684_v;
  wire n_161_v;
  wire n_160_v;
  wire n_163_v;
  wire n_169_v;
  wire n_168_v;
  wire n_785_v;
  wire n_781_v;
  wire n_783_v;
  wire n_782_v;
  wire n_789_v;
  wire __AxB_6_v;
  wire __AxB_4_v;
  wire __AxB_2_v;
  wire __AxB_0_v;
  wire n_1318_v;
  wire n_1319_v;
  wire n_1312_v;
  wire n_1315_v;
  wire n_1316_v;
  wire dpc2_XSB_v;
  wire n_1175_v;
  wire n_1177_v;
  wire n_1170_v;
  wire n_1178_v;
  wire n_1179_v;
  wire n_578_v;
  wire n_572_v;
  wire n_570_v;
  wire n_571_v;
  wire n_318_v;
  wire n_319_v;
  wire n_312_v;
  wire n_310_v;
  wire n_311_v;
  wire n_317_v;
  wire PD_n_0xx0xx0x_v;
  wire C23_v;
  wire PD_0xx0xx0x_v;
  wire op_T0_dex_v;
  wire C78_phi2_v;
  wire op_T__ora_and_eor_adc_v;
  wire dpc14_SRS_v;
  wire op_T2_ind_x_v;
  wire op_T2_ind_y_v;
  wire op_plp_pla_v;
  wire op_T0_txs_v;
  wire n_69_v;
  wire n_66_v;
  wire n_62_v;
  wire n_61_v;
  wire n_149_v;
  wire n_147_v;
  wire n_146_v;
  wire n_141_v;
  wire _op_set_C_v;
  wire op_T5_rti_v;
  wire op_T5_ind_y_v;
  wire op_T5_ind_x_v;
  wire op_T3_jsr_v;
  wire op_T5_brk_v;
  wire ADL_ABL_v;
  wire n_1371_v;
  wire n_1376_v;
  wire n_1377_v;
  wire n_1374_v;
  wire n_1375_v;
  wire n_1379_v;
  wire n_1724_v;
  wire n_1194_v;
  wire n_1195_v;
  wire n_1192_v;
  wire n_1190_v;
  wire n_1191_v;
  wire n_708_v;
  wire n_556_v;
  wire n_550_v;
  wire n_551_v;
  wire n_553_v;
  wire n_559_v;
  wire C45_v;
  wire x_op_T3_ind_y_v;
  wire op_T__asl_rol_a_v;
  wire n_882_v;
  wire n_883_v;
  wire n_880_v;
  wire n_334_v;
  wire n_335_v;
  wire n_336_v;
  wire n_885_v;
  wire n_888_v;
  wire n_889_v;
  wire _AxB_4__C34_v;
  wire dpc28_0ADH0_v;
  wire fetch_v;
  wire op_ANDS_v;
  wire n_47_v;
  wire n_46_v;
  wire n_43_v;
  wire n_42_v;
  wire op_T__cpx_cpy_abs_v;
  wire n_1153_v;
  wire n_0_ADL1_v;
  wire n_0_ADL0_v;
  wire n_0_ADL2_v;
  wire op_T3_abs_idx_v;
  wire op_jsr_v;
  wire n_590_v;
  wire dpc40_ADLPCL_v;
  wire n_593_v;
  wire n_929_v;
  wire n_598_v;
  wire n_1255_v;
  wire n_1358_v;
  wire n_1427_v;
  wire n_1357_v;
  wire n_533_v;
  wire n_531_v;
  wire n_538_v;
  wire C67_v;
  wire C1x5Reset_v;
  wire op_T__adc_sbc_v;
  wire op_T0_cmp_v;
  wire pipeBRtaken_v;
  wire n_1218_v;
  wire dpc30_ADHPCH_v;
  wire pipeUNK41_v;
  wire pipeUNK40_v;
  wire pipeUNK42_v;
  wire dpc43_DL_DB_v;
  wire n_23_v;
  wire n_21_v;
  wire n_20_v;
  wire n_27_v;
  wire aluanorb0_v;
  wire n_25_v;
  wire n_24_v;
  wire n_29_v;
  wire n_1693_v;
  wire n_1694_v;
  wire a1_v;
  wire a0_v;
  wire a2_v;
  wire a5_v;
  wire a4_v;
  wire a7_v;
  wire pipephi2Reset0x_v;
  wire n_275_v;
  wire n_270_v;
  wire n_272_v;
  wire n_278_v;
  wire n_1486_v;
  wire n_638_v;
  wire n_1408_v;
  wire n_1409_v;
  wire n_188_v;
  wire n_1400_v;
  wire n_1402_v;
  wire op_T0_ora_v;
  wire n_518_v;
  wire n_519_v;
  wire n_510_v;
  wire n_512_v;
  wire n_513_v;
  wire n_515_v;
  wire n_1463_v;
  wire n_453_v;
  wire n_1467_v;
  wire n_980_v;
  wire n_1464_v;
  wire alucout_v;
  wire op_brk_rti_v;
  wire DBZ_v;
  wire pipeVectorA0_v;
  wire pipeVectorA1_v;
  wire n_1602_v;
  wire pipeT5out_v;
  wire n_1600_v;
  wire n_1093_v;
  wire n_1091_v;
  wire n_1090_v;
  wire n_1097_v;
  wire n_1094_v;
  wire n_1099_v;
  wire n_1679_v;
  wire n_1677_v;
  wire n_1676_v;
  wire n_1675_v;
  wire n_1674_v;
  wire n_1673_v;
  wire op_T5_rts_v;
  wire n_253_v;
  wire n_251_v;
  wire n_709_v;
  wire n_256_v;
  wire n_255_v;
  wire n_254_v;
  wire n_700_v;
  wire n_1462_v;
  wire n_1469_v;
  wire n_714_v;
  wire n_1286_v;
  wire n_1281_v;
  wire n_1289_v;
  wire A_B7_v;
  wire A_B5_v;
  wire A_B3_v;
  wire A_B1_v;
  wire n_392_v;
  wire n_393_v;
  wire n_390_v;
  wire n_396_v;
  wire n_397_v;
  wire n_398_v;
  wire n_1497_v;
  wire n_936_v;
  wire n_937_v;
  wire n_935_v;
  wire n_933_v;
  wire n_931_v;
  wire op_T2_php_pha_v;
  wire ONEBYTE_v;
  wire pipeUNK09_v;
  wire pipeUNK08_v;
  wire pipeUNK05_v;
  wire pipeUNK04_v;
  wire pipeUNK07_v;
  wire pipeUNK06_v;
  wire pipeUNK01_v;
  wire pipeUNK03_v;
  wire pipeUNK02_v;
  wire n_1075_v;
  wire n_1076_v;
  wire n_1070_v;
  wire n_1073_v;
  wire n_1072_v;
  wire n_1149_v;
  wire abl2_v;
  wire abl5_v;
  wire abl6_v;
  wire n_1619_v;
  wire notaluvout_v;
  wire n_1140_v;
  wire n_1614_v;
  wire n_1145_v;
  wire dpc34_PCLC_v;
  wire aluanorb1_v;
  wire H1x1_v;
  wire n_238_v;
  wire n_728_v;
  wire n_723_v;
  wire n_721_v;
  wire n_720_v;
  wire n_726_v;
  wire dpc1_SBY_v;
  wire op_T2_abs_v;
  wire op_T0_plp_v;
  wire op_T0_pla_v;
  wire op_T2_jmp_abs_v;
  wire pipe_T0_v;
  wire _C34_v;
  wire DA_C01_v;
  wire n_1448_v;
  wire n_1449_v;
  wire cclk_v;
  wire n_1446_v;
  wire n_1447_v;
  wire n_1440_v;
  wire n_1441_v;
  wire notRnWprepad_v;
  wire n_1511_v;
  wire n_918_v;
  wire n_919_v;
  wire n_916_v;
  wire n_917_v;
  wire RnWstretched_v;
  wire n_913_v;
  wire op_T0_tay_ldy_not_idx_v;
  wire op_T0_v;
  wire op_T3_v;
  wire op_T2_v;
  wire op_T4_v;
  wire n_1224_v;
  wire op_T3_stack_bit_jmp_v;
  wire op_T5_jsr_v;
  wire op_T2_stack_access_v;
  wire pipeUNK23_v;
  wire pipeUNK22_v;
  wire pipeUNK21_v;
  wire pipeUNK20_v;
  wire pipeUNK27_v;
  wire pipeUNK26_v;
  wire pipeUNK29_v;
  wire pipeUNK28_v;
  wire n_1056_v;
  wire n_1055_v;
  wire n_1054_v;
  wire op_T4_mem_abs_idx_v;
  wire n_1588_v;
  wire n_1581_v;
  wire n_1580_v;
  wire n_1633_v;
  wire n_1639_v;
  wire n_1638_v;
  wire C34_v;
  wire _DA_ADD2_v;
  wire _DA_ADD1_v;
  wire n_743_v;
  wire n_213_v;
  wire n_212_v;
  wire n_747_v;
  wire n_210_v;
  wire n_748_v;
  wire n_218_v;
  wire notRdy0_v;
  wire notalucout_v;
  wire dpc36_IPC_v;
  wire op_T0_cpx_cpy_inx_iny_v;
  wire n_624_v;
  wire op_T2_zp_zp_idx_v;
  wire _C12_v;
  wire clk2out_v;
  wire n_688_v;
  wire n_689_v;
  wire n_680_v;
  wire n_681_v;
  wire n_1471_v;
  wire op_T4_ind_x_v;
  wire n_979_v;
  wire n_973_v;
  wire n_976_v;
  wire op_T__bit_v;
  wire op_T0_iny_dey_v;
  wire n_1270_v;
  wire op_T__cmp_v;
  wire n_1618_v;
  wire op_T0_jsr_v;
  wire n_1610_v;
  wire op_T2_abs_access_v;
  wire n_1613_v;
  wire n_1033_v;
  wire n_1034_v;
  wire n_1037_v;
  wire alub3_v;
  wire n_1038_v;
  wire alub1_v;
  wire alub0_v;
  wire alub7_v;
  wire alub6_v;
  wire alub5_v;
  wire alub4_v;
  wire notalu4_v;
  wire notalu5_v;
  wire notalu6_v;
  wire notalu7_v;
  wire notalu0_v;
  wire notalu1_v;
  wire notalu2_v;
  wire notalu3_v;
  wire x_op_T4_rti_v;
  wire dpc42_DL_ADH_v;
  wire n_769_v;
  wire n_767_v;
  wire n_763_v;
  wire n_762_v;
  wire n_761_v;
  wire n_760_v;
  wire notidl4_v;
  wire notidl3_v;
  wire notidl1_v;
  wire op_T3_abs_idx_ind_v;
  wire op_T2_jsr_v;
  wire DA_C45_v;
  wire n_231_v;
  wire _C78_v;
  wire n_233_v;
  wire n_232_v;
  wire n_236_v;
  wire n_951_v;
  wire n_952_v;
  wire n_953_v;
  wire n_402_v;
  wire n_958_v;
  wire n_959_v;
  wire n_408_v;
  wire n_409_v;
  wire op_T0_eor_v;
  wire pd1_clearIR_v;
  wire abl3_v;
  wire op_T0_jmp_v;
  wire n_1018_v;
  wire n_1549_v;
  wire n_1548_v;
  wire n_1016_v;
  wire p1_v;
  wire p4_v;
  wire __AxB1__C01_v;
  wire op_T2_idx_x_xy_v;
  wire _TWOCYCLE_phi1_v;
  wire op_clv_v;
  wire op_T0_and_v;
  wire n_171_v;
  wire op_T0_clc_sec_v;
  wire _C56_v;
  wire n_1209_v;
  wire n_1206_v;
  wire n_1205_v;
  wire n_1202_v;
  wire n_1500_v;
  wire _ABH2_v;
  wire _ABH4_v;
  wire n_1507_v;
  wire notidl5_v;
  wire n_428_v;
  wire n_424_v;
  wire n_420_v;
  wire n_423_v;
  wire op_sty_cpy_mem_v;
  wire n_1254_v;
  wire dpc18__DAA_v;
  wire n_1720_v;
  wire AxB5_v;
  wire AxB7_v;
  wire AxB1_v;
  wire AxB3_v;
  wire op_T3_ind_y_v;
  wire op_T3_ind_x_v;
  wire n_1566_v;
  wire n_1565_v;
  wire n_1561_v;
  wire n_1560_v;
  wire dpc38_PCLADL_v;
  wire n_1691_v;
  wire n_1697_v;
  wire n_1696_v;
  wire n_1699_v;
  wire x_op_T3_abs_idx_v;
  wire op_from_x_v;
  wire n_855_v;
  wire n_850_v;
  wire n_853_v;
  wire n_852_v;
  wire op_T0_cli_sei_v;
  wire op_T0_ldx_tax_tsx_v;
  wire n_1049_v;
  wire n_1229_v;
  wire n_1593_v;
  wire n_1221_v;
  wire n_1222_v;
  wire n_1223_v;
  wire n_1225_v;
  wire n_1044_v;
  wire n_1594_v;
  wire n_1047_v;
  wire n_198_v;
  wire n_628_v;
  wire n_629_v;
  wire n_626_v;
  wire n_196_v;
  wire n_625_v;
  wire n_190_v;
  wire n_191_v;
  wire n_192_v;
  wire n_621_v;
  wire n_442_v;
  wire n_440_v;
  wire n_441_v;
  wire n_445_v;
  wire DBNeg_v;
  wire op_T0_tsx_v;
  wire notidl7_v;
  wire notidl6_v;
  wire notidl2_v;
  wire n_994_v;
  wire n_995_v;
  wire n_990_v;
  wire n_992_v;
  wire n_993_v;
  wire n_998_v;
  wire n_999_v;
  wire _op_store_v;
  wire n_1501_v;
  wire n_1505_v;
  wire n_1509_v;
  wire op_T0_cpx_inx_v;
  wire n_299_v;
  wire n_298_v;
  wire n_293_v;
  wire n_291_v;
  wire n_871_v;
  wire n_877_v;
  wire n_876_v;
  wire n_875_v;
  wire n_878_v;
  wire n_956_v;

  spice_pin_input pin_4286(nmi, nmi_v, nmi_port_2);
  spice_pin_input pin_4287(irq, irq_v, irq_port_2);
  spice_pin_input pin_4285(rdy, rdy_v, rdy_port_3);
  spice_pin_input pin_4282(clk0, clk0_v, clk0_port_3);
  spice_pin_input pin_4281(so, so_v, so_port_3);
  spice_pin_input pin_4278(res, res_v, res_port_2);

  spice_pin_output pin_4284(clk2out, a(clk2out_v));
  spice_pin_output pin_4283(clk1out, a(clk1out_v));
  spice_pin_output pin_4280(sync, a(sync_v));
  spice_pin_output pin_4268(ab14, a(ab14_v));
  spice_pin_output pin_4264(ab10, a(ab10_v));
  spice_pin_output pin_4266(ab12, a(ab12_v));
  spice_pin_output pin_4260(ab6, a(ab6_v));
  spice_pin_output pin_4261(ab7, a(ab7_v));
  spice_pin_output pin_4262(ab8, a(ab8_v));
  spice_pin_output pin_4263(ab9, a(ab9_v));
  spice_pin_output pin_4269(ab15, a(ab15_v));
  spice_pin_output pin_4265(ab11, a(ab11_v));
  spice_pin_output pin_4267(ab13, a(ab13_v));
  spice_pin_output pin_4279(rw, a(rw_v));
  spice_pin_output pin_4255(ab1, a(ab1_v));
  spice_pin_output pin_4254(ab0, a(ab0_v));
  spice_pin_output pin_4257(ab3, a(ab3_v));
  spice_pin_output pin_4256(ab2, a(ab2_v));
  spice_pin_output pin_4259(ab5, a(ab5_v));
  spice_pin_output pin_4258(ab4, a(ab4_v));

  spice_pin_bidirectional pin_4277(db7_i, db7_o, db7_t, db7_v, db7_port_5);
  spice_pin_bidirectional pin_4276(db6_i, db6_o, db6_t, db6_v, db6_port_5);
  spice_pin_bidirectional pin_4275(db5_i, db5_o, db5_t, db5_v, db5_port_5);
  spice_pin_bidirectional pin_4274(db4_i, db4_o, db4_t, db4_v, db4_port_5);
  spice_pin_bidirectional pin_4273(db3_i, db3_o, db3_t, db3_v, db3_port_5);
  spice_pin_bidirectional pin_4272(db2_i, db2_o, db2_t, db2_v, db2_port_5);
  spice_pin_bidirectional pin_4271(db1_i, db1_o, db1_t, db1_v, db1_port_5);
  spice_pin_bidirectional pin_4270(db0_i, db0_o, db0_t, db0_v, db0_port_5);

  wire [`W-1:0] temp_6390;
  spice_transistor_nmos t989(dpc37_PCLDB_v, idb0_v, a(n_488_v), idb0_port_6, temp_6390);
  wire [`W-1:0] temp_6391;
  spice_transistor_nmos t2363(dpc24_ACSB_v, sb0_v, a(n_146_v), sb0_port_10, temp_6391);
  wire [`W-1:0] temp_6392;
  spice_transistor_nmos t2366(dpc24_ACSB_v, sb3_v, a(n_1654_v), sb3_port_10, temp_6392);
  wire [`W-1:0] temp_6393;
  spice_transistor_nmos t2367(dpc24_ACSB_v, sb4_v, a(n_1344_v), sb4_port_11, temp_6393);
  wire [`W-1:0] temp_6394;
  spice_transistor_nmos t2364(dpc24_ACSB_v, sb1_v, a(n_929_v), sb1_port_9, temp_6394);
  wire [`W-1:0] temp_6395;
  spice_transistor_nmos t2365(dpc24_ACSB_v, a(n_1618_v), sb2_v, temp_6395, sb2_port_9);
  wire [`W-1:0] temp_6396;
  spice_transistor_nmos t2368(dpc24_ACSB_v, sb5_v, a(n_831_v), sb5_port_8, temp_6396);
  wire [`W-1:0] temp_6397;
  spice_transistor_nmos t2369(dpc24_ACSB_v, a(n_326_v), sb6_v, temp_6397, sb6_port_11);
  spice_transistor_nmos_gnd t1184(n_0_ADL1_v, adl1_v, adl1_port_1);
  spice_transistor_nmos t2197(dpc27_SBADH_v, adh4_v, sb4_v, adh4_port_4, sb4_port_9);
  wire [`W-1:0] temp_6398;
  spice_transistor_nmos t374(dpc4_SSB_v, a(n_694_v), sb1_v, temp_6398, sb1_port_2);
  wire [`W-1:0] temp_6399;
  spice_transistor_nmos t2526(dpc38_PCLADL_v, a(n_72_v), adl5_v, temp_6399, adl5_port_4);
  wire [`W-1:0] temp_6400;
  spice_transistor_nmos t2527(dpc38_PCLADL_v, adl6_v, a(n_1458_v), adl6_port_4, temp_6400);
  wire [`W-1:0] temp_6401;
  spice_transistor_nmos t3118(dpc2_XSB_v, a(n_1694_v), sb2_v, temp_6401, sb2_port_10);
  wire [`W-1:0] temp_6402;
  spice_transistor_nmos t3119(dpc2_XSB_v, a(n_242_v), sb3_v, temp_6402, sb3_port_11);
  wire [`W-1:0] temp_6403;
  spice_transistor_nmos t3116(dpc2_XSB_v, a(n_1724_v), sb6_v, temp_6403, sb6_port_12);
  wire [`W-1:0] temp_6404;
  spice_transistor_nmos t3115(dpc2_XSB_v, a(n_578_v), sb5_v, temp_6404, sb5_port_10);
  spice_transistor_nmos_vdd t961(cclk_v, idb3_v, idb3_port_1);
  wire [`W-1:0] temp_6405;
  spice_transistor_nmos t3342(cp1_v, n_1095_v, a(idl4_v), n_1095_port_3, temp_6405);
  spice_transistor_nmos_vdd t3340(cclk_v, sb5_v, sb5_port_12);
  spice_transistor_nmos_vdd t1536(n_520_v, db2_v, db2_port_3);
  wire [`W-1:0] temp_6406;
  spice_transistor_nmos t142(cp1_v, n_1424_v, a(idl2_v), n_1424_port_0, temp_6406);
  spice_transistor_nmos t2254(dpc27_SBADH_v, sb1_v, adh1_v, sb1_port_8, adh1_port_4);
  wire [`W-1:0] temp_6407;
  spice_transistor_nmos g_4819((cp1_v&ADH_ABH_v), a(n_1668_v), _ABH0_v, temp_6407, _ABH0_port_3);
  wire [`W-1:0] temp_6408;
  spice_transistor_nmos t941(dpc16_EORS_v, a(n_1469_v), n_277_v, temp_6408, n_277_port_1);
  wire [`W-1:0] temp_6409;
  spice_transistor_nmos t940(dpc16_EORS_v, a(__AxB_4_v), n_296_v, temp_6409, n_296_port_0);
  wire [`W-1:0] temp_6410;
  spice_transistor_nmos t943(dpc16_EORS_v, n_304_v, a(n_177_v), n_304_port_1, temp_6410);
  wire [`W-1:0] temp_6411;
  spice_transistor_nmos t942(dpc16_EORS_v, a(__AxB_6_v), n_722_v, temp_6411, n_722_port_1);
  wire [`W-1:0] temp_6412;
  spice_transistor_nmos t128(dpc4_SSB_v, a(n_1389_v), sb2_v, temp_6412, sb2_port_1);
  wire [`W-1:0] temp_6413;
  spice_transistor_nmos t127(dpc4_SSB_v, a(n_998_v), sb3_v, temp_6413, sb3_port_1);
  wire [`W-1:0] temp_6414;
  spice_transistor_nmos t1723(dpc5_SADL_v, adl3_v, a(n_998_v), adl3_port_3, temp_6414);
  wire [`W-1:0] temp_6415;
  spice_transistor_nmos t1722(dpc5_SADL_v, adl4_v, a(n_3_v), adl4_port_4, temp_6415);
  wire [`W-1:0] temp_6416;
  spice_transistor_nmos t1721(dpc5_SADL_v, adl5_v, a(n_280_v), adl5_port_3, temp_6416);
  wire [`W-1:0] temp_6417;
  spice_transistor_nmos t1727(dpc5_SADL_v, a(n_721_v), adl7_v, temp_6417, adl7_port_2);
  wire [`W-1:0] temp_6418;
  spice_transistor_nmos t1724(dpc5_SADL_v, adl2_v, a(n_1389_v), adl2_port_3, temp_6418);
  wire [`W-1:0] temp_6419;
  spice_transistor_nmos g_4857((ADH_ABH_v&cp1_v), _ABH6_v, a(n_880_v), _ABH6_port_3, temp_6419);
  wire [`W-1:0] temp_6420;
  spice_transistor_nmos g_4858((ADH_ABH_v&cp1_v), _ABH3_v, a(n_883_v), _ABH3_port_3, temp_6420);
  wire [`W-1:0] temp_6421;
  spice_transistor_nmos t83(H1x1_v, idb2_v, a(Pout2_v), idb2_port_0, temp_6421);
  wire [`W-1:0] temp_6422;
  spice_transistor_nmos t2257(dpc0_YSB_v, a(n_1251_v), sb7_v, temp_6422, sb7_port_8);
  wire [`W-1:0] temp_6423;
  spice_transistor_nmos t2745(dpc37_PCLDB_v, a(n_723_v), idb3_v, temp_6423, idb3_port_9);
  wire [`W-1:0] temp_6424;
  spice_transistor_nmos t2746(dpc37_PCLDB_v, a(n_976_v), idb1_v, temp_6424, idb1_port_8);
  spice_transistor_nmos_vdd t2598(cclk_v, idb6_v, idb6_port_9);
  wire [`W-1:0] temp_6425;
  spice_transistor_nmos t2592(dpc13_ORS_v, a(n_404_v), n_296_v, temp_6425, n_296_port_5);
  spice_transistor_nmos_gnd t1024(n_471_v, db6_v, db6_port_0);
  wire [`W-1:0] temp_6426;
  spice_transistor_nmos t1505(dpc0_YSB_v, a(n_1491_v), sb2_v, temp_6426, sb2_port_3);
  spice_transistor_nmos_vdd t3504(cclk_v, idb4_v, idb4_port_10);
  spice_transistor_nmos_vdd t3502(cclk_v, sb2_v, sb2_port_12);
  spice_transistor_nmos_vdd t1760(cclk_v, idb2_v, idb2_port_4);
  wire [`W-1:0] temp_6427;
  spice_transistor_nmos t3195(dpc4_SSB_v, a(n_332_v), sb0_v, temp_6427, sb0_port_12);
  spice_transistor_nmos_vdd t2028(cclk_v, adh7_v, adh7_port_2);
  wire [`W-1:0] temp_6428;
  spice_transistor_nmos t521(dpc21_ADDADL_v, adl3_v, a(alu3_v), adl3_port_0, temp_6428);
  wire [`W-1:0] temp_6429;
  spice_transistor_nmos t520(cp1_v, n_87_v, a(idl1_v), n_87_port_1, temp_6429);
  wire [`W-1:0] temp_6430;
  spice_transistor_nmos t1590(dpc14_SRS_v, a(aluanandb1_v), notaluoutmux0_v, temp_6430, notaluoutmux0_port_2);
  wire [`W-1:0] temp_6431;
  spice_transistor_nmos t1591(dpc14_SRS_v, notaluoutmux1_v, a(n_681_v), notaluoutmux1_port_2, temp_6431);
  wire [`W-1:0] temp_6432;
  spice_transistor_nmos t1592(dpc14_SRS_v, a(n_350_v), n_740_v, temp_6432, n_740_port_3);
  wire [`W-1:0] temp_6433;
  spice_transistor_nmos t1593(dpc14_SRS_v, n_1071_v, a(n_1063_v), n_1071_port_4, temp_6433);
  wire [`W-1:0] temp_6434;
  spice_transistor_nmos t1594(dpc14_SRS_v, n_296_v, a(n_477_v), n_296_port_3, temp_6434);
  wire [`W-1:0] temp_6435;
  spice_transistor_nmos t1595(dpc14_SRS_v, n_277_v, a(n_336_v), n_277_port_3, temp_6435);
  wire [`W-1:0] temp_6436;
  spice_transistor_nmos t1596(dpc14_SRS_v, n_722_v, a(n_1318_v), n_722_port_4, temp_6436);
  spice_transistor_nmos t588(dpc43_DL_DB_v, idb3_v, n_1661_v, idb3_port_0, n_1661_port_1);
  spice_transistor_nmos t585(dpc43_DL_DB_v, idb0_v, n_719_v, idb0_port_5, n_719_port_2);
  spice_transistor_nmos_gnd t3038(n_147_v, db4_v, db4_port_3);
  wire [`W-1:0] temp_6437;
  spice_transistor_nmos t1961(dpc5_SADL_v, adl0_v, a(n_332_v), adl0_port_4, temp_6437);
  wire [`W-1:0] temp_6438;
  spice_transistor_nmos g_4726((ADH_ABH_v&cp1_v), _ABH7_v, a(n_494_v), _ABH7_port_3, temp_6438);
  wire [`W-1:0] temp_6439;
  spice_transistor_nmos t2551(dpc32_PCHADH_v, adh3_v, a(n_141_v), adh3_port_6, temp_6439);
  wire [`W-1:0] temp_6440;
  spice_transistor_nmos t2550(dpc32_PCHADH_v, adh4_v, a(n_27_v), adh4_port_6, temp_6440);
  wire [`W-1:0] temp_6441;
  spice_transistor_nmos t2553(dpc32_PCHADH_v, adh1_v, a(n_209_v), adh1_port_6, temp_6441);
  wire [`W-1:0] temp_6442;
  spice_transistor_nmos t2552(dpc32_PCHADH_v, adh2_v, a(n_1496_v), adh2_port_6, temp_6442);
  wire [`W-1:0] temp_6443;
  spice_transistor_nmos t1208(dpc20_ADDSB06_v, a(alu6_v), sb6_v, temp_6443, sb6_port_6);
  wire [`W-1:0] temp_6444;
  spice_transistor_nmos t1209(dpc20_ADDSB06_v, a(alu5_v), sb5_v, temp_6444, sb5_port_3);
  spice_transistor_nmos_vdd t2353(n_298_v, db7_v, db7_port_3);
  wire [`W-1:0] temp_6445;
  spice_transistor_nmos t3225(dpc2_XSB_v, a(n_1709_v), sb1_v, temp_6445, sb1_port_12);
  wire [`W-1:0] temp_6446;
  spice_transistor_nmos t3489(dpc13_ORS_v, a(aluanorb1_v), notaluoutmux1_v, temp_6446, notaluoutmux1_port_5);
  spice_transistor_nmos_gnd t1887(n_643_v, db3_v, db3_port_3);
  spice_transistor_nmos_gnd t1089(n_37_v, db2_v, db2_port_2);
  spice_transistor_nmos_gnd g_4913((v(n_975_v)|(n_312_v&cclk_v)), n_854_v, n_854_port_6);
  wire [`W-1:0] temp_6447;
  spice_transistor_nmos t2218(dpc15_ANDS_v, a(n_336_v), n_722_v, temp_6447, n_722_port_5);
  wire [`W-1:0] temp_6448;
  spice_transistor_nmos t2219(dpc15_ANDS_v, n_304_v, a(n_1318_v), n_304_port_4, temp_6448);
  wire [`W-1:0] temp_6449;
  spice_transistor_nmos t2216(dpc15_ANDS_v, a(n_1063_v), n_296_v, temp_6449, n_296_port_4);
  wire [`W-1:0] temp_6450;
  spice_transistor_nmos t2217(dpc15_ANDS_v, n_277_v, a(n_477_v), n_277_port_4, temp_6450);
  wire [`W-1:0] temp_6451;
  spice_transistor_nmos t2214(dpc15_ANDS_v, a(n_681_v), n_740_v, temp_6451, n_740_port_4);
  wire [`W-1:0] temp_6452;
  spice_transistor_nmos t2747(dpc37_PCLDB_v, idb7_v, a(n_1647_v), idb7_port_9, temp_6452);
  wire [`W-1:0] temp_6453;
  spice_transistor_nmos t2212(dpc15_ANDS_v, a(aluanandb0_v), notaluoutmux0_v, temp_6453, notaluoutmux0_port_5);
  wire [`W-1:0] temp_6454;
  spice_transistor_nmos t2213(dpc15_ANDS_v, a(aluanandb1_v), notaluoutmux1_v, temp_6454, notaluoutmux1_port_4);
  wire [`W-1:0] temp_6455;
  spice_transistor_nmos t2554(dpc32_PCHADH_v, adh0_v, a(n_1722_v), adh0_port_6, temp_6455);
  spice_transistor_nmos_gnd g_4937(((n_284_v&cclk_v)|v(n_297_v)), NMIP_v, NMIP_port_7);
  wire [`W-1:0] temp_6456;
  spice_transistor_nmos t2235(dpc26_ACDB_v, a(n_146_v), idb0_v, temp_6456, idb0_port_8);
  wire [`W-1:0] temp_6457;
  spice_transistor_nmos t2236(dpc26_ACDB_v, a(n_929_v), idb1_v, temp_6457, idb1_port_5);
  wire [`W-1:0] temp_6458;
  spice_transistor_nmos t2237(dpc26_ACDB_v, a(n_1618_v), idb2_v, temp_6458, idb2_port_6);
  wire [`W-1:0] temp_6459;
  spice_transistor_nmos t2238(dpc26_ACDB_v, a(n_1654_v), idb3_v, temp_6459, idb3_port_6);
  wire [`W-1:0] temp_6460;
  spice_transistor_nmos t2239(dpc26_ACDB_v, idb4_v, a(n_1344_v), idb4_port_6, temp_6460);
  wire [`W-1:0] temp_6461;
  spice_transistor_nmos t2724(cp1_v, n_1147_v, a(idl7_v), n_1147_port_3, temp_6461);
  spice_transistor_nmos_vdd t426(cclk_v, adh4_v, adh4_port_2);
  spice_transistor_nmos_vdd t427(cclk_v, adl5_v, adl5_port_0);
  spice_transistor_nmos_vdd t227(cclk_v, idb0_v, idb0_port_1);
  spice_transistor_nmos_gnd t2537(n_0_ADL2_v, adl2_v, adl2_port_6);
  wire [`W-1:0] temp_6462;
  spice_transistor_nmos t2532(dpc38_PCLADL_v, a(n_723_v), adl3_v, temp_6462, adl3_port_4);
  wire [`W-1:0] temp_6463;
  spice_transistor_nmos t2531(dpc38_PCLADL_v, adl2_v, a(n_481_v), adl2_port_5, temp_6463);
  wire [`W-1:0] temp_6464;
  spice_transistor_nmos t2530(dpc38_PCLADL_v, a(n_976_v), adl1_v, temp_6464, adl1_port_5);
  spice_transistor_nmos t1860(dpc25_SBDB_v, idb5_v, sb5_v, idb5_port_4, sb5_port_6);
  spice_transistor_nmos t1861(dpc25_SBDB_v, idb6_v, sb6_v, idb6_port_5, sb6_port_8);
  spice_transistor_nmos t1862(dpc25_SBDB_v, sb7_v, idb7_v, sb7_port_5, idb7_port_4);
  spice_transistor_nmos t589(dpc43_DL_DB_v, idb4_v, n_1095_v, idb4_port_0, n_1095_port_1);
  spice_transistor_nmos t587(dpc43_DL_DB_v, idb2_v, n_1424_v, idb2_port_1, n_1424_port_2);
  spice_transistor_nmos t586(dpc43_DL_DB_v, idb1_v, n_87_v, idb1_port_0, n_87_port_2);
  spice_transistor_nmos_vdd t2270(cclk_v, idb5_v, idb5_port_6);
  wire [`W-1:0] temp_6465;
  spice_transistor_nmos t268(H1x1_v, idb0_v, a(Pout0_v), idb0_port_2, temp_6465);
  wire [`W-1:0] temp_6466;
  spice_transistor_nmos t2130(H1x1_v, a(p6_v), idb6_v, temp_6466, idb6_port_6);
  spice_transistor_nmos_vdd t1118(cclk_v, sb3_v, sb3_port_3);
  wire [`W-1:0] temp_6467;
  spice_transistor_nmos t1110(dpc17_SUMS_v, a(__AxBxC_4_v), n_296_v, temp_6467, n_296_port_1);
  wire [`W-1:0] temp_6468;
  spice_transistor_nmos t1111(dpc17_SUMS_v, a(__AxBxC_5_v), n_277_v, temp_6468, n_277_port_2);
  wire [`W-1:0] temp_6469;
  spice_transistor_nmos t1112(dpc17_SUMS_v, n_722_v, a(__AxBxC_6_v), n_722_port_2, temp_6469);
  wire [`W-1:0] temp_6470;
  spice_transistor_nmos t1113(dpc17_SUMS_v, n_304_v, a(__AxBxC_7_v), n_304_port_2, temp_6470);
  wire [`W-1:0] temp_6471;
  spice_transistor_nmos t2762(cp1_v, n_1661_v, a(idl3_v), n_1661_port_3, temp_6471);
  spice_transistor_nmos_gnd t2487(dpc29_0ADH17_v, adh5_v, adh5_port_3);
  spice_transistor_nmos_gnd t2486(dpc29_0ADH17_v, adh2_v, adh2_port_5);
  spice_transistor_nmos_gnd t2485(dpc29_0ADH17_v, adh3_v, adh3_port_5);
  wire [`W-1:0] temp_6472;
  spice_transistor_nmos t2334(dpc37_PCLDB_v, idb4_v, a(n_208_v), idb4_port_7, temp_6472);
  spice_transistor_nmos_gnd t2488(dpc29_0ADH17_v, adh4_v, adh4_port_5);
  spice_transistor_nmos_vdd t382(n_1076_v, db4_v, db4_port_0);
  wire [`W-1:0] temp_6473;
  spice_transistor_nmos t385(dpc4_SSB_v, a(n_280_v), sb5_v, temp_6473, sb5_port_2);
  wire [`W-1:0] temp_6474;
  spice_transistor_nmos t3142(dpc0_YSB_v, a(n_767_v), sb1_v, temp_6474, sb1_port_11);
  spice_transistor_nmos_gnd t2819(n_0_ADL0_v, adl0_v, adl0_port_7);
  spice_transistor_nmos_vdd t1548(cclk_v, sb7_v, sb7_port_3);
  wire [`W-1:0] temp_6475;
  spice_transistor_nmos t993(dpc37_PCLDB_v, idb2_v, a(n_481_v), idb2_port_3, temp_6475);
  wire [`W-1:0] temp_6476;
  spice_transistor_nmos t2371(dpc5_SADL_v, adl1_v, a(n_694_v), adl1_port_4, temp_6476);
  wire [`W-1:0] temp_6477;
  spice_transistor_nmos t2370(dpc24_ACSB_v, a(n_1592_v), sb7_v, temp_6477, sb7_port_9);
  spice_transistor_nmos t2199(dpc27_SBADH_v, adh2_v, sb2_v, adh2_port_4, sb2_port_8);
  spice_transistor_nmos t2198(dpc27_SBADH_v, adh3_v, sb3_v, adh3_port_3, sb3_port_9);
  spice_transistor_nmos t2191(dpc27_SBADH_v, sb6_v, adh6_v, sb6_port_9, adh6_port_3);
  spice_transistor_nmos t2190(dpc27_SBADH_v, adh7_v, sb7_v, adh7_port_3, sb7_port_7);
  spice_transistor_nmos t2193(dpc27_SBADH_v, adh0_v, sb0_v, adh0_port_2, sb0_port_9);
  wire [`W-1:0] temp_6478;
  spice_transistor_nmos t1508(dpc0_YSB_v, sb3_v, a(n_1531_v), sb3_port_5, temp_6478);
  spice_transistor_nmos_vdd t154(n_798_v, db1_v, db1_port_1);
  wire [`W-1:0] temp_6479;
  spice_transistor_nmos t1333(H1x1_v, a(Pout1_v), idb1_v, temp_6479, idb1_port_3);
  wire [`W-1:0] temp_6480;
  spice_transistor_nmos g_4803((ADH_ABH_v&cp1_v), _ABH5_v, a(n_254_v), _ABH5_port_3, temp_6480);
  wire [`W-1:0] temp_6481;
  spice_transistor_nmos t3120(dpc2_XSB_v, a(n_436_v), sb4_v, temp_6481, sb4_port_12);
  spice_transistor_nmos_vdd t3352(cclk_v, adh6_v, adh6_port_6);
  spice_transistor_nmos_vdd t3353(cclk_v, adl7_v, adl7_port_7);
  wire [`W-1:0] temp_6482;
  spice_transistor_nmos t132(dpc4_SSB_v, a(n_721_v), sb7_v, temp_6482, sb7_port_0);
  wire [`W-1:0] temp_6483;
  spice_transistor_nmos t133(dpc4_SSB_v, a(n_618_v), sb6_v, temp_6483, sb6_port_2);
  wire [`W-1:0] temp_6484;
  spice_transistor_nmos t136(dpc4_SSB_v, a(n_3_v), sb4_v, temp_6484, sb4_port_3);
  wire [`W-1:0] temp_6485;
  spice_transistor_nmos t546(dpc13_ORS_v, a(n_649_v), n_1071_v, temp_6485, n_1071_port_0);
  spice_transistor_nmos_vdd t1712(n_1325_v, db0_v, db0_port_1);
  spice_transistor_nmos_gnd t301(n_612_v, db5_v, db5_port_0);
  wire [`W-1:0] temp_6486;
  spice_transistor_nmos t936(dpc16_EORS_v, a(__AxB_0_v), notaluoutmux0_v, temp_6486, notaluoutmux0_port_0);
  wire [`W-1:0] temp_6487;
  spice_transistor_nmos t937(dpc16_EORS_v, notaluoutmux1_v, a(n_953_v), notaluoutmux1_port_0, temp_6487);
  wire [`W-1:0] temp_6488;
  spice_transistor_nmos t938(dpc16_EORS_v, a(__AxB_2_v), n_740_v, temp_6488, n_740_port_1);
  wire [`W-1:0] temp_6489;
  spice_transistor_nmos t939(dpc16_EORS_v, a(n_884_v), n_1071_v, temp_6489, n_1071_port_2);
  wire [`W-1:0] temp_6490;
  spice_transistor_nmos t2895(dpc20_ADDSB06_v, a(alu1_v), sb1_v, temp_6490, sb1_port_10);
  wire [`W-1:0] temp_6491;
  spice_transistor_nmos t2897(dpc20_ADDSB06_v, a(alu0_v), sb0_v, temp_6491, sb0_port_11);
  spice_transistor_nmos_vdd t2336(cclk_v, adh3_v, adh3_port_4);
  spice_transistor_nmos t1484(dpc41_DL_ADL_v, adl2_v, n_1424_v, adl2_port_2, n_1424_port_3);
  spice_transistor_nmos_vdd t1739(cclk_v, sb1_v, sb1_port_6);
  wire [`W-1:0] temp_6492;
  spice_transistor_nmos t329(dpc0_YSB_v, a(n_564_v), sb0_v, temp_6492, sb0_port_1);
  wire [`W-1:0] temp_6493;
  spice_transistor_nmos t321(dpc21_ADDADL_v, a(alu2_v), adl2_v, temp_6493, adl2_port_0);
  wire [`W-1:0] temp_6494;
  spice_transistor_nmos t323(dpc21_ADDADL_v, adl0_v, a(alu0_v), adl0_port_0, temp_6494);
  wire [`W-1:0] temp_6495;
  spice_transistor_nmos t322(dpc21_ADDADL_v, adl1_v, a(alu1_v), adl1_port_0, temp_6495);
  wire [`W-1:0] temp_6496;
  spice_transistor_nmos t2215(dpc15_ANDS_v, a(n_350_v), n_1071_v, temp_6496, n_1071_port_5);
  spice_transistor_nmos_gnd t2442(dpc28_0ADH0_v, adh0_v, adh0_port_3);
  wire [`W-1:0] temp_6497;
  spice_transistor_nmos t2918(dpc33_PCHDB_v, idb7_v, a(n_1206_v), idb7_port_10, temp_6497);
  wire [`W-1:0] temp_6498;
  spice_transistor_nmos t2915(dpc33_PCHDB_v, a(n_27_v), idb4_v, temp_6498, idb4_port_9);
  wire [`W-1:0] temp_6499;
  spice_transistor_nmos t2914(dpc33_PCHDB_v, a(n_141_v), idb3_v, temp_6499, idb3_port_10);
  wire [`W-1:0] temp_6500;
  spice_transistor_nmos t2917(dpc33_PCHDB_v, idb6_v, a(n_652_v), idb6_port_11, temp_6500);
  wire [`W-1:0] temp_6501;
  spice_transistor_nmos t2916(dpc33_PCHDB_v, a(n_1301_v), idb5_v, temp_6501, idb5_port_9);
  wire [`W-1:0] temp_6502;
  spice_transistor_nmos t2911(dpc33_PCHDB_v, a(n_1722_v), idb0_v, temp_6502, idb0_port_10);
  wire [`W-1:0] temp_6503;
  spice_transistor_nmos t2913(dpc33_PCHDB_v, idb2_v, a(n_1496_v), idb2_port_10, temp_6503);
  wire [`W-1:0] temp_6504;
  spice_transistor_nmos t2912(dpc33_PCHDB_v, idb1_v, a(n_209_v), idb1_port_9, temp_6504);
  wire [`W-1:0] temp_6505;
  spice_transistor_nmos t499(dpc13_ORS_v, n_722_v, a(n_1084_v), n_722_port_0, temp_6505);
  wire [`W-1:0] temp_6506;
  spice_transistor_nmos t1752(cp1_v, n_1014_v, a(idl6_v), n_1014_port_3, temp_6506);
  spice_transistor_nmos_vdd t1750(cclk_v, adl2_v, adl2_port_4);
  spice_transistor_nmos_vdd t1757(n_373_v, db5_v, db5_port_4);
  spice_transistor_nmos t3181(dpc27_SBADH_v, adh5_v, sb5_v, adh5_port_5, sb5_port_11);
  wire [`W-1:0] temp_6507;
  spice_transistor_nmos t3182(dpc5_SADL_v, a(n_618_v), adl6_v, temp_6507, adl6_port_5);
  spice_transistor_nmos_vdd t1587(cclk_v, sb0_v, sb0_port_4);
  spice_transistor_nmos_vdd t1911(cclk_v, adh2_v, adh2_port_3);
  spice_transistor_nmos t1485(dpc41_DL_ADL_v, adl0_v, n_719_v, adl0_port_3, n_719_port_3);
  spice_transistor_nmos t1482(dpc41_DL_ADL_v, adl4_v, n_1095_v, adl4_port_3, n_1095_port_2);
  spice_transistor_nmos t1483(dpc41_DL_ADL_v, adl1_v, n_87_v, adl1_port_2, n_87_port_3);
  spice_transistor_nmos t1481(dpc41_DL_ADL_v, adl3_v, n_1661_v, adl3_port_2, n_1661_port_2);
  wire [`W-1:0] temp_6508;
  spice_transistor_nmos t1211(dpc20_ADDSB06_v, a(alu3_v), sb3_v, temp_6508, sb3_port_4);
  wire [`W-1:0] temp_6509;
  spice_transistor_nmos t1210(dpc20_ADDSB06_v, sb4_v, a(alu4_v), sb4_port_5, temp_6509);
  spice_transistor_nmos_gnd t2490(dpc29_0ADH17_v, adh7_v, adh7_port_4);
  spice_transistor_nmos_gnd t2491(dpc29_0ADH17_v, adh6_v, adh6_port_4);
  wire [`W-1:0] temp_6510;
  spice_transistor_nmos t2320(dpc37_PCLDB_v, a(n_72_v), idb5_v, temp_6510, idb5_port_7);
  spice_transistor_nmos_gnd g_4944((v(n_807_v)|(cclk_v&n_538_v)), n_330_v, n_330_port_7);
  spice_transistor_nmos_gnd t1792(n_1501_v, db7_v, db7_port_1);
  wire [`W-1:0] temp_6511;
  spice_transistor_nmos g_4717((ADH_ABH_v&cp1_v), _ABH1_v, a(n_1267_v), _ABH1_port_3, temp_6511);
  spice_transistor_nmos_vdd t299(cclk_v, adh0_v, adh0_port_1);
  wire [`W-1:0] temp_6512;
  spice_transistor_nmos t296(cp1_v, n_719_v, a(idl0_v), n_719_port_1, temp_6512);
  wire [`W-1:0] temp_6513;
  spice_transistor_nmos t2548(dpc32_PCHADH_v, adh6_v, a(n_652_v), adh6_port_5, temp_6513);
  wire [`W-1:0] temp_6514;
  spice_transistor_nmos t2549(dpc32_PCHADH_v, adh5_v, a(n_1301_v), adh5_port_4, temp_6514);
  wire [`W-1:0] temp_6515;
  spice_transistor_nmos t2547(dpc32_PCHADH_v, adh7_v, a(n_1206_v), adh7_port_5, temp_6515);
  wire [`W-1:0] temp_6516;
  spice_transistor_nmos t1958(dpc13_ORS_v, a(aluanorb0_v), notaluoutmux0_v, temp_6516, notaluoutmux0_port_3);
  wire [`W-1:0] temp_6517;
  spice_transistor_nmos t1957(dpc13_ORS_v, n_304_v, a(n_1398_v), n_304_port_3, temp_6517);
  spice_transistor_nmos_vdd t75(dpc14_SRS_v, n_304_v, n_304_port_0);
  spice_transistor_nmos_vdd t1602(cclk_v, idb7_v, idb7_port_3);
  spice_transistor_nmos_gnd g_4907((v(n_330_v)|(cclk_v&n_1599_v)), n_807_v, n_807_port_5);
  spice_transistor_nmos_gnd g_4906((v(NMIP_v)|(n_1392_v&cclk_v)), n_297_v, n_297_port_5);
  spice_transistor_nmos_vdd t3442(n_7_v, db6_v, db6_port_4);
  spice_transistor_nmos_vdd t3331(cclk_v, idb1_v, idb1_port_10);
  spice_transistor_nmos_vdd t2221(cclk_v, adl1_v, adl1_port_3);
  spice_transistor_nmos_vdd t2736(cclk_v, adl0_v, adl0_port_6);
  spice_transistor_nmos_vdd t416(cclk_v, sb6_v, sb6_port_4);
  spice_transistor_nmos t1859(dpc25_SBDB_v, idb4_v, sb4_v, idb4_port_4, sb4_port_8);
  spice_transistor_nmos t1858(dpc25_SBDB_v, sb3_v, idb3_v, sb3_port_7, idb3_port_3);
  spice_transistor_nmos t1855(dpc25_SBDB_v, sb0_v, idb0_v, sb0_port_6, idb0_port_7);
  spice_transistor_nmos t1857(dpc25_SBDB_v, idb2_v, sb2_v, idb2_port_5, sb2_port_7);
  spice_transistor_nmos t1856(dpc25_SBDB_v, sb1_v, idb1_v, sb1_port_7, idb1_port_4);
  spice_transistor_nmos t1677(dpc41_DL_ADL_v, adl5_v, n_1387_v, adl5_port_2, n_1387_port_2);
  spice_transistor_nmos_gnd g_4923((v(n_854_v)|(cclk_v&n_995_v)), n_975_v, n_975_port_6);
  wire [`W-1:0] temp_6518;
  spice_transistor_nmos t528(dpc21_ADDADL_v, adl6_v, a(alu6_v), adl6_port_1, temp_6518);
  wire [`W-1:0] temp_6519;
  spice_transistor_nmos t527(dpc21_ADDADL_v, adl5_v, a(alu5_v), adl5_port_1, temp_6519);
  wire [`W-1:0] temp_6520;
  spice_transistor_nmos t526(dpc21_ADDADL_v, a(alu7_v), adl7_v, temp_6520, adl7_port_0);
  wire [`W-1:0] temp_6521;
  spice_transistor_nmos t522(dpc21_ADDADL_v, adl4_v, a(alu4_v), adl4_port_1, temp_6521);
  wire [`W-1:0] temp_6522;
  spice_transistor_nmos t2241(dpc26_ACDB_v, a(n_326_v), idb6_v, temp_6522, idb6_port_7);
  wire [`W-1:0] temp_6523;
  spice_transistor_nmos t2240(dpc26_ACDB_v, a(n_831_v), idb5_v, temp_6523, idb5_port_5);
  wire [`W-1:0] temp_6524;
  spice_transistor_nmos t432(dpc2_XSB_v, a(n_1169_v), sb0_v, temp_6524, sb0_port_2);
  spice_transistor_nmos t2863(cclk_v, n_633_v, n_1059_v, n_633_port_0, n_1059_port_0);
  spice_transistor_nmos t238(dpc42_DL_ADH_v, adh7_v, n_1147_v, adh7_port_0, n_1147_port_0);
  spice_transistor_nmos t237(dpc42_DL_ADH_v, adh6_v, n_1014_v, adh6_port_0, n_1014_port_0);
  spice_transistor_nmos t236(dpc42_DL_ADH_v, adh5_v, n_1387_v, adh5_port_0, n_1387_port_0);
  spice_transistor_nmos t235(dpc42_DL_ADH_v, adh4_v, n_1095_v, adh4_port_0, n_1095_port_0);
  spice_transistor_nmos t234(dpc42_DL_ADH_v, adh3_v, n_1661_v, adh3_port_0, n_1661_port_0);
  spice_transistor_nmos t233(dpc42_DL_ADH_v, adh2_v, n_1424_v, adh2_port_0, n_1424_port_1);
  spice_transistor_nmos t232(dpc42_DL_ADH_v, adh1_v, n_87_v, adh1_port_0, n_87_port_0);
  spice_transistor_nmos t231(dpc42_DL_ADH_v, adh0_v, n_719_v, adh0_port_0, n_719_port_0);
  spice_transistor_nmos_vdd t36(cclk_v, sb4_v, sb4_port_0);
  wire [`W-1:0] temp_6525;
  spice_transistor_nmos t2528(dpc38_PCLADL_v, a(n_1647_v), adl7_v, temp_6525, adl7_port_5);
  wire [`W-1:0] temp_6526;
  spice_transistor_nmos t2529(dpc38_PCLADL_v, adl0_v, a(n_488_v), adl0_port_5, temp_6526);
  wire [`W-1:0] temp_6527;
  spice_transistor_nmos t3384(dpc20_ADDSB06_v, a(alu2_v), sb2_v, temp_6527, sb2_port_11);
  spice_transistor_nmos t1876(dpc41_DL_ADL_v, n_1147_v, adl7_v, n_1147_port_2, adl7_port_3);
  wire [`W-1:0] temp_6528;
  spice_transistor_nmos t1384(dpc37_PCLDB_v, a(n_1458_v), idb6_v, temp_6528, idb6_port_3);
  spice_transistor_nmos t592(dpc43_DL_DB_v, idb7_v, n_1147_v, idb7_port_2, n_1147_port_1);
  spice_transistor_nmos t590(dpc43_DL_DB_v, idb5_v, n_1387_v, idb5_port_2, n_1387_port_1);
  spice_transistor_nmos t591(dpc43_DL_DB_v, idb6_v, n_1014_v, idb6_port_0, n_1014_port_1);
  wire [`W-1:0] temp_6529;
  spice_transistor_nmos t82(H1x1_v, a(p7_v), idb7_v, temp_6529, idb7_port_0);
  wire [`W-1:0] temp_6530;
  spice_transistor_nmos t2263(dpc0_YSB_v, a(n_733_v), sb5_v, temp_6530, sb5_port_7);
  wire [`W-1:0] temp_6531;
  spice_transistor_nmos t2262(dpc0_YSB_v, a(n_518_v), sb6_v, temp_6531, sb6_port_10);
  wire [`W-1:0] temp_6532;
  spice_transistor_nmos t2260(dpc0_YSB_v, a(n_658_v), sb4_v, temp_6532, sb4_port_10);
  spice_transistor_nmos_vdd t456(cclk_v, adh1_v, adh1_port_2);
  wire [`W-1:0] temp_6533;
  spice_transistor_nmos t455(dpc2_XSB_v, a(n_871_v), sb7_v, temp_6533, sb7_port_1);
  spice_transistor_nmos_gnd t3410(n_794_v, db1_v, db1_port_4);
  spice_transistor_nmos_vdd t1679(n_42_v, db3_v, db3_port_2);
  wire [`W-1:0] temp_6534;
  spice_transistor_nmos t2595(dpc13_ORS_v, a(n_1632_v), n_277_v, temp_6534, n_277_port_5);
  spice_transistor_nmos t1676(dpc41_DL_ADL_v, adl6_v, n_1014_v, adl6_port_2, n_1014_port_2);
  wire [`W-1:0] temp_6535;
  spice_transistor_nmos t2108(cp1_v, n_1387_v, a(idl5_v), n_1387_port_3, temp_6535);
  spice_transistor_nmos_vdd t1101(cclk_v, adl3_v, adl3_port_1);
  wire [`W-1:0] temp_6536;
  spice_transistor_nmos t1107(dpc17_SUMS_v, a(__AxBxC_1_v), notaluoutmux1_v, temp_6536, notaluoutmux1_port_1);
  wire [`W-1:0] temp_6537;
  spice_transistor_nmos t1106(dpc17_SUMS_v, a(__AxBxC_0_v), notaluoutmux0_v, temp_6537, notaluoutmux0_port_1);
  wire [`W-1:0] temp_6538;
  spice_transistor_nmos t1109(dpc17_SUMS_v, a(__AxBxC_3_v), n_1071_v, temp_6538, n_1071_port_3);
  wire [`W-1:0] temp_6539;
  spice_transistor_nmos t1108(dpc17_SUMS_v, a(__AxBxC_2_v), n_740_v, temp_6539, n_740_port_2);
  spice_transistor_nmos_vdd t279(cclk_v, adl4_v, adl4_port_0);
  wire [`W-1:0] temp_6540;
  spice_transistor_nmos t2525(dpc38_PCLADL_v, adl4_v, a(n_208_v), adl4_port_5, temp_6540);
  spice_transistor_nmos_gnd t3473(n_1072_v, db0_v, db0_port_4);
  wire [`W-1:0] temp_6541;
  spice_transistor_nmos t2129(H1x1_v, a(Pout3_v), idb3_v, temp_6541, idb3_port_5);
  wire [`W-1:0] temp_6542;
  spice_transistor_nmos t2127(H1x1_v, a(p4_v), idb4_v, temp_6542, idb4_port_5);
  spice_transistor_nmos_gnd t398(dpc29_0ADH17_v, adh1_v, adh1_port_1);
  wire [`W-1:0] temp_6543;
  spice_transistor_nmos t2242(dpc26_ACDB_v, a(n_1592_v), idb7_v, temp_6543, idb7_port_7);
  wire [`W-1:0] temp_6544;
  spice_transistor_nmos t538(dpc13_ORS_v, n_740_v, a(n_1691_v), n_740_port_0, temp_6544);
  spice_transistor_nmos_vdd t2148(cclk_v, adh5_v, adh5_port_2);
  spice_transistor_nmos_vdd t2149(cclk_v, adl6_v, adl6_port_3);
  wire [`W-1:0] temp_6545;
  spice_transistor_nmos t2053(dpc19_ADDSB7_v, a(alu7_v), sb7_v, temp_6545, sb7_port_6);

  spice_pullup pullup_3283(rdy_v, rdy_port_2);
  spice_pullup pullup_3714(n_807_v, n_807_port_3);
  spice_pullup pullup_4226(so_v, so_port_2);
  spice_pullup pullup_3815(n_975_v, n_975_port_3);
  spice_pullup pullup_3412(n_297_v, n_297_port_3);
  spice_pullup pullup_3435(n_330_v, n_330_port_4);
  spice_pullup pullup_3746(n_854_v, n_854_port_4);
  spice_pullup pullup_3848(NMIP_v, NMIP_port_4);

  spice_latch latch_5130(eclk,ereset, cclk_v, op_EORS_v, n_982_v);
  spice_latch latch_5131(eclk,ereset, cclk_v, n_1110_v, pipeUNK01_v);
  spice_latch latch_5132(eclk,ereset, cp1_v, n_533_v, n_599_v);
  spice_latch latch_5133(eclk,ereset, cp1_v, n_920_v, n_785_v);
  spice_latch latch_5134(eclk,ereset, cclk_v, VEC1_v, n_1452_v);
  spice_latch latch_5135(eclk,ereset, cclk_v, n_896_v, notidl3_v);
  spice_latch latch_5138(eclk,ereset, cclk_v, n_1187_v, nots6_v);
  spice_latch latch_5109(eclk,ereset, cclk_v, v(n_722_v), notalu6_v);
  spice_latch latch_5107(eclk,ereset, cp1_v, n_566_v, p1_v);
  spice_latch latch_5106(eclk,ereset, cp1_v, notRnWprepad_v, n_1579_v);
  spice_latch latch_5045(eclk,ereset, cp1_v, n_1215_v, n_223_v);
  spice_latch latch_5047(eclk,ereset, cp1_v, n_931_v, n_1674_v);
  spice_latch latch_4972(eclk,ereset, cclk_v, n_862_v, pipeUNK11_v);
  spice_latch latch_5088(eclk,ereset, cp1_v, n_1497_v, n_653_v);
  spice_latch latch_5089(eclk,ereset, cclk_v, n_616_v, n_460_v);
  spice_latch latch_5084(eclk,ereset, cclk_v, n_1281_v, pd3_v);
  spice_latch latch_5085(eclk,ereset, cclk_v, n_1588_v, pd5_v);
  spice_latch latch_5086(eclk,ereset, cclk_v, n_1075_v, pd4_v);
  spice_latch latch_5087(eclk,ereset, cclk_v, n_1638_v, notidl6_v);
  spice_latch latch_5080(eclk,ereset, cclk_v, v(notaluoutmux0_v), notalu0_v);
  spice_latch latch_5081(eclk,ereset, cclk_v, v(n_296_v), notalu4_v);
  spice_latch latch_5082(eclk,ereset, cclk_v, n_340_v, pipeUNK12_v);
  spice_latch latch_5083(eclk,ereset, cp1_v, notRnWprepad_v, n_759_v);
  spice_latch latch_5136(eclk,ereset, cp1_v, n_720_v, n_1338_v);
  spice_latch latch_5137(eclk,ereset, cclk_v, n_1229_v, pchp0_v);
  spice_latch latch_5139(eclk,ereset, cp1_v, n_1082_v, p0_v);
  spice_latch latch_5054(eclk,ereset, cp1_v, n_1376_v, notdor2_v);
  spice_latch latch_4959(eclk,ereset, cclk_v, n_1194_v, pipeUNK04_v);
  spice_latch latch_4958(eclk,ereset, cclk_v, n_1106_v, n_1404_v);
  spice_latch latch_4955(eclk,ereset, cp1_v, n_1275_v, n_1581_v);
  spice_latch latch_4954(eclk,ereset, cclk_v, n_718_v, notidl0_v);
  spice_latch latch_4957(eclk,ereset, cclk_v, n_1391_v, pipeUNK15_v);
  spice_latch latch_4956(eclk,ereset, cp1_v, D1x1_v, n_1472_v);
  spice_latch latch_4951(eclk,ereset, cclk_v, n_548_v, nots7_v);
  spice_latch latch_4950(eclk,ereset, cclk_v, n_695_v, n_1341_v);
  spice_latch latch_4953(eclk,ereset, cclk_v, v(n_740_v), notalu2_v);
  spice_latch latch_4952(eclk,ereset, cclk_v, n_795_v, n_360_v);
  spice_latch latch_4977(eclk,ereset, cclk_v, n_182_v, n_265_v);
  spice_latch latch_4976(eclk,ereset, cp1_v, notRdy0_v, n_902_v);
  spice_latch latch_4975(eclk,ereset, cp1_v, n_789_v, notdor7_v);
  spice_latch latch_4974(eclk,ereset, cclk_v, n_213_v, notidl1_v);
  spice_latch latch_4971(eclk,ereset, cp1_v, n_299_v, n_1625_v);
  spice_latch latch_4970(eclk,ereset, cp1_v, n_1687_v, notdor0_v);
  spice_latch latch_5022(eclk,ereset, cp1_v, n_845_v, p2_v);
  spice_latch latch_5023(eclk,ereset, cclk_v, n_318_v, pipeUNK14_v);
  spice_latch latch_5020(eclk,ereset, cclk_v, notaluvout_v, n_408_v);
  spice_latch latch_5021(eclk,ereset, cclk_v, n_462_v, n_878_v);
  spice_latch latch_5026(eclk,ereset, cclk_v, C78_v, C78_phi2_v);
  spice_latch latch_5027(eclk,ereset, cclk_v, n_1090_v, n_1683_v);
  spice_latch latch_5024(eclk,ereset, cclk_v, n_188_v, pipeT4out_v);
  spice_latch latch_5025(eclk,ereset, cp1_v, n_1087_v, n_1132_v);
  spice_latch latch_5028(eclk,ereset, cclk_v, n_586_v, pipeBRtaken_v);
  spice_latch latch_5029(eclk,ereset, cclk_v, n_983_v, nots0_v);
  spice_latch latch_5123(eclk,ereset, cclk_v, n_1175_v, pipeUNK28_v);
  spice_latch latch_5122(eclk,ereset, cclk_v, n_1085_v, pipeUNK23_v);
  spice_latch latch_5129(eclk,ereset, cclk_v, n_484_v, pclp7_v);
  spice_latch latch_5128(eclk,ereset, cp1_v, n_916_v, n_1409_v);
  spice_latch latch_5004(eclk,ereset, cclk_v, _WR_v, pipe_WR_phi2_v);
  spice_latch latch_5005(eclk,ereset, cp1_v, n_1375_v, n_95_v);
  spice_latch latch_5006(eclk,ereset, cp1_v, n_1089_v, n_1529_v);
  spice_latch latch_5007(eclk,ereset, cclk_v, n_1631_v, pclp3_v);
  spice_latch latch_5000(eclk,ereset, cclk_v, n_875_v, n_469_v);
  spice_latch latch_5001(eclk,ereset, cp1_v, n_913_v, n_1274_v);
  spice_latch latch_5002(eclk,ereset, cclk_v, n_1688_v, n_680_v);
  spice_latch latch_5003(eclk,ereset, cclk_v, VEC0_v, n_1126_v);
  spice_latch latch_5008(eclk,ereset, cp1_v, brk_done_v, n_1291_v);
  spice_latch latch_5009(eclk,ereset, cp1_v, n_428_v, n_644_v);
  spice_latch latch_5068(eclk,ereset, cclk_v, n_1705_v, n_1020_v);
  spice_latch latch_5069(eclk,ereset, cclk_v, n_944_v, pipeUNK37_v);
  spice_latch latch_5066(eclk,ereset, cp1_v, INTG_v, n_50_v);
  spice_latch latch_5067(eclk,ereset, cclk_v, n_396_v, n_796_v);
  spice_latch latch_5064(eclk,ereset, cclk_v, op_ORS_v, n_88_v);
  spice_latch latch_5065(eclk,ereset, cclk_v, n_629_v, n_760_v);
  spice_latch latch_5062(eclk,ereset, cclk_v, n_515_v, n_1411_v);
  spice_latch latch_5063(eclk,ereset, cclk_v, n_1211_v, n_897_v);
  spice_latch latch_5060(eclk,ereset, cclk_v, n_504_v, pipeUNK41_v);
  spice_latch latch_5061(eclk,ereset, cclk_v, op_ANDS_v, n_1574_v);
  spice_latch latch_5071(eclk,ereset, cclk_v, n_17_v, pipe_T0_v);
  spice_latch latch_5040(eclk,ereset, cclk_v, n_62_v, pd7_v);
  spice_latch latch_5041(eclk,ereset, cp1_v, n_1290_v, n_698_v);
  spice_latch latch_5042(eclk,ereset, cclk_v, n_374_v, pd6_v);
  spice_latch latch_5043(eclk,ereset, cp1_v, n_1718_v, n_671_v);
  spice_latch latch_5044(eclk,ereset, cp1_v, notRdy0_v, n_1679_v);
  spice_latch latch_5046(eclk,ereset, cclk_v, n_440_v, pipeUNK39_v);
  spice_latch latch_5048(eclk,ereset, cp1_v, n_1526_v, n_1450_v);
  spice_latch latch_5049(eclk,ereset, cclk_v, n_604_v, n_1477_v);
  spice_latch latch_5118(eclk,ereset, cclk_v, n_80_v, n_1333_v);
  spice_latch latch_4973(eclk,ereset, cclk_v, n_862_v, pipeT_SYNC_v);
  spice_latch latch_4979(eclk,ereset, cclk_v, op_T__bit_v, n_1673_v);
  spice_latch latch_4978(eclk,ereset, cclk_v, n_490_v, notidl4_v);
  spice_latch latch_5141(eclk,ereset, cclk_v, n_844_v, n_459_v);
  spice_latch latch_5140(eclk,ereset, cclk_v, n_1486_v, n_126_v);
  spice_latch latch_5143(eclk,ereset, cclk_v, n_1575_v, pipeT2out_v);
  spice_latch latch_5142(eclk,ereset, cclk_v, n_474_v, n_15_v);
  spice_latch latch_5145(eclk,ereset, cp1_v, n_1339_v, n_597_v);
  spice_latch latch_5144(eclk,ereset, cclk_v, n_973_v, nots4_v);
  spice_latch latch_5149(eclk,ereset, cclk_v, n_29_v, pipeUNK22_v);
  spice_latch latch_5157(eclk,ereset, cp1_v, n_1650_v, n_94_v);
  spice_latch latch_4989(eclk,ereset, cp1_v, n_1178_v, n_590_v);
  spice_latch latch_4980(eclk,ereset, cclk_v, n_513_v, pipeUNK06_v);
  spice_latch latch_4981(eclk,ereset, cp1_v, v(n_854_v), n_1395_v);
  spice_latch latch_4986(eclk,ereset, cclk_v, nnT2BR_v, n_1269_v);
  spice_latch latch_4984(eclk,ereset, cclk_v, n_20_v, n_993_v);
  spice_latch latch_4985(eclk,ereset, cclk_v, n_1101_v, n_190_v);
  spice_latch latch_5169(eclk,ereset, cclk_v, n_588_v, notidl7_v);
  spice_latch latch_5168(eclk,ereset, cp1_v, n_1180_v, n_1533_v);
  spice_latch latch_5163(eclk,ereset, cclk_v, n_958_v, n_865_v);
  spice_latch latch_5162(eclk,ereset, cclk_v, n_889_v, pipeUNK42_v);
  spice_latch latch_5161(eclk,ereset, cclk_v, n_90_v, pipeUNK05_v);
  spice_latch latch_5160(eclk,ereset, cp1_v, n_472_v, n_1606_v);
  spice_latch latch_5167(eclk,ereset, cclk_v, n_1455_v, n_1505_v);
  spice_latch latch_5166(eclk,ereset, cclk_v, n_1037_v, n_266_v);
  spice_latch latch_5165(eclk,ereset, cclk_v, n_1649_v, n_1027_v);
  spice_latch latch_5164(eclk,ereset, cclk_v, Reset0_v, pipephi2Reset0_v);
  spice_latch latch_5105(eclk,ereset, cclk_v, _op_set_C_v, pipeUNK08_v);
  spice_latch latch_5104(eclk,ereset, cclk_v, n_678_v, pipeT3out_v);
  spice_latch latch_5101(eclk,ereset, cclk_v, n_1225_v, n_1121_v);
  spice_latch latch_5100(eclk,ereset, cclk_v, n_1402_v, pchp2_v);
  spice_latch latch_5103(eclk,ereset, cclk_v, n_1024_v, n_1699_v);
  spice_latch latch_5102(eclk,ereset, cclk_v, v(n_277_v), notalu5_v);
  spice_latch latch_5152(eclk,ereset, cclk_v, x_op_T__adc_sbc_v, pipeUNK03_v);
  spice_latch latch_5153(eclk,ereset, cclk_v, DC78_v, DC78_phi2_v);
  spice_latch latch_5150(eclk,ereset, cclk_v, n_14_v, pipeUNK20_v);
  spice_latch latch_5151(eclk,ereset, cclk_v, n_696_v, n_610_v);
  spice_latch latch_5154(eclk,ereset, cclk_v, n_207_v, n_1061_v);
  spice_latch latch_5155(eclk,ereset, cclk_v, n_31_v, pipeUNK16_v);
  spice_latch latch_5127(eclk,ereset, cclk_v, n_1319_v, pd1_v);
  spice_latch latch_5126(eclk,ereset, cclk_v, n_93_v, pd0_v);
  spice_latch latch_5125(eclk,ereset, cclk_v, op_SRS_v, pipeUNK27_v);
  spice_latch latch_5124(eclk,ereset, cclk_v, n_160_v, n_1049_v);
  spice_latch latch_5121(eclk,ereset, cclk_v, n_378_v, pipeT5out_v);
  spice_latch latch_5120(eclk,ereset, cp1_v, n_1215_v, n_1528_v);
  spice_latch latch_5146(eclk,ereset, cp1_v, notRnWprepad_v, n_402_v);
  spice_latch latch_5148(eclk,ereset, cclk_v, n_1717_v, n_1113_v);
  spice_latch latch_5093(eclk,ereset, cclk_v, n_1069_v, n_1177_v);
  spice_latch latch_5092(eclk,ereset, cclk_v, n_1045_v, pipeUNK13_v);
  spice_latch latch_5091(eclk,ereset, cclk_v, n_728_v, pipeVectorA0_v);
  spice_latch latch_5090(eclk,ereset, cp1_v, n_109_v, n_1161_v);
  spice_latch latch_5097(eclk,ereset, cclk_v, n_1711_v, nots1_v);
  spice_latch latch_5096(eclk,ereset, cclk_v, n_1586_v, n_621_v);
  spice_latch latch_5095(eclk,ereset, cclk_v, n_1225_v, pipedpc28_v);
  spice_latch latch_5094(eclk,ereset, cclk_v, Reset0_v, pipephi2Reset0x_v);
  spice_latch latch_5099(eclk,ereset, cclk_v, n_1073_v, pclp5_v);
  spice_latch latch_5098(eclk,ereset, cclk_v, n_1358_v, n_521_v);
  spice_latch latch_4948(eclk,ereset, cp1_v, n_645_v, n_562_v);
  spice_latch latch_4949(eclk,ereset, cp1_v, n_262_v, n_1447_v);
  spice_latch latch_4947(eclk,ereset, cclk_v, n_11_v, n_55_v);
  spice_latch latch_4960(eclk,ereset, cclk_v, n_385_v, pipeUNK30_v);
  spice_latch latch_4961(eclk,ereset, cclk_v, n_442_v, n_509_v);
  spice_latch latch_4962(eclk,ereset, cp1_v, n_1368_v, n_1149_v);
  spice_latch latch_4963(eclk,ereset, cclk_v, n_1179_v, n_393_v);
  spice_latch latch_4964(eclk,ereset, cp1_v, n_430_v, n_1570_v);
  spice_latch latch_4965(eclk,ereset, cclk_v, _VEC_v, pipe_VEC_v);
  spice_latch latch_4966(eclk,ereset, cclk_v, n_261_v, pipeUNK36_v);
  spice_latch latch_4967(eclk,ereset, cp1_v, n_959_v, n_323_v);
  spice_latch latch_4968(eclk,ereset, cclk_v, n_176_v, n_598_v);
  spice_latch latch_4969(eclk,ereset, cclk_v, n_169_v, pipeUNK29_v);
  spice_latch latch_5031(eclk,ereset, cp1_v, n_1495_v, p3_v);
  spice_latch latch_5030(eclk,ereset, cclk_v, n_272_v, n_1162_v);
  spice_latch latch_5033(eclk,ereset, cclk_v, n_1500_v, n_526_v);
  spice_latch latch_5032(eclk,ereset, cclk_v, n_191_v, pipeUNK40_v);
  spice_latch latch_5035(eclk,ereset, cclk_v, n_264_v, n_1693_v);
  spice_latch latch_5034(eclk,ereset, cclk_v, n_264_v, n_799_v);
  spice_latch latch_5037(eclk,ereset, cclk_v, n_824_v, n_398_v);
  spice_latch latch_5036(eclk,ereset, cclk_v, n_334_v, pipeUNK17_v);
  spice_latch latch_5039(eclk,ereset, cclk_v, n_111_v, pd2_v);
  spice_latch latch_5038(eclk,ereset, cclk_v, n_1065_v, n_1124_v);
  spice_latch latch_5019(eclk,ereset, cclk_v, n_779_v, n_805_v);
  spice_latch latch_5018(eclk,ereset, cp1_v, n_1141_v, n_101_v);
  spice_latch latch_5013(eclk,ereset, cclk_v, n_1374_v, n_1252_v);
  spice_latch latch_5012(eclk,ereset, cclk_v, n_1347_v, n_1527_v);
  spice_latch latch_5011(eclk,ereset, cp1_v, n_1380_v, n_666_v);
  spice_latch latch_5010(eclk,ereset, cp1_v, n_1474_v, notdor1_v);
  spice_latch latch_5017(eclk,ereset, cclk_v, n_132_v, pipeUNK26_v);
  spice_latch latch_5016(eclk,ereset, cclk_v, n_1209_v, n_663_v);
  spice_latch latch_5015(eclk,ereset, cp1_v, n_1181_v, n_69_v);
  spice_latch latch_5014(eclk,ereset, cclk_v, n_1594_v, n_688_v);
  spice_latch latch_4982(eclk,ereset, cp1_v, n_468_v, n_18_v);
  spice_latch latch_4983(eclk,ereset, cp1_v, n_1039_v, n_24_v);
  spice_latch latch_4987(eclk,ereset, cclk_v, n_327_v, pipeUNK09_v);
  spice_latch latch_5079(eclk,ereset, cclk_v, v(n_1071_v), notalu3_v);
  spice_latch latch_5078(eclk,ereset, cclk_v, n_473_v, pipeUNK33_v);
  spice_latch latch_5075(eclk,ereset, cclk_v, n_1199_v, notidl2_v);
  spice_latch latch_5074(eclk,ereset, cclk_v, n_1081_v, pipeUNK32_v);
  spice_latch latch_5077(eclk,ereset, cclk_v, n_389_v, pipeUNK31_v);
  spice_latch latch_5076(eclk,ereset, cclk_v, n_824_v, pipeUNK34_v);
  spice_latch latch_5070(eclk,ereset, cp1_v, n_1684_v, notdor6_v);
  spice_latch latch_5073(eclk,ereset, cclk_v, v(notaluoutmux1_v), notalu1_v);
  spice_latch latch_5072(eclk,ereset, cp1_v, _TWOCYCLE_v, _TWOCYCLE_phi1_v);
  spice_latch latch_5108(eclk,ereset, cclk_v, n_306_v, n_581_v);
  spice_latch latch_5057(eclk,ereset, cp1_v, n_797_v, notdor4_v);
  spice_latch latch_5056(eclk,ereset, cclk_v, n_1117_v, pipeVectorA1_v);
  spice_latch latch_5055(eclk,ereset, cclk_v, n_34_v, nots3_v);
  spice_latch latch_5053(eclk,ereset, cclk_v, n_952_v, n_1509_v);
  spice_latch latch_5052(eclk,ereset, cp1_v, n_961_v, notdor5_v);
  spice_latch latch_5051(eclk,ereset, cp1_v, notRdy0_v, n_1276_v);
  spice_latch latch_5050(eclk,ereset, cclk_v, n_501_v, pipeUNK35_v);
  spice_latch latch_5059(eclk,ereset, cp1_v, n_1091_v, n_1360_v);
  spice_latch latch_5058(eclk,ereset, cclk_v, n_700_v, n_1565_v);
  spice_latch latch_5156(eclk,ereset, cclk_v, n_506_v, n_1602_v);
  spice_latch latch_5158(eclk,ereset, cp1_v, notRdy0_v, n_1272_v);
  spice_latch latch_5159(eclk,ereset, cp1_v, n_1093_v, n_226_v);
  spice_latch latch_5147(eclk,ereset, cclk_v, n_568_v, notidl5_v);
  spice_latch latch_5119(eclk,ereset, cclk_v, n_1657_v, pchp4_v);
  spice_latch latch_5112(eclk,ereset, cp1_v, n_626_v, n_756_v);
  spice_latch latch_5113(eclk,ereset, cclk_v, n_104_v, n_1221_v);
  spice_latch latch_5170(eclk,ereset, cp1_v, notRdy0_v, n_1624_v);
  spice_latch latch_5171(eclk,ereset, cp1_v, v(n_330_v), n_675_v);
  spice_latch latch_5172(eclk,ereset, cclk_v, n_1712_v, pipeVectorA2_v);
  spice_latch latch_5173(eclk,ereset, cclk_v, n_496_v, nots5_v);
  spice_latch latch_4999(eclk,ereset, cclk_v, op_SUMS_v, n_415_v);
  spice_latch latch_4998(eclk,ereset, cclk_v, op_SRS_v, n_968_v);
  spice_latch latch_4991(eclk,ereset, cclk_v, n_632_v, n_339_v);
  spice_latch latch_4990(eclk,ereset, cclk_v, n_1192_v, pchp6_v);
  spice_latch latch_4993(eclk,ereset, cclk_v, n_1379_v, pipeUNK07_v);
  spice_latch latch_4992(eclk,ereset, cclk_v, n_1190_v, nots2_v);
  spice_latch latch_4995(eclk,ereset, cclk_v, n_1130_v, n_512_v);
  spice_latch latch_4994(eclk,ereset, cclk_v, n_1099_v, pclp1_v);
  spice_latch latch_4997(eclk,ereset, cclk_v, n_774_v, pipeUNK02_v);
  spice_latch latch_4996(eclk,ereset, cclk_v, n_674_v, n_745_v);
  spice_latch latch_5116(eclk,ereset, cclk_v, n_19_v, pipeUNK18_v);
  spice_latch latch_5117(eclk,ereset, cclk_v, v(n_304_v), notalu7_v);
  spice_latch latch_5114(eclk,ereset, cp1_v, n_420_v, n_47_v);
  spice_latch latch_5115(eclk,ereset, cclk_v, n_1231_v, pipeUNK21_v);
  spice_latch latch_5110(eclk,ereset, cclk_v, n_608_v, n_559_v);
  spice_latch latch_5111(eclk,ereset, cp1_v, n_457_v, notdor3_v);

  assign n_951_v = ~(abl2_v);
  assign op_T__cpx_cpy_abs_v = ~((notir3_v|ir4_v|irline3_v|notir6_v|notir2_v|clock2_v|notir7_v));
  assign n_1219_v = ~(op_T5_jsr_v);
  assign AxB5_v = ~((n_1632_v|n_647_v));
  assign n_1222_v = ~(n_1225_v);
  assign n_1694_v = ~(n_890_v);
  assign n_1691_v = ~((alub2_v|alua2_v));
  assign dpc34_PCLC_v = ~((n_641_v|n_783_v|n_937_v|n_329_v|n_386_v|n_1643_v|n_232_v|dpc36_IPC_v|n_249_v));
  assign C12_v = ~(_C12_v);
  assign n_506_v = ~((n_236_v|n_192_v));
  assign n_578_v = ~(n_1017_v);
  assign n_565_v = ~(y4_v);
  assign n_1209_v = ~((n_1213_v|(n_609_v&n_453_v)));
  assign op_T2_ind_y_v = ~((_t2_v|notir0_v|notir4_v|ir3_v|ir2_v));
  assign n_141_v = ~(pchp3_v);
  assign C45_v = ~(((n_1063_v&_C34_v)|n_404_v));
  assign op_T5_ind_x_v = ~((ir3_v|ir4_v|notir0_v|_t5_v|ir2_v));
  assign n_1211_v = ~((n_1286_v|n_862_v|op_T2_abs_access_v|nnT2BR_v|n_1002_v));
  assign n_1457_v = ~((n_781_v|n_1492_v));
  assign n_1441_v = ~(n_1277_v);
  assign Pout1_v = ~(n_318_v);
  assign n_1446_v = ~((n_850_v|n_771_v));
  assign n_755_v = ~(pipeUNK06_v);
  assign dor5_v = ~(notdor5_v);
  assign n_1455_v = ~((op_T__ora_and_eor_adc_v|op_T__shift_a_v|op_T0_tya_v|op_T0_pla_v|op_T0_txa_v|op_T0_lda_v|op_T__adc_sbc_v));
  assign n_761_v = ~(alu5_v);
  assign n_1347_v = ~((n_782_v|op_T0_shift_a_v|n_550_v|n_862_v|nnT2BR_v|n_979_v));
  assign n_1344_v = ~(n_556_v);
  assign n_1345_v = ~((n_937_v|dpc36_IPC_v));
  assign op_T0_acc_v = ~((notir0_v|clock1_v));
  assign n_1343_v = ~((n_152_v|notRdy0_v));
  assign n_1433_v = ~((_op_branch_bit6_v|n_201_v|n_90_v));
  assign abl5_v = ~(_ABL5_v);
  assign n_231_v = ~(PD_xxxx10x0_v);
  assign n_227_v = ~(pd4_clearIR_v);
  assign n_233_v = ~((n_761_v&n_149_v));
  assign dpc28_0ADH0_v = ~(pipedpc28_v);
  assign n_225_v = ~(n_1223_v);
  assign _DA_ADD1_v = ~(alu1_v);
  assign op_T2_zp_zp_idx_v = ~((ir3_v|notir2_v|_t2_v));
  assign n_284_v = ~(n_1392_v);
  assign n_1717_v = ~(((op_T2_idx_x_xy_v&op_xy_v)|(x_op_T0_tya_v|op_T2_abs_y_v|op_T0_cpy_iny_v|op_T3_ind_y_v|op_T0_iny_dey_v)|(n_335_v&op_sty_cpy_mem_v)));
  assign n_1709_v = ~(n_1434_v);
  assign op_T__cpx_cpy_imm_zp_v = ~((irline3_v|notir7_v|clock2_v|notir6_v|ir3_v|ir4_v));
  assign n_1711_v = ~(s1_v);
  assign n_1719_v = ~(a5_v);
  assign n_1714_v = ~(pipeUNK26_v);
  assign n_1715_v = ~(n_358_v);
  assign n_1716_v = ~((n_510_v|op_T3_branch_v|n_1258_v|n_218_v));
  assign n_1712_v = ~((C1x5Reset_v|_VEC_v|n_264_v));
  assign op_T0_jmp_v = ~((clock1_v|notir3_v|notir2_v|notir6_v|ir7_v|ir4_v|irline3_v));
  assign n_928_v = ~(pd5_clearIR_v);
  assign n_930_v = ~((n_134_v|n_1276_v));
  assign n_929_v = ~(n_1549_v);
  assign n_327_v = ~((x_op_T4_rti_v|op_T0_plp_v));
  assign n_931_v = ~(n_415_v);
  assign op_inc_nop_v = ~((notir1_v|notir7_v|notir5_v|notir6_v));
  assign n_329_v = ~(pcl1_v);
  assign n_326_v = ~(n_1356_v);
  assign n_709_v = ~(n_1499_v);
  assign op_T2_jsr_v = ~((ir3_v|ir4_v|ir2_v|notir5_v|irline3_v|_t2_v|ir6_v|ir7_v));
  assign abh1_v = ~(v(_ABH1_v));
  assign n_714_v = ~(n_906_v);
  assign n_700_v = ~(dpc18__DAA_v);
  assign __AxB_2_v = ~((n_681_v&n_110_v));
  assign notir1_v = ~(ir1_v);
  assign n_708_v = ~(n_1230_v);
  assign n_715_v = ~(n_641_v);
  assign n_717_v = ~((n_1132_v|pipephi2Reset0x_v));
  assign op_T2_ADL_ADD_v = ~((_t2_v|ir3_v));
  assign n_206_v = ~(alucout_v);
  assign n_213_v = ~(v(db1_v));
  assign n_209_v = ~(pchp1_v);
  assign n_637_v = ~((n_1318_v|C67_v));
  assign n_638_v = ~(op_T0_v);
  assign n_632_v = ~((op_T2_stack_v|(op_T0_jsr_v&n_1289_v)));
  assign n_636_v = ~(op_T2_branch_v);
  assign n_624_v = ~(v(idb0_v));
  assign DA_C01_v = ~((aluanorb0_v|(notalucin_v&aluanandb0_v)));
  assign n_254_v = ~(v(adh5_v));
  assign n_261_v = ~((x_op_T3_abs_idx_v|x_op_T4_ind_y_v));
  assign n_256_v = ~((op_T5_rti_v|op_T3_v|op_T5_rts_v|op_T5_ind_x_v|op_T0_jmp_v|op_T4_v|op_T0_brk_rti_v));
  assign n_255_v = ~(n_611_v);
  assign n_488_v = ~(pclp0_v);
  assign op_T0_tya_v = ~((ir5_v|ir2_v|notir7_v|clock1_v|ir6_v|notir4_v|irline3_v|notir3_v));
  assign n_478_v = ~(v(idb4_v));
  assign abh7_v = ~(v(_ABH7_v));
  assign n_479_v = ~((n_61_v|n_739_v));
  assign n_953_v = ~(AxB1_v);
  assign n_954_v = ~(pipeUNK08_v);
  assign n_956_v = ~(n_476_v);
  assign n_959_v = ~((pipeUNK20_v|n_430_v));
  assign n_961_v = ~(v(idb5_v));
  assign n_992_v = ~(n_595_v);
  assign n_986_v = ~((_DA_ADD2_v&_DA_ADD1_v));
  assign n_990_v = ~(abl3_v);
  assign n_988_v = ~(n_350_v);
  assign irline3_v = ~(n_1133_v);
  assign op_T0_ldx_tax_tsx_v = ~((notir5_v|notir1_v|ir6_v|clock1_v|notir7_v));
  assign n_983_v = ~(s0_v);
  assign n_987_v = ~(x0_v);
  assign n_1069_v = ~((n_1024_v|n_1274_v));
  assign n_1070_v = ~(pch1_v);
  assign n_1368_v = ~((n_645_v|n_1578_v|n_1374_v));
  assign n_1364_v = ~(n_101_v);
  assign n_1358_v = ~((n_1109_v|n_917_v|op_T0_txs_v));
  assign n_1357_v = ~(n_223_v);
  assign DC34_v = ~((dpc18__DAA_v|((n_319_v|n_1691_v)&(n_388_v|n_1610_v))));
  assign n_1371_v = ~((n_1045_v|n_201_v|n_846_v));
  assign p7_v = ~(n_1045_v);
  assign n_1369_v = ~(n_897_v);
  assign pd3_clearIR_v = ~((pd3_v|clearIR_v));
  assign n_1586_v = ~(op_T0_tsx_v);
  assign n_1588_v = ~(v(db5_v));
  assign n_845_v = ~(((n_1573_v&n_781_v)|(pipeUNK17_v&n_553_v)|(n_270_v&n_1662_v)));
  assign n_846_v = ~(_op_branch_bit6_v);
  assign n_838_v = ~(n_581_v);
  assign n_839_v = ~(cp1_v);
  assign n_834_v = ~(n_402_v);
  assign n_1585_v = ~(cclk_v);
  assign op_T2_stack_v = ~((ir7_v|ir2_v|irline3_v|_t2_v|ir4_v));
  assign n_228_v = ~(n_21_v);
  assign alu0_v = ~(notalu0_v);
  assign op_T0_ora_v = ~((ir6_v|notir0_v|clock1_v|ir5_v|ir7_v));
  assign op_T0_tsx_v = ~((ir6_v|notir4_v|notir5_v|ir2_v|clock1_v|notir1_v|notir7_v|notir3_v));
  assign n_0_ADL1_v = ~(pipeVectorA1_v);
  assign __AxB3__C23_v = ~((AxB3_v|_C23_v));
  assign n_1265_v = ~(pch2_v);
  assign n_1267_v = ~(v(adh1_v));
  assign n_1260_v = ~(n_598_v);
  assign n_1262_v = ~(n_1679_v);
  assign n_1258_v = ~(n_390_v);
  assign n_1256_v = ~(n_91_v);
  assign n_1257_v = ~((notalucout_v|n_1218_v));
  assign n_1253_v = ~((n_1542_v|n_783_v));
  assign n_1413_v = ~(n_1260_v);
  assign n_1412_v = ~(n_1455_v);
  assign Pout2_v = ~(n_334_v);
  assign op_T0_lda_v = ~((clock1_v|notir0_v|notir5_v|notir7_v|ir6_v));
  assign n_397_v = ~(op_T0_lda_v);
  assign n_104_v = ~((n_440_v|nnT2BR_v|n_275_v|op_T4_jmp_v|n_847_v));
  assign n_105_v = ~(notalucin_v);
  assign op_T2_ind_x_v = ~((ir2_v|_t2_v|ir3_v|notir0_v|ir4_v));
  assign pd7_clearIR_v = ~((pd7_v|clearIR_v));
  assign n_1408_v = ~((n_1044_v&(op_rol_ror_v|op_T0_adc_sbc_v)));
  assign n_595_v = ~((op_T4_abs_idx_v|op_T5_ind_y_v));
  assign n_583_v = ~(v(idb1_v));
  assign n_586_v = ~(((BRtaken_v&nnT2BR_v)|n_1619_v));
  assign op_T3_jsr_v = ~((irline3_v|ir6_v|notir5_v|ir3_v|ir2_v|ir7_v|_t3_v|ir4_v));
  assign n_582_v = ~(n_610_v);
  assign _C67_v = ~(C67_v);
  assign n_593_v = ~(n_355_v);
  assign n_587_v = ~(pipeUNK12_v);
  assign n_588_v = ~(v(db7_v));
  assign n_72_v = ~(pclp5_v);
  assign n_871_v = ~(n_1561_v);
  assign alu1_v = ~(notalu1_v);
  assign n_877_v = ~((n_933_v|n_506_v));
  assign n_1720_v = ~((RnWstretched_v|dor5_v));
  assign n_875_v = ~(((n_523_v&n_499_v)|n_743_v));
  assign n_876_v = ~(n_867_v);
  assign n_457_v = ~(v(idb3_v));
  assign n_453_v = ~(pch7_v);
  assign idl3_v = ~(notidl3_v);
  assign n_462_v = ~(n_1338_v);
  assign aluanorb1_v = ~((alua1_v|alub1_v));
  assign clock2_v = ~(n_1533_v);
  assign n_1205_v = ~(((n_1018_v&n_811_v)|(n_1257_v&n_233_v)));
  assign n_38_v = ~(cp1_v);
  assign alu5_v = ~(notalu5_v);
  assign n_973_v = ~(s4_v);
  assign n_320_v = ~(v(sb1_v));
  assign n_317_v = ~(n_445_v);
  assign _t3_v = ~(n_678_v);
  assign n_321_v = ~(n_398_v);
  assign n_23_v = ~((dor7_v|RnWstretched_v));
  assign n_1552_v = ~(n_1593_v);
  assign n_976_v = ~(pclp1_v);
  assign n_1055_v = ~((n_1708_v|n_771_v));
  assign n_1063_v = ~((alub4_v&alua4_v));
  assign n_1386_v = ~((n_715_v&n_1316_v));
  assign op_T5_mem_ind_idx_v = ~((ir3_v|_t5_v|ir2_v|notir0_v));
  assign n_1380_v = ~((n_819_v|n_1154_v));
  assign n_1379_v = ~(x_op_T0_bit_v);
  assign n_1065_v = ~(op_T0_cli_sei_v);
  assign n_1464_v = ~((op_T5_brk_v|op_T5_rti_v|op_T0_php_pha_v|op_T4_rts_v|op_T3_plp_pla_v|op_T0_jsr_v));
  assign n_1491_v = ~(n_1484_v);
  assign n_385_v = ~((n_604_v|n_1377_v));
  assign n_1449_v = ~(n_958_v);
  assign n_754_v = ~((n_1673_v|(pipeUNK09_v&pipeUNK06_v)));
  assign n_551_v = ~(n_393_v);
  assign n_550_v = ~((op_ANDS_v|n_384_v));
  assign ir1_v = ~(n_119_v);
  assign op_T0_eor_v = ~((notir0_v|ir5_v|clock1_v|notir6_v|ir7_v));
  assign n_544_v = ~(op_ror_v);
  assign n_543_v = ~(n_339_v);
  assign n_553_v = ~((n_781_v|n_1662_v));
  assign op_T0_php_pha_v = ~((ir4_v|ir7_v|notir3_v|clock1_v|ir2_v|ir5_v|irline3_v));
  assign n_548_v = ~(s7_v);
  assign op_shift_v = ~((ir7_v|ir6_v|notir1_v));
  assign n_1423_v = ~(abh5_v);
  assign n_1427_v = ~((nnT2BR_v|n_236_v));
  assign n_1542_v = ~((n_1166_v&n_1345_v));
  assign x_op_T0_txa_v = ~((notir7_v|ir4_v|notir3_v|ir5_v|ir2_v|notir1_v|clock1_v|ir6_v));
  assign n_811_v = ~((n_838_v|alucout_v));
  assign n_1541_v = ~((n_1477_v|n_43_v));
  assign C78_v = ~(_C78_v);
  assign n_812_v = ~((n_440_v|n_646_v));
  assign n_810_v = ~((n_923_v|n_293_v));
  assign pd1_clearIR_v = ~((pd1_v|clearIR_v));
  assign BRtaken_v = ~(((n_270_v&n_620_v)|n_1115_v));
  assign n_1526_v = ~(n_680_v);
  assign n_212_v = ~(v(adh4_v));
  assign n_689_v = ~(op_T5_brk_v);
  assign Pout0_v = ~(n_31_v);
  assign op_asl_rol_v = ~((ir6_v|notir1_v|ir7_v));
  assign _t4_v = ~(n_188_v);
  assign aluaorb0_v = ~(aluanorb0_v);
  assign n_692_v = ~((n_43_v|n_460_v));
  assign n_695_v = ~((C34_v&n_700_v));
  assign n_694_v = ~(nots1_v);
  assign n_1722_v = ~(pchp0_v);
  assign n_1724_v = ~(n_730_v);
  assign op_T3_mem_abs_v = ~((_t3_v|ir4_v|notir2_v|notir3_v));
  assign op_branch_done_v = ~((n_603_v|irline3_v|notir4_v|ir2_v|clock1_v|ir3_v));
  assign n_609_v = ~((n_743_v&n_1488_v));
  assign op_T3_ind_y_v = ~((ir2_v|_t3_v|ir3_v|notir0_v|notir4_v));
  assign n_602_v = ~(n_133_v);
  assign n_608_v = ~(n_1272_v);
  assign n_604_v = ~(((op_T2_ADL_ADD_v&n_638_v)|(op_T4_rti_v|op_T4_brk_jsr_v|op_T3_ind_x_v|op_T2_stack_v|notRdy0_v|op_T3_stack_bit_jmp_v)));
  assign pclp4_v = ~(n_15_v);
  assign n_1521_v = ~(x3_v);
  assign _WR_v = ~((op_T2_php_pha_v|n_1258_v|op_T4_brk_v|n_440_v|n_335_v|n_1642_v));
  assign n_1346_v = ~(abh3_v);
  assign n_35_v = ~((n_43_v|n_796_v));
  assign pchp5_v = ~(n_469_v);
  assign op_T__dex_v = ~((notir7_v|ir4_v|notir3_v|clock2_v|ir5_v|notir6_v|ir2_v|notir1_v));
  assign op_T5_rti_v = ~((notir6_v|ir4_v|ir3_v|ir7_v|ir2_v|irline3_v|_t5_v|ir5_v));
  assign op_T2_v = ~(_t2_v);
  assign op_T0_sbc_v = ~((clock1_v|notir5_v|notir6_v|notir7_v|notir0_v));
  assign n_790_v = ~((op_asl_rol_v|op_lsr_ror_dec_inc_v));
  assign n_789_v = ~(v(idb7_v));
  assign n_795_v = ~(n_1649_v);
  assign op_push_pull_v = ~((notir3_v|irline3_v|ir2_v|ir7_v|ir4_v));
  assign _C45_v = ~(C45_v);
  assign n_1573_v = ~(v(idb2_v));
  assign op_T2_php_v = ~((irline3_v|ir6_v|ir4_v|ir5_v|ir7_v|_t2_v|ir2_v|notir3_v));
  assign n_1054_v = ~(C1x5Reset_v);
  assign op_T2_abs_v = ~((_t2_v|notir2_v|ir4_v|notir3_v));
  assign n_1056_v = ~(n_761_v);
  assign _op_branch_done_v = ~(op_branch_done_v);
  assign n_1275_v = ~((pipeBRtaken_v|notRdy0_v|ONEBYTE_v));
  assign C01_v = ~(((notalucin_v&aluanandb0_v)|aluanorb0_v));
  assign n_1281_v = ~(v(db3_v));
  assign n_1270_v = ~((n_43_v|n_509_v));
  assign _DBZ_v = ~(DBZ_v);
  assign op_T0_v = ~(clock1_v);
  assign n_1271_v = ~(n_1596_v);
  assign n_1657_v = ~(((n_83_v|dpc35_PCHC_v)&n_523_v));
  assign n_1286_v = ~((n_930_v|n_470_v));
  assign n_1277_v = ~(n_1020_v);
  assign n_198_v = ~(pipeUNK37_v);
  assign n_600_v = ~(n_1341_v);
  assign n_46_v = ~((n_992_v|notRdy0_v));
  assign n_1389_v = ~(nots2_v);
  assign n_1391_v = ~((op_T2_php_v|op_T4_brk_v));
  assign n_1401_v = ~(n_1269_v);
  assign n_1402_v = ~(((n_1202_v|n_200_v)&n_293_v));
  assign alu4_v = ~(notalu4_v);
  assign n_61_v = ~(v(sb6_v));
  assign op_lsr_ror_dec_inc_v = ~((notir6_v|notir1_v));
  assign op_T3_abs_idx_v = ~((_t3_v|notir3_v|notir4_v));
  assign n_494_v = ~(v(adh7_v));
  assign n_503_v = ~(notir5_v);
  assign n_504_v = ~((n_1120_v&n_440_v));
  assign n_264_v = ~((n_1149_v|n_1312_v));
  assign n_267_v = ~((n_1175_v|n_785_v|n_544_v));
  assign n_269_v = ~((AxB7_v|n_1038_v));
  assign n_270_v = ~(n_503_v);
  assign op_T0_jsr_v = ~((ir2_v|irline3_v|clock1_v|ir4_v|ir6_v|ir7_v|notir5_v|ir3_v));
  assign n_491_v = ~(n_1541_v);
  assign op_T4_ind_y_v = ~((_t4_v|ir2_v|notir0_v|notir4_v|ir3_v));
  assign n_773_v = ~((op_T2_abs_access_v|n_646_v));
  assign n_770_v = ~(n_559_v);
  assign abh5_v = ~(v(_ABH5_v));
  assign n_772_v = ~(n_1674_v);
  assign n_781_v = ~((pipeUNK09_v|notRdy0_v));
  assign _C12_v = ~(((C01_v&A_B1_v)|n_936_v));
  assign n_771_v = ~(n_1110_v);
  assign n_779_v = ~((n_1440_v&(n_1081_v|op_T0_sbc_v|n_1002_v)));
  assign notir3_v = ~(ir3_v);
  assign p4_v = ~(n_1471_v);
  assign n_1440_v = ~(notRdy0_v);
  assign n_1439_v = ~(y6_v);
  assign n_652_v = ~(pchp6_v);
  assign n_649_v = ~((alub3_v|alua3_v));
  assign pd5_clearIR_v = ~((pd5_v|clearIR_v));
  assign n_420_v = ~(n_865_v);
  assign n_885_v = ~(n_384_v);
  assign n_884_v = ~(AxB3_v);
  assign notir6_v = ~(ir6_v);
  assign n_889_v = ~(op_T0_clc_sec_v);
  assign n_888_v = ~(n_675_v);
  assign C67_v = ~(((_C56_v&n_336_v)|n_1084_v));
  assign A_B3_v = ~(n_649_v);
  assign n_1316_v = ~((n_232_v|n_344_v));
  assign n_1315_v = ~(abh0_v);
  assign abh6_v = ~(v(_ABH6_v));
  assign n_1660_v = ~(abl0_v);
  assign op_T__asl_rol_a_v = ~((ir4_v|ir6_v|ir2_v|notir3_v|notir1_v|clock2_v|ir7_v));
  assign op_T__inx_v = ~((notir5_v|notir6_v|ir2_v|clock2_v|notir7_v|ir4_v|notir3_v|irline3_v));
  assign n_1682_v = ~(_DA_ADD1_v);
  assign PD_xxx010x1_v = ~((n_409_v|n_1083_v|pd4_clearIR_v|pd2_clearIR_v));
  assign n_307_v = ~((n_31_v|_op_branch_bit7_v|n_846_v));
  assign n_306_v = ~(dpc22__DSA_v);
  assign n_1293_v = ~((n_318_v|_op_branch_bit6_v|_op_branch_bit7_v));
  assign PD_1xx000x0_v = ~((pd2_clearIR_v|pd3_clearIR_v|pd4_clearIR_v|pd0_clearIR_v|n_1605_v));
  assign n_1290_v = ~((n_1126_v|(VEC1_v&notRdy0_v)));
  assign n_571_v = ~(pd2_clearIR_v);
  assign n_572_v = ~(pipeUNK21_v);
  assign n_1596_v = ~(n_1602_v);
  assign idl0_v = ~(notidl0_v);
  assign op_sty_cpy_mem_v = ~((ir5_v|notir2_v|notir7_v|irline3_v|ir6_v));
  assign n_1605_v = ~(pd7_clearIR_v);
  assign n_1593_v = ~(n_226_v);
  assign n_1600_v = ~(v(idb3_v));
  assign n_1495_v = ~(((n_1457_v&pipeUNK04_v)|(n_1492_v&n_270_v)|(n_781_v&n_1600_v)));
  assign abl2_v = ~(_ABL2_v);
  assign n_409_v = ~(pd0_clearIR_v);
  assign n_404_v = ~((alub4_v|alua4_v));
  assign abh3_v = ~(v(_ABH3_v));
  assign n_419_v = ~(a2_v);
  assign AxB1_v = ~((n_936_v|aluanorb1_v));
  assign n_1496_v = ~(pchp2_v);
  assign n_1497_v = ~(pipeUNK41_v);
  assign dasb7_v = ~((n_260_v|(n_852_v&n_1205_v)));
  assign n_1649_v = ~((brk_done_v|notRdy0_v|n_389_v|op_T4_ind_x_v|op_jmp_v|op_T2_jsr_v|op_rti_rts_v|op_T2_abs_v|n_1109_v));
  assign n_1650_v = ~(v(so_v));
  assign n_1642_v = ~((n_462_v&n_824_v));
  assign n_1643_v = ~(pcl4_v);
  assign op_ORS_v = ~(n_1145_v);
  assign n_523_v = ~((dpc35_PCHC_v&n_83_v));
  assign n_538_v = ~(n_1599_v);
  assign pd4_clearIR_v = ~((clearIR_v|pd4_v));
  assign n_525_v = ~((cclk_v|n_266_v));
  assign xx_op_T5_jsr_v = ~((_t5_v|ir6_v|irline3_v|ir2_v|ir3_v|ir7_v|ir4_v|notir5_v));
  assign dor0_v = ~(notdor0_v);
  assign n_83_v = ~(n_1400_v);
  assign DA_AB2_v = ~(n_681_v);
  assign DA_AxB2_v = ~((n_1691_v|DA_AB2_v));
  assign n_519_v = ~(v(clk0_v));
  assign n_513_v = ~((op_T__bit_v|n_954_v|n_885_v));
  assign op_store_v = ~((ir6_v|ir5_v|notir7_v));
  assign op_T0_tay_v = ~((notir3_v|clock1_v|ir4_v|notir7_v|ir2_v|irline3_v|ir6_v|notir5_v));
  assign H1x1_v = ~(pipeUNK15_v);
  assign n_518_v = ~(n_1439_v);
  assign n_5_v = ~(a0_v);
  assign n_507_v = ~(n_1049_v);
  assign n_515_v = ~((n_1253_v|(n_783_v&n_1542_v)));
  assign n_465_v = ~(n_206_v);
  assign n_466_v = ~((dor6_v|RnWstretched_v));
  assign n_473_v = ~((n_1408_v&n_980_v));
  assign n_474_v = ~(((n_1643_v&n_1184_v)|n_410_v));
  assign n_830_v = ~((n_1505_v|n_43_v));
  assign n_1613_v = ~((RnWstretched_v|dor3_v));
  assign n_467_v = ~((n_470_v|n_134_v));
  assign n_468_v = ~(((n_16_v&pipeT4out_v)|(notRdy0_v&pipeT5out_v)));
  assign __AxB5__C45_v = ~((AxB5_v|_C45_v));
  assign n_831_v = ~(n_1719_v);
  assign n_1154_v = ~((notRdy0_v|n_959_v));
  assign notalucin_v = ~(alucin_v);
  assign alucout_v = ~(notalucout_v);
  assign n_1153_v = ~(abh7_v);
  assign op_clv_v = ~((ir6_v|irline3_v|notir4_v|notir3_v|notir7_v|notir5_v|ir2_v));
  assign n_1145_v = ~((notRdy0_v|op_T0_ora_v));
  assign n_1157_v = ~(n_291_v);
  assign n_1159_v = ~((n_1580_v|n_613_v));
  assign op_T2_stack_access_v = ~((irline3_v|ir4_v|ir2_v|_t2_v|ir7_v));
  assign x_op_T__adc_sbc_v = ~((notir0_v|notir6_v|clock2_v|notir5_v));
  assign n_1523_v = ~(abh6_v);
  assign n_442_v = ~(n_182_v);
  assign dor3_v = ~(notdor3_v);
  assign Pout3_v = ~(n_1194_v);
  assign n_441_v = ~(n_692_v);
  assign op_rmw_v = ~(n_790_v);
  assign n_436_v = ~(n_485_v);
  assign op_plp_pla_v = ~((notir3_v|ir7_v|notir5_v|irline3_v|ir2_v|ir4_v));
  assign n_1519_v = ~(v(adl4_v));
  assign C1x5Reset_v = ~(n_717_v);
  assign ir0_v = ~(n_310_v);
  assign n_916_v = ~((n_1517_v|(n_206_v&n_853_v)));
  assign n_917_v = ~((notRdy0_v|n_383_v));
  assign op_T3_mem_zp_idx_v = ~((notir2_v|ir3_v|notir4_v|_t3_v));
  assign n_905_v = ~((n_440_v&op_shift_v));
  assign n_1251_v = ~(n_1640_v);
  assign abl3_v = ~(_ABL3_v);
  assign alucin_v = ~(n_590_v);
  assign n_913_v = ~(n_1699_v);
  assign n_906_v = ~(n_1333_v);
  assign _t5_v = ~(n_378_v);
  assign op_T0_iny_dey_v = ~((ir2_v|clock1_v|ir4_v|ir5_v|irline3_v|notir3_v|notir7_v));
  assign dpc36_IPC_v = ~((n_1472_v&(n_1581_v|n_1570_v)));
  assign n_384_v = ~((n_946_v|n_1412_v|n_1258_v|op_ANDS_v));
  assign n_383_v = ~(op_T2_jsr_v);
  assign n_374_v = ~(v(db6_v));
  assign n_372_v = ~(notRdy0_v);
  assign n_378_v = ~((n_1357_v|n_18_v));
  assign abl1_v = ~(_ABL1_v);
  assign n_1474_v = ~(v(idb1_v));
  assign dasb3_v = ~(((n_432_v&n_345_v)|n_1097_v));
  assign n_1047_v = ~(n_830_v);
  assign x_op_jmp_v = ~((notir3_v|ir4_v|irline3_v|ir7_v|notir2_v|notir6_v));
  assign x_op_push_pull_v = ~((ir4_v|ir7_v|notir3_v|irline3_v|ir2_v));
  assign n_340_v = ~(op_clv_v);
  assign op_T4_v = ~(_t4_v);
  assign op_SUMS_v = ~((op_SRS_v|op_ANDS_v|op_ORS_v|op_EORS_v));
  assign n_1195_v = ~(abl6_v);
  assign n_1192_v = ~(((n_743_v|n_1488_v)&n_609_v));
  assign n_1190_v = ~(s2_v);
  assign x_op_T3_ind_y_v = ~((ir3_v|notir4_v|_t3_v|ir2_v|notir0_v));
  assign n_344_v = ~((n_410_v&n_392_v));
  assign n_345_v = ~(((n_8_v&n_876_v)|(n_986_v&n_600_v)));
  assign n_423_v = ~(v(idb7_v));
  assign n_91_v = ~(n_1529_v);
  assign n_109_v = ~(n_1380_v);
  assign n_118_v = ~(n_334_v);
  assign n_625_v = ~((n_43_v|n_459_v));
  assign n_122_v = ~(__AxB_6_v);
  assign op_T2_mem_zp_v = ~((ir4_v|notir2_v|_t2_v|ir3_v));
  assign n_626_v = ~(((pipeUNK01_v&n_1401_v)|(DBNeg_v&n_1269_v)));
  assign n_111_v = ~(v(db2_v));
  assign n_108_v = ~(n_1364_v);
  assign n_123_v = ~(v(adl0_v));
  assign n_110_v = ~(n_1691_v);
  assign n_762_v = ~((n_149_v|n_761_v));
  assign alu7_v = ~(notalu7_v);
  assign n_757_v = ~((DA_C45_v&n_647_v));
  assign n_763_v = ~(n_1534_v);
  assign n_767_v = ~(n_1138_v);
  assign DA_C45_v = ~(_C45_v);
  assign op_jmp_v = ~((irline3_v|notir3_v|ir7_v|ir4_v|notir6_v|notir2_v));
  assign n_769_v = ~((RnWstretched_v|dor0_v));
  assign abh4_v = ~(_ABH4_v);
  assign n_1130_v = ~((n_1109_v|n_1258_v|n_192_v|n_1002_v|n_862_v));
  assign n_1084_v = ~((alub6_v|alua6_v));
  assign n_1085_v = ~(((n_862_v&notRdy0_v)|(((nnT2BR_v&BRtaken_v)|n_646_v)&n_372_v)));
  assign n_1082_v = ~(((n_253_v&n_270_v)|(pipeUNK16_v&n_279_v)|(n_954_v&n_206_v)|(n_507_v&n_1224_v)));
  assign n_1083_v = ~(pd3_clearIR_v);
  assign op_T0_pla_v = ~((notir5_v|irline3_v|clock1_v|ir7_v|ir4_v|ir2_v|notir3_v|notir6_v));
  assign n_130_v = ~(n_220_v);
  assign n_133_v = ~((cclk_v|n_1404_v));
  assign n_132_v = ~(n_31_v);
  assign PD_n_0xx0xx0x_v = ~(PD_0xx0xx0x_v);
  assign pchp3_v = ~(n_1061_v);
  assign n_1335_v = ~(n_628_v);
  assign dpc35_PCHC_v = ~((n_1070_v|n_1007_v|n_1010_v|n_1265_v|n_923_v));
  assign n_1339_v = ~(n_799_v);
  assign op_T0_cpx_cpy_inx_iny_v = ~((notir7_v|clock1_v|ir4_v|irline3_v|notir6_v));
  assign _AxB_0__C0in_v = ~((__AxB_0_v|n_105_v));
  assign n_556_v = ~(a4_v);
  assign n_1323_v = ~(n_631_v);
  assign notir7_v = ~(ir7_v);
  assign _C78_v = ~((n_748_v|(C67_v&A_B7_v)));
  assign op_T__shift_a_v = ~((notir3_v|clock2_v|notir1_v|ir2_v|ir4_v|ir7_v));
  assign idl5_v = ~(notidl5_v);
  assign n_243_v = ~(v(idb1_v));
  assign n_242_v = ~(n_1521_v);
  assign A_B5_v = ~(n_1632_v);
  assign op_T0_cpy_iny_v = ~((ir5_v|irline3_v|clock1_v|notir7_v|ir4_v|notir6_v));
  assign op_ANDS_v = ~(n_669_v);
  assign pclp0_v = ~(n_526_v);
  assign op_T0_plp_v = ~((ir6_v|ir7_v|notir3_v|ir4_v|notir5_v|clock1_v|ir2_v|irline3_v));
  assign n_1225_v = ~((op_T2_ind_v|op_T2_zp_zp_idx_v));
  assign abl4_v = ~(_ABL4_v);
  assign n_1488_v = ~(n_278_v);
  assign op_T3_plp_pla_v = ~((ir7_v|ir2_v|irline3_v|ir4_v|notir3_v|_t3_v|notir5_v));
  assign n_396_v = ~(n_1358_v);
  assign n_390_v = ~(n_653_v);
  assign idl7_v = ~(notidl7_v);
  assign n_388_v = ~((DA_C01_v|n_936_v|DA_AxB2_v|AxB1_v));
  assign n_389_v = ~(n_1107_v);
  assign n_1492_v = ~(pipeUNK02_v);
  assign n_1486_v = ~((n_200_v|(n_1070_v&n_919_v)));
  assign n_1484_v = ~(y2_v);
  assign n_11_v = ~(((op_T0_tay_v|op_ANDS_v|op_T0_shift_a_v|op_T0_tax_v)|(op_T0_acc_v&n_397_v)));
  assign n_6_v = ~((n_43_v|n_521_v));
  assign n_16_v = ~(notRdy0_v);
  assign n_10_v = ~((n_467_v|n_1211_v|op_branch_done_v));
  assign n_19_v = ~((n_1708_v|n_770_v));
  assign op_T0_cmp_v = ~((notir6_v|notir7_v|clock1_v|notir0_v|ir5_v));
  assign aluvout_v = ~(n_408_v);
  assign n_944_v = ~((n_759_v|n_1449_v));
  assign n_946_v = ~((n_844_v&n_616_v));
  assign n_947_v = ~(a3_v);
  assign op_SRS_v = ~(n_366_v);
  assign n_935_v = ~(v(adl2_v));
  assign n_936_v = ~(aluanandb1_v);
  assign n_937_v = ~(pcl0_v);
  assign n_318_v = ~(p1_v);
  assign n_319_v = ~((DA_C01_v&n_936_v));
  assign n_149_v = ~(alu6_v);
  assign n_146_v = ~(n_5_v);
  assign n_154_v = ~(n_512_v);
  assign n_152_v = ~((op_T2_v|n_630_v|n_952_v|n_1002_v));
  assign DC78_v = ~((dpc18__DAA_v|((n_570_v|n_269_v)&(n_757_v|__AxB_6_v))));
  assign n_334_v = ~((p2_v|brk_done_v));
  assign alu6_v = ~(notalu6_v);
  assign n_332_v = ~(nots0_v);
  assign op_sta_cmp_v = ~((notir0_v|ir5_v|ir6_v|notir7_v));
  assign aluanorb0_v = ~((alub0_v|alua0_v));
  assign notRnWprepad_v = ~((notRdy0_v|C1x5Reset_v|pipe_WR_phi2_v));
  assign n_1179_v = ~((C34_v|dpc22__DSA_v));
  assign n_182_v = ~(((n_1262_v&n_236_v)|(n_1655_v|op_T5_rts_v|n_646_v)));
  assign n_188_v = ~((n_1606_v|n_1357_v));
  assign n_180_v = ~((notRdy0_v|n_1716_v));
  assign n_184_v = ~(y3_v);
  assign abl6_v = ~(_ABL6_v);
  assign n_177_v = ~(AxB7_v);
  assign n_192_v = ~((n_595_v&_op_branch_done_v));
  assign n_191_v = ~((n_790_v|notRdy0_v|n_347_v));
  assign n_673_v = ~((Pout3_v&op_T0_adc_sbc_v));
  assign n_964_v = ~((n_1533_v|pipe_T0_v));
  assign __AxBxC_1_v = ~((__AxB1__C01_v|(AxB1_v&_C01_v)));
  assign n_952_v = ~(n_272_v);
  assign n_958_v = ~(v(rdy_v));
  assign n_962_v = ~(n_1585_v);
  assign n_670_v = ~(n_519_v);
  assign n_681_v = ~((alua2_v&alub2_v));
  assign dasb6_v = ~(((n_739_v&n_61_v)|n_479_v));
  assign n_1218_v = ~(n_1565_v);
  assign __AxB7__C67_v = ~((_C67_v|AxB7_v));
  assign n_1213_v = ~((n_609_v|n_453_v));
  assign n_1224_v = ~(v(idb0_v));
  assign n_1215_v = ~((n_238_v|short_circuit_idx_add_v|brk_done_v));
  assign n_1214_v = ~(pipeUNK11_v);
  assign n_236_v = ~(n_1708_v);
  assign n_232_v = ~(pcl6_v);
  assign n_1223_v = ~((n_43_v|n_688_v));
  assign n_238_v = ~(pipeUNK35_v);
  assign n_720_v = ~((notRdy0_v|pipeUNK34_v));
  assign n_721_v = ~(nots7_v);
  assign n_723_v = ~(pclp3_v);
  assign pclp6_v = ~(n_993_v);
  assign n_726_v = ~((x_op_T4_ind_y_v|op_T5_ind_x_v|op_T3_abs_idx_ind_v|op_T5_rts_v));
  assign n_728_v = ~(VEC0_v);
  assign n_730_v = ~(x6_v);
  assign n_718_v = ~(v(db0_v));
  assign n_1718_v = ~(notRdy0_v);
  assign dpc22__DSA_v = ~(n_599_v);
  assign n_923_v = ~(pch3_v);
  assign _op_store_v = ~(op_store_v);
  assign DBNeg_v = ~(v(idb7_v));
  assign op_T2_php_pha_v = ~((ir2_v|notir3_v|ir5_v|ir4_v|ir7_v|_t2_v|irline3_v));
  assign n_933_v = ~((n_572_v&n_1262_v));
  assign n_920_v = ~(pipeUNK27_v);
  assign n_1206_v = ~(pchp7_v);
  assign n_1199_v = ~(v(db2_v));
  assign __AxBxC_6_v = ~((_AxB_6__C56_v|(__AxB_6_v&C56_v)));
  assign n_1202_v = ~(n_1265_v);
  assign op_T4_abs_idx_v = ~((notir3_v|notir4_v|_t4_v));
  assign n_355_v = ~(n_621_v);
  assign __AxBxC_0_v = ~(((n_105_v&__AxB_0_v)|_AxB_0__C0in_v));
  assign __AxB_6_v = ~((n_803_v&n_336_v));
  assign PD_0xx0xx0x_v = ~((pd1_clearIR_v|pd4_clearIR_v|pd7_clearIR_v));
  assign n_366_v = ~(((n_440_v&op_shift_right_v)|op_T0_shift_right_a_v));
  assign n_351_v = ~(v(idb6_v));
  assign op_T4_brk_v = ~((ir4_v|irline3_v|ir7_v|ir5_v|ir2_v|ir3_v|ir6_v|_t4_v));
  assign n_1458_v = ~(pclp6_v);
  assign n_1448_v = ~(n_1427_v);
  assign alu2_v = ~(notalu2_v);
  assign op_T3_ind_x_v = ~((_t3_v|notir0_v|ir2_v|ir4_v|ir3_v));
  assign n_1641_v = ~(pd1_clearIR_v);
  assign n_1640_v = ~(y7_v);
  assign abh0_v = ~(v(_ABH0_v));
  assign x_op_T3_plp_pla_v = ~((notir3_v|notir5_v|ir7_v|_t3_v|ir4_v|irline3_v|ir2_v));
  assign _C34_v = ~(((DC34_v|n_988_v)|(A_B3_v&C23_v)));
  assign n_1434_v = ~(x1_v);
  assign n_93_v = ~(v(db0_v));
  assign n_90_v = ~(n_1625_v);
  assign n_80_v = ~((n_267_v|n_1130_v));
  assign n_288_v = ~((RnWstretched_v|dor1_v));
  assign n_291_v = ~(n_1121_v);
  assign n_0_ADL0_v = ~(pipeVectorA0_v);
  assign n_218_v = ~(n_368_v);
  assign n_279_v = ~((n_253_v|n_954_v|n_507_v));
  assign n_280_v = ~(nots5_v);
  assign op_T4_mem_abs_idx_v = ~((notir4_v|_t4_v|notir3_v));
  assign n_282_v = ~(n_6_v);
  assign op_T0_tay_ldy_not_idx_v = ~((notir5_v|ir4_v|notir7_v|clock1_v|ir6_v|irline3_v));
  assign abh2_v = ~(_ABH2_v);
  assign n_1099_v = ~((n_1542_v&(n_1345_v|n_1166_v)));
  assign n_1101_v = ~((n_813_v&n_46_v));
  assign n_1109_v = ~((n_902_v|n_1464_v));
  assign n_1110_v = ~(n_756_v);
  assign n_1093_v = ~(n_968_v);
  assign n_1094_v = ~(v(adl5_v));
  assign n_1106_v = ~(((x_op_T0_txa_v|op_T0_txs_v|op_T0_dex_v|op_T0_cpx_inx_v|op_T2_ind_x_v)|(op_T2_idx_x_xy_v&n_1244_v)|(op_from_x_v&n_335_v)));
  assign n_1107_v = ~(((op_plp_pla_v|op_T3_ind_x_v|op_T2_ind_y_v|op_T3_abs_idx_v|op_T4_ind_y_v)|(n_440_v&op_inc_nop_v)));
  assign abl0_v = ~(_ABL0_v);
  assign n_1097_v = ~((n_345_v|n_432_v));
  assign n_480_v = ~(((n_888_v|n_118_v)&n_264_v));
  assign n_674_v = ~(n_25_v);
  assign n_678_v = ~((n_644_v|n_1357_v));
  assign op_T3_abs_idx_ind_v = ~((op_push_pull_v|notir3_v|_t3_v));
  assign n_1684_v = ~(v(idb6_v));
  assign n_1687_v = ~(v(idb0_v));
  assign n_669_v = ~((op_T0_and_v|op_T0_bit_v));
  assign n_696_v = ~((((n_1343_v|n_877_v)&n_79_v)|n_0_ADL0_v));
  assign _DA_ADD2_v = ~(alu2_v);
  assign n_1067_v = ~(n_582_v);
  assign idl2_v = ~(notidl2_v);
  assign clearIR_v = ~((fetch_v&D1x1_v));
  assign n_1075_v = ~(v(db4_v));
  assign op_T0_shift_right_a_v = ~((ir2_v|clock1_v|notir1_v|notir6_v|notir3_v|ir7_v|ir4_v));
  assign n_1073_v = ~((n_344_v&(n_410_v|n_392_v)));
  assign n_1081_v = ~(n_1560_v);
  assign pclp2_v = ~(n_1411_v);
  assign n_424_v = ~(n_198_v);
  assign n_1187_v = ~(s6_v);
  assign n_139_v = ~(op_SRS_v);
  assign op_from_x_v = ~((ir6_v|notir7_v|ir5_v|notir1_v));
  assign n_1548_v = ~(v(adl6_v));
  assign n_1531_v = ~(n_184_v);
  assign n_1534_v = ~((n_805_v|n_43_v));
  assign dasb5_v = ~((n_1629_v|(n_753_v&n_1135_v)));
  assign op_T2_idx_x_xy_v = ~((_t2_v|notir2_v|notir4_v));
  assign n_1549_v = ~(a1_v);
  assign n_262_v = ~(((pipeUNK29_v&n_1714_v)|(n_1511_v&pipeUNK28_v)));
  assign op_jsr_v = ~((ir7_v|irline3_v|ir3_v|notir5_v|ir4_v|ir2_v|ir6_v));
  assign n_260_v = ~((n_1205_v|n_852_v));
  assign n_1697_v = ~(n_664_v);
  assign n_995_v = ~(n_312_v);
  assign n_1374_v = ~((n_882_v|n_562_v));
  assign n_1375_v = ~(n_88_v);
  assign n_79_v = ~(n_236_v);
  assign C34_v = ~(_C34_v);
  assign n_71_v = ~(n_35_v);
  assign Reset0_v = ~(n_1395_v);
  assign _AxB_4__C34_v = ~((C34_v|__AxB_4_v));
  assign p6_v = ~(n_90_v);
  assign op_T0_dex_v = ~((notir1_v|clock1_v|notir6_v|ir2_v|notir7_v|ir4_v|notir3_v|ir5_v));
  assign n_75_v = ~(n_154_v);
  assign n_815_v = ~(pipeVectorA2_v);
  assign n_842_v = ~(abl1_v);
  assign n_837_v = ~(op_T0_eor_v);
  assign n_481_v = ~(pclp2_v);
  assign n_484_v = ~(((n_715_v|n_1316_v)&n_1386_v));
  assign n_485_v = ~(x4_v);
  assign __AxBxC_5_v = ~((__AxB5__C45_v|(AxB5_v&_C45_v)));
  assign op_T2_brk_v = ~((_t2_v|ir3_v|ir7_v|ir5_v|ir4_v|irline3_v|ir2_v|ir6_v));
  assign aluanandb1_v = ~((alub1_v&alua1_v));
  assign _op_branch_bit6_v = ~(ir6_v);
  assign n_844_v = ~((op_T0_ldx_tax_tsx_v|op_T__inx_v|op_T__dex_v));
  assign n_852_v = ~(v(sb7_v));
  assign n_853_v = ~(n_770_v);
  assign op_rti_rts_v = ~((ir4_v|ir7_v|notir6_v|ir3_v|ir2_v|irline3_v));
  assign n_847_v = ~(n_300_v);
  assign n_849_v = ~(n_321_v);
  assign n_850_v = ~(pipeUNK18_v);
  assign _TWOCYCLE_v = ~(((PD_n_0xx0xx0x_v&PD_xxxx10x0_v)|(PD_1xx000x0_v|PD_xxx010x1_v)));
  assign n_1647_v = ~(pclp7_v);
  assign op_T__bit_v = ~((irline3_v|ir6_v|ir7_v|clock2_v|notir5_v|notir2_v|ir4_v));
  assign AxB3_v = ~((n_649_v|n_988_v));
  assign n_641_v = ~(pcl7_v);
  assign n_1416_v = ~(v(idb6_v));
  assign op_T0_cld_sed_v = ~((notir6_v|ir2_v|irline3_v|notir7_v|notir3_v|notir4_v|clock1_v));
  assign alu3_v = ~(notalu3_v);
  assign dor6_v = ~(notdor6_v);
  assign n_207_v = ~((n_810_v|(n_923_v&n_293_v)));
  assign n_208_v = ~(pclp4_v);
  assign n_645_v = ~(v(NMIP_v));
  assign n_646_v = ~(n_17_v);
  assign n_981_v = ~(y5_v);
  assign n_980_v = ~(op_T3_jmp_v);
  assign n_662_v = ~(n_625_v);
  assign n_664_v = ~(op_implied_v);
  assign nnT2BR_v = ~(n_636_v);
  assign n_966_v = ~(n_1683_v);
  assign _t2_v = ~(n_1575_v);
  assign n_969_v = ~(n_161_v);
  assign n_658_v = ~(n_565_v);
  assign op_T3_branch_v = ~((ir2_v|_t3_v|notir4_v|irline3_v|ir3_v));
  assign n_1026_v = ~(n_567_v);
  assign n_1025_v = ~(y0_v);
  assign n_458_v = ~(v(idb2_v));
  assign x_op_T4_ind_y_v = ~((_t4_v|ir3_v|ir2_v|notir0_v|notir4_v));
  assign n_445_v = ~(n_862_v);
  assign op_T5_rti_rts_v = ~((_t5_v|notir6_v|ir2_v|ir3_v|irline3_v|ir4_v|ir7_v));
  assign x_op_T3_abs_idx_v = ~((_t3_v|notir4_v|notir3_v));
  assign dasb2_v = ~((n_1159_v|(n_1580_v&n_613_v)));
  assign n_1575_v = ~((n_1360_v|n_1357_v));
  assign ir3_v = ~(n_1620_v);
  assign n_1578_v = ~(pipe_VEC_v);
  assign n_1580_v = ~(v(sb2_v));
  assign n_440_v = ~(n_24_v);
  assign n_1507_v = ~(v(adl3_v));
  assign n_803_v = ~(n_1084_v);
  assign op_T4_brk_jsr_v = ~((irline3_v|ir6_v|ir2_v|ir3_v|ir7_v|_t4_v|ir4_v));
  assign n_1499_v = ~(n_1450_v);
  assign op_T0_and_v = ~((notir0_v|clock1_v|notir5_v|ir6_v|ir7_v));
  assign _C01_v = ~(C01_v);
  assign n_1500_v = ~(((dpc36_IPC_v&n_937_v)|n_1345_v));
  assign n_797_v = ~(v(idb4_v));
  assign n_800_v = ~(n_525_v);
  assign __AxBxC_2_v = ~((_AxB_2__C12_v|(__AxB_2_v&C12_v)));
  assign notir4_v = ~(ir4_v);
  assign n_31_v = ~(p0_v);
  assign n_34_v = ~(s3_v);
  assign op_T3_jmp_v = ~((ir7_v|notir6_v|notir2_v|_t3_v|notir3_v|ir4_v|irline3_v));
  assign n_25_v = ~((n_256_v|n_192_v));
  assign n_29_v = ~((Pout3_v&op_T0_sbc_v));
  assign n_27_v = ~(pchp4_v);
  assign n_753_v = ~((n_1257_v|n_811_v));
  assign n_733_v = ~(n_981_v);
  assign n_1610_v = ~((DA_AB2_v|AxB3_v));
  assign op_T4_rts_v = ~((ir2_v|ir3_v|notir6_v|ir4_v|notir5_v|irline3_v|_t4_v|ir7_v));
  assign n_1618_v = ~(n_419_v);
  assign n_1619_v = ~((n_1448_v|n_182_v));
  assign idl1_v = ~(notidl1_v);
  assign n_867_v = ~((_DA_ADD1_v|_DA_ADD2_v));
  assign n_862_v = ~(n_666_v);
  assign n_275_v = ~((n_773_v|n_1697_v));
  assign n_1621_v = ~(v(idb3_v));
  assign pd0_clearIR_v = ~((clearIR_v|pd0_v));
  assign n_1614_v = ~((pipeUNK03_v|n_1177_v|n_1111_v));
  assign op_T2_branch_v = ~((ir2_v|_t2_v|irline3_v|notir4_v|ir3_v));
  assign ir7_v = ~(n_541_v);
  assign n_611_v = ~((n_43_v|n_1509_v));
  assign dor7_v = ~(notdor7_v);
  assign n_36_v = ~((n_8_v|n_600_v));
  assign n_613_v = ~(((_DA_ADD1_v&n_600_v)|(n_8_v&n_1682_v)));
  assign n_1383_v = ~(v(idb5_v));
  assign ir2_v = ~(n_1300_v);
  assign n_62_v = ~(v(db7_v));
  assign brk_done_v = ~((notRdy0_v|n_861_v));
  assign n_1376_v = ~(v(idb2_v));
  assign n_1377_v = ~(op_rti_rts_v);
  assign op_ror_v = ~((ir7_v|notir5_v|notir6_v|notir1_v));
  assign __AxBxC_4_v = ~((_AxB_4__C34_v|(__AxB_4_v&C34_v)));
  assign n_647_v = ~(n_477_v);
  assign op_T0_ldy_mem_v = ~((irline3_v|notir7_v|notir2_v|ir6_v|notir5_v|clock1_v));
  assign n_1560_v = ~((op_T0_cmp_v|op_T0_cpx_cpy_inx_iny_v|n_1055_v));
  assign n_1566_v = ~(n_1221_v);
  assign op_brk_rti_v = ~((ir5_v|ir3_v|ir4_v|irline3_v|ir2_v|ir7_v));
  assign n_1561_v = ~(x7_v);
  assign n_477_v = ~((alua5_v&alub5_v));
  assign n_476_v = ~((n_1027_v|n_43_v));
  assign op_xy_v = ~((ir6_v|notir7_v|notir1_v));
  assign x_op_T4_rti_v = ~((ir2_v|irline3_v|ir5_v|ir7_v|notir6_v|ir4_v|ir3_v|_t4_v));
  assign n_472_v = ~(((pipeT3out_v&n_16_v)|(pipeT4out_v&notRdy0_v)));
  assign n_470_v = ~(n_646_v);
  assign n_1462_v = ~(n_1369_v);
  assign pd6_clearIR_v = ~((pd6_v|clearIR_v));
  assign VEC0_v = ~((notRdy0_v|n_689_v));
  assign n_1463_v = ~((RnWstretched_v|dor4_v));
  assign n_1469_v = ~(AxB5_v);
  assign op_rol_ror_v = ~((notir1_v|notir5_v|ir6_v|ir7_v));
  assign op_T5_jsr_v = ~((ir4_v|ir6_v|irline3_v|_t5_v|ir3_v|notir5_v|ir2_v|ir7_v));
  assign n_1471_v = ~(D1x1_v);
  assign n_774_v = ~(op_T0_cld_sed_v);
  assign ONEBYTE_v = ~(n_231_v);
  assign _C23_v = ~(C23_v);
  assign dasb1_v = ~((n_735_v|(n_36_v&n_320_v)));
  assign n_1007_v = ~(dpc34_PCLC_v);
  assign n_1016_v = ~(v(adl1_v));
  assign n_1010_v = ~(pch0_v);
  assign n_1018_v = ~(n_762_v);
  assign n_1017_v = ~(x5_v);
  assign n_70_v = ~((_VEC_v|n_1054_v));
  assign n_998_v = ~(nots3_v);
  assign op_implied_v = ~((x_op_push_pull_v|ir0_v|notir3_v|ir2_v));
  assign n_1289_v = ~(n_902_v);
  assign n_1033_v = ~(n_241_v);
  assign n_1024_v = ~(n_94_v);
  assign C23_v = ~((n_1691_v|(_C12_v&n_681_v)));
  assign A_B1_v = ~(aluanorb1_v);
  assign PD_xxxx10x0_v = ~((pd0_clearIR_v|pd2_clearIR_v|n_1083_v));
  assign op_T3_stack_bit_jmp_v = ~((_t3_v|ir4_v|ir7_v|irline3_v));
  assign n_1028_v = ~(n_251_v);
  assign n_890_v = ~(x2_v);
  assign n_1044_v = ~((n_31_v|n_812_v));
  assign n_732_v = ~(((n_1528_v&_TWOCYCLE_phi1_v)|n_1161_v));
  assign n_1034_v = ~(abh2_v);
  assign _DBE_v = ~((cclk_v|n_962_v));
  assign n_603_v = ~(n_47_v);
  assign n_1045_v = ~(n_69_v);
  assign n_1039_v = ~(((pipeUNK39_v&notRdy0_v)|pipeUNK40_v));
  assign n_1043_v = ~(n_818_v);
  assign n_1037_v = ~((op_T2_pha_v|(op_sta_cmp_v&n_335_v)));
  assign n_1038_v = ~(n_336_v);
  assign n_782_v = ~((n_383_v&n_1303_v));
  assign n_490_v = ~(v(db4_v));
  assign n_501_v = ~((n_180_v|Reset0_v|n_819_v));
  assign C56_v = ~(_C56_v);
  assign n_499_v = ~(pch5_v);
  assign n_496_v = ~(s5_v);
  assign op_T5_ind_y_v = ~((_t5_v|notir4_v|ir2_v|ir3_v|notir0_v));
  assign n_880_v = ~(v(adh6_v));
  assign fetch_v = ~((notRdy0_v|n_1214_v));
  assign n_1677_v = ~(abh4_v);
  assign ir4_v = ~(n_927_v);
  assign n_1111_v = ~((pipeUNK07_v&pipeUNK09_v));
  assign n_1115_v = ~((n_620_v|n_270_v));
  assign op_T0_clc_sec_v = ~((irline3_v|ir6_v|ir2_v|ir7_v|notir3_v|clock1_v|notir4_v));
  assign n_1117_v = ~(n_70_v);
  assign idl6_v = ~(notidl6_v);
  assign n_1120_v = ~(notRdy0_v);
  assign n_410_v = ~((n_1184_v|n_1643_v));
  assign notalucout_v = ~((DC78_phi2_v|C78_phi2_v));
  assign n_783_v = ~(pcl2_v);
  assign n_1654_v = ~(n_947_v);
  assign op_T0_cpx_inx_v = ~((notir6_v|notir5_v|clock1_v|irline3_v|notir7_v|ir4_v));
  assign n_1705_v = ~((n_467_v|n_630_v));
  assign n_1655_v = ~(n_1211_v);
  assign n_1688_v = ~(n_1304_v);
  assign n_1708_v = ~(op_T3_branch_v);
  assign n_896_v = ~(v(db3_v));
  assign op_EORS_v = ~(n_837_v);
  assign n_882_v = ~((n_597_v|n_1252_v));
  assign n_883_v = ~(v(adh3_v));
  assign n_1662_v = ~(n_1124_v);
  assign n_1676_v = ~(abl4_v);
  assign n_1668_v = ~(v(adh0_v));
  assign pd2_clearIR_v = ~((clearIR_v|pd2_v));
  assign n_1400_v = ~(pch4_v);
  assign n_1399_v = ~(n_1715_v);
  assign n_1398_v = ~((alua7_v|alub7_v));
  assign op_T0_shift_a_v = ~((ir4_v|notir3_v|clock1_v|ir7_v|ir2_v|notir1_v));
  assign notir5_v = ~(ir5_v);
  assign n_1392_v = ~(v(nmi_v));
  assign n_160_v = ~((op_SRS_v|n_781_v));
  assign n_1255_v = ~(n_531_v);
  assign op_T0_adc_sbc_v = ~((notir0_v|clock1_v|notir6_v|notir5_v));
  assign n_564_v = ~(n_1025_v);
  assign n_567_v = ~(_ABL7_v);
  assign n_566_v = ~(((n_243_v&n_781_v)|(n_755_v&_DBZ_v)|(n_1170_v&pipeUNK14_v)));
  assign n_570_v = ~((DA_C45_v|n_647_v|AxB5_v|n_122_v));
  assign n_568_v = ~(v(db5_v));
  assign n_163_v = ~(n_249_v);
  assign n_161_v = ~((n_1113_v|cclk_v));
  assign n_172_v = ~(abl5_v);
  assign n_169_v = ~((n_1624_v|n_139_v));
  assign n_168_v = ~(v(adh2_v));
  assign op_T0_tax_v = ~((ir2_v|notir5_v|notir1_v|ir4_v|notir7_v|notir3_v|ir6_v|clock1_v));
  assign n_347_v = ~((op_T2_mem_zp_v|op_T3_mem_zp_idx_v|op_T3_mem_abs_v|op_T4_mem_abs_idx_v|op_T5_mem_ind_idx_v));
  assign ir6_v = ~(n_1675_v);
  assign n_176_v = ~((n_10_v|n_236_v));
  assign _AxB_6__C56_v = ~((__AxB_6_v|C56_v));
  assign op_T4_ind_x_v = ~((ir2_v|notir0_v|_t4_v|ir4_v|ir3_v));
  assign n_1318_v = ~((alua7_v&alub7_v));
  assign n_1319_v = ~(v(db1_v));
  assign notaluvout_v = ~((n_637_v|(n_1398_v&C67_v)));
  assign n_1309_v = ~(pd6_clearIR_v);
  assign __AxBxC_7_v = ~((__AxB7__C67_v|(_C67_v&AxB7_v)));
  assign n_531_v = ~(n_95_v);
  assign pchp7_v = ~(n_663_v);
  assign n_533_v = ~(pipeUNK22_v);
  assign op_T4_rti_v = ~((notir6_v|ir4_v|irline3_v|_t4_v|ir2_v|ir3_v|ir5_v|ir7_v));
  assign n_1312_v = ~((n_1291_v|n_1693_v));
  assign op_T2_ind_v = ~((ir3_v|ir2_v|notir0_v|_t2_v));
  assign __AxB_0_v = ~((aluaorb0_v&aluanandb0_v));
  assign __AxBxC_3_v = ~((__AxB3__C23_v|(_C23_v&AxB3_v)));
  assign n_278_v = ~(pch6_v);
  assign n_1517_v = ~((n_572_v|n_853_v));
  assign n_1518_v = ~(n_1270_v);
  assign n_1511_v = ~(pipeUNK29_v);
  assign op_T2_abs_y_v = ~((notir4_v|ir2_v|notir0_v|notir3_v|_t2_v));
  assign n_272_v = ~((n_646_v|nnT2BR_v|op_T5_rts_v|op_T2_abs_access_v|n_862_v|n_236_v));
  assign op_T2_abs_access_v = ~((_t2_v|op_push_pull_v|notir3_v));
  assign n_1295_v = ~(n_1527_v);
  assign n_1304_v = ~((op_T0_sbc_v|n_673_v));
  assign n_1305_v = ~(n_772_v);
  assign n_1301_v = ~(pchp5_v);
  assign n_3_v = ~(nots4_v);
  assign idl4_v = ~(notidl4_v);
  assign n_510_v = ~((x_op_jmp_v|op_rmw_v|n_347_v));
  assign op_T5_rts_v = ~((ir7_v|notir6_v|ir4_v|ir2_v|notir5_v|_t5_v|irline3_v|ir3_v));
  assign n_1303_v = ~(((op_sty_cpy_mem_v&n_335_v)|(op_from_x_v&n_335_v)));
  assign op_T0_cli_sei_v = ~((ir7_v|ir2_v|notir6_v|clock1_v|notir3_v|irline3_v|notir4_v));
  assign n_819_v = ~((pipeUNK23_v|pipephi2Reset0_v));
  assign op_T__adc_sbc_v = ~((notir6_v|notir5_v|clock2_v|notir0_v));
  assign n_368_v = ~((xx_op_T5_jsr_v|x_op_T3_plp_pla_v|op_T4_jmp_v|op_T5_rti_rts_v|op_T2_jmp_abs_v|op_T2_php_pha_v));
  assign op_T5_brk_v = ~((ir7_v|ir3_v|ir5_v|ir2_v|irline3_v|_t5_v|ir6_v|ir4_v));
  assign n_818_v = ~((n_43_v|n_265_v));
  assign n_813_v = ~((n_1258_v|n_440_v));
  assign n_824_v = ~((op_T2_brk_v|op_T3_jsr_v));
  assign n_1595_v = ~(n_754_v);
  assign n_1594_v = ~((n_779_v&n_604_v));
  assign n_196_v = ~(n_543_v);
  assign notir0_v = ~(ir0_v);
  assign _AxB_2__C12_v = ~((C12_v|__AxB_2_v));
  assign n_1166_v = ~(n_329_v);
  assign n_630_v = ~(n_726_v);
  assign n_201_v = ~(_op_branch_bit7_v);
  assign n_200_v = ~((n_919_v|n_1070_v));
  assign n_386_v = ~(pcl5_v);
  assign n_631_v = ~(n_878_v);
  assign INTG_v = ~((n_760_v|brk_done_v));
  assign n_1356_v = ~(a6_v);
  assign n_14_v = ~((n_671_v|n_323_v|Reset0_v));
  assign n_17_v = ~((n_964_v|n_732_v));
  assign n_1638_v = ~(v(db6_v));
  assign n_1046_v = ~(v(adl7_v));
  assign n_1631_v = ~(((n_1253_v|n_163_v)&n_1184_v));
  assign n_1632_v = ~((alua5_v|alub5_v));
  assign dor2_v = ~(notdor2_v);
  assign n_1635_v = ~(n_966_v);
  assign n_919_v = ~((n_311_v&dpc34_PCLC_v));
  assign n_918_v = ~(n_404_v);
  assign aluanandb0_v = ~((alub0_v&alua0_v));
  assign n_1629_v = ~((n_1135_v|n_753_v));
  assign n_1592_v = ~(n_128_v);
  assign n_1599_v = ~(v(irq_v));
  assign n_220_v = ~(n_190_v);
  assign n_618_v = ~(nots6_v);
  assign n_629_v = ~((n_50_v|((n_646_v|nnT2BR_v)&n_480_v)));
  assign n_1002_v = ~(n_1219_v);
  assign n_224_v = ~((RnWstretched_v|dor2_v));
  assign n_628_v = ~((n_55_v|cclk_v));
  assign n_617_v = ~(abh1_v);
  assign n_221_v = ~(n_1579_v);
  assign n_620_v = ~((n_1371_v|n_1433_v|n_1293_v|n_307_v));
  assign n_616_v = ~((op_T0_tay_ldy_not_idx_v|op_T__iny_dey_v|op_T0_ldy_mem_v));
  assign _VEC_v = ~((VEC0_v|VEC1_v));
  assign n_1129_v = ~((cp1_v|n_358_v));
  assign n_1137_v = ~((n_790_v&_op_store_v));
  assign n_1133_v = ~((ir0_v|ir1_v));
  assign n_1141_v = ~(n_982_v);
  assign n_1135_v = ~(v(sb5_v));
  assign op_T0_txa_v = ~((ir4_v|ir5_v|notir3_v|notir1_v|notir7_v|ir2_v|ir6_v|clock1_v));
  assign n_1138_v = ~(y1_v);
  assign n_392_v = ~(n_386_v);
  assign n_400_v = ~(n_834_v);
  assign n_0_ADL2_v = ~(n_815_v);
  assign n_1194_v = ~(p3_v);
  assign short_circuit_idx_add_v = ~((notRdy0_v|n_1137_v|n_916_v|pipeUNK36_v));
  assign notir2_v = ~(ir2_v);
  assign n_1184_v = ~((n_163_v&n_1253_v));
  assign n_127_v = ~((n_519_v|cp1_v));
  assign n_128_v = ~(a7_v);
  assign n_134_v = ~((op_jsr_v|op_brk_rti_v|x_op_jmp_v));
  assign n_861_v = ~(n_1452_v);
  assign n_1238_v = ~(n_1295_v);
  assign ir5_v = ~(n_1609_v);
  assign op_shift_right_v = ~((notir1_v|notir6_v|ir7_v));
  assign n_1245_v = ~(aluvout_v);
  assign n_1244_v = ~(op_xy_v);
  assign op_T__ora_and_eor_adc_v = ~((ir7_v|clock2_v|notir0_v));
  assign AxB7_v = ~((n_1398_v|n_748_v));
  assign n_1240_v = ~(n_1566_v);
  assign n_241_v = ~(n_745_v);
  assign n_249_v = ~(pcl3_v);
  assign n_251_v = ~((n_221_v|_DBE_v));
  assign op_T0_txs_v = ~((notir3_v|notir4_v|ir5_v|ir6_v|notir7_v|ir2_v|notir1_v|clock1_v));
  assign _op_set_C_v = ~(((op_T__cpx_cpy_abs_v|op_T__asl_rol_a_v|op_T__cpx_cpy_imm_zp_v|x_op_T__adc_sbc_v|op_T__cmp_v)|(op_asl_rol_v&n_1258_v)));
  assign n_253_v = ~(pipeUNK42_v);
  assign A_B7_v = ~(n_1398_v);
  assign pchp1_v = ~(n_126_v);
  assign op_T3_v = ~(_t3_v);
  assign _C56_v = ~(((A_B5_v&C45_v)|n_647_v));
  assign n_350_v = ~((alub3_v&alua3_v));
  assign n_335_v = ~((n_347_v|_op_store_v));
  assign n_336_v = ~((alua6_v&alub6_v));
  assign VEC1_v = ~(n_698_v);
  assign op_T__iny_dey_v = ~((ir5_v|notir7_v|clock2_v|irline3_v|notir3_v|ir2_v|ir4_v));
  assign x_op_T0_bit_v = ~((ir7_v|ir4_v|clock1_v|notir5_v|notir2_v|irline3_v|ir6_v));
  assign op_T0_brk_rti_v = ~((irline3_v|ir5_v|ir2_v|ir3_v|ir7_v|ir4_v|clock1_v));
  assign n_432_v = ~(v(sb3_v));
  assign n_428_v = ~(((n_16_v&pipeT2out_v)|(pipeT3out_v&notRdy0_v)));
  assign op_T__cmp_v = ~((notir7_v|notir6_v|clock2_v|notir0_v|ir5_v));
  assign n_312_v = ~(v(res_v));
  assign n_311_v = ~(n_1010_v);
  assign op_T2_jmp_abs_v = ~((ir5_v|irline3_v|ir4_v|_t2_v|notir2_v|ir7_v|notir6_v|notir3_v));
  assign __AxB_4_v = ~((n_918_v&n_1063_v));
  assign n_1089_v = ~(n_1574_v);
  assign dor4_v = ~(notdor4_v);
  assign n_1091_v = ~(((n_16_v&pipeT_SYNC_v)|(notRdy0_v&pipeT2out_v)));
  assign n_1090_v = ~((op_T2_stack_access_v|n_1222_v));
  assign n_1087_v = ~((n_717_v|brk_done_v));
  assign op_T2_pha_v = ~((ir4_v|ir5_v|notir6_v|notir3_v|irline3_v|ir7_v|_t2_v|ir2_v));
  assign n_979_v = ~(n_905_v);
  assign n_20_v = ~((n_1316_v|(n_344_v&n_232_v)));
  assign n_739_v = ~(((n_1056_v&n_811_v)|(n_761_v&n_1257_v)));
  assign n_748_v = ~(n_1318_v);
  assign __AxB1__C01_v = ~((AxB1_v|_C01_v));
  assign n_293_v = ~((n_200_v&n_1202_v));
  assign n_300_v = ~((brk_done_v|op_T2_jsr_v|n_389_v|op_rti_rts_v|x_op_T3_ind_y_v|op_T4_ind_x_v));
  assign n_299_v = ~(((pipeUNK05_v&n_1614_v)|(n_1416_v&n_1111_v)|(n_1245_v&pipeUNK03_v)|n_587_v));
  assign n_1230_v = ~((n_360_v|n_43_v));
  assign n_1231_v = ~(n_1409_v);
  assign op_T4_jmp_v = ~((notir6_v|ir4_v|_t4_v|notir3_v|ir7_v|irline3_v|notir2_v));
  assign n_1229_v = ~(((n_311_v|dpc34_PCLC_v)&n_919_v));
  assign op_T0_bit_v = ~((ir6_v|clock1_v|notir5_v|ir4_v|notir2_v|irline3_v|ir7_v));
  assign n_358_v = ~(v(clk0_v));
  assign D1x1_v = ~((C1x5Reset_v|INTG_v));
  assign n_1169_v = ~(n_987_v);
  assign n_1170_v = ~((n_755_v|n_781_v));
  assign n_1180_v = ~((pipe_T0_v|notRdy0_v));
  assign n_1181_v = ~(((n_1595_v&pipeUNK13_v)|(DBNeg_v&n_754_v)));
  assign n_1175_v = ~(n_1447_v);
  assign n_1178_v = ~((pipeUNK30_v|pipeUNK32_v|pipeUNK31_v|pipeUNK33_v));
  assign x_op_T0_tya_v = ~((notir3_v|ir6_v|ir2_v|notir4_v|clock1_v|notir7_v|ir5_v|irline3_v));
  assign _op_branch_bit7_v = ~(ir7_v);
  assign n_8_v = ~(n_551_v);
  assign n_743_v = ~((n_523_v|n_499_v));
  assign DBZ_v = ~((v(idb7_v)|v(idb6_v)|v(idb5_v)|v(idb2_v)|v(idb1_v)|v(idb0_v)|v(idb4_v)|v(idb3_v)));
  assign n_735_v = ~((n_320_v|n_36_v));
  assign n_21_v = ~((n_43_v|n_1162_v));
  assign dor1_v = ~(notdor1_v);
  assign n_747_v = ~(n_670_v);

  spice_mux_2 mux_6281(eclk, ereset, dpc11_SBADD_v,dpc12_0ADD_v, v(sb0_v),1'b0, alua0_v);
  spice_mux_2 mux_6280(eclk, ereset, dpc11_SBADD_v,dpc12_0ADD_v, v(sb3_v),1'b0, alua3_v);
  spice_mux_2 mux_6283(eclk, ereset, n_1157_v,n_291_v, 1'b0,1'b1, dpc41_DL_ADL_v);
  spice_mux_2 mux_6282(eclk, ereset, dpc11_SBADD_v,dpc12_0ADD_v, v(sb1_v),1'b0, alua1_v);
  spice_mux_2 mux_6285(eclk, ereset, n_476_v,(cclk_v|n_1247_v|n_956_v), 1'b1,1'b0, dpc12_0ADD_v);
  spice_mux_2 mux_6284(eclk, ereset, n_631_v,n_1323_v, 1'b1,1'b0, dpc37_PCLDB_v);
  spice_mux_2 mux_6287(eclk, ereset, n_445_v,n_317_v, 1'b0,1'b1, n_417_v);
  spice_mux_2 mux_6286(eclk, ereset, n_355_v,n_593_v, 1'b1,1'b0, dpc4_SSB_v);
  spice_mux_2 mux_6289(eclk, ereset, cclk_v,dpc1_SBY_v, n_564_v,v(sb0_v), y0_v);
  spice_mux_2 mux_6288(eclk, ereset, dpc1_SBY_v,cclk_v, v(sb1_v),n_767_v, y1_v);
  spice_mux_2 mux_6362(eclk, ereset, n_692_v,(n_441_v|cclk_v|n_1247_v), 1'b1,1'b0, dpc1_SBY_v);
  spice_mux_2 mux_6363(eclk, ereset, n_1467_v,n_1129_v, 1'b0,1'b1, cclk_v);
  spice_mux_2 mux_6360(eclk, ereset, n_769_v,(dor0_v|RnWstretched_v), 1'b1,1'b0, n_1072_v);
  spice_mux_2 mux_6361(eclk, ereset, n_617_v,abh1_v, 1'b0,1'b1, n_1140_v);
  spice_mux_2 mux_6366(eclk, ereset, n_1153_v,abh7_v, 1'b0,1'b1, n_1639_v);
  spice_mux_2 mux_6367(eclk, ereset, abl5_v,n_172_v, 1'b0,1'b1, n_210_v);
  spice_mux_2 mux_6364(eclk, ereset, n_1028_v,n_251_v, 1'b1,1'b0, RnWstretched_v);
  spice_mux_2 mux_6365(eclk, ereset, abl5_v,n_172_v, 1'b1,1'b0, n_1633_v);
  spice_mux_2 mux_6368(eclk, ereset, n_424_v,n_198_v, 1'b1,1'b0, notRdy0_v);
  spice_mux_2 mux_6369(eclk, ereset, n_127_v,n_135_v, 1'b1,1'b0, clk2out_v);
  spice_mux_2 mux_6223(eclk, ereset, n_1545_v,n_994_v, 1'b1,1'b0, ab10_v);
  spice_mux_2 mux_6222(eclk, ereset, n_1608_v,n_869_v, 1'b1,1'b0, ab13_v);
  spice_mux_2 mux_6221(eclk, ereset, n_999_v,n_475_v, 1'b0,1'b1, ab12_v);
  spice_mux_2 mux_6220(eclk, ereset, dor0_v,(RnWstretched_v|n_769_v), 1'b1,1'b0, n_1325_v);
  spice_mux_2 mux_6227(eclk, ereset, n_288_v,(dor1_v|RnWstretched_v), 1'b1,1'b0, n_794_v);
  spice_mux_2 mux_6225(eclk, ereset, n_963_v,n_635_v, 1'b1,1'b0, ab14_v);
  spice_mux_2 mux_6224(eclk, ereset, n_1296_v,n_359_v, 1'b1,1'b0, ab11_v);
  spice_mux_2 mux_6229(eclk, ereset, cclk_v,(cp1_v&fetch_v), notir2_v,n_571_v, n_1300_v);
  spice_mux_2 mux_6228(eclk, ereset, dor1_v,(RnWstretched_v|n_288_v), 1'b1,1'b0, n_798_v);
  spice_mux_2 mux_6209(eclk, ereset, n_1256_v,n_91_v, 1'b0,1'b1, dpc15_ANDS_v);
  spice_mux_2 mux_6208(eclk, ereset, dpc6_SBS_v,dpc7_SS_v, v(sb4_v),n_3_v, s4_v);
  spice_mux_2 mux_6253(eclk, ereset, (cp1_v&fetch_v),cclk_v, n_928_v,notir5_v, n_1609_v);
  spice_mux_2 mux_6255(eclk, ereset, n_35_v,(n_1247_v|cclk_v|n_71_v), 1'b1,1'b0, dpc7_SS_v);
  spice_mux_2 mux_6259(eclk, ereset, cclk_v,dpc3_SBX_v, n_242_v,v(sb3_v), x3_v);
  spice_mux_2 mux_6269(eclk, ereset, dpc40_ADLPCL_v,dpc39_PCLPCL_v, v(adl0_v),n_488_v, pcl0_v);
  spice_mux_2 mux_6268(eclk, ereset, dpc40_ADLPCL_v,dpc39_PCLPCL_v, v(adl1_v),n_976_v, pcl1_v);
  spice_mux_2 mux_6267(eclk, ereset, dpc40_ADLPCL_v,dpc39_PCLPCL_v, v(adl2_v),n_481_v, pcl2_v);
  spice_mux_2 mux_6266(eclk, ereset, dpc40_ADLPCL_v,dpc39_PCLPCL_v, v(adl3_v),n_723_v, pcl3_v);
  spice_mux_2 mux_6265(eclk, ereset, abh6_v,n_1523_v, 1'b1,1'b0, n_963_v);
  spice_mux_2 mux_6264(eclk, ereset, cclk_v,dpc3_SBX_v, n_578_v,v(sb5_v), x5_v);
  spice_mux_2 mux_6263(eclk, ereset, dpc3_SBX_v,cclk_v, v(sb4_v),n_436_v, x4_v);
  spice_mux_2 mux_6262(eclk, ereset, cclk_v,dpc3_SBX_v, n_871_v,v(sb7_v), x7_v);
  spice_mux_2 mux_6261(eclk, ereset, cclk_v,dpc3_SBX_v, n_1709_v,v(sb1_v), x1_v);
  spice_mux_2 mux_6260(eclk, ereset, dpc3_SBX_v,cclk_v, v(sb0_v),n_1169_v, x0_v);
  spice_mux_3 mux_6375(eclk, ereset, dpc9_DBADD_v,dpc8_nDBADD_v,dpc10_ADLADD_v, v(idb5_v),n_1383_v,v(adl5_v), alub5_v);
  spice_mux_2 mux_6377(eclk, ereset, n_1441_v,n_1277_v, 1'b0,1'b1, dpc42_DL_ADH_v);
  spice_mux_3 mux_6376(eclk, ereset, dpc9_DBADD_v,dpc8_nDBADD_v,dpc10_ADLADD_v, v(idb4_v),n_478_v,v(adl4_v), alub4_v);
  spice_mux_2 mux_6245(eclk, ereset, dpc31_PCHPCH_v,dpc30_ADHPCH_v, n_1301_v,v(adh5_v), pch5_v);
  spice_mux_2 mux_6247(eclk, ereset, dpc31_PCHPCH_v,dpc30_ADHPCH_v, n_141_v,v(adh3_v), pch3_v);
  spice_mux_2 mux_6246(eclk, ereset, dpc31_PCHPCH_v,dpc30_ADHPCH_v, n_27_v,v(adh4_v), pch4_v);
  spice_mux_3 mux_6242(eclk, ereset, dpc8_nDBADD_v,dpc10_ADLADD_v,dpc9_DBADD_v, n_458_v,v(adl2_v),v(idb2_v), alub2_v);
  spice_mux_2 mux_6249(eclk, ereset, dpc31_PCHPCH_v,dpc30_ADHPCH_v, n_209_v,v(adh1_v), pch1_v);
  spice_mux_2 mux_6248(eclk, ereset, dpc30_ADHPCH_v,dpc31_PCHPCH_v, v(adh2_v),n_1496_v, pch2_v);
  spice_mux_2 mux_6188(eclk, ereset, (ADL_ABL_v&cp1_v),cclk_v, n_1507_v,n_138_v, _ABL3_v);
  spice_mux_2 mux_6189(eclk, ereset, cclk_v,(ADL_ABL_v&cp1_v), n_642_v,n_935_v, _ABL2_v);
  spice_mux_2 mux_6186(eclk, ereset, (ADL_ABL_v&cp1_v),cclk_v, n_1548_v,n_1254_v, _ABL6_v);
  spice_mux_2 mux_6187(eclk, ereset, (ADL_ABL_v&cp1_v),cclk_v, n_1094_v,n_210_v, _ABL5_v);
  spice_mux_2 mux_6184(eclk, ereset, cp1_v,n_38_v, 1'b0,1'b1, n_1247_v);
  spice_mux_2 mux_6185(eclk, ereset, (ADL_ABL_v&cp1_v),cclk_v, n_1046_v,n_171_v, _ABL7_v);
  spice_mux_2 mux_6244(eclk, ereset, dpc31_PCHPCH_v,dpc30_ADHPCH_v, n_652_v,v(adh6_v), pch6_v);
  spice_mux_2 mux_6241(eclk, ereset, (cp1_v&fetch_v),cclk_v, n_227_v,notir4_v, n_927_v);
  spice_mux_3 mux_6240(eclk, ereset, cclk_v,n_1315_v,abh0_v, v(_ABH0_v),1'b1,1'b0, n_381_v);
  spice_mux_2 mux_6243(eclk, ereset, dpc31_PCHPCH_v,dpc30_ADHPCH_v, n_1206_v,v(adh7_v), pch7_v);
  spice_mux_2 mux_6354(eclk, ereset, dpc23_SBAC_v,cclk_v, dasb5_v,n_831_v, a5_v);
  spice_mux_2 mux_6313(eclk, ereset, n_611_v,(cclk_v|n_1247_v|n_255_v), 1'b1,1'b0, dpc31_PCHPCH_v);
  spice_mux_2 mux_6312(eclk, ereset, n_625_v,(n_1247_v|n_662_v|cclk_v), 1'b1,1'b0, dpc3_SBX_v);
  spice_mux_2 mux_6311(eclk, ereset, n_1305_v,n_772_v, 1'b0,1'b1, dpc17_SUMS_v);
  spice_mux_3 mux_6310(eclk, ereset, n_1423_v,cclk_v,abh5_v, 1'b1,v(_ABH5_v),1'b0, n_869_v);
  spice_mux_2 mux_6317(eclk, ereset, n_1223_v,(cclk_v|n_1247_v|n_225_v), 1'b1,1'b0, dpc9_DBADD_v);
  spice_mux_2 mux_6316(eclk, ereset, n_1315_v,abh0_v, 1'b0,1'b1, n_826_v);
  spice_mux_3 mux_6315(eclk, ereset, n_1153_v,cclk_v,abh7_v, 1'b1,v(_ABH7_v),1'b0, n_659_v);
  spice_mux_3 mux_6314(eclk, ereset, abh1_v,n_617_v,cclk_v, 1'b0,1'b1,v(_ABH1_v), n_676_v);
  spice_mux_2 mux_6319(eclk, ereset, n_321_v,n_849_v, 1'b1,1'b0, dpc33_PCHDB_v);
  spice_mux_3 mux_6318(eclk, ereset, n_1346_v,abh3_v,cclk_v, 1'b1,1'b0,v(_ABH3_v), n_359_v);
  spice_mux_2 mux_6279(eclk, ereset, dpc11_SBADD_v,dpc12_0ADD_v, v(sb2_v),1'b0, alua2_v);
  spice_mux_2 mux_6339(eclk, ereset, n_133_v,(n_602_v|cclk_v|n_1247_v), 1'b1,1'b0, dpc2_XSB_v);
  spice_mux_2 mux_6338(eclk, ereset, abl4_v,n_1676_v, 1'b0,1'b1, n_86_v);
  spice_mux_2 mux_6331(eclk, ereset, n_1041_v,n_138_v, 1'b1,1'b0, ab3_v);
  spice_mux_2 mux_6330(eclk, ereset, n_1152_v,n_642_v, 1'b1,1'b0, ab2_v);
  spice_mux_2 mux_6333(eclk, ereset, n_210_v,n_1633_v, 1'b0,1'b1, ab5_v);
  spice_mux_2 mux_6332(eclk, ereset, n_86_v,n_634_v, 1'b0,1'b1, ab4_v);
  spice_mux_2 mux_6335(eclk, ereset, n_322_v,n_171_v, 1'b1,1'b0, ab7_v);
  spice_mux_2 mux_6334(eclk, ereset, n_1191_v,n_1254_v, 1'b1,1'b0, ab6_v);
  spice_mux_2 mux_6337(eclk, ereset, n_1140_v,n_676_v, 1'b1,1'b0, ab9_v);
  spice_mux_2 mux_6336(eclk, ereset, n_826_v,n_381_v, 1'b1,1'b0, ab8_v);
  spice_mux_2 mux_6302(eclk, ereset, n_1676_v,abl4_v, 1'b0,1'b1, n_634_v);
  spice_mux_2 mux_6298(eclk, ereset, n_966_v,n_1635_v, 1'b1,1'b0, dpc29_0ADH17_v);
  spice_mux_2 mux_6299(eclk, ereset, n_525_v,(n_800_v|cclk_v|n_1247_v), 1'b1,1'b0, dpc26_ACDB_v);
  spice_mux_2 mux_6296(eclk, ereset, n_1230_v,(n_708_v|cclk_v|n_1247_v), 1'b1,1'b0, dpc11_SBADD_v);
  spice_mux_2 mux_6297(eclk, ereset, n_1541_v,(n_1247_v|n_491_v|cclk_v), 1'b1,1'b0, dpc10_ADLADD_v);
  spice_mux_2 mux_6294(eclk, ereset, cclk_v,dpc1_SBY_v, n_1251_v,v(sb7_v), y7_v);
  spice_mux_2 mux_6295(eclk, ereset, cclk_v,dpc1_SBY_v, n_518_v,v(sb6_v), y6_v);
  spice_mux_2 mux_6292(eclk, ereset, dpc1_SBY_v,cclk_v, v(sb5_v),n_733_v, y5_v);
  spice_mux_2 mux_6290(eclk, ereset, dpc1_SBY_v,cclk_v, v(sb3_v),n_1531_v, y3_v);
  spice_mux_2 mux_6291(eclk, ereset, dpc1_SBY_v,cclk_v, v(sb2_v),n_1491_v, y2_v);
  spice_mux_2 mux_6359(eclk, ereset, dor4_v,(n_1463_v|RnWstretched_v), 1'b1,1'b0, n_1076_v);
  spice_mux_2 mux_6358(eclk, ereset, (cp1_v&fetch_v),cclk_v, n_1309_v,notir6_v, n_1675_v);
  spice_mux_2 mux_6357(eclk, ereset, n_358_v,n_1129_v, 1'b1,1'b0, n_1467_v);
  spice_mux_2 mux_6356(eclk, ereset, dpc23_SBAC_v,cclk_v, dasb7_v,n_1592_v, a7_v);
  spice_mux_2 mux_6355(eclk, ereset, cclk_v,dpc23_SBAC_v, n_1344_v,v(sb4_v), a4_v);
  spice_mux_2 mux_6353(eclk, ereset, cclk_v,dpc23_SBAC_v, n_1618_v,dasb2_v, a2_v);
  spice_mux_2 mux_6352(eclk, ereset, cclk_v,dpc23_SBAC_v, n_146_v,v(sb0_v), a0_v);
  spice_mux_2 mux_6351(eclk, ereset, cclk_v,dpc23_SBAC_v, n_929_v,dasb1_v, a1_v);
  spice_mux_2 mux_6350(eclk, ereset, n_1566_v,n_1240_v, 1'b1,1'b0, dpc43_DL_DB_v);
  spice_mux_3 mux_6374(eclk, ereset, dpc9_DBADD_v,dpc8_nDBADD_v,dpc10_ADLADD_v, v(idb6_v),n_351_v,v(adl6_v), alub6_v);
  spice_mux_3 mux_6371(eclk, ereset, dpc8_nDBADD_v,dpc9_DBADD_v,dpc10_ADLADD_v, n_583_v,v(idb1_v),v(adl1_v), alub1_v);
  spice_mux_3 mux_6370(eclk, ereset, dpc8_nDBADD_v,dpc9_DBADD_v,dpc10_ADLADD_v, n_1621_v,v(idb3_v),v(adl3_v), alub3_v);
  spice_mux_3 mux_6373(eclk, ereset, dpc8_nDBADD_v,dpc9_DBADD_v,dpc10_ADLADD_v, n_423_v,v(idb7_v),v(adl7_v), alub7_v);
  spice_mux_3 mux_6372(eclk, ereset, dpc10_ADLADD_v,dpc9_DBADD_v,dpc8_nDBADD_v, v(adl0_v),v(idb0_v),n_624_v, alub0_v);
  spice_mux_2 mux_6379(eclk, ereset, cclk_v,(ADH_ABH_v&cp1_v), n_994_v,n_168_v, _ABH2_v);
  spice_mux_2 mux_6378(eclk, ereset, n_1026_v,n_567_v, 1'b1,1'b0, n_171_v);
  spice_mux_2 mux_6230(eclk, ereset, (cp1_v&fetch_v),cclk_v, n_1605_v,notir7_v, n_541_v);
  spice_mux_2 mux_6231(eclk, ereset, n_1026_v,n_567_v, 1'b0,1'b1, n_322_v);
  spice_mux_2 mux_6232(eclk, ereset, n_628_v,(n_1247_v|n_1335_v|cclk_v), 1'b1,1'b0, dpc24_ACSB_v);
  spice_mux_2 mux_6233(eclk, ereset, dor2_v,(RnWstretched_v|n_224_v), 1'b1,1'b0, n_520_v);
  spice_mux_2 mux_6234(eclk, ereset, n_1033_v,n_241_v, 1'b0,1'b1, dpc21_ADDADL_v);
  spice_mux_2 mux_6235(eclk, ereset, n_224_v,(dor2_v|RnWstretched_v), 1'b1,1'b0, n_37_v);
  spice_mux_2 mux_6236(eclk, ereset, n_1417_v,n_747_v, 1'b0,1'b1, clk1out_v);
  spice_mux_2 mux_6237(eclk, ereset, n_17_v,(n_732_v|n_964_v), 1'b1,1'b0, clock1_v);
  spice_mux_2 mux_6238(eclk, ereset, n_1413_v,n_1260_v, 1'b0,1'b1, dpc32_PCHADH_v);
  spice_mux_2 mux_6239(eclk, ereset, n_747_v,n_670_v, 1'b0,1'b1, n_1417_v);
  spice_mux_2 mux_6216(eclk, ereset, cclk_v,dpc23_SBAC_v, n_1654_v,dasb3_v, a3_v);
  spice_mux_2 mux_6217(eclk, ereset, dpc23_SBAC_v,cclk_v, dasb6_v,n_326_v, a6_v);
  spice_mux_2 mux_6214(eclk, ereset, (cp1_v&fetch_v),cclk_v, n_1641_v,notir1_v, n_119_v);
  spice_mux_2 mux_6215(eclk, ereset, n_1399_v,n_1105_v, 1'b1,1'b0, cp1_v);
  spice_mux_2 mux_6212(eclk, ereset, n_951_v,abl2_v, 1'b1,1'b0, n_642_v);
  spice_mux_2 mux_6213(eclk, ereset, n_1613_v,(dor3_v|RnWstretched_v), 1'b1,1'b0, n_643_v);
  spice_mux_2 mux_6210(eclk, ereset, n_1271_v,n_1596_v, 1'b0,1'b1, dpc27_SBADH_v);
  spice_mux_2 mux_6211(eclk, ereset, abl3_v,n_990_v, 1'b0,1'b1, n_138_v);
  spice_mux_2 mux_6218(eclk, ereset, abl1_v,n_842_v, 1'b1,1'b0, n_1479_v);
  spice_mux_2 mux_6219(eclk, ereset, n_445_v,n_417_v, 1'b0,1'b1, sync_v);
  spice_mux_2 mux_6278(eclk, ereset, dpc11_SBADD_v,dpc12_0ADD_v, v(sb5_v),1'b0, alua5_v);
  spice_mux_2 mux_6226(eclk, ereset, n_659_v,n_1639_v, 1'b0,1'b1, ab15_v);
  spice_mux_2 mux_6276(eclk, ereset, dpc11_SBADD_v,dpc12_0ADD_v, v(sb7_v),1'b0, alua7_v);
  spice_mux_2 mux_6277(eclk, ereset, dpc11_SBADD_v,dpc12_0ADD_v, v(sb4_v),1'b0, alua4_v);
  spice_mux_2 mux_6270(eclk, ereset, dpc39_PCLPCL_v,dpc40_ADLPCL_v, n_1647_v,v(adl7_v), pcl7_v);
  spice_mux_2 mux_6271(eclk, ereset, dpc40_ADLPCL_v,dpc39_PCLPCL_v, v(adl6_v),n_1458_v, pcl6_v);
  spice_mux_2 mux_6273(eclk, ereset, dpc40_ADLPCL_v,dpc39_PCLPCL_v, v(adl4_v),n_208_v, pcl4_v);
  spice_mux_2 mux_6321(eclk, ereset, n_834_v,n_400_v, 1'b1,1'b0, n_102_v);
  spice_mux_2 mux_6328(eclk, ereset, n_1100_v,n_855_v, 1'b0,1'b1, ab0_v);
  spice_mux_2 mux_6329(eclk, ereset, n_66_v,n_1479_v, 1'b0,1'b1, ab1_v);
  spice_mux_2 mux_6252(eclk, ereset, n_1423_v,abh5_v, 1'b0,1'b1, n_1608_v);
  spice_mux_2 mux_6250(eclk, ereset, dpc31_PCHPCH_v,dpc30_ADHPCH_v, n_1722_v,v(adh0_v), pch0_v);
  spice_mux_2 mux_6251(eclk, ereset, n_531_v,n_1255_v, 1'b1,1'b0, dpc13_ORS_v);
  spice_mux_2 mux_6256(eclk, ereset, abl3_v,n_990_v, 1'b1,1'b0, n_1041_v);
  spice_mux_2 mux_6257(eclk, ereset, (cp1_v&fetch_v),cclk_v, n_1083_v,notir3_v, n_1620_v);
  spice_mux_2 mux_6254(eclk, ereset, n_1346_v,abh3_v, 1'b0,1'b1, n_1296_v);
  spice_mux_2 mux_6258(eclk, ereset, cclk_v,dpc3_SBX_v, n_1694_v,v(sb2_v), x2_v);
  spice_mux_2 mux_6199(eclk, ereset, n_1660_v,abl0_v, 1'b1,1'b0, n_1100_v);
  spice_mux_2 mux_6198(eclk, ereset, n_1399_v,n_1715_v, 1'b0,1'b1, n_1105_v);
  spice_mux_2 mux_6195(eclk, ereset, cclk_v,dpc3_SBX_v, n_1724_v,v(sb6_v), x6_v);
  spice_mux_2 mux_6194(eclk, ereset, n_154_v,n_75_v, 1'b1,1'b0, dpc20_ADDSB06_v);
  spice_mux_2 mux_6197(eclk, ereset, (ADL_ABL_v&cp1_v),cclk_v, n_1519_v,n_86_v, _ABL4_v);
  spice_mux_2 mux_6196(eclk, ereset, dor6_v,(n_466_v|RnWstretched_v), 1'b1,1'b0, n_7_v);
  spice_mux_2 mux_6191(eclk, ereset, cclk_v,(ADL_ABL_v&cp1_v), n_1100_v,n_123_v, _ABL0_v);
  spice_mux_2 mux_6190(eclk, ereset, cclk_v,(cp1_v&ADL_ABL_v), n_66_v,n_1016_v, _ABL1_v);
  spice_mux_2 mux_6193(eclk, ereset, n_102_v,n_1696_v, 1'b1,1'b0, rw_v);
  spice_mux_2 mux_6192(eclk, ereset, n_543_v,n_196_v, 1'b1,1'b0, dpc5_SADL_v);
  spice_mux_2 mux_6388(eclk, ereset, n_23_v,(dor7_v|RnWstretched_v), 1'b1,1'b0, n_1501_v);
  spice_mux_2 mux_6389(eclk, ereset, dor7_v,(n_23_v|RnWstretched_v), 1'b1,1'b0, n_298_v);
  spice_mux_2 mux_6380(eclk, ereset, cclk_v,(cp1_v&ADH_ABH_v), n_999_v,n_212_v, _ABH4_v);
  spice_mux_2 mux_6381(eclk, ereset, abl6_v,n_1195_v, 1'b0,1'b1, n_1254_v);
  spice_mux_2 mux_6382(eclk, ereset, n_709_v,n_1499_v, 1'b0,1'b1, dpc18__DAA_v);
  spice_mux_2 mux_6383(eclk, ereset, n_1462_v,n_1369_v, 1'b0,1'b1, dpc38_PCLADL_v);
  spice_mux_2 mux_6384(eclk, ereset, n_400_v,n_834_v, 1'b1,1'b0, n_1696_v);
  spice_mux_2 mux_6385(eclk, ereset, n_1660_v,abl0_v, 1'b0,1'b1, n_855_v);
  spice_mux_2 mux_6386(eclk, ereset, n_1034_v,abh2_v, 1'b1,1'b0, n_994_v);
  spice_mux_2 mux_6387(eclk, ereset, abh4_v,n_1677_v, 1'b0,1'b1, n_999_v);
  spice_mux_2 mux_6201(eclk, ereset, dpc6_SBS_v,dpc7_SS_v, v(sb3_v),n_998_v, s3_v);
  spice_mux_2 mux_6203(eclk, ereset, dpc6_SBS_v,dpc7_SS_v, v(sb1_v),n_694_v, s1_v);
  spice_mux_2 mux_6202(eclk, ereset, dpc6_SBS_v,dpc7_SS_v, v(sb2_v),n_1389_v, s2_v);
  spice_mux_2 mux_6207(eclk, ereset, dpc6_SBS_v,dpc7_SS_v, v(sb5_v),n_280_v, s5_v);
  spice_mux_2 mux_6206(eclk, ereset, dpc6_SBS_v,dpc7_SS_v, v(sb6_v),n_618_v, s6_v);
  spice_mux_2 mux_6293(eclk, ereset, cclk_v,dpc1_SBY_v, n_658_v,v(sb4_v), y4_v);
  spice_mux_3 mux_6300(eclk, ereset, n_850_v,n_771_v,n_1446_v, 1'b0,n_465_v,n_206_v, n_430_v);
  spice_mux_3 mux_6301(eclk, ereset, cclk_v,n_1523_v,abh6_v, v(_ABH6_v),1'b1,1'b0, n_635_v);
  spice_mux_2 mux_6303(eclk, ereset, n_108_v,n_1364_v, 1'b0,1'b1, dpc16_EORS_v);
  spice_mux_2 mux_6304(eclk, ereset, n_1720_v,(dor5_v|RnWstretched_v), 1'b1,1'b0, n_612_v);
  spice_mux_2 mux_6305(eclk, ereset, n_1034_v,abh2_v, 1'b0,1'b1, n_1545_v);
  spice_mux_2 mux_6306(eclk, ereset, n_906_v,n_714_v, 1'b0,1'b1, dpc19_ADDSB7_v);
  spice_mux_2 mux_6307(eclk, ereset, abh4_v,n_1677_v, 1'b1,1'b0, n_475_v);
  spice_mux_2 mux_6308(eclk, ereset, n_466_v,(dor6_v|RnWstretched_v), 1'b1,1'b0, n_471_v);
  spice_mux_2 mux_6309(eclk, ereset, n_127_v,n_519_v, 1'b0,1'b1, n_135_v);
  spice_mux_2 mux_6326(eclk, ereset, n_951_v,abl2_v, 1'b0,1'b1, n_1152_v);
  spice_mux_2 mux_6327(eclk, ereset, dor5_v,(RnWstretched_v|n_1720_v), 1'b1,1'b0, n_373_v);
  spice_mux_2 mux_6324(eclk, ereset, n_1295_v,n_1238_v, 1'b1,1'b0, dpc25_SBDB_v);
  spice_mux_2 mux_6325(eclk, ereset, n_830_v,(n_1047_v|cclk_v|n_1247_v), 1'b1,1'b0, dpc23_SBAC_v);
  spice_mux_2 mux_6322(eclk, ereset, n_1270_v,(cclk_v|n_1247_v|n_1518_v), 1'b1,1'b0, dpc39_PCLPCL_v);
  spice_mux_2 mux_6323(eclk, ereset, n_1067_v,n_582_v, 1'b0,1'b1, ADH_ABH_v);
  spice_mux_2 mux_6320(eclk, ereset, n_1534_v,(n_763_v|cclk_v|n_1247_v), 1'b1,1'b0, dpc8_nDBADD_v);
  spice_mux_2 mux_6274(eclk, ereset, n_161_v,(n_969_v|n_1247_v|cclk_v), 1'b1,1'b0, dpc0_YSB_v);
  spice_mux_2 mux_6275(eclk, ereset, dpc11_SBADD_v,dpc12_0ADD_v, v(sb6_v),1'b0, alua6_v);
  spice_mux_2 mux_6272(eclk, ereset, dpc40_ADLPCL_v,dpc39_PCLPCL_v, v(adl5_v),n_72_v, pcl5_v);
  spice_mux_2 mux_6200(eclk, ereset, n_6_v,(n_1247_v|n_282_v|cclk_v), 1'b1,1'b0, dpc6_SBS_v);
  spice_mux_2 mux_6205(eclk, ereset, dpc6_SBS_v,dpc7_SS_v, v(sb7_v),n_721_v, s7_v);
  spice_mux_2 mux_6204(eclk, ereset, dpc7_SS_v,dpc6_SBS_v, n_332_v,v(sb0_v), s0_v);
  spice_mux_2 mux_6348(eclk, ereset, n_818_v,(cclk_v|n_1043_v|n_1247_v), 1'b1,1'b0, dpc40_ADLPCL_v);
  spice_mux_2 mux_6349(eclk, ereset, n_21_v,(n_228_v|n_1247_v|cclk_v), 1'b1,1'b0, dpc30_ADHPCH_v);
  spice_mux_2 mux_6344(eclk, ereset, n_220_v,n_130_v, 1'b1,1'b0, ADL_ABL_v);
  spice_mux_2 mux_6345(eclk, ereset, abl6_v,n_1195_v, 1'b1,1'b0, n_1191_v);
  spice_mux_2 mux_6346(eclk, ereset, n_839_v,cp1_v, 1'b1,1'b0, n_43_v);
  spice_mux_2 mux_6347(eclk, ereset, dor3_v,(n_1613_v|RnWstretched_v), 1'b1,1'b0, n_42_v);
  spice_mux_2 mux_6340(eclk, ereset, (cp1_v&fetch_v),cclk_v, n_409_v,notir0_v, n_310_v);
  spice_mux_2 mux_6341(eclk, ereset, n_1552_v,n_1593_v, 1'b0,1'b1, dpc14_SRS_v);
  spice_mux_2 mux_6342(eclk, ereset, n_842_v,abl1_v, 1'b1,1'b0, n_66_v);
  spice_mux_2 mux_6343(eclk, ereset, n_1463_v,(dor4_v|RnWstretched_v), 1'b1,1'b0, n_147_v);

  spice_node_4 n_n_1387(eclk, ereset, n_1387_port_2,n_1387_port_3,n_1387_port_0,n_1387_port_1, n_1387_v);
  spice_node_1 n_irq(eclk, ereset, irq_port_2, irq_v);
  spice_node_2 n_so(eclk, ereset, so_port_2,so_port_3, so_v);
  spice_node_5 n_n_304(eclk, ereset, n_304_port_2,n_304_port_3,n_304_port_0,n_304_port_1,n_304_port_4, n_304_v);
  spice_node_2 n_n_330(eclk, ereset, n_330_port_7,n_330_port_4, n_330_v);
  spice_node_2 n_rdy(eclk, ereset, rdy_port_2,rdy_port_3, rdy_v);
  spice_node_3 n_db1(eclk, ereset, db1_port_1,db1_port_4,db1_port_5, db1_v);
  spice_node_3 n_db0(eclk, ereset, db0_port_1,db0_port_4,db0_port_5, db0_v);
  spice_node_3 n_db3(eclk, ereset, db3_port_2,db3_port_3,db3_port_5, db3_v);
  spice_node_3 n_db2(eclk, ereset, db2_port_2,db2_port_3,db2_port_5, db2_v);
  spice_node_3 n_db5(eclk, ereset, db5_port_0,db5_port_4,db5_port_5, db5_v);
  spice_node_3 n_db4(eclk, ereset, db4_port_3,db4_port_0,db4_port_5, db4_v);
  spice_node_3 n_db7(eclk, ereset, db7_port_3,db7_port_1,db7_port_5, db7_v);
  spice_node_3 n_db6(eclk, ereset, db6_port_0,db6_port_4,db6_port_5, db6_v);
  spice_node_4 n_n_1661(eclk, ereset, n_1661_port_2,n_1661_port_3,n_1661_port_0,n_1661_port_1, n_1661_v);
  spice_node_7 n_idb1(eclk, ereset, idb1_port_8,idb1_port_9,idb1_port_3,idb1_port_0,idb1_port_4,idb1_port_5,idb1_port_10, idb1_v);
  spice_node_7 n_idb0(eclk, ereset, idb0_port_8,idb0_port_2,idb0_port_1,idb0_port_6,idb0_port_7,idb0_port_5,idb0_port_10, idb0_v);
  spice_node_7 n_idb3(eclk, ereset, idb3_port_9,idb3_port_3,idb3_port_0,idb3_port_1,idb3_port_6,idb3_port_5,idb3_port_10, idb3_v);
  spice_node_7 n_idb2(eclk, ereset, idb2_port_3,idb2_port_0,idb2_port_1,idb2_port_6,idb2_port_4,idb2_port_5,idb2_port_10, idb2_v);
  spice_node_6 n_idb5(eclk, ereset, idb5_port_9,idb5_port_2,idb5_port_6,idb5_port_7,idb5_port_4,idb5_port_5, idb5_v);
  spice_node_7 n_idb4(eclk, ereset, idb4_port_9,idb4_port_0,idb4_port_6,idb4_port_7,idb4_port_4,idb4_port_5,idb4_port_10, idb4_v);
  spice_node_7 n_idb7(eclk, ereset, idb7_port_9,idb7_port_2,idb7_port_3,idb7_port_0,idb7_port_7,idb7_port_4,idb7_port_10, idb7_v);
  spice_node_7 n_idb6(eclk, ereset, idb6_port_9,idb6_port_3,idb6_port_0,idb6_port_6,idb6_port_7,idb6_port_5,idb6_port_11, idb6_v);
  spice_node_4 n_n_719(eclk, ereset, n_719_port_2,n_719_port_3,n_719_port_0,n_719_port_1, n_719_v);
  spice_node_1 n_nmi(eclk, ereset, nmi_port_2, nmi_v);
  spice_node_1 n_n_633(eclk, ereset, n_633_port_0, n_633_v);
  spice_node_0 n_n_866(eclk, ereset,  n_866_v);
  spice_node_0 n_n_806(eclk, ereset,  n_806_v);
  spice_node_2 n_n_807(eclk, ereset, n_807_port_3,n_807_port_5, n_807_v);
  spice_node_4 n_n_87(eclk, ereset, n_87_port_2,n_87_port_3,n_87_port_0,n_87_port_1, n_87_v);
  spice_node_8 n_sb2(eclk, ereset, sb2_port_8,sb2_port_9,sb2_port_3,sb2_port_1,sb2_port_7,sb2_port_10,sb2_port_11,sb2_port_12, sb2_v);
  spice_node_8 n_sb3(eclk, ereset, sb3_port_9,sb3_port_3,sb3_port_1,sb3_port_7,sb3_port_4,sb3_port_5,sb3_port_10,sb3_port_11, sb3_v);
  spice_node_8 n_sb0(eclk, ereset, sb0_port_9,sb0_port_2,sb0_port_1,sb0_port_6,sb0_port_4,sb0_port_10,sb0_port_11,sb0_port_12, sb0_v);
  spice_node_8 n_sb1(eclk, ereset, sb1_port_8,sb1_port_9,sb1_port_2,sb1_port_6,sb1_port_7,sb1_port_10,sb1_port_11,sb1_port_12, sb1_v);
  spice_node_8 n_sb6(eclk, ereset, sb6_port_8,sb6_port_9,sb6_port_2,sb6_port_6,sb6_port_4,sb6_port_10,sb6_port_11,sb6_port_12, sb6_v);
  spice_node_8 n_sb7(eclk, ereset, sb7_port_8,sb7_port_9,sb7_port_3,sb7_port_0,sb7_port_1,sb7_port_6,sb7_port_7,sb7_port_5, sb7_v);
  spice_node_8 n_sb4(eclk, ereset, sb4_port_8,sb4_port_9,sb4_port_3,sb4_port_0,sb4_port_5,sb4_port_10,sb4_port_11,sb4_port_12, sb4_v);
  spice_node_8 n_sb5(eclk, ereset, sb5_port_8,sb5_port_2,sb5_port_3,sb5_port_6,sb5_port_7,sb5_port_10,sb5_port_11,sb5_port_12, sb5_v);
  spice_node_1 n_res(eclk, ereset, res_port_2, res_v);
  spice_node_5 n_adl7(eclk, ereset, adl7_port_2,adl7_port_3,adl7_port_0,adl7_port_7,adl7_port_5, adl7_v);
  spice_node_5 n_adl6(eclk, ereset, adl6_port_2,adl6_port_3,adl6_port_1,adl6_port_4,adl6_port_5, adl6_v);
  spice_node_5 n_adl5(eclk, ereset, adl5_port_2,adl5_port_3,adl5_port_0,adl5_port_1,adl5_port_4, adl5_v);
  spice_node_5 n_adl4(eclk, ereset, adl4_port_3,adl4_port_0,adl4_port_1,adl4_port_4,adl4_port_5, adl4_v);
  spice_node_5 n_adl3(eclk, ereset, adl3_port_2,adl3_port_3,adl3_port_0,adl3_port_1,adl3_port_4, adl3_v);
  spice_node_6 n_adl2(eclk, ereset, adl2_port_2,adl2_port_3,adl2_port_0,adl2_port_6,adl2_port_4,adl2_port_5, adl2_v);
  spice_node_6 n_adl1(eclk, ereset, adl1_port_2,adl1_port_3,adl1_port_0,adl1_port_1,adl1_port_4,adl1_port_5, adl1_v);
  spice_node_6 n_adl0(eclk, ereset, adl0_port_3,adl0_port_0,adl0_port_6,adl0_port_7,adl0_port_4,adl0_port_5, adl0_v);
  spice_node_4 n_n_1014(eclk, ereset, n_1014_port_2,n_1014_port_3,n_1014_port_0,n_1014_port_1, n_1014_v);
  spice_node_4 n_n_1424(eclk, ereset, n_1424_port_2,n_1424_port_3,n_1424_port_0,n_1424_port_1, n_1424_v);
  spice_node_5 n_notaluoutmux0(eclk, ereset, notaluoutmux0_port_2,notaluoutmux0_port_3,notaluoutmux0_port_0,notaluoutmux0_port_1,notaluoutmux0_port_5, notaluoutmux0_v);
  spice_node_5 n_notaluoutmux1(eclk, ereset, notaluoutmux1_port_2,notaluoutmux1_port_0,notaluoutmux1_port_1,notaluoutmux1_port_4,notaluoutmux1_port_5, notaluoutmux1_v);
  spice_node_5 n_n_277(eclk, ereset, n_277_port_2,n_277_port_3,n_277_port_1,n_277_port_4,n_277_port_5, n_277_v);
  spice_node_4 n_n_1095(eclk, ereset, n_1095_port_2,n_1095_port_3,n_1095_port_0,n_1095_port_1, n_1095_v);
  spice_node_5 n_adh3(eclk, ereset, adh3_port_3,adh3_port_0,adh3_port_6,adh3_port_4,adh3_port_5, adh3_v);
  spice_node_5 n_adh2(eclk, ereset, adh2_port_3,adh2_port_0,adh2_port_6,adh2_port_4,adh2_port_5, adh2_v);
  spice_node_5 n_adh1(eclk, ereset, adh1_port_2,adh1_port_0,adh1_port_1,adh1_port_6,adh1_port_4, adh1_v);
  spice_node_5 n_adh0(eclk, ereset, adh0_port_2,adh0_port_3,adh0_port_0,adh0_port_1,adh0_port_6, adh0_v);
  spice_node_5 n_adh7(eclk, ereset, adh7_port_2,adh7_port_3,adh7_port_0,adh7_port_4,adh7_port_5, adh7_v);
  spice_node_5 n_adh6(eclk, ereset, adh6_port_3,adh6_port_0,adh6_port_6,adh6_port_4,adh6_port_5, adh6_v);
  spice_node_5 n_adh5(eclk, ereset, adh5_port_2,adh5_port_3,adh5_port_0,adh5_port_4,adh5_port_5, adh5_v);
  spice_node_5 n_adh4(eclk, ereset, adh4_port_2,adh4_port_0,adh4_port_6,adh4_port_4,adh4_port_5, adh4_v);
  spice_node_2 n_NMIP(eclk, ereset, NMIP_port_7,NMIP_port_4, NMIP_v);
  spice_node_5 n_n_1071(eclk, ereset, n_1071_port_2,n_1071_port_3,n_1071_port_0,n_1071_port_4,n_1071_port_5, n_1071_v);
  spice_node_4 n_n_1147(eclk, ereset, n_1147_port_2,n_1147_port_3,n_1147_port_0,n_1147_port_1, n_1147_v);
  spice_node_5 n_n_722(eclk, ereset, n_722_port_2,n_722_port_0,n_722_port_1,n_722_port_4,n_722_port_5, n_722_v);
  spice_node_1 n_n_1059(eclk, ereset, n_1059_port_0, n_1059_v);
  spice_node_5 n_n_740(eclk, ereset, n_740_port_2,n_740_port_3,n_740_port_0,n_740_port_1,n_740_port_4, n_740_v);
  spice_node_2 n_n_975(eclk, ereset, n_975_port_3,n_975_port_6, n_975_v);
  spice_node_1 n_clk0(eclk, ereset, clk0_port_3, clk0_v);
  spice_node_1 n__ABH3(eclk, ereset, _ABH3_port_3, _ABH3_v);
  spice_node_1 n__ABH1(eclk, ereset, _ABH1_port_3, _ABH1_v);
  spice_node_1 n__ABH0(eclk, ereset, _ABH0_port_3, _ABH0_v);
  spice_node_1 n__ABH7(eclk, ereset, _ABH7_port_3, _ABH7_v);
  spice_node_1 n__ABH6(eclk, ereset, _ABH6_port_3, _ABH6_v);
  spice_node_1 n__ABH5(eclk, ereset, _ABH5_port_3, _ABH5_v);
  spice_node_2 n_n_854(eclk, ereset, n_854_port_6,n_854_port_4, n_854_v);
  spice_node_2 n_n_297(eclk, ereset, n_297_port_3,n_297_port_5, n_297_v);
  spice_node_5 n_n_296(eclk, ereset, n_296_port_3,n_296_port_0,n_296_port_1,n_296_port_4,n_296_port_5, n_296_v);

endmodule

module spice_node_0(input eclk,ereset, output signed [`W-1:0] v);
  assign v = 0;
endmodule

module spice_node_1(input eclk,ereset, input signed [`W-1:0] i0, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_2(input eclk,ereset, input signed [`W-1:0] i0,i1, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_3(input eclk,ereset, input signed [`W-1:0] i0,i1,i2, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_4(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_5(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_6(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_7(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_8(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6,i7, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6+i7;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_mux_2(input eclk,ereset, input clk0,clk1, input x0,x1, output reg y);
  wire c0,z0;
  wire c1,z1;

  assign c0 = clk0;
  assign z0 = x0;

  mux_cascade m0(c0, z0, clk1, x1, c1, z1);

  wire clk = c1;
  wire x = z1;

  always @(posedge eclk)
    if (ereset)
      y <= 0;
    else begin
      if (clk)
        y <= x;
    end

endmodule

module spice_mux_3(input eclk,ereset, input clk0,clk1,clk2, input x0,x1,x2, output reg y);
  wire c0,z0;
  wire c1,z1;
  wire c2,z2;

  assign c0 = clk0;
  assign z0 = x0;

  mux_cascade m0(c0, z0, clk1, x1, c1, z1);
  mux_cascade m1(c1, z1, clk2, x2, c2, z2);

  wire clk = c2;
  wire x = z2;

  always @(posedge eclk)
    if (ereset)
      y <= 0;
    else begin
      if (clk)
        y <= x;
    end

endmodule

