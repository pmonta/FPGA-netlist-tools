* SPICE3 file created from 4003.ext - technology: nmos

.option scale=0.001u

M1000 Vdd Vdd diff_258130_451520# GND efet w=10790 l=9960
+ ad=-1.73615e+09 pd=5.68882e+06 as=-1.17478e+08 ps=665660 
M1001 Vdd Vdd Vdd GND efet w=2075 l=5395
+ ad=0 pd=0 as=0 ps=0 
M1002 Vdd Vdd Vdd GND efet w=2905 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1003 Vdd Vdd diff_1540480_996000# GND efet w=6640 l=143590
+ ad=0 pd=0 as=4.1334e+08 ps=112880 
M1004 diff_1540480_996000# diff_232400_451520# GND GND efet w=14940 l=7470
+ ad=0 pd=0 as=-3.63212e+08 ps=1.71777e+07 
M1005 GND diff_1466610_1008450# diff_258130_451520# GND efet w=247340 l=14110
+ ad=0 pd=0 as=0 ps=0 
M1006 Vdd Vdd diff_1466610_1008450# GND efet w=6640 l=146080
+ ad=0 pd=0 as=2.14179e+09 ps=353580 
M1007 diff_1466610_1008450# diff_1540480_996000# GND GND efet w=174300 l=22410
+ ad=0 pd=0 as=0 ps=0 
M1008 GND diff_273900_560250# diff_232400_451520# GND efet w=150230 l=7470
+ ad=0 pd=0 as=9.35161e+08 ps=811740 
M1009 diff_273900_560250# diff_232400_451520# GND GND efet w=61420 l=7470
+ ad=-1.96855e+09 pd=463140 as=0 ps=0 
M1010 q4 diff_404210_938730# GND GND efet w=351505 l=7885
+ ad=6.85091e+08 pd=833320 as=0 ps=0 
M1011 GND diff_312080_771900# diff_296310_846600# GND efet w=66815 l=7885
+ ad=0 pd=0 as=1.77805e+09 ps=328680 
M1012 diff_296310_846600# diff_207500_451520# GND GND efet w=37765 l=7885
+ ad=0 pd=0 as=0 ps=0 
M1013 diff_296310_846600# diff_296310_846600# diff_296310_846600# GND efet w=2490 l=2490
+ ad=0 pd=0 as=0 ps=0 
M1014 diff_296310_846600# diff_296310_846600# diff_296310_846600# GND efet w=1660 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1015 diff_312080_771900# diff_312080_771900# diff_312080_771900# GND efet w=3320 l=3320
+ ad=9.44482e+08 pd=215800 as=0 ps=0 
M1016 diff_312080_771900# diff_312080_771900# diff_312080_771900# GND efet w=1660 l=4980
+ ad=0 pd=0 as=0 ps=0 
M1017 diff_296310_846600# Vdd Vdd GND efet w=8300 l=24900
+ ad=0 pd=0 as=0 ps=0 
M1018 Vdd Vdd Vdd GND efet w=2075 l=7055
+ ad=0 pd=0 as=0 ps=0 
M1019 Vdd Vdd Vdd GND efet w=3320 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1020 q3 diff_644910_939560# GND GND efet w=350260 l=7470
+ ad=8.22182e+08 pd=830000 as=0 ps=0 
M1021 GND diff_551950_771900# diff_536180_846600# GND efet w=67645 l=7885
+ ad=0 pd=0 as=1.83454e+09 ps=333660 
M1022 diff_536180_846600# diff_207500_451520# GND GND efet w=39010 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1023 diff_536180_846600# diff_536180_846600# diff_536180_846600# GND efet w=2905 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1024 diff_536180_846600# diff_536180_846600# diff_536180_846600# GND efet w=2490 l=4150
+ ad=0 pd=0 as=0 ps=0 
M1025 diff_404210_938730# diff_296310_846600# GND GND efet w=54780 l=7470
+ ad=6.94411e+08 pd=167660 as=0 ps=0 
M1026 diff_404210_938730# diff_404210_938730# diff_404210_938730# GND efet w=2905 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1027 diff_404210_938730# diff_404210_938730# diff_404210_938730# GND efet w=2075 l=5395
+ ad=0 pd=0 as=0 ps=0 
M1028 diff_551950_771900# diff_551950_771900# diff_551950_771900# GND efet w=2490 l=2490
+ ad=1.01819e+09 pd=217460 as=0 ps=0 
M1029 diff_551950_771900# diff_551950_771900# diff_551950_771900# GND efet w=2075 l=4150
+ ad=0 pd=0 as=0 ps=0 
M1030 q4 diff_296310_846600# Vdd GND efet w=24900 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1031 diff_404210_938730# Vdd Vdd GND efet w=9960 l=19920
+ ad=0 pd=0 as=0 ps=0 
M1032 diff_536180_846600# Vdd Vdd GND efet w=8300 l=24070
+ ad=0 pd=0 as=0 ps=0 
M1033 Vdd Vdd Vdd GND efet w=2075 l=6225
+ ad=0 pd=0 as=0 ps=0 
M1034 Vdd Vdd Vdd GND efet w=4150 l=4150
+ ad=0 pd=0 as=0 ps=0 
M1035 Vdd Vdd Vdd GND efet w=2075 l=7055
+ ad=0 pd=0 as=0 ps=0 
M1036 Vdd Vdd Vdd GND efet w=3320 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1037 Vdd Vdd Vdd GND efet w=2075 l=6225
+ ad=0 pd=0 as=0 ps=0 
M1038 Vdd Vdd Vdd GND efet w=3320 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1039 diff_312080_771900# diff_258130_451520# diff_278050_567720# GND efet w=14110 l=8300
+ ad=0 pd=0 as=1.79252e+09 ps=345280 
M1040 diff_292990_681430# diff_258130_451520# diff_278050_567720# GND efet w=14110 l=7470
+ ad=2.03914e+08 pd=64740 as=0 ps=0 
M1041 diff_292990_681430# diff_292990_681430# diff_292990_681430# GND efet w=2905 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1042 diff_292990_681430# diff_292990_681430# diff_292990_681430# GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1043 diff_278050_567720# diff_273900_607560# GND GND efet w=21995 l=7885
+ ad=0 pd=0 as=0 ps=0 
M1044 Vdd Vdd diff_278050_567720# GND efet w=8300 l=40670
+ ad=0 pd=0 as=0 ps=0 
M1045 q2 diff_884780_939560# GND GND efet w=350260 l=7470
+ ad=8.63516e+08 pd=831660 as=0 ps=0 
M1046 GND diff_792650_771900# diff_776880_846600# GND efet w=68060 l=7470
+ ad=0 pd=0 as=1.84281e+09 ps=335320 
M1047 diff_776880_846600# diff_207500_451520# GND GND efet w=39010 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1048 diff_776880_846600# diff_776880_846600# diff_776880_846600# GND efet w=3320 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1049 diff_776880_846600# diff_776880_846600# diff_776880_846600# GND efet w=2490 l=4150
+ ad=0 pd=0 as=0 ps=0 
M1050 diff_644910_939560# diff_536180_846600# GND GND efet w=54780 l=7470
+ ad=6.86833e+08 pd=166000 as=0 ps=0 
M1051 diff_644910_939560# diff_644910_939560# diff_644910_939560# GND efet w=2905 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1052 diff_644910_939560# diff_644910_939560# diff_644910_939560# GND efet w=2075 l=5395
+ ad=0 pd=0 as=0 ps=0 
M1053 diff_792650_771900# diff_792650_771900# diff_792650_771900# GND efet w=2490 l=3320
+ ad=9.57571e+08 pd=217460 as=0 ps=0 
M1054 diff_792650_771900# diff_792650_771900# diff_792650_771900# GND efet w=2075 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1055 q3 diff_536180_846600# Vdd GND efet w=24070 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1056 diff_644910_939560# Vdd Vdd GND efet w=9960 l=20750
+ ad=0 pd=0 as=0 ps=0 
M1057 diff_776880_846600# Vdd Vdd GND efet w=8300 l=24070
+ ad=0 pd=0 as=0 ps=0 
M1058 Vdd Vdd Vdd GND efet w=2075 l=7055
+ ad=0 pd=0 as=0 ps=0 
M1059 Vdd Vdd Vdd GND efet w=3320 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1060 Vdd Vdd Vdd GND efet w=1660 l=5810
+ ad=0 pd=0 as=0 ps=0 
M1061 Vdd Vdd Vdd GND efet w=3735 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1062 Vdd Vdd Vdd GND efet w=2075 l=7055
+ ad=0 pd=0 as=0 ps=0 
M1063 Vdd Vdd Vdd GND efet w=3320 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1064 diff_551950_771900# diff_258130_451520# diff_510450_712970# GND efet w=14110 l=7470
+ ad=0 pd=0 as=1.7877e+09 ps=345280 
M1065 diff_390930_703840# diff_390930_703840# diff_390930_703840# GND efet w=3735 l=4150
+ ad=2.35604e+08 pd=84660 as=0 ps=0 
M1066 diff_390930_703840# diff_390930_703840# diff_390930_703840# GND efet w=4150 l=4150
+ ad=0 pd=0 as=0 ps=0 
M1067 diff_278050_567720# diff_232400_451520# diff_395080_711310# GND efet w=48970 l=7470
+ ad=0 pd=0 as=6.67544e+08 ps=151060 
M1068 diff_510450_738700# diff_273900_560250# diff_390930_703840# GND efet w=14110 l=7470
+ ad=1.84625e+09 pd=373500 as=0 ps=0 
M1069 diff_510450_738700# diff_510450_738700# diff_510450_738700# GND efet w=2905 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1070 diff_510450_738700# diff_510450_738700# diff_510450_738700# GND efet w=2905 l=4150
+ ad=0 pd=0 as=0 ps=0 
M1071 GND diff_292990_681430# diff_273900_607560# GND efet w=37350 l=7470
+ ad=0 pd=0 as=-1.91275e+09 ps=493020 
M1072 diff_395080_711310# diff_390930_703840# GND GND efet w=78020 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1073 GND diff_390930_685580# diff_395080_673960# GND efet w=78020 l=7470
+ ad=0 pd=0 as=8.28058e+08 ps=182600 
M1074 diff_390930_685580# diff_390930_685580# diff_390930_685580# GND efet w=3735 l=4150
+ ad=2.39737e+08 pd=84660 as=0 ps=0 
M1075 diff_390930_685580# diff_390930_685580# diff_390930_685580# GND efet w=3735 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1076 diff_510450_712970# diff_273900_560250# diff_390930_685580# GND efet w=14110 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1077 diff_532860_681430# diff_258130_451520# diff_510450_712970# GND efet w=14110 l=7470
+ ad=2.03914e+08 pd=64740 as=0 ps=0 
M1078 diff_532860_681430# diff_532860_681430# diff_532860_681430# GND efet w=2905 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1079 diff_532860_681430# diff_532860_681430# diff_532860_681430# GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1080 diff_510450_712970# diff_510450_738700# GND GND efet w=22410 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1081 Vdd Vdd diff_510450_712970# GND efet w=8300 l=39840
+ ad=0 pd=0 as=0 ps=0 
M1082 q1 diff_1125480_939560# GND GND efet w=351090 l=7470
+ ad=9.15183e+08 pd=833320 as=0 ps=0 
M1083 GND diff_1032520_771900# diff_1016750_846600# GND efet w=68060 l=7470
+ ad=0 pd=0 as=1.82972e+09 ps=335320 
M1084 diff_1016750_846600# diff_207500_451520# GND GND efet w=39010 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1085 diff_1016750_846600# diff_1016750_846600# diff_1016750_846600# GND efet w=3320 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1086 diff_1016750_846600# diff_1016750_846600# diff_1016750_846600# GND efet w=2490 l=4150
+ ad=0 pd=0 as=0 ps=0 
M1087 diff_884780_939560# diff_776880_846600# GND GND efet w=54780 l=7470
+ ad=6.86833e+08 pd=166000 as=0 ps=0 
M1088 diff_884780_939560# diff_884780_939560# diff_884780_939560# GND efet w=2905 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1089 diff_884780_939560# diff_884780_939560# diff_884780_939560# GND efet w=2075 l=5395
+ ad=0 pd=0 as=0 ps=0 
M1090 diff_1032520_771900# diff_1032520_771900# diff_1032520_771900# GND efet w=2490 l=2490
+ ad=1.01062e+09 pd=219120 as=0 ps=0 
M1091 diff_1032520_771900# diff_1032520_771900# diff_1032520_771900# GND efet w=2490 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1092 q2 diff_776880_846600# Vdd GND efet w=24900 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1093 diff_884780_939560# Vdd Vdd GND efet w=9960 l=19920
+ ad=0 pd=0 as=0 ps=0 
M1094 diff_1016750_846600# Vdd Vdd GND efet w=8300 l=24070
+ ad=0 pd=0 as=0 ps=0 
M1095 Vdd Vdd Vdd GND efet w=3320 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1096 Vdd Vdd Vdd GND efet w=1660 l=6640
+ ad=0 pd=0 as=0 ps=0 
M1097 Vdd Vdd Vdd GND efet w=2075 l=6225
+ ad=0 pd=0 as=0 ps=0 
M1098 Vdd Vdd Vdd GND efet w=3735 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1099 Vdd Vdd Vdd GND efet w=2075 l=6225
+ ad=0 pd=0 as=0 ps=0 
M1100 Vdd Vdd Vdd GND efet w=3320 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1101 diff_792650_771900# diff_258130_451520# diff_751150_712970# GND efet w=14110 l=7470
+ ad=0 pd=0 as=1.79527e+09 ps=346940 
M1102 diff_630800_705500# diff_630800_705500# diff_630800_705500# GND efet w=3735 l=3735
+ ad=2.30093e+08 pd=81340 as=0 ps=0 
M1103 diff_630800_705500# diff_630800_705500# diff_630800_705500# GND efet w=3735 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1104 diff_510450_712970# diff_232400_451520# diff_634950_712140# GND efet w=49800 l=7470
+ ad=0 pd=0 as=6.5101e+08 ps=151060 
M1105 diff_751150_738700# diff_273900_560250# diff_630800_705500# GND efet w=14110 l=7470
+ ad=1.8683e+09 pd=373500 as=0 ps=0 
M1106 diff_751150_738700# diff_751150_738700# diff_751150_738700# GND efet w=2490 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1107 diff_751150_738700# diff_751150_738700# diff_751150_738700# GND efet w=2905 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1108 diff_395080_673960# diff_232400_451520# diff_273900_607560# GND efet w=48970 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1109 GND diff_341130_652380# diff_273900_607560# GND efet w=27390 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1110 diff_273900_607560# diff_273900_607560# diff_273900_607560# GND efet w=3735 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1111 diff_273900_607560# diff_273900_607560# diff_273900_607560# GND efet w=3735 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1112 diff_273900_607560# Vdd Vdd GND efet w=8300 l=43160
+ ad=0 pd=0 as=0 ps=0 
M1113 GND diff_532860_681430# diff_510450_738700# GND efet w=37350 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1114 diff_634950_712140# diff_630800_705500# GND GND efet w=78020 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1115 GND diff_630800_686410# diff_634950_673960# GND efet w=78850 l=7470
+ ad=0 pd=0 as=8.36325e+08 ps=184260 
M1116 diff_630800_686410# diff_630800_686410# diff_630800_686410# GND efet w=3735 l=3735
+ ad=2.33537e+08 pd=81340 as=0 ps=0 
M1117 diff_630800_686410# diff_630800_686410# diff_630800_686410# GND efet w=3320 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1118 diff_751150_712970# diff_273900_560250# diff_630800_686410# GND efet w=14110 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1119 diff_773560_682260# diff_258130_451520# diff_751150_712970# GND efet w=14110 l=6640
+ ad=2.03914e+08 pd=64740 as=0 ps=0 
M1120 diff_773560_682260# diff_773560_682260# diff_773560_682260# GND efet w=2905 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1121 diff_773560_682260# diff_773560_682260# diff_773560_682260# GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1122 diff_751150_712970# diff_751150_738700# GND GND efet w=22410 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1123 diff_634950_673960# diff_232400_451520# diff_510450_738700# GND efet w=49800 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1124 GND diff_341130_652380# diff_510450_738700# GND efet w=22410 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1125 diff_510450_738700# Vdd Vdd GND efet w=8300 l=42330
+ ad=0 pd=0 as=0 ps=0 
M1126 Vdd Vdd diff_751150_712970# GND efet w=8300 l=39840
+ ad=0 pd=0 as=0 ps=0 
M1127 q0 diff_1365350_939560# GND GND efet w=350260 l=7470
+ ad=8.30449e+08 pd=828340 as=0 ps=0 
M1128 GND diff_1273220_771900# diff_1257450_846600# GND efet w=67645 l=7055
+ ad=0 pd=0 as=1.84074e+09 ps=335320 
M1129 diff_1257450_846600# diff_207500_451520# GND GND efet w=39010 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1130 diff_1257450_846600# diff_1257450_846600# diff_1257450_846600# GND efet w=2905 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1131 diff_1257450_846600# diff_1257450_846600# diff_1257450_846600# GND efet w=2490 l=4150
+ ad=0 pd=0 as=0 ps=0 
M1132 diff_1125480_939560# diff_1016750_846600# GND GND efet w=55195 l=7055
+ ad=7.16456e+08 pd=166000 as=0 ps=0 
M1133 diff_1125480_939560# diff_1125480_939560# diff_1125480_939560# GND efet w=2490 l=2490
+ ad=0 pd=0 as=0 ps=0 
M1134 diff_1125480_939560# diff_1125480_939560# diff_1125480_939560# GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1135 diff_1273220_771900# diff_1273220_771900# diff_1273220_771900# GND efet w=2075 l=2075
+ ad=9.63082e+08 pd=220780 as=0 ps=0 
M1136 diff_1273220_771900# diff_1273220_771900# diff_1273220_771900# GND efet w=3320 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1137 q1 diff_1016750_846600# Vdd GND efet w=24900 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1138 diff_1125480_939560# Vdd Vdd GND efet w=10790 l=19920
+ ad=0 pd=0 as=0 ps=0 
M1139 diff_1257450_846600# Vdd Vdd GND efet w=8300 l=24070
+ ad=0 pd=0 as=0 ps=0 
M1140 Vdd Vdd Vdd GND efet w=3320 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1141 Vdd Vdd Vdd GND efet w=2075 l=5395
+ ad=0 pd=0 as=0 ps=0 
M1142 Vdd Vdd Vdd GND efet w=2075 l=6225
+ ad=0 pd=0 as=0 ps=0 
M1143 Vdd Vdd Vdd GND efet w=2905 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1144 Vdd Vdd Vdd GND efet w=2075 l=7055
+ ad=0 pd=0 as=0 ps=0 
M1145 Vdd Vdd Vdd GND efet w=3320 l=4980
+ ad=0 pd=0 as=0 ps=0 
M1146 diff_1032520_771900# diff_258130_451520# diff_991020_712970# GND efet w=14110 l=7470
+ ad=0 pd=0 as=1.78701e+09 ps=345280 
M1147 diff_871500_704670# diff_871500_704670# diff_871500_704670# GND efet w=3735 l=3735
+ ad=2.30782e+08 pd=81340 as=0 ps=0 
M1148 diff_871500_704670# diff_871500_704670# diff_871500_704670# GND efet w=3735 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1149 diff_751150_712970# diff_232400_451520# diff_875650_712140# GND efet w=48970 l=7470
+ ad=0 pd=0 as=6.4481e+08 ps=149400 
M1150 diff_991020_738700# diff_273900_560250# diff_871500_704670# GND efet w=14110 l=7470
+ ad=1.87932e+09 pd=373500 as=0 ps=0 
M1151 diff_991020_738700# diff_991020_738700# diff_991020_738700# GND efet w=2490 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1152 diff_991020_738700# diff_991020_738700# diff_991020_738700# GND efet w=2905 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1153 GND diff_773560_682260# diff_751150_738700# GND efet w=38180 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1154 diff_875650_712140# diff_871500_704670# GND GND efet w=77190 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1155 GND diff_871500_685580# diff_875650_674790# GND efet w=77605 l=7055
+ ad=0 pd=0 as=8.36325e+08 ps=182600 
M1156 diff_871500_685580# diff_871500_685580# diff_871500_685580# GND efet w=3735 l=4150
+ ad=2.43871e+08 pd=84660 as=0 ps=0 
M1157 diff_871500_685580# diff_871500_685580# diff_871500_685580# GND efet w=3320 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1158 diff_991020_712970# diff_273900_560250# diff_871500_685580# GND efet w=14110 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1159 diff_1013430_682260# diff_258130_451520# diff_991020_712970# GND efet w=14110 l=7470
+ ad=2.03914e+08 pd=64740 as=0 ps=0 
M1160 diff_1013430_682260# diff_1013430_682260# diff_1013430_682260# GND efet w=2905 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1161 diff_1013430_682260# diff_1013430_682260# diff_1013430_682260# GND efet w=2075 l=5395
+ ad=0 pd=0 as=0 ps=0 
M1162 diff_991020_712970# diff_991020_738700# GND GND efet w=22410 l=6640
+ ad=0 pd=0 as=0 ps=0 
M1163 Vdd Vdd diff_991020_712970# GND efet w=8300 l=39840
+ ad=0 pd=0 as=0 ps=0 
M1164 diff_1365350_939560# diff_1257450_846600# GND GND efet w=55610 l=7470
+ ad=7.21278e+08 pd=166000 as=0 ps=0 
M1165 diff_1365350_939560# diff_1365350_939560# diff_1365350_939560# GND efet w=2075 l=2075
+ ad=0 pd=0 as=0 ps=0 
M1166 diff_1365350_939560# diff_1365350_939560# diff_1365350_939560# GND efet w=2075 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1167 q0 diff_1257450_846600# Vdd GND efet w=24900 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1168 diff_1365350_939560# Vdd Vdd GND efet w=10375 l=20335
+ ad=0 pd=0 as=0 ps=0 
M1169 Vdd Vdd Vdd GND efet w=2490 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1170 Vdd Vdd Vdd GND efet w=2075 l=6225
+ ad=0 pd=0 as=0 ps=0 
M1171 Vdd Vdd Vdd GND efet w=2075 l=7055
+ ad=0 pd=0 as=0 ps=0 
M1172 Vdd Vdd Vdd GND efet w=2490 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1173 GND diff_1621820_879800# diff_232400_451520# GND efet w=149400 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1174 GND diff_1505620_931260# diff_273900_560250# GND efet w=64740 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1175 diff_273900_560250# Vdd Vdd GND efet w=10790 l=20750
+ ad=0 pd=0 as=0 ps=0 
M1176 diff_232400_451520# Vdd Vdd GND efet w=10790 l=9960
+ ad=0 pd=0 as=0 ps=0 
M1177 diff_1621820_879800# diff_1621820_879800# diff_1621820_879800# GND efet w=2075 l=6225
+ ad=6.765e+08 pd=132800 as=0 ps=0 
M1178 diff_1621820_879800# diff_1621820_879800# diff_1621820_879800# GND efet w=3320 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1179 diff_1621820_879800# Vdd Vdd GND efet w=8300 l=24070
+ ad=0 pd=0 as=0 ps=0 
M1180 GND diff_1505620_931260# diff_1621820_879800# GND efet w=34030 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1181 Vdd Vdd Vdd GND efet w=2905 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1182 Vdd Vdd Vdd GND efet w=2490 l=6640
+ ad=0 pd=0 as=0 ps=0 
M1183 GND diff_1588620_812570# diff_1505620_931260# GND efet w=34030 l=8300
+ ad=0 pd=0 as=5.16675e+08 ps=112880 
M1184 diff_1588620_812570# diff_1566210_789330# GND GND efet w=170150 l=22410
+ ad=1.09811e+09 pd=194220 as=0 ps=0 
M1185 diff_1273220_771900# diff_258130_451520# diff_1231720_712970# GND efet w=14110 l=7470
+ ad=0 pd=0 as=1.73878e+09 ps=343620 
M1186 diff_1111370_704670# diff_1111370_704670# diff_1111370_704670# GND efet w=3735 l=3735
+ ad=2.33537e+08 pd=81340 as=0 ps=0 
M1187 diff_1111370_704670# diff_1111370_704670# diff_1111370_704670# GND efet w=3320 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1188 diff_991020_712970# diff_232400_451520# diff_1115520_712140# GND efet w=49385 l=7055
+ ad=0 pd=0 as=6.58588e+08 ps=152720 
M1189 diff_1231720_738700# diff_273900_560250# diff_1111370_704670# GND efet w=14110 l=7470
+ ad=1.93236e+09 pd=378480 as=0 ps=0 
M1190 diff_1231720_738700# diff_1231720_738700# diff_1231720_738700# GND efet w=2905 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1191 diff_1231720_738700# diff_1231720_738700# diff_1231720_738700# GND efet w=2905 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1192 diff_875650_674790# diff_232400_451520# diff_751150_738700# GND efet w=49385 l=7055
+ ad=0 pd=0 as=0 ps=0 
M1193 GND diff_341130_652380# diff_751150_738700# GND efet w=22410 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1194 diff_751150_738700# Vdd Vdd GND efet w=8300 l=41500
+ ad=0 pd=0 as=0 ps=0 
M1195 GND diff_1013430_682260# diff_991020_738700# GND efet w=38180 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1196 diff_1115520_712140# diff_1111370_704670# GND GND efet w=78020 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1197 GND diff_1111370_685580# diff_1115520_674790# GND efet w=78435 l=7885
+ ad=0 pd=0 as=8.21169e+08 ps=184260 
M1198 diff_1111370_685580# diff_1111370_685580# diff_1111370_685580# GND efet w=2490 l=4150
+ ad=2.34915e+08 pd=74700 as=0 ps=0 
M1199 diff_1111370_685580# diff_1111370_685580# diff_1111370_685580# GND efet w=2905 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1200 diff_1231720_712970# diff_273900_560250# diff_1111370_685580# GND efet w=14110 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1201 diff_1254960_682260# diff_258130_451520# diff_1231720_712970# GND efet w=14110 l=7470
+ ad=2.01848e+08 pd=59760 as=0 ps=0 
M1202 diff_1254960_682260# diff_1254960_682260# diff_1254960_682260# GND efet w=2075 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1203 diff_1254960_682260# diff_1254960_682260# diff_1254960_682260# GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1204 diff_1231720_712970# diff_1231720_738700# GND GND efet w=22410 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1205 Vdd Vdd diff_1231720_712970# GND efet w=8300 l=39840
+ ad=0 pd=0 as=0 ps=0 
M1206 diff_1477400_740360# Vdd Vdd GND efet w=6640 l=180940
+ ad=4.0094e+08 pd=107900 as=0 ps=0 
M1207 diff_1505620_931260# Vdd Vdd GND efet w=8300 l=24900
+ ad=0 pd=0 as=0 ps=0 
M1208 Vdd Vdd diff_1588620_812570# GND efet w=8300 l=24070
+ ad=0 pd=0 as=0 ps=0 
M1209 Vdd Vdd Vdd GND efet w=1660 l=5810
+ ad=0 pd=0 as=0 ps=0 
M1210 Vdd Vdd Vdd GND efet w=2075 l=4150
+ ad=0 pd=0 as=0 ps=0 
M1211 data_in GND GND GND efet w=112880 l=8300
+ ad=-6.44486e+08 pd=655700 as=0 ps=0 
M1212 cp GND GND GND efet w=112880 l=8300
+ ad=-1.27001e+09 pd=610880 as=0 ps=0 
M1213 diff_1231720_712970# diff_232400_451520# diff_1355390_712140# GND efet w=50215 l=7885
+ ad=0 pd=0 as=7.68124e+08 ps=185920 
M1214 diff_1115520_674790# diff_232400_451520# diff_991020_738700# GND efet w=49385 l=7055
+ ad=0 pd=0 as=0 ps=0 
M1215 GND diff_341130_652380# diff_991020_738700# GND efet w=22410 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1216 diff_991020_738700# Vdd Vdd GND efet w=8300 l=41500
+ ad=0 pd=0 as=0 ps=0 
M1217 GND diff_1254960_682260# diff_1231720_738700# GND efet w=38180 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1218 diff_1355390_712140# diff_1352070_704670# GND GND efet w=79680 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1219 diff_1566210_789330# diff_1477400_740360# GND GND efet w=164340 l=23240
+ ad=-1.01098e+09 pd=585980 as=0 ps=0 
M1220 GND cp diff_1477400_740360# GND efet w=14110 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1221 GND diff_1352070_685580# diff_1355390_674790# GND efet w=80925 l=7885
+ ad=0 pd=0 as=6.86833e+08 ps=152720 
M1222 diff_1355390_674790# diff_232400_451520# diff_1231720_738700# GND efet w=49800 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1223 GND diff_341130_652380# diff_1231720_738700# GND efet w=21580 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1224 diff_1466610_655700# Vdd Vdd GND efet w=8300 l=22410
+ ad=9.12104e+08 pd=179280 as=0 ps=0 
M1225 GND data_in diff_1466610_629970# GND efet w=163095 l=7885
+ ad=0 pd=0 as=1.71949e+09 ps=317060 
M1226 GND diff_1466610_629970# diff_1466610_655700# GND efet w=50630 l=8300
+ ad=0 pd=0 as=0 ps=0 
M1227 diff_1352070_704670# diff_1352070_704670# diff_1352070_704670# GND efet w=2075 l=4980
+ ad=2.18381e+08 pd=71380 as=0 ps=0 
M1228 diff_1352070_704670# diff_1352070_704670# diff_1352070_704670# GND efet w=3320 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1229 diff_1466610_655700# diff_273900_560250# diff_1352070_704670# GND efet w=14110 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1230 diff_1231720_738700# Vdd Vdd GND efet w=8300 l=41500
+ ad=0 pd=0 as=0 ps=0 
M1231 diff_1352070_685580# diff_1352070_685580# diff_1352070_685580# GND efet w=2075 l=4150
+ ad=2.18381e+08 pd=71380 as=0 ps=0 
M1232 diff_1352070_685580# diff_1352070_685580# diff_1352070_685580# GND efet w=3320 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1233 diff_1466610_629970# diff_273900_560250# diff_1352070_685580# GND efet w=14110 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1234 diff_1466610_629970# diff_1466610_629970# diff_1466610_629970# GND efet w=2075 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1235 diff_1466610_629970# diff_1466610_629970# diff_1466610_629970# GND efet w=2490 l=2490
+ ad=0 pd=0 as=0 ps=0 
M1236 diff_1466610_629970# Vdd Vdd GND efet w=10790 l=19920
+ ad=0 pd=0 as=0 ps=0 
M1237 Vdd Vdd Vdd GND efet w=2490 l=4980
+ ad=0 pd=0 as=0 ps=0 
M1238 Vdd Vdd diff_336150_519580# GND efet w=7885 l=42745
+ ad=0 pd=0 as=-2.06293e+09 ps=507960 
M1239 Vdd Vdd Vdd GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1240 Vdd Vdd Vdd GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1241 Vdd Vdd Vdd GND efet w=2075 l=7055
+ ad=0 pd=0 as=0 ps=0 
M1242 Vdd Vdd Vdd GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1243 Vdd Vdd Vdd GND efet w=2490 l=2490
+ ad=0 pd=0 as=0 ps=0 
M1244 Vdd Vdd Vdd GND efet w=3735 l=4150
+ ad=0 pd=0 as=0 ps=0 
M1245 Vdd Vdd Vdd GND efet w=2075 l=6225
+ ad=0 pd=0 as=0 ps=0 
M1246 Vdd Vdd Vdd GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1247 Vdd Vdd Vdd GND efet w=2490 l=2490
+ ad=0 pd=0 as=0 ps=0 
M1248 Vdd Vdd Vdd GND efet w=2075 l=4150
+ ad=0 pd=0 as=0 ps=0 
M1249 Vdd Vdd Vdd GND efet w=2075 l=6225
+ ad=0 pd=0 as=0 ps=0 
M1250 Vdd Vdd Vdd GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1251 Vdd Vdd Vdd GND efet w=2490 l=2490
+ ad=0 pd=0 as=0 ps=0 
M1252 Vdd Vdd Vdd GND efet w=2075 l=4980
+ ad=0 pd=0 as=0 ps=0 
M1253 Vdd Vdd Vdd GND efet w=2075 l=7055
+ ad=0 pd=0 as=0 ps=0 
M1254 Vdd Vdd Vdd GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1255 Vdd Vdd Vdd GND efet w=2490 l=2490
+ ad=0 pd=0 as=0 ps=0 
M1256 diff_278050_567720# diff_273900_560250# diff_278050_543650# GND efet w=14110 l=7470
+ ad=0 pd=0 as=2.33537e+08 ps=61420 
M1257 diff_273900_607560# diff_273900_560250# diff_289670_464800# GND efet w=14110 l=7470
+ ad=0 pd=0 as=2.08737e+08 ps=64740 
M1258 diff_289670_464800# diff_289670_464800# diff_289670_464800# GND efet w=2905 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1259 diff_289670_464800# diff_289670_464800# diff_289670_464800# GND efet w=2075 l=4150
+ ad=0 pd=0 as=0 ps=0 
M1260 diff_336150_519580# diff_232400_451520# diff_322040_502150# GND efet w=48970 l=7470
+ ad=0 pd=0 as=6.45499e+08 ps=147740 
M1261 diff_336150_519580# diff_341130_652380# GND GND efet w=21580 l=8300
+ ad=0 pd=0 as=0 ps=0 
M1262 diff_322040_502150# diff_278050_543650# GND GND efet w=77605 l=7885
+ ad=0 pd=0 as=0 ps=0 
M1263 GND diff_289670_464800# diff_305440_456500# GND efet w=78020 l=7470
+ ad=0 pd=0 as=7.66057e+08 ps=180940 
M1264 diff_336150_519580# diff_415830_432430# GND GND efet w=37350 l=8300
+ ad=0 pd=0 as=0 ps=0 
M1265 diff_336150_427450# diff_232400_451520# diff_305440_456500# GND efet w=49385 l=7885
+ ad=1.72707e+09 pd=338640 as=0 ps=0 
M1266 diff_336150_427450# Vdd Vdd GND efet w=8300 l=39840
+ ad=0 pd=0 as=0 ps=0 
M1267 Vdd Vdd diff_576020_519580# GND efet w=8300 l=42330
+ ad=0 pd=0 as=1.76358e+09 ps=375160 
M1268 diff_576020_519580# diff_232400_451520# diff_544480_499660# GND efet w=49800 l=7470
+ ad=0 pd=0 as=7.81213e+08 ps=184260 
M1269 diff_576020_519580# diff_341130_652380# GND GND efet w=22410 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1270 diff_544480_499660# diff_512940_454840# GND GND efet w=79680 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1271 GND diff_336150_519580# diff_336150_427450# GND efet w=21580 l=8300
+ ad=0 pd=0 as=0 ps=0 
M1272 diff_415830_432430# diff_415830_432430# diff_415830_432430# GND efet w=2075 l=7055
+ ad=2.13559e+08 pd=73040 as=0 ps=0 
M1273 diff_415830_432430# diff_415830_432430# diff_415830_432430# GND efet w=3735 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1274 diff_336150_427450# diff_258130_451520# diff_415830_432430# GND efet w=14110 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1275 diff_512940_454840# diff_273900_560250# diff_336150_427450# GND efet w=12450 l=7470
+ ad=1.9427e+08 pd=63080 as=0 ps=0 
M1276 diff_512940_454840# diff_512940_454840# diff_512940_454840# GND efet w=2905 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1277 diff_563570_456500# diff_512940_429940# GND GND efet w=76775 l=7885
+ ad=6.39988e+08 pd=146080 as=0 ps=0 
M1278 diff_576020_519580# diff_656530_432430# GND GND efet w=38595 l=7885
+ ad=0 pd=0 as=0 ps=0 
M1279 diff_576020_427450# diff_232400_451520# diff_563570_456500# GND efet w=49800 l=7470
+ ad=1.80078e+09 pd=345280 as=0 ps=0 
M1280 diff_512940_454840# diff_512940_454840# diff_512940_454840# GND efet w=830 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1281 diff_336150_519580# diff_336150_519580# diff_336150_519580# GND efet w=1660 l=6640
+ ad=0 pd=0 as=0 ps=0 
M1282 diff_336150_519580# diff_336150_519580# diff_336150_519580# GND efet w=3735 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1283 diff_512940_429940# diff_273900_560250# diff_336150_519580# GND efet w=12450 l=7470
+ ad=1.92203e+08 pd=63080 as=0 ps=0 
M1284 diff_512940_429940# diff_512940_429940# diff_512940_429940# GND efet w=1660 l=4150
+ ad=0 pd=0 as=0 ps=0 
M1285 diff_512940_429940# diff_512940_429940# diff_512940_429940# GND efet w=2490 l=2490
+ ad=0 pd=0 as=0 ps=0 
M1286 diff_336150_427450# diff_258130_451520# diff_444050_322040# GND efet w=14110 l=7470
+ ad=0 pd=0 as=9.65149e+08 ps=220780 
M1287 Vdd Vdd Vdd GND efet w=2075 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1288 Vdd Vdd Vdd GND efet w=2075 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1289 Vdd Vdd Vdd GND efet w=2075 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1290 Vdd Vdd Vdd GND efet w=2075 l=2075
+ ad=0 pd=0 as=0 ps=0 
M1291 Vdd Vdd diff_275560_234060# GND efet w=10375 l=19920
+ ad=0 pd=0 as=6.88211e+08 ps=161020 
M1292 Vdd diff_314570_311250# q5 GND efet w=24900 l=8300
+ ad=0 pd=0 as=9.94407e+08 ps=831660 
M1293 diff_275560_234060# diff_275560_234060# diff_275560_234060# GND efet w=2075 l=6225
+ ad=0 pd=0 as=0 ps=0 
M1294 diff_275560_234060# diff_275560_234060# diff_275560_234060# GND efet w=1660 l=5810
+ ad=0 pd=0 as=0 ps=0 
M1295 diff_275560_234060# diff_314570_311250# GND GND efet w=56025 l=7885
+ ad=0 pd=0 as=0 ps=0 
M1296 GND diff_275560_234060# q5 GND efet w=347355 l=7885
+ ad=0 pd=0 as=0 ps=0 
M1297 diff_576020_427450# Vdd Vdd GND efet w=8300 l=39840
+ ad=0 pd=0 as=0 ps=0 
M1298 Vdd Vdd diff_816720_520410# GND efet w=9130 l=42330
+ ad=0 pd=0 as=1.73052e+09 ps=373500 
M1299 diff_816720_520410# diff_232400_451520# diff_786010_499660# GND efet w=49800 l=7470
+ ad=0 pd=0 as=8.07391e+08 ps=184260 
M1300 diff_816720_520410# diff_341130_652380# GND GND efet w=22410 l=6640
+ ad=0 pd=0 as=0 ps=0 
M1301 diff_786010_499660# diff_754470_454010# GND GND efet w=78850 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1302 GND diff_576020_519580# diff_576020_427450# GND efet w=21580 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1303 diff_656530_432430# diff_656530_432430# diff_656530_432430# GND efet w=2075 l=6225
+ ad=2.18381e+08 pd=71380 as=0 ps=0 
M1304 diff_656530_432430# diff_656530_432430# diff_656530_432430# GND efet w=3320 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1305 diff_576020_427450# diff_258130_451520# diff_656530_432430# GND efet w=14110 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1306 diff_754470_454010# diff_273900_560250# diff_576020_427450# GND efet w=13280 l=7470
+ ad=1.99092e+08 pd=59760 as=0 ps=0 
M1307 diff_754470_454010# diff_754470_454010# diff_754470_454010# GND efet w=2075 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1308 diff_804270_456500# diff_754470_429110# GND GND efet w=77190 l=7470
+ ad=6.62722e+08 pd=147740 as=0 ps=0 
M1309 diff_816720_520410# diff_896400_434090# GND GND efet w=38180 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1310 diff_816720_427450# diff_232400_451520# diff_804270_456500# GND efet w=49800 l=7470
+ ad=1.80492e+09 pd=345280 as=0 ps=0 
M1311 diff_754470_454010# diff_754470_454010# diff_754470_454010# GND efet w=1245 l=1660
+ ad=0 pd=0 as=0 ps=0 
M1312 diff_576020_519580# diff_576020_519580# diff_576020_519580# GND efet w=1660 l=6640
+ ad=0 pd=0 as=0 ps=0 
M1313 diff_576020_519580# diff_576020_519580# diff_576020_519580# GND efet w=3735 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1314 diff_754470_429110# diff_273900_560250# diff_576020_519580# GND efet w=13280 l=7470
+ ad=1.99092e+08 pd=61420 as=0 ps=0 
M1315 diff_754470_429110# diff_754470_429110# diff_754470_429110# GND efet w=1660 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1316 diff_754470_429110# diff_754470_429110# diff_754470_429110# GND efet w=2075 l=2075
+ ad=0 pd=0 as=0 ps=0 
M1317 diff_576020_427450# diff_258130_451520# diff_684750_321210# GND efet w=14110 l=7470
+ ad=0 pd=0 as=9.65838e+08 ps=220780 
M1318 Vdd Vdd Vdd GND efet w=2075 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1319 Vdd Vdd Vdd GND efet w=2075 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1320 Vdd Vdd Vdd GND efet w=2075 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1321 Vdd Vdd Vdd GND efet w=2075 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1322 Vdd Vdd Vdd GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1323 Vdd Vdd Vdd GND efet w=2490 l=2490
+ ad=0 pd=0 as=0 ps=0 
M1324 Vdd Vdd diff_314570_311250# GND efet w=7885 l=24485
+ ad=0 pd=0 as=1.72087e+09 ps=336980 
M1325 Vdd Vdd diff_517090_234060# GND efet w=10790 l=19920
+ ad=0 pd=0 as=7.20589e+08 ps=166000 
M1326 Vdd diff_556100_312080# q6 GND efet w=24900 l=7470
+ ad=0 pd=0 as=1.05572e+09 ps=833320 
M1327 diff_444050_322040# diff_444050_322040# diff_444050_322040# GND efet w=2905 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1328 diff_444050_322040# diff_444050_322040# diff_444050_322040# GND efet w=2075 l=6225
+ ad=0 pd=0 as=0 ps=0 
M1329 diff_517090_234060# diff_517090_234060# diff_517090_234060# GND efet w=2490 l=6640
+ ad=0 pd=0 as=0 ps=0 
M1330 diff_517090_234060# diff_517090_234060# diff_517090_234060# GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1331 diff_517090_234060# diff_556100_312080# GND GND efet w=56440 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1332 diff_314570_311250# diff_314570_311250# diff_314570_311250# GND efet w=2490 l=7055
+ ad=0 pd=0 as=0 ps=0 
M1333 diff_314570_311250# diff_314570_311250# diff_314570_311250# GND efet w=3735 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1334 GND diff_207500_451520# diff_314570_311250# GND efet w=39010 l=8300
+ ad=0 pd=0 as=0 ps=0 
M1335 diff_314570_311250# diff_444050_322040# GND GND efet w=67230 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1336 GND diff_517090_234060# q6 GND efet w=347355 l=7885
+ ad=0 pd=0 as=0 ps=0 
M1337 diff_816720_427450# Vdd Vdd GND efet w=8300 l=39840
+ ad=0 pd=0 as=0 ps=0 
M1338 Vdd Vdd diff_1056590_520410# GND efet w=9130 l=42330
+ ad=0 pd=0 as=1.73534e+09 ps=373500 
M1339 diff_1056590_520410# diff_232400_451520# diff_1025050_499660# GND efet w=49800 l=7470
+ ad=0 pd=0 as=8.19791e+08 ps=185920 
M1340 diff_1056590_520410# diff_341130_652380# GND GND efet w=22410 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1341 diff_1025050_499660# diff_993510_454010# GND GND efet w=79680 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1342 GND diff_816720_520410# diff_816720_427450# GND efet w=21580 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1343 diff_896400_434090# diff_896400_434090# diff_896400_434090# GND efet w=2075 l=7055
+ ad=2.17004e+08 pd=73040 as=0 ps=0 
M1344 diff_896400_434090# diff_896400_434090# diff_896400_434090# GND efet w=3320 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1345 diff_816720_427450# diff_258130_451520# diff_896400_434090# GND efet w=14110 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1346 diff_993510_454010# diff_273900_560250# diff_816720_427450# GND efet w=13280 l=6640
+ ad=2.05981e+08 pd=63080 as=0 ps=0 
M1347 diff_993510_454010# diff_993510_454010# diff_993510_454010# GND efet w=2490 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1348 diff_1043310_456500# diff_993510_429110# GND GND efet w=77605 l=7055
+ ad=6.765e+08 pd=149400 as=0 ps=0 
M1349 diff_1056590_520410# diff_1137100_433260# GND GND efet w=38180 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1350 diff_1056590_427450# diff_232400_451520# diff_1043310_456500# GND efet w=49800 l=7470
+ ad=1.82421e+09 pd=346940 as=0 ps=0 
M1351 diff_993510_454010# diff_993510_454010# diff_993510_454010# GND efet w=1245 l=2075
+ ad=0 pd=0 as=0 ps=0 
M1352 diff_816720_520410# diff_816720_520410# diff_816720_520410# GND efet w=1660 l=6640
+ ad=0 pd=0 as=0 ps=0 
M1353 diff_816720_520410# diff_816720_520410# diff_816720_520410# GND efet w=3735 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1354 diff_993510_429110# diff_273900_560250# diff_816720_520410# GND efet w=13280 l=6640
+ ad=2.10114e+08 pd=63080 as=0 ps=0 
M1355 diff_993510_429110# diff_993510_429110# diff_993510_429110# GND efet w=1660 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1356 diff_993510_429110# diff_993510_429110# diff_993510_429110# GND efet w=2075 l=2075
+ ad=0 pd=0 as=0 ps=0 
M1357 diff_816720_427450# diff_258130_451520# diff_924620_321210# GND efet w=14110 l=7470
+ ad=0 pd=0 as=9.65838e+08 ps=220780 
M1358 Vdd Vdd Vdd GND efet w=2075 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1359 Vdd Vdd Vdd GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1360 Vdd Vdd Vdd GND efet w=2075 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1361 Vdd Vdd Vdd GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1362 Vdd Vdd Vdd GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1363 Vdd Vdd Vdd GND efet w=2490 l=2490
+ ad=0 pd=0 as=0 ps=0 
M1364 Vdd Vdd diff_556100_312080# GND efet w=7885 l=25315
+ ad=0 pd=0 as=1.76083e+09 ps=346940 
M1365 Vdd Vdd diff_756130_234890# GND efet w=10790 l=20750
+ ad=0 pd=0 as=6.98545e+08 ps=162680 
M1366 Vdd diff_795140_312080# q7 GND efet w=24900 l=7470
+ ad=0 pd=0 as=1.05641e+09 ps=833320 
M1367 diff_684750_321210# diff_684750_321210# diff_684750_321210# GND efet w=2905 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1368 diff_684750_321210# diff_684750_321210# diff_684750_321210# GND efet w=2075 l=6225
+ ad=0 pd=0 as=0 ps=0 
M1369 diff_756130_234890# diff_756130_234890# diff_756130_234890# GND efet w=2075 l=6225
+ ad=0 pd=0 as=0 ps=0 
M1370 diff_756130_234890# diff_756130_234890# diff_756130_234890# GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1371 diff_756130_234890# diff_795140_312080# GND GND efet w=56025 l=7885
+ ad=0 pd=0 as=0 ps=0 
M1372 diff_556100_312080# diff_556100_312080# diff_556100_312080# GND efet w=4565 l=5395
+ ad=0 pd=0 as=0 ps=0 
M1373 diff_556100_312080# diff_556100_312080# diff_556100_312080# GND efet w=3735 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1374 GND diff_207500_451520# diff_556100_312080# GND efet w=39010 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1375 diff_556100_312080# diff_684750_321210# GND GND efet w=66815 l=7885
+ ad=0 pd=0 as=0 ps=0 
M1376 GND diff_756130_234890# q7 GND efet w=347355 l=7885
+ ad=0 pd=0 as=0 ps=0 
M1377 diff_1056590_427450# Vdd Vdd GND efet w=8300 l=39840
+ ad=0 pd=0 as=0 ps=0 
M1378 Vdd Vdd diff_1297290_520410# GND efet w=8300 l=42330
+ ad=0 pd=0 as=1.28962e+09 ps=255640 
M1379 diff_341130_652380# Vdd Vdd GND efet w=8300 l=16600
+ ad=7.32301e+08 pd=151060 as=0 ps=0 
M1380 GND diff_1483210_498830# diff_341130_652380# GND efet w=61835 l=7885
+ ad=0 pd=0 as=0 ps=0 
M1381 Vdd Vdd diff_1509770_516260# GND efet w=8300 l=62250
+ ad=0 pd=0 as=1.06986e+09 ps=189240 
M1382 Vdd Vdd diff_1483210_498830# GND efet w=8715 l=23655
+ ad=0 pd=0 as=4.84297e+08 ps=114540 
M1383 diff_1297290_520410# diff_232400_451520# diff_1266580_499660# GND efet w=48970 l=7470
+ ad=0 pd=0 as=7.97746e+08 ps=182600 
M1384 diff_1297290_520410# diff_341130_652380# GND GND efet w=22410 l=8300
+ ad=0 pd=0 as=0 ps=0 
M1385 diff_1266580_499660# diff_1235040_454010# GND GND efet w=78020 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1386 GND diff_1056590_520410# diff_1056590_427450# GND efet w=22410 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1387 diff_1137100_433260# diff_1137100_433260# diff_1137100_433260# GND efet w=2075 l=7885
+ ad=2.27337e+08 pd=76360 as=0 ps=0 
M1388 diff_1137100_433260# diff_1137100_433260# diff_1137100_433260# GND efet w=3320 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1389 diff_1056590_427450# diff_258130_451520# diff_1137100_433260# GND efet w=14110 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1390 diff_1235040_454010# diff_273900_560250# diff_1056590_427450# GND efet w=13280 l=7470
+ ad=2.05292e+08 pd=63080 as=0 ps=0 
M1391 diff_1235040_454010# diff_1235040_454010# diff_1235040_454010# GND efet w=2075 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1392 diff_1284840_456500# diff_1235040_429110# GND GND efet w=76360 l=7470
+ ad=6.55833e+08 pd=146080 as=0 ps=0 
M1393 diff_1297290_520410# diff_1376970_433260# GND GND efet w=39840 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1394 diff_1297290_428280# diff_232400_451520# diff_1284840_456500# GND efet w=48970 l=7470
+ ad=1.55623e+09 pd=278880 as=0 ps=0 
M1395 diff_1235040_454010# diff_1235040_454010# diff_1235040_454010# GND efet w=1660 l=2075
+ ad=0 pd=0 as=0 ps=0 
M1396 diff_1056590_520410# diff_1056590_520410# diff_1056590_520410# GND efet w=1660 l=6640
+ ad=0 pd=0 as=0 ps=0 
M1397 diff_1056590_520410# diff_1056590_520410# diff_1056590_520410# GND efet w=3320 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1398 diff_1235040_429110# diff_273900_560250# diff_1056590_520410# GND efet w=13280 l=7470
+ ad=2.08048e+08 pd=64740 as=0 ps=0 
M1399 diff_1235040_429110# diff_1235040_429110# diff_1235040_429110# GND efet w=1660 l=4150
+ ad=0 pd=0 as=0 ps=0 
M1400 diff_1235040_429110# diff_1235040_429110# diff_1235040_429110# GND efet w=2075 l=2075
+ ad=0 pd=0 as=0 ps=0 
M1401 diff_1056590_427450# diff_258130_451520# diff_1165320_321210# GND efet w=14110 l=7470
+ ad=0 pd=0 as=9.66527e+08 ps=220780 
M1402 Vdd Vdd Vdd GND efet w=2075 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1403 Vdd Vdd Vdd GND efet w=2075 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1404 Vdd Vdd Vdd GND efet w=2075 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1405 Vdd Vdd Vdd GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1406 Vdd Vdd Vdd GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1407 Vdd Vdd Vdd GND efet w=2490 l=2490
+ ad=0 pd=0 as=0 ps=0 
M1408 Vdd Vdd diff_795140_312080# GND efet w=8300 l=24900
+ ad=0 pd=0 as=1.7567e+09 ps=338640 
M1409 Vdd Vdd diff_994340_234060# GND efet w=9960 l=20750
+ ad=0 pd=0 as=6.96478e+08 ps=162680 
M1410 Vdd diff_1033350_312080# q8 GND efet w=24900 l=7470
+ ad=0 pd=0 as=1.11083e+09 ps=836640 
M1411 diff_924620_321210# diff_924620_321210# diff_924620_321210# GND efet w=2905 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1412 diff_924620_321210# diff_924620_321210# diff_924620_321210# GND efet w=2075 l=4150
+ ad=0 pd=0 as=0 ps=0 
M1413 diff_994340_234060# diff_994340_234060# diff_994340_234060# GND efet w=2075 l=6225
+ ad=0 pd=0 as=0 ps=0 
M1414 diff_994340_234060# diff_994340_234060# diff_994340_234060# GND efet w=2075 l=6225
+ ad=0 pd=0 as=0 ps=0 
M1415 diff_994340_234060# diff_1033350_312080# GND GND efet w=55610 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1416 diff_795140_312080# diff_795140_312080# diff_795140_312080# GND efet w=2490 l=7885
+ ad=0 pd=0 as=0 ps=0 
M1417 diff_795140_312080# diff_795140_312080# diff_795140_312080# GND efet w=3735 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1418 GND diff_207500_451520# diff_795140_312080# GND efet w=38595 l=7885
+ ad=0 pd=0 as=0 ps=0 
M1419 diff_795140_312080# diff_924620_321210# GND GND efet w=67230 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1420 GND diff_994340_234060# q8 GND efet w=347770 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1421 diff_1297290_428280# Vdd Vdd GND efet w=8300 l=40670
+ ad=0 pd=0 as=0 ps=0 
M1422 GND diff_1297290_520410# diff_1297290_428280# GND efet w=22410 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1423 diff_1483210_498830# diff_1509770_516260# GND GND efet w=38180 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1424 Vdd Vdd diff_1566210_789330# GND efet w=7885 l=180525
+ ad=0 pd=0 as=0 ps=0 
M1425 GND diff_1505620_931260# diff_1509770_516260# GND efet w=20335 l=7885
+ ad=0 pd=0 as=0 ps=0 
M1426 diff_1509770_516260# diff_1483210_498830# diff_1552100_502150# GND efet w=28220 l=7470
+ ad=0 pd=0 as=3.04494e+08 ps=78020 
M1427 diff_1552100_502150# diff_1548780_494680# GND GND efet w=28220 l=8300
+ ad=0 pd=0 as=0 ps=0 
M1428 GND diff_1505620_352750# diff_1472420_424130# GND efet w=27805 l=7885
+ ad=0 pd=0 as=1.33715e+09 ps=267260 
M1429 GND diff_273900_560250# diff_1472420_449860# GND efet w=68890 l=7470
+ ad=0 pd=0 as=1.73878e+09 ps=287180 
M1430 GND diff_1472420_424130# diff_1505620_352750# GND efet w=34030 l=7470
+ ad=0 pd=0 as=-1.97337e+09 ps=448200 
M1431 diff_1472420_424130# diff_1472420_424130# diff_1472420_424130# GND efet w=2075 l=7055
+ ad=0 pd=0 as=0 ps=0 
M1432 diff_1376970_433260# diff_1376970_433260# diff_1376970_433260# GND efet w=2075 l=7055
+ ad=2.21137e+08 pd=73040 as=0 ps=0 
M1433 diff_1376970_433260# diff_1376970_433260# diff_1376970_433260# GND efet w=2905 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1434 diff_1297290_428280# diff_258130_451520# diff_1376970_433260# GND efet w=14110 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1435 diff_1472420_449860# diff_1297290_520410# diff_1472420_424130# GND efet w=43990 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1436 diff_1472420_449860# diff_1297290_428280# diff_1505620_352750# GND efet w=76360 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1437 diff_1472420_424130# diff_1472420_424130# diff_1472420_424130# GND efet w=3320 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1438 diff_1297290_428280# diff_258130_451520# diff_1405190_321210# GND efet w=14110 l=7470
+ ad=0 pd=0 as=9.77549e+08 ps=222440 
M1439 Vdd Vdd diff_1505620_352750# GND efet w=8715 l=21995
+ ad=0 pd=0 as=0 ps=0 
M1440 diff_1472420_424130# Vdd Vdd GND efet w=8715 l=40255
+ ad=0 pd=0 as=0 ps=0 
M1441 Vdd Vdd Vdd GND efet w=2075 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1442 Vdd Vdd Vdd GND efet w=2075 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1443 Vdd Vdd Vdd GND efet w=2075 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1444 Vdd Vdd Vdd GND efet w=1660 l=4980
+ ad=0 pd=0 as=0 ps=0 
M1445 Vdd Vdd Vdd GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1446 Vdd Vdd Vdd GND efet w=2490 l=2490
+ ad=0 pd=0 as=0 ps=0 
M1447 Vdd Vdd diff_1033350_312080# GND efet w=8300 l=24900
+ ad=0 pd=0 as=1.78701e+09 ps=340300 
M1448 Vdd Vdd diff_1236700_234890# GND efet w=10790 l=20750
+ ad=0 pd=0 as=7.02678e+08 ps=162680 
M1449 Vdd diff_1276540_312080# q9 GND efet w=24900 l=7470
+ ad=0 pd=0 as=1.12599e+09 ps=838300 
M1450 diff_1165320_321210# diff_1165320_321210# diff_1165320_321210# GND efet w=2905 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1451 diff_1165320_321210# diff_1165320_321210# diff_1165320_321210# GND efet w=2075 l=6225
+ ad=0 pd=0 as=0 ps=0 
M1452 diff_1236700_234890# diff_1236700_234890# diff_1236700_234890# GND efet w=1660 l=5810
+ ad=0 pd=0 as=0 ps=0 
M1453 diff_1236700_234890# diff_1236700_234890# diff_1236700_234890# GND efet w=2075 l=4150
+ ad=0 pd=0 as=0 ps=0 
M1454 diff_1236700_234890# diff_1276540_312080# GND GND efet w=55610 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1455 diff_1033350_312080# diff_1033350_312080# diff_1033350_312080# GND efet w=2075 l=7055
+ ad=0 pd=0 as=0 ps=0 
M1456 diff_1033350_312080# diff_1033350_312080# diff_1033350_312080# GND efet w=3735 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1457 GND diff_207500_451520# diff_1033350_312080# GND efet w=39010 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1458 diff_1033350_312080# diff_1165320_321210# GND GND efet w=66400 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1459 GND diff_1236700_234890# q9 GND efet w=349015 l=7885
+ ad=0 pd=0 as=0 ps=0 
M1460 Vdd Vdd Vdd GND efet w=2490 l=4150
+ ad=0 pd=0 as=0 ps=0 
M1461 Vdd Vdd Vdd GND efet w=2075 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1462 Vdd Vdd Vdd GND efet w=1660 l=3320
+ ad=0 pd=0 as=0 ps=0 
M1463 Vdd Vdd Vdd GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1464 diff_1548780_494680# Vdd Vdd GND efet w=6640 l=120350
+ ad=2.30782e+08 pd=64740 as=0 ps=0 
M1465 Vdd Vdd Vdd GND efet w=2075 l=7055
+ ad=0 pd=0 as=0 ps=0 
M1466 Vdd Vdd Vdd GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1467 Vdd Vdd Vdd GND efet w=2490 l=2490
+ ad=0 pd=0 as=0 ps=0 
M1468 Vdd Vdd Vdd GND efet w=3735 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1469 Vdd Vdd diff_1276540_312080# GND efet w=8300 l=24900
+ ad=0 pd=0 as=1.76772e+09 ps=338640 
M1470 Vdd Vdd diff_207500_451520# GND efet w=9960 l=18260
+ ad=0 pd=0 as=-1.98233e+09 ps=408360 
M1471 diff_1505620_352750# diff_1505620_352750# diff_1505620_352750# GND efet w=2490 l=2490
+ ad=0 pd=0 as=0 ps=0 
M1472 diff_1505620_352750# diff_1505620_352750# diff_1505620_352750# GND efet w=2075 l=6225
+ ad=0 pd=0 as=0 ps=0 
M1473 Vdd diff_1505620_352750# serial_out GND efet w=49800 l=7470
+ ad=0 pd=0 as=6.86469e+08 ps=654040 
M1474 diff_1405190_321210# diff_1405190_321210# diff_1405190_321210# GND efet w=2905 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1475 diff_1405190_321210# diff_1405190_321210# diff_1405190_321210# GND efet w=2075 l=6225
+ ad=0 pd=0 as=0 ps=0 
M1476 diff_207500_451520# e GND GND efet w=166830 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1477 diff_1276540_312080# diff_1276540_312080# diff_1276540_312080# GND efet w=2075 l=7055
+ ad=0 pd=0 as=0 ps=0 
M1478 diff_1276540_312080# diff_1276540_312080# diff_1276540_312080# GND efet w=2905 l=2905
+ ad=0 pd=0 as=0 ps=0 
M1479 GND diff_207500_451520# diff_1276540_312080# GND efet w=39425 l=7885
+ ad=0 pd=0 as=0 ps=0 
M1480 diff_1276540_312080# diff_1405190_321210# GND GND efet w=67230 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1481 Vdd Vdd Vdd GND efet w=1660 l=1660
+ ad=0 pd=0 as=0 ps=0 
M1482 Vdd Vdd Vdd GND efet w=2075 l=4565
+ ad=0 pd=0 as=0 ps=0 
M1483 diff_1534670_282200# Vdd Vdd GND efet w=8300 l=16600
+ ad=1.07951e+09 pd=185920 as=0 ps=0 
M1484 diff_1534670_282200# diff_1534670_282200# diff_1534670_282200# GND efet w=2075 l=3735
+ ad=0 pd=0 as=0 ps=0 
M1485 serial_out diff_1534670_282200# GND GND efet w=228665 l=7885
+ ad=0 pd=0 as=0 ps=0 
M1486 diff_1534670_282200# diff_1534670_282200# diff_1534670_282200# GND efet w=1660 l=1660
+ ad=0 pd=0 as=0 ps=0 
M1487 diff_1534670_282200# diff_1505620_352750# GND GND efet w=53120 l=7470
+ ad=0 pd=0 as=0 ps=0 
M1488 e GND GND GND efet w=111220 l=9130
+ ad=-1.50079e+09 pd=529540 as=0 ps=0 
C0 metal_567720_25730# gnd! 13.7fF ;**FLOATING
C1 metal_530370_44820# gnd! 7.5fF ;**FLOATING
C2 metal_530370_63910# gnd! 65.6fF ;**FLOATING
C3 metal_505470_64740# gnd! 27.5fF ;**FLOATING
C4 metal_605900_125330# gnd! 175.9fF ;**FLOATING
C5 metal_505470_151060# gnd! 4.6fF ;**FLOATING
C6 metal_649060_1066550# gnd! 54.9fF ;**FLOATING
C7 metal_597600_1064890# gnd! 55.7fF ;**FLOATING
C8 metal_546140_1082320# gnd! 46.9fF ;**FLOATING
C9 metal_700520_1115520# gnd! 46.5fF ;**FLOATING
C10 metal_281370_1115520# gnd! 8.7fF ;**FLOATING
C11 metal_302120_1144570# gnd! 8.9fF ;**FLOATING
C12 diff_1538820_21580# gnd! 1030.2fF ;**FLOATING
C13 diff_1534670_282200# gnd! 257.3fF
C14 serial_out gnd! 666.4fF
C15 e gnd! 803.6fF
C16 q9 gnd! 895.1fF
C17 diff_1236700_234890# gnd! 254.5fF
C18 diff_1276540_312080# gnd! 313.8fF
C19 diff_1405190_321210# gnd! 161.1fF
C20 diff_1472420_449860# gnd! 202.6fF
C21 diff_1472420_424130# gnd! 243.6fF
C22 diff_1505620_352750# gnd! 444.6fF
C23 diff_1552100_502150# gnd! 38.3fF
C24 diff_1548780_494680# gnd! 94.2fF
C25 q8 gnd! 841.2fF
C26 diff_994340_234060# gnd! 251.4fF
C27 diff_1033350_312080# gnd! 321.7fF
C28 diff_1165320_321210# gnd! 159.2fF
C29 diff_1297290_428280# gnd! 310.0fF
C30 diff_1376970_433260# gnd! 81.9fF
C31 diff_1284840_456500# gnd! 80.2fF
C32 diff_1235040_429110# gnd! 87.2fF
C33 diff_1235040_454010# gnd! 88.0fF
C34 diff_1266580_499660# gnd! 98.0fF
C35 diff_1509770_516260# gnd! 180.8fF
C36 diff_1297290_520410# gnd! 277.8fF
C37 diff_1483210_498830# gnd! 154.8fF
C38 q7 gnd! 773.2fF
C39 diff_756130_234890# gnd! 254.7fF
C40 diff_795140_312080# gnd! 312.7fF
C41 diff_924620_321210# gnd! 158.9fF
C42 diff_1056590_427450# gnd! 275.1fF
C43 diff_1137100_433260# gnd! 81.7fF
C44 diff_1043310_456500# gnd! 82.6fF
C45 diff_993510_429110# gnd! 85.1fF
C46 diff_993510_454010# gnd! 89.8fF
C47 diff_1025050_499660# gnd! 100.6fF
C48 diff_1056590_520410# gnd! 327.6fF
C49 q6 gnd! 955.5fF
C50 diff_517090_234060# gnd! 259.4fF
C51 diff_556100_312080# gnd! 312.6fF
C52 diff_684750_321210# gnd! 161.4fF
C53 diff_816720_427450# gnd! 271.8fF
C54 diff_896400_434090# gnd! 82.6fF
C55 diff_804270_456500# gnd! 81.0fF
C56 diff_754470_429110# gnd! 84.8fF
C57 diff_754470_454010# gnd! 87.0fF
C58 diff_786010_499660# gnd! 99.2fF
C59 diff_816720_520410# gnd! 325.8fF
C60 q5 gnd! 968.7fF
C61 diff_275560_234060# gnd! 259.8fF
C62 diff_314570_311250# gnd! 311.6fF
C63 diff_444050_322040# gnd! 160.1fF
C64 diff_576020_427450# gnd! 271.0fF
C65 diff_656530_432430# gnd! 81.5fF
C66 diff_563570_456500# gnd! 78.6fF
C67 diff_512940_429940# gnd! 85.7fF
C68 diff_512940_454840# gnd! 87.0fF
C69 diff_544480_499660# gnd! 96.5fF
C70 diff_576020_519580# gnd! 328.1fF
C71 diff_336150_427450# gnd! 263.6fF
C72 diff_415830_432430# gnd! 83.7fF
C73 diff_305440_456500# gnd! 94.7fF
C74 diff_322040_502150# gnd! 79.3fF
C75 diff_289670_464800# gnd! 109.5fF
C76 diff_278050_543650# gnd! 98.1fF
C77 diff_336150_519580# gnd! 392.3fF
C78 diff_1466610_629970# gnd! 279.9fF
C79 diff_1466610_655700# gnd! 109.1fF
C80 diff_1355390_674790# gnd! 84.0fF
C81 diff_1352070_685580# gnd! 92.7fF
C82 diff_1352070_704670# gnd! 89.5fF
C83 diff_1355390_712140# gnd! 95.4fF
C84 diff_1477400_740360# gnd! 299.0fF
C85 cp gnd! 674.9fF
C86 diff_1115520_674790# gnd! 100.5fF
C87 diff_1254960_682260# gnd! 77.9fF
C88 diff_1231720_712970# gnd! 266.0fF
C89 diff_1111370_685580# gnd! 93.6fF
C90 diff_1231720_738700# gnd! 349.8fF
C91 diff_1115520_712140# gnd! 81.1fF
C92 diff_1111370_704670# gnd! 90.0fF
C93 diff_1566210_789330# gnd! 657.4fF
C94 diff_1588620_812570# gnd! 188.7fF
C95 diff_1505620_931260# gnd! 322.3fF
C96 diff_875650_674790# gnd! 101.9fF
C97 diff_1013430_682260# gnd! 78.8fF
C98 diff_991020_712970# gnd! 270.5fF
C99 diff_871500_685580# gnd! 90.9fF
C100 diff_991020_738700# gnd! 340.3fF
C101 diff_875650_712140# gnd! 79.4fF
C102 diff_871500_704670# gnd! 89.0fF
C103 diff_1257450_846600# gnd! 318.6fF
C104 diff_1273220_771900# gnd! 158.8fF
C105 diff_1365350_939560# gnd! 254.2fF
C106 diff_634950_673960# gnd! 102.1fF
C107 diff_773560_682260# gnd! 79.7fF
C108 diff_751150_712970# gnd! 270.6fF
C109 diff_341130_652380# gnd! 901.3fF
C110 diff_630800_686410# gnd! 91.9fF
C111 diff_751150_738700# gnd! 340.0fF
C112 diff_634950_712140# gnd! 80.2fF
C113 diff_630800_705500# gnd! 90.0fF
C114 diff_1016750_846600# gnd! 317.4fF
C115 diff_1032520_771900# gnd! 164.9fF
C116 diff_1125480_939560# gnd! 253.0fF
C117 diff_395080_673960# gnd! 101.1fF
C118 diff_532860_681430# gnd! 82.4fF
C119 diff_510450_712970# gnd! 270.1fF
C120 diff_390930_685580# gnd! 93.9fF
C121 diff_510450_738700# gnd! 339.2fF
C122 diff_395080_711310# gnd! 81.9fF
C123 diff_390930_703840# gnd! 91.0fF
C124 diff_776880_846600# gnd! 318.9fF
C125 diff_792650_771900# gnd! 157.8fF
C126 diff_884780_939560# gnd! 252.2fF
C127 diff_273900_607560# gnd! 407.5fF
C128 diff_292990_681430# gnd! 79.5fF
C129 diff_278050_567720# gnd! 315.5fF
C130 diff_536180_846600# gnd! 319.4fF
C131 diff_551950_771900# gnd! 165.3fF
C132 diff_644910_939560# gnd! 252.3fF
C133 diff_207500_451520# gnd! 866.3fF
C134 diff_296310_846600# gnd! 314.5fF
C135 diff_312080_771900# gnd! 158.3fF
C136 diff_404210_938730# gnd! 257.7fF
C137 q0 gnd! 697.2fF
C138 q1 gnd! 705.2fF
C139 q2 gnd! 800.0fF
C140 q3 gnd! 974.7fF
C141 q4 gnd! 982.8fF
C142 diff_1621820_879800# gnd! 155.6fF
C143 data_in gnd! 829.0fF
C144 diff_273900_560250# gnd! 1764.9fF
C145 diff_232400_451520# gnd! 2418.5fF
C146 diff_1466610_1008450# gnd! 509.3fF
C147 diff_1540480_996000# gnd! 287.7fF
C148 diff_258130_451520# gnd! 1817.0fF
C149 Vdd gnd! 7800.5fF
C150 diff_291330_1124650# gnd! 13.9fF ;**FLOATING
C151 diff_283030_1135440# gnd! 20.0fF ;**FLOATING
C152 diff_282200_1144570# gnd! 74.3fF ;**FLOATING
C153 diff_283030_1154530# gnd! 39.8fF ;**FLOATING
