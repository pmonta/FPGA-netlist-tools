* SPICE3 file created from 4004.ext - technology: nmos

.option scale=0.001u

M1000 GND diff_622050_2844900# diff_627850_2752100# GND efet w=89900 l=11600
+ ad=-1.11604e+09 pd=2.81947e+08 as=-1.02724e+09 ps=2.0793e+06 
M1001 GND GND test GND efet w=119625 l=15225
+ ad=0 pd=0 as=-4.04902e+08 ps=1.827e+06 
M1002 reset GND GND GND efet w=118175 l=15225
+ ad=-2.6824e+08 pd=1.9343e+06 as=0 ps=0 
M1003 GND diff_443700_3526400# diff_507500_3552500# GND efet w=26100 l=13050
+ ad=0 pd=0 as=-6.7236e+08 ps=884500 
M1004 GND diff_916400_3567000# diff_909150_3567000# GND efet w=30450 l=12325
+ ad=0 pd=0 as=1.5979e+08 ps=66700 
M1005 diff_909150_3567000# diff_887400_2863750# diff_622050_2844900# GND efet w=26100 l=13050
+ ad=0 pd=0 as=-1.39806e+09 ps=5.2983e+06 
M1006 GND diff_345100_3549600# diff_443700_3526400# GND efet w=21750 l=11600
+ ad=0 pd=0 as=6.66492e+08 ps=139200 
M1007 diff_507500_3552500# diff_345100_3549600# diff_493000_3507550# GND efet w=78300 l=11600
+ ad=0 pd=0 as=1.0113e+09 ps=266800 
M1008 diff_443700_3526400# GND GND GND efet w=7250 l=69600
+ ad=0 pd=0 as=0 ps=0 
M1009 diff_443700_3526400# GND GND GND efet w=23925 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1010 GND GND diff_507500_3552500# GND efet w=8700 l=30450
+ ad=0 pd=0 as=0 ps=0 
M1011 diff_493000_3507550# GND GND GND efet w=126150 l=30450
+ ad=0 pd=0 as=0 ps=0 
M1012 GND diff_629300_2881150# diff_606100_2879700# GND efet w=44225 l=13775
+ ad=0 pd=0 as=-1.96241e+09 ps=2.8043e+06 
M1013 diff_627850_2752100# diff_627850_2752100# GND GND efet w=44225 l=17400
+ ad=0 pd=0 as=0 ps=0 
M1014 diff_622050_2844900# diff_784450_2863750# diff_507500_3552500# GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1015 GND GND diff_333500_3384300# GND efet w=15225 l=12325
+ ad=0 pd=0 as=8.9146e+08 ps=255200 
M1016 GND GND diff_345100_3549600# GND efet w=5075 l=18125
+ ad=0 pd=0 as=4.4573e+08 ps=153700 
M1017 GND diff_320450_2669450# GND GND efet w=21025 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1018 diff_606100_2879700# diff_606100_2879700# GND GND efet w=34075 l=21750
+ ad=0 pd=0 as=0 ps=0 
M1019 diff_329150_3371250# diff_320450_2669450# GND GND efet w=20300 l=11600
+ ad=3.23785e+08 pd=87000 as=0 ps=0 
M1020 diff_333500_3384300# diff_329150_3371250# diff_298700_3108800# GND efet w=14500 l=12325
+ ad=0 pd=0 as=1.005e+09 ps=246500 
M1021 diff_345100_3549600# diff_329150_3371250# diff_323350_3108800# GND efet w=26100 l=11600
+ ad=0 pd=0 as=6.53878e+08 ps=165300 
M1022 GND diff_329150_3371250# diff_493000_3316150# GND efet w=123250 l=11600
+ ad=0 pd=0 as=9.71355e+08 ps=243600 
M1023 GND diff_50750_3136350# GND GND efet w=1224525 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1024 diff_50750_3136350# diff_50750_3136350# diff_50750_3136350# GND efet w=63075 l=20300
+ ad=1.66938e+09 pd=539400 as=0 ps=0 
M1025 GND GND diff_50750_3136350# GND efet w=5800 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1026 GND diff_50750_3136350# diff_50750_3136350# GND efet w=10150 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1027 GND GND GND GND efet w=66700 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1028 GND GND GND GND efet w=11600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1029 GND GND GND GND efet w=6525 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1030 GND GND GND GND efet w=620600 l=71775
+ ad=0 pd=0 as=0 ps=0 
M1031 diff_606100_2879700# diff_606100_2879700# GND GND efet w=31175 l=22475
+ ad=0 pd=0 as=0 ps=0 
M1032 GND GND diff_361050_3108800# GND efet w=7975 l=19575
+ ad=0 pd=0 as=4.39422e+08 ps=133400 
M1033 diff_507500_3274100# diff_361050_3108800# diff_493000_3316150# GND efet w=68150 l=11600
+ ad=-7.92202e+08 pd=896100 as=0 ps=0 
M1034 GND diff_329150_3371250# GND GND efet w=23200 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1035 GND GND GND GND efet w=7250 l=68150
+ ad=0 pd=0 as=0 ps=0 
M1036 GND GND diff_507500_3274100# GND efet w=7250 l=27550
+ ad=0 pd=0 as=0 ps=0 
M1037 GND diff_361050_3108800# GND GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1038 diff_507500_3274100# GND GND GND efet w=23200 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1039 GND diff_442250_3204500# diff_507500_3229150# GND efet w=26100 l=11600
+ ad=0 pd=0 as=-8.84712e+08 ps=881600 
M1040 GND diff_378450_3143600# diff_442250_3204500# GND efet w=23925 l=11600
+ ad=0 pd=0 as=7.50593e+08 ps=145000 
M1041 diff_507500_3229150# diff_378450_3143600# diff_491550_3187100# GND efet w=70325 l=12325
+ ad=0 pd=0 as=9.27202e+08 ps=249400 
M1042 diff_442250_3204500# GND GND GND efet w=7975 l=67425
+ ad=0 pd=0 as=0 ps=0 
M1043 diff_442250_3204500# GND GND GND efet w=21025 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1044 GND GND diff_507500_3229150# GND efet w=7975 l=29725
+ ad=0 pd=0 as=0 ps=0 
M1045 diff_491550_3187100# GND GND GND efet w=116000 l=21750
+ ad=0 pd=0 as=0 ps=0 
M1046 diff_361050_3108800# GND diff_359600_3089950# GND efet w=23200 l=18850
+ ad=0 pd=0 as=1.2615e+08 ps=49300 
M1047 diff_298700_3108800# GND diff_298700_3089950# GND efet w=13050 l=11600
+ ad=0 pd=0 as=9.46125e+07 ps=40600 
M1048 diff_323350_3108800# GND diff_323350_3089950# GND efet w=23200 l=11600
+ ad=0 pd=0 as=1.682e+08 ps=60900 
M1049 GND GND diff_378450_3143600# GND efet w=9425 l=13775
+ ad=0 pd=0 as=8.38897e+08 ps=229100 
M1050 GND diff_320450_2669450# GND GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1051 diff_507500_3552500# diff_727900_2842000# diff_622050_2844900# GND efet w=14500 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1052 diff_622050_2844900# diff_622050_2844900# diff_507500_3552500# GND efet w=9425 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1053 diff_622050_2844900# diff_622050_2844900# diff_507500_3274100# GND efet w=15950 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1054 diff_507500_3274100# diff_727900_2842000# diff_622050_2844900# GND efet w=15950 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1055 GND diff_629300_2881150# diff_655400_3288600# GND efet w=44225 l=12325
+ ad=0 pd=0 as=1.86492e+09 ps=464000 
M1056 diff_627850_2752100# diff_627850_2752100# GND GND efet w=42050 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1057 GND diff_629300_2881150# diff_655400_3188550# GND efet w=44225 l=14500
+ ad=0 pd=0 as=1.91958e+09 ps=464000 
M1058 diff_627850_2752100# diff_627850_2752100# GND GND efet w=51475 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1059 diff_606100_2879700# diff_606100_2879700# GND GND efet w=31900 l=23200
+ ad=0 pd=0 as=0 ps=0 
M1060 diff_298700_3089950# diff_292900_3079800# diff_298700_3069650# GND efet w=13050 l=11600
+ ad=0 pd=0 as=1.09961e+09 ps=304500 
M1061 diff_323350_3089950# diff_292900_3079800# diff_323350_3071100# GND efet w=23200 l=11600
+ ad=0 pd=0 as=1.36242e+09 ps=298700 
M1062 diff_359600_3089950# diff_292900_3079800# diff_323350_3071100# GND efet w=17400 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1063 diff_378450_3143600# diff_292900_3079800# diff_323350_3071100# GND efet w=8700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1064 diff_292900_3079800# diff_320450_2669450# GND GND efet w=23200 l=12325
+ ad=1.89225e+08 pd=63800 as=0 ps=0 
M1065 GND diff_292900_3079800# diff_491550_2995700# GND efet w=125425 l=12325
+ ad=0 pd=0 as=9.56638e+08 ps=249400 
M1066 diff_298700_3069650# GND GND GND efet w=7975 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1067 diff_606100_2879700# diff_606100_2879700# GND GND efet w=33350 l=23925
+ ad=0 pd=0 as=0 ps=0 
M1068 GND GND diff_436450_2937700# GND efet w=10875 l=14500
+ ad=0 pd=0 as=3.04862e+08 ps=113100 
M1069 diff_507500_2950750# diff_436450_2937700# diff_491550_2995700# GND efet w=69600 l=11600
+ ad=-7.9851e+08 pd=881600 as=0 ps=0 
M1070 GND diff_292900_3079800# GND GND efet w=29000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1071 GND GND GND GND efet w=7975 l=67425
+ ad=0 pd=0 as=0 ps=0 
M1072 GND GND diff_507500_2950750# GND efet w=7250 l=27550
+ ad=0 pd=0 as=0 ps=0 
M1073 GND GND diff_323350_3071100# GND efet w=26100 l=18850
+ ad=0 pd=0 as=0 ps=0 
M1074 GND diff_436450_2937700# GND GND efet w=21750 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1075 diff_436450_2937700# GND GND GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1076 diff_507500_2950750# GND GND GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1077 GND GND diff_50750_3136350# GND efet w=90625 l=23925
+ ad=0 pd=0 as=0 ps=0 
M1078 diff_298700_3069650# GND diff_342200_2886950# GND efet w=14500 l=11600
+ ad=0 pd=0 as=4.56242e+08 ps=133400 
M1079 GND GND GND GND efet w=98600 l=27550
+ ad=0 pd=0 as=0 ps=0 
M1080 GND diff_1051250_3567000# diff_1044000_3564100# GND efet w=26100 l=14500
+ ad=0 pd=0 as=1.38765e+08 ps=66700 
M1081 diff_1000500_3543800# diff_978750_3526400# GND GND efet w=19575 l=10875
+ ad=1.7661e+08 pd=66700 as=0 ps=0 
M1082 diff_622050_2844900# diff_622050_2844900# diff_1000500_3543800# GND efet w=26825 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1083 diff_1044000_3564100# diff_1032400_2863750# diff_622050_2844900# GND efet w=26100 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1084 diff_622050_2844900# diff_622050_2844900# diff_1135350_3543800# GND efet w=27550 l=13050
+ ad=0 pd=0 as=1.7661e+08 ps=72500 
M1085 diff_1135350_3543800# diff_1115050_3526400# GND GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1086 diff_606100_2879700# diff_622050_2844900# GND GND efet w=72500 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1087 diff_627850_2752100# diff_914950_2865200# diff_916400_3567000# GND efet w=6525 l=12325
+ ad=0 pd=0 as=5.25625e+07 ps=31900 
M1088 diff_978750_3526400# diff_943950_2878250# diff_627850_2752100# GND efet w=7975 l=10875
+ ad=4.6255e+07 pd=31900 as=0 ps=0 
M1089 diff_606100_2879700# diff_914950_2865200# diff_916400_3472750# GND efet w=6525 l=12325
+ ad=0 pd=0 as=5.046e+07 ps=29000 
M1090 diff_978750_3509000# diff_943950_2878250# diff_606100_2879700# GND efet w=5800 l=10150
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M1091 diff_907700_3474200# diff_887400_2863750# diff_622050_2844900# GND efet w=27550 l=11600
+ ad=1.70302e+08 pd=69600 as=0 ps=0 
M1092 GND diff_916400_3472750# diff_907700_3474200# GND efet w=25375 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1093 diff_627850_2752100# diff_606100_2879700# diff_1051250_3567000# GND efet w=6525 l=12325
+ ad=0 pd=0 as=5.25625e+07 ps=31900 
M1094 diff_1115050_3526400# diff_622050_2844900# diff_627850_2752100# GND efet w=5800 l=11600
+ ad=4.41525e+07 pd=29000 as=0 ps=0 
M1095 diff_606100_2879700# diff_606100_2879700# diff_1051250_3474200# GND efet w=5075 l=13775
+ ad=0 pd=0 as=5.046e+07 ps=29000 
M1096 GND diff_622050_2844900# diff_606100_2879700# GND efet w=72500 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1097 diff_909150_3456800# diff_887400_2863750# diff_622050_2844900# GND efet w=24650 l=10875
+ ad=1.53482e+08 pd=66700 as=0 ps=0 
M1098 GND diff_916400_3459700# diff_909150_3456800# GND efet w=24650 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1099 diff_1000500_3474200# diff_978750_3509000# GND GND efet w=22475 l=13775
+ ad=1.87122e+08 pd=72500 as=0 ps=0 
M1100 diff_622050_2844900# diff_622050_2844900# diff_1000500_3474200# GND efet w=22475 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1101 diff_1044000_3472750# diff_1032400_2863750# diff_622050_2844900# GND efet w=26825 l=10875
+ ad=2.0184e+08 pd=69600 as=0 ps=0 
M1102 GND diff_1051250_3474200# diff_1044000_3472750# GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1103 diff_606100_2879700# diff_622050_2844900# GND GND efet w=71050 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1104 diff_606100_2879700# diff_914950_2865200# diff_916400_3459700# GND efet w=7975 l=12325
+ ad=0 pd=0 as=5.67675e+07 ps=37700 
M1105 diff_1000500_3436500# diff_978750_3419100# GND GND efet w=23925 l=15225
+ ad=1.87122e+08 pd=69600 as=0 ps=0 
M1106 diff_1115050_3509000# diff_622050_2844900# diff_606100_2879700# GND efet w=5800 l=13050
+ ad=5.25625e+07 pd=34800 as=0 ps=0 
M1107 GND diff_1048350_2488200# diff_622050_2844900# GND efet w=8700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1108 GND diff_320450_2669450# GND GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1109 GND diff_1489150_3117500# diff_1425350_3181300# GND efet w=17400 l=13050
+ ad=0 pd=0 as=1.11408e+09 ps=1.03936e+07 
M1110 GND diff_1425350_3181300# diff_1423900_3514800# GND efet w=63800 l=11600
+ ad=0 pd=0 as=-2.1336e+09 ps=580000 
M1111 GND GND diff_627850_2752100# GND efet w=6525 l=31175
+ ad=0 pd=0 as=0 ps=0 
M1112 GND GND GND GND efet w=101500 l=20300
+ ad=0 pd=0 as=0 ps=0 
M1113 GND GND diff_606100_2879700# GND efet w=6525 l=31175
+ ad=0 pd=0 as=0 ps=0 
M1114 GND diff_1052700_3456800# diff_1044000_3456800# GND efet w=25375 l=12325
+ ad=0 pd=0 as=1.91328e+08 ps=69600 
M1115 diff_622050_2844900# diff_622050_2844900# diff_1000500_3436500# GND efet w=19575 l=17400
+ ad=0 pd=0 as=0 ps=0 
M1116 diff_1044000_3456800# diff_1032400_2863750# diff_622050_2844900# GND efet w=26825 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1117 diff_1135350_3480000# diff_1115050_3509000# GND GND efet w=23925 l=13775
+ ad=1.82918e+08 pd=66700 as=0 ps=0 
M1118 diff_622050_2844900# diff_622050_2844900# diff_1135350_3480000# GND efet w=26825 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1119 GND diff_1048350_2488200# diff_622050_2844900# GND efet w=9425 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1120 GND GND diff_1423900_3514800# GND efet w=43500 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1121 diff_1425350_3181300# diff_1425350_3181300# GND GND efet w=41325 l=17400
+ ad=0 pd=0 as=0 ps=0 
M1122 GND GND GND GND efet w=7975 l=22475
+ ad=0 pd=0 as=0 ps=0 
M1123 diff_1135350_3436500# diff_1115050_3419100# GND GND efet w=23925 l=13775
+ ad=1.89225e+08 pd=69600 as=0 ps=0 
M1124 diff_622050_2844900# diff_622050_2844900# diff_1135350_3436500# GND efet w=28275 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1125 diff_978750_3419100# diff_943950_2878250# diff_606100_2879700# GND efet w=6525 l=10150
+ ad=5.4665e+07 pd=31900 as=0 ps=0 
M1126 diff_606100_2879700# diff_914950_2865200# diff_916400_3365450# GND efet w=5800 l=10150
+ ad=0 pd=0 as=5.046e+07 ps=29000 
M1127 diff_978750_3401700# diff_943950_2878250# diff_606100_2879700# GND efet w=5800 l=10150
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M1128 diff_907700_3365450# diff_887400_2863750# diff_622050_2844900# GND efet w=28275 l=10875
+ ad=1.72405e+08 pd=72500 as=0 ps=0 
M1129 GND diff_916400_3365450# diff_907700_3365450# GND efet w=24650 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1130 diff_606100_2879700# diff_606100_2879700# diff_1052700_3456800# GND efet w=4350 l=14500
+ ad=0 pd=0 as=5.4665e+07 ps=34800 
M1131 GND diff_1048350_2488200# diff_622050_2844900# GND efet w=9425 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1132 GND GND GND GND efet w=7975 l=21025
+ ad=0 pd=0 as=0 ps=0 
M1133 diff_1115050_3419100# diff_622050_2844900# diff_606100_2879700# GND efet w=5800 l=11600
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M1134 diff_606100_2879700# diff_606100_2879700# diff_1051250_3365450# GND efet w=5075 l=11600
+ ad=0 pd=0 as=5.046e+07 ps=29000 
M1135 diff_1115050_3401700# diff_622050_2844900# diff_606100_2879700# GND efet w=5800 l=11600
+ ad=5.4665e+07 pd=31900 as=0 ps=0 
M1136 GND diff_622050_2844900# diff_655400_3288600# GND efet w=63800 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1137 GND diff_622050_2844900# diff_627850_2752100# GND efet w=68875 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1138 diff_622050_2844900# diff_784450_2863750# diff_507500_3274100# GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1139 diff_909150_3349500# diff_887400_2863750# diff_622050_2844900# GND efet w=24650 l=10875
+ ad=1.53482e+08 pd=63800 as=0 ps=0 
M1140 GND diff_916400_3350950# diff_909150_3349500# GND efet w=24650 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1141 diff_999050_3374150# diff_978750_3401700# GND GND efet w=23925 l=13775
+ ad=1.7661e+08 pd=69600 as=0 ps=0 
M1142 diff_622050_2844900# diff_622050_2844900# diff_999050_3374150# GND efet w=21025 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1143 diff_1044000_3365450# diff_1032400_2863750# diff_622050_2844900# GND efet w=26825 l=10875
+ ad=1.97635e+08 pd=69600 as=0 ps=0 
M1144 GND diff_1051250_3365450# diff_1044000_3365450# GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1145 GND GND GND GND efet w=110925 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1146 GND GND diff_606100_2879700# GND efet w=7250 l=31900
+ ad=0 pd=0 as=0 ps=0 
M1147 GND GND diff_606100_2879700# GND efet w=6525 l=31175
+ ad=0 pd=0 as=0 ps=0 
M1148 diff_1135350_3372700# diff_1115050_3401700# GND GND efet w=23925 l=18125
+ ad=1.87122e+08 pd=69600 as=0 ps=0 
M1149 diff_1000500_3330650# diff_978750_3311800# GND GND efet w=22475 l=15225
+ ad=1.63995e+08 pd=66700 as=0 ps=0 
M1150 GND diff_1051250_3350950# diff_1044000_3346600# GND efet w=23925 l=12325
+ ad=0 pd=0 as=1.87122e+08 ps=66700 
M1151 diff_622050_2844900# diff_622050_2844900# diff_1000500_3330650# GND efet w=21750 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1152 diff_1044000_3346600# diff_1032400_2863750# diff_622050_2844900# GND efet w=25375 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1153 diff_622050_2844900# diff_622050_2844900# diff_1135350_3372700# GND efet w=21750 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1154 GND diff_1048350_2488200# diff_622050_2844900# GND efet w=8700 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1155 GND GND diff_1425350_3394450# GND efet w=43500 l=13050
+ ad=0 pd=0 as=2.07937e+09 ps=559700 
M1156 diff_1425350_3181300# diff_1425350_3181300# GND GND efet w=41325 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1157 diff_1425350_3181300# diff_1425350_3181300# GND GND efet w=8700 l=18125
+ ad=0 pd=0 as=0 ps=0 
M1158 diff_1425350_3181300# diff_1425350_3181300# GND GND efet w=59450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1159 diff_1673300_3561200# diff_1425350_3181300# diff_1425350_3181300# GND efet w=18850 l=18850
+ ad=1.40868e+08 pd=63800 as=0 ps=0 
M1160 GND GND diff_1673300_3561200# GND efet w=25375 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1161 diff_1764650_3543800# diff_1742900_3524950# GND GND efet w=24650 l=14500
+ ad=1.3456e+08 pd=60900 as=0 ps=0 
M1162 diff_1425350_3181300# diff_1425350_3181300# diff_1764650_3543800# GND efet w=19575 l=18125
+ ad=0 pd=0 as=0 ps=0 
M1163 diff_1808150_3561200# diff_1425350_3181300# diff_1425350_3181300# GND efet w=21750 l=17400
+ ad=1.682e+08 pd=63800 as=0 ps=0 
M1164 GND diff_1815400_3526400# diff_1808150_3561200# GND efet w=23925 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1165 diff_1899500_3543800# diff_1877750_3524950# GND GND efet w=25375 l=16675
+ ad=1.30355e+08 pd=60900 as=0 ps=0 
M1166 diff_1425350_3181300# diff_1425350_3181300# diff_1899500_3543800# GND efet w=20300 l=18125
+ ad=0 pd=0 as=0 ps=0 
M1167 diff_1943000_3564100# diff_1425350_3181300# diff_1425350_3181300# GND efet w=21025 l=19575
+ ad=1.36662e+08 pd=66700 as=0 ps=0 
M1168 GND diff_1948800_3562650# diff_1943000_3564100# GND efet w=26825 l=19575
+ ad=0 pd=0 as=0 ps=0 
M1169 diff_2034350_3542350# diff_2012600_3524950# GND GND efet w=25375 l=13775
+ ad=1.2615e+08 pd=69600 as=0 ps=0 
M1170 diff_1423900_3514800# diff_1687800_3075450# GND GND efet w=5800 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1171 diff_1742900_3524950# diff_1718250_3075450# diff_1423900_3514800# GND efet w=5800 l=11600
+ ad=4.41525e+07 pd=29000 as=0 ps=0 
M1172 diff_1423900_3514800# diff_1829900_3075450# diff_1815400_3526400# GND efet w=6525 l=12325
+ ad=0 pd=0 as=4.6255e+07 ps=31900 
M1173 diff_1425350_3181300# diff_1687800_3075450# diff_1679100_3471300# GND efet w=5800 l=11600
+ ad=0 pd=0 as=4.205e+07 ps=26100 
M1174 diff_1742900_3507550# diff_1718250_3075450# diff_1425350_3181300# GND efet w=5800 l=11600
+ ad=4.6255e+07 pd=31900 as=0 ps=0 
M1175 diff_1671850_3471300# diff_1425350_3181300# diff_1425350_3181300# GND efet w=27550 l=13050
+ ad=1.7661e+08 pd=69600 as=0 ps=0 
M1176 GND diff_1679100_3471300# diff_1671850_3471300# GND efet w=24650 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1177 diff_1877750_3524950# diff_1858900_3075450# diff_1423900_3514800# GND efet w=5800 l=11600
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M1178 GND diff_1679100_3456800# diff_1671850_3456800# GND efet w=23925 l=13775
+ ad=0 pd=0 as=1.63995e+08 ps=66700 
M1179 GND diff_320450_2669450# GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1180 diff_1135350_3330650# diff_1113600_3311800# GND GND efet w=24650 l=16675
+ ad=1.7661e+08 pd=66700 as=0 ps=0 
M1181 diff_622050_2844900# diff_622050_2844900# diff_1135350_3330650# GND efet w=19575 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1182 diff_655400_3288600# diff_914950_2865200# diff_916400_3350950# GND efet w=7975 l=12325
+ ad=0 pd=0 as=6.728e+07 ps=34800 
M1183 diff_978750_3311800# diff_943950_2878250# diff_655400_3288600# GND efet w=5800 l=12325
+ ad=5.887e+07 pd=37700 as=0 ps=0 
M1184 diff_627850_2752100# diff_914950_2865200# diff_916400_3258150# GND efet w=5800 l=10150
+ ad=0 pd=0 as=5.887e+07 ps=31900 
M1185 diff_978750_3294400# diff_943950_2878250# diff_627850_2752100# GND efet w=5800 l=10150
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M1186 diff_907700_3258150# diff_887400_2863750# diff_622050_2844900# GND efet w=27550 l=10875
+ ad=1.74508e+08 pd=69600 as=0 ps=0 
M1187 GND diff_916400_3258150# diff_907700_3258150# GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1188 diff_655400_3288600# diff_606100_2879700# diff_1051250_3350950# GND efet w=6525 l=10875
+ ad=0 pd=0 as=5.4665e+07 ps=34800 
M1189 diff_1113600_3311800# diff_622050_2844900# diff_655400_3288600# GND efet w=5800 l=10150
+ ad=5.887e+07 pd=31900 as=0 ps=0 
M1190 diff_627850_2752100# diff_606100_2879700# diff_1051250_3258150# GND efet w=5800 l=10150
+ ad=0 pd=0 as=5.046e+07 ps=29000 
M1191 diff_1113600_3294400# diff_622050_2844900# diff_627850_2752100# GND efet w=5800 l=10150
+ ad=5.887e+07 pd=31900 as=0 ps=0 
M1192 GND diff_622050_2844900# diff_627850_2752100# GND efet w=73225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1193 diff_622050_2844900# diff_784450_2863750# diff_507500_3229150# GND efet w=14500 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1194 diff_507500_3229150# diff_727900_2842000# diff_622050_2844900# GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1195 diff_907700_3243650# diff_887400_2863750# diff_622050_2844900# GND efet w=26825 l=10875
+ ad=1.5979e+08 pd=66700 as=0 ps=0 
M1196 GND diff_916400_3243650# diff_907700_3243650# GND efet w=24650 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1197 diff_1000500_3261050# diff_978750_3294400# GND GND efet w=23200 l=14500
+ ad=1.82918e+08 pd=66700 as=0 ps=0 
M1198 diff_622050_2844900# diff_622050_2844900# diff_1000500_3261050# GND efet w=26100 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1199 diff_1044000_3258150# diff_1032400_2863750# diff_622050_2844900# GND efet w=27550 l=11600
+ ad=1.99738e+08 pd=69600 as=0 ps=0 
M1200 GND diff_1051250_3258150# diff_1044000_3258150# GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1201 GND diff_1048350_2488200# diff_622050_2844900# GND efet w=8700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1202 GND diff_320450_2669450# GND GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1203 diff_622050_2844900# diff_622050_2844900# diff_507500_3229150# GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1204 diff_622050_2844900# diff_622050_2844900# diff_507500_2950750# GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1205 diff_655400_3188550# diff_622050_2844900# GND GND efet w=65975 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1206 diff_627850_2752100# diff_914950_2865200# diff_916400_3243650# GND efet w=6525 l=13050
+ ad=0 pd=0 as=5.67675e+07 ps=34800 
M1207 diff_999050_3223350# diff_978750_3204500# GND GND efet w=23200 l=14500
+ ad=1.95532e+08 pd=66700 as=0 ps=0 
M1208 GND diff_1051250_3243650# diff_1042550_3242200# GND efet w=26100 l=13050
+ ad=0 pd=0 as=1.82918e+08 ps=69600 
M1209 diff_622050_2844900# diff_622050_2844900# diff_999050_3223350# GND efet w=24650 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1210 diff_1042550_3242200# diff_1032400_2863750# diff_622050_2844900# GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1211 diff_1135350_3263950# diff_1113600_3294400# GND GND efet w=24650 l=13050
+ ad=1.80815e+08 pd=66700 as=0 ps=0 
M1212 diff_622050_2844900# diff_622050_2844900# diff_1135350_3263950# GND efet w=21750 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1213 GND GND diff_655400_3288600# GND efet w=6525 l=29725
+ ad=0 pd=0 as=0 ps=0 
M1214 GND GND diff_1425350_3181300# GND efet w=43500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1215 GND GND GND GND efet w=100775 l=19575
+ ad=0 pd=0 as=0 ps=0 
M1216 GND GND diff_627850_2752100# GND efet w=6525 l=29725
+ ad=0 pd=0 as=0 ps=0 
M1217 GND diff_1048350_2488200# diff_622050_2844900# GND efet w=10150 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1218 diff_1425350_3181300# diff_1425350_3181300# GND GND efet w=7975 l=18125
+ ad=0 pd=0 as=0 ps=0 
M1219 GND diff_1489150_3117500# diff_1425350_3181300# GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1220 GND diff_1489150_3117500# diff_1425350_3181300# GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1221 diff_1135350_3221900# diff_1113600_3204500# GND GND efet w=25375 l=13775
+ ad=1.78712e+08 pd=66700 as=0 ps=0 
M1222 diff_978750_3204500# diff_943950_2878250# diff_627850_2752100# GND efet w=5800 l=11600
+ ad=5.25625e+07 pd=31900 as=0 ps=0 
M1223 diff_978750_3187100# diff_943950_2878250# diff_655400_3188550# GND efet w=5800 l=13050
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M1224 diff_655400_3188550# diff_914950_2865200# diff_916400_3150850# GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.046e+07 ps=29000 
M1225 diff_907700_3150850# diff_887400_2863750# diff_622050_2844900# GND efet w=28275 l=10875
+ ad=1.80815e+08 pd=69600 as=0 ps=0 
M1226 GND diff_916400_3150850# diff_907700_3150850# GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1227 diff_627850_2752100# diff_606100_2879700# diff_1051250_3243650# GND efet w=5800 l=10150
+ ad=0 pd=0 as=5.25625e+07 ps=31900 
M1228 diff_622050_2844900# diff_622050_2844900# diff_1135350_3221900# GND efet w=21025 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1229 diff_1113600_3204500# diff_622050_2844900# diff_627850_2752100# GND efet w=5800 l=10150
+ ad=5.25625e+07 pd=31900 as=0 ps=0 
M1230 diff_655400_3188550# diff_606100_2879700# diff_1051250_3150850# GND efet w=5800 l=10150
+ ad=0 pd=0 as=5.046e+07 ps=29000 
M1231 diff_999050_3156650# diff_978750_3187100# GND GND efet w=23925 l=12325
+ ad=2.03942e+08 pd=72500 as=0 ps=0 
M1232 GND diff_916400_3134900# diff_907700_3136350# GND efet w=25375 l=13775
+ ad=0 pd=0 as=1.61892e+08 ps=66700 
M1233 GND diff_622050_2844900# diff_606100_2879700# GND efet w=69600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1234 diff_907700_3136350# diff_887400_2863750# diff_622050_2844900# GND efet w=25375 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1235 diff_622050_2844900# diff_622050_2844900# diff_999050_3156650# GND efet w=26825 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1236 diff_1044000_3150850# diff_1032400_2863750# diff_622050_2844900# GND efet w=26100 l=11600
+ ad=1.87122e+08 pd=72500 as=0 ps=0 
M1237 GND diff_1051250_3150850# diff_1044000_3150850# GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1238 diff_1113600_3187100# diff_622050_2844900# diff_655400_3188550# GND efet w=5800 l=11600
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M1239 diff_1135350_3156650# diff_1113600_3187100# GND GND efet w=23925 l=13775
+ ad=1.682e+08 pd=63800 as=0 ps=0 
M1240 diff_622050_2844900# diff_622050_2844900# diff_1135350_3156650# GND efet w=19575 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1241 diff_606100_2879700# diff_622050_2844900# GND GND efet w=68150 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1242 diff_606100_2879700# diff_914950_2865200# diff_916400_3134900# GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.046e+07 ps=29000 
M1243 diff_999050_3120400# diff_978750_3097200# GND GND efet w=24650 l=13050
+ ad=1.91328e+08 pd=72500 as=0 ps=0 
M1244 GND diff_1051250_3136350# diff_1044000_3132000# GND efet w=23925 l=12325
+ ad=0 pd=0 as=1.89225e+08 ps=66700 
M1245 diff_622050_2844900# diff_622050_2844900# diff_999050_3120400# GND efet w=25375 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1246 diff_1044000_3132000# diff_1032400_2863750# diff_622050_2844900# GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1247 GND GND GND GND efet w=7250 l=20300
+ ad=0 pd=0 as=0 ps=0 
M1248 GND diff_1048350_2488200# diff_622050_2844900# GND efet w=9425 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1249 GND GND diff_627850_2752100# GND efet w=5800 l=30450
+ ad=0 pd=0 as=0 ps=0 
M1250 diff_1328200_3190000# GND GND GND efet w=7975 l=20300
+ ad=1.98476e+09 pd=501700 as=0 ps=0 
M1251 GND diff_1328200_3190000# diff_1328200_3190000# GND efet w=110925 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1252 diff_1425350_3181300# diff_1425350_3181300# GND GND efet w=39875 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1253 GND diff_1425350_3181300# diff_1425350_3181300# GND efet w=59450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1254 diff_1425350_3394450# diff_1425350_3181300# GND GND efet w=60175 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1255 diff_1671850_3456800# diff_1425350_3181300# diff_1425350_3181300# GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1256 diff_1763200_3478550# diff_1742900_3507550# GND GND efet w=29000 l=14500
+ ad=1.63995e+08 pd=72500 as=0 ps=0 
M1257 diff_1425350_3181300# diff_1425350_3181300# diff_1763200_3478550# GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1258 diff_1806700_3472750# diff_1425350_3181300# diff_1425350_3181300# GND efet w=26100 l=13050
+ ad=1.682e+08 pd=66700 as=0 ps=0 
M1259 diff_1425350_3181300# diff_1829900_3075450# diff_1815400_3469850# GND efet w=5800 l=11600
+ ad=0 pd=0 as=4.205e+07 ps=26100 
M1260 GND diff_1815400_3469850# diff_1806700_3472750# GND efet w=21750 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1261 diff_1763200_3436500# diff_1742900_3417650# GND GND efet w=26825 l=15225
+ ad=1.682e+08 pd=75400 as=0 ps=0 
M1262 diff_1425350_3181300# diff_1687800_3075450# diff_1679100_3456800# GND efet w=5800 l=11600
+ ad=0 pd=0 as=4.83575e+07 ps=31900 
M1263 diff_1877750_3507550# diff_1858900_3075450# diff_1425350_3181300# GND efet w=5800 l=11600
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M1264 diff_1899500_3477100# diff_1877750_3507550# GND GND efet w=24650 l=15950
+ ad=1.3456e+08 pd=63800 as=0 ps=0 
M1265 diff_1425350_3181300# diff_2025650_3074000# diff_2034350_3542350# GND efet w=30450 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1266 diff_2077850_3561200# diff_1425350_3181300# diff_1425350_3181300# GND efet w=27550 l=13050
+ ad=1.30355e+08 pd=66700 as=0 ps=0 
M1267 GND diff_2083650_3562650# diff_2077850_3561200# GND efet w=26825 l=18850
+ ad=0 pd=0 as=0 ps=0 
M1268 diff_2169200_3542350# diff_2148900_3524950# GND GND efet w=27550 l=13050
+ ad=1.19842e+08 pd=66700 as=0 ps=0 
M1269 diff_1425350_3181300# diff_2166300_3074000# diff_2169200_3542350# GND efet w=29000 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1270 diff_1425350_3181300# diff_1425350_3181300# diff_1899500_3477100# GND efet w=23925 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1271 diff_1423900_3514800# diff_1425350_3181300# diff_1948800_3562650# GND efet w=5800 l=13050
+ ad=0 pd=0 as=4.41525e+07 ps=29000 
M1272 diff_2012600_3524950# diff_1425350_3181300# diff_1423900_3514800# GND efet w=7975 l=12325
+ ad=3.99475e+07 pd=29000 as=0 ps=0 
M1273 diff_1425350_3181300# diff_1425350_3181300# diff_1950250_3469850# GND efet w=7250 l=13050
+ ad=0 pd=0 as=4.205e+07 ps=26100 
M1274 GND diff_1950250_3469850# diff_1943000_3471300# GND efet w=21750 l=14500
+ ad=0 pd=0 as=1.682e+08 ps=63800 
M1275 diff_2012600_3507550# diff_1425350_3181300# diff_1425350_3181300# GND efet w=6525 l=12325
+ ad=4.6255e+07 pd=29000 as=0 ps=0 
M1276 diff_1943000_3471300# diff_1425350_3181300# diff_1425350_3181300# GND efet w=20300 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1277 GND diff_1815400_3456800# diff_1806700_3456800# GND efet w=23200 l=15225
+ ad=0 pd=0 as=1.70302e+08 ps=69600 
M1278 diff_1425350_3181300# diff_1425350_3181300# diff_1763200_3436500# GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1279 diff_1806700_3456800# diff_1425350_3181300# diff_1425350_3181300# GND efet w=25375 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1280 diff_1423900_3514800# diff_2106850_3184200# diff_2083650_3562650# GND efet w=5800 l=13050
+ ad=0 pd=0 as=4.205e+07 ps=26100 
M1281 diff_2148900_3524950# diff_1425350_3181300# diff_1423900_3514800# GND efet w=5800 l=14500
+ ad=3.364e+07 pd=23200 as=0 ps=0 
M1282 diff_1425350_3181300# diff_2106850_3184200# diff_2086550_3468400# GND efet w=7250 l=13775
+ ad=0 pd=0 as=4.6255e+07 ps=29000 
M1283 diff_1898050_3435050# diff_1877750_3417650# GND GND efet w=25375 l=16675
+ ad=1.66098e+08 pd=75400 as=0 ps=0 
M1284 diff_1425350_3181300# diff_1425350_3181300# diff_1898050_3435050# GND efet w=27550 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1285 diff_1742900_3417650# diff_1718250_3075450# diff_1425350_3181300# GND efet w=5800 l=11600
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M1286 diff_1425350_3394450# diff_1687800_3075450# diff_1680550_3362550# GND efet w=5800 l=11600
+ ad=0 pd=0 as=4.205e+07 ps=26100 
M1287 diff_1742900_3400250# diff_1718250_3075450# diff_1425350_3394450# GND efet w=5800 l=11600
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M1288 diff_1671850_3366900# diff_1425350_3181300# diff_1425350_3181300# GND efet w=27550 l=11600
+ ad=1.66098e+08 pd=66700 as=0 ps=0 
M1289 GND diff_1680550_3362550# diff_1671850_3366900# GND efet w=23200 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1290 diff_1425350_3181300# diff_1829900_3075450# diff_1815400_3456800# GND efet w=6525 l=10875
+ ad=0 pd=0 as=4.83575e+07 ps=31900 
M1291 diff_1943000_3453900# diff_1425350_3181300# diff_1425350_3181300# GND efet w=21025 l=17400
+ ad=1.74508e+08 pd=66700 as=0 ps=0 
M1292 GND diff_1950250_3456800# diff_1943000_3453900# GND efet w=22475 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1293 diff_2034350_3475650# diff_2012600_3507550# GND GND efet w=26825 l=13775
+ ad=1.28252e+08 pd=63800 as=0 ps=0 
M1294 diff_1425350_3181300# diff_2025650_3074000# diff_2034350_3475650# GND efet w=25375 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1295 diff_2077850_3471300# diff_1425350_3181300# diff_1425350_3181300# GND efet w=21025 l=16675
+ ad=1.7661e+08 pd=63800 as=0 ps=0 
M1296 GND diff_2086550_3468400# diff_2077850_3471300# GND efet w=20300 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1297 GND diff_1425350_3181300# diff_1425350_3181300# GND efet w=7975 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1298 diff_2034350_3435050# diff_2012600_3417650# GND GND efet w=26100 l=13050
+ ad=1.36662e+08 pd=66700 as=0 ps=0 
M1299 diff_1425350_3181300# diff_2025650_3074000# diff_2034350_3435050# GND efet w=26100 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1300 diff_2169200_3475650# GND GND GND efet w=25375 l=13775
+ ad=1.24048e+08 pd=63800 as=0 ps=0 
M1301 diff_1425350_3181300# diff_2166300_3074000# diff_2169200_3475650# GND efet w=26100 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1302 diff_1877750_3417650# diff_1858900_3075450# diff_1425350_3181300# GND efet w=5800 l=11600
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M1303 diff_1425350_3394450# diff_1829900_3075450# diff_1815400_3362550# GND efet w=5800 l=10875
+ ad=0 pd=0 as=4.205e+07 ps=26100 
M1304 diff_1877750_3400250# diff_1858900_3075450# diff_1425350_3394450# GND efet w=5800 l=11600
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M1305 diff_1763200_3387200# diff_1742900_3400250# GND GND efet w=24650 l=13050
+ ad=1.61892e+08 pd=72500 as=0 ps=0 
M1306 GND diff_1680550_3348050# diff_1673300_3346600# GND efet w=23925 l=13775
+ ad=0 pd=0 as=1.63995e+08 ps=63800 
M1307 GND diff_1425350_3181300# diff_1425350_3181300# GND efet w=53650 l=17400
+ ad=0 pd=0 as=0 ps=0 
M1308 diff_1673300_3346600# diff_1425350_3181300# diff_1425350_3181300# GND efet w=25375 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1309 diff_1425350_3181300# diff_1425350_3181300# diff_1763200_3387200# GND efet w=28275 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1310 diff_1808150_3364000# diff_1425350_3181300# diff_1425350_3181300# GND efet w=26100 l=11600
+ ad=1.7661e+08 pd=66700 as=0 ps=0 
M1311 GND diff_1815400_3362550# diff_1808150_3364000# GND efet w=23200 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1312 diff_1425350_3181300# diff_1425350_3181300# diff_1950250_3456800# GND efet w=5800 l=13050
+ ad=0 pd=0 as=4.41525e+07 ps=29000 
M1313 diff_2077850_3453900# diff_1425350_3181300# diff_1425350_3181300# GND efet w=20300 l=15950
+ ad=1.74508e+08 pd=66700 as=0 ps=0 
M1314 GND diff_2086550_3417650# diff_2077850_3453900# GND efet w=21025 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1315 GND diff_2072050_2521550# diff_1425350_3181300# GND efet w=11600 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1316 GND GND diff_1423900_3514800# GND efet w=8700 l=33350
+ ad=0 pd=0 as=0 ps=0 
M1317 GND GND diff_1425350_3181300# GND efet w=8700 l=33350
+ ad=0 pd=0 as=0 ps=0 
M1318 GND diff_2072050_2521550# diff_1425350_3181300# GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1319 diff_2169200_3435050# diff_2148900_3417650# GND GND efet w=26100 l=13050
+ ad=1.32458e+08 pd=63800 as=0 ps=0 
M1320 diff_2012600_3417650# diff_1425350_3181300# diff_1425350_3181300# GND efet w=5800 l=11600
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M1321 diff_1425350_3394450# diff_1425350_3181300# diff_1950250_3362550# GND efet w=5800 l=14500
+ ad=0 pd=0 as=4.205e+07 ps=26100 
M1322 diff_1425350_3181300# diff_1425350_3181300# GND GND efet w=62350 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1323 diff_1425350_3181300# diff_1425350_3181300# GND GND efet w=7975 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1324 diff_1764650_3329200# diff_1742900_3310350# GND GND efet w=23200 l=13050
+ ad=1.66098e+08 pd=63800 as=0 ps=0 
M1325 diff_1425350_3181300# diff_1425350_3181300# diff_1764650_3329200# GND efet w=25375 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1326 diff_1808150_3346600# diff_1425350_3181300# diff_1425350_3181300# GND efet w=24650 l=11600
+ ad=1.66098e+08 pd=63800 as=0 ps=0 
M1327 GND diff_1815400_3348050# diff_1808150_3346600# GND efet w=23200 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1328 diff_1899500_3369800# diff_1877750_3400250# GND GND efet w=23925 l=13775
+ ad=1.5138e+08 pd=69600 as=0 ps=0 
M1329 diff_1425350_3181300# diff_1425350_3181300# diff_1899500_3369800# GND efet w=26825 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1330 diff_1943000_3364000# diff_1425350_3181300# diff_1425350_3181300# GND efet w=21750 l=15950
+ ad=1.82918e+08 pd=66700 as=0 ps=0 
M1331 GND diff_1950250_3362550# diff_1943000_3364000# GND efet w=23200 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1332 diff_2012600_3400250# diff_1425350_3181300# diff_1425350_3394450# GND efet w=7250 l=13050
+ ad=5.046e+07 pd=31900 as=0 ps=0 
M1333 diff_1425350_3181300# diff_2106850_3184200# diff_2086550_3417650# GND efet w=5800 l=13050
+ ad=0 pd=0 as=4.205e+07 ps=26100 
M1334 diff_1425350_3181300# diff_2166300_3074000# diff_2169200_3435050# GND efet w=26100 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1335 diff_2148900_3417650# diff_1425350_3181300# diff_1425350_3181300# GND efet w=6525 l=13775
+ ad=4.205e+07 pd=26100 as=0 ps=0 
M1336 diff_1425350_3394450# diff_2106850_3184200# diff_2086550_3362550# GND efet w=7250 l=13050
+ ad=0 pd=0 as=5.25625e+07 ps=29000 
M1337 diff_2034350_3369800# diff_2012600_3400250# GND GND efet w=23200 l=13775
+ ad=1.36662e+08 pd=66700 as=0 ps=0 
M1338 diff_1425350_3181300# diff_2025650_3074000# diff_2034350_3369800# GND efet w=25375 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1339 diff_2077850_3364000# diff_1425350_3181300# diff_1425350_3181300# GND efet w=20300 l=16675
+ ad=1.78712e+08 pd=66700 as=0 ps=0 
M1340 GND diff_2086550_3362550# diff_2077850_3364000# GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1341 diff_1899500_3329200# diff_1877750_3314700# GND GND efet w=23200 l=14500
+ ad=1.61892e+08 pd=63800 as=0 ps=0 
M1342 diff_1425350_3181300# diff_1687800_3075450# diff_1680550_3348050# GND efet w=5800 l=12325
+ ad=0 pd=0 as=3.7845e+07 ps=29000 
M1343 diff_1742900_3310350# diff_1718250_3075450# diff_1425350_3181300# GND efet w=6525 l=12325
+ ad=5.4665e+07 pd=34800 as=0 ps=0 
M1344 diff_1425350_3181300# diff_1687800_3075450# diff_1680550_3256700# GND efet w=7975 l=10875
+ ad=0 pd=0 as=4.6255e+07 ps=31900 
M1345 diff_1742900_3292950# diff_1718250_3075450# diff_1425350_3181300# GND efet w=5800 l=11600
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M1346 diff_1673300_3258150# diff_1425350_3181300# diff_1425350_3181300# GND efet w=24650 l=11600
+ ad=1.63995e+08 pd=63800 as=0 ps=0 
M1347 GND diff_1680550_3256700# diff_1673300_3258150# GND efet w=23200 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1348 diff_1425350_3181300# diff_1425350_3181300# diff_1899500_3329200# GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1349 diff_1943000_3346600# diff_1425350_3181300# diff_1425350_3181300# GND efet w=20300 l=15950
+ ad=1.682e+08 pd=63800 as=0 ps=0 
M1350 GND diff_1950250_3349500# diff_1943000_3346600# GND efet w=23925 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1351 diff_2148900_3398800# diff_1425350_3181300# diff_1425350_3394450# GND efet w=7975 l=15225
+ ad=5.4665e+07 pd=31900 as=0 ps=0 
M1352 diff_2169200_3368350# diff_2148900_3398800# GND GND efet w=27550 l=14500
+ ad=1.2615e+08 pd=63800 as=0 ps=0 
M1353 diff_2034350_3329200# diff_2014050_3310350# GND GND efet w=23200 l=14500
+ ad=1.53482e+08 pd=63800 as=0 ps=0 
M1354 diff_1425350_3181300# diff_1829900_3075450# diff_1815400_3348050# GND efet w=5800 l=13050
+ ad=0 pd=0 as=4.41525e+07 ps=29000 
M1355 diff_1877750_3314700# diff_1858900_3075450# diff_1425350_3181300# GND efet w=7250 l=10875
+ ad=4.41525e+07 pd=29000 as=0 ps=0 
M1356 diff_1425350_3181300# diff_1829900_3075450# diff_1816850_3255250# GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.046e+07 ps=29000 
M1357 GND diff_1680550_3242200# diff_1673300_3240750# GND efet w=23925 l=13775
+ ad=0 pd=0 as=1.61892e+08 ps=63800 
M1358 GND GND diff_655400_3188550# GND efet w=5800 l=30450
+ ad=0 pd=0 as=0 ps=0 
M1359 GND diff_1048350_2488200# diff_622050_2844900# GND efet w=10875 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1360 diff_1328200_3190000# diff_320450_2669450# GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1361 GND GND diff_1425350_3181300# GND efet w=46400 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1362 diff_1425350_3181300# diff_1425350_3181300# GND GND efet w=39875 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1363 diff_1135350_3116050# diff_1113600_3097200# GND GND efet w=23925 l=15225
+ ad=1.72405e+08 pd=66700 as=0 ps=0 
M1364 diff_978750_3097200# diff_943950_2878250# diff_606100_2879700# GND efet w=5800 l=11600
+ ad=5.25625e+07 pd=31900 as=0 ps=0 
M1365 diff_622050_2844900# diff_622050_2844900# diff_1135350_3116050# GND efet w=20300 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1366 diff_606100_2879700# diff_606100_2879700# diff_1051250_3136350# GND efet w=5800 l=10150
+ ad=0 pd=0 as=5.4665e+07 ps=31900 
M1367 diff_1113600_3097200# diff_622050_2844900# diff_606100_2879700# GND efet w=5800 l=10150
+ ad=5.25625e+07 pd=31900 as=0 ps=0 
M1368 diff_606100_2879700# diff_914950_2865200# diff_916400_3043550# GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.046e+07 ps=29000 
M1369 diff_907700_3043550# diff_887400_2863750# diff_622050_2844900# GND efet w=27550 l=10875
+ ad=1.80815e+08 pd=69600 as=0 ps=0 
M1370 GND diff_916400_3043550# diff_907700_3043550# GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1371 diff_978750_3079800# diff_943950_2878250# diff_606100_2879700# GND efet w=5800 l=11600
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M1372 diff_999050_3049350# diff_978750_3079800# GND GND efet w=23925 l=13775
+ ad=1.78712e+08 pd=69600 as=0 ps=0 
M1373 diff_606100_2879700# diff_606100_2879700# diff_1051250_3043550# GND efet w=5800 l=10150
+ ad=0 pd=0 as=5.046e+07 ps=29000 
M1374 GND diff_622050_2844900# diff_655400_2966700# GND efet w=68150 l=11600
+ ad=0 pd=0 as=1.97215e+09 ps=475600 
M1375 GND diff_916400_3029050# diff_907700_3027600# GND efet w=24650 l=14500
+ ad=0 pd=0 as=1.682e+08 ps=66700 
M1376 diff_507500_2950750# diff_727900_2842000# diff_622050_2844900# GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1377 GND diff_629300_2881150# diff_655400_2966700# GND efet w=43500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1378 diff_627850_2752100# diff_627850_2752100# GND GND efet w=43500 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1379 GND GND diff_342200_2886950# GND efet w=7250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1380 diff_488650_2876800# diff_342200_2886950# GND GND efet w=29000 l=11600
+ ad=5.7188e+08 pd=162400 as=0 ps=0 
M1381 diff_907700_3027600# diff_887400_2863750# diff_622050_2844900# GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1382 diff_622050_2844900# diff_622050_2844900# diff_999050_3049350# GND efet w=25375 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1383 diff_1044000_3043550# diff_1032400_2863750# diff_622050_2844900# GND efet w=26100 l=11600
+ ad=1.74508e+08 pd=72500 as=0 ps=0 
M1384 GND diff_1051250_3043550# diff_1044000_3043550# GND efet w=23925 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1385 diff_1113600_3079800# diff_622050_2844900# diff_606100_2879700# GND efet w=5800 l=10875
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M1386 diff_1135350_3047900# diff_1113600_3079800# GND GND efet w=22475 l=15225
+ ad=1.70302e+08 pd=63800 as=0 ps=0 
M1387 diff_1000500_3008750# diff_978750_2989900# GND GND efet w=21750 l=14500
+ ad=1.63995e+08 pd=63800 as=0 ps=0 
M1388 diff_622050_2844900# diff_622050_2844900# diff_1000500_3008750# GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1389 GND diff_622050_2844900# diff_627850_2752100# GND efet w=68875 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1390 diff_622050_2844900# diff_784450_2863750# diff_507500_2950750# GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1391 diff_655400_2966700# diff_914950_2865200# diff_916400_3029050# GND efet w=6525 l=13775
+ ad=0 pd=0 as=5.25625e+07 ps=31900 
M1392 diff_1044000_3024700# diff_1032400_2863750# diff_622050_2844900# GND efet w=24650 l=11600
+ ad=1.61892e+08 pd=66700 as=0 ps=0 
M1393 GND diff_1051250_3029050# diff_1044000_3024700# GND efet w=23200 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1394 diff_622050_2844900# diff_622050_2844900# diff_1135350_3047900# GND efet w=20300 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1395 GND diff_1048350_2488200# diff_622050_2844900# GND efet w=8700 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1396 diff_1425350_3181300# diff_1425350_3181300# diff_1328200_3190000# GND efet w=8700 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1397 diff_1328200_3190000# diff_1489150_3117500# diff_1425350_3181300# GND efet w=15225 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1398 GND diff_1425350_3181300# diff_1425350_3181300# GND efet w=59450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1399 diff_1673300_3240750# diff_1425350_3181300# diff_1425350_3181300# GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1400 diff_1764650_3262500# diff_1742900_3292950# GND GND efet w=23925 l=13775
+ ad=1.66098e+08 pd=63800 as=0 ps=0 
M1401 diff_1425350_3181300# diff_1425350_3181300# diff_1764650_3262500# GND efet w=21025 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1402 diff_1808150_3258150# diff_1425350_3181300# diff_1425350_3181300# GND efet w=24650 l=13050
+ ad=1.78712e+08 pd=69600 as=0 ps=0 
M1403 GND diff_1816850_3255250# diff_1808150_3258150# GND efet w=25375 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1404 diff_1764650_3221900# diff_1742900_3204500# GND GND efet w=23200 l=13050
+ ad=1.70302e+08 pd=63800 as=0 ps=0 
M1405 diff_1879200_3292950# diff_1858900_3075450# diff_1425350_3181300# GND efet w=5800 l=11600
+ ad=4.41525e+07 pd=29000 as=0 ps=0 
M1406 diff_1425350_3181300# diff_2025650_3074000# diff_2034350_3329200# GND efet w=25375 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1407 diff_2077850_3346600# diff_1425350_3181300# diff_1425350_3181300# GND efet w=22475 l=16675
+ ad=1.78712e+08 pd=69600 as=0 ps=0 
M1408 GND diff_2086550_3310350# diff_2077850_3346600# GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1409 diff_1425350_3181300# diff_1425350_3181300# diff_1950250_3349500# GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.046e+07 ps=29000 
M1410 diff_2014050_3310350# diff_1425350_3181300# diff_1425350_3181300# GND efet w=6525 l=13050
+ ad=4.205e+07 pd=26100 as=0 ps=0 
M1411 diff_1425350_3181300# diff_2166300_3074000# diff_2169200_3368350# GND efet w=25375 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1412 GND diff_2072050_2521550# diff_1425350_3181300# GND efet w=11600 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1413 GND GND diff_1425350_3181300# GND efet w=7250 l=37700
+ ad=0 pd=0 as=0 ps=0 
M1414 GND GND diff_1425350_3394450# GND efet w=7975 l=35525
+ ad=0 pd=0 as=0 ps=0 
M1415 GND diff_2072050_2521550# diff_1425350_3181300# GND efet w=12325 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1416 diff_2169200_3327750# diff_2148900_3310350# GND GND efet w=27550 l=14500
+ ad=1.36662e+08 pd=66700 as=0 ps=0 
M1417 diff_1425350_3181300# diff_2166300_3074000# diff_2169200_3327750# GND efet w=26100 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1418 diff_1425350_3181300# diff_1425350_3181300# diff_1950250_3256700# GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.046e+07 ps=29000 
M1419 diff_1425350_3181300# diff_1425350_3181300# GND GND efet w=59450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1420 diff_1425350_3181300# diff_1425350_3181300# diff_1764650_3221900# GND efet w=21025 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1421 diff_1808150_3240750# diff_1425350_3181300# diff_1425350_3181300# GND efet w=24650 l=11600
+ ad=1.682e+08 pd=66700 as=0 ps=0 
M1422 GND diff_1815400_3242200# diff_1808150_3240750# GND efet w=26825 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1423 diff_1899500_3262500# diff_1879200_3292950# GND GND efet w=23925 l=15225
+ ad=1.72405e+08 pd=69600 as=0 ps=0 
M1424 diff_1425350_3181300# diff_1425350_3181300# diff_1899500_3262500# GND efet w=28275 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1425 diff_1943000_3256700# diff_1425350_3181300# diff_1425350_3181300# GND efet w=29000 l=11600
+ ad=1.78712e+08 pd=75400 as=0 ps=0 
M1426 GND diff_1950250_3256700# diff_1943000_3256700# GND efet w=25375 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1427 diff_2014050_3292950# diff_1425350_3181300# diff_1425350_3181300# GND efet w=5800 l=11600
+ ad=4.41525e+07 pd=29000 as=0 ps=0 
M1428 diff_1425350_3181300# diff_2106850_3184200# diff_2086550_3310350# GND efet w=5800 l=12325
+ ad=0 pd=0 as=4.205e+07 ps=26100 
M1429 diff_2148900_3310350# diff_1425350_3181300# diff_1425350_3181300# GND efet w=3625 l=16675
+ ad=4.205e+07 pd=26100 as=0 ps=0 
M1430 diff_1425350_3181300# diff_2106850_3184200# diff_2086550_3255250# GND efet w=6525 l=13775
+ ad=0 pd=0 as=4.6255e+07 ps=29000 
M1431 diff_2148900_3292950# diff_1425350_3181300# diff_1425350_3181300# GND efet w=3625 l=18125
+ ad=4.41525e+07 pd=29000 as=0 ps=0 
M1432 diff_2034350_3262500# diff_2014050_3292950# GND GND efet w=24650 l=13050
+ ad=1.5979e+08 pd=66700 as=0 ps=0 
M1433 diff_1425350_3181300# diff_2025650_3074000# diff_2034350_3262500# GND efet w=26825 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1434 diff_2077850_3256700# diff_1425350_3181300# diff_1425350_3181300# GND efet w=26100 l=14500
+ ad=1.5979e+08 pd=69600 as=0 ps=0 
M1435 diff_1899500_3221900# diff_1879200_3203050# GND GND efet w=23200 l=13775
+ ad=1.682e+08 pd=66700 as=0 ps=0 
M1436 diff_1425350_3181300# diff_1687800_3075450# diff_1680550_3242200# GND efet w=6525 l=13775
+ ad=0 pd=0 as=5.67675e+07 ps=37700 
M1437 diff_1742900_3204500# diff_1718250_3075450# diff_1425350_3181300# GND efet w=4350 l=12325
+ ad=3.7845e+07 pd=26100 as=0 ps=0 
M1438 diff_1425350_3181300# diff_1687800_3075450# diff_1680550_3149400# GND efet w=7250 l=11600
+ ad=0 pd=0 as=4.6255e+07 ps=31900 
M1439 diff_1742900_3185650# diff_1718250_3075450# diff_1425350_3181300# GND efet w=5800 l=11600
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M1440 diff_1673300_3150850# diff_1425350_3181300# diff_1425350_3181300# GND efet w=24650 l=13775
+ ad=1.61892e+08 pd=63800 as=0 ps=0 
M1441 GND diff_1680550_3149400# diff_1673300_3150850# GND efet w=23200 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1442 diff_1425350_3181300# diff_1829900_3075450# diff_1815400_3242200# GND efet w=7250 l=11600
+ ad=0 pd=0 as=6.09725e+07 ps=31900 
M1443 diff_1425350_3181300# diff_1425350_3181300# diff_1899500_3221900# GND efet w=26825 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1444 diff_1943000_3239300# diff_1425350_3181300# diff_1425350_3181300# GND efet w=24650 l=14500
+ ad=1.53482e+08 pd=69600 as=0 ps=0 
M1445 GND diff_1951700_3203050# diff_1943000_3239300# GND efet w=26100 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1446 GND diff_2086550_3255250# diff_2077850_3256700# GND efet w=21025 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1447 diff_2034350_3220450# diff_2014050_3203050# GND GND efet w=24650 l=14500
+ ad=1.63995e+08 pd=66700 as=0 ps=0 
M1448 diff_1879200_3203050# diff_1858900_3075450# diff_1425350_3181300# GND efet w=6525 l=13775
+ ad=4.41525e+07 pd=29000 as=0 ps=0 
M1449 diff_1425350_3181300# diff_1829900_3075450# diff_1816850_3147950# GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.046e+07 ps=29000 
M1450 GND GND diff_606100_2879700# GND efet w=5800 l=30450
+ ad=0 pd=0 as=0 ps=0 
M1451 GND diff_1329650_2830400# diff_1326750_3091400# GND efet w=13050 l=13050
+ ad=0 pd=0 as=5.5506e+08 ps=179800 
M1452 diff_1326750_3091400# GND GND GND efet w=8700 l=65250
+ ad=0 pd=0 as=0 ps=0 
M1453 diff_1329650_2830400# diff_1326750_3091400# GND GND efet w=11600 l=11600
+ ad=1.35191e+09 pd=353800 as=0 ps=0 
M1454 diff_1764650_3155200# diff_1742900_3185650# GND GND efet w=23925 l=13775
+ ad=1.7661e+08 pd=69600 as=0 ps=0 
M1455 diff_1425350_3181300# diff_1425350_3181300# diff_1764650_3155200# GND efet w=24650 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1456 diff_1808150_3149400# diff_1425350_3181300# diff_1425350_3181300# GND efet w=26100 l=14500
+ ad=1.8502e+08 pd=69600 as=0 ps=0 
M1457 GND diff_1816850_3147950# diff_1808150_3149400# GND efet w=27550 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1458 diff_1879200_3185650# diff_1858900_3075450# diff_1425350_3181300# GND efet w=5800 l=11600
+ ad=4.41525e+07 pd=29000 as=0 ps=0 
M1459 diff_1425350_3181300# diff_2025650_3074000# diff_2034350_3220450# GND efet w=26100 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1460 diff_2077850_3240750# diff_1425350_3181300# diff_1425350_3181300# GND efet w=27550 l=17400
+ ad=1.55585e+08 pd=66700 as=0 ps=0 
M1461 GND diff_2085100_3242200# diff_2077850_3240750# GND efet w=22475 l=17400
+ ad=0 pd=0 as=0 ps=0 
M1462 diff_2169200_3262500# diff_2148900_3292950# GND GND efet w=29725 l=15225
+ ad=1.2615e+08 pd=69600 as=0 ps=0 
M1463 diff_1425350_3181300# diff_2166300_3074000# diff_2169200_3262500# GND efet w=27550 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1464 GND diff_2072050_2521550# diff_1425350_3181300# GND efet w=14500 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1465 GND GND diff_1425350_3181300# GND efet w=8700 l=34075
+ ad=0 pd=0 as=0 ps=0 
M1466 GND GND diff_1425350_3181300# GND efet w=7975 l=32625
+ ad=0 pd=0 as=0 ps=0 
M1467 GND diff_2072050_2521550# diff_1425350_3181300# GND efet w=11600 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1468 diff_2169200_3220450# diff_2148900_3203050# GND GND efet w=29000 l=13050
+ ad=1.57688e+08 pd=75400 as=0 ps=0 
M1469 diff_1425350_3181300# diff_2166300_3074000# diff_2169200_3220450# GND efet w=29000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1470 diff_1425350_3181300# diff_1425350_3181300# diff_1951700_3203050# GND efet w=5800 l=11600
+ ad=0 pd=0 as=4.83575e+07 ps=29000 
M1471 diff_2014050_3203050# diff_1425350_3181300# diff_1425350_3181300# GND efet w=5075 l=14500
+ ad=4.205e+07 pd=26100 as=0 ps=0 
M1472 diff_1425350_3181300# diff_1425350_3181300# diff_1951700_3147950# GND efet w=5800 l=11600
+ ad=0 pd=0 as=4.83575e+07 ps=29000 
M1473 diff_1899500_3155200# diff_1879200_3185650# GND GND efet w=23925 l=13775
+ ad=1.78712e+08 pd=69600 as=0 ps=0 
M1474 diff_1425350_3181300# diff_1425350_3181300# diff_1899500_3155200# GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1475 diff_1943000_3149400# diff_1425350_3181300# diff_1425350_3181300# GND efet w=27550 l=11600
+ ad=1.7661e+08 pd=72500 as=0 ps=0 
M1476 GND diff_1951700_3147950# diff_1943000_3149400# GND efet w=25375 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1477 diff_2014050_3185650# diff_1425350_3181300# diff_1425350_3181300# GND efet w=5800 l=11600
+ ad=4.41525e+07 pd=29000 as=0 ps=0 
M1478 diff_2034350_3163900# diff_2014050_3185650# GND GND efet w=26825 l=14500
+ ad=1.47175e+08 pd=69600 as=0 ps=0 
M1479 diff_1425350_3181300# diff_2106850_3184200# diff_2085100_3242200# GND efet w=5800 l=11600
+ ad=0 pd=0 as=4.41525e+07 ps=29000 
M1480 GND diff_2072050_2521550# diff_1425350_3181300# GND efet w=11600 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1481 diff_2148900_3203050# diff_1425350_3181300# diff_1425350_3181300# GND efet w=3625 l=15225
+ ad=4.205e+07 pd=26100 as=0 ps=0 
M1482 diff_1425350_3181300# diff_2106850_3184200# diff_2086550_3147950# GND efet w=5800 l=13050
+ ad=0 pd=0 as=4.83575e+07 ps=31900 
M1483 diff_2148900_3184200# diff_1425350_3181300# diff_1425350_3181300# GND efet w=4350 l=17400
+ ad=5.25625e+07 pd=31900 as=0 ps=0 
M1484 diff_1425350_3181300# diff_2025650_3074000# diff_2034350_3163900# GND efet w=26100 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1485 diff_2079300_3149400# diff_1425350_3181300# diff_1425350_3181300# GND efet w=26100 l=13050
+ ad=1.5979e+08 pd=69600 as=0 ps=0 
M1486 GND diff_2086550_3147950# diff_2079300_3149400# GND efet w=27550 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1487 GND GND diff_1425350_3181300# GND efet w=8700 l=34075
+ ad=0 pd=0 as=0 ps=0 
M1488 GND GND GND GND efet w=118175 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1489 GND GND GND GND efet w=108025 l=18125
+ ad=0 pd=0 as=0 ps=0 
M1490 GND GND diff_1425350_3181300# GND efet w=8700 l=34075
+ ad=0 pd=0 as=0 ps=0 
M1491 diff_2169200_3155200# diff_2148900_3184200# GND GND efet w=26100 l=15950
+ ad=1.38765e+08 pd=63800 as=0 ps=0 
M1492 diff_1425350_3181300# diff_2166300_3074000# diff_2169200_3155200# GND efet w=26825 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1493 GND diff_2072050_2521550# diff_1425350_3181300# GND efet w=11600 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1494 GND GND diff_606100_2879700# GND efet w=5800 l=29000
+ ad=0 pd=0 as=0 ps=0 
M1495 GND GND diff_1329650_2830400# GND efet w=5800 l=65250
+ ad=0 pd=0 as=0 ps=0 
M1496 diff_1136800_2630300# GND GND GND efet w=8700 l=66700
+ ad=1.71144e+09 pd=490100 as=0 ps=0 
M1497 GND diff_1329650_2830400# diff_1136800_2630300# GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1498 diff_1415200_3075450# diff_1326750_3091400# GND GND efet w=14500 l=11600
+ ad=5.31933e+08 pd=162400 as=0 ps=0 
M1499 GND diff_1629800_3060950# diff_1425350_3181300# GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1500 GND diff_1629800_3060950# diff_1687800_3075450# GND efet w=11600 l=11600
+ ad=0 pd=0 as=1.8502e+08 ps=55100 
M1501 GND diff_1711000_3092850# diff_1718250_3075450# GND efet w=11600 l=11600
+ ad=0 pd=0 as=1.8502e+08 ps=55100 
M1502 GND diff_1711000_3092850# diff_1425350_3181300# GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1503 GND GND diff_1415200_3075450# GND efet w=9425 l=65975
+ ad=0 pd=0 as=0 ps=0 
M1504 GND diff_1048350_2488200# diff_622050_2844900# GND efet w=9425 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1505 diff_1629800_3060950# GND GND GND efet w=6525 l=61625
+ ad=6.85415e+08 pd=223300 as=0 ps=0 
M1506 diff_1425350_3181300# diff_1613850_2840550# diff_1613850_2840550# GND efet w=15950 l=11600
+ ad=0 pd=0 as=1.39107e+09 ps=3.7903e+06 
M1507 diff_1687800_3075450# diff_1613850_2840550# diff_1687800_3033400# GND efet w=13775 l=13050
+ ad=0 pd=0 as=-2.02803e+09 ps=1.3456e+06 
M1508 diff_1718250_3075450# diff_1613850_2840550# diff_1687800_3033400# GND efet w=12325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1509 diff_1425350_3181300# diff_1613850_2840550# diff_1613850_2840550# GND efet w=15950 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1510 diff_1135350_3008750# diff_1113600_2989900# GND GND efet w=22475 l=18125
+ ad=1.63995e+08 pd=63800 as=0 ps=0 
M1511 diff_1136800_2630300# diff_1270200_2518650# diff_1336900_3020350# GND efet w=8700 l=10150
+ ad=0 pd=0 as=6.93825e+07 ps=34800 
M1512 diff_1415200_3075450# diff_1270200_2518650# diff_1390550_2979750# GND efet w=8700 l=13050
+ ad=0 pd=0 as=7.569e+07 ps=34800 
M1513 diff_978750_2989900# diff_943950_2878250# diff_655400_2966700# GND efet w=6525 l=12325
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M1514 diff_627850_2752100# diff_914950_2865200# diff_916400_2936250# GND efet w=5800 l=11600
+ ad=0 pd=0 as=5.046e+07 ps=29000 
M1515 diff_907700_2937700# diff_887400_2863750# diff_622050_2844900# GND efet w=27550 l=13050
+ ad=1.682e+08 pd=66700 as=0 ps=0 
M1516 GND GND diff_488650_2876800# GND efet w=7250 l=65250
+ ad=0 pd=0 as=0 ps=0 
M1517 GND diff_136300_2602750# diff_423400_2781100# GND efet w=24650 l=11600
+ ad=0 pd=0 as=6.9803e+08 ps=165300 
M1518 diff_488650_2876800# GND diff_477050_2855050# GND efet w=13050 l=14500
+ ad=0 pd=0 as=8.41e+07 ps=49300 
M1519 GND GND GND GND efet w=401650 l=27550
+ ad=0 pd=0 as=0 ps=0 
M1520 GND GND GND GND efet w=563325 l=55100
+ ad=0 pd=0 as=0 ps=0 
M1521 diff_423400_2781100# diff_258100_694550# GND GND efet w=26825 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1522 GND GND GND GND efet w=29725 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1523 GND GND diff_727900_2842000# GND efet w=5800 l=27550
+ ad=0 pd=0 as=5.90802e+08 ps=191400 
M1524 GND diff_258100_549550# diff_387150_2801400# GND efet w=13050 l=12325
+ ad=0 pd=0 as=7.1485e+08 ps=200100 
M1525 diff_490100_2813000# diff_477050_2855050# GND GND efet w=20300 l=11600
+ ad=5.52958e+08 pd=121800 as=0 ps=0 
M1526 diff_622050_2844900# GND GND GND efet w=7250 l=27550
+ ad=0 pd=0 as=0 ps=0 
M1527 GND diff_536500_2711500# diff_622050_2844900# GND efet w=29000 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1528 GND GND diff_490100_2813000# GND efet w=6525 l=51475
+ ad=0 pd=0 as=0 ps=0 
M1529 diff_387150_2801400# GND GND GND efet w=6525 l=67425
+ ad=0 pd=0 as=0 ps=0 
M1530 diff_477050_2791250# GND diff_490100_2813000# GND efet w=8700 l=11600
+ ad=2.14455e+08 pd=78300 as=0 ps=0 
M1531 GND GND diff_622050_2844900# GND efet w=33350 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1532 GND diff_916400_2936250# diff_907700_2937700# GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1533 diff_978750_2972500# diff_943950_2878250# diff_627850_2752100# GND efet w=5800 l=11600
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M1534 diff_622050_2844900# diff_622050_2844900# diff_1135350_3008750# GND efet w=19575 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1535 diff_655400_2966700# diff_606100_2879700# diff_1051250_3029050# GND efet w=6525 l=10875
+ ad=0 pd=0 as=5.67675e+07 ps=34800 
M1536 diff_1113600_2989900# diff_622050_2844900# diff_655400_2966700# GND efet w=5800 l=10150
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M1537 diff_627850_2752100# diff_606100_2879700# diff_1051250_2936250# GND efet w=5800 l=10150
+ ad=0 pd=0 as=5.046e+07 ps=29000 
M1538 diff_1113600_2972500# diff_622050_2844900# diff_627850_2752100# GND efet w=5800 l=10150
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M1539 diff_999050_2946400# diff_978750_2972500# GND GND efet w=26100 l=13050
+ ad=1.8502e+08 pd=75400 as=0 ps=0 
M1540 diff_622050_2844900# diff_622050_2844900# diff_999050_2946400# GND efet w=23200 l=17400
+ ad=0 pd=0 as=0 ps=0 
M1541 diff_1044000_2936250# diff_1032400_2863750# diff_622050_2844900# GND efet w=25375 l=12325
+ ad=1.72405e+08 pd=72500 as=0 ps=0 
M1542 diff_784450_2863750# GND GND GND efet w=7975 l=31175
+ ad=8.72537e+08 pd=182700 as=0 ps=0 
M1543 GND diff_1051250_2936250# diff_1044000_2936250# GND efet w=25375 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1544 diff_1135350_2940600# diff_1113600_2972500# GND GND efet w=23925 l=15225
+ ad=1.74508e+08 pd=66700 as=0 ps=0 
M1545 diff_622050_2844900# diff_622050_2844900# diff_1135350_2940600# GND efet w=21025 l=19575
+ ad=0 pd=0 as=0 ps=0 
M1546 GND diff_1048350_2488200# diff_622050_2844900# GND efet w=8700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1547 diff_1355750_2985550# diff_1329650_2830400# diff_1326750_3091400# GND efet w=21750 l=12325
+ ad=2.24968e+08 pd=81200 as=0 ps=0 
M1548 GND GND diff_655400_2966700# GND efet w=6525 l=32625
+ ad=0 pd=0 as=0 ps=0 
M1549 GND diff_1336900_3020350# diff_1355750_2985550# GND efet w=34075 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1550 diff_1402150_2984100# diff_1390550_2979750# GND GND efet w=34800 l=11600
+ ad=2.29172e+08 pd=84100 as=0 ps=0 
M1551 diff_1329650_2830400# diff_1329650_2830400# diff_1402150_2984100# GND efet w=13050 l=18850
+ ad=0 pd=0 as=0 ps=0 
M1552 GND GND diff_627850_2752100# GND efet w=6525 l=31175
+ ad=0 pd=0 as=0 ps=0 
M1553 GND diff_1782050_3013100# diff_1425350_3181300# GND efet w=14500 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1554 GND diff_1782050_3013100# diff_1829900_3075450# GND efet w=11600 l=10150
+ ad=0 pd=0 as=1.8502e+08 ps=55100 
M1555 GND diff_1425350_3181300# diff_1858900_3075450# GND efet w=13050 l=10150
+ ad=0 pd=0 as=2.08148e+08 ps=58000 
M1556 GND diff_1425350_3181300# diff_1425350_3181300# GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1557 GND diff_1425350_3181300# diff_1425350_3181300# GND efet w=10150 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1558 diff_1425350_3181300# diff_1613850_2840550# diff_1613850_2840550# GND efet w=13775 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1559 diff_1829900_3075450# diff_1613850_2840550# diff_1687800_3033400# GND efet w=12325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1560 diff_1858900_3075450# diff_1613850_2840550# diff_1687800_3033400# GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1561 diff_1425350_3181300# diff_1613850_2840550# diff_1613850_2840550# GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1562 GND diff_1613850_2840550# diff_1629800_3060950# GND efet w=11600 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1563 diff_1711000_3092850# diff_1613850_2840550# GND GND efet w=10150 l=11600
+ ad=4.26807e+08 pd=121800 as=0 ps=0 
M1564 GND diff_1613850_2840550# diff_1782050_3013100# GND efet w=10875 l=12325
+ ad=0 pd=0 as=4.41525e+08 ps=121800 
M1565 diff_1425350_3181300# diff_1613850_2840550# GND GND efet w=10150 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1566 GND diff_1425350_3181300# diff_1425350_3181300# GND efet w=7975 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1567 GND diff_1425350_3181300# diff_1425350_3181300# GND efet w=10875 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1568 GND diff_1425350_3181300# diff_2025650_3074000# GND efet w=13050 l=12325
+ ad=0 pd=0 as=2.08148e+08 ps=58000 
M1569 diff_1425350_3181300# diff_1893700_2785450# diff_1613850_2840550# GND efet w=14500 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1570 diff_1687800_3033400# diff_1893700_2785450# diff_1425350_3181300# GND efet w=12325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1571 diff_1425350_3181300# diff_1947350_2814450# diff_1687800_3033400# GND efet w=12325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1572 diff_2025650_3074000# diff_1947350_2814450# diff_1613850_2840550# GND efet w=13050 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1573 GND diff_1893700_2785450# diff_1425350_3181300# GND efet w=12325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1574 GND diff_1552950_2965250# GND GND efet w=77575 l=6525
+ ad=0 pd=0 as=0 ps=0 
M1575 GND diff_1552950_2965250# GND GND efet w=10150 l=23200
+ ad=0 pd=0 as=0 ps=0 
M1576 diff_1552950_2965250# GND GND GND efet w=6525 l=13775
+ ad=3.364e+07 pd=23200 as=0 ps=0 
M1577 GND diff_1048350_2488200# diff_622050_2844900# GND efet w=10150 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1578 diff_1329650_2830400# GND GND GND efet w=6525 l=71775
+ ad=0 pd=0 as=0 ps=0 
M1579 GND diff_1270200_2518650# diff_1329650_2830400# GND efet w=11600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1580 diff_1270200_2518650# diff_1329650_2830400# GND GND efet w=13050 l=11600
+ ad=1.38555e+09 pd=356700 as=0 ps=0 
M1581 diff_1711000_3092850# GND GND GND efet w=6525 l=45675
+ ad=0 pd=0 as=0 ps=0 
M1582 GND GND diff_1782050_3013100# GND efet w=6525 l=52925
+ ad=0 pd=0 as=0 ps=0 
M1583 diff_1425350_3181300# diff_1947350_2814450# GND GND efet w=11600 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1584 GND diff_1425350_3181300# diff_1425350_3181300# GND efet w=10150 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1585 GND diff_1425350_3181300# diff_2106850_3184200# GND efet w=11600 l=11600
+ ad=0 pd=0 as=1.8502e+08 ps=55100 
M1586 GND diff_2134400_3091400# diff_1425350_3181300# GND efet w=11600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1587 GND diff_2134400_3091400# diff_2166300_3074000# GND efet w=14500 l=11600
+ ad=0 pd=0 as=2.24968e+08 ps=63800 
M1588 diff_1425350_3181300# diff_2002450_2731800# diff_1613850_2840550# GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1589 diff_2106850_3184200# diff_2002450_2731800# diff_1687800_3033400# GND efet w=12325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1590 diff_1425350_3181300# diff_1613850_2840550# diff_1687800_3033400# GND efet w=12325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1591 diff_2166300_3074000# diff_1613850_2840550# diff_1613850_2840550# GND efet w=10150 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1592 diff_1425350_3181300# GND GND GND efet w=5800 l=47850
+ ad=0 pd=0 as=0 ps=0 
M1593 GND GND diff_1425350_3181300# GND efet w=6525 l=52925
+ ad=0 pd=0 as=0 ps=0 
M1594 GND diff_2002450_2731800# diff_1425350_3181300# GND efet w=10150 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1595 diff_2134400_3091400# diff_1613850_2840550# GND GND efet w=10150 l=13050
+ ad=3.93167e+08 pd=116000 as=0 ps=0 
M1596 GND GND GND GND efet w=13050 l=45675
+ ad=0 pd=0 as=0 ps=0 
M1597 diff_1425350_3181300# GND GND GND efet w=6525 l=48575
+ ad=0 pd=0 as=0 ps=0 
M1598 GND GND diff_1425350_3181300# GND efet w=5800 l=47850
+ ad=0 pd=0 as=0 ps=0 
M1599 diff_2134400_3091400# GND GND GND efet w=5800 l=47850
+ ad=0 pd=0 as=0 ps=0 
M1600 diff_1613850_2840550# diff_1613850_2840550# GND GND efet w=22475 l=18125
+ ad=0 pd=0 as=0 ps=0 
M1601 GND GND diff_1613850_2840550# GND efet w=7250 l=29000
+ ad=0 pd=0 as=0 ps=0 
M1602 GND GND diff_1270200_2518650# GND efet w=6525 l=68875
+ ad=0 pd=0 as=0 ps=0 
M1603 diff_1136800_2604200# GND GND GND efet w=9425 l=73950
+ ad=1.66518e+09 pd=484300 as=0 ps=0 
M1604 GND diff_1270200_2518650# diff_1136800_2604200# GND efet w=13775 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1605 diff_1415200_2920300# diff_1329650_2830400# GND GND efet w=13050 l=11600
+ ad=5.23522e+08 pd=159500 as=0 ps=0 
M1606 GND GND diff_1415200_2920300# GND efet w=8700 l=66700
+ ad=0 pd=0 as=0 ps=0 
M1607 diff_1552950_2940600# GND GND GND efet w=6525 l=13775
+ ad=3.99475e+07 pd=31900 as=0 ps=0 
M1608 diff_1425350_3181300# diff_1552950_2940600# diff_1425350_3181300# GND efet w=57275 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1609 diff_1425350_3181300# diff_1552950_2940600# GND GND efet w=7250 l=21750
+ ad=0 pd=0 as=0 ps=0 
M1610 diff_727900_2842000# GND GND GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1611 GND diff_501700_2402650# diff_784450_2863750# GND efet w=29000 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1612 GND diff_536500_2711500# diff_727900_2842000# GND efet w=27550 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1613 diff_784450_2863750# diff_536500_2711500# GND GND efet w=29725 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1614 GND diff_867100_2815900# diff_887400_2863750# GND efet w=15950 l=10150
+ ad=0 pd=0 as=2.54402e+08 ps=63800 
M1615 GND diff_867100_2815900# diff_914950_2865200# GND efet w=11600 l=10150
+ ad=0 pd=0 as=1.82918e+08 ps=55100 
M1616 GND diff_938150_2881150# diff_943950_2878250# GND efet w=11600 l=11600
+ ad=0 pd=0 as=1.87122e+08 ps=58000 
M1617 GND diff_938150_2881150# diff_622050_2844900# GND efet w=15950 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1618 diff_887400_2863750# diff_880150_2855050# diff_772850_2547650# GND efet w=15950 l=11600
+ ad=0 pd=0 as=-1.06973e+09 ps=896100 
M1619 diff_914950_2865200# diff_880150_2855050# diff_839550_2504150# GND efet w=10150 l=11600
+ ad=0 pd=0 as=-1.25685e+09 ps=626400 
M1620 diff_943950_2878250# diff_938150_2853600# diff_839550_2504150# GND efet w=12325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1621 diff_622050_2844900# diff_938150_2853600# diff_772850_2547650# GND efet w=15950 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1622 GND GND GND GND efet w=9425 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1623 diff_387150_2801400# diff_417600_2791250# diff_423400_2781100# GND efet w=23200 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1624 GND diff_606100_2879700# diff_1032400_2863750# GND efet w=15950 l=10150
+ ad=0 pd=0 as=2.54402e+08 ps=63800 
M1625 diff_606100_2879700# diff_606100_2879700# GND GND efet w=9425 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1626 GND diff_622050_2844900# diff_622050_2844900# GND efet w=7975 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1627 diff_622050_2844900# diff_622050_2844900# GND GND efet w=15225 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1628 diff_1136800_2604200# GND diff_1336900_2865200# GND efet w=7250 l=11600
+ ad=0 pd=0 as=5.4665e+07 ps=31900 
M1629 diff_1613850_2840550# diff_1613850_2840550# GND GND efet w=14500 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1630 diff_1613850_2840550# diff_1613850_2840550# GND GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1631 diff_1613850_2840550# diff_1613850_2840550# GND GND efet w=13775 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1632 diff_1893700_2785450# GND GND GND efet w=13775 l=13775
+ ad=1.3477e+09 pd=371200 as=0 ps=0 
M1633 GND GND diff_1613850_2840550# GND efet w=29000 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1634 diff_1947350_2814450# GND GND GND efet w=15225 l=12325
+ ad=1.28042e+09 pd=365400 as=0 ps=0 
M1635 diff_2002450_2731800# GND GND GND efet w=13775 l=13775
+ ad=1.53062e+09 pd=437900 as=0 ps=0 
M1636 diff_1613850_2840550# GND GND GND efet w=16675 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1637 GND diff_2215600_2913050# GND GND efet w=52925 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1638 diff_1613850_2840550# diff_1668950_2924650# GND GND efet w=27550 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1639 diff_1613850_2840550# diff_1668950_2924650# GND GND efet w=14500 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1640 GND diff_1668950_2924650# diff_1893700_2785450# GND efet w=13775 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1641 GND diff_1668950_2924650# diff_1947350_2814450# GND efet w=13775 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1642 diff_1613850_2840550# diff_1789300_2900000# GND GND efet w=13775 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1643 GND diff_1613850_2840550# diff_1613850_2840550# GND efet w=24650 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1644 diff_1613850_2840550# diff_1789300_2900000# GND GND efet w=13775 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1645 diff_1415200_2920300# GND diff_1390550_2837650# GND efet w=7250 l=13050
+ ad=0 pd=0 as=5.4665e+07 ps=31900 
M1646 diff_2002450_2731800# diff_1789300_2900000# GND GND efet w=13050 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1647 diff_1613850_2840550# diff_1789300_2900000# GND GND efet w=15950 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1648 GND GND diff_1668950_2924650# GND efet w=5075 l=42775
+ ad=0 pd=0 as=5.73983e+08 ps=165300 
M1649 diff_1613850_2840550# diff_1613850_2840550# GND GND efet w=13050 l=17400
+ ad=0 pd=0 as=0 ps=0 
M1650 diff_1032400_2863750# diff_1004850_2637550# diff_772850_2547650# GND efet w=15950 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1651 diff_606100_2879700# diff_1004850_2637550# diff_839550_2504150# GND efet w=10875 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1652 diff_622050_2844900# diff_772850_2547650# diff_839550_2504150# GND efet w=11600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1653 diff_622050_2844900# diff_772850_2547650# diff_772850_2547650# GND efet w=15950 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1654 GND diff_1336900_2865200# diff_1355750_2828950# GND efet w=40600 l=11600
+ ad=0 pd=0 as=2.29172e+08 ps=89900 
M1655 GND diff_880150_2855050# diff_867100_2815900# GND efet w=12325 l=12325
+ ad=0 pd=0 as=5.02498e+08 ps=145000 
M1656 diff_938150_2881150# diff_938150_2853600# GND GND efet w=11600 l=11600
+ ad=2.81735e+08 pd=75400 as=0 ps=0 
M1657 diff_1355750_2828950# diff_1270200_2518650# diff_1329650_2830400# GND efet w=21750 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1658 diff_1402150_2830400# diff_1390550_2837650# GND GND efet w=38425 l=12325
+ ad=2.2707e+08 pd=87000 as=0 ps=0 
M1659 GND diff_1613850_2840550# diff_1893700_2785450# GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1660 GND diff_1613850_2840550# diff_2002450_2731800# GND efet w=13050 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1661 diff_1668950_2924650# diff_1789300_2900000# GND GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1662 diff_1789300_2900000# diff_1983600_2676700# GND GND efet w=52200 l=13050
+ ad=6.62287e+08 pd=182700 as=0 ps=0 
M1663 diff_1270200_2518650# diff_1270200_2518650# diff_1402150_2830400# GND efet w=11600 l=21025
+ ad=0 pd=0 as=0 ps=0 
M1664 diff_1613850_2840550# GND diff_1613850_2840550# GND efet w=41325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1665 diff_1613850_2840550# GND GND GND efet w=8700 l=40600
+ ad=0 pd=0 as=0 ps=0 
M1666 GND GND diff_1613850_2840550# GND efet w=19575 l=21025
+ ad=0 pd=0 as=0 ps=0 
M1667 GND GND diff_622050_2844900# GND efet w=5800 l=60900
+ ad=0 pd=0 as=0 ps=0 
M1668 GND diff_1004850_2637550# diff_606100_2879700# GND efet w=11600 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1669 diff_622050_2844900# diff_772850_2547650# GND GND efet w=11600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1670 diff_417600_2791250# diff_477050_2791250# GND GND efet w=19575 l=12325
+ ad=3.23785e+08 pd=92800 as=0 ps=0 
M1671 GND GND diff_417600_2791250# GND efet w=8700 l=65250
+ ad=0 pd=0 as=0 ps=0 
M1672 GND diff_387150_2801400# GND GND efet w=13775 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1673 GND diff_703250_2691200# diff_606100_2879700# GND efet w=43500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1674 diff_627850_2752100# GND GND GND efet w=7975 l=23200
+ ad=0 pd=0 as=0 ps=0 
M1675 diff_536500_2711500# GND GND GND efet w=26100 l=13050
+ ad=1.89646e+09 pd=490100 as=0 ps=0 
M1676 GND GND GND GND efet w=10150 l=50750
+ ad=0 pd=0 as=0 ps=0 
M1677 GND GND GND GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1678 GND GND diff_536500_2711500# GND efet w=6525 l=29725
+ ad=0 pd=0 as=0 ps=0 
M1679 GND GND GND GND efet w=79750 l=27550
+ ad=0 pd=0 as=0 ps=0 
M1680 diff_320450_2669450# diff_275500_2569400# GND GND efet w=23925 l=15225
+ ad=1.77451e+09 pd=391500 as=0 ps=0 
M1681 GND diff_282750_2514300# diff_320450_2669450# GND efet w=20300 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1682 diff_275500_2569400# diff_250850_2582450# diff_275500_2569400# GND efet w=57275 l=14500
+ ad=7.35875e+08 pd=310300 as=0 ps=0 
M1683 diff_250850_2582450# GND GND GND efet w=7250 l=11600
+ ad=5.25625e+07 pd=29000 as=0 ps=0 
M1684 GND diff_282750_2514300# diff_275500_2569400# GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1685 diff_468350_2653500# GND GND GND efet w=7975 l=60900
+ ad=7.2326e+08 pd=197200 as=0 ps=0 
M1686 GND GND diff_468350_2653500# GND efet w=15950 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1687 diff_629300_2881150# GND GND GND efet w=7975 l=26825
+ ad=6.09725e+08 pd=168200 as=0 ps=0 
M1688 diff_606100_2879700# GND GND GND efet w=8700 l=21750
+ ad=0 pd=0 as=0 ps=0 
M1689 diff_629300_2881150# GND GND GND efet w=50750 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1690 GND diff_749650_2701350# diff_629300_2881150# GND efet w=42775 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1691 diff_627850_2752100# GND GND GND efet w=53650 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1692 GND diff_794600_2701350# diff_627850_2752100# GND efet w=50025 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1693 GND GND diff_867100_2815900# GND efet w=5800 l=62350
+ ad=0 pd=0 as=0 ps=0 
M1694 GND GND diff_938150_2881150# GND efet w=6525 l=50025
+ ad=0 pd=0 as=0 ps=0 
M1695 diff_606100_2879700# GND GND GND efet w=5800 l=52200
+ ad=0 pd=0 as=0 ps=0 
M1696 GND GND GND GND efet w=23925 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1697 GND diff_1729850_2853600# diff_1613850_2840550# GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1698 diff_1613850_2840550# diff_1729850_2853600# GND GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1699 diff_1947350_2814450# diff_1729850_2853600# GND GND efet w=14500 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1700 diff_1613850_2840550# diff_1729850_2853600# GND GND efet w=14500 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1701 diff_1613850_2840550# diff_1613850_2840550# GND GND efet w=10150 l=18125
+ ad=0 pd=0 as=0 ps=0 
M1702 diff_1613850_2840550# diff_1613850_2840550# GND GND efet w=11600 l=17400
+ ad=0 pd=0 as=0 ps=0 
M1703 diff_1613850_2840550# diff_1613850_2840550# GND GND efet w=13775 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1704 diff_1893700_2785450# diff_1613850_2840550# GND GND efet w=16675 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1705 diff_1947350_2814450# diff_1613850_2840550# GND GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1706 diff_2002450_2731800# diff_1613850_2840550# GND GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1707 diff_1613850_2840550# diff_1613850_2840550# GND GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1708 diff_1613850_2840550# diff_1719700_2741950# diff_1613850_2840550# GND efet w=58725 l=29725
+ ad=0 pd=0 as=0 ps=0 
M1709 GND GND GND GND efet w=8700 l=65250
+ ad=0 pd=0 as=0 ps=0 
M1710 diff_1613850_2840550# diff_1660250_2731800# diff_1613850_2840550# GND efet w=15950 l=50750
+ ad=0 pd=0 as=0 ps=0 
M1711 diff_1004850_2637550# GND GND GND efet w=8700 l=15950
+ ad=1.0891e+09 pd=266800 as=0 ps=0 
M1712 diff_1329650_2769500# GND GND GND efet w=7250 l=65250
+ ad=5.48753e+08 pd=165300 as=0 ps=0 
M1713 GND diff_1329650_2521550# diff_1329650_2769500# GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1714 diff_1200600_2627400# GND GND GND efet w=8700 l=68150
+ ad=1.73666e+09 pd=449500 as=0 ps=0 
M1715 GND diff_1329650_2521550# diff_1200600_2627400# GND efet w=15225 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1716 diff_1329650_2521550# diff_1329650_2769500# GND GND efet w=13050 l=11600
+ ad=1.21945e+09 pd=345100 as=0 ps=0 
M1717 GND GND diff_1329650_2521550# GND efet w=6525 l=67425
+ ad=0 pd=0 as=0 ps=0 
M1718 diff_1415200_2753550# diff_1329650_2769500# GND GND efet w=14500 l=13050
+ ad=5.2142e+08 pd=162400 as=0 ps=0 
M1719 GND GND diff_1415200_2753550# GND efet w=8700 l=66700
+ ad=0 pd=0 as=0 ps=0 
M1720 diff_772850_2547650# GND GND GND efet w=16675 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1721 diff_1200600_2627400# diff_1331100_2717300# diff_1336900_2698450# GND efet w=8700 l=11600
+ ad=0 pd=0 as=6.51775e+07 ps=34800 
M1722 diff_1415200_2753550# diff_1331100_2717300# diff_1390550_2670900# GND efet w=9425 l=12325
+ ad=0 pd=0 as=6.09725e+07 ps=40600 
M1723 diff_468350_2653500# GND diff_703250_2691200# GND efet w=7250 l=13050
+ ad=0 pd=0 as=5.67675e+07 ps=34800 
M1724 diff_749650_2701350# GND diff_423400_2592600# GND efet w=7250 l=11600
+ ad=5.4665e+07 pd=31900 as=5.31933e+08 ps=150800 
M1725 diff_794600_2701350# GND diff_368300_2570850# GND efet w=7975 l=13775
+ ad=5.4665e+07 pd=31900 as=9.12485e+08 ps=237800 
M1726 diff_275500_2569400# diff_250850_2582450# GND GND efet w=7975 l=37700
+ ad=0 pd=0 as=0 ps=0 
M1727 diff_423400_2592600# diff_258100_549550# GND GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1728 GND diff_258100_694550# diff_368300_2570850# GND efet w=15950 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1729 GND GND diff_368300_2570850# GND efet w=9425 l=55825
+ ad=0 pd=0 as=0 ps=0 
M1730 GND GND diff_282750_2514300# GND efet w=6525 l=36975
+ ad=0 pd=0 as=1.07648e+09 ps=435000 
M1731 diff_282750_2514300# GND diff_265350_2463550# GND efet w=48575 l=15225
+ ad=0 pd=0 as=3.25887e+08 ps=104400 
M1732 diff_265350_2463550# diff_230550_2438900# GND GND efet w=44225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1733 GND GND diff_204450_2418600# GND efet w=6525 l=41325
+ ad=0 pd=0 as=8.03155e+08 ps=269700 
M1734 GND GND diff_282750_2514300# GND efet w=17400 l=18125
+ ad=0 pd=0 as=0 ps=0 
M1735 diff_282750_2514300# diff_249400_1373150# GND GND efet w=23200 l=8700
+ ad=0 pd=0 as=0 ps=0 
M1736 GND GND diff_423400_2592600# GND efet w=6525 l=52925
+ ad=0 pd=0 as=0 ps=0 
M1737 diff_230550_2438900# GND diff_204450_2418600# GND efet w=14500 l=11600
+ ad=2.4389e+08 pd=75400 as=0 ps=0 
M1738 GND GND diff_204450_2418600# GND efet w=21025 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1739 diff_606100_2879700# GND GND GND efet w=43500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1740 diff_880150_2855050# GND GND GND efet w=13050 l=10150
+ ad=1.36032e+09 pd=330600 as=0 ps=0 
M1741 diff_938150_2853600# GND GND GND efet w=20300 l=10150
+ ad=1.03864e+09 pd=368300 as=0 ps=0 
M1742 diff_880150_2855050# diff_904800_2683950# GND GND efet w=12325 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1743 diff_938150_2853600# diff_904800_2683950# GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1744 GND diff_1007750_2685400# diff_1004850_2637550# GND efet w=20300 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1745 diff_772850_2547650# diff_1007750_2685400# GND GND efet w=20300 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1746 diff_880150_2855050# diff_884500_2589700# diff_880150_2855050# GND efet w=30450 l=35525
+ ad=0 pd=0 as=0 ps=0 
M1747 GND diff_136300_2602750# diff_204450_2418600# GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1748 GND GND diff_501700_2402650# GND efet w=7250 l=69600
+ ad=0 pd=0 as=1.99317e+09 ps=548100 
M1749 diff_880150_2855050# diff_884500_2589700# GND GND efet w=7250 l=56550
+ ad=0 pd=0 as=0 ps=0 
M1750 diff_938150_2853600# diff_943950_2649150# diff_938150_2853600# GND efet w=60900 l=30450
+ ad=0 pd=0 as=0 ps=0 
M1751 diff_1004850_2637550# diff_999050_2583900# diff_1004850_2637550# GND efet w=29725 l=60175
+ ad=0 pd=0 as=0 ps=0 
M1752 GND diff_1336900_2698450# diff_1355750_2662200# GND efet w=39150 l=11600
+ ad=0 pd=0 as=2.31275e+08 ps=87000 
M1753 diff_772850_2547650# diff_1058500_2582450# diff_772850_2547650# GND efet w=62350 l=31900
+ ad=0 pd=0 as=0 ps=0 
M1754 diff_938150_2853600# diff_943950_2649150# GND GND efet w=7250 l=55100
+ ad=0 pd=0 as=0 ps=0 
M1755 diff_1004850_2637550# diff_999050_2583900# GND GND efet w=7250 l=56550
+ ad=0 pd=0 as=0 ps=0 
M1756 diff_904800_2683950# diff_1007750_2685400# GND GND efet w=24650 l=11600
+ ad=4.07885e+08 pd=113100 as=0 ps=0 
M1757 GND GND diff_904800_2683950# GND efet w=8700 l=66700
+ ad=0 pd=0 as=0 ps=0 
M1758 diff_1355750_2662200# diff_1329650_2521550# diff_1329650_2769500# GND efet w=21750 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1759 diff_1402150_2665100# diff_1390550_2670900# GND GND efet w=39150 l=13050
+ ad=2.24968e+08 pd=81200 as=0 ps=0 
M1760 diff_1329650_2521550# diff_1329650_2521550# diff_1402150_2665100# GND efet w=13050 l=20300
+ ad=0 pd=0 as=0 ps=0 
M1761 diff_1613850_2840550# diff_1660250_2731800# GND GND efet w=10150 l=55825
+ ad=0 pd=0 as=0 ps=0 
M1762 diff_1613850_2840550# diff_1773350_2733250# diff_1613850_2840550# GND efet w=28275 l=31175
+ ad=0 pd=0 as=0 ps=0 
M1763 diff_1613850_2840550# diff_1719700_2741950# GND GND efet w=7975 l=60175
+ ad=0 pd=0 as=0 ps=0 
M1764 diff_1613850_2840550# diff_1773350_2733250# GND GND efet w=7250 l=56550
+ ad=0 pd=0 as=0 ps=0 
M1765 diff_1613850_2840550# diff_1832800_2763700# diff_1613850_2840550# GND efet w=29725 l=55100
+ ad=0 pd=0 as=0 ps=0 
M1766 diff_1893700_2785450# diff_1886450_2740500# diff_1893700_2785450# GND efet w=29725 l=52925
+ ad=0 pd=0 as=0 ps=0 
M1767 diff_1947350_2814450# diff_1945900_2772400# diff_1947350_2814450# GND efet w=29725 l=52925
+ ad=0 pd=0 as=0 ps=0 
M1768 diff_2002450_2731800# diff_2002450_2731800# diff_2002450_2731800# GND efet w=29000 l=32625
+ ad=0 pd=0 as=0 ps=0 
M1769 diff_1613850_2840550# diff_1832800_2763700# GND GND efet w=7250 l=56550
+ ad=0 pd=0 as=0 ps=0 
M1770 diff_1893700_2785450# diff_1886450_2740500# GND GND efet w=8700 l=59450
+ ad=0 pd=0 as=0 ps=0 
M1771 diff_1947350_2814450# diff_1945900_2772400# GND GND efet w=9425 l=54375
+ ad=0 pd=0 as=0 ps=0 
M1772 diff_2002450_2731800# diff_2002450_2731800# GND GND efet w=9425 l=55825
+ ad=0 pd=0 as=0 ps=0 
M1773 GND GND diff_1789300_2900000# GND efet w=5075 l=41325
+ ad=0 pd=0 as=0 ps=0 
M1774 GND GND diff_1613850_2840550# GND efet w=11600 l=42775
+ ad=0 pd=0 as=0 ps=0 
M1775 diff_1613850_2840550# diff_2061900_2756450# diff_1613850_2840550# GND efet w=30450 l=31175
+ ad=0 pd=0 as=0 ps=0 
M1776 diff_1613850_2840550# diff_1729850_2853600# GND GND efet w=26100 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1777 diff_1729850_2853600# diff_1613850_2688300# GND GND efet w=48575 l=10875
+ ad=5.99212e+08 pd=179800 as=0 ps=0 
M1778 GND GND diff_1729850_2853600# GND efet w=10150 l=44225
+ ad=0 pd=0 as=0 ps=0 
M1779 diff_1613850_2840550# diff_2061900_2756450# GND GND efet w=7250 l=53650
+ ad=0 pd=0 as=0 ps=0 
M1780 GND diff_2282300_2737600# diff_1613850_2688300# GND efet w=8700 l=13050
+ ad=0 pd=0 as=1.46965e+09 ps=446600 
M1781 GND diff_2282300_2737600# diff_1983600_2676700# GND efet w=7250 l=13050
+ ad=0 pd=0 as=1.56006e+09 ps=336400 
M1782 diff_1660250_2731800# GND GND GND efet w=8700 l=11600
+ ad=9.04075e+07 pd=43500 as=0 ps=0 
M1783 diff_1719700_2741950# GND GND GND efet w=8700 l=12325
+ ad=7.77925e+07 pd=37700 as=0 ps=0 
M1784 diff_1773350_2733250# GND GND GND efet w=10150 l=10150
+ ad=9.251e+07 pd=40600 as=0 ps=0 
M1785 diff_1832800_2763700# GND GND GND efet w=10150 l=10150
+ ad=9.04075e+07 pd=40600 as=0 ps=0 
M1786 diff_1886450_2740500# GND GND GND efet w=8700 l=10150
+ ad=7.77925e+07 pd=37700 as=0 ps=0 
M1787 diff_1945900_2772400# GND GND GND efet w=9425 l=10875
+ ad=7.569e+07 pd=34800 as=0 ps=0 
M1788 diff_2002450_2731800# GND GND GND efet w=10875 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1789 diff_2061900_2756450# GND GND GND efet w=10150 l=11600
+ ad=8.8305e+07 pd=37700 as=0 ps=0 
M1790 GND GND diff_1629800_2623050# GND efet w=5800 l=68875
+ ad=0 pd=0 as=1.14166e+09 ps=234900 
M1791 GND GND diff_1699400_2604200# GND efet w=6525 l=65975
+ ad=0 pd=0 as=1.25519e+09 ps=287100 
M1792 GND GND diff_1790750_2624500# GND efet w=5800 l=66700
+ ad=0 pd=0 as=3.84758e+08 ps=130500 
M1793 GND GND diff_1919800_2605650# GND efet w=5800 l=63800
+ ad=0 pd=0 as=1.07648e+09 ps=208800 
M1794 diff_1613850_2688300# diff_1668950_2660750# diff_1693600_2615800# GND efet w=8700 l=11600
+ ad=0 pd=0 as=1.02602e+09 ps=234900 
M1795 GND GND diff_1693600_2615800# GND efet w=5800 l=33350
+ ad=0 pd=0 as=0 ps=0 
M1796 GND GND diff_1987950_2604200# GND efet w=5800 l=72500
+ ad=0 pd=0 as=1.30776e+09 ps=292900 
M1797 GND GND diff_2079300_2623050# GND efet w=5800 l=63800
+ ad=0 pd=0 as=3.99475e+08 ps=124700 
M1798 GND GND diff_1982150_2614350# GND efet w=6525 l=41325
+ ad=0 pd=0 as=1.08069e+09 ps=232000 
M1799 diff_1983600_2676700# diff_1668950_2660750# diff_1982150_2614350# GND efet w=10875 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1800 diff_772850_2547650# diff_1058500_2582450# GND GND efet w=7250 l=53650
+ ad=0 pd=0 as=0 ps=0 
M1801 GND diff_249400_1373150# diff_1136800_2630300# GND efet w=8700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1802 diff_1200600_2627400# GND GND GND efet w=8700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1803 diff_1007750_2685400# diff_249400_1373150# diff_1136800_2604200# GND efet w=8700 l=11600
+ ad=1.30355e+08 pd=78300 as=0 ps=0 
M1804 diff_1200600_2607100# GND diff_1007750_2685400# GND efet w=7975 l=13050
+ ad=2.03312e+09 pd=501700 as=0 ps=0 
M1805 diff_688750_2531700# diff_682950_2483850# diff_688750_2531700# GND efet w=73950 l=29000
+ ad=1.92589e+09 pd=623500 as=0 ps=0 
M1806 GND GND diff_774300_2469350# GND efet w=6525 l=60175
+ ad=0 pd=0 as=1.70302e+08 ps=81200 
M1807 diff_884500_2589700# GND GND GND efet w=10150 l=11600
+ ad=8.8305e+07 pd=37700 as=0 ps=0 
M1808 diff_943950_2649150# GND GND GND efet w=11600 l=10150
+ ad=8.62025e+07 pd=37700 as=0 ps=0 
M1809 diff_999050_2583900# GND GND GND efet w=10875 l=10150
+ ad=8.8305e+07 pd=40600 as=0 ps=0 
M1810 diff_1058500_2582450# GND GND GND efet w=11600 l=11600
+ ad=8.19975e+07 pd=40600 as=0 ps=0 
M1811 diff_772850_2547650# diff_688750_2531700# GND GND efet w=41325 l=21025
+ ad=0 pd=0 as=0 ps=0 
M1812 GND GND diff_682950_2483850# GND efet w=7975 l=12325
+ ad=0 pd=0 as=4.83575e+07 ps=31900 
M1813 GND GND diff_595950_2407000# GND efet w=34075 l=13775
+ ad=0 pd=0 as=2.20762e+08 ps=75400 
M1814 GND diff_682950_2483850# diff_688750_2531700# GND efet w=5800 l=43500
+ ad=0 pd=0 as=0 ps=0 
M1815 GND diff_774300_2469350# diff_772850_2547650# GND efet w=29725 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1816 GND GND GND GND efet w=6525 l=68875
+ ad=0 pd=0 as=0 ps=0 
M1817 diff_568400_2407000# GND diff_501700_2402650# GND efet w=30450 l=11600
+ ad=4.85678e+08 pd=92800 as=0 ps=0 
M1818 diff_595950_2407000# diff_552450_2137300# diff_568400_2407000# GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1819 diff_614800_2349000# GND GND GND efet w=32625 l=12325
+ ad=6.728e+08 pd=237800 as=0 ps=0 
M1820 diff_501700_2402650# diff_136300_2602750# GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1821 diff_614800_2349000# GND diff_595950_2349000# GND efet w=36975 l=20300
+ ad=0 pd=0 as=2.1025e+08 ps=72500 
M1822 diff_529250_2347550# GND GND GND efet w=30450 l=13050
+ ad=2.58608e+08 pd=78300 as=0 ps=0 
M1823 diff_549550_2349000# diff_537950_2248950# diff_529250_2347550# GND efet w=29000 l=13050
+ ad=2.1866e+08 pd=75400 as=0 ps=0 
M1824 GND GND diff_549550_2349000# GND efet w=25375 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1825 diff_595950_2349000# diff_552450_2137300# GND GND efet w=29000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1826 diff_633650_2347550# diff_622050_2318550# diff_614800_2349000# GND efet w=30450 l=11600
+ ad=2.20762e+08 pd=75400 as=0 ps=0 
M1827 GND diff_640900_2343200# diff_633650_2347550# GND efet w=31175 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1828 diff_774300_2469350# diff_688750_2531700# GND GND efet w=13050 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1829 GND GND diff_855500_2512850# GND efet w=8700 l=51475
+ ad=0 pd=0 as=2.20762e+08 ps=107300 
M1830 GND diff_855500_2512850# diff_839550_2504150# GND efet w=20300 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1831 GND diff_974400_2502700# diff_855500_2492550# GND efet w=7250 l=40600
+ ad=0 pd=0 as=1.38344e+09 ps=580000 
M1832 GND GND diff_974400_2502700# GND efet w=5800 l=10150
+ ad=0 pd=0 as=5.046e+07 ps=29000 
M1833 diff_1046900_2517200# GND GND GND efet w=5800 l=11600
+ ad=5.67675e+07 pd=34800 as=0 ps=0 
M1834 GND diff_1046900_2517200# diff_1048350_2488200# GND efet w=7975 l=18125
+ ad=0 pd=0 as=-1.383e+09 ps=754000 
M1835 diff_855500_2492550# diff_974400_2502700# diff_855500_2492550# GND efet w=48575 l=23200
+ ad=0 pd=0 as=0 ps=0 
M1836 GND diff_855500_2492550# diff_839550_2504150# GND efet w=21025 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1837 GND diff_855500_2492550# diff_855500_2512850# GND efet w=13775 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1838 diff_1048350_2488200# diff_1046900_2517200# diff_1048350_2488200# GND efet w=81925 l=22475
+ ad=0 pd=0 as=0 ps=0 
M1839 diff_1048350_2488200# diff_1120850_2447600# GND GND efet w=35525 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1840 GND GND diff_1048350_2488200# GND efet w=22475 l=25375
+ ad=0 pd=0 as=0 ps=0 
M1841 GND diff_1158550_2475150# diff_1048350_2488200# GND efet w=34800 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1842 GND GND diff_807650_2418600# GND efet w=5800 l=50750
+ ad=0 pd=0 as=1.78712e+08 ps=92800 
M1843 diff_688750_2531700# GND GND GND efet w=13775 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1844 diff_855500_2492550# diff_935250_2476600# GND GND efet w=13775 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1845 diff_855500_2492550# diff_907700_2450500# diff_894650_2441800# GND efet w=29725 l=10875
+ ad=0 pd=0 as=3.5322e+08 ps=113100 
M1846 diff_688750_2531700# GND GND GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1847 GND diff_784450_2395400# diff_688750_2531700# GND efet w=14500 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1848 diff_688750_2531700# diff_807650_2418600# GND GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1849 diff_894650_2441800# diff_537950_2248950# GND GND efet w=29725 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1850 GND diff_884500_2331600# diff_855500_2492550# GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1851 GND diff_258100_694550# GND GND efet w=18125 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1852 diff_807650_2418600# GND GND GND efet w=14500 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1853 GND diff_537950_1786400# diff_640900_2343200# GND efet w=34075 l=13775
+ ad=0 pd=0 as=1.24678e+09 ps=406000 
M1854 diff_640900_2343200# GND GND GND efet w=26825 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1855 diff_551000_2193850# GND GND GND efet w=32625 l=10150
+ ad=2.64915e+08 pd=78300 as=0 ps=0 
M1856 GND diff_258100_549550# GND GND efet w=12325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1857 diff_569850_2193850# diff_537950_2248950# diff_551000_2193850# GND efet w=31900 l=10150
+ ad=2.54402e+08 pd=81200 as=0 ps=0 
M1858 GND GND diff_569850_2193850# GND efet w=23925 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1859 GND GND GND GND efet w=7975 l=64525
+ ad=0 pd=0 as=0 ps=0 
M1860 diff_633650_2205450# diff_552450_2137300# diff_614800_2167750# GND efet w=36250 l=11600
+ ad=2.88042e+08 pd=92800 as=1.63364e+09 ps=382800 
M1861 GND GND diff_633650_2205450# GND efet w=38425 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1862 diff_680050_2190950# diff_622050_2318550# GND GND efet w=33350 l=11600
+ ad=2.41788e+08 pd=81200 as=0 ps=0 
M1863 diff_614800_2167750# diff_640900_2343200# diff_680050_2190950# GND efet w=33350 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1864 GND diff_249400_1373150# diff_614800_2167750# GND efet w=34800 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1865 GND GND diff_552450_2137300# GND efet w=27550 l=10875
+ ad=0 pd=0 as=2.98555e+08 ps=104400 
M1866 diff_552450_2137300# GND GND GND efet w=5800 l=27550
+ ad=0 pd=0 as=0 ps=0 
M1867 diff_640900_2343200# GND GND GND efet w=6525 l=28275
+ ad=0 pd=0 as=0 ps=0 
M1868 diff_532150_2082200# diff_595950_2080750# GND GND efet w=6525 l=28275
+ ad=8.5782e+08 pd=362500 as=0 ps=0 
M1869 GND diff_532150_2082200# GND GND efet w=37700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1870 GND GND diff_595950_2080750# GND efet w=5800 l=13775
+ ad=0 pd=0 as=4.6255e+07 ps=29000 
M1871 GND diff_249400_1373150# diff_784450_2395400# GND efet w=15225 l=12325
+ ad=0 pd=0 as=9.251e+08 ps=298700 
M1872 GND GND diff_784450_2395400# GND efet w=12325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1873 GND GND diff_935250_2476600# GND efet w=6525 l=51475
+ ad=0 pd=0 as=3.46913e+08 ps=98600 
M1874 diff_784450_2395400# GND GND GND efet w=5800 l=66700
+ ad=0 pd=0 as=0 ps=0 
M1875 diff_935250_2476600# GND GND GND efet w=14500 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1876 GND GND diff_872900_2288100# GND efet w=5800 l=27550
+ ad=0 pd=0 as=7.1485e+08 ps=223300 
M1877 GND GND GND GND efet w=5800 l=29000
+ ad=0 pd=0 as=0 ps=0 
M1878 diff_1097650_2396850# GND GND GND efet w=7975 l=54375
+ ad=1.39185e+09 pd=339300 as=0 ps=0 
M1879 diff_1120850_2447600# GND diff_1097650_2396850# GND efet w=9425 l=15225
+ ad=1.49278e+08 pd=66700 as=0 ps=0 
M1880 diff_1329650_2521550# GND GND GND efet w=6525 l=73225
+ ad=0 pd=0 as=0 ps=0 
M1881 GND diff_1331100_2717300# diff_1329650_2521550# GND efet w=11600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1882 GND diff_1331100_2717300# diff_1200600_2607100# GND efet w=18850 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1883 diff_1200600_2607100# GND GND GND efet w=7975 l=68875
+ ad=0 pd=0 as=0 ps=0 
M1884 diff_1331100_2717300# diff_1329650_2521550# GND GND efet w=13050 l=11600
+ ad=-1.68576e+09 pd=806200 as=0 ps=0 
M1885 GND GND diff_1331100_2717300# GND efet w=6525 l=65250
+ ad=0 pd=0 as=0 ps=0 
M1886 diff_1415200_2605650# diff_1329650_2521550# GND GND efet w=14500 l=11600
+ ad=5.17215e+08 pd=165300 as=0 ps=0 
M1887 GND GND diff_1415200_2605650# GND efet w=9425 l=76125
+ ad=0 pd=0 as=0 ps=0 
M1888 diff_1336900_2549100# GND diff_1200600_2607100# GND efet w=8700 l=10875
+ ad=6.09725e+07 pd=34800 as=0 ps=0 
M1889 diff_1415200_2605650# GND diff_1390550_2521550# GND efet w=7250 l=10150
+ ad=0 pd=0 as=6.3075e+07 ps=31900 
M1890 diff_1693600_2615800# GND diff_1619650_2578100# GND efet w=7975 l=15225
+ ad=0 pd=0 as=5.046e+07 ps=29000 
M1891 diff_1629800_2623050# diff_1610950_2605650# diff_1626900_2588250# GND efet w=24650 l=12325
+ ad=0 pd=0 as=2.39685e+08 ps=87000 
M1892 diff_1626900_2588250# diff_1619650_2578100# GND GND efet w=34075 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1893 GND diff_1699400_2604200# diff_1693600_2615800# GND efet w=21750 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1894 GND diff_1699400_2604200# diff_1629800_2623050# GND efet w=12325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1895 GND GND diff_1790750_2624500# GND efet w=7975 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1896 diff_1790750_2624500# diff_1629800_2623050# GND GND efet w=12325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1897 diff_1699400_2604200# diff_1629800_2623050# GND GND efet w=12325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1898 diff_1982150_2614350# diff_1629800_2623050# diff_1908200_2576650# GND efet w=10150 l=12325
+ ad=0 pd=0 as=3.99475e+07 ps=29000 
M1899 GND diff_1336900_2549100# diff_1355750_2514300# GND efet w=39150 l=13050
+ ad=0 pd=0 as=2.24968e+08 ps=84100 
M1900 GND GND diff_1239750_2443250# GND efet w=7250 l=65250
+ ad=0 pd=0 as=4.205e+08 ps=171100 
M1901 diff_1270200_2518650# GND GND GND efet w=6525 l=28275
+ ad=0 pd=0 as=0 ps=0 
M1902 diff_1355750_2514300# diff_1331100_2717300# diff_1329650_2521550# GND efet w=19575 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1903 diff_1402150_2514300# diff_1390550_2521550# GND GND efet w=39150 l=11600
+ ad=2.24968e+08 pd=81200 as=0 ps=0 
M1904 diff_1331100_2717300# diff_1331100_2717300# diff_1402150_2514300# GND efet w=16675 l=16675
+ ad=0 pd=0 as=0 ps=0 
M1905 GND diff_1500750_2386700# GND GND efet w=40600 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1906 GND diff_1239750_2443250# diff_1270200_2518650# GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1907 GND GND diff_1158550_2475150# GND efet w=5800 l=36250
+ ad=0 pd=0 as=5.67675e+08 ps=182700 
M1908 diff_1331100_2717300# diff_1325300_2459200# GND GND efet w=26825 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1909 GND diff_1075900_2275050# GND GND efet w=31175 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1910 diff_1699400_2604200# diff_1610950_2605650# diff_1840050_2588250# GND efet w=21025 l=12325
+ ad=0 pd=0 as=2.4389e+08 ps=84100 
M1911 diff_2117000_2625950# diff_1629800_2623050# diff_2079300_2623050# GND efet w=8700 l=13050
+ ad=5.887e+07 pd=34800 as=0 ps=0 
M1912 GND diff_1919800_2605650# diff_2079300_2623050# GND efet w=13050 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1913 diff_1919800_2605650# diff_1699400_2604200# diff_1915450_2589700# GND efet w=21750 l=13050
+ ad=0 pd=0 as=2.45992e+08 ps=84100 
M1914 GND diff_1987950_2604200# diff_1982150_2614350# GND efet w=21750 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1915 diff_1919800_2605650# diff_1987950_2604200# GND GND efet w=11600 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1916 diff_1840050_2588250# GND GND GND efet w=25375 l=23200
+ ad=0 pd=0 as=0 ps=0 
M1917 diff_1915450_2589700# diff_1908200_2576650# GND GND efet w=33350 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1918 GND GND GND GND efet w=29000 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1919 GND GND diff_1331100_2717300# GND efet w=9425 l=30450
+ ad=0 pd=0 as=0 ps=0 
M1920 GND GND diff_1289050_2415700# GND efet w=29725 l=15225
+ ad=0 pd=0 as=2.96453e+08 ps=89900 
M1921 diff_1289050_2415700# GND diff_1270200_2417150# GND efet w=31175 l=12325
+ ad=0 pd=0 as=2.14455e+08 ps=75400 
M1922 GND GND diff_872900_2288100# GND efet w=26100 l=13775
+ ad=0 pd=0 as=0 ps=0 
M1923 GND diff_1023700_2175000# GND GND efet w=26100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1924 GND diff_249400_1373150# diff_1097650_2396850# GND efet w=18850 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1925 diff_1158550_2475150# GND GND GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1926 diff_1270200_2417150# diff_872900_2288100# diff_1239750_2443250# GND efet w=29000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1927 diff_867100_2254750# diff_249400_1373150# GND GND efet w=21750 l=13050
+ ad=1.57688e+08 pd=58000 as=0 ps=0 
M1928 diff_884500_2331600# GND diff_865650_2222850# GND efet w=7975 l=12325
+ ad=7.569e+07 pd=49300 as=8.41e+08 ps=272600 
M1929 diff_865650_2222850# diff_872900_2288100# diff_867100_2254750# GND efet w=21750 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1930 diff_907700_2450500# GND GND GND efet w=14500 l=10875
+ ad=4.81473e+08 pd=165300 as=0 ps=0 
M1931 GND GND diff_1003400_2257650# GND efet w=5800 l=52200
+ ad=0 pd=0 as=3.04862e+08 ps=113100 
M1932 diff_865650_2222850# GND GND GND efet w=5800 l=65250
+ ad=0 pd=0 as=0 ps=0 
M1933 diff_865650_2222850# diff_136300_2602750# GND GND efet w=14500 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1934 diff_907700_2450500# GND GND GND efet w=7250 l=47850
+ ad=0 pd=0 as=0 ps=0 
M1935 GND GND diff_1097650_2396850# GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1936 GND diff_1075900_2275050# diff_1023700_2217050# GND efet w=29725 l=12325
+ ad=0 pd=0 as=1.56426e+09 ps=423400 
M1937 GND diff_537950_1786400# diff_1003400_2257650# GND efet w=16675 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1938 GND GND diff_1094750_2248950# GND efet w=21750 l=11600
+ ad=0 pd=0 as=1.57688e+08 ps=58000 
M1939 diff_1094750_2248950# diff_537950_2248950# diff_1023700_2175000# GND efet w=25375 l=10875
+ ad=0 pd=0 as=1.65467e+09 ps=414700 
M1940 diff_1023700_2217050# diff_1003400_2257650# diff_1023700_2198200# GND efet w=29725 l=12325
+ ad=0 pd=0 as=2.1025e+08 ps=72500 
M1941 diff_1325300_2459200# GND diff_1325300_2459200# GND efet w=2900 l=66700
+ ad=1.70933e+09 pd=591600 as=0 ps=0 
M1942 diff_1318050_2322900# GND GND GND efet w=30450 l=11600
+ ad=2.20762e+08 pd=75400 as=0 ps=0 
M1943 diff_1336900_2322900# diff_249400_1373150# diff_1318050_2322900# GND efet w=31900 l=11600
+ ad=2.1866e+08 pd=78300 as=0 ps=0 
M1944 diff_1325300_2459200# diff_1075900_2275050# diff_1336900_2322900# GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1945 GND GND diff_1392000_2341750# GND efet w=5800 l=33350
+ ad=0 pd=0 as=3.5322e+08 ps=130500 
M1946 GND GND diff_1448550_2322900# GND efet w=5800 l=70325
+ ad=0 pd=0 as=9.90278e+08 ps=275500 
M1947 diff_1500750_2386700# GND diff_1448550_2322900# GND efet w=13050 l=13050
+ ad=9.04075e+07 pd=43500 as=0 ps=0 
M1948 GND GND diff_1392000_2341750# GND efet w=21750 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1949 diff_1987950_2604200# diff_1919800_2605650# GND GND efet w=12325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M1950 diff_1987950_2604200# diff_1699400_2604200# diff_2134400_2586800# GND efet w=21750 l=13050
+ ad=0 pd=0 as=2.41788e+08 ps=87000 
M1951 diff_2134400_2586800# diff_2117000_2625950# GND GND efet w=36250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1952 GND diff_2282300_2737600# diff_2215600_2913050# GND efet w=10150 l=13050
+ ad=0 pd=0 as=1.3435e+09 ps=327700 
M1953 GND GND diff_2212700_2604200# GND efet w=5800 l=65250
+ ad=0 pd=0 as=1.10381e+09 ps=214600 
M1954 GND GND diff_2280850_2602750# GND efet w=6525 l=67425
+ ad=0 pd=0 as=1.35401e+09 ps=290000 
M1955 GND GND diff_2373650_2621600# GND efet w=7250 l=69600
+ ad=0 pd=0 as=3.9527e+08 ps=124700 
M1956 diff_2215600_2913050# diff_1668950_2660750# diff_2275050_2614350# GND efet w=7250 l=11600
+ ad=0 pd=0 as=1.02602e+09 ps=223300 
M1957 GND GND diff_2275050_2614350# GND efet w=5075 l=34075
+ ad=0 pd=0 as=0 ps=0 
M1958 diff_2275050_2614350# diff_1919800_2605650# diff_2201100_2576650# GND efet w=7975 l=12325
+ ad=0 pd=0 as=3.99475e+07 ps=34800 
M1959 diff_2212700_2604200# diff_1987950_2604200# diff_2209800_2586800# GND efet w=21025 l=12325
+ ad=0 pd=0 as=2.75427e+08 ps=87000 
M1960 GND diff_2280850_2602750# diff_2275050_2614350# GND efet w=21750 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1961 diff_2212700_2604200# diff_2280850_2602750# GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1962 diff_2209800_2586800# diff_2201100_2576650# GND GND efet w=36250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1963 GND diff_1919800_2605650# diff_2373650_2621600# GND efet w=10875 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1964 diff_2373650_2621600# diff_2212700_2604200# GND GND efet w=11600 l=10150
+ ad=0 pd=0 as=0 ps=0 
M1965 diff_2280850_2602750# diff_2212700_2604200# GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1966 GND GND GND GND efet w=5800 l=51475
+ ad=0 pd=0 as=0 ps=0 
M1967 GND diff_1969100_2514300# diff_1489150_3117500# GND efet w=24650 l=11600
+ ad=0 pd=0 as=1.22576e+09 ps=272600 
M1968 GND diff_2021300_2420050# diff_1610950_2605650# GND efet w=21025 l=12325
+ ad=0 pd=0 as=6.87518e+08 ps=208800 
M1969 diff_2072050_2521550# diff_2063350_2495450# diff_2072050_2521550# GND efet w=55825 l=27550
+ ad=-1.64792e+09 pd=875800 as=0 ps=0 
M1970 diff_1425350_3181300# diff_1075900_2275050# GND GND efet w=39150 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1971 GND GND diff_1660250_2388150# GND efet w=5800 l=71050
+ ad=0 pd=0 as=9.62945e+08 ps=261000 
M1972 GND diff_1706650_2405550# diff_1425350_3181300# GND efet w=36975 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1973 GND diff_1392000_2341750# diff_1331100_2717300# GND efet w=29725 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1974 diff_1660250_2388150# GND diff_1706650_2405550# GND efet w=16675 l=10875
+ ad=0 pd=0 as=1.15638e+08 ps=55100 
M1975 diff_1429700_2322900# GND GND GND efet w=22475 l=12325
+ ad=1.55585e+08 pd=58000 as=0 ps=0 
M1976 diff_1470300_2340300# diff_1452900_2244600# diff_1448550_2322900# GND efet w=32625 l=13775
+ ad=2.1866e+08 pd=78300 as=0 ps=0 
M1977 diff_1448550_2322900# GND diff_1429700_2322900# GND efet w=21750 l=12325
+ ad=0 pd=0 as=0 ps=0 
M1978 diff_1492050_2322900# diff_249400_1373150# diff_1470300_2340300# GND efet w=29725 l=13775
+ ad=1.7661e+08 pd=72500 as=0 ps=0 
M1979 diff_249400_1373150# GND GND GND efet w=23925 l=12325
+ ad=-4.41867e+08 pd=3.9411e+06 as=0 ps=0 
M1980 diff_1023700_2198200# diff_622050_2318550# diff_1023700_2175000# GND efet w=29000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1981 diff_1023700_2175000# GND diff_1023700_2217050# GND efet w=21750 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1982 diff_249400_1373150# diff_249400_1373150# diff_1325300_2459200# GND efet w=23925 l=15225
+ ad=0 pd=0 as=0 ps=0 
M1983 diff_1325300_2459200# GND diff_249400_1373150# GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M1984 diff_1325300_2459200# diff_249400_1373150# diff_249400_1373150# GND efet w=21750 l=13050
+ ad=0 pd=0 as=0 ps=0 
M1985 GND GND diff_1492050_2322900# GND efet w=17400 l=26100
+ ad=0 pd=0 as=0 ps=0 
M1986 GND GND diff_1425350_3181300# GND efet w=34800 l=15950
+ ad=0 pd=0 as=0 ps=0 
M1987 diff_1660250_2388150# diff_249400_1373150# diff_1638500_2367850# GND efet w=31175 l=15225
+ ad=0 pd=0 as=1.31827e+09 ps=382800 
M1988 GND diff_249400_1373150# diff_1552950_2298250# GND efet w=42775 l=13775
+ ad=0 pd=0 as=7.21158e+08 ps=269700 
M1989 GND GND diff_1075900_2275050# GND efet w=8700 l=24650
+ ad=0 pd=0 as=1.02392e+09 ps=345100 
M1990 diff_1489150_3117500# GND GND GND efet w=5800 l=33350
+ ad=0 pd=0 as=0 ps=0 
M1991 diff_1892250_2309850# GND GND GND efet w=5800 l=69600
+ ad=7.27465e+08 pd=278400 as=0 ps=0 
M1992 GND GND diff_1425350_3181300# GND efet w=7250 l=29000
+ ad=0 pd=0 as=0 ps=0 
M1993 diff_1610950_2605650# GND GND GND efet w=5800 l=36250
+ ad=0 pd=0 as=0 ps=0 
M1994 diff_2072050_2521550# diff_2063350_2495450# GND GND efet w=10150 l=27550
+ ad=0 pd=0 as=0 ps=0 
M1995 diff_2072050_2521550# diff_2108300_2408450# GND GND efet w=37700 l=14500
+ ad=0 pd=0 as=0 ps=0 
M1996 diff_2280850_2602750# diff_1987950_2604200# diff_2427300_2585350# GND efet w=24650 l=15950
+ ad=0 pd=0 as=2.4389e+08 ps=84100 
M1997 diff_2427300_2585350# GND GND GND efet w=21750 l=23200
+ ad=0 pd=0 as=0 ps=0 
M1998 GND diff_2179350_2360600# diff_2201100_2537500# GND efet w=12325 l=12325
+ ad=0 pd=0 as=8.2418e+08 ps=298700 
M1999 diff_2201100_2537500# diff_2192400_2495450# diff_2201100_2537500# GND efet w=52925 l=29000
+ ad=0 pd=0 as=0 ps=0 
M2000 GND diff_2192400_2495450# diff_2201100_2537500# GND efet w=6525 l=54375
+ ad=0 pd=0 as=0 ps=0 
M2001 GND diff_2179350_2360600# diff_1687800_3033400# GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2002 GND diff_2322900_2508500# diff_2404100_2504150# GND efet w=11600 l=11600
+ ad=0 pd=0 as=3.42707e+08 ps=142100 
M2003 diff_2322900_2508500# diff_2314200_2449050# diff_2322900_2508500# GND efet w=52925 l=18125
+ ad=-1.94858e+09 pd=690200 as=0 ps=0 
M2004 diff_1687800_3033400# diff_2201100_2537500# GND GND efet w=18850 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2005 diff_1613850_2840550# diff_2404100_2504150# GND GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2006 diff_2063350_2495450# GND GND GND efet w=6525 l=10875
+ ad=5.67675e+07 pd=34800 as=0 ps=0 
M2007 diff_1425350_3181300# diff_1892250_2309850# GND GND efet w=33350 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2008 diff_1638500_2367850# diff_1080250_1561650# diff_1638500_2351900# GND efet w=52925 l=12325
+ ad=0 pd=0 as=3.72142e+08 ps=118900 
M2009 diff_1571800_2293900# diff_1080250_1561650# diff_1552950_2298250# GND efet w=80475 l=13050
+ ad=3.55322e+08 pd=133400 as=0 ps=0 
M2010 GND GND diff_1571800_2293900# GND efet w=38425 l=18125
+ ad=0 pd=0 as=0 ps=0 
M2011 GND GND diff_1638500_2351900# GND efet w=25375 l=16675
+ ad=0 pd=0 as=0 ps=0 
M2012 GND GND diff_1732750_2273600# GND efet w=29725 l=13775
+ ad=0 pd=0 as=6.24442e+08 ps=188500 
M2013 diff_1075900_2275050# GND GND GND efet w=60175 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2014 GND GND diff_1638500_2367850# GND efet w=21750 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2015 diff_1452900_2244600# diff_1080250_1561650# GND GND efet w=55100 l=11600
+ ad=9.71355e+08 pd=255200 as=0 ps=0 
M2016 GND diff_1075900_2275050# diff_1850200_2324350# GND efet w=30450 l=11600
+ ad=0 pd=0 as=2.20762e+08 ps=75400 
M2017 diff_1850200_2324350# GND diff_1850200_2308400# GND efet w=31175 l=10875
+ ad=0 pd=0 as=7.21158e+08 ps=205900 
M2018 diff_2021300_2420050# GND GND GND efet w=5800 l=71050
+ ad=4.2891e+08 pd=130500 as=0 ps=0 
M2019 GND GND diff_2108300_2408450# GND efet w=5800 l=71050
+ ad=0 pd=0 as=1.19842e+09 ps=345100 
M2020 diff_2192400_2495450# GND GND GND efet w=7250 l=11600
+ ad=6.3075e+07 pd=31900 as=0 ps=0 
M2021 diff_2108300_2408450# GND diff_2108300_2347550# GND efet w=30450 l=10150
+ ad=0 pd=0 as=5.15113e+08 ps=165300 
M2022 diff_2021300_2420050# GND diff_2045950_2335950# GND efet w=30450 l=11600
+ ad=0 pd=0 as=4.35218e+08 ps=162400 
M2023 diff_2322900_2508500# diff_2314200_2449050# GND GND efet w=5800 l=52200
+ ad=0 pd=0 as=0 ps=0 
M2024 diff_1732750_2273600# GND diff_1732750_2256200# GND efet w=36975 l=12325
+ ad=0 pd=0 as=7.1485e+08 ps=258100 
M2025 diff_1811050_2224300# diff_1796550_2237350# GND GND efet w=29725 l=14500
+ ad=7.19055e+08 pd=176900 as=0 ps=0 
M2026 diff_1023700_2175000# GND GND GND efet w=5800 l=60900
+ ad=0 pd=0 as=0 ps=0 
M2027 GND GND GND GND efet w=31900 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2028 diff_991800_1986500# GND GND GND efet w=32625 l=10875
+ ad=1.9322e+09 pd=614800 as=0 ps=0 
M2029 GND diff_1075900_2275050# diff_1077350_1464500# GND efet w=24650 l=11600
+ ad=0 pd=0 as=-1.95488e+09 ps=704700 
M2030 diff_1452900_2244600# GND GND GND efet w=5800 l=27550
+ ad=0 pd=0 as=0 ps=0 
M2031 GND diff_1754500_2189500# diff_1712450_2234450# GND efet w=28275 l=14500
+ ad=0 pd=0 as=4.56242e+08 ps=159500 
M2032 diff_1850200_2308400# diff_1080250_1561650# diff_1796550_2237350# GND efet w=54375 l=12325
+ ad=0 pd=0 as=5.5506e+08 ps=176900 
M2033 diff_1712450_2234450# GND GND GND efet w=5800 l=27550
+ ad=0 pd=0 as=0 ps=0 
M2034 diff_1932850_2308400# diff_1811050_2224300# diff_1914000_2251850# GND efet w=34075 l=15950
+ ad=1.80815e+08 pd=78300 as=6.0552e+08 ps=261000 
M2035 GND GND diff_1932850_2308400# GND efet w=34075 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2036 diff_1979250_2308400# diff_249400_1373150# GND GND efet w=31175 l=13775
+ ad=1.7661e+08 pd=72500 as=0 ps=0 
M2037 diff_1998100_2237350# diff_1811050_2224300# diff_1979250_2308400# GND efet w=30450 l=13050
+ ad=6.728e+08 pd=229100 as=0 ps=0 
M2038 diff_1914000_2251850# GND diff_1892250_2309850# GND efet w=34075 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2039 diff_1932850_2225750# diff_1080250_1561650# diff_1914000_2251850# GND efet w=53650 l=13775
+ ad=2.523e+08 pd=113100 as=0 ps=0 
M2040 diff_1754500_2189500# GND diff_1732750_2256200# GND efet w=31175 l=12325
+ ad=2.92247e+08 pd=101500 as=0 ps=0 
M2041 GND GND diff_1754500_2189500# GND efet w=6525 l=64525
+ ad=0 pd=0 as=0 ps=0 
M2042 diff_1811050_2224300# GND GND GND efet w=5800 l=27550
+ ad=0 pd=0 as=0 ps=0 
M2043 diff_1979250_2237350# diff_1712450_2234450# GND GND efet w=31175 l=13775
+ ad=1.7661e+08 pd=72500 as=0 ps=0 
M2044 GND diff_1712450_2234450# diff_1932850_2225750# GND efet w=30450 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2045 diff_1998100_2237350# diff_1452900_2244600# diff_1979250_2237350# GND efet w=30450 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2046 diff_2127150_2344650# GND diff_2108300_2347550# GND efet w=32625 l=15225
+ ad=6.26545e+08 pd=185600 as=0 ps=0 
M2047 diff_2064800_2330150# diff_258100_549550# diff_2045950_2335950# GND efet w=32625 l=13775
+ ad=1.7661e+08 pd=72500 as=0 ps=0 
M2048 GND GND diff_2064800_2330150# GND efet w=30450 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2049 GND diff_249400_1373150# diff_2127150_2344650# GND efet w=31175 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2050 GND GND diff_2179350_2360600# GND efet w=7250 l=68150
+ ad=0 pd=0 as=1.63995e+09 ps=501700 
M2051 diff_2314200_2449050# GND GND GND efet w=6525 l=10875
+ ad=5.046e+07 pd=29000 as=0 ps=0 
M2052 GND GND diff_2404100_2504150# GND efet w=5800 l=52200
+ ad=0 pd=0 as=0 ps=0 
M2053 diff_2179350_2360600# GND diff_2179350_2344650# GND efet w=36975 l=10875
+ ad=0 pd=0 as=3.88962e+08 ps=174000 
M2054 GND GND diff_2176450_2302600# GND efet w=30450 l=11600
+ ad=0 pd=0 as=1.61893e+09 ps=348000 
M2055 diff_2218500_2198200# diff_249400_1373150# diff_2172100_2192400# GND efet w=84825 l=16675
+ ad=-1.8813e+09 pd=672800 as=-1.98011e+09 ps=667000 
M2056 diff_2176450_2302600# diff_258100_549550# GND GND efet w=36250 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2057 GND diff_258100_694550# diff_2127150_2344650# GND efet w=29725 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2058 diff_1969100_2514300# GND diff_1998100_2237350# GND efet w=31900 l=13050
+ ad=4.47833e+08 pd=118900 as=0 ps=0 
M2059 GND GND diff_1969100_2514300# GND efet w=7975 l=67425
+ ad=0 pd=0 as=0 ps=0 
M2060 diff_1796550_2237350# GND GND GND efet w=5800 l=65250
+ ad=0 pd=0 as=0 ps=0 
M2061 diff_2176450_2302600# GND diff_2179350_2344650# GND efet w=34075 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2062 GND GND diff_2172100_2192400# GND efet w=86275 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2063 GND GND diff_1668950_2660750# GND efet w=5800 l=34800
+ ad=0 pd=0 as=-1.85607e+09 ps=600300 
M2064 diff_1613850_2840550# diff_2322900_2508500# GND GND efet w=21750 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2065 GND GND diff_2485300_2392500# GND efet w=9425 l=65975
+ ad=0 pd=0 as=3.25887e+08 ps=101500 
M2066 GND GND diff_2282300_2737600# GND efet w=7975 l=25375
+ ad=0 pd=0 as=8.2418e+08 ps=232000 
M2067 diff_2282300_2737600# diff_2485300_2392500# GND GND efet w=37700 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2068 diff_2322900_2508500# diff_2335950_2264900# GND GND efet w=13775 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2069 GND GND diff_2322900_2508500# GND efet w=16675 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2070 diff_2485300_2392500# diff_249400_1373150# diff_2485300_2375100# GND efet w=32625 l=12325
+ ad=0 pd=0 as=2.79633e+08 ps=95700 
M2071 GND diff_2430200_2244600# diff_1668950_2660750# GND efet w=25375 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2072 diff_2161950_1146950# GND diff_2218500_2198200# GND efet w=14500 l=13050
+ ad=-7.08102e+08 pd=783000 as=0 ps=0 
M2073 diff_2495450_2354800# GND diff_2485300_2375100# GND efet w=30450 l=11600
+ ad=2.20762e+08 pd=75400 as=0 ps=0 
M2074 diff_2495450_2354800# GND GND GND efet w=28275 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2075 diff_2379450_2250400# diff_249400_1373150# GND GND efet w=31175 l=12325
+ ad=7.54798e+08 pd=220400 as=0 ps=0 
M2076 diff_1181750_1322400# GND GND GND efet w=30450 l=15225
+ ad=-1.86868e+09 pd=730800 as=0 ps=0 
M2077 GND GND GND GND efet w=30450 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2078 GND GND GND GND efet w=52925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2079 GND GND diff_842450_2070600# GND efet w=47850 l=11600
+ ad=0 pd=0 as=-4.99955e+08 ps=1.0005e+06 
M2080 GND GND GND GND efet w=31175 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2081 GND GND GND GND efet w=30450 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2082 GND GND GND GND efet w=31175 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2083 diff_622050_2318550# GND GND GND efet w=50025 l=11600
+ ad=-1.30101e+09 pd=759800 as=0 ps=0 
M2084 GND GND GND GND efet w=25375 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2085 GND GND GND GND efet w=23925 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2086 diff_629300_1979250# GND GND GND efet w=6525 l=35525
+ ad=6.28647e+08 pd=226200 as=0 ps=0 
M2087 diff_532150_2082200# diff_595950_2080750# diff_532150_2082200# GND efet w=69600 l=5075
+ ad=0 pd=0 as=0 ps=0 
M2088 GND diff_569850_2003900# GND GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2089 diff_532150_2082200# diff_569850_2003900# GND GND efet w=29000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2090 GND GND diff_791700_1716800# GND efet w=24650 l=11600
+ ad=0 pd=0 as=1.88174e+09 ps=574200 
M2091 GND GND GND GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2092 GND GND diff_537950_2248950# GND efet w=44950 l=11600
+ ad=0 pd=0 as=-1.01717e+09 ps=756900 
M2093 GND GND GND GND efet w=44225 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2094 GND GND diff_1077350_1464500# GND efet w=23200 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2095 diff_791700_1716800# diff_842450_2070600# GND GND efet w=31175 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2096 GND diff_842450_2070600# GND GND efet w=29725 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2097 diff_991800_1986500# diff_842450_2070600# GND GND efet w=31175 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2098 GND diff_842450_2070600# GND GND efet w=55825 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2099 GND GND GND GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2100 GND GND GND GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2101 GND GND GND GND efet w=31900 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2102 GND diff_136300_2602750# diff_2379450_2250400# GND efet w=29725 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2103 diff_2379450_2250400# GND diff_2360600_2244600# GND efet w=34075 l=13775
+ ad=0 pd=0 as=2.31275e+08 ps=87000 
M2104 GND GND diff_2172100_2192400# GND efet w=81925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2105 GND diff_136300_2602750# diff_2218500_2198200# GND efet w=51475 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2106 diff_2218500_2198200# GND GND GND efet w=36975 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2107 GND diff_2161950_1146950# diff_2161950_1146950# GND efet w=47850 l=18850
+ ad=0 pd=0 as=0 ps=0 
M2108 diff_2161950_1146950# diff_2161950_1146950# GND GND efet w=60900 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2109 diff_2360600_2244600# GND diff_2335950_2264900# GND efet w=30450 l=8700
+ ad=0 pd=0 as=5.69777e+08 ps=185600 
M2110 GND GND diff_2505600_2279400# GND efet w=29725 l=10875
+ ad=0 pd=0 as=3.0276e+08 ps=81200 
M2111 diff_2505600_2279400# GND diff_2505600_2260550# GND efet w=29725 l=10875
+ ad=0 pd=0 as=2.58608e+08 ps=78300 
M2112 diff_2459200_2230100# diff_258100_694550# diff_2430200_2244600# GND efet w=23925 l=9425
+ ad=1.682e+08 pd=60900 as=3.7004e+08 ps=127600 
M2113 GND GND diff_2459200_2230100# GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2114 diff_2505600_2260550# GND diff_2505600_2241700# GND efet w=30450 l=10150
+ ad=0 pd=0 as=3.4481e+08 ps=116000 
M2115 diff_2218500_2198200# GND GND GND efet w=7250 l=37700
+ ad=0 pd=0 as=0 ps=0 
M2116 GND GND diff_2335950_2264900# GND efet w=6525 l=64525
+ ad=0 pd=0 as=0 ps=0 
M2117 GND GND GND GND efet w=42775 l=18125
+ ad=0 pd=0 as=0 ps=0 
M2118 diff_842450_2070600# GND GND GND efet w=35525 l=18125
+ ad=0 pd=0 as=0 ps=0 
M2119 GND diff_842450_2070600# diff_1149850_1992300# GND efet w=92075 l=10875
+ ad=0 pd=0 as=2.13193e+09 ps=426300 
M2120 diff_1077350_1464500# diff_842450_2070600# GND GND efet w=30450 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2121 GND diff_842450_2070600# GND GND efet w=30450 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2122 diff_703250_1961850# diff_622050_2318550# diff_677150_1960400# GND efet w=36250 l=15950
+ ad=1.53272e+09 pd=446600 as=1.37924e+09 ps=362500 
M2123 diff_677150_1960400# GND diff_703250_1961850# GND efet w=33350 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2124 GND diff_842450_2070600# GND GND efet w=31900 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2125 GND GND GND GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2126 GND GND GND GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2127 GND diff_842450_2070600# GND GND efet w=56550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2128 diff_842450_2070600# diff_842450_2070600# GND GND efet w=45675 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2129 GND diff_842450_2070600# GND GND efet w=32625 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2130 diff_1149850_1992300# GND diff_622050_2318550# GND efet w=98600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2131 GND GND GND GND efet w=18850 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2132 GND GND GND GND efet w=21025 l=16675
+ ad=0 pd=0 as=0 ps=0 
M2133 GND GND GND GND efet w=20300 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2134 GND diff_842450_2070600# GND GND efet w=32625 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2135 GND GND diff_537950_2248950# GND efet w=44950 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2136 GND GND GND GND efet w=31175 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2137 diff_791700_1716800# GND GND GND efet w=31900 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2138 GND GND diff_1181750_1322400# GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2139 GND GND GND GND efet w=21025 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2140 GND GND GND GND efet w=46400 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2141 GND diff_2093800_1972000# GND GND efet w=47850 l=20300
+ ad=0 pd=0 as=0 ps=0 
M2142 GND GND diff_842450_2070600# GND efet w=33350 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2143 diff_842450_2070600# GND GND GND efet w=36250 l=17400
+ ad=0 pd=0 as=0 ps=0 
M2144 GND GND GND GND efet w=22475 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2145 GND GND GND GND efet w=29725 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2146 GND GND GND GND efet w=29725 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2147 diff_991800_1986500# GND GND GND efet w=30450 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2148 diff_537950_2248950# GND GND GND efet w=53650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2149 diff_1077350_1464500# GND GND GND efet w=29725 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2150 diff_1149850_1992300# GND GND GND efet w=89175 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2151 diff_1181750_1322400# GND GND GND efet w=30450 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2152 GND GND GND GND efet w=20300 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2153 GND GND GND GND efet w=19575 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2154 GND GND GND GND efet w=21025 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2155 GND GND GND GND efet w=57275 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2156 GND GND diff_842450_2070600# GND efet w=45675 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2157 diff_629300_1979250# GND diff_569850_2003900# GND efet w=14500 l=13050
+ ad=0 pd=0 as=3.06965e+08 ps=87000 
M2158 diff_677150_1960400# GND GND GND efet w=37700 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2159 diff_529250_1925600# GND GND GND efet w=7975 l=64525
+ ad=1.4297e+08 pd=75400 as=0 ps=0 
M2160 GND diff_636550_1956050# diff_629300_1979250# GND efet w=22475 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2161 diff_703250_1961850# GND diff_677150_1960400# GND efet w=31900 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2162 diff_620600_1919800# GND diff_703250_1961850# GND efet w=34800 l=11600
+ ad=1.42339e+09 pd=379900 as=0 ps=0 
M2163 GND GND GND GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2164 GND GND GND GND efet w=41325 l=18125
+ ad=0 pd=0 as=0 ps=0 
M2165 GND GND GND GND efet w=23200 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2166 diff_1149850_1992300# GND diff_622050_2318550# GND efet w=96425 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2167 GND GND GND GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2168 GND GND GND GND efet w=21750 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2169 GND GND diff_842450_2070600# GND efet w=42775 l=16675
+ ad=0 pd=0 as=0 ps=0 
M2170 GND GND GND GND efet w=30450 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2171 GND GND GND GND efet w=31900 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2172 GND diff_2093800_1972000# diff_842450_2070600# GND efet w=32625 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2173 GND GND GND GND efet w=29725 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2174 diff_2161950_1146950# GND GND GND efet w=10150 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2175 GND diff_2208350_2030000# GND GND efet w=39150 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2176 GND diff_2201100_2086550# GND GND efet w=20300 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2177 GND GND diff_2430200_2244600# GND efet w=7250 l=60900
+ ad=0 pd=0 as=0 ps=0 
M2178 diff_2505600_2241700# GND GND GND efet w=6525 l=63075
+ ad=0 pd=0 as=0 ps=0 
M2179 GND diff_2505600_2241700# diff_2534600_2179350# GND efet w=36975 l=9425
+ ad=0 pd=0 as=3.6163e+08 ps=124700 
M2180 diff_2534600_2179350# GND GND GND efet w=6525 l=26100
+ ad=0 pd=0 as=0 ps=0 
M2181 GND diff_2534600_2179350# diff_2317100_1996650# GND efet w=11600 l=12325
+ ad=0 pd=0 as=2.79633e+08 ps=81200 
M2182 GND diff_2534600_2179350# diff_2382350_1993750# GND efet w=10875 l=11600
+ ad=0 pd=0 as=2.62812e+08 ps=84100 
M2183 GND diff_2201100_2086550# GND GND efet w=29725 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2184 GND diff_2208350_2030000# GND GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2185 GND GND GND GND efet w=8700 l=30450
+ ad=0 pd=0 as=0 ps=0 
M2186 GND GND GND GND efet w=10150 l=32625
+ ad=0 pd=0 as=0 ps=0 
M2187 GND diff_2317100_1996650# GND GND efet w=58725 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2188 GND diff_2518650_2030000# diff_2201100_2086550# GND efet w=62350 l=11600
+ ad=0 pd=0 as=6.53878e+08 ps=252300 
M2189 GND diff_2534600_2179350# diff_2447600_1993750# GND efet w=10875 l=12325
+ ad=0 pd=0 as=2.7753e+08 ps=81200 
M2190 diff_2153250_1870500# GND GND GND efet w=12325 l=29000
+ ad=5.78188e+08 pd=203000 as=0 ps=0 
M2191 GND diff_2382350_1993750# GND GND efet w=61625 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2192 diff_2201100_2086550# GND GND GND efet w=8700 l=33350
+ ad=0 pd=0 as=0 ps=0 
M2193 GND GND GND GND efet w=23925 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2194 GND GND GND GND efet w=22475 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2195 GND GND GND GND efet w=21750 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2196 diff_791700_1716800# GND GND GND efet w=31900 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2197 GND GND GND GND efet w=30450 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2198 diff_991800_1986500# GND GND GND efet w=30450 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2199 diff_537950_2248950# GND GND GND efet w=52200 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2200 GND GND diff_529250_1925600# GND efet w=12325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2201 diff_601750_1919800# diff_529250_1925600# GND GND efet w=21750 l=11600
+ ad=1.57688e+08 pd=58000 as=0 ps=0 
M2202 diff_620600_1919800# diff_569850_2003900# diff_601750_1919800# GND efet w=21750 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2203 diff_636550_1956050# GND diff_620600_1919800# GND efet w=8700 l=11600
+ ad=1.13535e+08 pd=43500 as=0 ps=0 
M2204 diff_620600_1919800# GND diff_620600_1919800# GND efet w=3625 l=70325
+ ad=0 pd=0 as=0 ps=0 
M2205 diff_1181750_1322400# GND GND GND efet w=29725 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2206 GND GND diff_622050_2318550# GND efet w=52925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2207 GND GND GND GND efet w=31175 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2208 GND GND GND GND efet w=21025 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2209 GND GND diff_842450_2070600# GND efet w=52200 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2210 GND GND GND GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2211 GND GND GND GND efet w=31175 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2212 GND GND GND GND efet w=39875 l=21750
+ ad=0 pd=0 as=0 ps=0 
M2213 GND diff_797500_1757400# GND GND efet w=21750 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2214 GND GND GND GND efet w=21750 l=18850
+ ad=0 pd=0 as=0 ps=0 
M2215 GND GND GND GND efet w=20300 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2216 GND GND diff_526350_1657350# GND efet w=6525 l=39875
+ ad=0 pd=0 as=3.23785e+08 ps=116000 
M2217 GND GND GND GND efet w=7975 l=22475
+ ad=0 pd=0 as=0 ps=0 
M2218 diff_537950_1786400# GND GND GND efet w=10150 l=28275
+ ad=6.58082e+08 pd=182700 as=0 ps=0 
M2219 diff_526350_1657350# diff_258100_549550# GND GND efet w=18125 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2220 GND GND GND GND efet w=5800 l=59450
+ ad=0 pd=0 as=0 ps=0 
M2221 GND GND GND GND efet w=18850 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2222 GND diff_2035800_1877750# GND GND efet w=20300 l=17400
+ ad=0 pd=0 as=0 ps=0 
M2223 GND GND GND GND efet w=24650 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2224 GND GND GND GND efet w=18850 l=16675
+ ad=0 pd=0 as=0 ps=0 
M2225 diff_791700_1716800# GND GND GND efet w=7250 l=63800
+ ad=0 pd=0 as=0 ps=0 
M2226 GND GND GND GND efet w=5800 l=62350
+ ad=0 pd=0 as=0 ps=0 
M2227 GND GND GND GND efet w=5800 l=63075
+ ad=0 pd=0 as=0 ps=0 
M2228 GND GND GND GND efet w=9425 l=73225
+ ad=0 pd=0 as=0 ps=0 
M2229 diff_665550_1548600# GND GND GND efet w=7250 l=72500
+ ad=4.83575e+08 pd=153700 as=0 ps=0 
M2230 GND GND diff_991800_1986500# GND efet w=7250 l=56550
+ ad=0 pd=0 as=0 ps=0 
M2231 diff_537950_2248950# GND GND GND efet w=7250 l=36975
+ ad=0 pd=0 as=0 ps=0 
M2232 GND GND diff_1025150_1793650# GND efet w=7250 l=50750
+ ad=0 pd=0 as=2.1866e+08 ps=89900 
M2233 GND GND GND GND efet w=8700 l=39150
+ ad=0 pd=0 as=0 ps=0 
M2234 diff_622050_2318550# GND GND GND efet w=8700 l=34800
+ ad=0 pd=0 as=0 ps=0 
M2235 diff_1077350_1464500# GND GND GND efet w=7250 l=55100
+ ad=0 pd=0 as=0 ps=0 
M2236 GND GND GND GND efet w=5800 l=63800
+ ad=0 pd=0 as=0 ps=0 
M2237 GND diff_797500_1757400# diff_903350_1763200# GND efet w=38425 l=10875
+ ad=0 pd=0 as=2.64915e+08 ps=95700 
M2238 diff_903350_1763200# GND diff_688750_1509450# GND efet w=23200 l=13050
+ ad=0 pd=0 as=7.46388e+08 ps=234900 
M2239 GND GND diff_740950_1728400# GND efet w=33350 l=10150
+ ad=0 pd=0 as=2.71222e+08 ps=87000 
M2240 GND reset diff_497350_1687800# GND efet w=35525 l=12325
+ ad=0 pd=0 as=9.77663e+08 ps=252300 
M2241 GND GND diff_537950_1786400# GND efet w=51475 l=18850
+ ad=0 pd=0 as=0 ps=0 
M2242 GND diff_497350_1687800# diff_526350_1657350# GND efet w=19575 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2243 GND diff_497350_1687800# GND GND efet w=55825 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2244 diff_668450_1715350# GND GND GND efet w=21750 l=13050
+ ad=2.523e+08 pd=89900 as=0 ps=0 
M2245 diff_674250_1700850# GND GND GND efet w=13775 l=12325
+ ad=1.7661e+08 pd=87000 as=0 ps=0 
M2246 diff_740950_1728400# GND diff_740950_1709550# GND efet w=34075 l=10875
+ ad=0 pd=0 as=2.64915e+08 ps=78300 
M2247 GND GND diff_665550_1548600# GND efet w=13775 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2248 diff_1025150_1793650# diff_991800_1986500# GND GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2249 GND diff_1025150_1793650# GND GND efet w=29000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2250 GND GND diff_665550_1548600# GND efet w=34800 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2251 diff_665550_1548600# diff_665550_1548600# GND GND efet w=7975 l=18125
+ ad=0 pd=0 as=0 ps=0 
M2252 GND diff_791700_1716800# diff_797500_1693600# GND efet w=13050 l=11600
+ ad=0 pd=0 as=3.99475e+08 ps=95700 
M2253 GND GND diff_826500_1682000# GND efet w=8700 l=17400
+ ad=0 pd=0 as=4.22602e+08 ps=147900 
M2254 GND diff_991800_1986500# GND GND efet w=29725 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2255 GND GND GND GND efet w=7250 l=53650
+ ad=0 pd=0 as=0 ps=0 
M2256 GND GND GND GND efet w=5800 l=65975
+ ad=0 pd=0 as=0 ps=0 
M2257 GND GND GND GND efet w=8700 l=43500
+ ad=0 pd=0 as=0 ps=0 
M2258 GND GND GND GND efet w=8700 l=43500
+ ad=0 pd=0 as=0 ps=0 
M2259 diff_1181750_1322400# GND GND GND efet w=5800 l=57275
+ ad=0 pd=0 as=0 ps=0 
M2260 GND GND GND GND efet w=6525 l=57275
+ ad=0 pd=0 as=0 ps=0 
M2261 GND GND GND GND efet w=7250 l=55100
+ ad=0 pd=0 as=0 ps=0 
M2262 GND GND GND GND efet w=6525 l=60900
+ ad=0 pd=0 as=0 ps=0 
M2263 GND GND GND GND efet w=10150 l=65250
+ ad=0 pd=0 as=0 ps=0 
M2264 GND GND diff_1286150_1331100# GND efet w=5800 l=56550
+ ad=0 pd=0 as=7.02235e+08 ps=188500 
M2265 GND GND diff_1400700_1510900# GND efet w=7250 l=55100
+ ad=0 pd=0 as=1.30565e+09 ps=400200 
M2266 GND GND GND GND efet w=6525 l=55100
+ ad=0 pd=0 as=0 ps=0 
M2267 GND GND GND GND efet w=6525 l=55825
+ ad=0 pd=0 as=0 ps=0 
M2268 GND GND GND GND efet w=7250 l=56550
+ ad=0 pd=0 as=0 ps=0 
M2269 GND GND GND GND efet w=5800 l=61625
+ ad=0 pd=0 as=0 ps=0 
M2270 GND GND GND GND efet w=5800 l=65250
+ ad=0 pd=0 as=0 ps=0 
M2271 GND GND GND GND efet w=6525 l=67425
+ ad=0 pd=0 as=0 ps=0 
M2272 GND GND GND GND efet w=7250 l=50750
+ ad=0 pd=0 as=0 ps=0 
M2273 diff_1286150_1331100# diff_665550_1548600# GND GND efet w=38425 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2274 GND GND GND GND efet w=7250 l=53650
+ ad=0 pd=0 as=0 ps=0 
M2275 GND GND GND GND efet w=6525 l=52925
+ ad=0 pd=0 as=0 ps=0 
M2276 GND GND GND GND efet w=5800 l=56550
+ ad=0 pd=0 as=0 ps=0 
M2277 GND GND GND GND efet w=7250 l=63075
+ ad=0 pd=0 as=0 ps=0 
M2278 GND GND GND GND efet w=7250 l=60900
+ ad=0 pd=0 as=0 ps=0 
M2279 GND GND GND GND efet w=7250 l=59450
+ ad=0 pd=0 as=0 ps=0 
M2280 GND GND GND GND efet w=7975 l=58725
+ ad=0 pd=0 as=0 ps=0 
M2281 GND GND GND GND efet w=7250 l=63800
+ ad=0 pd=0 as=0 ps=0 
M2282 GND GND GND GND efet w=7975 l=65250
+ ad=0 pd=0 as=0 ps=0 
M2283 GND GND GND GND efet w=7250 l=56550
+ ad=0 pd=0 as=0 ps=0 
M2284 GND GND GND GND efet w=5800 l=56550
+ ad=0 pd=0 as=0 ps=0 
M2285 GND GND GND GND efet w=21025 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2286 GND diff_2035800_1877750# GND GND efet w=29725 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2287 GND diff_2153250_1870500# GND GND efet w=38425 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2288 GND diff_2153250_1957500# GND GND efet w=24650 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2289 diff_2035800_1877750# GND GND GND efet w=21750 l=17400
+ ad=5.76085e+08 pd=188500 as=0 ps=0 
M2290 GND diff_2447600_1993750# diff_2153250_1870500# GND efet w=58000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2291 diff_2093800_1972000# GND GND GND efet w=23200 l=17400
+ ad=9.8397e+08 pd=263900 as=0 ps=0 
M2292 diff_2153250_1957500# diff_2153250_1870500# GND GND efet w=29000 l=10150
+ ad=6.58082e+08 pd=174000 as=0 ps=0 
M2293 GND diff_2534600_2179350# diff_2518650_2030000# GND efet w=10150 l=12325
+ ad=0 pd=0 as=2.6912e+08 ps=78300 
M2294 diff_2208350_2030000# diff_2201100_2086550# GND GND efet w=26825 l=10875
+ ad=6.20238e+08 pd=179800 as=0 ps=0 
M2295 diff_2035800_1877750# diff_2295350_1931400# diff_2035800_1877750# GND efet w=3625 l=51475
+ ad=0 pd=0 as=0 ps=0 
M2296 GND diff_2153250_1957500# GND GND efet w=34075 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2297 GND diff_2153250_1870500# GND GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2298 diff_2093800_1972000# GND diff_2093800_1972000# GND efet w=4350 l=53650
+ ad=0 pd=0 as=0 ps=0 
M2299 diff_2153250_1957500# GND diff_2153250_1957500# GND efet w=3625 l=42775
+ ad=0 pd=0 as=0 ps=0 
M2300 diff_2208350_2030000# GND diff_2208350_2030000# GND efet w=2900 l=51475
+ ad=0 pd=0 as=0 ps=0 
M2301 GND diff_1999550_1331100# GND GND efet w=58725 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2302 GND GND GND GND efet w=10875 l=41325
+ ad=0 pd=0 as=0 ps=0 
M2303 GND diff_665550_1548600# GND GND efet w=31900 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2304 GND diff_665550_1548600# GND GND efet w=31900 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2305 GND GND diff_1925600_1133900# GND efet w=5800 l=49300
+ ad=0 pd=0 as=6.62287e+08 ps=188500 
M2306 GND diff_846800_1278900# diff_2157600_1809600# GND efet w=13775 l=12325
+ ad=0 pd=0 as=3.1958e+08 ps=121800 
M2307 diff_2157600_1809600# GND GND GND efet w=7250 l=67425
+ ad=0 pd=0 as=0 ps=0 
M2308 diff_2218500_1796550# diff_2157600_1809600# diff_1925600_1133900# GND efet w=27550 l=11600
+ ad=1.8502e+08 pd=69600 as=0 ps=0 
M2309 diff_2179350_1790750# GND GND GND efet w=7250 l=77575
+ ad=2.1025e+08 pd=89900 as=0 ps=0 
M2310 diff_2218500_1796550# diff_2179350_1790750# GND GND efet w=26825 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2311 diff_2179350_1790750# GND GND GND efet w=9425 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2312 diff_668450_1715350# diff_674250_1700850# diff_681500_1692150# GND efet w=20300 l=11600
+ ad=0 pd=0 as=7.16953e+08 ps=188500 
M2313 diff_740950_1709550# diff_733700_1700850# diff_681500_1692150# GND efet w=30450 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2314 GND diff_526350_1657350# diff_497350_1687800# GND efet w=33350 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2315 diff_362500_1632700# GND GND GND efet w=26100 l=11600
+ ad=1.32247e+09 pd=411800 as=0 ps=0 
M2316 diff_362500_1632700# diff_371200_1631250# diff_362500_1632700# GND efet w=74675 l=5075
+ ad=0 pd=0 as=0 ps=0 
M2317 GND GND diff_314650_1616750# GND efet w=10875 l=15225
+ ad=0 pd=0 as=1.38765e+08 ps=58000 
M2318 GND diff_371200_1631250# diff_362500_1632700# GND efet w=7975 l=32625
+ ad=0 pd=0 as=0 ps=0 
M2319 GND GND diff_371200_1631250# GND efet w=5800 l=13050
+ ad=0 pd=0 as=4.6255e+07 ps=29000 
M2320 GND diff_362500_1632700# diff_332050_1580500# GND efet w=27550 l=11600
+ ad=0 pd=0 as=1.04704e+09 ps=284200 
M2321 diff_332050_1580500# diff_314650_1616750# GND GND efet w=62350 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2322 GND GND diff_332050_1580500# GND efet w=7975 l=21025
+ ad=0 pd=0 as=0 ps=0 
M2323 GND GND diff_332050_1580500# GND efet w=11600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2324 diff_633650_1644300# GND GND GND efet w=14500 l=11600
+ ad=3.8686e+08 pd=116000 as=0 ps=0 
M2325 GND diff_640900_1654450# diff_633650_1644300# GND efet w=26825 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2326 diff_681500_1692150# GND diff_640900_1654450# GND efet w=8700 l=11600
+ ad=0 pd=0 as=1.4297e+08 ps=63800 
M2327 GND GND diff_674250_1700850# GND efet w=7250 l=84100
+ ad=0 pd=0 as=0 ps=0 
M2328 GND test diff_519100_1629800# GND efet w=36250 l=10150
+ ad=0 pd=0 as=1.54744e+09 ps=420500 
M2329 GND GND diff_519100_1629800# GND efet w=4350 l=58000
+ ad=0 pd=0 as=0 ps=0 
M2330 diff_497350_1687800# GND GND GND efet w=5800 l=26100
+ ad=0 pd=0 as=0 ps=0 
M2331 GND GND diff_633650_1644300# GND efet w=7250 l=36250
+ ad=0 pd=0 as=0 ps=0 
M2332 GND GND diff_559700_1464500# GND efet w=5800 l=50750
+ ad=0 pd=0 as=3.49015e+08 ps=124700 
M2333 diff_336400_1510900# GND GND GND efet w=31900 l=10875
+ ad=1.14166e+09 pd=362500 as=0 ps=0 
M2334 GND GND GND GND efet w=8700 l=20300
+ ad=0 pd=0 as=0 ps=0 
M2335 diff_681500_1692150# GND GND GND efet w=6525 l=63075
+ ad=0 pd=0 as=0 ps=0 
M2336 diff_797500_1693600# GND GND GND efet w=10875 l=65975
+ ad=0 pd=0 as=0 ps=0 
M2337 GND diff_826500_1682000# diff_852600_1702300# GND efet w=23200 l=11600
+ ad=0 pd=0 as=-2.12729e+09 ps=649600 
M2338 GND GND GND GND efet w=19575 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2339 GND GND GND GND efet w=20300 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2340 GND GND GND GND efet w=23925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2341 GND GND GND GND efet w=38425 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2342 GND GND GND GND efet w=34075 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2343 diff_1400700_1510900# GND GND GND efet w=23925 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2344 GND GND GND GND efet w=23925 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2345 GND GND GND GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2346 diff_852600_1702300# diff_916400_1668950# diff_935250_1697950# GND efet w=44225 l=15225
+ ad=0 pd=0 as=1.06176e+09 ps=330600 
M2347 diff_852600_1702300# GND diff_935250_1697950# GND efet w=63800 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2348 diff_852600_1702300# diff_797500_1693600# diff_733700_1700850# GND efet w=41325 l=13775
+ ad=0 pd=0 as=8.2418e+08 ps=185600 
M2349 GND diff_665550_1548600# GND GND efet w=59450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2350 diff_826500_1682000# GND GND GND efet w=5800 l=58000
+ ad=0 pd=0 as=0 ps=0 
M2351 diff_852600_1702300# diff_871450_1602250# diff_733700_1700850# GND efet w=47125 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2352 diff_733700_1700850# GND GND GND efet w=5800 l=50025
+ ad=0 pd=0 as=0 ps=0 
M2353 GND GND diff_688750_1509450# GND efet w=5800 l=68875
+ ad=0 pd=0 as=0 ps=0 
M2354 GND GND GND GND efet w=30450 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2355 GND GND GND GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2356 GND GND GND GND efet w=40600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2357 GND GND GND GND efet w=40600 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2358 GND GND diff_935250_1697950# GND efet w=46400 l=18850
+ ad=0 pd=0 as=0 ps=0 
M2359 GND GND diff_935250_1697950# GND efet w=75400 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2360 GND GND GND GND efet w=18850 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2361 GND GND GND GND efet w=19575 l=16675
+ ad=0 pd=0 as=0 ps=0 
M2362 GND GND GND GND efet w=19575 l=16675
+ ad=0 pd=0 as=0 ps=0 
M2363 GND GND GND GND efet w=18850 l=17400
+ ad=0 pd=0 as=0 ps=0 
M2364 GND GND GND GND efet w=19575 l=16675
+ ad=0 pd=0 as=0 ps=0 
M2365 GND diff_665550_1548600# GND GND efet w=39875 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2366 diff_1925600_1133900# diff_258100_549550# diff_2041600_1738550# GND efet w=31900 l=11600
+ ad=0 pd=0 as=3.32195e+08 ps=101500 
M2367 GND diff_1999550_1331100# GND GND efet w=61625 l=16675
+ ad=0 pd=0 as=0 ps=0 
M2368 GND GND diff_2041600_1738550# GND efet w=29000 l=17400
+ ad=0 pd=0 as=0 ps=0 
M2369 GND GND GND GND efet w=19575 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2370 GND GND GND GND efet w=19575 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2371 GND GND GND GND efet w=31175 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2372 GND GND GND GND efet w=29725 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2373 GND GND GND GND efet w=32625 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2374 GND GND GND GND efet w=30450 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2375 GND GND GND GND efet w=41325 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2376 GND diff_2085100_1422450# GND GND efet w=29725 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2377 GND GND GND GND efet w=56550 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2378 GND GND GND GND efet w=19575 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2379 GND GND diff_1286150_1331100# GND efet w=31900 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2380 GND GND diff_1400700_1510900# GND efet w=24650 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2381 GND GND GND GND efet w=23925 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2382 GND GND GND GND efet w=23200 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2383 GND GND GND GND efet w=23200 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2384 GND GND GND GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2385 GND GND GND GND efet w=19575 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2386 GND GND diff_916400_1668950# GND efet w=13050 l=11600
+ ad=0 pd=0 as=3.23785e+08 ps=127600 
M2387 GND diff_1080250_1657350# GND GND efet w=30450 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2388 GND GND diff_1016450_1635600# GND efet w=44950 l=14500
+ ad=0 pd=0 as=5.65572e+08 ps=147900 
M2389 diff_1016450_1635600# diff_925100_1455800# GND GND efet w=29000 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2390 diff_916400_1668950# GND GND GND efet w=5800 l=50750
+ ad=0 pd=0 as=0 ps=0 
M2391 GND GND diff_781550_1535550# GND efet w=6525 l=26100
+ ad=0 pd=0 as=7.35875e+08 ps=249400 
M2392 GND diff_1080250_1657350# GND GND efet w=30450 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2393 diff_1400700_1510900# diff_1080250_1657350# GND GND efet w=31900 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2394 GND diff_1080250_1657350# GND GND efet w=31175 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2395 GND GND GND GND efet w=18850 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2396 GND GND GND GND efet w=20300 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2397 GND diff_1080250_1657350# GND GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2398 GND diff_1080250_1657350# GND GND efet w=31175 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2399 GND GND GND GND efet w=5800 l=47850
+ ad=0 pd=0 as=0 ps=0 
M2400 GND GND GND GND efet w=31175 l=16675
+ ad=0 pd=0 as=0 ps=0 
M2401 GND GND GND GND efet w=30450 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2402 GND diff_2215600_1422450# diff_1080250_1657350# GND efet w=36975 l=15225
+ ad=0 pd=0 as=8.2418e+08 ps=226200 
M2403 GND GND GND GND efet w=48575 l=21750
+ ad=0 pd=0 as=0 ps=0 
M2404 GND GND GND GND efet w=22475 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2405 GND diff_2085100_1422450# GND GND efet w=25375 l=9425
+ ad=0 pd=0 as=0 ps=0 
M2406 GND GND GND GND efet w=19575 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2407 GND GND GND GND efet w=21750 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2408 GND GND GND GND efet w=22475 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2409 GND GND GND GND efet w=25375 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2410 GND GND GND GND efet w=25375 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2411 GND GND GND GND efet w=18125 l=18125
+ ad=0 pd=0 as=0 ps=0 
M2412 GND diff_1232500_1610950# GND GND efet w=43500 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2413 GND GND diff_781550_1535550# GND efet w=47850 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2414 GND GND diff_497350_1464500# GND efet w=6525 l=67425
+ ad=0 pd=0 as=1.60631e+09 ps=481400 
M2415 diff_336400_1510900# diff_345100_1497850# diff_336400_1510900# GND efet w=72500 l=5800
+ ad=0 pd=0 as=0 ps=0 
M2416 GND diff_345100_1497850# diff_336400_1510900# GND efet w=6525 l=26825
+ ad=0 pd=0 as=0 ps=0 
M2417 GND GND diff_345100_1497850# GND efet w=5800 l=13050
+ ad=0 pd=0 as=5.25625e+07 ps=34800 
M2418 GND GND GND GND efet w=31175 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2419 GND diff_497350_1464500# diff_559700_1464500# GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2420 GND diff_336400_1510900# GND GND efet w=36250 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2421 diff_858400_1561650# GND diff_258100_694550# GND efet w=8700 l=11600
+ ad=6.93825e+07 pd=34800 as=1.10303e+09 ps=2.9841e+06 
M2422 diff_497350_1464500# diff_688750_1509450# GND GND efet w=13050 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2423 diff_846800_1510900# diff_858400_1561650# GND GND efet w=14500 l=11600
+ ad=4.77267e+08 pd=156600 as=0 ps=0 
M2424 diff_846800_1510900# diff_781550_1535550# diff_810550_1503650# GND efet w=8700 l=13050
+ ad=0 pd=0 as=1.72405e+08 ps=69600 
M2425 GND GND diff_896100_1570350# GND efet w=6525 l=11600
+ ad=0 pd=0 as=3.21682e+08 ps=107300 
M2426 GND diff_896100_1570350# GND GND efet w=5800 l=16675
+ ad=0 pd=0 as=0 ps=0 
M2427 GND diff_896100_1570350# GND GND efet w=69600 l=26825
+ ad=0 pd=0 as=0 ps=0 
M2428 diff_1015000_1583400# diff_667000_980200# GND GND efet w=27550 l=11600
+ ad=4.6255e+08 pd=156600 as=0 ps=0 
M2429 diff_1400700_1510900# diff_1232500_1610950# GND GND efet w=31175 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2430 GND diff_1232500_1610950# GND GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2431 GND GND diff_1015000_1583400# GND efet w=45675 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2432 GND diff_1232500_1610950# GND GND efet w=31900 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2433 GND diff_1232500_1610950# GND GND efet w=31175 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2434 GND diff_1232500_1610950# GND GND efet w=31900 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2435 GND GND GND GND efet w=28275 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2436 GND GND GND GND efet w=21750 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2437 GND diff_1232500_1610950# GND GND efet w=29725 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2438 GND diff_497350_1464500# GND GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2439 GND diff_559700_1464500# GND GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2440 diff_630750_1461600# diff_526350_1077350# diff_497350_1464500# GND efet w=30450 l=10150
+ ad=1.99738e+08 pd=69600 as=0 ps=0 
M2441 GND GND diff_630750_1461600# GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2442 diff_677150_1461600# diff_552450_1347050# GND GND efet w=27550 l=11600
+ ad=5.3824e+08 pd=156600 as=0 ps=0 
M2443 diff_497350_1464500# diff_497350_1464500# diff_677150_1461600# GND efet w=23925 l=18125
+ ad=0 pd=0 as=0 ps=0 
M2444 GND diff_733700_1481900# diff_497350_1464500# GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2445 GND GND diff_785900_1464500# GND efet w=16675 l=12325
+ ad=0 pd=0 as=8.95665e+08 ps=307400 
M2446 diff_733700_1481900# diff_810550_1503650# GND GND efet w=20300 l=12325
+ ad=2.92247e+08 pd=92800 as=0 ps=0 
M2447 GND GND diff_733700_1481900# GND efet w=7975 l=55100
+ ad=0 pd=0 as=0 ps=0 
M2448 GND diff_336400_1363000# GND GND efet w=39150 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2449 GND diff_290000_1419550# GND GND efet w=36975 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2450 GND GND diff_249400_1373150# GND efet w=25375 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2451 diff_336400_1363000# diff_290000_1419550# GND GND efet w=30450 l=11600
+ ad=1.16899e+09 pd=342200 as=0 ps=0 
M2452 diff_336400_1363000# diff_345100_1370250# diff_336400_1363000# GND efet w=70325 l=5800
+ ad=0 pd=0 as=0 ps=0 
M2453 GND GND diff_345100_1370250# GND efet w=6525 l=13775
+ ad=0 pd=0 as=3.57425e+07 ps=26100 
M2454 GND diff_345100_1370250# diff_336400_1363000# GND efet w=7250 l=27550
+ ad=0 pd=0 as=0 ps=0 
M2455 diff_365400_1315150# diff_337850_1312250# GND GND efet w=26825 l=10875
+ ad=7.00132e+08 pd=211700 as=0 ps=0 
M2456 diff_337850_1312250# GND diff_249400_1373150# GND efet w=13050 l=13775
+ ad=1.63995e+08 pd=60900 as=0 ps=0 
M2457 diff_290000_1419550# GND diff_365400_1315150# GND efet w=14500 l=11600
+ ad=1.45072e+08 pd=60900 as=0 ps=0 
M2458 GND GND diff_365400_1315150# GND efet w=8700 l=37700
+ ad=0 pd=0 as=0 ps=0 
M2459 diff_767050_1451450# GND GND GND efet w=14500 l=11600
+ ad=2.6071e+08 pd=95700 as=0 ps=0 
M2460 diff_497350_1464500# diff_661200_1406500# diff_497350_1464500# GND efet w=15950 l=58000
+ ad=0 pd=0 as=0 ps=0 
M2461 diff_249400_1373150# diff_249400_1373150# GND GND efet w=18125 l=17400
+ ad=0 pd=0 as=0 ps=0 
M2462 GND GND diff_249400_1373150# GND efet w=28275 l=19575
+ ad=0 pd=0 as=0 ps=0 
M2463 diff_249400_1373150# diff_291450_1273100# GND GND efet w=36975 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2464 GND diff_345100_1226700# GND GND efet w=75400 l=5800
+ ad=0 pd=0 as=0 ps=0 
M2465 GND diff_291450_1273100# GND GND efet w=26100 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2466 GND GND diff_345100_1226700# GND efet w=5800 l=11600
+ ad=0 pd=0 as=4.6255e+07 ps=29000 
M2467 GND diff_345100_1226700# GND GND efet w=7975 l=26825
+ ad=0 pd=0 as=0 ps=0 
M2468 GND diff_661200_1406500# diff_497350_1464500# GND efet w=5800 l=39875
+ ad=0 pd=0 as=0 ps=0 
M2469 diff_787350_1442750# GND diff_767050_1451450# GND efet w=8700 l=11600
+ ad=5.887e+07 pd=31900 as=0 ps=0 
M2470 GND GND diff_846800_1510900# GND efet w=5800 l=49300
+ ad=0 pd=0 as=0 ps=0 
M2471 GND GND GND GND efet w=19575 l=18125
+ ad=0 pd=0 as=0 ps=0 
M2472 GND GND GND GND efet w=25375 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2473 GND GND GND GND efet w=31175 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2474 GND GND GND GND efet w=20300 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2475 GND GND GND GND efet w=20300 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2476 GND GND GND GND efet w=18850 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2477 GND GND GND GND efet w=20300 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2478 GND GND GND GND efet w=24650 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2479 GND GND GND GND efet w=19575 l=17400
+ ad=0 pd=0 as=0 ps=0 
M2480 diff_1048350_1547150# diff_519100_1629800# GND GND efet w=27550 l=11600
+ ad=5.25625e+08 pd=168200 as=0 ps=0 
M2481 GND diff_797500_1757400# diff_1048350_1547150# GND efet w=49300 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2482 GND diff_1080250_1561650# GND GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2483 GND diff_1080250_1561650# GND GND efet w=42050 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2484 GND diff_1080250_1561650# GND GND efet w=41325 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2485 GND diff_1080250_1561650# GND GND efet w=31175 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2486 GND diff_1080250_1561650# GND GND efet w=30450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2487 GND diff_1080250_1561650# GND GND efet w=31900 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2488 GND diff_1080250_1561650# GND GND efet w=31175 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2489 GND diff_1080250_1561650# GND GND efet w=29725 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2490 GND diff_797500_1757400# GND GND efet w=24650 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2491 GND diff_797500_1757400# diff_1400700_1510900# GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2492 GND diff_797500_1757400# GND GND efet w=26100 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2493 GND GND diff_1080250_1657350# GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2494 GND GND GND GND efet w=68875 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2495 GND diff_797500_1757400# GND GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2496 GND diff_797500_1757400# GND GND efet w=23200 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2497 GND diff_797500_1757400# GND GND efet w=23200 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2498 GND diff_797500_1757400# GND GND efet w=24650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2499 GND diff_797500_1757400# GND GND efet w=24650 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2500 GND GND GND GND efet w=44225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2501 GND diff_1016450_1492050# diff_535050_885950# GND efet w=22475 l=10875
+ ad=0 pd=0 as=2.0228e+08 ps=1.0266e+06 
M2502 diff_535050_885950# GND GND GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2503 GND GND diff_1016450_1492050# GND efet w=14500 l=10150
+ ad=0 pd=0 as=3.09067e+08 ps=127600 
M2504 diff_1194800_1497850# GND GND GND efet w=14500 l=10150
+ ad=-3.65395e+08 pd=1.2383e+06 as=0 ps=0 
M2505 GND GND GND GND efet w=44225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2506 GND GND diff_767050_1451450# GND efet w=5800 l=47850
+ ad=0 pd=0 as=0 ps=0 
M2507 diff_785900_1464500# diff_787350_1442750# GND GND efet w=21750 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2508 GND GND diff_846800_1278900# GND efet w=5800 l=15950
+ ad=0 pd=0 as=1.83548e+09 ps=498800 
M2509 diff_1016450_1492050# GND GND GND efet w=6525 l=64525
+ ad=0 pd=0 as=0 ps=0 
M2510 GND GND diff_1194800_1497850# GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2511 diff_1194800_1497850# GND GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2512 diff_661200_1406500# GND GND GND efet w=5800 l=11600
+ ad=1.19842e+08 pd=55100 as=0 ps=0 
M2513 GND GND GND GND efet w=6525 l=18850
+ ad=0 pd=0 as=0 ps=0 
M2514 diff_846800_1278900# diff_785900_1464500# GND GND efet w=65250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2515 diff_785900_1464500# GND GND GND efet w=5800 l=36250
+ ad=0 pd=0 as=0 ps=0 
M2516 diff_598850_1270200# GND GND GND efet w=5800 l=56550
+ ad=4.85678e+08 pd=188500 as=0 ps=0 
M2517 diff_655400_1313700# GND GND GND efet w=5800 l=29000
+ ad=9.18793e+08 pd=272600 as=0 ps=0 
M2518 GND GND diff_733700_1262950# GND efet w=6525 l=64525
+ ad=0 pd=0 as=9.37715e+08 ps=324800 
M2519 diff_365400_1168700# diff_337850_1168700# GND GND efet w=26825 l=10875
+ ad=6.95927e+08 pd=203000 as=0 ps=0 
M2520 diff_337850_1168700# GND diff_249400_1373150# GND efet w=15950 l=11600
+ ad=1.7661e+08 pd=60900 as=0 ps=0 
M2521 diff_291450_1273100# GND diff_365400_1168700# GND efet w=14500 l=11600
+ ad=1.63995e+08 pd=60900 as=0 ps=0 
M2522 GND GND diff_365400_1168700# GND efet w=7250 l=30450
+ ad=0 pd=0 as=0 ps=0 
M2523 diff_655400_1313700# diff_617700_1270200# GND GND efet w=34800 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2524 GND GND diff_655400_1313700# GND efet w=21750 l=18850
+ ad=0 pd=0 as=0 ps=0 
M2525 GND diff_655400_1313700# GND GND efet w=53650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2526 GND GND diff_733700_1262950# GND efet w=10150 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2527 diff_733700_1262950# GND GND GND efet w=11600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2528 diff_667000_1268750# GND GND GND efet w=29000 l=13050
+ ad=2.1025e+08 pd=72500 as=0 ps=0 
M2529 GND GND diff_667000_1268750# GND efet w=29725 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2530 diff_598850_1270200# diff_249400_1373150# GND GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2531 diff_617700_1270200# GND diff_598850_1270200# GND efet w=9425 l=12325
+ ad=1.15638e+08 pd=52200 as=0 ps=0 
M2532 diff_706150_1268750# GND GND GND efet w=31175 l=12325
+ ad=2.33378e+08 pd=81200 as=0 ps=0 
M2533 diff_725000_1268750# diff_655400_1313700# diff_706150_1268750# GND efet w=31175 l=10875
+ ad=2.45992e+08 pd=75400 as=0 ps=0 
M2534 diff_710500_1136800# diff_733700_1262950# diff_725000_1268750# GND efet w=29725 l=12325
+ ad=1.98266e+09 pd=774300 as=0 ps=0 
M2535 GND GND diff_710500_1136800# GND efet w=27550 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2536 GND GND diff_564050_1106350# GND efet w=21750 l=13050
+ ad=0 pd=0 as=6.11828e+08 ps=165300 
M2537 diff_710500_1136800# GND GND GND efet w=29000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2538 diff_535050_885950# GND GND GND efet w=7250 l=43500
+ ad=0 pd=0 as=0 ps=0 
M2539 GND diff_1077350_1464500# diff_1057050_1325300# GND efet w=15950 l=10150
+ ad=0 pd=0 as=2.523e+08 ps=75400 
M2540 diff_1057050_1325300# GND GND GND efet w=6525 l=58725
+ ad=0 pd=0 as=0 ps=0 
M2541 GND GND GND GND efet w=11600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2542 GND GND diff_1197700_1436950# GND efet w=12325 l=12325
+ ad=0 pd=0 as=1.04074e+09 ps=365400 
M2543 diff_1267300_1444200# GND GND GND efet w=13050 l=11600
+ ad=1.7619e+09 pd=600300 as=0 ps=0 
M2544 GND diff_1141150_1415200# diff_1109250_1280350# GND efet w=76125 l=10875
+ ad=0 pd=0 as=-2.1399e+09 ps=565500 
M2545 GND diff_710500_1136800# GND GND efet w=21025 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2546 GND GND diff_564050_1106350# GND efet w=6525 l=31175
+ ad=0 pd=0 as=0 ps=0 
M2547 GND diff_249400_1373150# diff_249400_1373150# GND efet w=17400 l=18850
+ ad=0 pd=0 as=0 ps=0 
M2548 GND diff_336400_1125200# diff_249400_1373150# GND efet w=40600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2549 diff_249400_1373150# diff_291450_1128100# GND GND efet w=34800 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2550 diff_336400_1125200# diff_345100_1081700# diff_336400_1125200# GND efet w=70325 l=5800
+ ad=1.12694e+09 pd=339300 as=0 ps=0 
M2551 diff_336400_1125200# diff_291450_1128100# GND GND efet w=27550 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2552 GND GND diff_345100_1081700# GND efet w=5800 l=11600
+ ad=0 pd=0 as=6.728e+07 ps=34800 
M2553 GND diff_345100_1081700# diff_336400_1125200# GND efet w=4350 l=31175
+ ad=0 pd=0 as=0 ps=0 
M2554 GND GND diff_577100_1051250# GND efet w=5800 l=49300
+ ad=0 pd=0 as=6.3075e+08 ps=208800 
M2555 diff_709050_1219450# GND diff_709050_1219450# GND efet w=4350 l=75400
+ ad=4.14193e+08 pd=127600 as=0 ps=0 
M2556 diff_577100_1051250# diff_564050_1106350# diff_546650_1088950# GND efet w=10150 l=10875
+ ad=0 pd=0 as=5.887e+07 ps=40600 
M2557 diff_365400_1023700# diff_339300_1022250# GND GND efet w=26825 l=10875
+ ad=6.79108e+08 pd=211700 as=0 ps=0 
M2558 diff_339300_1022250# GND GND GND efet w=13775 l=15225
+ ad=1.61892e+08 pd=58000 as=0 ps=0 
M2559 diff_291450_1128100# GND diff_365400_1023700# GND efet w=14500 l=11600
+ ad=1.5979e+08 pd=66700 as=0 ps=0 
M2560 GND GND diff_582900_1045450# GND efet w=8700 l=12325
+ ad=0 pd=0 as=6.3075e+07 ps=37700 
M2561 GND diff_709050_1219450# GND GND efet w=20300 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2562 GND diff_710500_1136800# diff_709050_1219450# GND efet w=11600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2563 GND diff_713400_1139700# diff_710500_1136800# GND efet w=6525 l=52925
+ ad=0 pd=0 as=0 ps=0 
M2564 diff_713400_1139700# GND GND GND efet w=6525 l=12325
+ ad=1.38765e+08 pd=63800 as=0 ps=0 
M2565 diff_710500_1136800# diff_713400_1139700# diff_710500_1136800# GND efet w=70325 l=5075
+ ad=0 pd=0 as=0 ps=0 
M2566 GND GND diff_552450_1347050# GND efet w=11600 l=54375
+ ad=0 pd=0 as=-4.01137e+08 ps=988900 
M2567 GND GND GND GND efet w=3625 l=71775
+ ad=0 pd=0 as=0 ps=0 
M2568 diff_249400_1373150# GND diff_803300_1059950# GND efet w=7975 l=13050
+ ad=0 pd=0 as=1.38765e+08 ps=55100 
M2569 diff_751100_1103450# GND GND GND efet w=5800 l=56550
+ ad=7.77925e+08 pd=208800 as=0 ps=0 
M2570 diff_751100_1103450# diff_564050_1106350# GND GND efet w=10875 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2571 GND GND diff_552450_1347050# GND efet w=26825 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2572 GND diff_249400_1373150# GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2573 GND diff_582900_1045450# diff_577100_1051250# GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2574 GND diff_803300_1059950# diff_751100_1103450# GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2575 diff_526350_1077350# GND GND GND efet w=6525 l=51475
+ ad=1.34981e+09 pd=406000 as=0 ps=0 
M2576 GND GND diff_365400_1023700# GND efet w=7975 l=38425
+ ad=0 pd=0 as=0 ps=0 
M2577 GND diff_546650_1088950# diff_526350_1077350# GND efet w=23925 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2578 diff_249400_1373150# GND GND GND efet w=21750 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2579 GND GND GND GND efet w=34800 l=26100
+ ad=0 pd=0 as=0 ps=0 
M2580 GND diff_681500_959900# GND GND efet w=24650 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2581 GND diff_291450_967150# GND GND efet w=38425 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2582 GND diff_495900_936700# GND GND efet w=65975 l=7250
+ ad=0 pd=0 as=0 ps=0 
M2583 GND GND GND GND efet w=70325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2584 GND diff_495900_936700# GND GND efet w=10150 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2585 GND diff_345100_925100# GND GND efet w=78300 l=8700
+ ad=0 pd=0 as=0 ps=0 
M2586 GND diff_754000_974400# GND GND efet w=21750 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2587 GND GND diff_1109250_1280350# GND efet w=73950 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2588 GND diff_1181750_1322400# diff_1194800_1497850# GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2589 diff_1194800_1497850# GND GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2590 diff_1305000_1400700# diff_1077350_1464500# GND GND efet w=11600 l=12325
+ ad=6.11828e+08 pd=194300 as=0 ps=0 
M2591 GND GND GND GND efet w=14500 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2592 GND GND diff_1194800_1497850# GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2593 diff_1194800_1497850# GND GND GND efet w=13775 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2594 GND GND diff_1194800_1497850# GND efet w=11600 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2595 diff_1194800_1497850# GND GND GND efet w=11600 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2596 GND diff_2150350_1422450# diff_1232500_1610950# GND efet w=34075 l=15225
+ ad=0 pd=0 as=6.5598e+08 ps=205900 
M2597 diff_1194800_1497850# GND GND GND efet w=12325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2598 GND GND diff_1232500_1610950# GND efet w=30450 l=26100
+ ad=0 pd=0 as=0 ps=0 
M2599 GND diff_2150350_1422450# GND GND efet w=26825 l=16675
+ ad=0 pd=0 as=0 ps=0 
M2600 GND GND diff_1194800_1497850# GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2601 diff_1194800_1497850# GND GND GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2602 GND GND diff_1194800_1497850# GND efet w=13775 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2603 diff_1194800_1497850# GND GND GND efet w=13775 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2604 GND GND GND GND efet w=16675 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2605 GND GND GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2606 GND GND GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2607 GND GND GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2608 GND GND GND GND efet w=13775 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2609 GND GND GND GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2610 GND GND GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2611 GND GND GND GND efet w=13775 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2612 GND GND GND GND efet w=13050 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2613 GND GND GND GND efet w=13775 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2614 GND diff_1400700_1510900# diff_1267300_1444200# GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2615 diff_1267300_1444200# GND GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2616 diff_1109250_1280350# diff_1141150_1351400# diff_1087500_571300# GND efet w=74675 l=10875
+ ad=0 pd=0 as=-1.88785e+08 ps=951200 
M2617 diff_1087500_571300# diff_846800_1278900# diff_1109250_1280350# GND efet w=76125 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2618 GND diff_1057050_1325300# diff_1055600_1228150# GND efet w=39150 l=12325
+ ad=0 pd=0 as=-1.42295e+09 ps=791700 
M2619 GND diff_1181750_1322400# diff_1141150_1351400# GND efet w=21750 l=11600
+ ad=0 pd=0 as=2.79633e+08 ps=116000 
M2620 GND diff_1141150_1415200# diff_1177400_1117950# GND efet w=14500 l=11600
+ ad=0 pd=0 as=6.28647e+08 ps=171100 
M2621 GND diff_1286150_1331100# diff_1141150_1415200# GND efet w=21750 l=11600
+ ad=0 pd=0 as=4.73062e+08 ps=162400 
M2622 diff_1197700_1436950# GND GND GND efet w=13050 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2623 diff_1267300_1444200# GND GND GND efet w=12325 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2624 GND GND diff_1267300_1444200# GND efet w=12325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2625 GND GND diff_1267300_1444200# GND efet w=11600 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2626 GND diff_1592100_1387650# GND GND efet w=65250 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2627 GND GND diff_1305000_1400700# GND efet w=11600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2628 diff_1349950_1289050# GND GND GND efet w=15225 l=10875
+ ad=4.4573e+08 pd=150800 as=0 ps=0 
M2629 diff_1177400_1117950# diff_846800_1278900# GND GND efet w=15950 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2630 GND GND GND GND efet w=23925 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2631 GND diff_1592100_1387650# GND GND efet w=5800 l=40600
+ ad=0 pd=0 as=0 ps=0 
M2632 diff_1305000_1400700# GND GND GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2633 diff_1305000_1400700# GND GND GND efet w=7250 l=66700
+ ad=0 pd=0 as=0 ps=0 
M2634 diff_1267300_1444200# GND GND GND efet w=7250 l=69600
+ ad=0 pd=0 as=0 ps=0 
M2635 GND diff_1400700_1510900# diff_1419550_1315150# GND efet w=15225 l=15225
+ ad=0 pd=0 as=5.42445e+08 ps=188500 
M2636 GND diff_846800_1278900# diff_1332550_1297750# GND efet w=17400 l=10875
+ ad=0 pd=0 as=6.60185e+08 ps=188500 
M2637 GND diff_846800_1278900# diff_1055600_1228150# GND efet w=38425 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2638 diff_1055600_1228150# diff_1048350_1142600# diff_1055600_1228150# GND efet w=84100 l=28275
+ ad=0 pd=0 as=0 ps=0 
M2639 diff_1055600_1228150# diff_1048350_1142600# GND GND efet w=8700 l=24650
+ ad=0 pd=0 as=0 ps=0 
M2640 diff_1087500_571300# diff_1113600_1132450# diff_1087500_571300# GND efet w=74675 l=50025
+ ad=0 pd=0 as=0 ps=0 
M2641 diff_1141150_1351400# GND diff_1141150_1351400# GND efet w=3625 l=46400
+ ad=0 pd=0 as=0 ps=0 
M2642 GND diff_1349950_1289050# diff_1332550_1297750# GND efet w=13050 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2643 diff_1177400_1117950# GND GND GND efet w=5800 l=72500
+ ad=0 pd=0 as=0 ps=0 
M2644 diff_1141150_1415200# GND GND GND efet w=8700 l=43500
+ ad=0 pd=0 as=0 ps=0 
M2645 GND diff_846800_1278900# diff_1426800_1106350# GND efet w=14500 l=11600
+ ad=0 pd=0 as=-1.95068e+09 ps=638000 
M2646 diff_1426800_1106350# diff_1419550_1315150# GND GND efet w=15950 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2647 GND GND diff_1525400_1289050# GND efet w=11600 l=11600
+ ad=0 pd=0 as=1.57688e+08 ps=78300 
M2648 GND GND diff_1592100_1387650# GND efet w=6525 l=13775
+ ad=0 pd=0 as=1.5979e+08 ps=66700 
M2649 diff_1087500_571300# diff_1113600_1132450# GND GND efet w=10875 l=29725
+ ad=0 pd=0 as=0 ps=0 
M2650 GND GND diff_1332550_1297750# GND efet w=8700 l=65250
+ ad=0 pd=0 as=0 ps=0 
M2651 diff_1349950_1289050# GND GND GND efet w=5800 l=60900
+ ad=0 pd=0 as=0 ps=0 
M2652 GND GND diff_1419550_1315150# GND efet w=7975 l=84825
+ ad=0 pd=0 as=0 ps=0 
M2653 diff_1426800_1106350# GND GND GND efet w=7250 l=65250
+ ad=0 pd=0 as=0 ps=0 
M2654 diff_1547150_726450# diff_1525400_1289050# GND GND efet w=13775 l=11600
+ ad=-2.1399e+09 pd=748200 as=0 ps=0 
M2655 GND GND diff_1547150_726450# GND efet w=13050 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2656 GND GND GND GND efet w=6525 l=63800
+ ad=0 pd=0 as=0 ps=0 
M2657 diff_1525400_1289050# GND diff_1525400_1289050# GND efet w=3625 l=87725
+ ad=0 pd=0 as=0 ps=0 
M2658 GND GND diff_1197700_311750# GND efet w=19575 l=13775
+ ad=0 pd=0 as=2.08989e+09 ps=696000 
M2659 diff_1267300_1444200# GND GND GND efet w=13050 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2660 diff_1197700_1436950# GND GND GND efet w=12325 l=16675
+ ad=0 pd=0 as=0 ps=0 
M2661 GND GND GND GND efet w=21750 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2662 diff_1197700_1436950# GND diff_1197700_1436950# GND efet w=2900 l=63800
+ ad=0 pd=0 as=0 ps=0 
M2663 GND GND GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2664 diff_1267300_1444200# GND GND GND efet w=13050 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2665 GND GND diff_1194800_1497850# GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2666 GND GND diff_1267300_1444200# GND efet w=13775 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2667 GND GND diff_1197700_1436950# GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2668 GND GND GND GND efet w=17400 l=17400
+ ad=0 pd=0 as=0 ps=0 
M2669 diff_2085100_1422450# GND diff_2085100_1422450# GND efet w=5800 l=44950
+ ad=5.8029e+08 pd=171100 as=0 ps=0 
M2670 GND diff_2215600_1422450# GND GND efet w=32625 l=25375
+ ad=0 pd=0 as=0 ps=0 
M2671 diff_2085100_1422450# GND GND GND efet w=25375 l=16675
+ ad=0 pd=0 as=0 ps=0 
M2672 GND GND diff_2150350_1422450# GND efet w=7975 l=38425
+ ad=0 pd=0 as=5.57162e+08 ps=162400 
M2673 GND diff_1999550_1331100# GND GND efet w=58725 l=18125
+ ad=0 pd=0 as=0 ps=0 
M2674 GND GND diff_1624000_314650# GND efet w=54375 l=12325
+ ad=0 pd=0 as=-1.58274e+09 ps=823600 
M2675 diff_1624000_314650# diff_2654950_1667500# diff_1624000_314650# GND efet w=65250 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2676 diff_2654950_1667500# GND GND GND efet w=8700 l=15950
+ ad=5.4665e+07 pd=34800 as=0 ps=0 
M2677 GND GND diff_2578100_1628350# GND efet w=13050 l=33350
+ ad=0 pd=0 as=1.47175e+09 ps=292900 
M2678 GND diff_1999550_1331100# diff_797500_1757400# GND efet w=65250 l=13050
+ ad=0 pd=0 as=-1.42295e+09 ps=646700 
M2679 GND diff_2280850_1441300# diff_1080250_1561650# GND efet w=37700 l=14500
+ ad=0 pd=0 as=-1.78458e+09 ps=652500 
M2680 diff_797500_1757400# diff_2269250_1429700# GND GND efet w=70325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2681 diff_1624000_314650# diff_2654950_1667500# GND GND efet w=13050 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2682 diff_2578100_1628350# diff_1624000_314650# GND GND efet w=27550 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2683 diff_2578100_1628350# GND GND GND efet w=48575 l=18125
+ ad=0 pd=0 as=0 ps=0 
M2684 GND diff_2269250_1429700# diff_1080250_1561650# GND efet w=52925 l=25375
+ ad=0 pd=0 as=0 ps=0 
M2685 diff_797500_1757400# diff_2280850_1441300# GND GND efet w=29000 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2686 GND GND diff_2215600_1422450# GND efet w=7250 l=40600
+ ad=0 pd=0 as=6.2234e+08 ps=191400 
M2687 diff_2150350_1422450# GND GND GND efet w=21750 l=19575
+ ad=0 pd=0 as=0 ps=0 
M2688 GND diff_2108300_1347050# GND GND efet w=56550 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2689 GND diff_2173550_1360100# GND GND efet w=55825 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2690 GND GND diff_1999550_1331100# GND efet w=15225 l=12325
+ ad=0 pd=0 as=1.58949e+09 ps=464000 
M2691 diff_2215600_1422450# GND GND GND efet w=21025 l=20300
+ ad=0 pd=0 as=0 ps=0 
M2692 GND GND diff_2280850_1441300# GND efet w=9425 l=35525
+ ad=0 pd=0 as=4.7937e+08 ps=147900 
M2693 diff_2280850_1441300# diff_2269250_1429700# GND GND efet w=34800 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2694 GND diff_2238800_1378950# GND GND efet w=57275 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2695 GND diff_2324350_1402150# diff_2269250_1429700# GND efet w=64525 l=12325
+ ad=0 pd=0 as=4.7937e+08 ps=229100 
M2696 GND GND GND GND efet w=8700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2697 diff_2637550_1542800# GND GND GND efet w=8700 l=17400
+ ad=5.4665e+07 pd=43500 as=0 ps=0 
M2698 GND diff_2637550_1542800# GND GND efet w=68875 l=7250
+ ad=0 pd=0 as=0 ps=0 
M2699 GND diff_2637550_1542800# GND GND efet w=10150 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2700 GND GND GND GND efet w=10150 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2701 GND GND GND GND efet w=49300 l=39875
+ ad=0 pd=0 as=0 ps=0 
M2702 GND GND GND GND efet w=42050 l=23200
+ ad=0 pd=0 as=0 ps=0 
M2703 GND GND GND GND efet w=250850 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2704 GND GND GND GND efet w=227650 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2705 GND GND GND GND efet w=72500 l=37700
+ ad=0 pd=0 as=0 ps=0 
M2706 GND GND GND GND efet w=58000 l=22475
+ ad=0 pd=0 as=0 ps=0 
M2707 GND diff_2282300_2737600# diff_2324350_1402150# GND efet w=10150 l=13050
+ ad=0 pd=0 as=6.51775e+07 ps=40600 
M2708 GND GND GND GND efet w=47125 l=16675
+ ad=0 pd=0 as=0 ps=0 
M2709 GND GND GND GND efet w=19575 l=42050
+ ad=0 pd=0 as=0 ps=0 
M2710 diff_1999550_1331100# GND GND GND efet w=10875 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2711 diff_1194800_1497850# GND diff_1194800_1497850# GND efet w=3625 l=74675
+ ad=0 pd=0 as=0 ps=0 
M2712 GND GND GND GND efet w=11600 l=30450
+ ad=0 pd=0 as=0 ps=0 
M2713 GND GND GND GND efet w=12325 l=49300
+ ad=0 pd=0 as=0 ps=0 
M2714 diff_2269250_1429700# GND GND GND efet w=9425 l=51475
+ ad=0 pd=0 as=0 ps=0 
M2715 GND diff_2282300_2737600# diff_2238800_1378950# GND efet w=10875 l=13775
+ ad=0 pd=0 as=5.4665e+07 ps=40600 
M2716 GND GND GND GND efet w=1227425 l=25375
+ ad=0 pd=0 as=0 ps=0 
M2717 GND diff_1999550_1331100# diff_1999550_1331100# GND efet w=39150 l=18850
+ ad=0 pd=0 as=0 ps=0 
M2718 GND GND diff_1999550_1331100# GND efet w=7250 l=69600
+ ad=0 pd=0 as=0 ps=0 
M2719 diff_1999550_1331100# GND GND GND efet w=36975 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2720 GND diff_2282300_2737600# diff_2173550_1360100# GND efet w=10875 l=13775
+ ad=0 pd=0 as=5.67675e+07 ps=40600 
M2721 GND GND GND GND efet w=657575 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2722 diff_1999550_1331100# diff_2096700_1296300# diff_1999550_1331100# GND efet w=37700 l=47850
+ ad=0 pd=0 as=0 ps=0 
M2723 GND diff_2282300_2737600# diff_2108300_1347050# GND efet w=10150 l=11600
+ ad=0 pd=0 as=6.93825e+07 ps=40600 
M2724 GND diff_2096700_1296300# diff_1999550_1331100# GND efet w=8700 l=20300
+ ad=0 pd=0 as=0 ps=0 
M2725 GND GND GND GND efet w=46400 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2726 GND GND GND GND efet w=39875 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2727 GND GND diff_2096700_1296300# GND efet w=7250 l=11600
+ ad=0 pd=0 as=5.25625e+07 ps=29000 
M2728 GND GND GND GND efet w=7975 l=36250
+ ad=0 pd=0 as=0 ps=0 
M2729 GND GND GND GND efet w=11600 l=21025
+ ad=0 pd=0 as=0 ps=0 
M2730 GND GND GND GND efet w=53650 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2731 GND GND diff_2105400_1174500# GND efet w=11600 l=37700
+ ad=0 pd=0 as=6.9803e+08 ps=165300 
M2732 GND diff_1305000_1400700# diff_2002450_1074450# GND efet w=11600 l=12325
+ ad=0 pd=0 as=3.65835e+08 ps=87000 
M2733 diff_2206900_1222350# GND GND GND efet w=7250 l=20300
+ ad=1.50119e+09 pd=440800 as=0 ps=0 
M2734 GND diff_2161950_1146950# diff_2338850_1251350# GND efet w=57275 l=15225
+ ad=0 pd=0 as=3.55322e+08 ps=118900 
M2735 GND diff_2161950_1146950# diff_2206900_1222350# GND efet w=42775 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2736 GND GND diff_2002450_1074450# GND efet w=13050 l=87000
+ ad=0 pd=0 as=0 ps=0 
M2737 diff_2002450_1074450# GND GND GND efet w=12325 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2738 GND GND diff_1612400_1041100# GND efet w=14500 l=11600
+ ad=0 pd=0 as=1.14166e+09 ps=336400 
M2739 GND diff_1197700_1436950# diff_1592100_1117950# GND efet w=11600 l=10875
+ ad=0 pd=0 as=9.90278e+08 ps=400200 
M2740 GND GND diff_2077850_1148400# GND efet w=8700 l=34075
+ ad=0 pd=0 as=3.63733e+08 ps=95700 
M2741 GND GND diff_2206900_1222350# GND efet w=21025 l=18850
+ ad=0 pd=0 as=0 ps=0 
M2742 diff_667000_980200# diff_1426800_1106350# diff_1426800_1106350# GND efet w=10150 l=15950
+ ad=-1.71686e+09 pd=1.8676e+06 as=0 ps=0 
M2743 diff_1048350_1142600# GND GND GND efet w=5800 l=11600
+ ad=5.887e+07 pd=31900 as=0 ps=0 
M2744 diff_1113600_1132450# GND diff_1113600_1132450# GND efet w=2900 l=18850
+ ad=5.887e+07 pd=31900 as=0 ps=0 
M2745 diff_1284700_1093300# GND diff_1238300_1142600# GND efet w=15950 l=10150
+ ad=1.57057e+09 pd=466900 as=3.67938e+08 ps=107300 
M2746 diff_1238300_1142600# GND GND GND efet w=9425 l=17400
+ ad=0 pd=0 as=0 ps=0 
M2747 diff_1612400_1041100# diff_1726950_1144050# diff_1612400_1041100# GND efet w=60175 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2748 diff_1284700_1093300# GND diff_1262950_1112150# GND efet w=7975 l=12325
+ ad=0 pd=0 as=-1.31993e+09 ps=800400 
M2749 diff_1603700_1123750# diff_1592100_1117950# diff_1262950_1112150# GND efet w=14500 l=11600
+ ad=7.12748e+08 pd=226200 as=0 ps=0 
M2750 diff_1262950_1112150# GND GND GND efet w=10150 l=34800
+ ad=0 pd=0 as=0 ps=0 
M2751 diff_1262950_1112150# GND GND GND efet w=37700 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2752 diff_1426800_1106350# diff_1332550_1297750# diff_1284700_1093300# GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2753 GND diff_1177400_1117950# diff_667000_980200# GND efet w=57275 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2754 GND GND diff_1612400_1041100# GND efet w=13775 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2755 diff_1592100_1117950# diff_1786400_1088950# diff_1592100_1117950# GND efet w=79750 l=20300
+ ad=0 pd=0 as=0 ps=0 
M2756 diff_1448550_1090400# diff_1436950_1083150# diff_1284700_1093300# GND efet w=10150 l=13050
+ ad=1.48857e+09 pd=319000 as=0 ps=0 
M2757 GND diff_1284700_1093300# GND GND efet w=59450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2758 GND GND GND GND efet w=10150 l=33350
+ ad=0 pd=0 as=0 ps=0 
M2759 diff_1090400_903350# diff_1426800_1106350# diff_1284700_1093300# GND efet w=7250 l=11600
+ ad=5.01275e+08 pd=2.1054e+06 as=0 ps=0 
M2760 diff_1612400_1041100# diff_1726950_1144050# GND GND efet w=6525 l=48575
+ ad=0 pd=0 as=0 ps=0 
M2761 GND GND diff_1592100_1117950# GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2762 GND diff_1267300_1444200# diff_1590650_513300# GND efet w=14500 l=11600
+ ad=0 pd=0 as=1.45913e+09 ps=510400 
M2763 GND GND diff_1590650_513300# GND efet w=15225 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2764 GND GND diff_1436950_1083150# GND efet w=13775 l=10875
+ ad=0 pd=0 as=5.36138e+08 ps=110200 
M2765 diff_1194800_1497850# diff_1194800_1497850# GND GND efet w=11600 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2766 diff_2105400_1174500# GND GND GND efet w=22475 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2767 GND GND diff_2338850_1251350# GND efet w=43500 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2768 GND diff_2105400_1174500# diff_2077850_1148400# GND efet w=29000 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2769 GND diff_2130050_1220900# diff_2105400_1174500# GND efet w=24650 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2770 diff_2206900_1222350# diff_1624000_314650# diff_2130050_1220900# GND efet w=10150 l=11600
+ ad=0 pd=0 as=2.06045e+08 ps=92800 
M2771 diff_1352850_295800# diff_2077850_1148400# GND GND efet w=41325 l=14500
+ ad=4.16735e+08 pd=954100 as=0 ps=0 
M2772 diff_2105400_1174500# GND GND GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2773 GND diff_2105400_1174500# diff_1352850_295800# GND efet w=45675 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2774 GND diff_1925600_1133900# diff_1436950_1083150# GND efet w=13050 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2775 GND diff_1925600_1133900# diff_1194800_1497850# GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2776 GND GND diff_1194800_1497850# GND efet w=5800 l=69600
+ ad=0 pd=0 as=0 ps=0 
M2777 GND diff_1786400_1088950# diff_1592100_1117950# GND efet w=5800 l=58000
+ ad=0 pd=0 as=0 ps=0 
M2778 diff_1436950_1083150# GND GND GND efet w=8700 l=79750
+ ad=0 pd=0 as=0 ps=0 
M2779 diff_1786400_1088950# GND GND GND efet w=7250 l=11600
+ ad=1.28252e+08 pd=63800 as=0 ps=0 
M2780 diff_1726950_1144050# GND GND GND efet w=7975 l=10150
+ ad=6.09725e+07 pd=37700 as=0 ps=0 
M2781 diff_2161950_1146950# GND diff_2243150_1175950# GND efet w=10875 l=13050
+ ad=0 pd=0 as=8.41e+07 ps=40600 
M2782 GND GND diff_2344650_1202050# GND efet w=44950 l=15950
+ ad=0 pd=0 as=4.31013e+08 ps=130500 
M2783 diff_2344650_1202050# GND GND GND efet w=49300 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2784 GND diff_2243150_1175950# GND GND efet w=59450 l=9425
+ ad=0 pd=0 as=0 ps=0 
M2785 GND diff_2161950_1146950# diff_2153250_1116500# GND efet w=126150 l=13050
+ ad=0 pd=0 as=9.62945e+08 ps=272600 
M2786 GND GND GND GND efet w=55825 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2787 diff_2153250_1116500# diff_1624000_314650# GND GND efet w=96425 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2788 GND GND GND GND efet w=15225 l=27550
+ ad=0 pd=0 as=0 ps=0 
M2789 GND GND diff_2272150_1090400# GND efet w=37700 l=15950
+ ad=0 pd=0 as=4.09987e+08 ps=150800 
M2790 GND GND diff_1603700_1123750# GND efet w=10150 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2791 diff_1603700_1123750# diff_2002450_1074450# GND GND efet w=9425 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2792 GND diff_1168700_1032400# diff_667000_980200# GND efet w=53650 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2793 diff_667000_980200# GND GND GND efet w=6525 l=29000
+ ad=0 pd=0 as=0 ps=0 
M2794 GND diff_1197700_311750# diff_1168700_1032400# GND efet w=8700 l=10150
+ ad=0 pd=0 as=4.68858e+08 ps=156600 
M2795 diff_1603700_1123750# diff_1612400_1041100# GND GND efet w=15950 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2796 GND GND diff_2122800_433550# GND efet w=13050 l=11600
+ ad=0 pd=0 as=1.49067e+09 ps=452400 
M2797 diff_2122800_433550# GND GND GND efet w=18125 l=9425
+ ad=0 pd=0 as=0 ps=0 
M2798 diff_2272150_1090400# GND GND GND efet w=9425 l=38425
+ ad=0 pd=0 as=0 ps=0 
M2799 GND diff_2272150_1090400# GND GND efet w=65975 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2800 GND GND GND GND efet w=13775 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2801 diff_1842950_996150# diff_1603700_1123750# diff_1824100_994700# GND efet w=59450 l=11600
+ ad=5.44548e+08 pd=179800 as=3.6163e+08 ps=124700 
M2802 GND diff_1603700_1123750# diff_1850200_999050# GND efet w=61625 l=10875
+ ad=0 pd=0 as=-1.57643e+09 ps=693100 
M2803 GND diff_1745800_945400# diff_1090400_903350# GND efet w=60900 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2804 GND GND GND GND efet w=7250 l=50750
+ ad=0 pd=0 as=0 ps=0 
M2805 GND diff_1160000_1010650# GND GND efet w=58725 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2806 diff_1290500_990350# diff_1197700_311750# diff_1160000_1010650# GND efet w=7975 l=12325
+ ad=-1.06763e+09 pd=733700 as=3.9527e+08 ps=127600 
M2807 GND GND GND GND efet w=6525 l=32625
+ ad=0 pd=0 as=0 ps=0 
M2808 GND diff_1547150_726450# diff_1290500_990350# GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2809 diff_1090400_903350# diff_1731300_991800# GND GND efet w=13050 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2810 diff_1824100_994700# GND GND GND efet w=44225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2811 GND diff_667000_980200# diff_681500_959900# GND efet w=14500 l=17400
+ ad=0 pd=0 as=5.61367e+08 ps=188500 
M2812 GND diff_291450_967150# GND GND efet w=29000 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2813 GND GND diff_345100_925100# GND efet w=6525 l=11600
+ ad=0 pd=0 as=6.728e+07 ps=34800 
M2814 diff_495900_936700# GND GND GND efet w=8700 l=13050
+ ad=6.51775e+07 pd=34800 as=0 ps=0 
M2815 GND GND GND GND efet w=77575 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2816 GND diff_345100_925100# GND GND efet w=5800 l=27550
+ ad=0 pd=0 as=0 ps=0 
M2817 diff_291450_967150# GND diff_365400_861300# GND efet w=15950 l=10150
+ ad=1.5138e+08 pd=63800 as=7.21158e+08 ps=214600 
M2818 diff_365400_861300# diff_339300_859850# GND GND efet w=27550 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2819 diff_339300_859850# GND diff_136300_2602750# GND efet w=14500 l=11600
+ ad=1.57688e+08 pd=58000 as=-1.77275e+09 ps=3.6801e+06 
M2820 GND GND diff_365400_861300# GND efet w=8700 l=40600
+ ad=0 pd=0 as=0 ps=0 
M2821 diff_249400_1373150# diff_136300_2602750# GND GND efet w=23200 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2822 GND GND diff_754000_974400# GND efet w=13050 l=11600
+ ad=0 pd=0 as=2.6071e+08 ps=75400 
M2823 diff_849700_965700# diff_681500_959900# GND GND efet w=28275 l=11600
+ ad=2.1025e+08 pd=72500 as=0 ps=0 
M2824 GND GND diff_849700_965700# GND efet w=29000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2825 GND GND GND GND efet w=10875 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2826 GND GND GND GND efet w=17400 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2827 diff_1290500_990350# GND GND GND efet w=10150 l=37700
+ ad=0 pd=0 as=0 ps=0 
M2828 diff_681500_959900# GND diff_681500_891750# GND efet w=28275 l=10150
+ ad=0 pd=0 as=1.24888e+09 ps=365400 
M2829 GND diff_337850_765600# diff_136300_2602750# GND efet w=38425 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2830 diff_136300_2602750# diff_291450_822150# GND GND efet w=39150 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2831 diff_337850_765600# diff_346550_772850# diff_337850_765600# GND efet w=68150 l=6525
+ ad=1.1753e+09 pd=348000 as=0 ps=0 
M2832 diff_337850_765600# diff_291450_822150# GND GND efet w=34800 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2833 GND GND diff_346550_772850# GND efet w=5800 l=13050
+ ad=0 pd=0 as=7.1485e+07 ps=37700 
M2834 GND diff_346550_772850# diff_337850_765600# GND efet w=7250 l=26100
+ ad=0 pd=0 as=0 ps=0 
M2835 GND GND diff_535050_885950# GND efet w=8700 l=43500
+ ad=0 pd=0 as=0 ps=0 
M2836 GND GND GND GND efet w=7975 l=45675
+ ad=0 pd=0 as=0 ps=0 
M2837 GND GND GND GND efet w=7250 l=44950
+ ad=0 pd=0 as=0 ps=0 
M2838 GND GND diff_681500_891750# GND efet w=33350 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2839 diff_681500_891750# GND GND GND efet w=37700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2840 diff_681500_959900# GND GND GND efet w=3625 l=52925
+ ad=0 pd=0 as=0 ps=0 
M2841 GND GND GND GND efet w=5800 l=34075
+ ad=0 pd=0 as=0 ps=0 
M2842 diff_754000_974400# GND GND GND efet w=5800 l=71050
+ ad=0 pd=0 as=0 ps=0 
M2843 GND GND GND GND efet w=6525 l=47125
+ ad=0 pd=0 as=0 ps=0 
M2844 GND GND GND GND efet w=8700 l=50750
+ ad=0 pd=0 as=0 ps=0 
M2845 GND GND GND GND efet w=5075 l=45675
+ ad=0 pd=0 as=0 ps=0 
M2846 GND GND diff_717750_555350# GND efet w=7975 l=51475
+ ad=0 pd=0 as=-2.11467e+09 ps=519100 
M2847 GND GND GND GND efet w=3625 l=51475
+ ad=0 pd=0 as=0 ps=0 
M2848 GND GND GND GND efet w=26825 l=19575
+ ad=0 pd=0 as=0 ps=0 
M2849 GND GND diff_925100_1455800# GND efet w=21750 l=11600
+ ad=0 pd=0 as=2.0163e+09 ps=458200 
M2850 diff_667000_980200# diff_1332550_1297750# GND GND efet w=7250 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2851 GND GND diff_1290500_990350# GND efet w=50750 l=22475
+ ad=0 pd=0 as=0 ps=0 
M2852 GND GND GND GND efet w=13050 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2853 diff_1262950_939600# GND GND GND efet w=9425 l=36975
+ ad=-1.3788e+09 pd=730800 as=0 ps=0 
M2854 GND diff_1087500_571300# GND GND efet w=43500 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2855 diff_925100_1455800# GND GND GND efet w=8700 l=44950
+ ad=0 pd=0 as=0 ps=0 
M2856 GND diff_1090400_903350# diff_871450_1602250# GND efet w=42775 l=10875
+ ad=0 pd=0 as=1.67149e+09 ps=449500 
M2857 GND GND diff_1262950_939600# GND efet w=7250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2858 diff_1090400_903350# diff_1194800_1497850# GND GND efet w=10150 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2859 GND diff_1745800_945400# diff_1731300_991800# GND efet w=12325 l=13775
+ ad=0 pd=0 as=2.6071e+08 ps=81200 
M2860 diff_1745800_945400# diff_1850200_999050# diff_1842950_996150# GND efet w=60900 l=12325
+ ad=9.251e+08 pd=284200 as=0 ps=0 
M2861 GND GND GND GND efet w=60175 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2862 diff_1850200_999050# diff_1850200_999050# GND GND efet w=46400 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2863 GND diff_1290500_990350# diff_1262950_939600# GND efet w=36250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2864 diff_1731300_991800# GND GND GND efet w=5800 l=59450
+ ad=0 pd=0 as=0 ps=0 
M2865 diff_1850200_999050# GND diff_1925600_946850# GND efet w=68875 l=17400
+ ad=0 pd=0 as=7.10645e+08 ps=205900 
M2866 diff_1925600_946850# diff_1850200_999050# GND GND efet w=55825 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2867 diff_2148900_1010650# diff_2209800_997600# GND GND efet w=22475 l=12325
+ ad=8.55718e+08 pd=226200 as=0 ps=0 
M2868 GND GND GND GND efet w=93525 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2869 diff_2148900_1010650# diff_2122800_433550# diff_1850200_999050# GND efet w=13775 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2870 GND diff_2144550_958450# diff_2148900_1010650# GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2871 GND GND diff_1925600_946850# GND efet w=5800 l=66700
+ ad=0 pd=0 as=0 ps=0 
M2872 diff_1090400_862750# diff_1426800_1106350# GND GND efet w=10150 l=11600
+ ad=-3.12392e+08 pd=1.9111e+06 as=0 ps=0 
M2873 diff_1745800_945400# GND GND GND efet w=7250 l=53650
+ ad=0 pd=0 as=0 ps=0 
M2874 diff_1798000_938150# diff_1784950_914950# diff_1745800_945400# GND efet w=36250 l=13050
+ ad=8.55718e+08 pd=229100 as=0 ps=0 
M2875 GND GND diff_1798000_938150# GND efet w=35525 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2876 diff_1798000_938150# diff_1603700_1123750# GND GND efet w=43500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2877 GND diff_1850200_999050# diff_1798000_938150# GND efet w=35525 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2878 diff_1996650_962800# diff_1925600_946850# GND GND efet w=11600 l=11600
+ ad=2.08148e+08 pd=92800 as=0 ps=0 
M2879 GND GND diff_1996650_962800# GND efet w=7250 l=63075
+ ad=0 pd=0 as=0 ps=0 
M2880 GND diff_1055600_1228150# diff_1090400_903350# GND efet w=40600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2881 GND diff_1590650_513300# diff_1262950_939600# GND efet w=14500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2882 diff_2209800_997600# GND GND GND efet w=4350 l=47850
+ ad=2.16558e+08 pd=104400 as=0 ps=0 
M2883 GND diff_2144550_958450# diff_2209800_997600# GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2884 diff_2144550_958450# GND diff_1850200_999050# GND efet w=15225 l=12325
+ ad=2.00578e+09 pd=574200 as=0 ps=0 
M2885 diff_2144550_958450# diff_2209800_997600# GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2886 GND diff_2144550_958450# diff_2144550_958450# GND efet w=18850 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2887 GND GND diff_2275050_913500# GND efet w=7250 l=11600
+ ad=0 pd=0 as=3.67938e+08 ps=113100 
M2888 diff_1784950_914950# diff_1996650_962800# GND GND efet w=20300 l=10150
+ ad=1.39606e+09 pd=435000 as=0 ps=0 
M2889 GND diff_2314200_884500# diff_2275050_913500# GND efet w=12325 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2890 GND diff_2275050_913500# diff_2144550_958450# GND efet w=42050 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2891 diff_2144550_958450# diff_2172100_899000# diff_2144550_958450# GND efet w=51475 l=19575
+ ad=0 pd=0 as=0 ps=0 
M2892 diff_2144550_958450# diff_2172100_899000# GND GND efet w=5800 l=47850
+ ad=0 pd=0 as=0 ps=0 
M2893 GND diff_1925600_946850# diff_1784950_914950# GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2894 GND diff_1740000_820700# diff_1090400_862750# GND efet w=63075 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2895 GND diff_1608050_883050# diff_1547150_726450# GND efet w=5800 l=45675
+ ad=0 pd=0 as=0 ps=0 
M2896 diff_1547150_726450# diff_1608050_883050# diff_1547150_726450# GND efet w=79025 l=5075
+ ad=0 pd=0 as=0 ps=0 
M2897 diff_871450_1602250# GND GND GND efet w=8700 l=46400
+ ad=0 pd=0 as=0 ps=0 
M2898 GND GND GND GND efet w=8700 l=43500
+ ad=0 pd=0 as=0 ps=0 
M2899 GND GND GND GND efet w=35525 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2900 diff_535050_885950# diff_535050_885950# GND GND efet w=21025 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2901 GND GND GND GND efet w=41325 l=16675
+ ad=0 pd=0 as=0 ps=0 
M2902 GND diff_535050_885950# diff_597400_767050# GND efet w=12325 l=12325
+ ad=0 pd=0 as=4.3732e+08 ps=153700 
M2903 GND GND GND GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2904 GND GND GND GND efet w=35525 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2905 GND diff_597400_767050# GND GND efet w=50750 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2906 diff_717750_555350# GND GND GND efet w=14500 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2907 GND GND GND GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2908 GND GND GND GND efet w=15950 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2909 GND GND GND GND efet w=18125 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2910 GND GND diff_716300_748200# GND efet w=5800 l=59450
+ ad=0 pd=0 as=7.75823e+08 ps=249400 
M2911 GND diff_1090400_862750# diff_871450_1602250# GND efet w=39875 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2912 diff_1090400_862750# diff_1055600_1228150# GND GND efet w=39875 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2913 GND GND diff_1608050_883050# GND efet w=5800 l=11600
+ ad=0 pd=0 as=4.205e+07 ps=26100 
M2914 diff_1090400_862750# diff_1719700_845350# GND GND efet w=15950 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2915 GND GND diff_2038700_881600# GND efet w=7975 l=12325
+ ad=0 pd=0 as=9.251e+07 ps=52200 
M2916 GND diff_1087500_571300# GND GND efet w=39875 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2917 diff_1584850_851150# diff_1547150_726450# diff_1262950_843900# GND efet w=14500 l=13050
+ ad=1.98266e+09 pd=490100 as=-1.70258e+09 ps=710500 
M2918 diff_1841500_870000# diff_1784950_914950# diff_1809600_885950# GND efet w=57275 l=10875
+ ad=5.92905e+08 pd=174000 as=4.7937e+08 ps=159500 
M2919 diff_1809600_885950# diff_1584850_851150# GND GND efet w=58000 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2920 diff_1719700_845350# diff_1850200_854050# diff_1841500_870000# GND efet w=60175 l=11600
+ ad=9.71355e+08 pd=258100 as=0 ps=0 
M2921 GND GND diff_925100_1455800# GND efet w=23200 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2922 diff_1262950_843900# GND GND GND efet w=10875 l=35525
+ ad=0 pd=0 as=0 ps=0 
M2923 diff_1262950_843900# GND diff_1302100_807650# GND efet w=8700 l=11600
+ ad=0 pd=0 as=1.24468e+09 ps=406000 
M2924 diff_1262950_843900# GND GND GND efet w=32625 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2925 diff_1090400_903350# diff_1332550_1297750# diff_1302100_807650# GND efet w=8700 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2926 GND diff_1719700_845350# diff_1740000_820700# GND efet w=12325 l=10875
+ ad=0 pd=0 as=3.0276e+08 ps=145000 
M2927 diff_1784950_914950# diff_1784950_914950# diff_1944450_801850# GND efet w=56550 l=14500
+ ad=0 pd=0 as=1.44021e+09 ps=374100 
M2928 diff_1784950_914950# diff_1584850_851150# GND GND efet w=65975 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2929 diff_1944450_801850# diff_1850200_854050# GND GND efet w=48575 l=10875
+ ad=0 pd=0 as=0 ps=0 
M2930 GND diff_716300_748200# GND GND efet w=17400 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2931 diff_716300_748200# GND GND GND efet w=10875 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2932 GND GND diff_690200_720650# GND efet w=6525 l=68875
+ ad=0 pd=0 as=6.0552e+08 ps=217500 
M2933 diff_365400_716300# diff_339300_716300# GND GND efet w=27550 l=11600
+ ad=6.8962e+08 pd=208800 as=0 ps=0 
M2934 diff_339300_716300# GND diff_258100_694550# GND efet w=13775 l=12325
+ ad=1.49278e+08 pd=55100 as=0 ps=0 
M2935 diff_291450_822150# GND diff_365400_716300# GND efet w=14500 l=11600
+ ad=1.5138e+08 pd=60900 as=0 ps=0 
M2936 diff_365400_716300# GND diff_365400_716300# GND efet w=3625 l=42050
+ ad=0 pd=0 as=0 ps=0 
M2937 GND diff_527800_677150# GND GND efet w=49300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2938 diff_716300_748200# diff_535050_885950# diff_597400_767050# GND efet w=12325 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2939 diff_1925600_801850# diff_1850200_854050# diff_1784950_914950# GND efet w=57275 l=13775
+ ad=1.52852e+09 pd=490100 as=0 ps=0 
M2940 diff_1944450_801850# diff_1584850_851150# diff_1925600_801850# GND efet w=67425 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2941 diff_1925600_801850# diff_2038700_881600# diff_1925600_801850# GND efet w=50025 l=23200
+ ad=0 pd=0 as=0 ps=0 
M2942 diff_2172100_899000# GND GND GND efet w=8700 l=11600
+ ad=1.91328e+08 pd=66700 as=0 ps=0 
M2943 GND GND diff_2314200_884500# GND efet w=21750 l=15950
+ ad=0 pd=0 as=5.7188e+08 ps=133400 
M2944 diff_2314200_884500# GND GND GND efet w=10875 l=35525
+ ad=0 pd=0 as=0 ps=0 
M2945 GND diff_1584850_851150# diff_1796550_791700# GND efet w=34800 l=14500
+ ad=0 pd=0 as=9.65047e+08 ps=234900 
M2946 GND diff_1302100_807650# GND GND efet w=59450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2947 diff_1090400_862750# diff_1194800_1497850# diff_1302100_807650# GND efet w=8700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2948 diff_1740000_820700# GND GND GND efet w=7250 l=50025
+ ad=0 pd=0 as=0 ps=0 
M2949 GND GND GND GND efet w=10150 l=33350
+ ad=0 pd=0 as=0 ps=0 
M2950 diff_1051250_652500# diff_1426800_1106350# diff_1302100_807650# GND efet w=7975 l=13775
+ ad=4.8866e+08 pd=2.0735e+06 as=0 ps=0 
M2951 GND GND GND GND efet w=7250 l=33350
+ ad=0 pd=0 as=0 ps=0 
M2952 GND GND GND GND efet w=55100 l=14500
+ ad=0 pd=0 as=0 ps=0 
M2953 GND diff_1197700_311750# GND GND efet w=8700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2954 GND GND diff_1584850_851150# GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2955 diff_1719700_845350# GND GND GND efet w=5075 l=68875
+ ad=0 pd=0 as=0 ps=0 
M2956 diff_1796550_791700# GND diff_1719700_845350# GND efet w=35525 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2957 diff_1796550_791700# diff_1784950_914950# GND GND efet w=43500 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2958 GND diff_1850200_854050# diff_1796550_791700# GND efet w=36250 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2959 diff_1584850_851150# diff_1590650_513300# GND GND efet w=15950 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2960 diff_717750_555350# GND GND GND efet w=18125 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2961 GND GND GND GND efet w=11600 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2962 GND GND GND GND efet w=18850 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2963 diff_249400_1373150# diff_258100_694550# GND GND efet w=23200 l=13050
+ ad=0 pd=0 as=0 ps=0 
M2964 GND diff_594500_717750# diff_527800_677150# GND efet w=39150 l=11600
+ ad=0 pd=0 as=1.05966e+09 ps=316100 
M2965 GND GND GND GND efet w=31900 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2966 GND diff_1744350_653950# diff_1051250_652500# GND efet w=60900 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2967 GND diff_2038700_881600# diff_1925600_801850# GND efet w=5800 l=51475
+ ad=0 pd=0 as=0 ps=0 
M2968 diff_2143100_796050# diff_2122800_433550# diff_1850200_854050# GND efet w=14500 l=11600
+ ad=-1.52387e+09 pd=765600 as=1.11432e+09 ps=295800 
M2969 diff_2143100_796050# diff_2201100_846800# GND GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2970 diff_2409900_877250# GND GND GND efet w=57275 l=12325
+ ad=1.13114e+09 pd=237800 as=0 ps=0 
M2971 GND GND GND GND efet w=29725 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2972 GND GND diff_2409900_877250# GND efet w=10875 l=40600
+ ad=0 pd=0 as=0 ps=0 
M2973 GND GND GND GND efet w=7250 l=15950
+ ad=0 pd=0 as=0 ps=0 
M2974 GND GND GND GND efet w=7250 l=15225
+ ad=0 pd=0 as=0 ps=0 
M2975 GND GND GND GND efet w=54375 l=26100
+ ad=0 pd=0 as=0 ps=0 
M2976 GND GND GND GND efet w=10150 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2977 GND GND GND GND efet w=12325 l=18125
+ ad=0 pd=0 as=0 ps=0 
M2978 GND diff_2143100_796050# diff_2143100_796050# GND efet w=7975 l=18125
+ ad=0 pd=0 as=0 ps=0 
M2979 GND diff_1624000_314650# diff_2409900_877250# GND efet w=27550 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2980 diff_2201100_846800# GND GND GND efet w=5075 l=48575
+ ad=2.56505e+08 pd=121800 as=0 ps=0 
M2981 diff_1995200_817800# diff_1925600_801850# GND GND efet w=13050 l=10150
+ ad=2.12352e+08 pd=95700 as=0 ps=0 
M2982 GND GND diff_1995200_817800# GND efet w=7250 l=63075
+ ad=0 pd=0 as=0 ps=0 
M2983 GND diff_2143100_796050# diff_2201100_846800# GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2984 GND GND GND GND efet w=21750 l=67425
+ ad=0 pd=0 as=0 ps=0 
M2985 GND GND diff_2273600_775750# GND efet w=7975 l=10150
+ ad=0 pd=0 as=3.1958e+08 ps=95700 
M2986 diff_2143100_796050# diff_2201100_846800# GND GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2987 diff_2143100_796050# GND diff_1850200_854050# GND efet w=18125 l=12325
+ ad=0 pd=0 as=0 ps=0 
M2988 GND diff_2143100_796050# diff_2143100_796050# GND efet w=14500 l=17400
+ ad=0 pd=0 as=0 ps=0 
M2989 GND GND GND GND efet w=251575 l=23925
+ ad=0 pd=0 as=0 ps=0 
M2990 GND diff_2314200_884500# diff_2273600_775750# GND efet w=12325 l=13775
+ ad=0 pd=0 as=0 ps=0 
M2991 GND diff_1995200_817800# GND GND efet w=20300 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2992 GND GND GND GND efet w=226925 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2993 GND diff_2273600_775750# diff_2143100_796050# GND efet w=41325 l=18125
+ ad=0 pd=0 as=0 ps=0 
M2994 GND diff_1925600_801850# GND GND efet w=14500 l=10150
+ ad=0 pd=0 as=0 ps=0 
M2995 diff_2143100_796050# diff_2172100_739500# diff_2143100_796050# GND efet w=50025 l=20300
+ ad=0 pd=0 as=0 ps=0 
M2996 diff_2143100_796050# diff_2172100_739500# GND GND efet w=5800 l=43500
+ ad=0 pd=0 as=0 ps=0 
M2997 GND diff_1161450_745300# GND GND efet w=56550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M2998 diff_1290500_722100# diff_1197700_311750# diff_1161450_745300# GND efet w=7250 l=13050
+ ad=-1.3788e+09 pd=669900 as=4.01578e+08 ps=127600 
M2999 GND GND GND GND efet w=8700 l=29000
+ ad=0 pd=0 as=0 ps=0 
M3000 GND diff_337850_655400# diff_258100_694550# GND efet w=41325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3001 diff_258100_694550# diff_292900_675700# GND GND efet w=37700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3002 GND GND diff_527800_677150# GND efet w=18850 l=15950
+ ad=0 pd=0 as=0 ps=0 
M3003 diff_527800_677150# GND GND GND efet w=7250 l=49300
+ ad=0 pd=0 as=0 ps=0 
M3004 diff_690200_720650# diff_535050_885950# diff_594500_717750# GND efet w=12325 l=15225
+ ad=0 pd=0 as=2.45992e+08 ps=124700 
M3005 GND diff_690200_720650# GND GND efet w=17400 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3006 GND GND diff_717750_555350# GND efet w=24650 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3007 GND GND GND GND efet w=10875 l=15225
+ ad=0 pd=0 as=0 ps=0 
M3008 diff_690200_720650# GND GND GND efet w=14500 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3009 GND diff_1547150_726450# diff_1290500_722100# GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3010 diff_1051250_652500# diff_1731300_701800# GND GND efet w=13775 l=15225
+ ad=0 pd=0 as=0 ps=0 
M3011 diff_1290500_722100# GND GND GND efet w=10150 l=41325
+ ad=0 pd=0 as=0 ps=0 
M3012 GND GND GND GND efet w=14500 l=14500
+ ad=0 pd=0 as=0 ps=0 
M3013 GND GND GND GND efet w=32625 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3014 GND diff_527800_677150# GND GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3015 GND GND GND GND efet w=7250 l=52200
+ ad=0 pd=0 as=0 ps=0 
M3016 diff_337850_655400# diff_346550_629300# diff_337850_655400# GND efet w=69600 l=5800
+ ad=1.04074e+09 pd=339300 as=0 ps=0 
M3017 diff_337850_655400# diff_292900_675700# GND GND efet w=32625 l=15225
+ ad=0 pd=0 as=0 ps=0 
M3018 GND GND diff_346550_629300# GND efet w=6525 l=13775
+ ad=0 pd=0 as=6.3075e+07 ps=40600 
M3019 GND diff_346550_629300# diff_337850_655400# GND efet w=5800 l=24650
+ ad=0 pd=0 as=0 ps=0 
M3020 GND diff_535050_885950# diff_594500_717750# GND efet w=10150 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3021 GND GND diff_711950_652500# GND efet w=6525 l=73225
+ ad=0 pd=0 as=3.97373e+08 ps=165300 
M3022 diff_711950_652500# diff_535050_885950# GND GND efet w=10150 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3023 GND diff_711950_652500# GND GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3024 diff_711950_652500# GND GND GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3025 GND GND diff_925100_1455800# GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3026 diff_1090400_862750# diff_1332550_1297750# GND GND efet w=7250 l=14500
+ ad=0 pd=0 as=0 ps=0 
M3027 GND GND diff_1290500_722100# GND efet w=54375 l=21750
+ ad=0 pd=0 as=0 ps=0 
M3028 diff_1262950_671350# GND GND GND efet w=12325 l=36975
+ ad=-1.37459e+09 pd=768500 as=0 ps=0 
M3029 GND diff_1051250_652500# diff_871450_1602250# GND efet w=42775 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3030 GND diff_1087500_571300# GND GND efet w=39150 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3031 diff_1051250_652500# diff_1194800_1497850# GND GND efet w=7975 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3032 GND GND diff_1262950_671350# GND efet w=7975 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3033 GND diff_1290500_722100# diff_1262950_671350# GND efet w=36250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3034 diff_1841500_707600# GND diff_1808150_742400# GND efet w=59450 l=11600
+ ad=6.43365e+08 pd=179800 as=5.15113e+08 ps=162400 
M3035 diff_1808150_742400# GND GND GND efet w=60900 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3036 diff_1744350_653950# diff_1796550_646700# diff_1841500_707600# GND efet w=65250 l=10875
+ ad=1.62944e+09 pd=420500 as=0 ps=0 
M3037 GND GND GND GND efet w=63075 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3038 GND diff_1744350_653950# diff_1731300_701800# GND efet w=10150 l=12325
+ ad=0 pd=0 as=2.33378e+08 ps=78300 
M3039 GND GND GND GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3040 diff_1051250_593050# diff_1426800_1106350# GND GND efet w=9425 l=12325
+ ad=-1.0798e+09 pd=1.6994e+06 as=0 ps=0 
M3041 diff_1796550_646700# diff_1796550_646700# GND GND efet w=50750 l=13050
+ ad=-5.02057e+08 pd=988900 as=0 ps=0 
M3042 diff_1796550_646700# GND diff_1925600_656850# GND efet w=68150 l=14500
+ ad=0 pd=0 as=9.3351e+08 ps=243600 
M3043 diff_1925600_656850# diff_1796550_646700# GND GND efet w=56550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3044 diff_1731300_701800# GND GND GND efet w=5800 l=68875
+ ad=0 pd=0 as=0 ps=0 
M3045 GND diff_1055600_1228150# diff_1051250_652500# GND efet w=42775 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3046 GND diff_1590650_513300# diff_1262950_671350# GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3047 diff_1744350_653950# GND GND GND efet w=7250 l=59450
+ ad=0 pd=0 as=0 ps=0 
M3048 GND GND GND GND efet w=40600 l=13050
+ ad=0 pd=0 as=0 ps=0 
M3049 diff_365400_569850# diff_339300_571300# GND GND efet w=27550 l=11600
+ ad=6.62287e+08 pd=208800 as=0 ps=0 
M3050 diff_292900_675700# GND diff_365400_569850# GND efet w=13775 l=12325
+ ad=1.30355e+08 pd=58000 as=0 ps=0 
M3051 diff_339300_571300# GND diff_258100_549550# GND efet w=15950 l=11600
+ ad=1.30355e+08 pd=55100 as=-2.04021e+09 ps=2.2794e+06 
M3052 GND GND GND GND efet w=40600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3053 GND GND diff_717750_555350# GND efet w=18850 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3054 GND GND GND GND efet w=19575 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3055 GND GND GND GND efet w=15950 l=14500
+ ad=0 pd=0 as=0 ps=0 
M3056 GND GND GND GND efet w=33350 l=13050
+ ad=0 pd=0 as=0 ps=0 
M3057 diff_1796550_646700# diff_1744350_653950# diff_1744350_653950# GND efet w=29725 l=17400
+ ad=0 pd=0 as=0 ps=0 
M3058 GND GND diff_1796550_646700# GND efet w=36250 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3059 diff_1796550_646700# GND GND GND efet w=38425 l=16675
+ ad=0 pd=0 as=0 ps=0 
M3060 GND diff_1796550_646700# diff_1796550_646700# GND efet w=36250 l=17400
+ ad=0 pd=0 as=0 ps=0 
M3061 diff_1590650_513300# diff_1616750_597400# diff_1590650_513300# GND efet w=81200 l=4350
+ ad=0 pd=0 as=0 ps=0 
M3062 GND GND diff_1796550_646700# GND efet w=56550 l=15950
+ ad=0 pd=0 as=0 ps=0 
M3063 GND GND GND GND efet w=68875 l=38425
+ ad=0 pd=0 as=0 ps=0 
M3064 GND diff_2314200_884500# GND GND efet w=19575 l=17400
+ ad=0 pd=0 as=0 ps=0 
M3065 GND GND GND GND efet w=60175 l=25375
+ ad=0 pd=0 as=0 ps=0 
M3066 diff_2172100_739500# GND GND GND efet w=9425 l=12325
+ ad=1.99738e+08 pd=63800 as=0 ps=0 
M3067 GND GND diff_1925600_656850# GND efet w=5800 l=58000
+ ad=0 pd=0 as=0 ps=0 
M3068 diff_2144550_636550# diff_2201100_690200# GND GND efet w=22475 l=11600
+ ad=-1.75515e+09 pd=707600 as=0 ps=0 
M3069 diff_2144550_636550# diff_2122800_433550# diff_1796550_646700# GND efet w=15950 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3070 GND diff_2144550_636550# diff_2144550_636550# GND efet w=8700 l=18850
+ ad=0 pd=0 as=0 ps=0 
M3071 GND GND GND GND efet w=1178125 l=31900
+ ad=0 pd=0 as=0 ps=0 
M3072 GND GND GND GND efet w=8700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3073 diff_2385250_669900# diff_1352850_295800# GND GND efet w=26100 l=13050
+ ad=8.38897e+08 pd=220400 as=0 ps=0 
M3074 diff_1995200_672800# diff_1925600_656850# GND GND efet w=13050 l=10875
+ ad=2.0184e+08 pd=92800 as=0 ps=0 
M3075 GND GND diff_1995200_672800# GND efet w=5800 l=63800
+ ad=0 pd=0 as=0 ps=0 
M3076 diff_1744350_653950# diff_1995200_672800# GND GND efet w=20300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3077 GND diff_1925600_656850# diff_1744350_653950# GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3078 GND GND diff_2041600_566950# GND efet w=5800 l=11600
+ ad=0 pd=0 as=4.41525e+07 ps=29000 
M3079 diff_2201100_690200# GND GND GND efet w=5075 l=47125
+ ad=2.31275e+08 pd=116000 as=0 ps=0 
M3080 GND diff_2144550_636550# diff_2201100_690200# GND efet w=13775 l=15225
+ ad=0 pd=0 as=0 ps=0 
M3081 diff_2144550_636550# diff_2201100_690200# GND GND efet w=15950 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3082 GND diff_2144550_636550# diff_2144550_636550# GND efet w=13775 l=19575
+ ad=0 pd=0 as=0 ps=0 
M3083 diff_2144550_636550# GND diff_1796550_646700# GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3084 GND GND GND GND efet w=599575 l=54375
+ ad=0 pd=0 as=0 ps=0 
M3085 GND GND diff_2385250_669900# GND efet w=11600 l=52200
+ ad=0 pd=0 as=0 ps=0 
M3086 diff_2385250_669900# GND GND GND efet w=10150 l=17400
+ ad=0 pd=0 as=0 ps=0 
M3087 diff_2144550_636550# diff_2177900_597400# GND GND efet w=8700 l=53650
+ ad=0 pd=0 as=0 ps=0 
M3088 GND GND GND GND efet w=3625 l=64525
+ ad=0 pd=0 as=0 ps=0 
M3089 GND diff_1616750_597400# diff_1590650_513300# GND efet w=6525 l=45675
+ ad=0 pd=0 as=0 ps=0 
M3090 GND GND diff_365400_569850# GND efet w=7250 l=38425
+ ad=0 pd=0 as=0 ps=0 
M3091 diff_249400_1373150# diff_258100_549550# GND GND efet w=22475 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3092 GND GND GND GND efet w=8700 l=43500
+ ad=0 pd=0 as=0 ps=0 
M3093 GND GND GND GND efet w=7250 l=43500
+ ad=0 pd=0 as=0 ps=0 
M3094 GND diff_337850_514750# diff_258100_549550# GND efet w=39150 l=13050
+ ad=0 pd=0 as=0 ps=0 
M3095 GND GND GND GND efet w=22475 l=14500
+ ad=0 pd=0 as=0 ps=0 
M3096 GND GND GND GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3097 diff_258100_549550# diff_292900_530700# GND GND efet w=38425 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3098 diff_337850_514750# diff_346550_482850# diff_337850_514750# GND efet w=68150 l=5800
+ ad=1.05966e+09 pd=345100 as=0 ps=0 
M3099 diff_337850_514750# diff_292900_530700# GND GND efet w=27550 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3100 GND GND diff_346550_482850# GND efet w=5800 l=12325
+ ad=0 pd=0 as=7.35875e+07 ps=37700 
M3101 GND diff_535050_885950# GND GND efet w=9425 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3102 GND GND diff_717750_555350# GND efet w=13775 l=18850
+ ad=0 pd=0 as=0 ps=0 
M3103 GND GND GND GND efet w=15225 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3104 GND GND GND GND efet w=11600 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3105 GND diff_1051250_593050# diff_871450_1602250# GND efet w=41325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3106 GND GND GND GND efet w=17400 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3107 GND GND GND GND efet w=16675 l=18125
+ ad=0 pd=0 as=0 ps=0 
M3108 GND GND GND GND efet w=33350 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3109 GND diff_346550_482850# diff_337850_514750# GND efet w=5800 l=26100
+ ad=0 pd=0 as=0 ps=0 
M3110 diff_1051250_593050# diff_1055600_1228150# GND GND efet w=40600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3111 GND GND diff_1616750_597400# GND efet w=5800 l=10150
+ ad=0 pd=0 as=3.364e+07 ps=23200 
M3112 diff_1051250_593050# diff_1718250_556800# GND GND efet w=19575 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3113 GND diff_1087500_571300# GND GND efet w=40600 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3114 diff_1584850_569850# diff_1547150_726450# diff_1262950_575650# GND efet w=15950 l=13775
+ ad=6.8165e+08 pd=1.5892e+06 as=-1.62269e+09 ps=727900 
M3115 GND GND GND GND efet w=62350 l=15950
+ ad=0 pd=0 as=0 ps=0 
M3116 GND diff_717750_555350# GND GND efet w=72500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3117 GND GND GND GND efet w=61625 l=16675
+ ad=0 pd=0 as=0 ps=0 
M3118 GND GND GND GND efet w=74675 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3119 GND GND GND GND efet w=54375 l=16675
+ ad=0 pd=0 as=0 ps=0 
M3120 GND GND GND GND efet w=5800 l=66700
+ ad=0 pd=0 as=0 ps=0 
M3121 GND diff_651050_437900# GND GND efet w=76850 l=7250
+ ad=0 pd=0 as=0 ps=0 
M3122 GND GND GND GND efet w=26825 l=31175
+ ad=0 pd=0 as=0 ps=0 
M3123 diff_292900_530700# GND diff_365400_424850# GND efet w=13775 l=10150
+ ad=1.38765e+08 pd=60900 as=6.2234e+08 ps=208800 
M3124 diff_365400_424850# diff_340750_424850# GND GND efet w=29000 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3125 GND GND diff_365400_424850# GND efet w=5075 l=42050
+ ad=0 pd=0 as=0 ps=0 
M3126 diff_340750_424850# GND diff_249400_1373150# GND efet w=13050 l=11600
+ ad=1.15638e+08 pd=49300 as=0 ps=0 
M3127 GND GND GND GND efet w=44225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3128 GND GND diff_651050_437900# GND efet w=4350 l=15950
+ ad=0 pd=0 as=6.51775e+07 ps=40600 
M3129 GND diff_651050_437900# GND GND efet w=10150 l=24650
+ ad=0 pd=0 as=0 ps=0 
M3130 GND GND GND GND efet w=5800 l=66700
+ ad=0 pd=0 as=0 ps=0 
M3131 GND GND diff_249400_1373150# GND efet w=4350 l=39150
+ ad=0 pd=0 as=0 ps=0 
M3132 GND diff_651050_353800# GND GND efet w=76850 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3133 GND GND GND GND efet w=35525 l=21025
+ ad=0 pd=0 as=0 ps=0 
M3134 GND GND GND GND efet w=115275 l=38425
+ ad=0 pd=0 as=0 ps=0 
M3135 GND GND GND GND efet w=47850 l=18850
+ ad=0 pd=0 as=0 ps=0 
M3136 GND GND GND GND efet w=43500 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3137 GND GND GND GND efet w=55100 l=17400
+ ad=0 pd=0 as=0 ps=0 
M3138 GND GND GND GND efet w=59450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3139 GND GND GND GND efet w=55825 l=15950
+ ad=0 pd=0 as=0 ps=0 
M3140 GND GND GND GND efet w=59450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3141 GND GND GND GND efet w=60900 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3142 GND GND diff_925100_1455800# GND efet w=23200 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3143 diff_1262950_575650# GND GND GND efet w=10875 l=35525
+ ad=0 pd=0 as=0 ps=0 
M3144 GND diff_1158550_546650# GND GND efet w=53650 l=13050
+ ad=0 pd=0 as=0 ps=0 
M3145 GND GND GND GND efet w=8700 l=34800
+ ad=0 pd=0 as=0 ps=0 
M3146 GND GND GND GND efet w=60175 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3147 GND GND diff_651050_353800# GND efet w=7975 l=12325
+ ad=0 pd=0 as=6.728e+07 ps=40600 
M3148 GND GND GND GND efet w=139925 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3149 GND GND GND GND efet w=5075 l=23925
+ ad=0 pd=0 as=0 ps=0 
M3150 GND GND GND GND efet w=6525 l=22475
+ ad=0 pd=0 as=0 ps=0 
M3151 GND GND GND GND efet w=40600 l=13050
+ ad=0 pd=0 as=0 ps=0 
M3152 GND diff_651050_353800# GND GND efet w=10150 l=24650
+ ad=0 pd=0 as=0 ps=0 
M3153 GND GND GND GND efet w=4350 l=63800
+ ad=0 pd=0 as=0 ps=0 
M3154 GND diff_717750_555350# GND GND efet w=61625 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3155 diff_772850_316100# GND GND GND efet w=6525 l=68150
+ ad=-2.28732e+08 pd=959900 as=0 ps=0 
M3156 GND diff_681500_266800# GND GND efet w=79025 l=6525
+ ad=0 pd=0 as=0 ps=0 
M3157 GND GND GND GND efet w=230550 l=47850
+ ad=0 pd=0 as=0 ps=0 
M3158 GND GND GND GND efet w=229825 l=45675
+ ad=0 pd=0 as=0 ps=0 
M3159 GND GND GND GND efet w=37700 l=18850
+ ad=0 pd=0 as=0 ps=0 
M3160 GND GND GND GND efet w=59450 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3161 GND GND GND GND efet w=74675 l=6525
+ ad=0 pd=0 as=0 ps=0 
M3162 GND GND GND GND efet w=7975 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3163 GND GND GND GND efet w=42775 l=15225
+ ad=0 pd=0 as=0 ps=0 
M3164 GND GND GND GND efet w=60175 l=18125
+ ad=0 pd=0 as=0 ps=0 
M3165 GND GND GND GND efet w=60175 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3166 GND GND GND GND efet w=48575 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3167 GND GND GND GND efet w=44950 l=18850
+ ad=0 pd=0 as=0 ps=0 
M3168 GND GND GND GND efet w=53650 l=17400
+ ad=0 pd=0 as=0 ps=0 
M3169 diff_681500_266800# GND diff_681500_266800# GND efet w=4350 l=15950
+ ad=5.67675e+07 pd=31900 as=0 ps=0 
M3170 GND diff_681500_266800# GND GND efet w=10875 l=23925
+ ad=0 pd=0 as=0 ps=0 
M3171 GND GND GND GND efet w=9425 l=22475
+ ad=0 pd=0 as=0 ps=0 
M3172 GND diff_717750_555350# diff_772850_316100# GND efet w=62350 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3173 GND GND diff_772850_316100# GND efet w=63800 l=15950
+ ad=0 pd=0 as=0 ps=0 
M3174 GND GND diff_772850_316100# GND efet w=60175 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3175 GND GND GND GND efet w=46400 l=15950
+ ad=0 pd=0 as=0 ps=0 
M3176 GND GND diff_772850_316100# GND efet w=51475 l=15950
+ ad=0 pd=0 as=0 ps=0 
M3177 diff_1262950_575650# GND diff_1302100_537950# GND efet w=8700 l=11600
+ ad=0 pd=0 as=1.27411e+09 ps=397300 
M3178 diff_1262950_575650# GND GND GND efet w=34075 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3179 diff_1051250_652500# diff_1332550_1297750# diff_1302100_537950# GND efet w=8700 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3180 GND diff_1738550_530700# diff_1051250_593050# GND efet w=65975 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3181 GND GND diff_2144550_636550# GND efet w=36250 l=18850
+ ad=0 pd=0 as=0 ps=0 
M3182 diff_1808150_595950# diff_1584850_569850# GND GND efet w=60175 l=10875
+ ad=5.17215e+08 pd=156600 as=0 ps=0 
M3183 GND diff_1718250_556800# diff_1738550_530700# GND efet w=13775 l=10150
+ ad=0 pd=0 as=3.17478e+08 ps=130500 
M3184 diff_1841500_561150# diff_1744350_653950# diff_1808150_595950# GND efet w=56550 l=11600
+ ad=6.53878e+08 pd=182700 as=0 ps=0 
M3185 diff_1718250_556800# diff_1584850_569850# diff_1841500_561150# GND efet w=65250 l=10150
+ ad=1.0092e+09 pd=281300 as=0 ps=0 
M3186 diff_1584850_569850# diff_1584850_569850# GND GND efet w=73950 l=21750
+ ad=0 pd=0 as=0 ps=0 
M3187 GND diff_1584850_569850# diff_1943000_511850# GND efet w=61625 l=28275
+ ad=0 pd=0 as=1.49488e+09 ps=371200 
M3188 GND diff_1302100_537950# GND GND efet w=58725 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3189 diff_1051250_593050# diff_1194800_1497850# diff_1302100_537950# GND efet w=9425 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3190 GND GND GND GND efet w=9425 l=35525
+ ad=0 pd=0 as=0 ps=0 
M3191 diff_1051250_593050# diff_1332550_1297750# diff_1426800_1106350# GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3192 GND diff_1197700_311750# diff_1158550_546650# GND efet w=7250 l=13050
+ ad=0 pd=0 as=3.93167e+08 ps=127600 
M3193 diff_1426800_1106350# diff_1426800_1106350# diff_1302100_537950# GND efet w=13050 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3194 diff_1584850_569850# diff_1584850_569850# diff_1584850_569850# GND efet w=55825 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3195 GND diff_1584850_569850# diff_1584850_569850# GND efet w=30450 l=17400
+ ad=0 pd=0 as=0 ps=0 
M3196 diff_1738550_530700# GND GND GND efet w=5800 l=58000
+ ad=0 pd=0 as=0 ps=0 
M3197 GND GND diff_1584850_569850# GND efet w=13775 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3198 diff_1584850_569850# diff_1448550_1090400# diff_1718250_556800# GND efet w=37700 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3199 diff_1718250_556800# GND GND GND efet w=7250 l=65250
+ ad=0 pd=0 as=0 ps=0 
M3200 diff_1584850_569850# diff_1590650_513300# GND GND efet w=15950 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3201 diff_1943000_511850# diff_1584850_569850# diff_1584850_569850# GND efet w=65250 l=17400
+ ad=0 pd=0 as=0 ps=0 
M3202 diff_1584850_569850# diff_1744350_653950# GND GND efet w=43500 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3203 GND diff_1584850_569850# diff_1584850_569850# GND efet w=35525 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3204 diff_1584850_569850# diff_1744350_653950# diff_1943000_511850# GND efet w=58000 l=10150
+ ad=0 pd=0 as=0 ps=0 
M3205 diff_2144550_636550# diff_2177900_597400# diff_2144550_636550# GND efet w=46400 l=21025
+ ad=0 pd=0 as=0 ps=0 
M3206 diff_1584850_569850# diff_2041600_566950# diff_1584850_569850# GND efet w=57275 l=34075
+ ad=0 pd=0 as=0 ps=0 
M3207 diff_2177900_597400# GND GND GND efet w=12325 l=13050
+ ad=1.19842e+08 pd=72500 as=0 ps=0 
M3208 GND GND GND GND efet w=42050 l=21025
+ ad=0 pd=0 as=0 ps=0 
M3209 GND diff_2385250_669900# GND GND efet w=39875 l=15225
+ ad=0 pd=0 as=0 ps=0 
M3210 GND diff_2041600_566950# diff_1584850_569850# GND efet w=5075 l=52200
+ ad=0 pd=0 as=0 ps=0 
M3211 GND GND GND GND efet w=10150 l=39150
+ ad=0 pd=0 as=0 ps=0 
M3212 diff_2144550_503150# diff_2199650_546650# GND GND efet w=21025 l=13050
+ ad=-1.49444e+09 pd=774300 as=0 ps=0 
M3213 GND GND GND GND efet w=66700 l=16675
+ ad=0 pd=0 as=0 ps=0 
M3214 diff_2144550_503150# GND diff_1584850_569850# GND efet w=14500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3215 GND diff_1352850_295800# GND GND efet w=44950 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3216 GND diff_2144550_503150# diff_2144550_503150# GND efet w=8700 l=17400
+ ad=0 pd=0 as=0 ps=0 
M3217 diff_1998100_527800# diff_1584850_569850# GND GND efet w=12325 l=12325
+ ad=1.55585e+08 pd=84100 as=0 ps=0 
M3218 GND GND diff_1998100_527800# GND efet w=5800 l=63800
+ ad=0 pd=0 as=0 ps=0 
M3219 diff_1448550_1090400# diff_1998100_527800# GND GND efet w=18850 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3220 diff_2199650_546650# GND GND GND efet w=6525 l=45675
+ ad=2.56505e+08 pd=118900 as=0 ps=0 
M3221 GND diff_2144550_503150# diff_2199650_546650# GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3222 GND GND diff_2304050_481400# GND efet w=9425 l=8700
+ ad=0 pd=0 as=3.09067e+08 ps=92800 
M3223 diff_2144550_503150# diff_2122800_433550# diff_1584850_569850# GND efet w=15225 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3224 diff_2144550_503150# diff_2199650_546650# GND GND efet w=13775 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3225 GND diff_1584850_569850# diff_1448550_1090400# GND efet w=13050 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3226 GND GND diff_2201100_484300# GND efet w=6525 l=9425
+ ad=0 pd=0 as=4.205e+07 ps=26100 
M3227 GND diff_2144550_503150# diff_2144550_503150# GND efet w=15950 l=15950
+ ad=0 pd=0 as=0 ps=0 
M3228 GND diff_2314200_884500# diff_2304050_481400# GND efet w=14500 l=14500
+ ad=0 pd=0 as=0 ps=0 
M3229 diff_2144550_503150# diff_2201100_484300# diff_2144550_503150# GND efet w=68150 l=5800
+ ad=0 pd=0 as=0 ps=0 
M3230 GND diff_2304050_481400# diff_2144550_503150# GND efet w=38425 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3231 GND GND GND GND efet w=116000 l=13050
+ ad=0 pd=0 as=0 ps=0 
M3232 diff_1197700_311750# diff_1196250_255200# diff_1197700_311750# GND efet w=57275 l=17400
+ ad=0 pd=0 as=0 ps=0 
M3233 GND GND diff_772850_316100# GND efet w=60175 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3234 GND GND diff_2083650_427750# GND efet w=7250 l=9425
+ ad=0 pd=0 as=5.25625e+07 ps=34800 
M3235 diff_2144550_503150# diff_2201100_484300# GND GND efet w=5800 l=40600
+ ad=0 pd=0 as=0 ps=0 
M3236 diff_2122800_433550# diff_2083650_427750# diff_2122800_433550# GND efet w=66700 l=5800
+ ad=0 pd=0 as=0 ps=0 
M3237 diff_1370250_332050# GND GND GND efet w=71775 l=12325
+ ad=1.75979e+09 pd=394400 as=0 ps=0 
M3238 GND diff_1370250_332050# GND GND efet w=49300 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3239 GND diff_1370250_332050# diff_1416650_342200# GND efet w=13775 l=11600
+ ad=0 pd=0 as=7.94745e+08 ps=229100 
M3240 GND GND GND GND efet w=114550 l=14500
+ ad=0 pd=0 as=0 ps=0 
M3241 diff_1197700_311750# diff_1196250_255200# GND GND efet w=7250 l=52200
+ ad=0 pd=0 as=0 ps=0 
M3242 GND GND diff_1196250_255200# GND efet w=8700 l=13050
+ ad=0 pd=0 as=1.36662e+08 ps=55100 
M3243 diff_1370250_332050# diff_1352850_295800# GND GND efet w=51475 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3244 GND diff_1352850_295800# diff_1416650_342200# GND efet w=25375 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3245 GND diff_1416650_342200# GND GND efet w=38425 l=13050
+ ad=0 pd=0 as=0 ps=0 
M3246 diff_1370250_332050# GND GND GND efet w=10150 l=36975
+ ad=0 pd=0 as=0 ps=0 
M3247 diff_1416650_342200# GND GND GND efet w=5800 l=50750
+ ad=0 pd=0 as=0 ps=0 
M3248 GND GND diff_1635600_343650# GND efet w=57275 l=12325
+ ad=0 pd=0 as=8.64127e+08 ps=217500 
M3249 diff_1635600_343650# GND GND GND efet w=13050 l=39150
+ ad=0 pd=0 as=0 ps=0 
M3250 diff_1635600_343650# diff_1624000_314650# diff_1558750_169650# GND efet w=27550 l=11600
+ ad=0 pd=0 as=3.25887e+08 ps=92800 
M3251 GND diff_1558750_169650# GND GND efet w=99325 l=10875
+ ad=0 pd=0 as=0 ps=0 
M3252 GND GND GND GND efet w=645250 l=31900
+ ad=0 pd=0 as=0 ps=0 
M3253 GND GND GND GND efet w=50025 l=19575
+ ad=0 pd=0 as=0 ps=0 
M3254 GND GND GND GND efet w=129775 l=23925
+ ad=0 pd=0 as=0 ps=0 
M3255 GND GND GND GND efet w=127600 l=26100
+ ad=0 pd=0 as=0 ps=0 
M3256 GND GND GND GND efet w=7250 l=23200
+ ad=0 pd=0 as=0 ps=0 
M3257 GND GND GND GND efet w=6525 l=23925
+ ad=0 pd=0 as=0 ps=0 
M3258 GND GND GND GND efet w=43500 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3259 GND GND GND GND efet w=230550 l=43500
+ ad=0 pd=0 as=0 ps=0 
M3260 GND GND GND GND efet w=216775 l=51475
+ ad=0 pd=0 as=0 ps=0 
M3261 GND GND GND GND efet w=1210750 l=14500
+ ad=0 pd=0 as=0 ps=0 
M3262 GND GND GND GND efet w=247950 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3263 GND GND GND GND efet w=9425 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3264 GND GND GND GND efet w=10875 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3265 GND GND GND GND efet w=65250 l=18850
+ ad=0 pd=0 as=0 ps=0 
M3266 GND GND GND GND efet w=81925 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3267 GND GND GND GND efet w=229100 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3268 GND diff_1644300_82650# GND GND efet w=10150 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3269 GND diff_1644300_82650# GND GND efet w=58000 l=34800
+ ad=0 pd=0 as=0 ps=0 
M3270 GND GND diff_1644300_82650# GND efet w=10150 l=13050
+ ad=0 pd=0 as=4.83575e+07 ps=34800 
M3271 GND GND GND GND efet w=66700 l=13050
+ ad=0 pd=0 as=0 ps=0 
M3272 diff_2122800_433550# diff_2083650_427750# GND GND efet w=6525 l=33350
+ ad=0 pd=0 as=0 ps=0 
M3273 GND GND GND GND efet w=99325 l=15225
+ ad=0 pd=0 as=0 ps=0 
M3274 GND GND GND GND efet w=44950 l=15950
+ ad=0 pd=0 as=0 ps=0 
M3275 diff_2096700_342200# GND GND GND efet w=16675 l=10875
+ ad=7.35875e+08 pd=194300 as=0 ps=0 
M3276 GND diff_1352850_295800# diff_2096700_342200# GND efet w=26825 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3277 GND diff_1352850_295800# GND GND efet w=44225 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3278 GND GND diff_2096700_342200# GND efet w=6525 l=55825
+ ad=0 pd=0 as=0 ps=0 
M3279 GND diff_2096700_342200# GND GND efet w=39150 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3280 GND GND GND GND efet w=6525 l=37700
+ ad=0 pd=0 as=0 ps=0 
M3281 GND GND diff_2311300_334950# GND efet w=50750 l=10875
+ ad=0 pd=0 as=9.31407e+08 ps=226200 
M3282 diff_2311300_334950# diff_1624000_314650# GND GND efet w=27550 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3283 diff_2311300_334950# GND GND GND efet w=10875 l=36975
+ ad=0 pd=0 as=0 ps=0 
M3284 GND diff_1352850_295800# GND GND efet w=49300 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3285 GND diff_2444700_139200# GND GND efet w=39875 l=12325
+ ad=0 pd=0 as=0 ps=0 
M3286 GND GND GND GND efet w=29000 l=14500
+ ad=0 pd=0 as=0 ps=0 
M3287 GND GND GND GND efet w=656125 l=36975
+ ad=0 pd=0 as=0 ps=0 
M3288 GND GND GND GND efet w=33350 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3289 GND GND GND GND efet w=73950 l=36250
+ ad=0 pd=0 as=0 ps=0 
M3290 GND GND GND GND efet w=243600 l=33350
+ ad=0 pd=0 as=0 ps=0 
M3291 GND GND GND GND efet w=7250 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3292 GND GND GND GND efet w=9425 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3293 GND GND GND GND efet w=1203500 l=20300
+ ad=0 pd=0 as=0 ps=0 
M3294 GND GND GND GND efet w=60900 l=21750
+ ad=0 pd=0 as=0 ps=0 
M3295 GND GND diff_2444700_139200# GND efet w=9425 l=49300
+ ad=0 pd=0 as=7.44285e+08 ps=220400 
M3296 GND GND diff_1352850_295800# GND efet w=8700 l=36250
+ ad=0 pd=0 as=0 ps=0 
M3297 GND diff_1352850_295800# diff_1352850_295800# GND efet w=50025 l=21025
+ ad=0 pd=0 as=0 ps=0 
M3298 GND GND GND GND efet w=75400 l=13050
+ ad=0 pd=0 as=0 ps=0 
M3299 GND GND GND GND efet w=217500 l=23200
+ ad=0 pd=0 as=0 ps=0 
M3300 GND GND GND GND efet w=10150 l=14500
+ ad=0 pd=0 as=0 ps=0 
M3301 GND GND GND GND efet w=35525 l=58725
+ ad=0 pd=0 as=0 ps=0 
M3302 GND GND GND GND efet w=7250 l=13775
+ ad=0 pd=0 as=0 ps=0 
M3303 GND diff_1352850_295800# diff_2444700_139200# GND efet w=23200 l=15950
+ ad=0 pd=0 as=0 ps=0 
M3304 diff_2444700_139200# diff_1352850_295800# GND GND efet w=23925 l=11600
+ ad=0 pd=0 as=0 ps=0 
M3305 GND GND diff_1352850_295800# GND efet w=86275 l=15225
+ ad=0 pd=0 as=0 ps=0 
M3306 GND GND GND GND efet w=110925 l=26825
+ ad=0 pd=0 as=0 ps=0 
M3307 GND GND GND GND efet w=30450 l=10875
+ ad=0 pd=0 as=0 ps=0 
C0 metal_2544750_3477100# gnd! 33.7fF ;**FLOATING
C1 metal_2525900_3472750# gnd! 73.8fF ;**FLOATING
C2 metal_2537500_3545250# gnd! 29.1fF ;**FLOATING
C3 metal_2511400_3548150# gnd! 4.4fF ;**FLOATING
C4 metal_2625950_3569900# gnd! 7.6fF ;**FLOATING
C5 metal_2670900_3567000# gnd! 26.0fF ;**FLOATING
C6 metal_2537500_3571350# gnd! 62.4fF ;**FLOATING
C7 metal_2670900_3626450# gnd! 17.9fF ;**FLOATING
C8 metal_2625950_3607600# gnd! 13.8fF ;**FLOATING
C9 metal_105850_3567000# gnd! 31.4fF ;**FLOATING
C10 metal_105850_3623550# gnd! 30.1fF ;**FLOATING
C11 metal_2511400_3772900# gnd! 195.8fF ;**FLOATING
C12 metal_2016950_3793200# gnd! 221.7fF ;**FLOATING
C13 metal_1299200_3830900# gnd! 54.9fF ;**FLOATING
C14 metal_1190450_3787400# gnd! 55.7fF ;**FLOATING
C15 metal_1119400_3830900# gnd! 55.5fF ;**FLOATING
C16 metal_1249900_3788850# gnd! 55.5fF ;**FLOATING
C17 diff_2311300_334950# gnd! 115.8fF
C18 diff_2096700_342200# gnd! 148.4fF
C19 diff_2444700_139200# gnd! 305.9fF
C20 diff_1644300_82650# gnd! 124.9fF
C21 diff_1558750_169650# gnd! 173.1fF
C22 diff_1635600_343650# gnd! 108.0fF
C23 diff_1416650_342200# gnd! 183.4fF
C24 diff_1370250_332050# gnd! 281.2fF
C25 diff_2083650_427750# gnd! 138.0fF
C26 diff_1196250_255200# gnd! 153.0fF
C27 diff_2201100_484300# gnd! 126.4fF
C28 diff_2304050_481400# gnd! 85.9fF
C29 diff_1998100_527800# gnd! 56.9fF
C30 diff_2144550_503150# gnd! 473.9fF
C31 diff_2199650_546650# gnd! 92.4fF
C32 diff_1943000_511850# gnd! 212.4fF
C33 diff_1841500_561150# gnd! 83.5fF
C34 diff_1808150_595950# gnd! 67.2fF
C35 diff_681500_266800# gnd! 128.9fF
C36 diff_772850_316100# gnd! 628.3fF
C37 diff_1158550_546650# gnd! 124.2fF
C38 diff_651050_353800# gnd! 132.5fF
C39 diff_365400_424850# gnd! 83.0fF
C40 diff_340750_424850# gnd! 48.7fF
C41 diff_651050_437900# gnd! 132.1fF
C42 diff_1302100_537950# gnd! 233.2fF
C43 diff_1584850_569850# gnd! 1487.9fF
C44 diff_1718250_556800# gnd! 245.3fF
C45 diff_1262950_575650# gnd! 340.0fF
C46 diff_346550_482850# gnd! 125.7fF
C47 diff_292900_530700# gnd! 124.5fF
C48 diff_337850_514750# gnd! 201.5fF
C49 diff_2177900_597400# gnd! 138.5fF
C50 diff_2041600_566950# gnd! 131.2fF
C51 diff_1995200_672800# gnd! 61.5fF
C52 diff_2385250_669900# gnd! 178.8fF
C53 diff_2144550_636550# gnd! 447.1fF
C54 diff_2201100_690200# gnd! 93.2fF
C55 diff_1925600_656850# gnd! 253.1fF
C56 diff_1738550_530700# gnd! 97.3fF
C57 diff_1616750_597400# gnd! 128.9fF
C58 diff_365400_569850# gnd! 84.6fF
C59 diff_339300_571300# gnd! 50.0fF
C60 diff_1051250_593050# gnd! 1091.8fF
C61 diff_1796550_646700# gnd! 803.5fF
C62 diff_1841500_707600# gnd! 82.0fF
C63 diff_1808150_742400# gnd! 67.8fF
C64 diff_1262950_671350# gnd! 368.7fF
C65 diff_711950_652500# gnd! 189.0fF
C66 diff_346550_629300# gnd! 122.2fF
C67 diff_292900_675700# gnd! 123.8fF
C68 diff_337850_655400# gnd! 202.3fF
C69 diff_1290500_722100# gnd! 418.5fF
C70 diff_1731300_701800# gnd! 68.7fF
C71 diff_1161450_745300# gnd! 102.7fF
C72 diff_2172100_739500# gnd! 148.9fF
C73 diff_2273600_775750# gnd! 93.2fF
C74 diff_1995200_817800# gnd! 59.0fF
C75 diff_2409900_877250# gnd! 136.5fF
C76 diff_2143100_796050# gnd! 506.6fF
C77 diff_690200_720650# gnd! 215.0fF
C78 diff_594500_717750# gnd! 174.3fF
C79 diff_1744350_653950# gnd! 373.9fF
C80 diff_1051250_652500# gnd! 1304.0fF
C81 diff_1796550_791700# gnd! 139.2fF
C82 diff_2201100_846800# gnd! 92.0fF
C83 diff_2038700_881600# gnd! 144.4fF
C84 diff_527800_677150# gnd! 225.5fF
C85 diff_365400_716300# gnd! 87.5fF
C86 diff_1944450_801850# gnd! 206.5fF
C87 diff_1302100_807650# gnd! 234.1fF
C88 diff_1850200_854050# gnd! 430.0fF
C89 diff_1841500_870000# gnd! 76.5fF
C90 diff_1809600_885950# gnd! 63.7fF
C91 diff_1925600_801850# gnd! 331.2fF
C92 diff_1584850_851150# gnd! 564.9fF
C93 diff_1262950_843900# gnd! 330.0fF
C94 diff_1719700_845350# gnd! 243.3fF
C95 diff_716300_748200# gnd! 228.3fF
C96 diff_339300_716300# gnd! 48.7fF
C97 diff_597400_767050# gnd! 144.3fF
C98 diff_1608050_883050# gnd! 125.9fF
C99 diff_1740000_820700# gnd! 99.0fF
C100 diff_2172100_899000# gnd! 146.9fF
C101 diff_2314200_884500# gnd! 336.1fF
C102 diff_2275050_913500# gnd! 101.5fF
C103 diff_1996650_962800# gnd! 58.4fF
C104 diff_1925600_946850# gnd! 240.5fF
C105 diff_1262950_939600# gnd! 364.6fF
C106 diff_1090400_862750# gnd! 1207.7fF
C107 diff_1784950_914950# gnd! 505.0fF
C108 diff_1798000_938150# gnd! 127.4fF
C109 diff_2144550_958450# gnd! 346.9fF
C110 diff_2148900_1010650# gnd! 132.0fF
C111 diff_2209800_997600# gnd! 86.0fF
C112 diff_1850200_999050# gnd! 641.7fF
C113 diff_717750_555350# gnd! 577.8fF
C114 diff_346550_772850# gnd! 128.7fF
C115 diff_291450_822150# gnd! 126.1fF
C116 diff_337850_765600# gnd! 218.0fF
C117 diff_681500_891750# gnd! 161.0fF
C118 diff_849700_965700# gnd! 28.3fF
C119 diff_365400_861300# gnd! 91.3fF
C120 diff_339300_859850# gnd! 51.6fF
C121 diff_1160000_1010650# gnd! 103.9fF
C122 diff_1290500_990350# gnd! 455.7fF
C123 diff_1745800_945400# gnd! 226.6fF
C124 diff_1842950_996150# gnd! 72.3fF
C125 diff_1731300_991800# gnd! 67.3fF
C126 diff_1824100_994700# gnd! 48.5fF
C127 diff_1168700_1032400# gnd! 111.3fF
C128 diff_2122800_433550# gnd! 485.1fF
C129 diff_2272150_1090400# gnd! 111.8fF
C130 diff_2153250_1116500# gnd! 123.3fF
C131 diff_2243150_1175950# gnd! 59.4fF
C132 diff_2344650_1202050# gnd! 55.9fF
C133 diff_1352850_295800# gnd! 2190.7fF
C134 diff_2077850_1148400# gnd! 86.1fF
C135 diff_2130050_1220900# gnd! 65.4fF
C136 diff_1090400_903350# gnd! 1288.3fF
C137 diff_1448550_1090400# gnd! 276.4fF
C138 diff_1786400_1088950# gnd! 174.4fF
C139 diff_1603700_1123750# gnd! 270.9fF
C140 diff_1262950_1112150# gnd! 377.3fF
C141 diff_1436950_1083150# gnd! 358.7fF
C142 diff_1726950_1144050# gnd! 142.8fF
C143 diff_1284700_1093300# gnd! 305.9fF
C144 diff_1238300_1142600# gnd! 47.4fF
C145 diff_1590650_513300# gnd! 649.8fF
C146 diff_1612400_1041100# gnd! 269.2fF
C147 diff_2338850_1251350# gnd! 47.3fF
C148 diff_1592100_1117950# gnd! 272.9fF
C149 diff_2002450_1074450# gnd! 135.7fF
C150 diff_2206900_1222350# gnd! 191.9fF
C151 diff_2105400_1174500# gnd! 197.9fF
C152 diff_2096700_1296300# gnd! 134.5fF
C153 diff_2637550_1542800# gnd! 116.5fF
C154 diff_2324350_1402150# gnd! 66.6fF
C155 diff_2238800_1378950# gnd! 163.1fF
C156 diff_2173550_1360100# gnd! 191.2fF
C157 diff_2578100_1628350# gnd! 175.4fF
C158 diff_2269250_1429700# gnd! 255.4fF
C159 diff_2280850_1441300# gnd! 279.1fF
C160 diff_2654950_1667500# gnd! 122.4fF
C161 diff_1624000_314650# gnd! 1178.5fF
C162 diff_2108300_1347050# gnd! 229.9fF
C163 diff_1547150_726450# gnd! 624.3fF
C164 diff_1197700_311750# gnd! 499.5fF
C165 diff_1525400_1289050# gnd! 56.2fF
C166 diff_1426800_1106350# gnd! 951.3fF
C167 diff_1419550_1315150# gnd! 102.3fF
C168 diff_1113600_1132450# gnd! 154.3fF
C169 diff_1048350_1142600# gnd! 139.1fF
C170 diff_1332550_1297750# gnd! 619.8fF
C171 diff_1177400_1117950# gnd! 255.2fF
C172 diff_1349950_1289050# gnd! 84.7fF
C173 diff_1592100_1387650# gnd! 144.7fF
C174 diff_1055600_1228150# gnd! 774.6fF
C175 diff_1087500_571300# gnd! 945.4fF
C176 diff_1141150_1351400# gnd! 100.7fF
C177 diff_1305000_1400700# gnd! 411.1fF
C178 diff_1109250_1280350# gnd! 272.1fF
C179 diff_345100_925100# gnd! 128.9fF
C180 diff_495900_936700# gnd! 110.4fF
C181 diff_291450_967150# gnd! 126.4fF
C182 diff_681500_959900# gnd! 172.9fF
C183 diff_754000_974400# gnd! 106.5fF
C184 diff_803300_1059950# gnd! 45.2fF
C185 diff_751100_1103450# gnd! 98.7fF
C186 diff_713400_1139700# gnd! 179.8fF
C187 diff_582900_1045450# gnd! 50.0fF
C188 diff_365400_1023700# gnd! 87.5fF
C189 diff_339300_1022250# gnd! 50.1fF
C190 diff_546650_1088950# gnd! 87.8fF
C191 diff_577100_1051250# gnd! 80.3fF
C192 diff_709050_1219450# gnd! 126.5fF
C193 diff_345100_1081700# gnd! 124.5fF
C194 diff_291450_1128100# gnd! 126.3fF
C195 diff_336400_1125200# gnd! 214.7fF
C196 diff_564050_1106350# gnd! 252.6fF
C197 diff_1141150_1415200# gnd! 228.0fF
C198 diff_1267300_1444200# gnd! 603.1fF
C199 diff_1197700_1436950# gnd! 468.3fF
C200 diff_1057050_1325300# gnd! 178.9fF
C201 diff_725000_1268750# gnd! 32.1fF
C202 diff_706150_1268750# gnd! 31.5fF
C203 diff_710500_1136800# gnd! 338.7fF
C204 diff_667000_1268750# gnd! 28.3fF
C205 diff_733700_1262950# gnd! 168.6fF
C206 diff_598850_1270200# gnd! 66.5fF
C207 diff_365400_1168700# gnd! 87.6fF
C208 diff_337850_1168700# gnd! 53.3fF
C209 diff_617700_1270200# gnd! 65.9fF
C210 diff_655400_1313700# gnd! 202.2fF
C211 diff_1194800_1497850# gnd! 1383.8fF
C212 diff_535050_885950# gnd! 1273.8fF
C213 diff_1016450_1492050# gnd! 72.8fF
C214 diff_1048350_1547150# gnd! 68.8fF
C215 diff_345100_1226700# gnd! 121.5fF
C216 diff_291450_1273100# gnd! 124.8fF
C217 diff_787350_1442750# gnd! 52.0fF
C218 diff_661200_1406500# gnd! 138.0fF
C219 diff_767050_1451450# gnd! 34.3fF
C220 diff_365400_1315150# gnd! 89.2fF
C221 diff_337850_1312250# gnd! 51.9fF
C222 diff_345100_1370250# gnd! 118.0fF
C223 diff_290000_1419550# gnd! 121.6fF
C224 diff_336400_1363000# gnd! 222.9fF
C225 diff_785900_1464500# gnd! 182.5fF
C226 diff_630750_1461600# gnd! 26.9fF
C227 diff_552450_1347050# gnd! 609.2fF
C228 diff_526350_1077350# gnd! 429.9fF
C229 diff_677150_1461600# gnd! 69.5fF
C230 diff_733700_1481900# gnd! 105.2fF
C231 diff_1015000_1583400# gnd! 61.9fF
C232 diff_810550_1503650# gnd! 51.1fF
C233 diff_846800_1510900# gnd! 62.8fF
C234 diff_858400_1561650# gnd! 44.8fF
C235 diff_345100_1497850# gnd! 123.3fF
C236 diff_559700_1464500# gnd! 76.5fF
C237 diff_497350_1464500# gnd! 391.2fF
C238 diff_781550_1535550# gnd! 139.3fF
C239 diff_896100_1570350# gnd! 164.3fF
C240 diff_1232500_1610950# gnd! 650.8fF
C241 diff_667000_980200# gnd! 1381.4fF
C242 diff_2150350_1422450# gnd! 333.0fF
C243 diff_1016450_1635600# gnd! 71.1fF
C244 diff_1080250_1657350# gnd! 786.4fF
C245 diff_925100_1455800# gnd! 830.8fF
C246 diff_2085100_1422450# gnd! 340.2fF
C247 diff_2215600_1422450# gnd! 361.8fF
C248 diff_2041600_1738550# gnd! 42.8fF
C249 diff_935250_1697950# gnd! 138.4fF
C250 diff_871450_1602250# gnd! 858.2fF
C251 diff_916400_1668950# gnd! 130.3fF
C252 diff_852600_1702300# gnd! 280.1fF
C253 diff_336400_1510900# gnd! 218.4fF
C254 diff_519100_1629800# gnd! 427.8fF
C255 diff_797500_1693600# gnd! 110.3fF
C256 diff_633650_1644300# gnd! 49.1fF
C257 diff_332050_1580500# gnd! 131.1fF
C258 diff_314650_1616750# gnd! 83.3fF
C259 diff_371200_1631250# gnd! 118.0fF
C260 diff_362500_1632700# gnd! 213.5fF
C261 diff_640900_1654450# gnd! 57.4fF
C262 diff_681500_1692150# gnd! 112.3fF
C263 diff_733700_1700850# gnd! 171.4fF
C264 diff_2218500_1796550# gnd! 25.5fF
C265 diff_2179350_1790750# gnd! 65.8fF
C266 diff_2157600_1809600# gnd! 78.6fF
C267 diff_1925600_1133900# gnd! 435.2fF
C268 diff_846800_1278900# gnd! 1047.7fF
C269 diff_1999550_1331100# gnd! 830.1fF
C270 diff_2295350_1931400# gnd! 84.1fF
C271 diff_2153250_1957500# gnd! 307.7fF
C272 diff_1400700_1510900# gnd! 388.7fF
C273 diff_1286150_1331100# gnd! 320.9fF
C274 diff_740950_1709550# gnd! 34.3fF
C275 diff_674250_1700850# gnd! 56.9fF
C276 diff_826500_1682000# gnd! 85.8fF
C277 diff_668450_1715350# gnd! 34.2fF
C278 diff_740950_1728400# gnd! 35.8fF
C279 diff_497350_1687800# gnd! 241.7fF
C280 diff_688750_1509450# gnd! 277.0fF
C281 diff_903350_1763200# gnd! 35.6fF
C282 diff_1025150_1793650# gnd! 82.3fF
C283 diff_665550_1548600# gnd! 937.5fF
C284 diff_526350_1657350# gnd! 75.8fF
C285 diff_797500_1757400# gnd! 1240.2fF
C286 diff_601750_1919800# gnd! 21.6fF
C287 diff_529250_1925600# gnd! 87.1fF
C288 diff_2035800_1877750# gnd! 442.1fF
C289 diff_2153250_1870500# gnd! 399.8fF
C290 diff_2518650_2030000# gnd! 101.7fF
C291 diff_2447600_1993750# gnd! 165.9fF
C292 diff_2382350_1993750# gnd! 207.1fF
C293 diff_2317100_1996650# gnd! 236.1fF
C294 diff_2534600_2179350# gnd! 162.4fF
C295 diff_2201100_2086550# gnd! 286.2fF
C296 diff_2208350_2030000# gnd! 327.3fF
C297 diff_620600_1919800# gnd! 199.7fF
C298 diff_2093800_1972000# gnd! 508.3fF
C299 diff_636550_1956050# gnd! 47.6fF
C300 diff_629300_1979250# gnd! 84.6fF
C301 diff_677150_1960400# gnd! 173.3fF
C302 diff_703250_1961850# gnd! 197.5fF
C303 diff_1149850_1992300# gnd! 286.5fF
C304 diff_2505600_2241700# gnd! 89.9fF
C305 diff_2459200_2230100# gnd! 22.9fF
C306 diff_2505600_2260550# gnd! 33.7fF
C307 diff_2505600_2279400# gnd! 38.4fF
C308 diff_2360600_2244600# gnd! 31.7fF
C309 diff_2379450_2250400# gnd! 122.4fF
C310 diff_791700_1716800# gnd! 383.8fF
C311 diff_842450_2070600# gnd! 1286.3fF
C312 diff_569850_2003900# gnd! 172.8fF
C313 diff_1181750_1322400# gnd! 645.4fF
C314 diff_2495450_2354800# gnd! 29.6fF
C315 diff_2161950_1146950# gnd! 1160.7fF
C316 diff_2430200_2244600# gnd! 123.2fF
C317 diff_2485300_2375100# gnd! 37.2fF
C318 diff_2485300_2392500# gnd! 93.4fF
C319 diff_2335950_2264900# gnd! 136.9fF
C320 diff_2179350_2344650# gnd! 56.2fF
C321 diff_2218500_2198200# gnd! 302.6fF
C322 diff_2172100_2192400# gnd! 318.8fF
C323 diff_2176450_2302600# gnd! 215.5fF
C324 diff_2127150_2344650# gnd! 80.8fF
C325 diff_2064800_2330150# gnd! 24.9fF
C326 diff_2045950_2335950# gnd! 59.6fF
C327 diff_1979250_2237350# gnd! 24.9fF
C328 diff_1932850_2225750# gnd! 36.5fF
C329 diff_1077350_1464500# gnd! 672.2fF
C330 diff_1998100_2237350# gnd! 84.1fF
C331 diff_1979250_2308400# gnd! 24.9fF
C332 diff_1932850_2308400# gnd! 25.9fF
C333 diff_1712450_2234450# gnd! 219.5fF
C334 diff_991800_1986500# gnd! 382.9fF
C335 diff_1754500_2189500# gnd! 82.3fF
C336 diff_1796550_2237350# gnd! 128.8fF
C337 diff_1732750_2256200# gnd! 97.0fF
C338 diff_1850200_2308400# gnd! 92.4fF
C339 diff_1914000_2251850# gnd! 86.1fF
C340 diff_2108300_2347550# gnd! 67.9fF
C341 diff_1811050_2224300# gnd! 241.3fF
C342 diff_1850200_2324350# gnd! 29.6fF
C343 diff_1732750_2273600# gnd! 81.1fF
C344 diff_1638500_2351900# gnd! 47.4fF
C345 diff_1571800_2293900# gnd! 48.6fF
C346 diff_1080250_1561650# gnd! 1828.5fF
C347 diff_1552950_2298250# gnd! 97.2fF
C348 diff_1638500_2367850# gnd! 169.5fF
C349 diff_2404100_2504150# gnd! 80.9fF
C350 diff_2314200_2449050# gnd! 151.0fF
C351 diff_2192400_2495450# gnd! 149.7fF
C352 diff_2201100_2537500# gnd! 141.2fF
C353 diff_2179350_2360600# gnd! 282.7fF
C354 diff_2322900_2508500# gnd! 453.1fF
C355 diff_2427300_2585350# gnd! 32.4fF
C356 diff_1892250_2309850# gnd! 227.8fF
C357 diff_1492050_2322900# gnd! 24.9fF
C358 diff_1023700_2198200# gnd! 28.3fF
C359 diff_1429700_2322900# gnd! 21.4fF
C360 diff_1470300_2340300# gnd! 29.7fF
C361 diff_1452900_2244600# gnd! 439.7fF
C362 diff_1660250_2388150# gnd! 122.4fF
C363 diff_1706650_2405550# gnd! 106.3fF
C364 diff_2063350_2495450# gnd! 141.0fF
C365 diff_1969100_2514300# gnd! 262.7fF
C366 diff_2021300_2420050# gnd! 172.7fF
C367 diff_2108300_2408450# gnd! 199.6fF
C368 diff_2373650_2621600# gnd! 51.7fF
C369 diff_2280850_2602750# gnd! 246.0fF
C370 diff_2209800_2586800# gnd! 35.7fF
C371 diff_2201100_2576650# gnd! 65.7fF
C372 diff_2212700_2604200# gnd! 256.0fF
C373 diff_2275050_2614350# gnd! 124.6fF
C374 diff_2134400_2586800# gnd! 32.2fF
C375 diff_1448550_2322900# gnd! 126.6fF
C376 diff_1392000_2341750# gnd! 91.7fF
C377 diff_1336900_2322900# gnd! 29.7fF
C378 diff_1318050_2322900# gnd! 29.6fF
C379 diff_1094750_2248950# gnd! 21.6fF
C380 diff_1023700_2217050# gnd! 198.3fF
C381 diff_1003400_2257650# gnd! 101.3fF
C382 diff_867100_2254750# gnd! 21.6fF
C383 diff_865650_2222850# gnd! 111.4fF
C384 diff_1270200_2417150# gnd! 29.0fF
C385 diff_1023700_2175000# gnd! 359.6fF
C386 diff_1289050_2415700# gnd! 38.2fF
C387 diff_1915450_2589700# gnd! 32.6fF
C388 diff_1840050_2588250# gnd! 32.4fF
C389 diff_2117000_2625950# gnd! 77.1fF
C390 diff_2079300_2623050# gnd! 50.8fF
C391 diff_1325300_2459200# gnd! 303.3fF
C392 diff_1075900_2275050# gnd! 934.8fF
C393 diff_1500750_2386700# gnd! 112.6fF
C394 diff_1402150_2514300# gnd! 30.2fF
C395 diff_1390550_2521550# gnd! 61.1fF
C396 diff_1239750_2443250# gnd! 126.7fF
C397 diff_1355750_2514300# gnd! 30.3fF
C398 diff_1908200_2576650# gnd! 70.0fF
C399 diff_1626900_2588250# gnd! 32.2fF
C400 diff_1987950_2604200# gnd! 394.6fF
C401 diff_1919800_2605650# gnd! 477.1fF
C402 diff_1790750_2624500# gnd! 50.2fF
C403 diff_1610950_2605650# gnd! 303.6fF
C404 diff_1619650_2578100# gnd! 67.8fF
C405 diff_1629800_2623050# gnd! 476.0fF
C406 diff_1336900_2549100# gnd! 51.7fF
C407 diff_1415200_2605650# gnd! 68.1fF
C408 diff_1097650_2396850# gnd! 170.1fF
C409 diff_872900_2288100# gnd! 364.0fF
C410 diff_532150_2082200# gnd! 166.9fF
C411 diff_595950_2080750# gnd! 117.5fF
C412 diff_680050_2190950# gnd! 32.3fF
C413 diff_614800_2167750# gnd! 223.6fF
C414 diff_633650_2205450# gnd! 38.1fF
C415 diff_569850_2193850# gnd! 33.6fF
C416 diff_551000_2193850# gnd! 34.3fF
C417 diff_537950_1786400# gnd! 616.1fF
C418 diff_884500_2331600# gnd! 86.8fF
C419 diff_894650_2441800# gnd! 45.3fF
C420 diff_784450_2395400# gnd! 159.0fF
C421 diff_807650_2418600# gnd! 62.8fF
C422 diff_907700_2450500# gnd! 185.8fF
C423 diff_935250_2476600# gnd! 97.5fF
C424 diff_1158550_2475150# gnd! 153.5fF
C425 diff_1120850_2447600# gnd! 87.1fF
C426 diff_1046900_2517200# gnd! 113.0fF
C427 diff_855500_2512850# gnd! 59.9fF
C428 diff_855500_2492550# gnd! 312.0fF
C429 diff_633650_2347550# gnd! 29.6fF
C430 diff_595950_2349000# gnd! 28.3fF
C431 diff_549550_2349000# gnd! 29.4fF
C432 diff_529250_2347550# gnd! 33.7fF
C433 diff_622050_2318550# gnd! 893.8fF
C434 diff_640900_2343200# gnd! 371.6fF
C435 diff_537950_2248950# gnd! 969.6fF
C436 diff_614800_2349000# gnd! 90.6fF
C437 diff_595950_2407000# gnd! 29.6fF
C438 diff_568400_2407000# gnd! 57.8fF
C439 diff_774300_2469350# gnd! 77.3fF
C440 diff_552450_2137300# gnd! 252.7fF
C441 diff_974400_2502700# gnd! 124.8fF
C442 diff_682950_2483850# gnd! 139.0fF
C443 diff_688750_2531700# gnd! 351.0fF
C444 diff_1200600_2607100# gnd! 253.2fF
C445 diff_1982150_2614350# gnd! 131.0fF
C446 diff_1699400_2604200# gnd! 270.2fF
C447 diff_1693600_2615800# gnd! 125.8fF
C448 diff_1668950_2660750# gnd! 715.6fF
C449 diff_2282300_2737600# gnd! 828.2fF
C450 diff_2061900_2756450# gnd! 172.9fF
C451 diff_1945900_2772400# gnd! 175.9fF
C452 diff_1886450_2740500# gnd! 174.3fF
C453 diff_1832800_2763700# gnd! 174.5fF
C454 diff_1773350_2733250# gnd! 173.6fF
C455 diff_1613850_2688300# gnd! 494.1fF
C456 diff_1402150_2665100# gnd! 30.0fF
C457 diff_1058500_2582450# gnd! 168.8fF
C458 diff_1355750_2662200# gnd! 31.2fF
C459 diff_999050_2583900# gnd! 167.6fF
C460 diff_943950_2649150# gnd! 169.4fF
C461 diff_884500_2589700# gnd! 174.8fF
C462 diff_1007750_2685400# gnd! 208.0fF
C463 diff_1390550_2670900# gnd! 64.2fF
C464 diff_1336900_2698450# gnd! 53.2fF
C465 diff_904800_2683950# gnd! 202.1fF
C466 diff_204450_2418600# gnd! 106.8fF
C467 diff_265350_2463550# gnd! 42.9fF
C468 diff_230550_2438900# gnd! 75.7fF
C469 diff_249400_1373150# gnd! 5802.4fF
C470 diff_368300_2570850# gnd! 244.5fF
C471 diff_423400_2592600# gnd! 177.1fF
C472 diff_1331100_2717300# gnd! 650.3fF
C473 diff_1415200_2753550# gnd! 68.2fF
C474 diff_1200600_2627400# gnd! 254.3fF
C475 diff_1329650_2521550# gnd! 445.2fF
C476 diff_1329650_2769500# gnd! 206.1fF
C477 diff_1719700_2741950# gnd! 173.6fF
C478 diff_1660250_2731800# gnd! 176.9fF
C479 diff_1729850_2853600# gnd! 373.6fF
C480 diff_468350_2653500# gnd! 164.6fF
C481 diff_250850_2582450# gnd! 125.3fF
C482 diff_282750_2514300# gnd! 210.8fF
C483 diff_275500_2569400# gnd! 141.3fF
C484 diff_703250_2691200# gnd! 51.8fF
C485 diff_794600_2701350# gnd! 53.1fF
C486 diff_749650_2701350# gnd! 51.4fF
C487 diff_1402150_2830400# gnd! 30.8fF
C488 diff_1983600_2676700# gnd! 382.6fF
C489 diff_1390550_2837650# gnd! 62.9fF
C490 diff_1355750_2828950# gnd! 31.3fF
C491 diff_1004850_2637550# gnd! 256.9fF
C492 diff_1336900_2865200# gnd! 52.1fF
C493 diff_1789300_2900000# gnd! 148.5fF
C494 diff_1668950_2924650# gnd! 411.6fF
C495 diff_2215600_2913050# gnd! 284.2fF
C496 diff_839550_2504150# gnd! 506.0fF
C497 diff_417600_2791250# gnd! 127.1fF
C498 diff_772850_2547650# gnd! 716.8fF
C499 diff_938150_2853600# gnd! 272.0fF
C500 diff_880150_2855050# gnd! 281.7fF
C501 diff_938150_2881150# gnd! 123.2fF
C502 diff_867100_2815900# gnd! 152.0fF
C503 diff_501700_2402650# gnd! 487.1fF
C504 diff_1415200_2920300# gnd! 67.9fF
C505 diff_1136800_2604200# gnd! 332.8fF
C506 diff_1552950_2940600# gnd! 133.3fF
C507 diff_2002450_2731800# gnd! 513.3fF
C508 diff_2134400_3091400# gnd! 139.6fF
C509 diff_1552950_2965250# gnd! 135.4fF
C510 diff_1947350_2814450# gnd! 324.9fF
C511 diff_1893700_2785450# gnd! 328.1fF
C512 diff_1402150_2984100# gnd! 30.9fF
C513 diff_1355750_2985550# gnd! 30.5fF
C514 diff_1390550_2979750# gnd! 72.0fF
C515 diff_1336900_3020350# gnd! 59.7fF
C516 diff_1135350_2940600# gnd! 23.8fF
C517 diff_1044000_2936250# gnd! 24.2fF
C518 diff_999050_2946400# gnd! 25.8fF
C519 diff_1113600_2972500# gnd! 39.2fF
C520 diff_1051250_2936250# gnd! 38.9fF
C521 diff_907700_2937700# gnd! 23.3fF
C522 diff_477050_2791250# gnd! 64.3fF
C523 diff_387150_2801400# gnd! 142.3fF
C524 diff_490100_2813000# gnd! 66.9fF
C525 diff_536500_2711500# gnd! 397.5fF
C526 diff_258100_549550# gnd! 3198.4fF
C527 diff_258100_694550# gnd! 3262.7fF
C528 diff_423400_2781100# gnd! 113.6fF
C529 diff_477050_2855050# gnd! 54.4fF
C530 diff_136300_2602750# gnd! 2988.4fF
C531 diff_978750_2972500# gnd! 37.6fF
C532 diff_916400_2936250# gnd! 37.4fF
C533 diff_1135350_3008750# gnd! 22.6fF
C534 diff_1113600_2989900# gnd! 39.1fF
C535 diff_1270200_2518650# gnd! 633.8fF
C536 diff_1687800_3033400# gnd! 1067.8fF
C537 diff_1782050_3013100# gnd! 136.1fF
C538 diff_1711000_3092850# gnd! 137.0fF
C539 diff_1415200_3075450# gnd! 69.3fF
C540 diff_1136800_2630300# gnd! 372.5fF
C541 diff_1629800_3060950# gnd! 153.4fF
C542 diff_1613850_2840550# gnd! 3633.5fF
C543 diff_2169200_3155200# gnd! 20.0fF
C544 diff_2079300_3149400# gnd! 22.5fF
C545 diff_2034350_3163900# gnd! 21.5fF
C546 diff_2148900_3184200# gnd! 44.1fF
C547 diff_2086550_3147950# gnd! 40.6fF
C548 diff_1943000_3149400# gnd! 24.9fF
C549 diff_1899500_3155200# gnd! 24.8fF
C550 diff_2014050_3185650# gnd! 39.9fF
C551 diff_1951700_3147950# gnd! 38.1fF
C552 diff_2169200_3220450# gnd! 22.9fF
C553 diff_2148900_3203050# gnd! 40.8fF
C554 diff_2169200_3262500# gnd! 19.6fF
C555 diff_2077850_3240750# gnd! 21.8fF
C556 diff_2034350_3220450# gnd! 22.9fF
C557 diff_1808150_3149400# gnd! 25.5fF
C558 diff_1764650_3155200# gnd! 24.6fF
C559 diff_1329650_2830400# gnd! 473.1fF
C560 diff_1326750_3091400# gnd! 214.9fF
C561 diff_1879200_3185650# gnd! 38.0fF
C562 diff_1816850_3147950# gnd! 37.2fF
C563 diff_2085100_3242200# gnd! 40.2fF
C564 diff_2014050_3203050# gnd! 38.9fF
C565 diff_1951700_3203050# gnd! 38.8fF
C566 diff_1943000_3239300# gnd! 22.2fF
C567 diff_1899500_3221900# gnd! 23.2fF
C568 diff_1673300_3150850# gnd! 22.6fF
C569 diff_1742900_3185650# gnd! 38.3fF
C570 diff_1680550_3149400# gnd! 38.6fF
C571 diff_1879200_3203050# gnd! 38.1fF
C572 diff_2077850_3256700# gnd! 22.5fF
C573 diff_2034350_3262500# gnd! 22.5fF
C574 diff_2148900_3292950# gnd! 40.8fF
C575 diff_2086550_3255250# gnd! 38.8fF
C576 diff_1943000_3256700# gnd! 24.8fF
C577 diff_1899500_3262500# gnd! 23.9fF
C578 diff_1808150_3240750# gnd! 23.3fF
C579 diff_1764650_3221900# gnd! 23.3fF
C580 diff_1815400_3242200# gnd! 41.4fF
C581 diff_2014050_3292950# gnd! 38.6fF
C582 diff_1950250_3256700# gnd! 38.1fF
C583 diff_2169200_3327750# gnd! 20.3fF
C584 diff_2148900_3310350# gnd! 40.8fF
C585 diff_2169200_3368350# gnd! 19.0fF
C586 diff_2077850_3346600# gnd! 24.5fF
C587 diff_2034350_3329200# gnd! 21.7fF
C588 diff_2086550_3310350# gnd! 36.5fF
C589 diff_1742900_3204500# gnd! 36.7fF
C590 diff_1808150_3258150# gnd! 24.5fF
C591 diff_1764650_3262500# gnd! 23.0fF
C592 diff_1673300_3240750# gnd! 22.6fF
C593 diff_1135350_3047900# gnd! 23.3fF
C594 diff_1044000_3024700# gnd! 22.7fF
C595 diff_1000500_3008750# gnd! 22.6fF
C596 diff_1051250_3029050# gnd! 39.9fF
C597 diff_978750_2989900# gnd! 38.2fF
C598 diff_907700_3027600# gnd! 23.5fF
C599 diff_488650_2876800# gnd! 73.3fF
C600 diff_655400_2966700# gnd! 411.2fF
C601 diff_916400_3029050# gnd! 38.3fF
C602 diff_999050_3049350# gnd! 24.7fF
C603 diff_1044000_3043550# gnd! 24.4fF
C604 diff_1113600_3079800# gnd! 38.9fF
C605 diff_1051250_3043550# gnd! 37.9fF
C606 diff_907700_3043550# gnd! 24.8fF
C607 diff_978750_3079800# gnd! 37.3fF
C608 diff_1135350_3116050# gnd! 23.9fF
C609 diff_916400_3043550# gnd! 38.1fF
C610 diff_1113600_3097200# gnd! 38.4fF
C611 diff_1680550_3242200# gnd! 39.9fF
C612 diff_1879200_3292950# gnd! 38.1fF
C613 diff_1816850_3255250# gnd! 38.6fF
C614 diff_2014050_3310350# gnd! 38.5fF
C615 diff_1943000_3346600# gnd! 23.1fF
C616 diff_1899500_3329200# gnd! 22.6fF
C617 diff_1950250_3349500# gnd! 37.6fF
C618 diff_1673300_3258150# gnd! 22.8fF
C619 diff_1742900_3292950# gnd! 38.6fF
C620 diff_1680550_3256700# gnd! 38.6fF
C621 diff_1877750_3314700# gnd! 37.8fF
C622 diff_2077850_3364000# gnd! 24.3fF
C623 diff_2034350_3369800# gnd! 20.2fF
C624 diff_2148900_3398800# gnd! 44.2fF
C625 diff_2086550_3362550# gnd! 38.1fF
C626 diff_2169200_3435050# gnd! 19.5fF
C627 diff_1943000_3364000# gnd! 24.5fF
C628 diff_1899500_3369800# gnd! 22.1fF
C629 diff_1808150_3346600# gnd! 22.7fF
C630 diff_1764650_3329200# gnd! 23.0fF
C631 diff_1815400_3348050# gnd! 37.1fF
C632 diff_1742900_3310350# gnd! 39.8fF
C633 diff_2012600_3400250# gnd! 39.5fF
C634 diff_1950250_3362550# gnd! 36.6fF
C635 diff_2148900_3417650# gnd! 41.6fF
C636 diff_1808150_3364000# gnd! 23.9fF
C637 diff_1673300_3346600# gnd! 22.6fF
C638 diff_1680550_3348050# gnd! 37.3fF
C639 diff_1763200_3387200# gnd! 23.1fF
C640 diff_1877750_3400250# gnd! 39.3fF
C641 diff_1815400_3362550# gnd! 36.9fF
C642 diff_2077850_3453900# gnd! 23.8fF
C643 diff_2169200_3475650# gnd! 18.6fF
C644 diff_2086550_3417650# gnd! 36.6fF
C645 diff_2034350_3435050# gnd! 20.3fF
C646 diff_2012600_3417650# gnd! 40.2fF
C647 diff_2077850_3471300# gnd! 23.9fF
C648 diff_2034350_3475650# gnd! 19.1fF
C649 diff_1943000_3453900# gnd! 24.0fF
C650 diff_1671850_3366900# gnd! 23.0fF
C651 diff_1742900_3400250# gnd! 38.3fF
C652 diff_1680550_3362550# gnd! 38.1fF
C653 diff_1898050_3435050# gnd! 24.1fF
C654 diff_1950250_3456800# gnd! 36.3fF
C655 diff_1877750_3417650# gnd! 38.6fF
C656 diff_2086550_3468400# gnd! 39.8fF
C657 diff_2106850_3184200# gnd! 329.3fF
C658 diff_1806700_3456800# gnd! 24.0fF
C659 diff_1763200_3436500# gnd! 24.4fF
C660 diff_1815400_3456800# gnd! 37.9fF
C661 diff_1943000_3471300# gnd! 23.1fF
C662 diff_1899500_3477100# gnd! 19.8fF
C663 diff_2012600_3507550# gnd! 42.1fF
C664 diff_1950250_3469850# gnd! 36.9fF
C665 diff_2169200_3542350# gnd! 18.7fF
C666 diff_2148900_3524950# gnd! 41.1fF
C667 diff_2083650_3562650# gnd! 41.8fF
C668 diff_2077850_3561200# gnd! 19.6fF
C669 diff_2034350_3542350# gnd! 19.6fF
C670 diff_2166300_3074000# gnd! 348.8fF
C671 diff_1742900_3417650# gnd! 37.7fF
C672 diff_1806700_3472750# gnd! 23.1fF
C673 diff_1763200_3478550# gnd! 23.5fF
C674 diff_1671850_3456800# gnd! 22.9fF
C675 diff_1328200_3190000# gnd! 374.5fF
C676 diff_1044000_3132000# gnd! 25.3fF
C677 diff_999050_3120400# gnd! 26.1fF
C678 diff_1051250_3136350# gnd! 37.3fF
C679 diff_978750_3097200# gnd! 37.3fF
C680 diff_1135350_3156650# gnd! 22.9fF
C681 diff_1044000_3150850# gnd! 25.8fF
C682 diff_907700_3136350# gnd! 22.7fF
C683 diff_916400_3134900# gnd! 38.5fF
C684 diff_999050_3156650# gnd! 27.5fF
C685 diff_1113600_3187100# gnd! 39.6fF
C686 diff_1051250_3150850# gnd! 38.2fF
C687 diff_907700_3150850# gnd! 24.9fF
C688 diff_978750_3187100# gnd! 35.2fF
C689 diff_916400_3150850# gnd! 37.7fF
C690 diff_1135350_3221900# gnd! 24.4fF
C691 diff_1113600_3204500# gnd! 39.0fF
C692 diff_1135350_3263950# gnd! 24.5fF
C693 diff_1042550_3242200# gnd! 25.3fF
C694 diff_999050_3223350# gnd! 26.1fF
C695 diff_1051250_3243650# gnd! 38.5fF
C696 diff_978750_3204500# gnd! 35.6fF
C697 diff_1044000_3258150# gnd! 26.9fF
C698 diff_1000500_3261050# gnd! 24.8fF
C699 diff_916400_3243650# gnd! 39.0fF
C700 diff_907700_3243650# gnd! 22.6fF
C701 diff_1113600_3294400# gnd! 38.5fF
C702 diff_1051250_3258150# gnd! 36.4fF
C703 diff_907700_3258150# gnd! 24.1fF
C704 diff_978750_3294400# gnd! 37.7fF
C705 diff_916400_3258150# gnd! 39.4fF
C706 diff_1135350_3330650# gnd! 24.0fF
C707 diff_1113600_3311800# gnd! 38.0fF
C708 diff_1679100_3456800# gnd! 38.8fF
C709 diff_1877750_3507550# gnd! 40.2fF
C710 diff_1815400_3469850# gnd! 37.7fF
C711 diff_1671850_3471300# gnd! 24.6fF
C712 diff_1742900_3507550# gnd! 39.6fF
C713 diff_1679100_3471300# gnd! 38.1fF
C714 diff_1858900_3075450# gnd! 314.1fF
C715 diff_1829900_3075450# gnd! 314.9fF
C716 diff_1718250_3075450# gnd! 313.5fF
C717 diff_1687800_3075450# gnd! 316.5fF
C718 diff_2012600_3524950# gnd! 42.8fF
C719 diff_2025650_3074000# gnd! 334.4fF
C720 diff_1943000_3564100# gnd! 19.9fF
C721 diff_1899500_3543800# gnd! 18.8fF
C722 diff_1948800_3562650# gnd! 40.2fF
C723 diff_1877750_3524950# gnd! 42.0fF
C724 diff_1808150_3561200# gnd! 23.2fF
C725 diff_1764650_3543800# gnd! 19.5fF
C726 diff_1815400_3526400# gnd! 38.6fF
C727 diff_1742900_3524950# gnd! 41.4fF
C728 diff_1673300_3561200# gnd! 20.3fF
C729 diff_1135350_3372700# gnd! 25.2fF
C730 diff_1044000_3346600# gnd! 25.4fF
C731 diff_1000500_3330650# gnd! 23.1fF
C732 diff_1051250_3350950# gnd! 37.9fF
C733 diff_978750_3311800# gnd! 38.6fF
C734 diff_1425350_3394450# gnd! 490.7fF
C735 diff_1044000_3365450# gnd! 26.7fF
C736 diff_999050_3374150# gnd! 24.6fF
C737 diff_916400_3350950# gnd! 40.3fF
C738 diff_909150_3349500# gnd! 21.7fF
C739 diff_1115050_3401700# gnd! 38.2fF
C740 diff_1051250_3365450# gnd! 36.5fF
C741 diff_907700_3365450# gnd! 24.3fF
C742 diff_978750_3401700# gnd! 37.5fF
C743 diff_916400_3365450# gnd! 39.8fF
C744 diff_1135350_3436500# gnd! 25.3fF
C745 diff_1115050_3419100# gnd! 36.9fF
C746 diff_1135350_3480000# gnd! 24.4fF
C747 diff_1044000_3456800# gnd! 26.1fF
C748 diff_1000500_3436500# gnd! 25.4fF
C749 diff_1052700_3456800# gnd! 37.4fF
C750 diff_1423900_3514800# gnd! 513.1fF
C751 diff_1489150_3117500# gnd! 729.8fF
C752 diff_1425350_3181300# gnd! 12502.5fF
C753 diff_2072050_2521550# gnd! 808.1fF
C754 diff_978750_3419100# gnd! 37.4fF
C755 diff_1044000_3472750# gnd! 26.9fF
C756 diff_1000500_3474200# gnd! 25.7fF
C757 diff_909150_3456800# gnd! 22.0fF
C758 diff_916400_3459700# gnd! 41.2fF
C759 diff_1115050_3509000# gnd! 38.8fF
C760 diff_1051250_3474200# gnd! 37.5fF
C761 diff_907700_3474200# gnd! 24.0fF
C762 diff_978750_3509000# gnd! 37.9fF
C763 diff_916400_3472750# gnd! 40.7fF
C764 diff_943950_2878250# gnd! 441.0fF
C765 diff_914950_2865200# gnd! 437.4fF
C766 diff_1135350_3543800# gnd! 24.6fF
C767 diff_1048350_2488200# gnd! 889.7fF
C768 diff_1115050_3526400# gnd! 34.7fF
C769 diff_1044000_3564100# gnd! 20.4fF
C770 diff_1000500_3543800# gnd! 24.0fF
C771 diff_1051250_3567000# gnd! 41.8fF
C772 diff_978750_3526400# gnd! 35.4fF
C773 diff_1032400_2863750# gnd! 437.6fF
C774 diff_342200_2886950# gnd! 195.8fF
C775 diff_507500_2950750# gnd! 488.9fF
C776 diff_436450_2937700# gnd! 149.2fF
C777 diff_491550_2995700# gnd! 120.2fF
C778 diff_323350_3071100# gnd! 212.2fF
C779 diff_298700_3069650# gnd! 184.2fF
C780 diff_292900_3079800# gnd! 304.0fF
C781 diff_655400_3188550# gnd! 403.5fF
C782 diff_655400_3288600# gnd! 401.9fF
C783 diff_727900_2842000# gnd! 476.2fF
C784 diff_359600_3089950# gnd! 17.5fF
C785 diff_323350_3089950# gnd! 22.9fF
C786 diff_298700_3089950# gnd! 13.5fF
C787 diff_491550_3187100# gnd! 117.4fF
C788 diff_507500_3229150# gnd! 483.0fF
C789 diff_378450_3143600# gnd! 275.4fF
C790 diff_442250_3204500# gnd! 140.5fF
C791 diff_507500_3274100# gnd! 490.1fF
C792 diff_361050_3108800# gnd! 252.9fF
C793 diff_493000_3316150# gnd! 120.9fF
C794 diff_50750_3136350# gnd! 1162.3fF
C795 diff_323350_3108800# gnd! 164.9fF
C796 diff_298700_3108800# gnd! 193.2fF
C797 diff_329150_3371250# gnd! 283.1fF
C798 diff_333500_3384300# gnd! 141.9fF
C799 diff_493000_3507550# gnd! 127.7fF
C800 diff_784450_2863750# gnd! 303.0fF
C801 diff_629300_2881150# gnd! 362.7fF
C802 diff_606100_2879700# gnd! 2911.6fF
C803 diff_507500_3552500# gnd! 504.8fF
C804 diff_909150_3567000# gnd! 22.6fF
C805 diff_916400_3567000# gnd! 41.8fF
C806 diff_887400_2863750# gnd! 446.8fF
C807 diff_627850_2752100# gnd! 2064.9fF
C808 diff_622050_2844900# gnd! 6682.6fF
C809 diff_345100_3549600# gnd! 284.4fF
C810 diff_443700_3526400# gnd! 137.1fF
C811 diff_320450_2669450# gnd! 1099.5fF
C812 test gnd! 1561.7fF
C813 reset gnd! 1482.3fF
