`include "common.h"

module chip_4004(
  input eclk, ereset,
  input clk1,
  input clk2,
  output sync,
  input reset,
  input test,
  input d0_i,
  output d0_o,
  output d0_t,
  input d1_i,
  output d1_o,
  output d1_t,
  input d2_i,
  output d2_o,
  output d2_t,
  input d3_i,
  output d3_o,
  output d3_t,
  output cm_rom,
  output cm_ram3,
  output cm_ram2,
  output cm_ram1,
  output cm_ram0
);

  function v;   // convert an analog node value to 2-level
  input [`W-1:0] x;
  begin
    v = ~x[`W-1];
  end
  endfunction

  function [`W-1:0] a;   // convert a 2-level node value to analog
  input x;
  begin
    a = x ? `HI2 : `LO2;
  end
  endfunction

  wire signed [`W-1:0] N0556_port_2, N0556_port_1, N0556_v;
  wire signed [`W-1:0] S00819_port_0, S00819_v;
  wire signed [`W-1:0] CY_ADA_port_3, CY_ADA_port_4, CY_ADA_v;
  wire signed [`W-1:0] N0449_port_1, N0449_port_7, N0449_v;
  wire signed [`W-1:0] N0440_port_6, N0440_port_5, N0440_v;
  wire signed [`W-1:0] N0444_port_12, N0444_port_13, N0444_v;
  wire signed [`W-1:0] N0883_port_0, N0883_port_10, N0883_port_19, N0883_v;
  wire signed [`W-1:0] N0880_port_0, N0880_port_10, N0880_port_19, N0880_v;
  wire signed [`W-1:0] N0887_port_3, N0887_port_5, N0887_v;
  wire signed [`W-1:0] N0530_port_4, N0530_port_5, N0530_v;
  wire signed [`W-1:0] S00579_port_1, S00579_v;
  wire signed [`W-1:0] S00578_port_1, S00578_v;
  wire signed [`W-1:0] N0939_port_3, N0939_port_4, N0939_v;
  wire signed [`W-1:0] S00757_port_1, S00757_v;
  wire signed [`W-1:0] S00817_port_0, S00817_v;
  wire signed [`W-1:0] SUB_GROUP_6__port_1, SUB_GROUP_6__port_12, SUB_GROUP_6__v;
  wire signed [`W-1:0] N0332_port_5, N0332_port_11, N0332_v;
  wire signed [`W-1:0] _TMP_1_port_2, _TMP_1_port_0, _TMP_1_port_1, _TMP_1_v;
  wire signed [`W-1:0] _TMP_0_port_2, _TMP_0_port_0, _TMP_0_port_1, _TMP_0_v;
  wire signed [`W-1:0] _TMP_3_port_2, _TMP_3_port_0, _TMP_3_port_1, _TMP_3_v;
  wire signed [`W-1:0] _TMP_2_port_2, _TMP_2_port_0, _TMP_2_port_1, _TMP_2_v;
  wire signed [`W-1:0] TMP_3_port_2, TMP_3_port_0, TMP_3_port_1, TMP_3_v;
  wire signed [`W-1:0] TMP_2_port_2, TMP_2_port_0, TMP_2_port_1, TMP_2_v;
  wire signed [`W-1:0] TMP_1_port_2, TMP_1_port_0, TMP_1_port_1, TMP_1_v;
  wire signed [`W-1:0] TMP_0_port_2, TMP_0_port_0, TMP_0_port_1, TMP_0_v;
  wire signed [`W-1:0] N0455_port_9, N0455_port_4, N0455_v;
  wire signed [`W-1:0] N0459_port_8, N0459_port_5, N0459_v;
  wire signed [`W-1:0] RRAB0_port_8, RRAB0_port_4, RRAB0_v;
  wire signed [`W-1:0] RRAB1_port_8, RRAB1_port_4, RRAB1_v;
  wire signed [`W-1:0] N0872_port_3, N0872_port_0, N0872_port_5, N0872_v;
  wire signed [`W-1:0] S00699_port_1, S00699_v;
  wire signed [`W-1:0] _OPR_1_port_15, _OPR_1_port_16, _OPR_1_v;
  wire signed [`W-1:0] _OPR_0_port_10, _OPR_0_port_11, _OPR_0_v;
  wire signed [`W-1:0] cm_rom_port_0, cm_rom_port_1, cm_rom_v;
  wire signed [`W-1:0] cm_ram0_port_0, cm_ram0_port_1, cm_ram0_v;
  wire signed [`W-1:0] N0344_port_2, N0344_port_0, N0344_v;
  wire signed [`W-1:0] d2_port_2, d2_port_6, d2_port_5, d2_v;
  wire signed [`W-1:0] d3_port_1, d3_port_6, d3_port_5, d3_v;
  wire signed [`W-1:0] N0617_port_2, N0617_port_1, N0617_v;
  wire signed [`W-1:0] N0610_port_0, N0610_port_10, N0610_v;
  wire signed [`W-1:0] ACC_ADA_port_7, ACC_ADA_port_5, ACC_ADA_v;
  wire signed [`W-1:0] __POC__CLK2_SC_A32_X12__port_8, __POC__CLK2_SC_A32_X12__port_9, __POC__CLK2_SC_A32_X12__port_2, __POC__CLK2_SC_A32_X12__port_3, __POC__CLK2_SC_A32_X12__port_0, __POC__CLK2_SC_A32_X12__port_1, __POC__CLK2_SC_A32_X12__port_6, __POC__CLK2_SC_A32_X12__port_7, __POC__CLK2_SC_A32_X12__port_4, __POC__CLK2_SC_A32_X12__port_5, __POC__CLK2_SC_A32_X12__v;
  wire signed [`W-1:0] N0342_port_0, N0342_port_1, N0342_v;
  wire signed [`W-1:0] N0420_port_3, N0420_port_4, N0420_v;
  wire signed [`W-1:0] N0424_port_12, N0424_port_13, N0424_v;
  wire signed [`W-1:0] N0427_port_6, N0427_port_5, N0427_v;
  wire signed [`W-1:0] N0426_port_12, N0426_port_13, N0426_v;
  wire signed [`W-1:0] S00582_port_1, S00582_v;
  wire signed [`W-1:0] S00583_port_1, S00583_v;
  wire signed [`W-1:0] N0738_port_3, N0738_port_0, N0738_v;
  wire signed [`W-1:0] CY_port_2, CY_port_3, CY_port_1, CY_port_6, CY_port_5, CY_v;
  wire signed [`W-1:0] S00685_port_0, S00685_v;
  wire signed [`W-1:0] S00687_port_0, S00687_v;
  wire signed [`W-1:0] S00689_port_0, S00689_v;
  wire signed [`W-1:0] N0559_port_2, N0559_port_1, N0559_v;
  wire signed [`W-1:0] N0558_port_2, N0558_port_0, N0558_port_1, N0558_v;
  wire signed [`W-1:0] N0882_port_1, N0882_port_10, N0882_port_19, N0882_v;
  wire signed [`W-1:0] N0881_port_0, N0881_port_10, N0881_port_19, N0881_v;
  wire signed [`W-1:0] S00731_port_1, S00731_v;
  wire signed [`W-1:0] S00836_port_0, S00836_v;
  wire signed [`W-1:0] S00724_port_1, S00724_v;
  wire signed [`W-1:0] N0642_port_0, N0642_port_6, N0642_v;
  wire signed [`W-1:0] S00833_port_0, S00833_v;
  wire signed [`W-1:0] N0891_port_4, N0891_port_5, N0891_v;
  wire signed [`W-1:0] N0436_port_8, N0436_port_0, N0436_v;
  wire signed [`W-1:0] N0434_port_12, N0434_port_13, N0434_v;
  wire signed [`W-1:0] N0439_port_12, N0439_port_13, N0439_v;
  wire signed [`W-1:0] reset_port_2, reset_v;
  wire signed [`W-1:0] N0943_port_3, N0943_port_4, N0943_v;
  wire signed [`W-1:0] N0893_port_4, N0893_port_5, N0893_v;
  wire signed [`W-1:0] N0548_port_2, N0548_port_0, N0548_port_1, N0548_v;
  wire signed [`W-1:0] N0549_port_2, N0549_port_0, N0549_port_1, N0549_v;
  wire signed [`W-1:0] S00839_port_1, S00839_v;
  wire signed [`W-1:0] N0543_port_8, N0543_port_9, N0543_v;
  wire signed [`W-1:0] N0544_port_8, N0544_port_9, N0544_v;
  wire signed [`W-1:0] N0545_port_8, N0545_port_7, N0545_v;
  wire signed [`W-1:0] N0466_port_2, N0466_port_11, N0466_v;
  wire signed [`W-1:0] _OPR_3_port_10, _OPR_3_port_11, _OPR_3_v;
  wire signed [`W-1:0] _OPR_2_port_12, _OPR_2_port_13, _OPR_2_v;
  wire signed [`W-1:0] N0513_port_2, N0513_port_3, N0513_port_0, N0513_port_1, N0513_v;
  wire signed [`W-1:0] M22_port_10, M22_port_11, M22_v;
  wire signed [`W-1:0] SC_A22_M22_CLK2_port_8, SC_A22_M22_CLK2_port_9, SC_A22_M22_CLK2_v;
  wire signed [`W-1:0] OPA_IB_port_6, OPA_IB_port_7, OPA_IB_v;
  wire signed [`W-1:0] S00654_port_1, S00654_v;
  wire signed [`W-1:0] S00818_port_0, S00818_v;
  wire signed [`W-1:0] S00729_port_1, S00729_v;
  wire signed [`W-1:0] N0409_port_3, N0409_port_4, N0409_v;
  wire signed [`W-1:0] N0406_port_12, N0406_port_13, N0406_v;
  wire signed [`W-1:0] S00678_port_1, S00678_v;
  wire signed [`W-1:0] N0713_port_2, N0713_port_5, N0713_v;
  wire signed [`W-1:0] N0710_port_2, N0710_port_1, N0710_v;
  wire signed [`W-1:0] N0717_port_3, N0717_port_5, N0717_v;
  wire signed [`W-1:0] N0715_port_4, N0715_port_5, N0715_v;
  wire signed [`W-1:0] N0714_port_2, N0714_port_5, N0714_v;
  wire signed [`W-1:0] N0574_port_0, N0574_port_11, N0574_v;
  wire signed [`W-1:0] N0571_port_9, N0571_port_0, N0571_v;
  wire signed [`W-1:0] N0570_port_8, N0570_port_7, N0570_v;
  wire signed [`W-1:0] S00825_port_0, S00825_v;
  wire signed [`W-1:0] S00531_port_0, S00531_v;
  wire signed [`W-1:0] S00536_port_1, S00536_v;
  wire signed [`W-1:0] N0889_port_4, N0889_port_5, N0889_v;
  wire signed [`W-1:0] N0514_port_2, N0514_port_3, N0514_port_0, N0514_port_6, N0514_port_4, N0514_port_5, N0514_v;
  wire signed [`W-1:0] N0848_port_2, N0848_port_0, N0848_port_1, N0848_port_6, N0848_port_4, N0848_port_5, N0848_v;
  wire signed [`W-1:0] M12_port_10, M12_port_11, M12_v;
  wire signed [`W-1:0] N0381_port_12, N0381_port_13, N0381_v;
  wire signed [`W-1:0] N0382_port_6, N0382_port_5, N0382_v;
  wire signed [`W-1:0] N0410_port_12, N0410_port_13, N0410_v;
  wire signed [`W-1:0] N0411_port_6, N0411_port_5, N0411_v;
  wire signed [`W-1:0] N0415_port_8, N0415_port_0, N0415_v;
  wire signed [`W-1:0] _COM_port_0, _COM_port_1, _COM_v;
  wire signed [`W-1:0] N0700_port_2, N0700_port_3, N0700_v;
  wire signed [`W-1:0] N0702_port_0, N0702_port_1, N0702_v;
  wire signed [`W-1:0] D2_port_13, D2_port_14, D2_port_15, D2_port_16, D2_port_17, D2_port_19, D2_port_9, D2_port_2, D2_port_3, D2_port_1, D2_port_6, D2_port_7, D2_port_5, D2_v;
  wire signed [`W-1:0] D3_port_13, D3_port_14, D3_port_15, D3_port_16, D3_port_17, D3_port_19, D3_port_9, D3_port_3, D3_port_0, D3_port_1, D3_port_6, D3_port_7, D3_port_5, D3_v;
  wire signed [`W-1:0] D0_port_11, D0_port_12, D0_port_13, D0_port_14, D0_port_15, D0_port_16, D0_port_19, D0_port_8, D0_port_3, D0_port_1, D0_port_6, D0_port_4, D0_port_5, D0_v;
  wire signed [`W-1:0] D1_port_12, D1_port_13, D1_port_14, D1_port_15, D1_port_16, D1_port_19, D1_port_9, D1_port_2, D1_port_3, D1_port_1, D1_port_7, D1_port_4, D1_port_5, D1_v;
  wire signed [`W-1:0] N0565_port_8, N0565_port_9, N0565_v;
  wire signed [`W-1:0] N0569_port_8, N0569_port_9, N0569_v;
  wire signed [`W-1:0] S00814_port_0, S00814_v;
  wire signed [`W-1:0] S00676_port_0, S00676_v;
  wire signed [`W-1:0] _OPA_0_port_13, _OPA_0_port_14, _OPA_0_v;
  wire signed [`W-1:0] _OPA_2_port_6, _OPA_2_port_7, _OPA_2_v;
  wire signed [`W-1:0] _OPA_3_port_10, _OPA_3_port_11, _OPA_3_v;
  wire signed [`W-1:0] N0646_port_2, N0646_port_1, N0646_v;
  wire signed [`W-1:0] ___SC__JIN_FIN__CLK1_M11_X21_INH__port_2, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_3, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_0, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_1, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_4, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_5, ___SC__JIN_FIN__CLK1_M11_X21_INH__v;
  wire signed [`W-1:0] N0941_port_3, N0941_port_4, N0941_v;
  wire signed [`W-1:0] N0861_port_2, N0861_port_3, N0861_port_0, N0861_v;
  wire signed [`W-1:0] N0866_port_0, N0866_port_10, N0866_port_19, N0866_v;
  wire signed [`W-1:0] N0911_port_2, N0911_port_0, N0911_port_1, N0911_v;
  wire signed [`W-1:0] N0621_port_0, N0621_port_1, N0621_v;
  wire signed [`W-1:0] N0771_port_1, N0771_port_6, N0771_port_11, N0771_v;
  wire signed [`W-1:0] N0770_port_2, N0770_port_6, N0770_port_11, N0770_v;
  wire signed [`W-1:0] N0773_port_1, N0773_port_6, N0773_port_11, N0773_v;
  wire signed [`W-1:0] N0772_port_1, N0772_port_6, N0772_port_11, N0772_v;
  wire signed [`W-1:0] N0775_port_0, N0775_port_6, N0775_port_11, N0775_v;
  wire signed [`W-1:0] N0774_port_0, N0774_port_6, N0774_port_11, N0774_v;
  wire signed [`W-1:0] N0777_port_1, N0777_port_6, N0777_port_11, N0777_v;
  wire signed [`W-1:0] N0776_port_0, N0776_port_6, N0776_port_11, N0776_v;
  wire signed [`W-1:0] N0779_port_0, N0779_port_6, N0779_port_11, N0779_v;
  wire signed [`W-1:0] N0778_port_0, N0778_port_6, N0778_port_11, N0778_v;
  wire signed [`W-1:0] N0626_port_1, N0626_port_5, N0626_v;
  wire signed [`W-1:0] N0914_port_2, N0914_port_0, N0914_port_1, N0914_v;
  wire signed [`W-1:0] test_port_2, test_v;
  wire signed [`W-1:0] S00834_port_0, S00834_v;
  wire signed [`W-1:0] S00804_port_0, S00804_v;
  wire signed [`W-1:0] N0599_port_8, N0599_port_7, N0599_v;
  wire signed [`W-1:0] N0598_port_8, N0598_port_9, N0598_v;
  wire signed [`W-1:0] S00801_port_1, S00801_v;
  wire signed [`W-1:0] S00800_port_0, S00800_v;
  wire signed [`W-1:0] N0591_port_8, N0591_port_9, N0591_v;
  wire signed [`W-1:0] N0606_port_0, N0606_port_1, N0606_v;
  wire signed [`W-1:0] N0600_port_9, N0600_port_0, N0600_v;
  wire signed [`W-1:0] __INH__X11_X31_CLK1_port_12, __INH__X11_X31_CLK1_port_16, __INH__X11_X31_CLK1_v;
  wire signed [`W-1:0] S00761_port_0, S00761_v;
  wire signed [`W-1:0] S00781_port_1, S00781_v;
  wire signed [`W-1:0] CY_ADAC_port_2, CY_ADAC_port_4, CY_ADAC_v;
  wire signed [`W-1:0] CLK2_SC_A12_M12__port_8, CLK2_SC_A12_M12__port_9, CLK2_SC_A12_M12__port_2, CLK2_SC_A12_M12__port_3, CLK2_SC_A12_M12__port_0, CLK2_SC_A12_M12__port_1, CLK2_SC_A12_M12__port_6, CLK2_SC_A12_M12__port_7, CLK2_SC_A12_M12__port_4, CLK2_SC_A12_M12__port_5, CLK2_SC_A12_M12__v;
  wire signed [`W-1:0] N0293_port_2, N0293_port_3, N0293_v;
  wire signed [`W-1:0] N0297_port_0, N0297_port_1, N0297_v;
  wire signed [`W-1:0] N0294_port_2, N0294_port_3, N0294_port_4, N0294_port_5, N0294_v;
  wire signed [`W-1:0] N0298_port_0, N0298_port_6, N0298_v;
  wire signed [`W-1:0] N0767_port_2, N0767_port_0, N0767_v;
  wire signed [`W-1:0] N0765_port_2, N0765_port_1, N0765_v;
  wire signed [`W-1:0] N0768_port_2, N0768_port_0, N0768_v;
  wire signed [`W-1:0] N0769_port_0, N0769_port_4, N0769_v;
  wire signed [`W-1:0] sync_port_0, sync_port_1, sync_v;
  wire signed [`W-1:0] N0584_port_8, N0584_port_7, N0584_v;
  wire signed [`W-1:0] N0582_port_2, N0582_port_1, N0582_v;
  wire signed [`W-1:0] N0583_port_8, N0583_port_9, N0583_v;
  wire signed [`W-1:0] N0581_port_8, N0581_port_9, N0581_v;
  wire signed [`W-1:0] N0619_port_8, N0619_port_9, N0619_v;
  wire signed [`W-1:0] N0616_port_8, N0616_port_9, N0616_v;
  wire signed [`W-1:0] S00612_port_1, S00612_v;
  wire signed [`W-1:0] S00613_port_0, S00613_v;
  wire signed [`W-1:0] S00580_port_1, S00580_v;
  wire signed [`W-1:0] S00581_port_1, S00581_v;
  wire signed [`W-1:0] S00584_port_1, S00584_v;
  wire signed [`W-1:0] S00585_port_1, S00585_v;
  wire signed [`W-1:0] cm_ram2_port_0, cm_ram2_port_1, cm_ram2_v;
  wire signed [`W-1:0] S00725_port_0, S00725_v;
  wire signed [`W-1:0] SC_port_13, SC_port_4, SC_v;
  wire signed [`W-1:0] N0620_port_8, N0620_port_7, N0620_v;
  wire signed [`W-1:0] N0854_port_0, N0854_port_6, N0854_v;
  wire signed [`W-1:0] _OPE_port_0, _OPE_port_1, _OPE_v;
  wire signed [`W-1:0] N0752_port_3, N0752_port_0, N0752_v;
  wire signed [`W-1:0] S00690_port_1, S00690_v;
  wire signed [`W-1:0] S00609_port_0, S00609_v;
  wire signed [`W-1:0] S00601_port_1, S00601_v;
  wire signed [`W-1:0] S00600_port_1, S00600_v;
  wire signed [`W-1:0] S00599_port_1, S00599_v;
  wire signed [`W-1:0] S00598_port_1, S00598_v;
  wire signed [`W-1:0] A32_port_8, A32_port_9, A32_v;
  wire signed [`W-1:0] S00734_port_1, S00734_v;
  wire signed [`W-1:0] S00732_port_1, S00732_v;
  wire signed [`W-1:0] __POC_CLK2_X12_X32__INH_port_2, __POC_CLK2_X12_X32__INH_port_3, __POC_CLK2_X12_X32__INH_port_0, __POC_CLK2_X12_X32__INH_port_1, __POC_CLK2_X12_X32__INH_port_4, __POC_CLK2_X12_X32__INH_port_5, __POC_CLK2_X12_X32__INH_v;
  wire signed [`W-1:0] M12_M22_CLK1__M11_M12__port_8, M12_M22_CLK1__M11_M12__port_9, M12_M22_CLK1__M11_M12__v;
  wire signed [`W-1:0] S00828_port_1, S00828_v;
  wire signed [`W-1:0] N0847_port_3, N0847_port_0, N0847_port_1, N0847_port_6, N0847_port_4, N0847_port_5, N0847_v;
  wire signed [`W-1:0] ACC_ADAC_port_3, ACC_ADAC_port_7, ACC_ADAC_v;
  wire signed [`W-1:0] _OPA_1_port_8, _OPA_1_port_7, _OPA_1_v;
  wire signed [`W-1:0] ACC_3_port_3, ACC_3_port_0, ACC_3_port_1, ACC_3_port_4, ACC_3_v;
  wire signed [`W-1:0] ACC_2_port_2, ACC_2_port_3, ACC_2_port_0, ACC_2_port_4, ACC_2_v;
  wire signed [`W-1:0] ACC_1_port_3, ACC_1_port_0, ACC_1_port_1, ACC_1_port_4, ACC_1_v;
  wire signed [`W-1:0] N0945_port_3, N0945_port_4, N0945_v;
  wire signed [`W-1:0] cm_ram1_port_0, cm_ram1_port_1, cm_ram1_v;
  wire signed [`W-1:0] cm_ram3_port_0, cm_ram3_port_1, cm_ram3_v;
  wire signed [`W-1:0] N0748_port_2, N0748_port_1, N0748_v;
  wire signed [`W-1:0] N0740_port_2, N0740_port_1, N0740_v;
  wire signed [`W-1:0] N0741_port_0, N0741_port_1, N0741_v;
  wire signed [`W-1:0] N0742_port_2, N0742_port_1, N0742_v;
  wire signed [`W-1:0] N0743_port_2, N0743_port_1, N0743_v;
  wire signed [`W-1:0] N0744_port_2, N0744_port_1, N0744_v;
  wire signed [`W-1:0] N0745_port_2, N0745_port_1, N0745_v;
  wire signed [`W-1:0] N0746_port_2, N0746_port_1, N0746_v;
  wire signed [`W-1:0] N0747_port_2, N0747_port_1, N0747_v;
  wire signed [`W-1:0] N0676_port_0, N0676_port_1, N0676_v;
  wire signed [`W-1:0] N0634_port_8, N0634_port_9, N0634_v;
  wire signed [`W-1:0] N0635_port_8, N0635_port_7, N0635_v;
  wire signed [`W-1:0] N0637_port_0, N0637_port_7, N0637_v;
  wire signed [`W-1:0] N0632_port_8, N0632_port_9, N0632_v;
  wire signed [`W-1:0] ACB_IB_port_8, ACB_IB_port_2, ACB_IB_v;
  wire signed [`W-1:0] A22_port_8, A22_port_9, A22_v;
  wire signed [`W-1:0] S00709_port_1, S00709_v;
  wire signed [`W-1:0] N0690_port_0, N0690_port_5, N0690_v;
  wire signed [`W-1:0] N0913_port_2, N0913_port_0, N0913_port_1, N0913_v;
  wire signed [`W-1:0] N0912_port_2, N0912_port_0, N0912_port_1, N0912_v;
  wire signed [`W-1:0] S00564_port_0, S00564_v;
  wire signed [`W-1:0] N0693_port_3, N0693_port_6, N0693_v;
  wire signed [`W-1:0] S00803_port_1, S00803_v;
  wire signed [`W-1:0] N0605_port_0, N0605_port_1, N0605_v;
  wire signed [`W-1:0] N0604_port_0, N0604_port_1, N0604_v;
  wire signed [`W-1:0] N0607_port_0, N0607_port_1, N0607_v;
  wire signed [`W-1:0] OPR_3_port_14, OPR_3_port_15, OPR_3_v;
  wire signed [`W-1:0] ADD_IB_port_2, ADD_IB_port_7, ADD_IB_v;
  wire signed [`W-1:0] clk1_port_28, clk1_v;
  wire signed [`W-1:0] clk2_port_51, clk2_v;
  wire signed [`W-1:0] N0645_port_8, N0645_port_9, N0645_v;
  wire signed [`W-1:0] N0647_port_8, N0647_port_9, N0647_v;
  wire signed [`W-1:0] N0648_port_8, N0648_port_7, N0648_v;
  wire signed [`W-1:0] S00840_port_1, S00840_v;
  wire signed [`W-1:0] N0869_port_0, N0869_port_10, N0869_port_19, N0869_v;
  wire signed [`W-1:0] N0868_port_0, N0868_port_10, N0868_port_19, N0868_v;
  wire signed [`W-1:0] N0867_port_0, N0867_port_10, N0867_port_19, N0867_v;
  wire signed [`W-1:0] A12_port_9, A12_port_10, A12_v;
  wire signed [`W-1:0] S00716_port_1, S00716_v;
  wire signed [`W-1:0] S00710_port_0, S00710_v;
  wire signed [`W-1:0] S00620_port_1, S00620_v;
  wire signed [`W-1:0] S00627_port_1, S00627_v;
  wire signed [`W-1:0] S00624_port_1, S00624_v;
  wire signed [`W-1:0] S00628_port_0, S00628_v;
  wire signed [`W-1:0] _I_O_port_0, _I_O_port_1, _I_O_v;
  wire signed [`W-1:0] d0_port_2, d0_port_6, d0_port_5, d0_v;
  wire signed [`W-1:0] d1_port_2, d1_port_7, d1_port_5, d1_v;
  wire signed [`W-1:0] N0937_port_6, N0937_port_7, N0937_v;
  wire signed [`W-1:0] OPR_1_port_9, OPR_1_port_10, OPR_1_v;
  wire signed [`W-1:0] OPR_0_port_3, OPR_0_port_6, OPR_0_v;
  wire signed [`W-1:0] OPR_2_port_14, OPR_2_port_8, OPR_2_v;
  wire signed [`W-1:0] N0780_port_0, N0780_port_6, N0780_port_11, N0780_v;
  wire signed [`W-1:0] N0781_port_0, N0781_port_6, N0781_port_11, N0781_v;
  wire signed [`W-1:0] N0782_port_8, N0782_port_5, N0782_v;
  wire signed [`W-1:0] N0301_port_2, N0301_port_7, N0301_v;
  wire signed [`W-1:0] N0305_port_2, N0305_port_1, N0305_port_4, N0305_v;
  wire signed [`W-1:0] N0306_port_0, N0306_port_1, N0306_v;
  wire signed [`W-1:0] X12_port_12, X12_port_13, X12_v;
  wire signed [`W-1:0] N0657_port_8, N0657_port_9, N0657_v;
  wire signed [`W-1:0] S00762_port_1, S00762_v;
  wire signed [`W-1:0] N0716_port_7, N0716_port_4, N0716_v;
  wire signed [`W-1:0] OPA_2_port_0, OPA_2_port_4, OPA_2_port_13, OPA_2_v;
  wire signed [`W-1:0] OPA_3_port_2, OPA_3_port_0, OPA_3_port_13, OPA_3_v;
  wire signed [`W-1:0] OPA_0_port_11, OPA_0_port_12, OPA_0_port_13, OPA_0_v;
  wire signed [`W-1:0] N0873_port_0, N0873_port_4, N0873_port_5, N0873_v;
  wire signed [`W-1:0] N0870_port_2, N0870_port_0, N0870_port_6, N0870_v;
  wire signed [`W-1:0] N0871_port_0, N0871_port_6, N0871_port_5, N0871_v;
  wire signed [`W-1:0] OPA_1_port_10, OPA_1_port_11, OPA_1_port_12, OPA_1_v;
  wire signed [`W-1:0] S00778_port_0, S00778_v;
  wire signed [`W-1:0] N0696_port_3, N0696_port_6, N0696_v;
  wire signed [`W-1:0] N0469_port_1, N0469_port_7, N0469_v;
  wire signed [`W-1:0] N0464_port_3, N0464_port_6, N0464_v;
  wire signed [`W-1:0] N0461_port_2, N0461_port_6, N0461_v;
  wire signed [`W-1:0] N0463_port_2, N0463_port_11, N0463_v;
  wire signed [`W-1:0] N0687_port_0, N0687_port_5, N0687_v;
  wire signed [`W-1:0] S00557_port_1, S00557_v;
  wire signed [`W-1:0] N0689_port_0, N0689_port_4, N0689_v;
  wire signed [`W-1:0] X22_port_6, X22_port_7, X22_v;
  wire signed [`W-1:0] N0846_port_2, N0846_port_0, N0846_port_1, N0846_port_6, N0846_port_4, N0846_port_5, N0846_v;
  wire signed [`W-1:0] N0692_port_0, N0692_port_5, N0692_v;
  wire signed [`W-1:0] N0695_port_3, N0695_port_4, N0695_v;
  wire signed [`W-1:0] N0475_port_0, N0475_port_7, N0475_v;
  wire signed [`W-1:0] X32_port_11, X32_port_12, X32_v;
  wire signed [`W-1:0] N0698_port_3, N0698_port_5, N0698_v;
  wire signed [`W-1:0] S00740_port_0, S00740_v;
  wire signed [`W-1:0] S00766_port_0, S00766_v;
  wire signed [`W-1:0] N0551_port_2, N0551_port_0, N0551_port_1, N0551_v;
  wire signed [`W-1:0] S00767_port_0, S00767_v;
  wire signed [`W-1:0] N0550_port_2, N0550_port_3, N0550_port_0, N0550_port_1, N0550_v;
  wire signed [`W-1:0] N0327_port_6, N0327_port_4, N0327_v;
  wire signed [`W-1:0] S00764_port_1, S00764_v;
  wire signed [`W-1:0] N0553_port_2, N0553_port_1, N0553_v;
  wire signed [`W-1:0] S00765_port_0, S00765_v;
  wire signed [`W-1:0] N0552_port_2, N0552_port_0, N0552_port_1, N0552_v;
  wire signed [`W-1:0] N0529_port_8, N0529_port_9, N0529_v;
  wire signed [`W-1:0] N0555_port_2, N0555_port_0, N0555_port_1, N0555_v;
  wire signed [`W-1:0] S00835_port_0, S00835_v;
  wire signed [`W-1:0] N0554_port_2, N0554_port_0, N0554_port_1, N0554_v;
  wire signed [`W-1:0] N0557_port_2, N0557_port_0, N0557_port_1, N0557_v;

  wire N0443_v;
  wire N0442_v;
  wire N0447_v;
  wire N0446_v;
  wire N0445_v;
  wire N0993_v;
  wire N0992_v;
  wire N0995_v;
  wire N0994_v;
  wire N0997_v;
  wire N0999_v;
  wire N0998_v;
  wire N0536_v;
  wire N0535_v;
  wire N0534_v;
  wire N0538_v;
  wire N0528_v;
  wire INC_ISZ_v;
  wire LD_v;
  wire INC_ISZ_XCH_v;
  wire R8_3_v;
  wire R8_2_v;
  wire R8_1_v;
  wire R8_0_v;
  wire N0668_v;
  wire N0337_v;
  wire JIN_FIN_v;
  wire N0454_v;
  wire N0456_v;
  wire N0457_v;
  wire N0450_v;
  wire N0451_v;
  wire N0452_v;
  wire N0453_v;
  wire N0458_v;
  wire JCN_ISZ_v;
  wire R3_0_v;
  wire R3_1_v;
  wire R3_3_v;
  wire LDM_BBL_v;
  wire N0983_v;
  wire R1_2_v;
  wire R1_3_v;
  wire N0366_v;
  wire R7_0_v;
  wire R7_1_v;
  wire R7_2_v;
  wire R7_3_v;
  wire N0902_v;
  wire R5_2_v;
  wire R5_0_v;
  wire N0524_v;
  wire N0522_v;
  wire BBL_v;
  wire N0964_v;
  wire POC_v;
  wire N0357_v;
  wire N0996_v;
  wire WRAB1_v;
  wire WRAB0_v;
  wire DCL_v;
  wire N0348_v;
  wire N0349_v;
  wire KBP_v;
  wire N0615_v;
  wire PC0_9_v;
  wire PC0_8_v;
  wire RADB2_v;
  wire RADB0_v;
  wire RADB1_v;
  wire PC0_1_v;
  wire PC0_0_v;
  wire PC0_3_v;
  wire PC0_2_v;
  wire PC0_5_v;
  wire PC0_4_v;
  wire PC0_7_v;
  wire PC0_6_v;
  wire N0421_v;
  wire N0423_v;
  wire N0422_v;
  wire N0425_v;
  wire N0428_v;
  wire N0343_v;
  wire O_IB_v;
  wire WRITE_CARRY_2__v;
  wire N0739_v;
  wire N0735_v;
  wire N0734_v;
  wire N0737_v;
  wire N0736_v;
  wire N0731_v;
  wire N0730_v;
  wire N0733_v;
  wire N0732_v;
  wire N0397_v;
  wire N0533_v;
  wire N0383_v;
  wire N0532_v;
  wire N0531_v;
  wire N0537_v;
  wire N0641_v;
  wire IOW_v;
  wire IOR_v;
  wire N0356_v;
  wire N0643_v;
  wire PC2_11_v;
  wire PC2_10_v;
  wire JMS_v;
  wire CY_IB_v;
  wire N0358_v;
  wire SUB_v;
  wire N0432_v;
  wire N0433_v;
  wire N0430_v;
  wire N0431_v;
  wire N0437_v;
  wire N0435_v;
  wire N0438_v;
  wire ADD_v;
  wire ADM_v;
  wire N0728_v;
  wire N0729_v;
  wire N0726_v;
  wire N0727_v;
  wire N0724_v;
  wire N0725_v;
  wire N0722_v;
  wire N0723_v;
  wire N0720_v;
  wire N0721_v;
  wire N0946_v;
  wire N0944_v;
  wire N0942_v;
  wire N0940_v;
  wire N0542_v;
  wire N0540_v;
  wire N0541_v;
  wire N0546_v;
  wire N0547_v;
  wire N0467_v;
  wire INC_GROUP_5__v;
  wire N0502_v;
  wire N0682_v;
  wire N0517_v;
  wire XCH_v;
  wire CMC_v;
  wire CMA_v;
  wire N0510_v;
  wire JUN2_JMS2_v;
  wire N0361_v;
  wire N0345_v;
  wire N0364_v;
  wire N0362_v;
  wire N0363_v;
  wire N0360_v;
  wire N0399_v;
  wire N0396_v;
  wire N0395_v;
  wire N0394_v;
  wire N0393_v;
  wire N0392_v;
  wire N0391_v;
  wire N0390_v;
  wire N0408_v;
  wire N0407_v;
  wire N0405_v;
  wire N0404_v;
  wire N0403_v;
  wire N0402_v;
  wire N0401_v;
  wire N0400_v;
  wire SBM_v;
  wire _CN_v;
  wire N0719_v;
  wire N0718_v;
  wire N0711_v;
  wire N0974_v;
  wire SC_M12_CLK2_v;
  wire N0577_v;
  wire N0573_v;
  wire N0578_v;
  wire N0379_v;
  wire PC1_0_v;
  wire R14_1_v;
  wire R14_0_v;
  wire R14_3_v;
  wire R14_2_v;
  wire R10_1_v;
  wire R10_0_v;
  wire R10_3_v;
  wire R10_2_v;
  wire N0515_v;
  wire N0511_v;
  wire N0371_v;
  wire N0849_v;
  wire ISZ_v;
  wire N0370_v;
  wire N0875_v;
  wire R12_3_v;
  wire CLB_v;
  wire CLC_v;
  wire __X21__CLK2__v;
  wire DC_v;
  wire N0388_v;
  wire N0389_v;
  wire N0380_v;
  wire N0384_v;
  wire N0385_v;
  wire N0386_v;
  wire N0387_v;
  wire R12_0_v;
  wire N0419_v;
  wire N0413_v;
  wire N0414_v;
  wire N0416_v;
  wire N0704_v;
  wire N0705_v;
  wire N0707_v;
  wire N0701_v;
  wire N0703_v;
  wire N0708_v;
  wire N0885_v;
  wire N0378_v;
  wire N0965_v;
  wire N0884_v;
  wire N0560_v;
  wire N0561_v;
  wire N0564_v;
  wire N0566_v;
  wire N0568_v;
  wire N0365_v;
  wire N0368_v;
  wire N0369_v;
  wire N0314_v;
  wire ADD_GROUP_4__v;
  wire N0486_v;
  wire N0863_v;
  wire N0862_v;
  wire N0865_v;
  wire N0864_v;
  wire WRITE_ACC_1__v;
  wire N0855_v;
  wire IO_v;
  wire N0280_v;
  wire N0284_v;
  wire N0286_v;
  wire N0289_v;
  wire N0288_v;
  wire N0919_v;
  wire N0918_v;
  wire N0915_v;
  wire N0590_v;
  wire N0593_v;
  wire N0592_v;
  wire N0609_v;
  wire N0359_v;
  wire N0603_v;
  wire N0917_v;
  wire N0292_v;
  wire N0290_v;
  wire N0291_v;
  wire N0296_v;
  wire N0295_v;
  wire N0762_v;
  wire N0763_v;
  wire N0760_v;
  wire N0761_v;
  wire N0766_v;
  wire N0764_v;
  wire SC_A12_CLK2_v;
  wire R3_2_v;
  wire N0588_v;
  wire N0586_v;
  wire N0580_v;
  wire N0613_v;
  wire N0833_v;
  wire R2_1_v;
  wire R2_0_v;
  wire R2_3_v;
  wire R2_2_v;
  wire R0_3_v;
  wire R0_2_v;
  wire R0_1_v;
  wire R0_0_v;
  wire R1_0_v;
  wire R1_1_v;
  wire R6_1_v;
  wire R6_0_v;
  wire R6_3_v;
  wire R6_2_v;
  wire N0851_v;
  wire R4_3_v;
  wire R4_2_v;
  wire R4_1_v;
  wire R4_0_v;
  wire N0622_v;
  wire N0627_v;
  wire N0625_v;
  wire N0803_v;
  wire ADSR_v;
  wire ADDR_PTR_1_v;
  wire ADDR_PTR_0_v;
  wire READ_ACC_3__v;
  wire L_v;
  wire N0856_v;
  wire N0857_v;
  wire N0858_v;
  wire N0758_v;
  wire N0756_v;
  wire N0754_v;
  wire N0751_v;
  wire N0750_v;
  wire N0802_v;
  wire N0801_v;
  wire N0805_v;
  wire N0804_v;
  wire ADSL_v;
  wire R9_2_v;
  wire R9_3_v;
  wire R9_0_v;
  wire R9_1_v;
  wire N0521_v;
  wire FIN_FIM_v;
  wire INC_ISZ_ADD_SUB_XCH_LD_v;
  wire IAC_v;
  wire ADD_ACC_v;
  wire N0281_v;
  wire N0283_v;
  wire N0282_v;
  wire ACC_0_v;
  wire N0285_v;
  wire N0287_v;
  wire TCS_v;
  wire SC_A22_v;
  wire TCC_v;
  wire REG_RFSH_2_v;
  wire REG_RFSH_1_v;
  wire REG_RFSH_0_v;
  wire N0749_v;
  wire N0670_v;
  wire CY_1_v;
  wire N0674_v;
  wire N0677_v;
  wire N0636_v;
  wire N0630_v;
  wire N0633_v;
  wire N0329_v;
  wire N0322_v;
  wire N0326_v;
  wire N0325_v;
  wire R5_3_v;
  wire N0473_v;
  wire N0928_v;
  wire N0697_v;
  wire R5_1_v;
  wire N0691_v;
  wire N0694_v;
  wire INH_v;
  wire N0916_v;
  wire N0820_v;
  wire PC1_1_v;
  wire PC1_2_v;
  wire PC1_3_v;
  wire PC1_4_v;
  wire PC1_5_v;
  wire PC1_6_v;
  wire PC1_7_v;
  wire PC1_8_v;
  wire PC1_9_v;
  wire PC3_6_v;
  wire PC3_7_v;
  wire PC3_4_v;
  wire PC3_5_v;
  wire PC3_2_v;
  wire PC3_3_v;
  wire PC3_0_v;
  wire PC3_1_v;
  wire PC3_8_v;
  wire PC3_9_v;
  wire N0353_v;
  wire N0352_v;
  wire N0351_v;
  wire N0350_v;
  wire N0608_v;
  wire N0355_v;
  wire N0354_v;
  wire ADC_CY_v;
  wire N0852_v;
  wire N0938_v;
  wire PC2_9_v;
  wire PC2_8_v;
  wire PC2_7_v;
  wire PC2_6_v;
  wire PC2_5_v;
  wire PC2_4_v;
  wire PC2_3_v;
  wire PC2_2_v;
  wire PC2_1_v;
  wire PC2_0_v;
  wire N0797_v;
  wire N0799_v;
  wire __X31__CLK2__v;
  wire N0317_v;
  wire N0316_v;
  wire N0315_v;
  wire N0310_v;
  wire N0649_v;
  wire N0318_v;
  wire N0487_v;
  wire N0480_v;
  wire WADB2_v;
  wire WADB1_v;
  wire WADB0_v;
  wire N0489_v;
  wire N0853_v;
  wire __INH__X32_CLK2_v;
  wire N0850_v;
  wire N0346_v;
  wire N0504_v;
  wire N0505_v;
  wire SC_M22_CLK2_v;
  wire N0503_v;
  wire N0500_v;
  wire ADD_0_v;
  wire N0347_v;
  wire N1013_v;
  wire N1012_v;
  wire N1011_v;
  wire N1010_v;
  wire N1015_v;
  wire N1014_v;
  wire R15_0_v;
  wire R15_1_v;
  wire R15_2_v;
  wire R15_3_v;
  wire R11_0_v;
  wire R11_1_v;
  wire R11_2_v;
  wire R11_3_v;
  wire R13_2_v;
  wire R13_3_v;
  wire R13_0_v;
  wire R13_1_v;
  wire N0340_v;
  wire N0859_v;
  wire N0688_v;
  wire N0784_v;
  wire N0783_v;
  wire N0300_v;
  wire N0304_v;
  wire N0307_v;
  wire N0658_v;
  wire N0659_v;
  wire N0490_v;
  wire N0492_v;
  wire N0493_v;
  wire N0494_v;
  wire N0497_v;
  wire N0498_v;
  wire N0499_v;
  wire N0878_v;
  wire N0879_v;
  wire N0653_v;
  wire N0655_v;
  wire RAL_v;
  wire RAR_v;
  wire _INH_v;
  wire STC_v;
  wire FIN_FIM_SRC_JIN_v;
  wire N0876_v;
  wire N0877_v;
  wire N0874_v;
  wire N1008_v;
  wire N1009_v;
  wire N1004_v;
  wire N1005_v;
  wire N1006_v;
  wire N1007_v;
  wire N1000_v;
  wire N1001_v;
  wire N1002_v;
  wire N1003_v;
  wire PC3_10_v;
  wire PC3_11_v;
  wire FIM_SRC_v;
  wire ADDR_RFSH_1_v;
  wire ADDR_RFSH_0_v;
  wire N0375_v;
  wire N0374_v;
  wire N0377_v;
  wire N0278_v;
  wire N0279_v;
  wire DCL_1_v;
  wire DCL_0_v;
  wire DCL_2_v;
  wire N0669_v;
  wire N0667_v;
  wire N0666_v;
  wire N0665_v;
  wire N0664_v;
  wire N0663_v;
  wire N0660_v;
  wire PC1_10_v;
  wire PC1_11_v;
  wire N0460_v;
  wire N0685_v;
  wire N0398_v;
  wire R12_2_v;
  wire R12_1_v;
  wire N0519_v;
  wire OPE_v;
  wire JCN_v;
  wire N0678_v;
  wire N0679_v;
  wire N0671_v;
  wire N0672_v;
  wire N0673_v;
  wire N0675_v;
  wire N0479_v;
  wire N0476_v;
  wire N0477_v;
  wire N0474_v;
  wire N0472_v;
  wire N0470_v;
  wire N0471_v;
  wire N0699_v;
  wire CLK2_JMS_DC_M22_BBL_M22_X12_X22___v;
  wire N0506_v;
  wire N0328_v;
  wire N0955_v;
  wire DAA_v;
  wire DAC_v;
  wire _SRC_v;
  wire __FIN_X12__v;
  wire JUN_JMS_v;
  wire PC0_11_v;
  wire PC0_10_v;

  spice_pin_input pin_2245(reset, reset_v, reset_port_2);
  spice_pin_input pin_2242(clk1, clk1_v, clk1_port_28);
  spice_pin_input pin_2246(test, test_v, test_port_2);
  spice_pin_input pin_2243(clk2, clk2_v, clk2_port_51);

  spice_pin_output pin_2253(cm_ram2, cm_ram2_v);
  spice_pin_output pin_2252(cm_ram3, cm_ram3_v);
  spice_pin_output pin_2251(cm_rom, cm_rom_v);
  spice_pin_output pin_2244(sync, sync_v);
  spice_pin_output pin_2255(cm_ram0, cm_ram0_v);
  spice_pin_output pin_2254(cm_ram1, cm_ram1_v);

  spice_pin_bidirectional pin_2247(d0_i, d0_o, d0_t, d0_v, d0_port_5);
  spice_pin_bidirectional pin_2248(d1_i, d1_o, d1_t, d1_v, d1_port_5);
  spice_pin_bidirectional pin_2249(d2_i, d2_o, d2_t, d2_v, d2_port_5);
  spice_pin_bidirectional pin_2250(d3_i, d3_o, d3_t, d3_v, d3_port_5);

  spice_transistor_nmos_vdd tM3268(v(S00839_v), N0698_v, N0698_port_3);
  spice_transistor_nmos_gnd g_2406((N0515_v|v(N0342_v)), ACC_ADAC_v, ACC_ADAC_port_7);
  spice_transistor_nmos_gnd g_2677((v(N0469_v)|(N0454_v&v(N0463_v))), N0461_v, N0461_port_6);
  spice_transistor_nmos_gnd tM3157(N0735_v, cm_ram2_v, cm_ram2_port_1);
  wire [`W-1:0] temp_3276;
  spice_transistor_nmos tM1203(WADB0_v, N0780_v, a(N0763_v), N0780_port_0, temp_3276);
  spice_transistor_nmos_vdd tM1201(v(__INH__X11_X31_CLK1_v), N0775_v, N0775_port_6);
  wire [`W-1:0] temp_3277;
  spice_transistor_nmos tM1204(WADB0_v, N0781_v, a(N0764_v), N0781_port_0, temp_3277);
  spice_transistor_nmos tM1561(v(N0584_v), N0591_v, __POC__CLK2_SC_A32_X12__v, N0591_port_9, __POC__CLK2_SC_A32_X12__port_3);
  spice_transistor_nmos_vdd tM1769(v(S00581_v), N0584_v, N0584_port_7);
  spice_transistor_nmos_vdd tM1761(v(S00578_v), N0530_v, N0530_port_4);
  spice_transistor_nmos_vdd tM1763(v(S00579_v), N0545_v, N0545_port_7);
  spice_transistor_nmos_vdd tM1764(v(S00580_v), N0570_v, N0570_port_7);
  spice_transistor_nmos_vdd tM2493(N1002_v, _OPA_2_v, _OPA_2_port_7);
  spice_transistor_nmos_gnd tM2494(N1004_v, OPA_1_v, OPA_1_port_10);
  spice_transistor_nmos_vdd tM1032(N0325_v, N0298_v, N0298_port_0);
  spice_transistor_nmos_vdd tM3252(v(N0696_v), d0_v, d0_port_2);
  spice_transistor_nmos_vdd tM2700(v(S00689_v), N0689_v, N0689_port_0);
  spice_transistor_nmos_gnd tM1615(N0783_v, N0381_v, N0381_port_12);
  spice_transistor_nmos_gnd tM1614(N0783_v, N0406_v, N0406_port_12);
  spice_transistor_nmos_gnd tM1617(N0804_v, N0424_v, N0424_port_12);
  spice_transistor_nmos_gnd tM1616(N0804_v, N0410_v, N0410_port_12);
  spice_transistor_nmos tM1619(v(N0382_v), N0381_v, ___SC__JIN_FIN__CLK1_M11_X21_INH__v, N0381_port_13, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_0);
  spice_transistor_nmos tM1618(v(N0382_v), N0406_v, __POC_CLK2_X12_X32__INH_v, N0406_port_13, __POC_CLK2_X12_X32__INH_port_0);
  spice_transistor_nmos_gnd tM2830(N0727_v, A32_v, A32_port_9);
  spice_transistor_nmos_gnd tM2832(N0727_v, N0746_v, N0746_port_1);
  spice_transistor_nmos_vdd tM2834(v(S00778_v), N0746_v, N0746_port_2);
  spice_transistor_nmos_gnd tM1079(N0295_v, N0738_v, N0738_port_3);
  spice_transistor_nmos_gnd g_2317((v(N0696_v)|v(N0700_v)), N0698_v, N0698_port_5);
  spice_transistor_nmos_gnd tM2773(N0678_v, N0676_v, N0676_port_1);
  spice_transistor_nmos tM1588(v(N0635_v), N0645_v, __POC__CLK2_SC_A32_X12__v, N0645_port_9, __POC__CLK2_SC_A32_X12__port_6);
  spice_transistor_nmos_gnd g_2356((v(_COM_v)|DCL_0_v|DCL_1_v|DCL_2_v), N0716_v, N0716_port_7);
  spice_transistor_nmos_gnd g_2354((POC_v|N0630_v), N0626_v, N0626_port_5);
  spice_transistor_nmos_gnd g_2353((DC_v|v(clk2_v)|N0592_v), RRAB1_v, RRAB1_port_8);
  spice_transistor_nmos_gnd g_2408((__X21__CLK2__v|v(_OPE_v)), N0415_v, N0415_port_8);
  spice_transistor_nmos_vdd tM1868(v(S00654_v), N0344_v, N0344_port_0);
  spice_transistor_nmos_vdd tM1869(v(N0344_v), SC_v, SC_port_4);
  spice_transistor_nmos_gnd g_2725((v(N0464_v)|(v(N0466_v)&N0492_v)), N0475_v, N0475_port_7);
  spice_transistor_nmos_gnd g_2724((v(N0642_v)|(N0633_v&v(N0610_v))), N0637_v, N0637_port_7);
  spice_transistor_nmos_gnd g_2722((v(N0475_v)|(v(N0466_v)&N0458_v)), N0464_v, N0464_port_6);
  spice_transistor_nmos_gnd g_2721(((v(N0434_v)&PC2_5_v)|(v(N0406_v)&PC0_5_v)|(PC1_5_v&v(N0424_v))|(v(N0444_v)&PC3_5_v)), N0776_v, N0776_port_11);
  spice_transistor_nmos_vdd tM2454(v(S00710_v), N0742_v, N0742_port_2);
  spice_transistor_nmos_vdd g_2287((N0659_v|N0667_v), D1_v, D1_port_19);
  wire [`W-1:0] temp_3278;
  spice_transistor_nmos tM1378(RADB2_v, a(N0396_v), D0_v, temp_3278, D0_port_6);
  wire [`W-1:0] temp_3279;
  spice_transistor_nmos tM1376(WADB1_v, a(N0764_v), N0777_v, temp_3279, N0777_port_1);
  wire [`W-1:0] temp_3280;
  spice_transistor_nmos tM1377(RADB1_v, D0_v, a(N0395_v), D0_port_5, temp_3280);
  spice_transistor_nmos_vdd tM1119(v(__INH__X11_X31_CLK1_v), N0774_v, N0774_port_6);
  spice_transistor_nmos tM2950(ADSR_v, N0848_v, ACC_1_v, N0848_port_0, ACC_1_port_4);
  wire [`W-1:0] temp_3281;
  spice_transistor_nmos tM2959(v(ACC_ADA_v), N0871_v, a(N0857_v), N0871_port_6, temp_3281);
  spice_transistor_nmos_vdd tM1575(v(S00557_v), RRAB1_v, RRAB1_port_4);
  spice_transistor_nmos_vdd tM1577(v(__INH__X11_X31_CLK1_v), N0773_v, N0773_port_6);
  spice_transistor_nmos tM1570(v(N0599_v), CLK2_SC_A12_M12__v, N0598_v, CLK2_SC_A12_M12__port_4, N0598_port_9);
  spice_transistor_nmos tM1571(v(N0620_v), N0619_v, CLK2_SC_A12_M12__v, N0619_port_9, CLK2_SC_A12_M12__port_5);
  spice_transistor_nmos_vdd tM1754(v(S00599_v), N0411_v, N0411_port_5);
  spice_transistor_nmos_vdd tM1755(v(S00600_v), N0427_v, N0427_port_5);
  spice_transistor_nmos_gnd tM1023(v(N0740_v), sync_v, sync_port_0);
  spice_transistor_nmos_gnd tM2005(N0627_v, __POC__CLK2_SC_A32_X12__v, __POC__CLK2_SC_A32_X12__port_8);
  spice_transistor_nmos_vdd tM1028(v(S00536_v), N0738_v, N0738_port_0);
  spice_transistor_nmos tM1591(v(N0648_v), N0657_v, __POC__CLK2_SC_A32_X12__v, N0657_port_9, __POC__CLK2_SC_A32_X12__port_7);
  spice_transistor_nmos tM1620(v(N0411_v), N0410_v, ___SC__JIN_FIN__CLK1_M11_X21_INH__v, N0410_port_13, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_1);
  spice_transistor_nmos tM1621(v(N0411_v), N0424_v, __POC_CLK2_X12_X32__INH_v, N0424_port_13, __POC_CLK2_X12_X32__INH_port_1);
  spice_transistor_nmos_gnd tM1624(N0820_v, N0434_v, N0434_port_12);
  spice_transistor_nmos_gnd tM1625(N0820_v, N0426_v, N0426_port_12);
  spice_transistor_nmos_gnd tM1626(N0833_v, N0439_v, N0439_port_12);
  spice_transistor_nmos_gnd tM1627(N0833_v, N0444_v, N0444_port_12);
  spice_transistor_nmos_vdd tM2829(v(N0746_v), A32_v, A32_port_8);
  spice_transistor_nmos tM3191(ADSL_v, N0514_v, N0513_v, N0514_port_6, N0513_port_2);
  spice_transistor_nmos tM3193(ADSR_v, N0513_v, ACC_3_v, N0513_port_3, ACC_3_port_4);
  spice_transistor_nmos tM3194(v(N0893_v), N0914_v, N0557_v, N0914_port_0, N0557_port_1);
  spice_transistor_nmos_vdd tM2222(N0999_v, OPR_0_v, OPR_0_port_3);
  wire [`W-1:0] temp_3282;
  spice_transistor_nmos tM2854(v(ACB_IB_v), a(N0346_v), D0_v, temp_3282, D0_port_12);
  spice_transistor_nmos_gnd tM3284(N0664_v, D3_v, D3_port_17);
  spice_transistor_nmos_vdd tM3287(v(N0693_v), d1_v, d1_port_2);
  spice_transistor_nmos tM3064(N0964_v, D2_v, N0606_v, D2_port_15, N0606_port_0);
  spice_transistor_nmos tM3062(v(N0556_v), N0554_v, N0555_v, N0554_port_2, N0555_port_2);
  spice_transistor_nmos_gnd tM3068(N0944_v, _TMP_2_v, _TMP_2_port_0);
  spice_transistor_nmos tM3069(v(N0937_v), _TMP_2_v, N0891_v, _TMP_2_port_1, N0891_port_4);
  spice_transistor_nmos_gnd tM3260(N0736_v, cm_ram0_v, cm_ram0_port_1);
  spice_transistor_nmos_gnd g_2344((v(N0695_v)|POC_v), d1_v, d1_port_7);
  spice_transistor_nmos_gnd g_2343((v(N0700_v)|v(N0693_v)), N0695_v, N0695_port_4);
  spice_transistor_nmos_gnd g_2342((v(N0327_v)|v(A12_v)), N0769_v, N0769_port_4);
  spice_transistor_nmos_gnd g_2349((v(SUB_GROUP_6__v)|v(M12_v)), N0937_v, N0937_port_7);
  spice_transistor_nmos_gnd g_2334((N0540_v|N0561_v|N0542_v|N0577_v), N0570_v, N0570_port_8);
  spice_transistor_nmos_vdd tM2799(N0704_v, N0700_v, N0700_port_2);
  wire [`W-1:0] temp_3283;
  spice_transistor_nmos tM1361(v(RRAB1_v), D3_v, a(N0538_v), D3_port_5, temp_3283);
  wire [`W-1:0] temp_3284;
  spice_transistor_nmos tM1362(v(RRAB0_v), a(N0537_v), D3_v, temp_3284, D3_port_6);
  wire [`W-1:0] temp_3285;
  spice_transistor_nmos tM1109(WRAB1_v, a(N0862_v), N0866_v, temp_3285, N0866_port_0);
  spice_transistor_nmos_vdd tM1107(v(__INH__X11_X31_CLK1_v), N0770_v, N0770_port_6);
  wire [`W-1:0] temp_3286;
  spice_transistor_nmos tM2923(v(M12_v), a(N0472_v), ACC_1_v, temp_3286, ACC_1_port_0);
  spice_transistor_nmos tM2927(v(N0553_v), N0551_v, N0552_v, N0551_port_0, N0552_port_0);
  spice_transistor_nmos tM2925(ADSL_v, N0846_v, ACC_1_v, N0846_port_6, ACC_1_port_1);
  spice_transistor_nmos_gnd tM2928(v(N0871_v), N0551_v, N0551_port_1);
  spice_transistor_nmos_gnd tM2929(v(N0889_v), N0552_v, N0552_port_1);
  spice_transistor_nmos tM1569(v(N0599_v), N0616_v, __POC__CLK2_SC_A32_X12__v, N0616_port_9, __POC__CLK2_SC_A32_X12__port_4);
  spice_transistor_nmos_gnd tM1568(N0965_v, N0632_v, N0632_port_8);
  spice_transistor_nmos_gnd g_2403((v(N0690_v)|v(N0700_v)), N0692_v, N0692_port_5);
  spice_transistor_nmos_gnd g_2400((SUB_v|SBM_v|CMC_v|v(M12_v)), SUB_GROUP_6__v, SUB_GROUP_6__port_12);
  spice_transistor_nmos tM1560(v(N0584_v), N0583_v, CLK2_SC_A12_M12__v, N0583_port_9, CLK2_SC_A12_M12__port_3);
  spice_transistor_nmos_gnd tM1567(N0965_v, N0619_v, N0619_port_8);
  spice_transistor_nmos_gnd tM1566(N0955_v, N0598_v, N0598_port_8);
  wire [`W-1:0] temp_3287;
  spice_transistor_nmos tM1031(RADB0_v, a(N0388_v), D2_v, temp_3287, D2_port_1);
  spice_transistor_nmos_vdd tM1030(v(N0738_v), sync_v, sync_port_1);
  spice_transistor_nmos_vdd tM1749(v(S00598_v), N0382_v, N0382_port_5);
  spice_transistor_nmos_gnd tM1585(N0974_v, N0634_v, N0634_port_8);
  spice_transistor_nmos_gnd tM1584(N0974_v, N0645_v, N0645_port_8);
  spice_transistor_nmos_gnd tM1587(N0983_v, N0657_v, N0657_port_8);
  spice_transistor_nmos_gnd tM1586(N0983_v, N0647_v, N0647_port_8);
  spice_transistor_nmos tM1589(v(N0635_v), N0634_v, CLK2_SC_A12_M12__v, N0634_port_9, CLK2_SC_A12_M12__port_6);
  spice_transistor_nmos_vdd tM2724(v(S00716_v), OPA_IB_v, OPA_IB_port_6);
  spice_transistor_nmos_vdd tM2721(v(N0687_v), d3_v, d3_port_1);
  wire [`W-1:0] temp_3288;
  spice_transistor_nmos tM2753(CY_IB_v, D0_v, a(CY_1_v), D0_port_11, temp_3288);
  spice_transistor_nmos_vdd tM1546(v(__INH__X11_X31_CLK1_v), N0777_v, N0777_port_6);
  wire [`W-1:0] temp_3289;
  spice_transistor_nmos tM2858(ADD_ACC_v, N0846_v, a(ACC_0_v), N0846_port_4, temp_3289);
  spice_transistor_nmos_gnd tM2581(N0725_v, M12_v, M12_port_11);
  wire [`W-1:0] temp_3290;
  wire [`W-1:0] temp_3291;
  spice_transistor_nmos tM2850(ADSL_v, a(CY_1_v), a(ACC_0_v), temp_3290, temp_3291);
  spice_transistor_nmos_vdd tM2584(v(S00757_v), N0717_v, N0717_port_3);
  wire [`W-1:0] temp_3292;
  wire [`W-1:0] temp_3293;
  spice_transistor_nmos tM2857(v(M12_v), a(ACC_0_v), a(N0471_v), temp_3292, temp_3293);
  spice_transistor_nmos_vdd tM3272(v(S00819_v), N0937_v, N0937_port_6);
  spice_transistor_nmos_gnd g_2713(((v(N0424_v)&PC1_8_v)|(v(N0444_v)&PC3_8_v)|(v(N0406_v)&PC0_8_v)|(v(N0434_v)&PC2_8_v)), N0773_v, N0773_port_11);
  spice_transistor_nmos_vdd tM2212(N0998_v, _OPR_0_v, _OPR_0_port_10);
  spice_transistor_nmos_vdd tM3292(v(S00836_v), N0693_v, N0693_port_3);
  wire [`W-1:0] temp_3294;
  spice_transistor_nmos tM3175(v(N0415_v), D1_v, a(N0359_v), D1_port_15, temp_3294);
  spice_transistor_nmos_vdd tM3072(v(M12_v), N0606_v, N0606_port_1);
  spice_transistor_nmos_vdd tM3070(v(N0943_v), _TMP_2_v, _TMP_2_port_2);
  spice_transistor_nmos_vdd tM3077(v(N0913_v), N0559_v, N0559_port_2);
  spice_transistor_nmos_gnd tM3076(N0917_v, N0559_v, N0559_port_1);
  spice_transistor_nmos_gnd tM3274(N0668_v, D1_v, D1_port_16);
  spice_transistor_nmos_vdd tM2870(v(N0939_v), _TMP_0_v, _TMP_0_port_2);
  spice_transistor_nmos_gnd tM3187(v(N0893_v), N0558_v, N0558_port_0);
  spice_transistor_nmos_gnd tM3186(v(N0873_v), N0557_v, N0557_port_0);
  spice_transistor_nmos tM3179(ADSL_v, N0848_v, ACC_3_v, N0848_port_6, ACC_3_port_1);
  spice_transistor_nmos tM3189(ADD_ACC_v, N0514_v, ACC_3_v, N0514_port_5, ACC_3_port_3);
  spice_transistor_nmos_gnd tM2403(N1002_v, OPA_2_v, OPA_2_port_4);
  spice_transistor_nmos_gnd tM3181(v(N0606_v), N0943_v, N0943_port_4);
  spice_transistor_nmos_gnd g_2395((v(_COM_v)|N0749_v), N0714_v, N0714_port_5);
  spice_transistor_nmos tM2884(v(SUB_GROUP_6__v), TMP_0_v, N0887_v, TMP_0_port_0, N0887_port_5);
  wire [`W-1:0] temp_3295;
  spice_transistor_nmos tM2881(v(ACC_ADA_v), N0870_v, a(N0471_v), N0870_port_6, temp_3295);
  spice_transistor_nmos_vdd tM1359(v(__INH__X11_X31_CLK1_v), N0776_v, N0776_port_6);
  spice_transistor_nmos tM2869(v(N0937_v), _TMP_0_v, N0887_v, _TMP_0_port_1, N0887_port_3);
  spice_transistor_nmos_gnd g_2568(((__X21__CLK2__v|N0446_v)&(N0445_v|__X31__CLK2__v)), ACB_IB_v, ACB_IB_port_8);
  wire [`W-1:0] temp_3296;
  spice_transistor_nmos tM1804(v(X32_v), a(ADDR_PTR_0_v), N0420_v, temp_3296, N0420_port_4);
  spice_transistor_nmos tM3228(N0964_v, D3_v, N0607_v, D3_port_16, N0607_port_1);
  spice_transistor_nmos tM2939(v(N0889_v), N0912_v, N0551_v, N0912_port_0, N0551_port_2);
  wire [`W-1:0] temp_3297;
  spice_transistor_nmos tM2938(N0351_v, a(N0371_v), N0767_v, temp_3297, N0767_port_2);
  spice_transistor_nmos_gnd g_2413((INH_v|N0451_v|POC_v|N0447_v), N0449_v, N0449_port_7);
  spice_transistor_nmos_vdd tM1131(v(__INH__X11_X31_CLK1_v), N0778_v, N0778_port_6);
  wire [`W-1:0] temp_3298;
  spice_transistor_nmos tM1138(WADB2_v, N0771_v, a(N0762_v), N0771_port_1, temp_3298);
  spice_transistor_nmos_gnd tM2449(N0719_v, X22_v, X22_port_7);
  spice_transistor_nmos_vdd tM2448(v(N0742_v), X22_v, X22_port_6);
  spice_transistor_nmos_gnd tM2561(N0340_v, N0342_v, N0342_port_1);
  spice_transistor_nmos_gnd tM2596(N1005_v, _OPA_1_v, _OPA_1_port_7);
  spice_transistor_nmos_vdd tM2599(N1005_v, OPA_1_v, OPA_1_port_11);
  spice_transistor_nmos_vdd tM2023(v(S00627_v), N0626_v, N0626_port_1);
  spice_transistor_nmos_vdd tM3089(v(S00803_v), ACC_ADA_v, ACC_ADA_port_5);
  spice_transistor_nmos_vdd tM3084(v(N0690_v), d2_v, d2_port_2);
  spice_transistor_nmos tM3083(v(SUB_GROUP_6__v), TMP_2_v, N0891_v, TMP_2_port_2, N0891_port_5);
  spice_transistor_nmos_vdd tM3081(N0944_v, TMP_2_v, TMP_2_port_0);
  spice_transistor_nmos_gnd g_2369((v(N0342_v)|ADD_GROUP_4__v), CY_ADA_v, CY_ADA_port_4);
  spice_transistor_nmos_gnd g_2368((N0517_v|INH_v|N0522_v), __INH__X11_X31_CLK1_v, __INH__X11_X31_CLK1_port_16);
  spice_transistor_nmos tM2912(v(ADD_IB_v), N0847_v, D1_v, N0847_port_3, D1_port_12);
  spice_transistor_nmos_vdd tM2681(v(S00676_v), N0702_v, N0702_port_1);
  spice_transistor_nmos_gnd tM2680(N1006_v, OPA_0_v, OPA_0_port_12);
  spice_transistor_nmos g_2555((N0292_v&N0291_v), N0294_v, N0298_v, N0294_port_4, N0298_port_6);
  spice_transistor_nmos g_2556((N0292_v&(N0290_v&N0291_v)), N0294_v, N0301_v, N0294_port_5, N0301_port_7);
  spice_transistor_nmos_vdd tM1834(v(S00628_v), __INH__X11_X31_CLK1_v, __INH__X11_X31_CLK1_port_12);
  spice_transistor_nmos_vdd tM1836(v(N0436_v), ___SC__JIN_FIN__CLK1_M11_X21_INH__v, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_5);
  spice_transistor_nmos_vdd tM1831(v(S00612_v), N0436_v, N0436_port_0);
  spice_transistor_nmos_gnd tM1830(N0437_v, ___SC__JIN_FIN__CLK1_M11_X21_INH__v, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_4);
  spice_transistor_nmos_vdd tM1066(N0325_v, N0305_v, N0305_port_1);
  wire [`W-1:0] temp_3299;
  spice_transistor_nmos tM1018(RADB0_v, a(N0387_v), D3_v, temp_3299, D3_port_3);
  spice_transistor_nmos_vdd tM1016(N0325_v, N0301_v, N0301_port_2);
  wire [`W-1:0] temp_3300;
  spice_transistor_nmos tM1014(WADB2_v, N0770_v, a(N0761_v), N0770_port_2, temp_3300);
  wire [`W-1:0] temp_3301;
  spice_transistor_nmos tM1012(RADB1_v, D3_v, a(N0386_v), D3_port_0, temp_3301);
  wire [`W-1:0] temp_3302;
  spice_transistor_nmos tM1121(v(RRAB0_v), a(N0532_v), D0_v, temp_3302, D0_port_4);
  wire [`W-1:0] temp_3303;
  spice_transistor_nmos tM1120(v(RRAB1_v), D0_v, a(N0531_v), D0_port_3, temp_3303);
  spice_transistor_nmos tM1651(v(N0427_v), N0426_v, ___SC__JIN_FIN__CLK1_M11_X21_INH__v, N0426_port_13, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_2);
  spice_transistor_nmos tM1650(v(N0427_v), N0434_v, __POC_CLK2_X12_X32__INH_v, N0434_port_13, __POC_CLK2_X12_X32__INH_port_2);
  spice_transistor_nmos tM1653(v(N0440_v), N0444_v, __POC_CLK2_X12_X32__INH_v, N0444_port_13, __POC_CLK2_X12_X32__INH_port_3);
  spice_transistor_nmos tM1652(v(N0440_v), N0439_v, ___SC__JIN_FIN__CLK1_M11_X21_INH__v, N0439_port_13, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_3);
  spice_transistor_nmos_vdd tM2791(N0546_v, N0550_v, N0550_port_2);
  spice_transistor_nmos_gnd tM3099(N0731_v, N0748_v, N0748_port_1);
  spice_transistor_nmos_vdd tM3094(v(N0748_v), A12_v, A12_port_9);
  spice_transistor_nmos_gnd tM3097(N0731_v, A12_v, A12_port_10);
  spice_transistor_nmos_gnd tM1520(N0737_v, cm_rom_v, cm_rom_port_1);
  spice_transistor_nmos_gnd tM2966(N0879_v, N0848_v, N0848_port_1);
  spice_transistor_nmos_gnd tM3259(N0733_v, cm_ram1_v, cm_ram1_port_1);
  spice_transistor_nmos tM2301(v(OPA_IB_v), D3_v, OPA_3_v, D3_port_9, OPA_3_port_0);
  spice_transistor_nmos_vdd tM3255(v(N0716_v), cm_ram0_v, cm_ram0_port_0);
  spice_transistor_nmos_vdd tM3254(v(N0713_v), cm_ram1_v, cm_ram1_port_0);
  spice_transistor_nmos_gnd g_2318((v(N0700_v)|N0697_v), N0696_v, N0696_port_6);
  spice_transistor_nmos_gnd g_2316((N0691_v|v(N0700_v)), N0690_v, N0690_port_5);
  spice_transistor_nmos_gnd g_2314((v(N0698_v)|POC_v), d0_v, d0_port_6);
  spice_transistor_nmos tM2940(v(N0871_v), N0552_v, N0912_v, N0552_port_2, N0912_port_1);
  spice_transistor_nmos_vdd tM2468(v(S00699_v), N0782_v, N0782_port_5);
  spice_transistor_nmos_gnd tM2463(N0721_v, X12_v, X12_port_13);
  spice_transistor_nmos_gnd tM2862(v(N0887_v), N0549_v, N0549_port_1);
  spice_transistor_nmos_vdd tM1800(v(S00601_v), N0440_v, N0440_port_5);
  wire [`W-1:0] temp_3304;
  spice_transistor_nmos tM1801(v(X12_v), N0409_v, a(ADDR_RFSH_1_v), N0409_port_3, temp_3304);
  wire [`W-1:0] temp_3305;
  spice_transistor_nmos tM1802(v(X32_v), a(ADDR_PTR_1_v), N0409_v, temp_3305, N0409_port_4);
  wire [`W-1:0] temp_3306;
  spice_transistor_nmos tM1803(v(X12_v), N0420_v, a(ADDR_RFSH_0_v), N0420_port_3, temp_3306);
  spice_transistor_nmos tM2947(ADD_ACC_v, N0847_v, ACC_1_v, N0847_port_5, ACC_1_port_3);
  spice_transistor_nmos_vdd tM2462(v(N0743_v), X12_v, X12_port_12);
  spice_transistor_nmos_gnd tM2868(N0705_v, N0700_v, N0700_port_3);
  spice_transistor_nmos_vdd tM1248(v(__INH__X11_X31_CLK1_v), N0772_v, N0772_port_6);
  wire [`W-1:0] temp_3307;
  spice_transistor_nmos tM2917(v(ACC_ADAC_v), N0871_v, a(N0472_v), N0871_port_0, temp_3307);
  wire [`W-1:0] temp_3308;
  spice_transistor_nmos tM2916(v(ACB_IB_v), D1_v, a(N0347_v), D1_port_13, temp_3308);
  spice_transistor_nmos_vdd tM2914(N0875_v, N0847_v, N0847_port_4);
  wire [`W-1:0] temp_3309;
  spice_transistor_nmos tM1799(SC_A22_v, N0617_v, a(REG_RFSH_1_v), N0617_port_2, temp_3309);
  spice_transistor_nmos_vdd tM1068(N0325_v, N0752_v, N0752_port_0);
  spice_transistor_nmos tM1063(N0292_v, N0293_v, N0294_v, N0293_port_3, N0294_port_2);
  wire [`W-1:0] temp_3310;
  spice_transistor_nmos tM1794(SC_A22_v, N0582_v, a(REG_RFSH_0_v), N0582_port_2, temp_3310);
  wire [`W-1:0] temp_3311;
  spice_transistor_nmos tM1067(RADB0_v, a(N0394_v), D0_v, temp_3311, D0_port_1);
  spice_transistor_nmos_gnd g_2330((N0613_v|N0561_v|N0577_v|N0542_v), N0635_v, N0635_port_8);
  spice_transistor_nmos_gnd g_2331((N0613_v|N0561_v|N0541_v|N0560_v), N0620_v, N0620_port_8);
  spice_transistor_nmos_vdd tM1480(v(SC_A22_M22_CLK2_v), N0883_v, N0883_port_10);
  spice_transistor_nmos_vdd tM2467(v(S00725_v), N0743_v, N0743_port_2);
  spice_transistor_nmos_gnd tM2465(N0721_v, N0743_v, N0743_port_1);
  spice_transistor_nmos_vdd tM1467(v(SC_A22_M22_CLK2_v), N0882_v, N0882_port_10);
  spice_transistor_nmos_vdd tM1464(v(SC_A22_M22_CLK2_v), N0868_v, N0868_port_10);
  spice_transistor_nmos_gnd tM2861(v(N0870_v), N0548_v, N0548_port_1);
  spice_transistor_nmos_gnd tM2867(N0940_v, _TMP_0_v, _TMP_0_port_0);
  spice_transistor_nmos tM2866(v(N0887_v), N0911_v, N0548_v, N0911_port_1, N0548_port_2);
  spice_transistor_nmos tM2865(v(N0870_v), N0549_v, N0911_v, N0549_port_2, N0911_port_0);
  spice_transistor_nmos_gnd tM2315(v(clk2_v), N0297_v, N0297_port_0);
  spice_transistor_nmos_vdd tM3222(v(M12_v), N0607_v, N0607_port_0);
  spice_transistor_nmos tM3223(v(N0937_v), TMP_3_v, N0893_v, TMP_3_port_0, N0893_port_5);
  spice_transistor_nmos_vdd tM2318(v(S00678_v), N0297_v, N0297_port_1);
  spice_transistor_nmos_vdd tM3224(N0946_v, TMP_3_v, TMP_3_port_1);
  spice_transistor_nmos_vdd tM3225(v(N0914_v), N0861_v, N0861_port_3);
  spice_transistor_nmos_gnd g_2301((N0658_v|__X21__CLK2__v), OPA_IB_v, OPA_IB_port_7);
  spice_transistor_nmos_gnd g_2303((N0540_v|N0561_v|N0560_v|N0541_v), N0545_v, N0545_port_8);
  spice_transistor_nmos_vdd tM1504(v(__INH__X11_X31_CLK1_v), N0781_v, N0781_port_6);
  spice_transistor_nmos_vdd tM3134(v(N0714_v), cm_ram3_v, cm_ram3_port_0);
  spice_transistor_nmos_gnd tM1502(N0919_v, N0565_v, N0565_port_8);
  spice_transistor_nmos_gnd tM2790(v(M12_v), N0550_v, N0550_port_1);
  spice_transistor_nmos_vdd tM2816(v(S00761_v), N0745_v, N0745_port_2);
  spice_transistor_nmos_vdd tM2545(v(N0332_v), N0342_v, N0342_port_0);
  spice_transistor_nmos_vdd tM2976(v(S00766_v), N0692_v, N0692_port_0);
  spice_transistor_nmos_gnd tM1815(N0450_v, __POC_CLK2_X12_X32__INH_v, __POC_CLK2_X12_X32__INH_port_5);
  spice_transistor_nmos_vdd tM1814(v(S00613_v), N0449_v, N0449_port_1);
  spice_transistor_nmos_vdd tM1811(v(N0449_v), __POC_CLK2_X12_X32__INH_v, __POC_CLK2_X12_X32__INH_port_4);
  wire [`W-1:0] temp_3312;
  spice_transistor_nmos tM1252(v(RRAB0_v), a(N0536_v), D2_v, temp_3312, D2_port_6);
  wire [`W-1:0] temp_3313;
  spice_transistor_nmos tM1323(WRAB0_v, N0882_v, a(N0864_v), N0882_port_1, temp_3313);
  spice_transistor_nmos tM1078(N0307_v, N0305_v, N0306_v, N0305_port_2, N0306_port_0);
  spice_transistor_nmos_gnd tM1073(N0307_v, N0294_v, N0294_port_3);
  spice_transistor_nmos_gnd tM1075(N0307_v, N0752_v, N0752_port_3);
  spice_transistor_nmos_gnd tM1077(v(N0738_v), N0740_v, N0740_port_2);
  spice_transistor_nmos_gnd tM3227(v(N0945_v), TMP_3_v, TMP_3_port_2);
  spice_transistor_nmos_gnd tM1499(N0902_v, N0543_v, N0543_port_8);
  spice_transistor_nmos_vdd tM1493(v(SC_A22_M22_CLK2_v), N0869_v, N0869_port_10);
  spice_transistor_nmos_gnd tM2418(N0739_v, X32_v, X32_port_11);
  spice_transistor_nmos_vdd tM2416(v(S00690_v), N0741_v, N0741_port_1);
  spice_transistor_nmos_gnd g_2541((N0289_v&(N0292_v&(N0290_v&N0291_v))), N0305_v, N0305_port_4);
  spice_transistor_nmos_vdd tM2893(v(N0911_v), N0553_v, N0553_port_2);
  spice_transistor_nmos_gnd tM2890(v(N0604_v), N0939_v, N0939_port_3);
  spice_transistor_nmos tM1781(SC_M22_CLK2_v, D2_v, N0617_v, D2_port_7, N0617_port_1);
  spice_transistor_nmos tM1780(SC_M22_CLK2_v, D1_v, N0582_v, D1_port_7, N0582_port_1);
  spice_transistor_nmos_gnd tM2254(OPE_v, _OPE_v, _OPE_port_1);
  spice_transistor_nmos_gnd tM2250(IO_v, _I_O_v, _I_O_port_0);
  spice_transistor_nmos_vdd tM2251(N0493_v, _I_O_v, _I_O_port_1);
  spice_transistor_nmos_vdd tM3300(v(S00840_v), N0695_v, N0695_port_3);
  spice_transistor_nmos_vdd tM2892(v(S00762_v), N0939_v, N0939_port_4);
  spice_transistor_nmos_gnd g_2333((N0540_v|N0561_v|N0577_v|N0560_v), N0584_v, N0584_port_8);
  spice_transistor_nmos_gnd tM3230(v(N0607_v), N0945_v, N0945_port_3);
  spice_transistor_nmos_vdd tM3129(v(S00818_v), N0714_v, N0714_port_2);
  spice_transistor_nmos_vdd tM2631(v(S00709_v), SUB_GROUP_6__v, SUB_GROUP_6__port_1);
  spice_transistor_nmos tM2968(v(N0937_v), TMP_1_v, N0889_v, TMP_1_port_0, N0889_port_4);
  spice_transistor_nmos_gnd tM2969(N0942_v, _TMP_1_v, _TMP_1_port_0);
  spice_transistor_nmos_vdd tM2639(v(S00729_v), ADD_IB_v, ADD_IB_port_2);
  spice_transistor_nmos_vdd tM2967(v(S00767_v), N0912_v, N0912_port_2);
  spice_transistor_nmos_gnd g_2337((POC_v|v(_COM_v)), N0717_v, N0717_port_5);
  spice_transistor_nmos_vdd tM2563(v(S00731_v), N0332_v, N0332_port_5);
  spice_transistor_nmos_gnd g_2676(((v(N0565_v)&R2_2_v)|(R8_2_v&v(N0616_v))|(R12_2_v&v(N0645_v))|(v(N0581_v)&R4_2_v)|(v(N0632_v)&R10_2_v)|(R14_2_v&v(N0657_v))|(R0_2_v&v(N0543_v))|(R6_2_v&v(N0591_v))), N0882_v, N0882_port_19);
  spice_transistor_nmos_vdd tM1379(N0325_v, N0306_v, N0306_port_1);
  spice_transistor_nmos_vdd tM1318(v(SC_A22_M22_CLK2_v), N0880_v, N0880_port_10);
  spice_transistor_nmos_vdd tM1315(v(SC_A22_M22_CLK2_v), N0866_v, N0866_port_10);
  spice_transistor_nmos_gnd tM1684(N0708_v, N0710_v, N0710_port_1);
  spice_transistor_nmos_gnd tM2402(N1003_v, _OPA_2_v, _OPA_2_port_6);
  spice_transistor_nmos_vdd tM2405(N1001_v, OPA_3_v, OPA_3_port_13);
  spice_transistor_nmos_vdd tM2404(N1000_v, _OPA_3_v, _OPA_3_port_11);
  spice_transistor_nmos_vdd tM1680(v(N0710_v), M12_M22_CLK1__M11_M12__v, M12_M22_CLK1__M11_M12__port_8);
  spice_transistor_nmos_gnd tM1681(N0708_v, M12_M22_CLK1__M11_M12__v, M12_M22_CLK1__M11_M12__port_9);
  spice_transistor_nmos_vdd tM2598(N1004_v, _OPA_1_v, _OPA_1_port_8);
  spice_transistor_nmos tM2889(N0964_v, D0_v, N0604_v, D0_port_14, N0604_port_1);
  spice_transistor_nmos_gnd tM2888(N0915_v, N0553_v, N0553_port_1);
  spice_transistor_nmos_vdd tM2885(N0940_v, TMP_0_v, TMP_0_port_1);
  spice_transistor_nmos_vdd tM2887(v(M12_v), N0604_v, N0604_port_0);
  spice_transistor_nmos_gnd tM2886(v(N0939_v), TMP_0_v, TMP_0_port_2);
  spice_transistor_nmos tM2880(v(ADD_IB_v), D0_v, N0846_v, D0_port_13, N0846_port_5);
  spice_transistor_nmos_vdd tM1049(N0325_v, N0293_v, N0293_port_2);
  spice_transistor_nmos_vdd g_2315((N0659_v|N0663_v), D3_v, D3_port_19);
  spice_transistor_nmos_vdd tM2064(v(N0626_v), __POC__CLK2_SC_A32_X12__v, __POC__CLK2_SC_A32_X12__port_9);
  spice_transistor_nmos_vdd tM2249(N0510_v, _OPE_v, _OPE_port_0);
  spice_transistor_nmos_gnd tM2089(N0343_v, N0344_v, N0344_port_2);
  spice_transistor_nmos_gnd tM2088(N0343_v, SC_v, SC_port_13);
  spice_transistor_nmos_gnd g_2421((READ_ACC_3__v|v(N0342_v)), ACC_ADA_v, ACC_ADA_port_7);
  spice_transistor_nmos_gnd tM2993(v(N0605_v), N0941_v, N0941_port_3);
  spice_transistor_nmos_gnd g_2302((POC_v|v(N0689_v)), d3_v, d3_port_6);
  spice_transistor_nmos_gnd tM2183(N0992_v, OPR_3_v, OPR_3_port_15);
  spice_transistor_nmos tM3204(v(N0559_v), N0557_v, N0558_v, N0557_port_2, N0558_port_2);
  wire [`W-1:0] temp_3314;
  spice_transistor_nmos tM3200(v(ACC_ADA_v), N0873_v, a(N0859_v), N0873_port_5, temp_3314);
  spice_transistor_nmos tM3201(v(N0873_v), N0558_v, N0914_v, N0558_port_1, N0914_port_1);
  spice_transistor_nmos_gnd tM3208(N0666_v, D2_v, D2_port_17);
  spice_transistor_nmos_gnd g_2323((N0400_v|v(N0420_v)), N0427_v, N0427_port_6);
  spice_transistor_nmos_gnd g_2322((v(N0409_v)|N0401_v), N0411_v, N0411_port_6);
  spice_transistor_nmos_gnd g_2329((N0613_v|N0561_v|N0560_v|N0577_v), N0648_v, N0648_port_8);
  spice_transistor_nmos_gnd tM2333(N0739_v, N0741_v, N0741_port_0);
  spice_transistor_nmos_gnd g_2269((v(N0687_v)|v(N0700_v)), N0689_v, N0689_port_4);
  spice_transistor_nmos tM3110(v(ADD_IB_v), N0514_v, D3_v, N0514_port_2, D3_port_13);
  spice_transistor_nmos_vdd tM3112(N0877_v, N0514_v, N0514_port_3);
  wire [`W-1:0] temp_3315;
  spice_transistor_nmos tM3113(v(ACB_IB_v), D3_v, a(N0356_v), D3_port_14, temp_3315);
  wire [`W-1:0] temp_3316;
  spice_transistor_nmos tM3114(v(ACC_ADAC_v), N0873_v, a(N0474_v), N0873_port_0, temp_3316);
  spice_transistor_nmos_gnd g_2332((N0613_v|N0561_v|N0542_v|N0541_v), N0599_v, N0599_port_8);
  spice_transistor_nmos_vdd g_2630((N0403_v&v(N0415_v)), CY_v, CY_port_6);
  spice_transistor_nmos_gnd g_2688((v(N0463_v)|(N0504_v&__INH__X32_CLK2_v)), N0455_v, N0455_port_9);
  spice_transistor_nmos_gnd g_2684(((v(N0444_v)&PC3_11_v)|(PC0_11_v&v(N0406_v))|(PC2_11_v&v(N0434_v))|(PC1_11_v&v(N0424_v))), N0770_v, N0770_port_11);
  spice_transistor_nmos_gnd g_2685((v(N0637_v)|(N0653_v&v(N0610_v))), N0642_v, N0642_port_6);
  spice_transistor_nmos_gnd g_2680(((SC_A12_CLK2_v&N0586_v)|v(N0571_v)), N0574_v, N0574_port_11);
  spice_transistor_nmos_gnd g_2681((v(N0610_v)|(v(N0574_v)&N0593_v)), N0600_v, N0600_port_9);
  spice_transistor_nmos_gnd g_2682((v(N0455_v)|(N0519_v&__INH__X32_CLK2_v)), N0463_v, N0463_port_11);
  spice_transistor_nmos_gnd tM2451(N0719_v, N0742_v, N0742_port_1);
  spice_transistor_nmos_vdd tM2954(v(M12_v), N0871_v, N0871_port_5);
  spice_transistor_nmos_gnd g_2289((N0615_v|v(clk2_v)|DC_v), RRAB0_v, RRAB0_port_8);
  spice_transistor_nmos_gnd g_2665(((v(clk1_v)&(N0328_v&N0337_v))|(v(clk2_v)&((POC_v|N0329_v)&v(X22_v)))), N0332_v, N0332_port_11);
  spice_transistor_nmos_gnd g_2662(((R9_2_v&v(N0616_v))|(v(N0543_v)&R1_2_v)|(R5_2_v&v(N0581_v))|(v(N0657_v)&R15_2_v)|(R11_2_v&v(N0632_v))|(R3_2_v&v(N0565_v))|(R7_2_v&v(N0591_v))|(R13_2_v&v(N0645_v))), N0868_v, N0868_port_19);
  spice_transistor_nmos_gnd g_2660(((v(N0565_v)&R3_3_v)|(v(N0645_v)&R13_3_v)|(v(N0591_v)&R7_3_v)|(v(N0657_v)&R15_3_v)|(v(N0632_v)&R11_3_v)|(v(N0616_v)&R9_3_v)|(R5_3_v&v(N0581_v))|(v(N0543_v)&R1_3_v)), N0869_v, N0869_port_19);
  spice_transistor_nmos_gnd g_2661(((v(N0574_v)&N0625_v)|v(N0600_v)), N0610_v, N0610_port_10);
  spice_transistor_nmos_gnd g_2668(((v(N0444_v)&PC3_6_v)|(v(N0434_v)&PC2_6_v)|(v(N0406_v)&PC0_6_v)|(v(N0424_v)&PC1_6_v)), N0775_v, N0775_port_11);
  spice_transistor_nmos_gnd tM3082(v(N0943_v), TMP_2_v, TMP_2_port_1);
  spice_transistor_nmos_vdd tM3241(v(S00828_v), N0854_v, N0854_port_6);
  wire [`W-1:0] temp_3317;
  spice_transistor_nmos tM1053(WADB0_v, N0779_v, a(N0762_v), N0779_port_0, temp_3317);
  wire [`W-1:0] temp_3318;
  spice_transistor_nmos tM1052(WADB0_v, N0778_v, a(N0761_v), N0778_port_0, temp_3318);
  wire [`W-1:0] temp_3319;
  spice_transistor_nmos tM1051(WADB1_v, a(N0761_v), N0774_v, temp_3319, N0774_port_0);
  wire [`W-1:0] temp_3320;
  spice_transistor_nmos tM1057(RADB1_v, D1_v, a(N0392_v), D1_port_1, temp_3320);
  wire [`W-1:0] temp_3321;
  spice_transistor_nmos tM1056(RADB2_v, a(N0390_v), D2_v, temp_3321, D2_port_3);
  wire [`W-1:0] temp_3322;
  spice_transistor_nmos tM1055(RADB1_v, D2_v, a(N0389_v), D2_port_2, temp_3322);
  wire [`W-1:0] temp_3323;
  spice_transistor_nmos tM1054(WADB1_v, a(N0762_v), N0775_v, temp_3323, N0775_port_0);
  wire [`W-1:0] temp_3324;
  spice_transistor_nmos tM1059(RADB0_v, a(N0393_v), D1_v, temp_3324, D1_port_3);
  wire [`W-1:0] temp_3325;
  spice_transistor_nmos tM1058(RADB2_v, a(N0391_v), D1_v, temp_3325, D1_port_2);
  spice_transistor_nmos_vdd tM1026(v(S00531_v), N0740_v, N0740_port_1);
  spice_transistor_nmos_gnd g_2702(((v(N0424_v)&PC1_0_v)|(v(N0434_v)&PC2_0_v)|(PC0_0_v&v(N0406_v))|(PC3_0_v&v(N0444_v))), N0781_v, N0781_port_11);
  wire [`W-1:0] temp_3326;
  spice_transistor_nmos tM3166(v(N0415_v), D2_v, a(N0366_v), D2_port_16, temp_3326);
  spice_transistor_nmos_vdd tM2438(v(N0782_v), _COM_v, _COM_port_0);
  spice_transistor_nmos_gnd tM2439(N0784_v, _COM_v, _COM_port_1);
  spice_transistor_nmos_gnd tM3212(N0946_v, _TMP_3_v, _TMP_3_port_0);
  spice_transistor_nmos_vdd tM3216(v(N0945_v), _TMP_3_v, _TMP_3_port_2);
  spice_transistor_nmos tM3214(v(SUB_GROUP_6__v), _TMP_3_v, N0893_v, _TMP_3_port_1, N0893_port_4);
  spice_transistor_nmos_gnd tM2001(N0622_v, CLK2_SC_A12_M12__v, CLK2_SC_A12_M12__port_8);
  spice_transistor_nmos_gnd tM3219(N0918_v, N0861_v, N0861_port_2);
  spice_transistor_nmos tM1590(v(N0648_v), N0647_v, CLK2_SC_A12_M12__v, N0647_port_9, CLK2_SC_A12_M12__port_7);
  spice_transistor_nmos_vdd tM3109(v(S00814_v), N0748_v, N0748_port_2);
  wire [`W-1:0] temp_3327;
  spice_transistor_nmos tM3101(N0766_v, N0768_v, a(N0749_v), N0768_port_2, temp_3327);
  spice_transistor_nmos_vdd g_2267((N0659_v|N0669_v), D0_v, D0_port_19);
  spice_transistor_nmos_gnd g_2426((v(N0700_v)|N0694_v), N0693_v, N0693_port_6);
  spice_transistor_nmos_gnd g_2698((v(N0574_v)|(SC_A12_CLK2_v&N0566_v)), N0571_v, N0571_port_9);
  spice_transistor_nmos_gnd g_2690(((v(N0406_v)&PC0_3_v)|(v(N0424_v)&PC1_3_v)|(PC3_3_v&v(N0444_v))|(v(N0434_v)&PC2_3_v)), N0778_v, N0778_port_11);
  spice_transistor_nmos_gnd g_2694(((N0443_v|N0438_v)|(JIN_FIN_v&N0435_v)), N0436_v, N0436_port_8);
  spice_transistor_nmos_gnd g_2675(((v(N0616_v)&R8_3_v)|(v(N0645_v)&R12_3_v)|(R10_3_v&v(N0632_v))|(R4_3_v&v(N0581_v))|(R0_3_v&v(N0543_v))|(v(N0591_v)&R6_3_v)|(R14_3_v&v(N0657_v))|(v(N0565_v)&R2_3_v)), N0883_v, N0883_port_19);
  spice_transistor_nmos_gnd g_2674(((R11_0_v&v(N0632_v))|(R5_0_v&v(N0581_v))|(v(N0565_v)&R3_0_v)|(R9_0_v&v(N0616_v))|(v(N0591_v)&R7_0_v)|(R15_0_v&v(N0657_v))|(R1_0_v&v(N0543_v))|(v(N0645_v)&R13_0_v)), N0866_v, N0866_port_19);
  spice_transistor_nmos_gnd tM1998(N0622_v, N0621_v, N0621_port_0);
  spice_transistor_nmos_gnd g_2671((v(N0466_v)|(N0506_v&CLK2_JMS_DC_M22_BBL_M22_X12_X22___v)), N0459_v, N0459_port_8);
  spice_transistor_nmos_gnd g_2673(((v(N0543_v)&R1_1_v)|(R15_1_v&v(N0657_v))|(R13_1_v&v(N0645_v))|(R5_1_v&v(N0581_v))|(v(N0591_v)&R7_1_v)|(R11_1_v&v(N0632_v))|(v(N0565_v)&R3_1_v)|(R9_1_v&v(N0616_v))), N0867_v, N0867_port_19);
  spice_transistor_nmos_gnd g_2672(((CLK2_JMS_DC_M22_BBL_M22_X12_X22___v&N0521_v)|v(N0459_v)), N0466_v, N0466_port_11);
  spice_transistor_nmos_vdd tM1519(v(N0717_v), cm_rom_v, cm_rom_port_0);
  wire [`W-1:0] temp_3328;
  spice_transistor_nmos tM1193(WADB2_v, N0772_v, a(N0763_v), N0772_port_1, temp_3328);
  wire [`W-1:0] temp_3329;
  spice_transistor_nmos tM1194(WADB1_v, a(N0763_v), N0776_v, temp_3329, N0776_port_0);
  spice_transistor_nmos_vdd tM2649(v(S00724_v), ACB_IB_v, ACB_IB_port_2);
  spice_transistor_nmos_vdd tM2420(v(N0741_v), X32_v, X32_port_12);
  spice_transistor_nmos_vdd tM2426(v(S00685_v), N0415_v, N0415_port_0);
  wire [`W-1:0] temp_3330;
  spice_transistor_nmos tM2795(v(CY_ADAC_v), N0550_v, a(N0855_v), N0550_port_3, temp_3330);
  spice_transistor_nmos_vdd tM3170(v(S00833_v), N0716_v, N0716_port_4);
  spice_transistor_nmos_vdd tM3171(v(S00834_v), N0713_v, N0713_port_2);
  wire [`W-1:0] temp_3331;
  spice_transistor_nmos tM3176(v(N0415_v), D0_v, a(N0357_v), D0_port_15, temp_3331);
  wire [`W-1:0] temp_3332;
  spice_transistor_nmos tM3177(v(M12_v), a(N0474_v), ACC_3_v, temp_3332, ACC_3_port_0);
  spice_transistor_nmos_vdd g_2270((N0659_v|N0665_v), D2_v, D2_port_19);
  wire [`W-1:0] temp_3333;
  spice_transistor_nmos tM3004(N0351_v, a(N0364_v), N0765_v, temp_3333, N0765_port_1);
  spice_transistor_nmos_vdd tM3000(v(N0747_v), A22_v, A22_port_8);
  spice_transistor_nmos_gnd tM3001(N0729_v, A22_v, A22_port_9);
  wire [`W-1:0] temp_3334;
  spice_transistor_nmos tM3009(v(ACC_ADAC_v), N0872_v, a(N0858_v), N0872_port_0, temp_3334);
  spice_transistor_nmos_vdd tM3197(v(M12_v), N0873_v, N0873_port_4);
  spice_transistor_nmos_gnd tM2674(v(clk2_v), N0702_v, N0702_port_0);
  spice_transistor_nmos tM1572(v(N0620_v), N0632_v, __POC__CLK2_SC_A32_X12__v, N0632_port_9, __POC__CLK2_SC_A32_X12__port_5);
  spice_transistor_nmos tM1509(v(N0545_v), N0565_v, __POC__CLK2_SC_A32_X12__v, N0565_port_9, __POC__CLK2_SC_A32_X12__port_1);
  spice_transistor_nmos tM1508(v(N0545_v), N0544_v, CLK2_SC_A12_M12__v, N0544_port_9, CLK2_SC_A12_M12__port_1);
  spice_transistor_nmos tM1507(v(N0530_v), N0529_v, CLK2_SC_A12_M12__v, N0529_port_9, CLK2_SC_A12_M12__port_0);
  spice_transistor_nmos tM1506(v(N0530_v), N0543_v, __POC__CLK2_SC_A32_X12__v, N0543_port_9, __POC__CLK2_SC_A32_X12__port_0);
  spice_transistor_nmos_gnd tM1501(N0919_v, N0544_v, N0544_port_8);
  spice_transistor_nmos_gnd tM1500(N0902_v, N0529_v, N0529_port_8);
  spice_transistor_nmos_gnd tM2658(N0853_v, N0854_v, N0854_port_0);
  wire [`W-1:0] temp_3335;
  spice_transistor_nmos tM1214(v(RRAB1_v), D2_v, a(N0535_v), D2_port_5, temp_3335);
  spice_transistor_nmos_vdd tM1217(v(__INH__X11_X31_CLK1_v), N0771_v, N0771_port_6);
  spice_transistor_nmos_vdd tM2978(v(N0941_v), _TMP_1_v, _TMP_1_port_1);
  wire [`W-1:0] temp_3336;
  spice_transistor_nmos tM1219(WRAB1_v, a(N0863_v), N0867_v, temp_3336, N0867_port_0);
  wire [`W-1:0] temp_3337;
  spice_transistor_nmos tM1218(WRAB0_v, N0881_v, a(N0863_v), N0881_port_0, temp_3337);
  wire [`W-1:0] temp_3338;
  spice_transistor_nmos tM2748(v(M12_v), CY_v, a(N0470_v), CY_port_1, temp_3338);
  wire [`W-1:0] temp_3339;
  spice_transistor_nmos tM2749(v(CY_ADA_v), N0550_v, a(N0470_v), N0550_port_0, temp_3339);
  wire [`W-1:0] temp_3340;
  spice_transistor_nmos tM2742(ADSR_v, a(CY_1_v), N0513_v, temp_3340, N0513_port_0);
  spice_transistor_nmos_vdd tM2985(v(M12_v), N0605_v, N0605_port_0);
  spice_transistor_nmos_gnd tM2988(v(N0941_v), TMP_1_v, TMP_1_port_2);
  spice_transistor_nmos_gnd tM2296(N0997_v, _OPR_1_v, _OPR_1_port_16);
  spice_transistor_nmos_gnd tM2297(N0996_v, OPR_1_v, OPR_1_port_10);
  spice_transistor_nmos_vdd tM1726(v(S00609_v), N0710_v, N0710_port_2);
  spice_transistor_nmos_gnd tM2184(N0993_v, _OPR_3_v, _OPR_3_port_11);
  spice_transistor_nmos tM2367(v(OPA_IB_v), D2_v, OPA_2_v, D2_port_9, OPA_2_port_0);
  spice_transistor_nmos_vdd tM2004(v(N0621_v), CLK2_SC_A12_M12__v, CLK2_SC_A12_M12__port_9);
  spice_transistor_nmos_gnd g_2268((N0688_v|v(N0700_v)), N0687_v, N0687_port_5);
  spice_transistor_nmos_gnd tM3017(N0729_v, N0747_v, N0747_port_1);
  spice_transistor_nmos_vdd tM3010(N0876_v, N0848_v, N0848_port_2);
  spice_transistor_nmos_vdd tM3019(v(S00800_v), N0747_v, N0747_port_2);
  spice_transistor_nmos_vdd tM3264(v(S00835_v), N0696_v, N0696_port_3);
  spice_transistor_nmos_gnd g_2264((v(N0409_v)|v(N0420_v)), N0440_v, N0440_port_6);
  spice_transistor_nmos_vdd tM2000(v(S00620_v), N0621_v, N0621_port_1);
  spice_transistor_nmos tM2759(ADSR_v, N0846_v, CY_v, N0846_port_0, CY_port_5);
  spice_transistor_nmos_gnd tM2376(N1001_v, _OPA_3_v, _OPA_3_port_10);
  spice_transistor_nmos_gnd tM2894(N0884_v, N0847_v, N0847_port_1);
  spice_transistor_nmos_vdd tM2895(v(S00764_v), ACC_ADAC_v, ACC_ADAC_port_3);
  spice_transistor_nmos_gnd g_2659(((v(N0543_v)&R0_1_v)|(v(N0616_v)&R8_1_v)|(v(N0632_v)&R10_1_v)|(R6_1_v&v(N0591_v))|(R4_1_v&v(N0581_v))|(R12_1_v&v(N0645_v))|(v(N0657_v)&R14_1_v)|(R2_1_v&v(N0565_v))), N0881_v, N0881_port_19);
  wire [`W-1:0] temp_3341;
  spice_transistor_nmos tM1220(WRAB1_v, a(N0864_v), N0868_v, temp_3341, N0868_port_0);
  wire [`W-1:0] temp_3342;
  spice_transistor_nmos tM1156(v(RRAB0_v), a(N0533_v), D1_v, temp_3342, D1_port_5);
  wire [`W-1:0] temp_3343;
  spice_transistor_nmos tM1157(WRAB0_v, N0880_v, a(N0862_v), N0880_port_0, temp_3343);
  spice_transistor_nmos_vdd tM1154(v(__INH__X11_X31_CLK1_v), N0779_v, N0779_port_6);
  wire [`W-1:0] temp_3344;
  spice_transistor_nmos tM1155(v(RRAB1_v), D1_v, a(N0534_v), D1_port_4, temp_3344);
  spice_transistor_nmos tM2756(ADC_CY_v, N0861_v, CY_v, N0861_port_0, CY_port_3);
  spice_transistor_nmos_gnd g_2347((POC_v|v(N0692_v)), d2_v, d2_port_6);
  spice_transistor_nmos_vdd tM2994(v(N0912_v), N0556_v, N0556_port_2);
  spice_transistor_nmos_vdd tM2579(v(N0745_v), M12_v, M12_port_10);
  spice_transistor_nmos_gnd tM2852(v(M12_v), N0870_v, N0870_port_2);
  spice_transistor_nmos tM2987(v(SUB_GROUP_6__v), _TMP_1_v, N0889_v, _TMP_1_port_2, N0889_port_5);
  spice_transistor_nmos_gnd tM2377(N1000_v, OPA_3_v, OPA_3_port_2);
  spice_transistor_nmos_vdd tM2175(N0993_v, OPR_3_v, OPR_3_port_14);
  spice_transistor_nmos_vdd tM2176(N0992_v, _OPR_3_v, _OPR_3_port_10);
  spice_transistor_nmos_gnd tM2173(N0994_v, OPR_2_v, OPR_2_port_14);
  spice_transistor_nmos_gnd tM2172(N0995_v, _OPR_2_v, _OPR_2_port_13);
  spice_transistor_nmos_vdd tM2287(N0996_v, _OPR_1_v, _OPR_1_port_15);
  spice_transistor_nmos_gnd tM2286(N0999_v, _OPR_0_v, _OPR_0_port_11);
  spice_transistor_nmos_gnd tM2285(N0998_v, OPR_0_v, OPR_0_port_6);
  spice_transistor_nmos_vdd tM2288(N0997_v, OPR_1_v, OPR_1_port_9);
  spice_transistor_nmos_vdd tM3152(v(S00825_v), N0715_v, N0715_port_4);
  spice_transistor_nmos_gnd tM3158(N0734_v, cm_ram3_v, cm_ram3_port_1);
  spice_transistor_nmos_vdd tM2986(N0942_v, TMP_1_v, TMP_1_port_1);
  wire [`W-1:0] temp_3345;
  spice_transistor_nmos tM3020(N0766_v, a(N0750_v), N0765_v, temp_3345, N0765_port_2);
  wire [`W-1:0] temp_3346;
  spice_transistor_nmos tM3022(N0351_v, a(N0355_v), N0768_v, temp_3346, N0768_port_0);
  spice_transistor_nmos tM3026(ADSL_v, N0847_v, ACC_2_v, N0847_port_6, ACC_2_port_0);
  spice_transistor_nmos_vdd tM3087(v(S00801_v), N0943_v, N0943_port_3);
  wire [`W-1:0] temp_3347;
  spice_transistor_nmos tM2902(N0766_v, a(N0751_v), N0767_v, temp_3347, N0767_port_0);
  wire [`W-1:0] temp_3348;
  spice_transistor_nmos tM3167(v(N0415_v), D3_v, a(N0358_v), D3_port_15, temp_3348);
  spice_transistor_nmos_gnd g_2697(((v(N0444_v)&PC3_2_v)|(PC0_2_v&v(N0406_v))|(PC1_2_v&v(N0424_v))|(PC2_2_v&v(N0434_v))), N0779_v, N0779_port_11);
  spice_transistor_nmos_gnd g_2715((N0797_v|(N0801_v&N0329_v)|(N0799_v&N0805_v)), N0782_v, N0782_port_8);
  spice_transistor_nmos_gnd g_2712(((PC1_9_v&v(N0424_v))|(v(N0444_v)&PC3_9_v)|(PC0_9_v&v(N0406_v))|(PC2_9_v&v(N0434_v))), N0772_v, N0772_port_11);
  spice_transistor_nmos_gnd g_2422((v(SUB_GROUP_6__v)|v(N0342_v)), CY_ADAC_v, CY_ADAC_port_4);
  spice_transistor_nmos_gnd g_2423((__X31__CLK2__v|N0442_v), ADD_IB_v, ADD_IB_port_7);
  spice_transistor_nmos_gnd tM3238(N0670_v, D0_v, D0_port_16);
  spice_transistor_nmos_gnd g_2425((v(_COM_v)|N0751_v), N0713_v, N0713_port_5);
  spice_transistor_nmos_vdd tM3235(v(S00817_v), N0945_v, N0945_port_4);
  spice_transistor_nmos_gnd g_2536(((N0542_v|N0540_v|N0541_v)&__FIN_X12__v), N0530_v, N0530_port_5);
  spice_transistor_nmos_vdd tM1412(v(SC_A22_M22_CLK2_v), N0881_v, N0881_port_10);
  spice_transistor_nmos_gnd g_2658(((v(N0657_v)&R14_0_v)|(v(N0565_v)&R2_0_v)|(R10_0_v&v(N0632_v))|(R6_0_v&v(N0591_v))|(v(N0645_v)&R12_0_v)|(v(N0616_v)&R8_0_v)|(v(N0543_v)&R0_0_v)|(v(N0581_v)&R4_0_v)), N0880_v, N0880_port_19);
  spice_transistor_nmos_vdd tM1415(v(SC_A22_M22_CLK2_v), N0867_v, N0867_port_10);
  spice_transistor_nmos_vdd tM2760(v(S00732_v), CY_ADAC_v, CY_ADAC_port_2);
  wire [`W-1:0] temp_3349;
  spice_transistor_nmos tM1013(RADB2_v, a(N0385_v), D3_v, temp_3349, D3_port_1);
  spice_transistor_nmos_vdd tM2699(v(S00687_v), N0687_v, N0687_port_0);
  spice_transistor_nmos tM2752(ADSL_v, N0513_v, CY_v, N0513_port_1, CY_port_2);
  spice_transistor_nmos_vdd tM2141(N0995_v, OPR_2_v, OPR_2_port_8);
  spice_transistor_nmos_vdd tM2142(N0994_v, _OPR_2_v, _OPR_2_port_12);
  spice_transistor_nmos_gnd tM2812(N0725_v, N0745_v, N0745_port_1);
  spice_transistor_nmos_vdd tM2548(v(N0744_v), M22_v, M22_port_10);
  spice_transistor_nmos_gnd tM2549(N0723_v, M22_v, M22_port_11);
  spice_transistor_nmos_gnd tM2991(N0916_v, N0556_v, N0556_port_1);
  spice_transistor_nmos tM2678(v(OPA_IB_v), D0_v, OPA_0_v, D0_port_8, OPA_0_port_11);
  spice_transistor_nmos tM2990(N0964_v, D1_v, N0605_v, D1_port_14, N0605_port_1);
  spice_transistor_nmos_vdd tM2996(v(S00781_v), N0941_v, N0941_port_4);
  spice_transistor_nmos_gnd tM2679(N1007_v, _OPA_0_v, _OPA_0_port_13);
  spice_transistor_nmos_gnd tM3039(v(M12_v), N0872_v, N0872_port_3);
  spice_transistor_nmos_gnd tM3037(v(N0872_v), N0554_v, N0554_port_0);
  wire [`W-1:0] temp_3350;
  spice_transistor_nmos tM3032(v(M12_v), ACC_2_v, a(N0473_v), ACC_2_port_3, temp_3350);
  spice_transistor_nmos tM3031(ADD_ACC_v, N0848_v, ACC_2_v, N0848_port_4, ACC_2_port_2);
  wire [`W-1:0] temp_3351;
  spice_transistor_nmos tM3030(v(ACB_IB_v), a(N0348_v), D2_v, temp_3351, D2_port_13);
  spice_transistor_nmos tM3042(v(N0872_v), N0555_v, N0913_v, N0555_port_1, N0913_port_0);
  spice_transistor_nmos_vdd tM2977(v(S00765_v), N0690_v, N0690_port_0);
  spice_transistor_nmos_gnd tM3041(v(N0891_v), N0555_v, N0555_port_0);
  wire [`W-1:0] temp_3352;
  spice_transistor_nmos tM3046(v(ACC_ADA_v), N0872_v, a(N0473_v), N0872_port_5, temp_3352);
  spice_transistor_nmos tM3045(v(ADD_IB_v), D2_v, N0848_v, D2_port_14, N0848_port_5);
  spice_transistor_nmos_gnd tM3180(N0885_v, N0514_v, N0514_port_4);
  spice_transistor_nmos_gnd g_2705(((v(N0434_v)&PC2_7_v)|(v(N0424_v)&PC1_7_v)|(PC0_7_v&v(N0406_v))|(v(N0444_v)&PC3_7_v)), N0774_v, N0774_port_11);
  spice_transistor_nmos_gnd g_2706(((PC2_10_v&v(N0434_v))|(PC1_10_v&v(N0424_v))|(v(N0406_v)&PC0_10_v)|(PC3_10_v&v(N0444_v))), N0771_v, N0771_port_11);
  spice_transistor_nmos_gnd g_2701((v(N0461_v)|(N0489_v&v(N0463_v))), N0469_v, N0469_port_7);
  spice_transistor_nmos_gnd g_2700(((v(N0424_v)&PC1_1_v)|(v(N0434_v)&PC2_1_v)|(PC0_1_v&v(N0406_v))|(v(N0444_v)&PC3_1_v)), N0780_v, N0780_port_11);
  spice_transistor_nmos_gnd g_2703(((v(N0406_v)&PC0_4_v)|(PC1_4_v&v(N0424_v))|(v(N0434_v)&PC2_4_v)|(PC3_4_v&v(N0444_v))), N0777_v, N0777_port_11);
  spice_transistor_nmos tM2673(v(OPA_IB_v), D1_v, OPA_1_v, D1_port_9, OPA_1_port_12);
  spice_transistor_nmos_vdd tM2670(N1003_v, OPA_2_v, OPA_2_port_13);
  wire [`W-1:0] temp_3353;
  spice_transistor_nmos tM1956(SC_A22_v, N0646_v, a(REG_RFSH_2_v), N0646_port_2, temp_3353);
  spice_transistor_nmos tM1952(SC_M22_CLK2_v, D3_v, N0646_v, D3_port_7, N0646_port_1);
  spice_transistor_nmos_vdd tM1395(v(__INH__X11_X31_CLK1_v), N0780_v, N0780_port_6);
  wire [`W-1:0] temp_3354;
  spice_transistor_nmos tM1396(WRAB0_v, N0883_v, a(N0865_v), N0883_port_0, temp_3354);
  wire [`W-1:0] temp_3355;
  spice_transistor_nmos tM1397(WRAB1_v, a(N0865_v), N0869_v, temp_3355, N0869_port_0);
  wire [`W-1:0] temp_3356;
  spice_transistor_nmos tM1390(WADB2_v, N0773_v, a(N0764_v), N0773_port_1, temp_3356);
  wire [`W-1:0] temp_3357;
  spice_transistor_nmos tM2872(ADSR_v, N0847_v, a(ACC_0_v), N0847_port_0, temp_3357);
  spice_transistor_nmos_vdd tM3210(v(S00804_v), N0914_v, N0914_port_2);
  spice_transistor_nmos_gnd tM1553(N0928_v, N0581_v, N0581_port_8);
  spice_transistor_nmos_gnd tM1556(N0938_v, N0591_v, N0591_port_8);
  spice_transistor_nmos_gnd tM1557(N0955_v, N0616_v, N0616_port_8);
  spice_transistor_nmos_gnd tM1554(N0928_v, N0569_v, N0569_port_8);
  spice_transistor_nmos_gnd tM1555(N0938_v, N0583_v, N0583_port_8);
  spice_transistor_nmos tM1558(v(N0570_v), N0581_v, __POC__CLK2_SC_A32_X12__v, N0581_port_9, __POC__CLK2_SC_A32_X12__port_2);
  spice_transistor_nmos tM1559(v(N0570_v), N0569_v, CLK2_SC_A12_M12__v, N0569_port_9, CLK2_SC_A12_M12__port_2);
  spice_transistor_nmos_vdd tM1779(v(S00585_v), N0648_v, N0648_port_7);
  spice_transistor_nmos_gnd g_2259((N0400_v|N0401_v), N0382_v, N0382_port_6);
  spice_transistor_nmos_vdd tM1772(v(S00584_v), N0635_v, N0635_port_7);
  spice_transistor_nmos_vdd tM1770(v(S00582_v), N0599_v, N0599_port_7);
  spice_transistor_nmos_vdd tM1771(v(S00583_v), N0620_v, N0620_port_7);
  spice_transistor_nmos_vdd tM2777(v(S00734_v), CY_ADA_v, CY_ADA_port_3);
  spice_transistor_nmos_vdd tM2771(N0677_v, N0676_v, N0676_port_0);
  spice_transistor_nmos_gnd g_2383((N0750_v|v(_COM_v)), N0715_v, N0715_port_5);
  spice_transistor_nmos_gnd g_2382((v(reset_v)|v(N0769_v)), N0327_v, N0327_port_6);
  spice_transistor_nmos_vdd tM1609(v(S00564_v), RRAB0_v, RRAB0_port_4);
  spice_transistor_nmos_vdd tM2553(v(S00740_v), N0744_v, N0744_port_2);
  spice_transistor_nmos_gnd tM2551(N0723_v, N0744_v, N0744_port_1);
  spice_transistor_nmos_gnd tM2803(N0878_v, N0846_v, N0846_port_1);
  spice_transistor_nmos tM2802(v(N0550_v), N0548_v, N0549_v, N0548_port_0, N0549_port_0);
  spice_transistor_nmos_vdd tM2809(N0874_v, N0846_v, N0846_port_2);
  wire [`W-1:0] temp_3358;
  spice_transistor_nmos tM2808(v(ACC_ADAC_v), N0870_v, a(N0856_v), N0870_port_0, temp_3358);
  spice_transistor_nmos_vdd tM1994(v(S00624_v), SC_A22_M22_CLK2_v, SC_A22_M22_CLK2_port_8);
  spice_transistor_nmos_gnd tM1995(N0655_v, SC_A22_M22_CLK2_v, SC_A22_M22_CLK2_port_9);
  spice_transistor_nmos tM3043(v(N0891_v), N0913_v, N0554_v, N0913_port_1, N0554_port_1);
  spice_transistor_nmos tM3040(ADSR_v, N0514_v, ACC_2_v, N0514_port_0, ACC_2_port_4);
  spice_transistor_nmos_vdd tM2685(N1007_v, OPA_0_v, OPA_0_port_13);
  spice_transistor_nmos_vdd tM2684(N1006_v, _OPA_0_v, _OPA_0_port_14);
  spice_transistor_nmos_vdd tM3148(v(N0715_v), cm_ram2_v, cm_ram2_port_0);

  spice_pullup pullup_493(N0461_v, N0461_port_2);
  spice_pullup pullup_705(N0475_v, N0475_port_0);
  spice_pullup pullup_814(S00612_v, S00612_port_1);
  spice_pullup pullup_815(S00628_v, S00628_port_0);
  spice_pullup pullup_1294(S00678_v, S00678_port_1);
  spice_pullup pullup_2148(S00801_v, S00801_port_1);
  spice_pullup pullup_2105(S00834_v, S00834_port_0);
  spice_pullup pullup_710(N0464_v, N0464_port_3);
  spice_pullup pullup_933(N0637_v, N0637_port_0);
  spice_pullup pullup_934(N0642_v, N0642_port_0);
  spice_pullup pullup_1827(N0911_v, N0911_port_2);
  spice_pullup pullup_776(N0600_v, N0600_port_0);
  spice_pullup pullup_774(N0574_v, N0574_port_0);
  spice_pullup pullup_773(N0571_v, N0571_port_0);
  spice_pullup pullup_772(S00585_v, S00585_port_1);
  spice_pullup pullup_771(S00584_v, S00584_port_1);
  spice_pullup pullup_2026(S00804_v, S00804_port_0);
  spice_pullup pullup_770(S00583_v, S00583_port_1);
  spice_pullup pullup_779(N0610_v, N0610_port_0);
  spice_pullup pullup_2112(S00833_v, S00833_port_0);
  spice_pullup pullup_2167(S00817_v, S00817_port_0);
  spice_pullup pullup_1638(S00676_v, S00676_port_0);
  spice_pullup pullup_1028(S00627_v, S00627_port_1);
  spice_pullup pullup_2227(S00836_v, S00836_port_0);
  spice_pullup pullup_2173(S00819_v, S00819_port_0);
  spice_pullup pullup_2236(S00840_v, S00840_port_1);
  spice_pullup pullup_1482(S00699_v, S00699_port_1);
  spice_pullup pullup_1926(S00765_v, S00765_port_0);
  spice_pullup pullup_1927(S00766_v, S00766_port_0);
  spice_pullup pullup_599(N0455_v, N0455_port_4);
  spice_pullup pullup_2206(S00839_v, S00839_port_1);
  spice_pullup pullup_2201(S00835_v, S00835_port_0);
  spice_pullup pullup_765(S00578_v, S00578_port_1);
  spice_pullup pullup_766(S00579_v, S00579_port_1);
  spice_pullup pullup_767(S00580_v, S00580_port_1);
  spice_pullup pullup_768(S00581_v, S00581_port_1);
  spice_pullup pullup_769(S00582_v, S00582_port_1);
  spice_pullup pullup_1771(S00757_v, S00757_port_1);
  spice_pullup pullup_1770(S00761_v, S00761_port_0);
  spice_pullup pullup_789(S00598_v, S00598_port_1);
  spice_pullup pullup_1737(S00732_v, S00732_port_1);
  spice_pullup pullup_1305(N0327_v, N0327_port_4);
  spice_pullup pullup_2092(S00825_v, S00825_port_0);
  spice_pullup pullup_573(S00557_v, S00557_port_1);
  spice_pullup pullup_575(N0463_v, N0463_port_2);
  spice_pullup pullup_791(S00600_v, S00600_port_1);
  spice_pullup pullup_790(S00599_v, S00599_port_1);
  spice_pullup pullup_792(S00601_v, S00601_port_1);
  spice_pullup pullup_794(S00613_v, S00613_port_0);
  spice_pullup pullup_1789(S00778_v, S00778_port_0);
  spice_pullup pullup_1686(S00716_v, S00716_port_1);
  spice_pullup pullup_1192(N0769_v, N0769_port_0);
  spice_pullup pullup_1611(S00709_v, S00709_port_1);
  spice_pullup pullup_2180(S00828_v, S00828_port_1);
  spice_pullup pullup_2058(S00803_v, S00803_port_1);
  spice_pullup pullup_678(S00609_v, S00609_port_0);
  spice_pullup pullup_27(S00536_v, S00536_port_1);
  spice_pullup pullup_24(S00531_v, S00531_port_0);
  spice_pullup pullup_2047(S00814_v, S00814_port_0);
  spice_pullup pullup_1425(S00710_v, S00710_port_0);
  spice_pullup pullup_1736(S00734_v, S00734_port_1);
  spice_pullup pullup_450(N0469_v, N0469_port_1);
  spice_pullup pullup_850(S00654_v, S00654_port_1);
  spice_pullup pullup_983(S00624_v, S00624_port_1);
  spice_pullup pullup_2074(S00818_v, S00818_port_0);
  spice_pullup pullup_1436(S00725_v, S00725_port_0);
  spice_pullup pullup_997(S00620_v, S00620_port_1);
  spice_pullup pullup_1658(S00689_v, S00689_port_0);
  spice_pullup pullup_1659(S00687_v, S00687_port_0);
  spice_pullup pullup_1967(S00800_v, S00800_port_0);
  spice_pullup pullup_1399(S00685_v, S00685_port_0);
  spice_pullup pullup_1391(S00690_v, S00690_port_1);
  spice_pullup pullup_1869(S00767_v, S00767_port_0);
  spice_pullup pullup_1867(S00764_v, S00764_port_1);
  spice_pullup pullup_1533(S00731_v, S00731_port_1);
  spice_pullup pullup_1895(S00762_v, S00762_port_1);
  spice_pullup pullup_2015(N0913_v, N0913_port_2);
  spice_pullup pullup_2014(S00781_v, S00781_port_1);
  spice_pullup pullup_1521(S00740_v, S00740_port_0);
  spice_pullup pullup_604(S00564_v, S00564_port_0);
  spice_pullup pullup_1702(S00729_v, S00729_port_1);
  spice_pullup pullup_1703(S00724_v, S00724_port_1);
  spice_pullup pullup_860(N0466_v, N0466_port_2);
  spice_pullup pullup_865(N0459_v, N0459_port_5);

  spice_latch latch_2768(eclk,ereset, v(N0569_v), N0533_v, R4_1_v);
  spice_latch latch_2769(eclk,ereset, v(N0647_v), N0532_v, R14_0_v);
  spice_latch latch_2760(eclk,ereset, v(N0702_v), N0673_v, N0694_v);
  spice_latch latch_2761(eclk,ereset, v(N0381_v), N0394_v, PC0_0_v);
  spice_latch latch_2762(eclk,ereset, v(N0410_v), N0393_v, PC1_1_v);
  spice_latch latch_2763(eclk,ereset, v(N0439_v), N0393_v, PC3_1_v);
  spice_latch latch_2764(eclk,ereset, v(N0426_v), N0393_v, PC2_1_v);
  spice_latch latch_2765(eclk,ereset, v(M12_M22_CLK1__M11_M12__v), v(D3_v), N0500_v);
  spice_latch latch_2766(eclk,ereset, v(M12_M22_CLK1__M11_M12__v), v(D0_v), N0497_v);
  spice_latch latch_2767(eclk,ereset, v(N0439_v), N0386_v, PC3_7_v);
  spice_latch latch_2830(eclk,ereset, v(N0529_v), N0533_v, R0_1_v);
  spice_latch latch_2831(eclk,ereset, v(N0583_v), N0532_v, R6_0_v);
  spice_latch latch_2832(eclk,ereset, v(clk1_v), N0503_v, N0504_v);
  spice_latch latch_2833(eclk,ereset, v(N0598_v), N0533_v, R8_1_v);
  spice_latch latch_2834(eclk,ereset, v(N0569_v), N0537_v, R4_3_v);
  spice_latch latch_2835(eclk,ereset, v(N0583_v), N0537_v, R6_3_v);
  spice_latch latch_2836(eclk,ereset, v(N0569_v), N0538_v, R5_3_v);
  spice_latch latch_2837(eclk,ereset, v(N0854_v), N0855_v, N0452_v);
  spice_latch latch_2838(eclk,ereset, v(clk2_v), v(X12_v), N0281_v);
  spice_latch latch_2839(eclk,ereset, v(clk2_v), N0511_v, N0517_v);
  spice_latch latch_2904(eclk,ereset, v(N0439_v), N0392_v, PC3_5_v);
  spice_latch latch_2905(eclk,ereset, v(N0426_v), N0392_v, PC2_5_v);
  spice_latch latch_2906(eclk,ereset, v(N0619_v), N0535_v, R11_2_v);
  spice_latch latch_2900(eclk,ereset, N0423_v, N0421_v, N0422_v);
  spice_latch latch_2896(eclk,ereset, v(clk1_v), N0720_v, N0721_v);
  spice_latch latch_2902(eclk,ereset, v(clk1_v), N0505_v, N0506_v);
  spice_latch latch_2903(eclk,ereset, v(N0583_v), N0536_v, R6_2_v);
  spice_latch latch_2908(eclk,ereset, v(N0426_v), N0386_v, PC2_7_v);
  spice_latch latch_2909(eclk,ereset, v(N0439_v), N0385_v, PC3_11_v);
  spice_latch latch_2777(eclk,ereset, v(clk1_v), N0726_v, N0727_v);
  spice_latch latch_2776(eclk,ereset, v(clk2_v), N0369_v, N0360_v);
  spice_latch latch_2775(eclk,ereset, v(N0569_v), N0536_v, R4_2_v);
  spice_latch latch_2774(eclk,ereset, v(N0583_v), N0535_v, R7_2_v);
  spice_latch latch_2773(eclk,ereset, v(N0569_v), N0535_v, R5_2_v);
  spice_latch latch_2772(eclk,ereset, v(N0647_v), N0534_v, R15_1_v);
  spice_latch latch_2770(eclk,ereset, SC_M22_CLK2_v, v(D1_v), N1014_v);
  spice_latch latch_2827(eclk,ereset, v(clk2_v), v(M12_v), N0433_v);
  spice_latch latch_2826(eclk,ereset, v(clk2_v), N0608_v, N0615_v);
  spice_latch latch_2825(eclk,ereset, v(clk1_v), N0730_v, N0731_v);
  spice_latch latch_2824(eclk,ereset, v(clk2_v), N0288_v, N0287_v);
  spice_latch latch_2823(eclk,ereset, v(clk2_v), N0413_v, N0405_v);
  spice_latch latch_2822(eclk,ereset, v(clk1_v), N0404_v, N0397_v);
  spice_latch latch_2821(eclk,ereset, v(clk1_v), N0296_v, N0739_v);
  spice_latch latch_2820(eclk,ereset, v(N0297_v), N0296_v, N0295_v);
  spice_latch latch_2829(eclk,ereset, v(clk2_v), N0402_v, N0416_v);
  spice_latch latch_2828(eclk,ereset, SC_M12_CLK2_v, v(D3_v), N1008_v);
  spice_latch latch_2919(eclk,ereset, v(N0569_v), N0531_v, R5_0_v);
  spice_latch latch_2918(eclk,ereset, v(N0544_v), N0531_v, R3_0_v);
  spice_latch latch_2910(eclk,ereset, v(N0426_v), N0385_v, PC2_11_v);
  spice_latch latch_2917(eclk,ereset, v(N0529_v), N0531_v, R1_0_v);
  spice_latch latch_2916(eclk,ereset, v(N0381_v), N0395_v, PC0_4_v);
  spice_latch latch_2915(eclk,ereset, v(N0600_v), REG_RFSH_2_v, N0633_v);
  spice_latch latch_2914(eclk,ereset, v(clk1_v), N0573_v, N0586_v);
  spice_latch latch_2907(eclk,ereset, v(N0598_v), N0536_v, R8_2_v);
  spice_latch latch_2901(eclk,ereset, v(clk1_v), ADDR_PTR_0_v, N0521_v);
  spice_latch latch_2746(eclk,ereset, SC_M22_CLK2_v, v(D3_v), N1012_v);
  spice_latch latch_2747(eclk,ereset, v(clk1_v), N0718_v, N0719_v);
  spice_latch latch_2744(eclk,ereset, v(clk2_v), v(A12_v), N0286_v);
  spice_latch latch_2749(eclk,ereset, v(N0410_v), N0394_v, PC1_0_v);
  spice_latch latch_2782(eclk,ereset, v(N0381_v), N0393_v, PC0_1_v);
  spice_latch latch_2783(eclk,ereset, v(clk2_v), N0368_v, N0362_v);
  spice_latch latch_2780(eclk,ereset, v(N0426_v), N0387_v, PC2_3_v);
  spice_latch latch_2781(eclk,ereset, v(N0439_v), N0387_v, PC3_3_v);
  spice_latch latch_2786(eclk,ereset, v(N0544_v), N0536_v, R2_2_v);
  spice_latch latch_2787(eclk,ereset, v(N0529_v), N0536_v, R0_2_v);
  spice_latch latch_2784(eclk,ereset, v(N0571_v), REG_RFSH_1_v, N0593_v);
  spice_latch latch_2785(eclk,ereset, v(clk1_v), REG_RFSH_0_v, N0566_v);
  spice_latch latch_2788(eclk,ereset, v(N0544_v), N0535_v, R3_2_v);
  spice_latch latch_2789(eclk,ereset, v(N0529_v), N0535_v, R1_2_v);
  spice_latch latch_2818(eclk,ereset, v(N0634_v), N0537_v, R12_3_v);
  spice_latch latch_2811(eclk,ereset, v(N0598_v), N0534_v, R9_1_v);
  spice_latch latch_2791(eclk,ereset, v(M12_M22_CLK1__M11_M12__v), v(D3_v), N0289_v);
  spice_latch latch_2790(eclk,ereset, v(M12_M22_CLK1__M11_M12__v), v(D2_v), N0290_v);
  spice_latch latch_2793(eclk,ereset, v(N0381_v), N0388_v, PC0_2_v);
  spice_latch latch_2792(eclk,ereset, v(N0410_v), N0388_v, PC1_2_v);
  spice_latch latch_2795(eclk,ereset, v(N0529_v), N0532_v, R0_0_v);
  spice_latch latch_2794(eclk,ereset, v(N0410_v), N0387_v, PC1_3_v);
  spice_latch latch_2797(eclk,ereset, v(clk2_v), N0383_v, N0380_v);
  spice_latch latch_2799(eclk,ereset, v(N0634_v), N0533_v, R12_1_v);
  spice_latch latch_2798(eclk,ereset, v(N0619_v), N0534_v, R11_1_v);
  spice_latch latch_2885(eclk,ereset, v(N0410_v), N0396_v, PC1_8_v);
  spice_latch latch_2884(eclk,ereset, v(clk1_v), N0316_v, N0317_v);
  spice_latch latch_2880(eclk,ereset, SC_M12_CLK2_v, v(D1_v), N1010_v);
  spice_latch latch_2883(eclk,ereset, v(N0439_v), N0396_v, PC3_8_v);
  spice_latch latch_2889(eclk,ereset, v(N0439_v), N0391_v, PC3_9_v);
  spice_latch latch_2888(eclk,ereset, v(N0426_v), N0396_v, PC2_8_v);
  spice_latch latch_2796(eclk,ereset, v(N0702_v), N0674_v, N0697_v);
  spice_latch latch_2897(eclk,ereset, v(N0410_v), N0385_v, PC1_11_v);
  spice_latch latch_2894(eclk,ereset, v(N0598_v), N0535_v, R9_2_v);
  spice_latch latch_2893(eclk,ereset, v(N0410_v), N0392_v, PC1_5_v);
  spice_latch latch_2898(eclk,ereset, v(N0381_v), N0386_v, PC0_7_v);
  spice_latch latch_2912(eclk,ereset, 1'b1, v(clk1_v), N0325_v);
  spice_latch latch_2911(eclk,ereset, v(N0410_v), N0386_v, PC1_7_v);
  spice_latch latch_2873(eclk,ereset, v(N0544_v), N0537_v, R2_3_v);
  spice_latch latch_2887(eclk,ereset, v(N0439_v), N0395_v, PC3_4_v);
  spice_latch latch_2886(eclk,ereset, v(N0426_v), N0395_v, PC2_4_v);
  spice_latch latch_2882(eclk,ereset, SC_M12_CLK2_v, v(D2_v), N1009_v);
  spice_latch latch_2779(eclk,ereset, v(N0439_v), N0388_v, PC3_2_v);
  spice_latch latch_2778(eclk,ereset, v(N0426_v), N0388_v, PC2_2_v);
  spice_latch latch_2771(eclk,ereset, v(N0571_v), N0609_v, N0625_v);
  spice_latch latch_2913(eclk,ereset, v(N0600_v), N0641_v, N0653_v);
  spice_latch latch_2871(eclk,ereset, v(N0647_v), N0536_v, R14_2_v);
  spice_latch latch_2851(eclk,ereset, v(N0455_v), ADDR_RFSH_1_v, N0489_v);
  spice_latch latch_2852(eclk,ereset, v(N0439_v), N0390_v, PC3_10_v);
  spice_latch latch_2853(eclk,ereset, v(M12_M22_CLK1__M11_M12__v), v(D2_v), N0499_v);
  spice_latch latch_2850(eclk,ereset, v(N0410_v), N0395_v, PC1_4_v);
  spice_latch latch_2856(eclk,ereset, v(N0619_v), N0536_v, R10_2_v);
  spice_latch latch_2857(eclk,ereset, v(clk2_v), N0279_v, N0278_v);
  spice_latch latch_2854(eclk,ereset, v(N0634_v), N0535_v, R13_2_v);
  spice_latch latch_2855(eclk,ereset, v(N0647_v), N0535_v, R15_2_v);
  spice_latch latch_2858(eclk,ereset, v(clk2_v), v(A22_v), N0414_v);
  spice_latch latch_2859(eclk,ereset, N0398_v, N0407_v, N0408_v);
  spice_latch latch_2891(eclk,ereset, v(N0426_v), N0391_v, PC2_9_v);
  spice_latch latch_2923(eclk,ereset, v(N0619_v), N0531_v, R11_0_v);
  spice_latch latch_2808(eclk,ereset, v(clk2_v), N0428_v, N0438_v);
  spice_latch latch_2841(eclk,ereset, v(N0583_v), N0533_v, R6_1_v);
  spice_latch latch_2840(eclk,ereset, v(N0569_v), N0534_v, R5_1_v);
  spice_latch latch_2843(eclk,ereset, v(N0619_v), N0532_v, R10_0_v);
  spice_latch latch_2842(eclk,ereset, v(N0583_v), N0534_v, R7_1_v);
  spice_latch latch_2845(eclk,ereset, v(N0583_v), N0538_v, R7_3_v);
  spice_latch latch_2847(eclk,ereset, v(clk2_v), N0314_v, N0315_v);
  spice_latch latch_2846(eclk,ereset, v(M12_M22_CLK1__M11_M12__v), v(D1_v), N0291_v);
  spice_latch latch_2849(eclk,ereset, v(N0455_v), N0453_v, N0454_v);
  spice_latch latch_2848(eclk,ereset, v(N0381_v), N0396_v, PC0_8_v);
  spice_latch latch_2874(eclk,ereset, v(N0529_v), N0537_v, R0_3_v);
  spice_latch latch_2875(eclk,ereset, v(clk2_v), v(X12_v), N0425_v);
  spice_latch latch_2876(eclk,ereset, v(clk2_v), N0365_v, N0374_v);
  spice_latch latch_2877(eclk,ereset, v(clk2_v), N0379_v, N0384_v);
  spice_latch latch_2870(eclk,ereset, v(N0529_v), N0538_v, R1_3_v);
  spice_latch latch_2872(eclk,ereset, v(N0634_v), N0536_v, R12_2_v);
  spice_latch latch_2878(eclk,ereset, v(N0459_v), ADDR_PTR_1_v, N0492_v);
  spice_latch latch_2879(eclk,ereset, v(N0459_v), N0457_v, N0458_v);
  spice_latch latch_2739(eclk,ereset, v(clk2_v), N0588_v, N0592_v);
  spice_latch latch_2738(eclk,ereset, v(N0426_v), N0390_v, PC2_10_v);
  spice_latch latch_2868(eclk,ereset, v(N0426_v), N0389_v, PC2_6_v);
  spice_latch latch_2863(eclk,ereset, v(N0410_v), N0389_v, PC1_6_v);
  spice_latch latch_2867(eclk,ereset, v(N0439_v), N0389_v, PC3_6_v);
  spice_latch latch_2866(eclk,ereset, v(N0381_v), N0390_v, PC0_10_v);
  spice_latch latch_2865(eclk,ereset, v(N0410_v), N0390_v, PC1_10_v);
  spice_latch latch_2864(eclk,ereset, v(N0381_v), N0389_v, PC0_6_v);
  spice_latch latch_2869(eclk,ereset, v(N0544_v), N0538_v, R3_3_v);
  spice_latch latch_2862(eclk,ereset, v(clk1_v), L_v, N0707_v);
  spice_latch latch_2861(eclk,ereset, v(clk1_v), N0724_v, N0725_v);
  spice_latch latch_2860(eclk,ereset, v(N0854_v), N0858_v, N0851_v);
  spice_latch latch_2745(eclk,ereset, v(clk1_v), N0728_v, N0729_v);
  spice_latch latch_2742(eclk,ereset, SC_M22_CLK2_v, v(D0_v), N1015_v);
  spice_latch latch_2743(eclk,ereset, v(clk2_v), v(A22_v), N0285_v);
  spice_latch latch_2740(eclk,ereset, v(N0439_v), N0394_v, PC3_0_v);
  spice_latch latch_2741(eclk,ereset, v(N0381_v), N0391_v, PC0_9_v);
  spice_latch latch_2748(eclk,ereset, v(N0426_v), N0394_v, PC2_0_v);
  spice_latch latch_2895(eclk,ereset, v(clk2_v), v(M22_v), N0282_v);
  spice_latch latch_2892(eclk,ereset, v(N0410_v), N0391_v, PC1_9_v);
  spice_latch latch_2890(eclk,ereset, v(N0381_v), N0392_v, PC0_5_v);
  spice_latch latch_2899(eclk,ereset, v(N0381_v), N0385_v, PC0_11_v);
  spice_latch latch_2819(eclk,ereset, v(clk2_v), N0682_v, N0703_v);
  spice_latch latch_2816(eclk,ereset, v(N0598_v), N0538_v, R9_3_v);
  spice_latch latch_2817(eclk,ereset, v(clk1_v), N0701_v, N0685_v);
  spice_latch latch_2814(eclk,ereset, v(N0619_v), N0537_v, R10_3_v);
  spice_latch latch_2815(eclk,ereset, v(N0598_v), N0537_v, R8_3_v);
  spice_latch latch_2812(eclk,ereset, v(N0619_v), N0533_v, R10_1_v);
  spice_latch latch_2813(eclk,ereset, v(N0619_v), N0538_v, R11_3_v);
  spice_latch latch_2810(eclk,ereset, v(N0569_v), N0532_v, R4_0_v);
  spice_latch latch_2922(eclk,ereset, v(M12_M22_CLK1__M11_M12__v), v(D1_v), N0498_v);
  spice_latch latch_2920(eclk,ereset, v(N0544_v), N0532_v, R2_0_v);
  spice_latch latch_2921(eclk,ereset, v(N0583_v), N0531_v, R7_0_v);
  spice_latch latch_2926(eclk,ereset, v(N0702_v), N0671_v, N0688_v);
  spice_latch latch_2927(eclk,ereset, v(clk1_v), N0361_v, N0343_v);
  spice_latch latch_2924(eclk,ereset, v(N0598_v), N0531_v, R9_0_v);
  spice_latch latch_2925(eclk,ereset, v(N0702_v), N0701_v, N0699_v);
  spice_latch latch_2928(eclk,ereset, v(N0854_v), N0856_v, N0849_v);
  spice_latch latch_2929(eclk,ereset, N0423_v, N0430_v, N0431_v);
  spice_latch latch_2755(eclk,ereset, v(N0544_v), N0533_v, R2_1_v);
  spice_latch latch_2754(eclk,ereset, v(N0544_v), N0534_v, R3_1_v);
  spice_latch latch_2757(eclk,ereset, SC_M22_CLK2_v, v(D2_v), N1013_v);
  spice_latch latch_2756(eclk,ereset, v(N0854_v), N0857_v, N0850_v);
  spice_latch latch_2751(eclk,ereset, v(N0634_v), N0531_v, R13_0_v);
  spice_latch latch_2750(eclk,ereset, v(N0634_v), N0532_v, R12_0_v);
  spice_latch latch_2753(eclk,ereset, v(N0529_v), N0534_v, R1_1_v);
  spice_latch latch_2752(eclk,ereset, v(N0647_v), N0531_v, R15_0_v);
  spice_latch latch_2759(eclk,ereset, v(N0854_v), N0859_v, N0852_v);
  spice_latch latch_2758(eclk,ereset, v(clk1_v), ADDR_RFSH_0_v, N0519_v);
  spice_latch latch_2809(eclk,ereset, v(clk2_v), v(A32_v), N0284_v);
  spice_latch latch_2805(eclk,ereset, v(N0647_v), N0538_v, R15_3_v);
  spice_latch latch_2804(eclk,ereset, v(N0634_v), N0538_v, R13_3_v);
  spice_latch latch_2807(eclk,ereset, v(N0702_v), N0672_v, N0691_v);
  spice_latch latch_2806(eclk,ereset, v(clk2_v), v(X22_v), N0280_v);
  spice_latch latch_2801(eclk,ereset, v(N0647_v), N0533_v, R14_1_v);
  spice_latch latch_2800(eclk,ereset, v(N0634_v), N0534_v, R13_1_v);
  spice_latch latch_2803(eclk,ereset, v(N0647_v), N0537_v, R14_3_v);
  spice_latch latch_2802(eclk,ereset, v(M12_M22_CLK1__M11_M12__v), v(D0_v), N0292_v);
  spice_latch latch_2931(eclk,ereset, v(clk2_v), v(M12_v), N0283_v);
  spice_latch latch_2930(eclk,ereset, v(clk1_v), N0722_v, N0723_v);
  spice_latch latch_2932(eclk,ereset, v(N0381_v), N0387_v, PC0_3_v);
  spice_latch latch_2844(eclk,ereset, v(N0598_v), N0532_v, R8_0_v);
  spice_latch latch_2881(eclk,ereset, SC_M12_CLK2_v, v(D0_v), N1011_v);

  assign N0391_v = ~(v(N0772_v));
  assign N0560_v = ~(v(N0582_v));
  assign INH_v = ~(N0524_v);
  assign N0443_v = ~(v(clk1_v));
  assign N0636_v = ~((v(_OPR_1_v)|v(OPR_3_v)|v(OPR_2_v)|v(_OPR_0_v)));
  assign CY_IB_v = ~((__X31__CLK2__v|N0446_v));
  assign N0446_v = ~(IOW_v);
  assign N0445_v = ~(XCH_v);
  assign ADDR_PTR_1_v = ~(v(N0464_v));
  assign N0400_v = ~(v(N0409_v));
  assign ADDR_RFSH_1_v = ~(v(N0461_v));
  assign N0394_v = ~(v(N0781_v));
  assign N0885_v = ~(N0877_v);
  assign N0756_v = ~((v(N0298_v)|N0290_v));
  assign N0655_v = ~((v(clk2_v)&((v(M22_v)|v(A22_v))&v(SC_v))));
  assign N0718_v = ~(N0281_v);
  assign N0393_v = ~(v(N0780_v));
  assign N0649_v = ~((v(SC_v)&(v(clk2_v)&v(A12_v))));
  assign N0322_v = ~((_CN_v|v(SC_v)));
  assign N1007_v = ~(N1006_v);
  assign N0603_v = ~((INC_ISZ_XCH_v&(v(SC_v)&v(X32_v))));
  assign N0310_v = ~(v(SC_v));
  assign LD_v = ~((v(_OPR_1_v)|v(OPR_2_v)|v(OPR_0_v)|v(_OPR_3_v)));
  assign FIN_FIM_SRC_JIN_v = ~((v(_OPR_1_v)|v(OPR_3_v)|v(OPR_2_v)));
  assign WRAB1_v = ~(N0578_v);
  assign DC_v = ~(v(SC_v));
  assign N0369_v = ~(v(X12_v));
  assign N0337_v = ~((N0360_v|v(clk2_v)));
  assign SC_M12_CLK2_v = ~(N0660_v);
  assign __X21__CLK2__v = ~(N0337_v);
  assign N0820_v = ~(v(N0427_v));
  assign N0660_v = ~((v(M12_v)&(v(SC_v)&v(clk2_v))));
  assign N0590_v = ~((v(_OPA_0_v)&(DC_v&FIN_FIM_SRC_JIN_v)));
  assign N0578_v = ~((v(clk2_v)&((N0568_v&N0580_v)|(v(M22_v)&N0564_v))));
  assign N0917_v = ~(v(N0913_v));
  assign DAA_v = ~((v(_OPA_3_v)|v(OPA_2_v)|v(_OPA_1_v)|v(_OPA_0_v)|v(_OPE_v)));
  assign XCH_v = ~((v(_OPR_3_v)|v(_OPR_1_v)|v(_OPR_0_v)|v(OPR_2_v)));
  assign BBL_v = ~((v(_OPR_2_v)|v(OPR_1_v)|v(_OPR_3_v)|v(OPR_0_v)));
  assign JMS_v = ~((v(_OPR_2_v)|v(OPR_1_v)|v(OPR_3_v)|v(_OPR_0_v)));
  assign N0761_v = ~((N0754_v|(v(N0301_v)&N0289_v)));
  assign N0288_v = ~((v(X12_v)|v(A22_v)|v(A32_v)|v(X22_v)|v(M12_v)|v(A12_v)|v(M22_v)));
  assign N0750_v = ~(DCL_1_v);
  assign N0351_v = ~((N0353_v|__X21__CLK2__v));
  assign N0366_v = ~((N0363_v|N0370_v|N0377_v|TCS_v|N0354_v));
  assign N0730_v = ~(N0287_v);
  assign N0375_v = ~((v(clk2_v)|N0380_v));
  assign N0855_v = ~(v(CY_v));
  assign IOR_v = ~((v(_I_O_v)|v(_OPA_3_v)));
  assign N0385_v = ~(v(N0770_v));
  assign N0389_v = ~(v(N0775_v));
  assign N0460_v = ~(v(clk2_v));
  assign N0328_v = ~((POC_v|N0329_v));
  assign N0390_v = ~(v(N0771_v));
  assign N0938_v = ~(v(N0584_v));
  assign N0511_v = ~((v(M22_v)|v(X22_v)));
  assign N0993_v = ~(N0992_v);
  assign N0480_v = ~(__X31__CLK2__v);
  assign N0396_v = ~(v(N0773_v));
  assign N0538_v = ~(v(N0869_v));
  assign N0361_v = ~(N0362_v);
  assign N0704_v = ~(N0705_v);
  assign N0370_v = ~((N0347_v|N0371_v|N0348_v|N0356_v|N0350_v));
  assign N0345_v = ~((N0346_v|N0347_v|N0350_v|N0349_v|N0348_v));
  assign N0659_v = ~(N0675_v);
  assign N0737_v = ~(v(N0717_v));
  assign N0304_v = ~((v(A32_v)|(JUN_JMS_v&(v(X22_v)&N0310_v))));
  assign N0401_v = ~(v(N0420_v));
  assign N0902_v = ~(v(N0530_v));
  assign N0453_v = ~(v(N0469_v));
  assign N0329_v = ~(v(_I_O_v));
  assign N0421_v = ~(N0425_v);
  assign N0853_v = ~(v(X12_v));
  assign CLB_v = ~((v(_OPE_v)|v(OPA_3_v)|v(OPA_1_v)|v(OPA_0_v)|v(OPA_2_v)));
  assign N1000_v = ~(N1012_v);
  assign N0395_v = ~(v(N0777_v));
  assign N0378_v = ~(((DAA_v&N0803_v)|O_IB_v));
  assign N0471_v = ~(N0856_v);
  assign N0916_v = ~(v(N0912_v));
  assign N0701_v = ~(L_v);
  assign N0678_v = ~((v(clk1_v)|N0699_v|N0685_v));
  assign N0435_v = ~(v(SC_v));
  assign N0622_v = ~((v(clk2_v)&((v(M12_v)|v(A12_v))&v(SC_v))));
  assign N0875_v = ~((((v(N0871_v)|v(N0889_v)|v(N0553_v))&v(N0556_v))|(v(N0871_v)&(v(N0889_v)&v(N0553_v)))));
  assign N0864_v = ~(N0499_v);
  assign N0641_v = ~(v(N0637_v));
  assign REG_RFSH_2_v = ~(v(N0642_v));
  assign ADD_0_v = ~((v(N0848_v)|v(N0846_v)|v(N0514_v)|v(N0847_v)));
  assign N0371_v = ~(N0346_v);
  assign N0358_v = ~((N0354_v|N0403_v|N0363_v|N0377_v|N0345_v|N0370_v));
  assign INC_ISZ_XCH_v = ~(((v(_OPR_2_v)|v(OPR_3_v)|v(_OPR_1_v))&(v(OPR_2_v)|v(_OPR_1_v)|v(_OPR_0_v)|v(_OPR_3_v))));
  assign STC_v = ~((v(OPA_2_v)|v(_OPA_3_v)|v(_OPA_1_v)|v(_OPE_v)|v(OPA_0_v)));
  assign TCC_v = ~((v(OPA_3_v)|v(_OPA_2_v)|v(_OPE_v)|v(_OPA_1_v)|v(_OPA_0_v)));
  assign CMA_v = ~((v(OPA_1_v)|v(_OPE_v)|v(_OPA_2_v)|v(OPA_0_v)|v(OPA_3_v)));
  assign RAL_v = ~((v(OPA_3_v)|v(_OPA_2_v)|v(OPA_1_v)|v(_OPE_v)|v(_OPA_0_v)));
  assign RAR_v = ~((v(_OPE_v)|v(_OPA_2_v)|v(OPA_0_v)|v(OPA_3_v)|v(_OPA_1_v)));
  assign IOW_v = ~((v(OPA_3_v)|v(_I_O_v)));
  assign N0364_v = ~(N0347_v);
  assign N0354_v = ~((N0346_v|N0347_v|N0356_v|N0355_v|N0350_v));
  assign N0802_v = ~(DAA_v);
  assign N0863_v = ~(N0498_v);
  assign N0541_v = ~(N0577_v);
  assign N0663_v = ~((N0664_v|v(N0676_v)));
  assign N0671_v = ~(v(D3_v));
  assign N1005_v = ~(N1004_v);
  assign N1001_v = ~(N1000_v);
  assign N0392_v = ~(v(N0776_v));
  assign N0627_v = ~(v(N0626_v));
  assign _INH_v = ~(INH_v);
  assign N0974_v = ~(v(N0635_v));
  assign N0983_v = ~(v(N0648_v));
  assign INC_ISZ_ADD_SUB_XCH_LD_v = ~(((v(OPR_3_v)|v(_OPR_2_v)|v(_OPR_1_v))&(v(OPR_2_v)|v(_OPR_3_v))));
  assign KBP_v = ~((v(_OPE_v)|v(OPA_1_v)|v(_OPA_3_v)|v(_OPA_2_v)|v(OPA_0_v)));
  assign N0447_v = ~((v(X12_v)|v(X32_v)));
  assign N0423_v = ~(v(clk2_v));
  assign N0764_v = ~((N0760_v|(v(N0752_v)&N0292_v)));
  assign ACC_0_v = ~((N0356_v|N0348_v|N0346_v|N0347_v));
  assign N0473_v = ~(N0858_v);
  assign O_IB_v = ~((v(OPA_3_v)|v(_OPE_v)));
  assign N0470_v = ~(N0855_v);
  assign ADDR_RFSH_0_v = ~(v(N0455_v));
  assign N0340_v = ~(v(N0332_v));
  assign N0472_v = ~(N0857_v);
  assign L_v = ~((N0703_v|N0703_v));
  assign N0430_v = ~(N0433_v);
  assign N0964_v = ~(v(N0342_v));
  assign N0682_v = ~(((v(X12_v)&(POC_v|IOR_v))|(v(A32_v)|v(M12_v))));
  assign N0799_v = ~(_SRC_v);
  assign N0726_v = ~(N0285_v);
  assign N0428_v = ~((v(A32_v)|(_INH_v&v(X12_v))));
  assign N0493_v = ~(IO_v);
  assign N0413_v = ~(((N0419_v&(v(SC_v)&v(X32_v)))|(N0399_v&N0397_v)));
  assign N0456_v = ~(ISZ_v);
  assign N0918_v = ~(v(N0914_v));
  assign DCL_1_v = ~((POC_v|v(N0765_v)));
  assign WRAB0_v = ~(N0547_v);
  assign N0580_v = ~(v(_OPA_0_v));
  assign SC_A12_CLK2_v = ~(N0649_v);
  assign N0547_v = ~((v(clk2_v)&((N0568_v&v(_OPA_0_v))|(N0564_v&v(M12_v)))));
  assign N0760_v = ~((v(N0752_v)|N0292_v));
  assign N0666_v = ~((v(d2_v)|v(N0676_v)));
  assign N0919_v = ~(v(N0545_v));
  assign N0928_v = ~(v(N0570_v));
  assign N0735_v = ~(v(N0715_v));
  assign N0314_v = ~(v(N0306_v));
  assign N0801_v = ~(N0431_v);
  assign N0356_v = ~(N0852_v);
  assign __X31__CLK2__v = ~(N0375_v);
  assign N0722_v = ~(N0283_v);
  assign N0573_v = ~(v(N0571_v));
  assign N0353_v = ~(DCL_v);
  assign N0995_v = ~(N0994_v);
  assign DCL_0_v = ~((POC_v|v(N0767_v)));
  assign N0403_v = ~((N0802_v|N0803_v));
  assign N0803_v = ~(((N0356_v&(N0348_v|N0347_v))|CY_1_v));
  assign N0667_v = ~((N0668_v|v(N0676_v)));
  assign REG_RFSH_0_v = ~(v(N0574_v));
  assign N0568_v = ~(N0603_v);
  assign N0534_v = ~(v(N0867_v));
  assign CLC_v = ~((v(OPA_3_v)|v(OPA_2_v)|v(_OPA_0_v)|v(_OPE_v)|v(OPA_1_v)));
  assign N0630_v = ~(((v(A32_v)|v(X12_v))&(v(SC_v)&v(clk2_v))));
  assign DAC_v = ~((v(OPA_1_v)|v(_OPE_v)|v(_OPA_3_v)|v(OPA_0_v)|v(OPA_2_v)));
  assign IAC_v = ~((v(_OPA_1_v)|v(_OPE_v)|v(OPA_2_v)|v(OPA_0_v)|v(OPA_3_v)));
  assign JUN2_JMS2_v = ~((v(OPR_1_v)|v(OPR_3_v)|v(_OPR_2_v)));
  assign CMC_v = ~((v(OPA_3_v)|v(OPA_2_v)|v(_OPA_0_v)|v(_OPA_1_v)|v(_OPE_v)));
  assign ADD_v = ~((v(OPR_2_v)|v(OPR_0_v)|v(_OPR_3_v)|v(OPR_1_v)));
  assign LDM_BBL_v = ~((v(OPR_1_v)|v(_OPR_3_v)|v(_OPR_2_v)));
  assign SBM_v = ~((v(OPA_2_v)|v(_I_O_v)|v(OPA_1_v)|v(_OPA_3_v)|v(OPA_0_v)));
  assign SUB_v = ~((v(OPR_1_v)|v(_OPR_0_v)|v(_OPR_3_v)|v(OPR_2_v)));
  assign N0402_v = ~(v(X32_v));
  assign N0804_v = ~(v(N0411_v));
  assign RADB0_v = ~((v(clk2_v)|N0416_v));
  assign N0955_v = ~(v(N0599_v));
  assign N0720_v = ~(N0282_v);
  assign N0965_v = ~(v(N0620_v));
  assign N0613_v = ~(v(N0646_v));
  assign N0783_v = ~(v(N0382_v));
  assign N0524_v = ~(((v(SC_v)&JIN_FIN_v)|(DC_v&(JUN_JMS_v|(N0528_v&JCN_ISZ_v)))));
  assign N0318_v = ~((((v(SC_v)&(v(X22_v)&JIN_FIN_v))|v(A22_v))|(v(M12_v)&((JCN_ISZ_v&N0322_v)|(N0310_v&JUN_JMS_v)))));
  assign N0859_v = ~(v(ACC_3_v));
  assign N0994_v = ~(N1009_v);
  assign N0998_v = ~(N1011_v);
  assign N0532_v = ~(v(N0880_v));
  assign N0531_v = ~(v(N0866_v));
  assign N0398_v = ~(v(clk2_v));
  assign N0608_v = ~((v(X12_v)&(FIN_FIM_SRC_JIN_v|(INC_ISZ_ADD_SUB_XCH_LD_v&v(_OPA_0_v)))));
  assign N0350_v = ~(KBP_v);
  assign N0346_v = ~(N0849_v);
  assign N0857_v = ~(v(ACC_1_v));
  assign N0884_v = ~(N0875_v);
  assign N0347_v = ~(N0850_v);
  assign N0996_v = ~(N1010_v);
  assign N0940_v = ~(v(N0939_v));
  assign N0664_v = ~((v(N0676_v)|v(d3_v)));
  assign N0805_v = ~(N0422_v);
  assign RADB2_v = ~((N0374_v|v(clk2_v)));
  assign N0490_v = ~(RAR_v);
  assign N0479_v = ~(IOR_v);
  assign N0477_v = ~(((v(A12_v)&IOR_v)|(N0480_v&N0479_v)));
  assign N0643_v = ~((v(SC_v)&v(A22_v)));
  assign N0540_v = ~(N0613_v);
  assign N0577_v = ~(v(N0617_v));
  assign N0542_v = ~(N0560_v);
  assign N0442_v = ~(INC_ISZ_v);
  assign IO_v = ~((v(_OPR_2_v)|v(_OPR_3_v)|v(OPR_0_v)|v(_OPR_1_v)));
  assign OPE_v = ~((v(_OPR_1_v)|v(_OPR_0_v)|v(_OPR_2_v)|v(_OPR_3_v)));
  assign JIN_FIN_v = ~((v(_OPR_1_v)|v(OPR_3_v)|v(_OPR_0_v)|v(OPR_2_v)));
  assign ISZ_v = ~((v(_OPR_1_v)|v(_OPR_0_v)|v(_OPR_2_v)|v(OPR_3_v)));
  assign JCN_v = ~((v(OPR_1_v)|v(OPR_2_v)|v(OPR_3_v)|v(_OPR_0_v)));
  assign FIM_SRC_v = ~((v(_OPR_1_v)|v(OPR_0_v)|v(OPR_2_v)|v(OPR_3_v)));
  assign N0766_v = ~(N0351_v);
  assign N0486_v = ~(((v(OPA_2_v)&ACC_0_v)|(v(OPA_1_v)&CY_1_v)|(v(OPA_0_v)&N0432_v)));
  assign N0942_v = ~(v(N0941_v));
  assign N0915_v = ~(v(N0911_v));
  assign N0992_v = ~(N1008_v);
  assign N0877_v = ~(((v(N0893_v)&(v(N0559_v)&v(N0873_v)))|(v(N0861_v)&(v(N0893_v)|v(N0873_v)|v(N0559_v)))));
  assign N0751_v = ~(DCL_0_v);
  assign N0326_v = ~((((v(SC_v)&(v(X32_v)&JIN_FIN_v))|v(A12_v))|(v(M22_v)&((N0310_v&JUN_JMS_v)|(JCN_ISZ_v&N0322_v)))));
  assign N0352_v = ~(v(X32_v));
  assign N0515_v = ~(CMA_v);
  assign N0379_v = ~(v(A12_v));
  assign N0365_v = ~(v(A22_v));
  assign N0708_v = ~(((N0278_v&v(clk1_v))|(v(M22_v)|v(M12_v))));
  assign N0724_v = ~(N0284_v);
  assign WRITE_ACC_1__v = ~((XCH_v|IAC_v|TCS_v|IOR_v|ADD_v|POC_v|KBP_v|TCC_v|CMA_v|SUB_v|LD_v|DAC_v|LDM_BBL_v|CLB_v|DAA_v));
  assign N1006_v = ~(N1015_v);
  assign N0658_v = ~((JUN2_JMS2_v|LDM_BBL_v));
  assign ADDR_PTR_0_v = ~(v(N0459_v));
  assign N0536_v = ~(v(N0882_v));
  assign N0535_v = ~(v(N0868_v));
  assign N1004_v = ~(N1014_v);
  assign N1002_v = ~(N1013_v);
  assign N0505_v = ~(v(N0466_v));
  assign ADM_v = ~((v(_OPA_3_v)|v(OPA_2_v)|v(_OPA_0_v)|v(_I_O_v)|v(_OPA_1_v)));
  assign N0946_v = ~(v(N0945_v));
  assign N0355_v = ~(N0348_v);
  assign JUN_JMS_v = ~((v(OPR_1_v)|v(OPR_3_v)|v(_OPR_2_v)));
  assign N0510_v = ~(OPE_v);
  assign N0876_v = ~(N0879_v);
  assign N0763_v = ~((N0758_v|(N0291_v&v(N0293_v))));
  assign N0537_v = ~(v(N0883_v));
  assign N0833_v = ~(v(N0440_v));
  assign N0377_v = ~((N0378_v&(N0347_v|N0346_v|N0348_v|N0350_v|N0356_v)));
  assign N0665_v = ~((N0666_v|v(N0676_v)));
  assign N0296_v = ~(N0280_v);
  assign N0357_v = ~((N0403_v|N0345_v|N0363_v|N0377_v));
  assign N0349_v = ~(N0356_v);
  assign N0561_v = ~(__FIN_X12__v);
  assign N0732_v = ~(N0317_v);
  assign N0502_v = ~(RAL_v);
  assign N0858_v = ~(v(ACC_2_v));
  assign N0734_v = ~(v(N0714_v));
  assign INC_ISZ_v = ~((v(_OPR_2_v)|v(_OPR_1_v)|v(OPR_3_v)|DC_v));
  assign N0528_v = ~(_CN_v);
  assign FIN_FIM_v = ~((v(OPR_2_v)|v(OPA_0_v)|v(_OPR_1_v)|v(OPR_3_v)));
  assign POC_v = ~(v(N0327_v));
  assign CY_1_v = ~(N0452_v);
  assign N0387_v = ~(v(N0778_v));
  assign WADB2_v = ~((N0304_v|N0300_v));
  assign CLK2_JMS_DC_M22_BBL_M22_X12_X22___v = ~((N0460_v|N0467_v));
  assign N0388_v = ~(v(N0779_v));
  assign _CN_v = ~(N0397_v);
  assign N0457_v = ~(v(N0475_v));
  assign N0588_v = ~(((INC_ISZ_ADD_SUB_XCH_LD_v&(N0580_v&v(X12_v)))|(FIN_FIM_SRC_JIN_v&v(X22_v))));
  assign N0754_v = ~((N0289_v|v(N0301_v)));
  assign N0437_v = ~(v(N0436_v));
  assign N0279_v = ~((v(M12_v)|v(A32_v)));
  assign ADD_GROUP_4__v = ~((ADD_v|ADM_v|TCS_v|TCC_v));
  assign N0467_v = ~(((JMS_v&(DC_v&v(M22_v)))|(BBL_v&(v(M22_v)|v(X22_v)|v(X12_v)))));
  assign N0997_v = ~(N0996_v);
  assign N0999_v = ~(N0998_v);
  assign TCS_v = ~((v(_OPA_3_v)|v(OPA_2_v)|v(_OPE_v)|v(OPA_1_v)|v(_OPA_0_v)));
  assign DCL_v = ~((v(_OPA_3_v)|v(_OPA_2_v)|v(_OPE_v)|v(_OPA_0_v)|v(OPA_1_v)));
  assign N0865_v = ~(N0500_v);
  assign JCN_ISZ_v = ~(((v(OPR_3_v)|v(_OPR_0_v))|((v(OPR_1_v)|v(OPR_2_v))&(v(_OPR_1_v)|v(_OPR_2_v)))));
  assign N0668_v = ~((v(N0676_v)|v(d1_v)));
  assign N0673_v = ~(v(D1_v));
  assign ADSR_v = ~((__X31__CLK2__v|N0490_v));
  assign N0359_v = ~((N0345_v|N0370_v|TCS_v|N0377_v));
  assign N0672_v = ~(v(D2_v));
  assign N0383_v = ~(v(X22_v));
  assign N0386_v = ~(v(N0774_v));
  assign N0419_v = ~(((N0456_v|ADD_0_v)&(((v(OPA_3_v)|N0486_v)&(v(_OPA_3_v)|N0487_v))|N0476_v)));
  assign READ_ACC_3__v = ~((ADD_v|DAA_v|RAR_v|DAC_v|IAC_v|SUB_v|RAL_v|ADM_v|SBM_v));
  assign N0862_v = ~(N0497_v);
  assign N0407_v = ~(N0414_v);
  assign N0307_v = ~((v(clk1_v)|N0711_v));
  assign N0300_v = ~(v(clk2_v));
  assign N0944_v = ~(v(N0943_v));
  assign N0546_v = ~((INC_GROUP_5__v|v(N0342_v)));
  assign N0878_v = ~(((v(N0870_v)&(v(N0887_v)&v(N0550_v)))|((v(N0550_v)|v(N0887_v)|v(N0870_v))&v(N0553_v))));
  assign ADC_CY_v = ~((WRITE_CARRY_2__v|N0477_v));
  assign N0879_v = ~(((v(N0872_v)&(v(N0891_v)&v(N0556_v)))|((v(N0556_v)|v(N0891_v)|v(N0872_v))&v(N0559_v))));
  assign N0474_v = ~(N0859_v);
  assign N0675_v = ~(((L_v&v(clk1_v))|(v(clk2_v)&N0685_v)));
  assign N0758_v = ~((v(N0293_v)|N0291_v));
  assign N0432_v = ~(v(test_v));
  assign N0784_v = ~(v(N0782_v));
  assign N0404_v = ~(N0405_v);
  assign N0399_v = ~(v(X32_v));
  assign REG_RFSH_1_v = ~(v(N0610_v));
  assign N0609_v = ~(v(N0600_v));
  assign N0450_v = ~(v(N0449_v));
  assign N0564_v = ~(N0590_v);
  assign N0348_v = ~(N0851_v);
  assign N0494_v = ~((v(clk2_v)&(v(X32_v)&_INH_v)));
  assign __INH__X32_CLK2_v = ~(N0494_v);
  assign N0674_v = ~(v(D0_v));
  assign N0670_v = ~((v(N0676_v)|v(d0_v)));
  assign N0669_v = ~((v(N0676_v)|N0670_v));
  assign ADSL_v = ~((__X31__CLK2__v|N0502_v));
  assign N0522_v = ~(v(clk1_v));
  assign N0677_v = ~(N0678_v);
  assign N0762_v = ~((N0756_v|(v(N0298_v)&N0290_v)));
  assign INC_GROUP_5__v = ~((IAC_v|INC_ISZ_v|STC_v));
  assign WRITE_CARRY_2__v = ~((CLC_v|POC_v|CMC_v|TCS_v|CLB_v|ADM_v|SUB_v|IAC_v|DAC_v|TCC_v|STC_v|SBM_v|ADD_v));
  assign N0856_v = ~(ACC_0_v);
  assign SC_A22_v = ~(N0643_v);
  assign SC_M22_CLK2_v = ~(N0679_v);
  assign N0679_v = ~((v(M22_v)&(v(SC_v)&v(clk2_v))));
  assign N0874_v = ~(N0878_v);
  assign N0533_v = ~(v(N0881_v));
  assign __FIN_X12__v = ~((v(X12_v)&(N0636_v&v(_OPA_0_v))));
  assign DCL_2_v = ~((POC_v|v(N0768_v)));
  assign N0749_v = ~(DCL_2_v);
  assign N0728_v = ~(N0286_v);
  assign N0487_v = ~(N0486_v);
  assign N0503_v = ~(v(N0463_v));
  assign N0368_v = ~(((N0343_v&N0352_v)|(v(SC_v)&((JUN_JMS_v|JCN_ISZ_v|FIN_FIM_v)&v(X32_v)))));
  assign N0705_v = ~(((POC_v|N0707_v)|(L_v&v(N0702_v))));
  assign N0733_v = ~(v(N0713_v));
  assign N0736_v = ~(v(N0716_v));
  assign N0797_v = ~(N0408_v);
  assign RADB1_v = ~((N0384_v|v(clk2_v)));
  assign _SRC_v = ~((v(OPA_0_v)&FIM_SRC_v));
  assign N0476_v = ~(JCN_v);
  assign N0316_v = ~(N0315_v);
  assign N0363_v = ~((N0346_v|N0364_v|N0356_v|N0350_v|N0348_v));
  assign WADB1_v = ~((N0300_v|N0318_v));
  assign N0711_v = ~(((N0732_v&(v(A32_v)|v(A22_v)))|v(A12_v)));
  assign N0451_v = ~(v(clk2_v));
  assign ADD_ACC_v = ~((WRITE_ACC_1__v|N0477_v));
  assign N1003_v = ~(N1002_v);
  assign WADB0_v = ~((N0300_v|N0326_v));


  spice_node_2 n_N0556(eclk, ereset, N0556_port_2,N0556_port_1, N0556_v);
  spice_node_1 n_S00819(eclk, ereset, S00819_port_0, S00819_v);
  spice_node_2 n_CY_ADA(eclk, ereset, CY_ADA_port_3,CY_ADA_port_4, CY_ADA_v);
  spice_node_2 n_N0449(eclk, ereset, N0449_port_1,N0449_port_7, N0449_v);
  spice_node_2 n_N0440(eclk, ereset, N0440_port_6,N0440_port_5, N0440_v);
  spice_node_2 n_N0444(eclk, ereset, N0444_port_12,N0444_port_13, N0444_v);
  spice_node_3 n_N0883(eclk, ereset, N0883_port_0,N0883_port_10,N0883_port_19, N0883_v);
  spice_node_3 n_N0880(eclk, ereset, N0880_port_0,N0880_port_10,N0880_port_19, N0880_v);
  spice_node_2 n_N0887(eclk, ereset, N0887_port_3,N0887_port_5, N0887_v);
  spice_node_2 n_N0530(eclk, ereset, N0530_port_4,N0530_port_5, N0530_v);
  spice_node_1 n_S00579(eclk, ereset, S00579_port_1, S00579_v);
  spice_node_1 n_S00578(eclk, ereset, S00578_port_1, S00578_v);
  spice_node_2 n_N0939(eclk, ereset, N0939_port_3,N0939_port_4, N0939_v);
  spice_node_1 n_S00757(eclk, ereset, S00757_port_1, S00757_v);
  spice_node_1 n_S00817(eclk, ereset, S00817_port_0, S00817_v);
  spice_node_2 n_SUB_GROUP_6_(eclk, ereset, SUB_GROUP_6__port_1,SUB_GROUP_6__port_12, SUB_GROUP_6__v);
  spice_node_2 n_N0332(eclk, ereset, N0332_port_5,N0332_port_11, N0332_v);
  spice_node_3 n__TMP_1(eclk, ereset, _TMP_1_port_2,_TMP_1_port_0,_TMP_1_port_1, _TMP_1_v);
  spice_node_3 n__TMP_0(eclk, ereset, _TMP_0_port_2,_TMP_0_port_0,_TMP_0_port_1, _TMP_0_v);
  spice_node_3 n__TMP_3(eclk, ereset, _TMP_3_port_2,_TMP_3_port_0,_TMP_3_port_1, _TMP_3_v);
  spice_node_3 n__TMP_2(eclk, ereset, _TMP_2_port_2,_TMP_2_port_0,_TMP_2_port_1, _TMP_2_v);
  spice_node_3 n_TMP_3(eclk, ereset, TMP_3_port_2,TMP_3_port_0,TMP_3_port_1, TMP_3_v);
  spice_node_3 n_TMP_2(eclk, ereset, TMP_2_port_2,TMP_2_port_0,TMP_2_port_1, TMP_2_v);
  spice_node_3 n_TMP_1(eclk, ereset, TMP_1_port_2,TMP_1_port_0,TMP_1_port_1, TMP_1_v);
  spice_node_3 n_TMP_0(eclk, ereset, TMP_0_port_2,TMP_0_port_0,TMP_0_port_1, TMP_0_v);
  spice_node_2 n_N0455(eclk, ereset, N0455_port_9,N0455_port_4, N0455_v);
  spice_node_2 n_N0459(eclk, ereset, N0459_port_8,N0459_port_5, N0459_v);
  spice_node_2 n_RRAB0(eclk, ereset, RRAB0_port_8,RRAB0_port_4, RRAB0_v);
  spice_node_2 n_RRAB1(eclk, ereset, RRAB1_port_8,RRAB1_port_4, RRAB1_v);
  spice_node_3 n_N0872(eclk, ereset, N0872_port_3,N0872_port_0,N0872_port_5, N0872_v);
  spice_node_1 n_S00699(eclk, ereset, S00699_port_1, S00699_v);
  spice_node_2 n__OPR_1(eclk, ereset, _OPR_1_port_15,_OPR_1_port_16, _OPR_1_v);
  spice_node_2 n__OPR_0(eclk, ereset, _OPR_0_port_10,_OPR_0_port_11, _OPR_0_v);
  spice_node_2 n_cm_rom(eclk, ereset, cm_rom_port_0,cm_rom_port_1, cm_rom_v);
  spice_node_2 n_cm_ram0(eclk, ereset, cm_ram0_port_0,cm_ram0_port_1, cm_ram0_v);
  spice_node_2 n_N0344(eclk, ereset, N0344_port_2,N0344_port_0, N0344_v);
  spice_node_3 n_d2(eclk, ereset, d2_port_2,d2_port_6,d2_port_5, d2_v);
  spice_node_3 n_d3(eclk, ereset, d3_port_1,d3_port_6,d3_port_5, d3_v);
  spice_node_2 n_N0617(eclk, ereset, N0617_port_2,N0617_port_1, N0617_v);
  spice_node_2 n_N0610(eclk, ereset, N0610_port_0,N0610_port_10, N0610_v);
  spice_node_2 n_ACC_ADA(eclk, ereset, ACC_ADA_port_7,ACC_ADA_port_5, ACC_ADA_v);
  spice_node_10 n___POC__CLK2_SC_A32_X12_(eclk, ereset, __POC__CLK2_SC_A32_X12__port_8,__POC__CLK2_SC_A32_X12__port_9,__POC__CLK2_SC_A32_X12__port_2,__POC__CLK2_SC_A32_X12__port_3,__POC__CLK2_SC_A32_X12__port_0,__POC__CLK2_SC_A32_X12__port_1,__POC__CLK2_SC_A32_X12__port_6,__POC__CLK2_SC_A32_X12__port_7,__POC__CLK2_SC_A32_X12__port_4,__POC__CLK2_SC_A32_X12__port_5, __POC__CLK2_SC_A32_X12__v);
  spice_node_2 n_N0342(eclk, ereset, N0342_port_0,N0342_port_1, N0342_v);
  spice_node_2 n_N0420(eclk, ereset, N0420_port_3,N0420_port_4, N0420_v);
  spice_node_2 n_N0424(eclk, ereset, N0424_port_12,N0424_port_13, N0424_v);
  spice_node_2 n_N0427(eclk, ereset, N0427_port_6,N0427_port_5, N0427_v);
  spice_node_2 n_N0426(eclk, ereset, N0426_port_12,N0426_port_13, N0426_v);
  spice_node_1 n_S00582(eclk, ereset, S00582_port_1, S00582_v);
  spice_node_1 n_S00583(eclk, ereset, S00583_port_1, S00583_v);
  spice_node_2 n_N0738(eclk, ereset, N0738_port_3,N0738_port_0, N0738_v);
  spice_node_5 n_CY(eclk, ereset, CY_port_2,CY_port_3,CY_port_1,CY_port_6,CY_port_5, CY_v);
  spice_node_1 n_S00685(eclk, ereset, S00685_port_0, S00685_v);
  spice_node_1 n_S00687(eclk, ereset, S00687_port_0, S00687_v);
  spice_node_1 n_S00689(eclk, ereset, S00689_port_0, S00689_v);
  spice_node_2 n_N0559(eclk, ereset, N0559_port_2,N0559_port_1, N0559_v);
  spice_node_3 n_N0558(eclk, ereset, N0558_port_2,N0558_port_0,N0558_port_1, N0558_v);
  spice_node_3 n_N0882(eclk, ereset, N0882_port_1,N0882_port_10,N0882_port_19, N0882_v);
  spice_node_3 n_N0881(eclk, ereset, N0881_port_0,N0881_port_10,N0881_port_19, N0881_v);
  spice_node_1 n_S00731(eclk, ereset, S00731_port_1, S00731_v);
  spice_node_1 n_S00836(eclk, ereset, S00836_port_0, S00836_v);
  spice_node_1 n_S00724(eclk, ereset, S00724_port_1, S00724_v);
  spice_node_2 n_N0642(eclk, ereset, N0642_port_0,N0642_port_6, N0642_v);
  spice_node_1 n_S00833(eclk, ereset, S00833_port_0, S00833_v);
  spice_node_2 n_N0891(eclk, ereset, N0891_port_4,N0891_port_5, N0891_v);
  spice_node_2 n_N0436(eclk, ereset, N0436_port_8,N0436_port_0, N0436_v);
  spice_node_2 n_N0434(eclk, ereset, N0434_port_12,N0434_port_13, N0434_v);
  spice_node_2 n_N0439(eclk, ereset, N0439_port_12,N0439_port_13, N0439_v);
  spice_node_1 n_reset(eclk, ereset, reset_port_2, reset_v);
  spice_node_2 n_N0943(eclk, ereset, N0943_port_3,N0943_port_4, N0943_v);
  spice_node_2 n_N0893(eclk, ereset, N0893_port_4,N0893_port_5, N0893_v);
  spice_node_3 n_N0548(eclk, ereset, N0548_port_2,N0548_port_0,N0548_port_1, N0548_v);
  spice_node_3 n_N0549(eclk, ereset, N0549_port_2,N0549_port_0,N0549_port_1, N0549_v);
  spice_node_1 n_S00839(eclk, ereset, S00839_port_1, S00839_v);
  spice_node_2 n_N0543(eclk, ereset, N0543_port_8,N0543_port_9, N0543_v);
  spice_node_2 n_N0544(eclk, ereset, N0544_port_8,N0544_port_9, N0544_v);
  spice_node_2 n_N0545(eclk, ereset, N0545_port_8,N0545_port_7, N0545_v);
  spice_node_2 n_N0466(eclk, ereset, N0466_port_2,N0466_port_11, N0466_v);
  spice_node_2 n__OPR_3(eclk, ereset, _OPR_3_port_10,_OPR_3_port_11, _OPR_3_v);
  spice_node_2 n__OPR_2(eclk, ereset, _OPR_2_port_12,_OPR_2_port_13, _OPR_2_v);
  spice_node_4 n_N0513(eclk, ereset, N0513_port_2,N0513_port_3,N0513_port_0,N0513_port_1, N0513_v);
  spice_node_2 n_M22(eclk, ereset, M22_port_10,M22_port_11, M22_v);
  spice_node_2 n_SC_A22_M22_CLK2(eclk, ereset, SC_A22_M22_CLK2_port_8,SC_A22_M22_CLK2_port_9, SC_A22_M22_CLK2_v);
  spice_node_2 n_OPA_IB(eclk, ereset, OPA_IB_port_6,OPA_IB_port_7, OPA_IB_v);
  spice_node_1 n_S00654(eclk, ereset, S00654_port_1, S00654_v);
  spice_node_1 n_S00818(eclk, ereset, S00818_port_0, S00818_v);
  spice_node_1 n_S00729(eclk, ereset, S00729_port_1, S00729_v);
  spice_node_2 n_N0409(eclk, ereset, N0409_port_3,N0409_port_4, N0409_v);
  spice_node_2 n_N0406(eclk, ereset, N0406_port_12,N0406_port_13, N0406_v);
  spice_node_1 n_S00678(eclk, ereset, S00678_port_1, S00678_v);
  spice_node_2 n_N0713(eclk, ereset, N0713_port_2,N0713_port_5, N0713_v);
  spice_node_2 n_N0710(eclk, ereset, N0710_port_2,N0710_port_1, N0710_v);
  spice_node_2 n_N0717(eclk, ereset, N0717_port_3,N0717_port_5, N0717_v);
  spice_node_2 n_N0715(eclk, ereset, N0715_port_4,N0715_port_5, N0715_v);
  spice_node_2 n_N0714(eclk, ereset, N0714_port_2,N0714_port_5, N0714_v);
  spice_node_2 n_N0574(eclk, ereset, N0574_port_0,N0574_port_11, N0574_v);
  spice_node_2 n_N0571(eclk, ereset, N0571_port_9,N0571_port_0, N0571_v);
  spice_node_2 n_N0570(eclk, ereset, N0570_port_8,N0570_port_7, N0570_v);
  spice_node_1 n_S00825(eclk, ereset, S00825_port_0, S00825_v);
  spice_node_1 n_S00531(eclk, ereset, S00531_port_0, S00531_v);
  spice_node_1 n_S00536(eclk, ereset, S00536_port_1, S00536_v);
  spice_node_2 n_N0889(eclk, ereset, N0889_port_4,N0889_port_5, N0889_v);
  spice_node_6 n_N0514(eclk, ereset, N0514_port_2,N0514_port_3,N0514_port_0,N0514_port_6,N0514_port_4,N0514_port_5, N0514_v);
  spice_node_6 n_N0848(eclk, ereset, N0848_port_2,N0848_port_0,N0848_port_1,N0848_port_6,N0848_port_4,N0848_port_5, N0848_v);
  spice_node_2 n_M12(eclk, ereset, M12_port_10,M12_port_11, M12_v);
  spice_node_2 n_N0381(eclk, ereset, N0381_port_12,N0381_port_13, N0381_v);
  spice_node_2 n_N0382(eclk, ereset, N0382_port_6,N0382_port_5, N0382_v);
  spice_node_2 n_N0410(eclk, ereset, N0410_port_12,N0410_port_13, N0410_v);
  spice_node_2 n_N0411(eclk, ereset, N0411_port_6,N0411_port_5, N0411_v);
  spice_node_2 n_N0415(eclk, ereset, N0415_port_8,N0415_port_0, N0415_v);
  spice_node_2 n__COM(eclk, ereset, _COM_port_0,_COM_port_1, _COM_v);
  spice_node_2 n_N0700(eclk, ereset, N0700_port_2,N0700_port_3, N0700_v);
  spice_node_2 n_N0702(eclk, ereset, N0702_port_0,N0702_port_1, N0702_v);
  spice_node_13 n_D2(eclk, ereset, D2_port_13,D2_port_14,D2_port_15,D2_port_16,D2_port_17,D2_port_19,D2_port_9,D2_port_2,D2_port_3,D2_port_1,D2_port_6,D2_port_7,D2_port_5, D2_v);
  spice_node_13 n_D3(eclk, ereset, D3_port_13,D3_port_14,D3_port_15,D3_port_16,D3_port_17,D3_port_19,D3_port_9,D3_port_3,D3_port_0,D3_port_1,D3_port_6,D3_port_7,D3_port_5, D3_v);
  spice_node_13 n_D0(eclk, ereset, D0_port_11,D0_port_12,D0_port_13,D0_port_14,D0_port_15,D0_port_16,D0_port_19,D0_port_8,D0_port_3,D0_port_1,D0_port_6,D0_port_4,D0_port_5, D0_v);
  spice_node_13 n_D1(eclk, ereset, D1_port_12,D1_port_13,D1_port_14,D1_port_15,D1_port_16,D1_port_19,D1_port_9,D1_port_2,D1_port_3,D1_port_1,D1_port_7,D1_port_4,D1_port_5, D1_v);
  spice_node_2 n_N0565(eclk, ereset, N0565_port_8,N0565_port_9, N0565_v);
  spice_node_2 n_N0569(eclk, ereset, N0569_port_8,N0569_port_9, N0569_v);
  spice_node_1 n_S00814(eclk, ereset, S00814_port_0, S00814_v);
  spice_node_1 n_S00676(eclk, ereset, S00676_port_0, S00676_v);
  spice_node_2 n__OPA_0(eclk, ereset, _OPA_0_port_13,_OPA_0_port_14, _OPA_0_v);
  spice_node_2 n__OPA_2(eclk, ereset, _OPA_2_port_6,_OPA_2_port_7, _OPA_2_v);
  spice_node_2 n__OPA_3(eclk, ereset, _OPA_3_port_10,_OPA_3_port_11, _OPA_3_v);
  spice_node_2 n_N0646(eclk, ereset, N0646_port_2,N0646_port_1, N0646_v);
  spice_node_6 n____SC__JIN_FIN__CLK1_M11_X21_INH_(eclk, ereset, ___SC__JIN_FIN__CLK1_M11_X21_INH__port_2,___SC__JIN_FIN__CLK1_M11_X21_INH__port_3,___SC__JIN_FIN__CLK1_M11_X21_INH__port_0,___SC__JIN_FIN__CLK1_M11_X21_INH__port_1,___SC__JIN_FIN__CLK1_M11_X21_INH__port_4,___SC__JIN_FIN__CLK1_M11_X21_INH__port_5, ___SC__JIN_FIN__CLK1_M11_X21_INH__v);
  spice_node_2 n_N0941(eclk, ereset, N0941_port_3,N0941_port_4, N0941_v);
  spice_node_3 n_N0861(eclk, ereset, N0861_port_2,N0861_port_3,N0861_port_0, N0861_v);
  spice_node_3 n_N0866(eclk, ereset, N0866_port_0,N0866_port_10,N0866_port_19, N0866_v);
  spice_node_3 n_N0911(eclk, ereset, N0911_port_2,N0911_port_0,N0911_port_1, N0911_v);
  spice_node_2 n_N0621(eclk, ereset, N0621_port_0,N0621_port_1, N0621_v);
  spice_node_3 n_N0771(eclk, ereset, N0771_port_1,N0771_port_6,N0771_port_11, N0771_v);
  spice_node_3 n_N0770(eclk, ereset, N0770_port_2,N0770_port_6,N0770_port_11, N0770_v);
  spice_node_3 n_N0773(eclk, ereset, N0773_port_1,N0773_port_6,N0773_port_11, N0773_v);
  spice_node_3 n_N0772(eclk, ereset, N0772_port_1,N0772_port_6,N0772_port_11, N0772_v);
  spice_node_3 n_N0775(eclk, ereset, N0775_port_0,N0775_port_6,N0775_port_11, N0775_v);
  spice_node_3 n_N0774(eclk, ereset, N0774_port_0,N0774_port_6,N0774_port_11, N0774_v);
  spice_node_3 n_N0777(eclk, ereset, N0777_port_1,N0777_port_6,N0777_port_11, N0777_v);
  spice_node_3 n_N0776(eclk, ereset, N0776_port_0,N0776_port_6,N0776_port_11, N0776_v);
  spice_node_3 n_N0779(eclk, ereset, N0779_port_0,N0779_port_6,N0779_port_11, N0779_v);
  spice_node_3 n_N0778(eclk, ereset, N0778_port_0,N0778_port_6,N0778_port_11, N0778_v);
  spice_node_2 n_N0626(eclk, ereset, N0626_port_1,N0626_port_5, N0626_v);
  spice_node_3 n_N0914(eclk, ereset, N0914_port_2,N0914_port_0,N0914_port_1, N0914_v);
  spice_node_1 n_test(eclk, ereset, test_port_2, test_v);
  spice_node_1 n_S00834(eclk, ereset, S00834_port_0, S00834_v);
  spice_node_1 n_S00804(eclk, ereset, S00804_port_0, S00804_v);
  spice_node_2 n_N0599(eclk, ereset, N0599_port_8,N0599_port_7, N0599_v);
  spice_node_2 n_N0598(eclk, ereset, N0598_port_8,N0598_port_9, N0598_v);
  spice_node_1 n_S00801(eclk, ereset, S00801_port_1, S00801_v);
  spice_node_1 n_S00800(eclk, ereset, S00800_port_0, S00800_v);
  spice_node_2 n_N0591(eclk, ereset, N0591_port_8,N0591_port_9, N0591_v);
  spice_node_2 n_N0606(eclk, ereset, N0606_port_0,N0606_port_1, N0606_v);
  spice_node_2 n_N0600(eclk, ereset, N0600_port_9,N0600_port_0, N0600_v);
  spice_node_2 n___INH__X11_X31_CLK1(eclk, ereset, __INH__X11_X31_CLK1_port_12,__INH__X11_X31_CLK1_port_16, __INH__X11_X31_CLK1_v);
  spice_node_1 n_S00761(eclk, ereset, S00761_port_0, S00761_v);
  spice_node_1 n_S00781(eclk, ereset, S00781_port_1, S00781_v);
  spice_node_2 n_CY_ADAC(eclk, ereset, CY_ADAC_port_2,CY_ADAC_port_4, CY_ADAC_v);
  spice_node_10 n_CLK2_SC_A12_M12_(eclk, ereset, CLK2_SC_A12_M12__port_8,CLK2_SC_A12_M12__port_9,CLK2_SC_A12_M12__port_2,CLK2_SC_A12_M12__port_3,CLK2_SC_A12_M12__port_0,CLK2_SC_A12_M12__port_1,CLK2_SC_A12_M12__port_6,CLK2_SC_A12_M12__port_7,CLK2_SC_A12_M12__port_4,CLK2_SC_A12_M12__port_5, CLK2_SC_A12_M12__v);
  spice_node_2 n_N0293(eclk, ereset, N0293_port_2,N0293_port_3, N0293_v);
  spice_node_2 n_N0297(eclk, ereset, N0297_port_0,N0297_port_1, N0297_v);
  spice_node_4 n_N0294(eclk, ereset, N0294_port_2,N0294_port_3,N0294_port_4,N0294_port_5, N0294_v);
  spice_node_2 n_N0298(eclk, ereset, N0298_port_0,N0298_port_6, N0298_v);
  spice_node_2 n_N0767(eclk, ereset, N0767_port_2,N0767_port_0, N0767_v);
  spice_node_2 n_N0765(eclk, ereset, N0765_port_2,N0765_port_1, N0765_v);
  spice_node_2 n_N0768(eclk, ereset, N0768_port_2,N0768_port_0, N0768_v);
  spice_node_2 n_N0769(eclk, ereset, N0769_port_0,N0769_port_4, N0769_v);
  spice_node_2 n_sync(eclk, ereset, sync_port_0,sync_port_1, sync_v);
  spice_node_2 n_N0584(eclk, ereset, N0584_port_8,N0584_port_7, N0584_v);
  spice_node_2 n_N0582(eclk, ereset, N0582_port_2,N0582_port_1, N0582_v);
  spice_node_2 n_N0583(eclk, ereset, N0583_port_8,N0583_port_9, N0583_v);
  spice_node_2 n_N0581(eclk, ereset, N0581_port_8,N0581_port_9, N0581_v);
  spice_node_2 n_N0619(eclk, ereset, N0619_port_8,N0619_port_9, N0619_v);
  spice_node_2 n_N0616(eclk, ereset, N0616_port_8,N0616_port_9, N0616_v);
  spice_node_1 n_S00612(eclk, ereset, S00612_port_1, S00612_v);
  spice_node_1 n_S00613(eclk, ereset, S00613_port_0, S00613_v);
  spice_node_1 n_S00580(eclk, ereset, S00580_port_1, S00580_v);
  spice_node_1 n_S00581(eclk, ereset, S00581_port_1, S00581_v);
  spice_node_1 n_S00584(eclk, ereset, S00584_port_1, S00584_v);
  spice_node_1 n_S00585(eclk, ereset, S00585_port_1, S00585_v);
  spice_node_2 n_cm_ram2(eclk, ereset, cm_ram2_port_0,cm_ram2_port_1, cm_ram2_v);
  spice_node_1 n_S00725(eclk, ereset, S00725_port_0, S00725_v);
  spice_node_2 n_SC(eclk, ereset, SC_port_13,SC_port_4, SC_v);
  spice_node_2 n_N0620(eclk, ereset, N0620_port_8,N0620_port_7, N0620_v);
  spice_node_2 n_N0854(eclk, ereset, N0854_port_0,N0854_port_6, N0854_v);
  spice_node_2 n__OPE(eclk, ereset, _OPE_port_0,_OPE_port_1, _OPE_v);
  spice_node_2 n_N0752(eclk, ereset, N0752_port_3,N0752_port_0, N0752_v);
  spice_node_1 n_S00690(eclk, ereset, S00690_port_1, S00690_v);
  spice_node_1 n_S00609(eclk, ereset, S00609_port_0, S00609_v);
  spice_node_1 n_S00601(eclk, ereset, S00601_port_1, S00601_v);
  spice_node_1 n_S00600(eclk, ereset, S00600_port_1, S00600_v);
  spice_node_1 n_S00599(eclk, ereset, S00599_port_1, S00599_v);
  spice_node_1 n_S00598(eclk, ereset, S00598_port_1, S00598_v);
  spice_node_2 n_A32(eclk, ereset, A32_port_8,A32_port_9, A32_v);
  spice_node_1 n_S00734(eclk, ereset, S00734_port_1, S00734_v);
  spice_node_1 n_S00732(eclk, ereset, S00732_port_1, S00732_v);
  spice_node_6 n___POC_CLK2_X12_X32__INH(eclk, ereset, __POC_CLK2_X12_X32__INH_port_2,__POC_CLK2_X12_X32__INH_port_3,__POC_CLK2_X12_X32__INH_port_0,__POC_CLK2_X12_X32__INH_port_1,__POC_CLK2_X12_X32__INH_port_4,__POC_CLK2_X12_X32__INH_port_5, __POC_CLK2_X12_X32__INH_v);
  spice_node_2 n_M12_M22_CLK1__M11_M12_(eclk, ereset, M12_M22_CLK1__M11_M12__port_8,M12_M22_CLK1__M11_M12__port_9, M12_M22_CLK1__M11_M12__v);
  spice_node_1 n_S00828(eclk, ereset, S00828_port_1, S00828_v);
  spice_node_6 n_N0847(eclk, ereset, N0847_port_3,N0847_port_0,N0847_port_1,N0847_port_6,N0847_port_4,N0847_port_5, N0847_v);
  spice_node_2 n_ACC_ADAC(eclk, ereset, ACC_ADAC_port_3,ACC_ADAC_port_7, ACC_ADAC_v);
  spice_node_2 n__OPA_1(eclk, ereset, _OPA_1_port_8,_OPA_1_port_7, _OPA_1_v);
  spice_node_4 n_ACC_3(eclk, ereset, ACC_3_port_3,ACC_3_port_0,ACC_3_port_1,ACC_3_port_4, ACC_3_v);
  spice_node_4 n_ACC_2(eclk, ereset, ACC_2_port_2,ACC_2_port_3,ACC_2_port_0,ACC_2_port_4, ACC_2_v);
  spice_node_4 n_ACC_1(eclk, ereset, ACC_1_port_3,ACC_1_port_0,ACC_1_port_1,ACC_1_port_4, ACC_1_v);
  spice_node_2 n_N0945(eclk, ereset, N0945_port_3,N0945_port_4, N0945_v);
  spice_node_2 n_cm_ram1(eclk, ereset, cm_ram1_port_0,cm_ram1_port_1, cm_ram1_v);
  spice_node_2 n_cm_ram3(eclk, ereset, cm_ram3_port_0,cm_ram3_port_1, cm_ram3_v);
  spice_node_2 n_N0748(eclk, ereset, N0748_port_2,N0748_port_1, N0748_v);
  spice_node_2 n_N0740(eclk, ereset, N0740_port_2,N0740_port_1, N0740_v);
  spice_node_2 n_N0741(eclk, ereset, N0741_port_0,N0741_port_1, N0741_v);
  spice_node_2 n_N0742(eclk, ereset, N0742_port_2,N0742_port_1, N0742_v);
  spice_node_2 n_N0743(eclk, ereset, N0743_port_2,N0743_port_1, N0743_v);
  spice_node_2 n_N0744(eclk, ereset, N0744_port_2,N0744_port_1, N0744_v);
  spice_node_2 n_N0745(eclk, ereset, N0745_port_2,N0745_port_1, N0745_v);
  spice_node_2 n_N0746(eclk, ereset, N0746_port_2,N0746_port_1, N0746_v);
  spice_node_2 n_N0747(eclk, ereset, N0747_port_2,N0747_port_1, N0747_v);
  spice_node_2 n_N0676(eclk, ereset, N0676_port_0,N0676_port_1, N0676_v);
  spice_node_2 n_N0634(eclk, ereset, N0634_port_8,N0634_port_9, N0634_v);
  spice_node_2 n_N0635(eclk, ereset, N0635_port_8,N0635_port_7, N0635_v);
  spice_node_2 n_N0637(eclk, ereset, N0637_port_0,N0637_port_7, N0637_v);
  spice_node_2 n_N0632(eclk, ereset, N0632_port_8,N0632_port_9, N0632_v);
  spice_node_2 n_ACB_IB(eclk, ereset, ACB_IB_port_8,ACB_IB_port_2, ACB_IB_v);
  spice_node_2 n_A22(eclk, ereset, A22_port_8,A22_port_9, A22_v);
  spice_node_1 n_S00709(eclk, ereset, S00709_port_1, S00709_v);
  spice_node_2 n_N0690(eclk, ereset, N0690_port_0,N0690_port_5, N0690_v);
  spice_node_3 n_N0913(eclk, ereset, N0913_port_2,N0913_port_0,N0913_port_1, N0913_v);
  spice_node_3 n_N0912(eclk, ereset, N0912_port_2,N0912_port_0,N0912_port_1, N0912_v);
  spice_node_1 n_S00564(eclk, ereset, S00564_port_0, S00564_v);
  spice_node_2 n_N0693(eclk, ereset, N0693_port_3,N0693_port_6, N0693_v);
  spice_node_1 n_S00803(eclk, ereset, S00803_port_1, S00803_v);
  spice_node_2 n_N0605(eclk, ereset, N0605_port_0,N0605_port_1, N0605_v);
  spice_node_2 n_N0604(eclk, ereset, N0604_port_0,N0604_port_1, N0604_v);
  spice_node_2 n_N0607(eclk, ereset, N0607_port_0,N0607_port_1, N0607_v);
  spice_node_2 n_OPR_3(eclk, ereset, OPR_3_port_14,OPR_3_port_15, OPR_3_v);
  spice_node_2 n_ADD_IB(eclk, ereset, ADD_IB_port_2,ADD_IB_port_7, ADD_IB_v);
  spice_node_1 n_clk1(eclk, ereset, clk1_port_28, clk1_v);
  spice_node_1 n_clk2(eclk, ereset, clk2_port_51, clk2_v);
  spice_node_2 n_N0645(eclk, ereset, N0645_port_8,N0645_port_9, N0645_v);
  spice_node_2 n_N0647(eclk, ereset, N0647_port_8,N0647_port_9, N0647_v);
  spice_node_2 n_N0648(eclk, ereset, N0648_port_8,N0648_port_7, N0648_v);
  spice_node_1 n_S00840(eclk, ereset, S00840_port_1, S00840_v);
  spice_node_3 n_N0869(eclk, ereset, N0869_port_0,N0869_port_10,N0869_port_19, N0869_v);
  spice_node_3 n_N0868(eclk, ereset, N0868_port_0,N0868_port_10,N0868_port_19, N0868_v);
  spice_node_3 n_N0867(eclk, ereset, N0867_port_0,N0867_port_10,N0867_port_19, N0867_v);
  spice_node_2 n_A12(eclk, ereset, A12_port_9,A12_port_10, A12_v);
  spice_node_1 n_S00716(eclk, ereset, S00716_port_1, S00716_v);
  spice_node_1 n_S00710(eclk, ereset, S00710_port_0, S00710_v);
  spice_node_1 n_S00620(eclk, ereset, S00620_port_1, S00620_v);
  spice_node_1 n_S00627(eclk, ereset, S00627_port_1, S00627_v);
  spice_node_1 n_S00624(eclk, ereset, S00624_port_1, S00624_v);
  spice_node_1 n_S00628(eclk, ereset, S00628_port_0, S00628_v);
  spice_node_2 n__I_O(eclk, ereset, _I_O_port_0,_I_O_port_1, _I_O_v);
  spice_node_3 n_d0(eclk, ereset, d0_port_2,d0_port_6,d0_port_5, d0_v);
  spice_node_3 n_d1(eclk, ereset, d1_port_2,d1_port_7,d1_port_5, d1_v);
  spice_node_2 n_N0937(eclk, ereset, N0937_port_6,N0937_port_7, N0937_v);
  spice_node_2 n_OPR_1(eclk, ereset, OPR_1_port_9,OPR_1_port_10, OPR_1_v);
  spice_node_2 n_OPR_0(eclk, ereset, OPR_0_port_3,OPR_0_port_6, OPR_0_v);
  spice_node_2 n_OPR_2(eclk, ereset, OPR_2_port_14,OPR_2_port_8, OPR_2_v);
  spice_node_3 n_N0780(eclk, ereset, N0780_port_0,N0780_port_6,N0780_port_11, N0780_v);
  spice_node_3 n_N0781(eclk, ereset, N0781_port_0,N0781_port_6,N0781_port_11, N0781_v);
  spice_node_2 n_N0782(eclk, ereset, N0782_port_8,N0782_port_5, N0782_v);
  spice_node_2 n_N0301(eclk, ereset, N0301_port_2,N0301_port_7, N0301_v);
  spice_node_3 n_N0305(eclk, ereset, N0305_port_2,N0305_port_1,N0305_port_4, N0305_v);
  spice_node_2 n_N0306(eclk, ereset, N0306_port_0,N0306_port_1, N0306_v);
  spice_node_2 n_X12(eclk, ereset, X12_port_12,X12_port_13, X12_v);
  spice_node_2 n_N0657(eclk, ereset, N0657_port_8,N0657_port_9, N0657_v);
  spice_node_1 n_S00762(eclk, ereset, S00762_port_1, S00762_v);
  spice_node_2 n_N0716(eclk, ereset, N0716_port_7,N0716_port_4, N0716_v);
  spice_node_3 n_OPA_2(eclk, ereset, OPA_2_port_0,OPA_2_port_4,OPA_2_port_13, OPA_2_v);
  spice_node_3 n_OPA_3(eclk, ereset, OPA_3_port_2,OPA_3_port_0,OPA_3_port_13, OPA_3_v);
  spice_node_3 n_OPA_0(eclk, ereset, OPA_0_port_11,OPA_0_port_12,OPA_0_port_13, OPA_0_v);
  spice_node_3 n_N0873(eclk, ereset, N0873_port_0,N0873_port_4,N0873_port_5, N0873_v);
  spice_node_3 n_N0870(eclk, ereset, N0870_port_2,N0870_port_0,N0870_port_6, N0870_v);
  spice_node_3 n_N0871(eclk, ereset, N0871_port_0,N0871_port_6,N0871_port_5, N0871_v);
  spice_node_3 n_OPA_1(eclk, ereset, OPA_1_port_10,OPA_1_port_11,OPA_1_port_12, OPA_1_v);
  spice_node_1 n_S00778(eclk, ereset, S00778_port_0, S00778_v);
  spice_node_2 n_N0696(eclk, ereset, N0696_port_3,N0696_port_6, N0696_v);
  spice_node_2 n_N0469(eclk, ereset, N0469_port_1,N0469_port_7, N0469_v);
  spice_node_2 n_N0464(eclk, ereset, N0464_port_3,N0464_port_6, N0464_v);
  spice_node_2 n_N0461(eclk, ereset, N0461_port_2,N0461_port_6, N0461_v);
  spice_node_2 n_N0463(eclk, ereset, N0463_port_2,N0463_port_11, N0463_v);
  spice_node_2 n_N0687(eclk, ereset, N0687_port_0,N0687_port_5, N0687_v);
  spice_node_1 n_S00557(eclk, ereset, S00557_port_1, S00557_v);
  spice_node_2 n_N0689(eclk, ereset, N0689_port_0,N0689_port_4, N0689_v);
  spice_node_2 n_X22(eclk, ereset, X22_port_6,X22_port_7, X22_v);
  spice_node_6 n_N0846(eclk, ereset, N0846_port_2,N0846_port_0,N0846_port_1,N0846_port_6,N0846_port_4,N0846_port_5, N0846_v);
  spice_node_2 n_N0692(eclk, ereset, N0692_port_0,N0692_port_5, N0692_v);
  spice_node_2 n_N0695(eclk, ereset, N0695_port_3,N0695_port_4, N0695_v);
  spice_node_2 n_N0475(eclk, ereset, N0475_port_0,N0475_port_7, N0475_v);
  spice_node_2 n_X32(eclk, ereset, X32_port_11,X32_port_12, X32_v);
  spice_node_2 n_N0698(eclk, ereset, N0698_port_3,N0698_port_5, N0698_v);
  spice_node_1 n_S00740(eclk, ereset, S00740_port_0, S00740_v);
  spice_node_1 n_S00766(eclk, ereset, S00766_port_0, S00766_v);
  spice_node_3 n_N0551(eclk, ereset, N0551_port_2,N0551_port_0,N0551_port_1, N0551_v);
  spice_node_1 n_S00767(eclk, ereset, S00767_port_0, S00767_v);
  spice_node_4 n_N0550(eclk, ereset, N0550_port_2,N0550_port_3,N0550_port_0,N0550_port_1, N0550_v);
  spice_node_2 n_N0327(eclk, ereset, N0327_port_6,N0327_port_4, N0327_v);
  spice_node_1 n_S00764(eclk, ereset, S00764_port_1, S00764_v);
  spice_node_2 n_N0553(eclk, ereset, N0553_port_2,N0553_port_1, N0553_v);
  spice_node_1 n_S00765(eclk, ereset, S00765_port_0, S00765_v);
  spice_node_3 n_N0552(eclk, ereset, N0552_port_2,N0552_port_0,N0552_port_1, N0552_v);
  spice_node_2 n_N0529(eclk, ereset, N0529_port_8,N0529_port_9, N0529_v);
  spice_node_3 n_N0555(eclk, ereset, N0555_port_2,N0555_port_0,N0555_port_1, N0555_v);
  spice_node_1 n_S00835(eclk, ereset, S00835_port_0, S00835_v);
  spice_node_3 n_N0554(eclk, ereset, N0554_port_2,N0554_port_0,N0554_port_1, N0554_v);
  spice_node_3 n_N0557(eclk, ereset, N0557_port_2,N0557_port_0,N0557_port_1, N0557_v);

endmodule

module spice_node_0(input eclk,ereset, output signed [`W-1:0] v);
  assign v = 0;
endmodule

module spice_node_1(input eclk,ereset, input signed [`W-1:0] i0, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_2(input eclk,ereset, input signed [`W-1:0] i0,i1, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_3(input eclk,ereset, input signed [`W-1:0] i0,i1,i2, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_4(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_5(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_6(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_10(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6+i7+i8+i9;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

module spice_node_13(input eclk,ereset, input signed [`W-1:0] i0,i1,i2,i3,i4,i5,i6,i7,i8,i9,i10,i11,i12, output reg signed [`W-1:0] v);
  wire signed [`W-1:0] i = i0+i1+i2+i3+i4+i5+i6+i7+i8+i9+i10+i11+i12;

  always @(posedge eclk)
    if (ereset)
      v <= 0;
    else
      v <= v + i;

endmodule

