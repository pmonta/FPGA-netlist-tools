module rom_6502(
  input eclk,ereset,
  input [15:0] ab,
  output reg [7:0] d
);

  reg [7:0] x;

  always @(posedge eclk)
    if (ereset)
      d <= 0;
    else
      d <= x;

  always @*
    case (ab[12:0])
      13'd0: x = 8'h4c;
      13'd1: x = 8'hb0;
      13'd2: x = 8'he2;
      13'd3: x = 8'had;
      13'd4: x = 8'h11;
      13'd5: x = 8'hd0;
      13'd6: x = 8'h10;
      13'd7: x = 8'hfb;
      13'd8: x = 8'had;
      13'd9: x = 8'h10;
      13'd10: x = 8'hd0;
      13'd11: x = 8'h60;
      13'd12: x = 8'h8a;
      13'd13: x = 8'h29;
      13'd14: x = 8'h20;
      13'd15: x = 8'hf0;
      13'd16: x = 8'h23;
      13'd17: x = 8'ha9;
      13'd18: x = 8'ha0;
      13'd19: x = 8'h85;
      13'd20: x = 8'he4;
      13'd21: x = 8'h4c;
      13'd22: x = 8'hc9;
      13'd23: x = 8'he3;
      13'd24: x = 8'ha9;
      13'd25: x = 8'h20;
      13'd26: x = 8'hc5;
      13'd27: x = 8'h24;
      13'd28: x = 8'hb0;
      13'd29: x = 8'h0c;
      13'd30: x = 8'ha9;
      13'd31: x = 8'h8d;
      13'd32: x = 8'ha0;
      13'd33: x = 8'h07;
      13'd34: x = 8'h20;
      13'd35: x = 8'hc9;
      13'd36: x = 8'he3;
      13'd37: x = 8'ha9;
      13'd38: x = 8'ha0;
      13'd39: x = 8'h88;
      13'd40: x = 8'hd0;
      13'd41: x = 8'hf8;
      13'd42: x = 8'ha0;
      13'd43: x = 8'h00;
      13'd44: x = 8'hb1;
      13'd45: x = 8'he2;
      13'd46: x = 8'he6;
      13'd47: x = 8'he2;
      13'd48: x = 8'hd0;
      13'd49: x = 8'h02;
      13'd50: x = 8'he6;
      13'd51: x = 8'he3;
      13'd52: x = 8'h60;
      13'd53: x = 8'h20;
      13'd54: x = 8'h15;
      13'd55: x = 8'he7;
      13'd56: x = 8'h20;
      13'd57: x = 8'h76;
      13'd58: x = 8'he5;
      13'd59: x = 8'ha5;
      13'd60: x = 8'he2;
      13'd61: x = 8'hc5;
      13'd62: x = 8'he6;
      13'd63: x = 8'ha5;
      13'd64: x = 8'he3;
      13'd65: x = 8'he5;
      13'd66: x = 8'he7;
      13'd67: x = 8'hb0;
      13'd68: x = 8'hef;
      13'd69: x = 8'h20;
      13'd70: x = 8'h6d;
      13'd71: x = 8'he0;
      13'd72: x = 8'h4c;
      13'd73: x = 8'h3b;
      13'd74: x = 8'he0;
      13'd75: x = 8'ha5;
      13'd76: x = 8'hca;
      13'd77: x = 8'h85;
      13'd78: x = 8'he2;
      13'd79: x = 8'ha5;
      13'd80: x = 8'hcb;
      13'd81: x = 8'h85;
      13'd82: x = 8'he3;
      13'd83: x = 8'ha5;
      13'd84: x = 8'h4c;
      13'd85: x = 8'h85;
      13'd86: x = 8'he6;
      13'd87: x = 8'ha5;
      13'd88: x = 8'h4d;
      13'd89: x = 8'h85;
      13'd90: x = 8'he7;
      13'd91: x = 8'hd0;
      13'd92: x = 8'hde;
      13'd93: x = 8'h20;
      13'd94: x = 8'h15;
      13'd95: x = 8'he7;
      13'd96: x = 8'h20;
      13'd97: x = 8'h6d;
      13'd98: x = 8'he5;
      13'd99: x = 8'ha5;
      13'd100: x = 8'he4;
      13'd101: x = 8'h85;
      13'd102: x = 8'he2;
      13'd103: x = 8'ha5;
      13'd104: x = 8'he5;
      13'd105: x = 8'h85;
      13'd106: x = 8'he3;
      13'd107: x = 8'hb0;
      13'd108: x = 8'hc7;
      13'd109: x = 8'h86;
      13'd110: x = 8'hd8;
      13'd111: x = 8'ha9;
      13'd112: x = 8'ha0;
      13'd113: x = 8'h85;
      13'd114: x = 8'hfa;
      13'd115: x = 8'h20;
      13'd116: x = 8'h2a;
      13'd117: x = 8'he0;
      13'd118: x = 8'h98;
      13'd119: x = 8'h85;
      13'd120: x = 8'he4;
      13'd121: x = 8'h20;
      13'd122: x = 8'h2a;
      13'd123: x = 8'he0;
      13'd124: x = 8'haa;
      13'd125: x = 8'h20;
      13'd126: x = 8'h2a;
      13'd127: x = 8'he0;
      13'd128: x = 8'h20;
      13'd129: x = 8'h1b;
      13'd130: x = 8'he5;
      13'd131: x = 8'h20;
      13'd132: x = 8'h18;
      13'd133: x = 8'he0;
      13'd134: x = 8'h84;
      13'd135: x = 8'hfa;
      13'd136: x = 8'haa;
      13'd137: x = 8'h10;
      13'd138: x = 8'h18;
      13'd139: x = 8'h0a;
      13'd140: x = 8'h10;
      13'd141: x = 8'he9;
      13'd142: x = 8'ha5;
      13'd143: x = 8'he4;
      13'd144: x = 8'hd0;
      13'd145: x = 8'h03;
      13'd146: x = 8'h20;
      13'd147: x = 8'h11;
      13'd148: x = 8'he0;
      13'd149: x = 8'h8a;
      13'd150: x = 8'h20;
      13'd151: x = 8'hc9;
      13'd152: x = 8'he3;
      13'd153: x = 8'ha9;
      13'd154: x = 8'h25;
      13'd155: x = 8'h20;
      13'd156: x = 8'h1a;
      13'd157: x = 8'he0;
      13'd158: x = 8'haa;
      13'd159: x = 8'h30;
      13'd160: x = 8'hf5;
      13'd161: x = 8'h85;
      13'd162: x = 8'he4;
      13'd163: x = 8'hc9;
      13'd164: x = 8'h01;
      13'd165: x = 8'hd0;
      13'd166: x = 8'h05;
      13'd167: x = 8'ha6;
      13'd168: x = 8'hd8;
      13'd169: x = 8'h4c;
      13'd170: x = 8'hcd;
      13'd171: x = 8'he3;
      13'd172: x = 8'h48;
      13'd173: x = 8'h84;
      13'd174: x = 8'hce;
      13'd175: x = 8'ha2;
      13'd176: x = 8'hed;
      13'd177: x = 8'h86;
      13'd178: x = 8'hcf;
      13'd179: x = 8'hc9;
      13'd180: x = 8'h51;
      13'd181: x = 8'h90;
      13'd182: x = 8'h04;
      13'd183: x = 8'hc6;
      13'd184: x = 8'hcf;
      13'd185: x = 8'he9;
      13'd186: x = 8'h50;
      13'd187: x = 8'h48;
      13'd188: x = 8'hb1;
      13'd189: x = 8'hce;
      13'd190: x = 8'haa;
      13'd191: x = 8'h88;
      13'd192: x = 8'hb1;
      13'd193: x = 8'hce;
      13'd194: x = 8'h10;
      13'd195: x = 8'hfa;
      13'd196: x = 8'he0;
      13'd197: x = 8'hc0;
      13'd198: x = 8'hb0;
      13'd199: x = 8'h04;
      13'd200: x = 8'he0;
      13'd201: x = 8'h00;
      13'd202: x = 8'h30;
      13'd203: x = 8'hf2;
      13'd204: x = 8'haa;
      13'd205: x = 8'h68;
      13'd206: x = 8'he9;
      13'd207: x = 8'h01;
      13'd208: x = 8'hd0;
      13'd209: x = 8'he9;
      13'd210: x = 8'h24;
      13'd211: x = 8'he4;
      13'd212: x = 8'h30;
      13'd213: x = 8'h03;
      13'd214: x = 8'h20;
      13'd215: x = 8'hf8;
      13'd216: x = 8'hef;
      13'd217: x = 8'hb1;
      13'd218: x = 8'hce;
      13'd219: x = 8'h10;
      13'd220: x = 8'h10;
      13'd221: x = 8'haa;
      13'd222: x = 8'h29;
      13'd223: x = 8'h3f;
      13'd224: x = 8'h85;
      13'd225: x = 8'he4;
      13'd226: x = 8'h18;
      13'd227: x = 8'h69;
      13'd228: x = 8'ha0;
      13'd229: x = 8'h20;
      13'd230: x = 8'hc9;
      13'd231: x = 8'he3;
      13'd232: x = 8'h88;
      13'd233: x = 8'he0;
      13'd234: x = 8'hc0;
      13'd235: x = 8'h90;
      13'd236: x = 8'hec;
      13'd237: x = 8'h20;
      13'd238: x = 8'h0c;
      13'd239: x = 8'he0;
      13'd240: x = 8'h68;
      13'd241: x = 8'hc9;
      13'd242: x = 8'h5d;
      13'd243: x = 8'hf0;
      13'd244: x = 8'ha4;
      13'd245: x = 8'hc9;
      13'd246: x = 8'h28;
      13'd247: x = 8'hd0;
      13'd248: x = 8'h8a;
      13'd249: x = 8'hf0;
      13'd250: x = 8'h9e;
      13'd251: x = 8'h20;
      13'd252: x = 8'h18;
      13'd253: x = 8'he1;
      13'd254: x = 8'h95;
      13'd255: x = 8'h50;
      13'd256: x = 8'hd5;
      13'd257: x = 8'h78;
      13'd258: x = 8'h90;
      13'd259: x = 8'h11;
      13'd260: x = 8'ha0;
      13'd261: x = 8'h2b;
      13'd262: x = 8'h4c;
      13'd263: x = 8'he0;
      13'd264: x = 8'he3;
      13'd265: x = 8'h20;
      13'd266: x = 8'h34;
      13'd267: x = 8'hee;
      13'd268: x = 8'hd5;
      13'd269: x = 8'h50;
      13'd270: x = 8'h90;
      13'd271: x = 8'hf4;
      13'd272: x = 8'h20;
      13'd273: x = 8'he4;
      13'd274: x = 8'hef;
      13'd275: x = 8'h95;
      13'd276: x = 8'h78;
      13'd277: x = 8'h4c;
      13'd278: x = 8'h23;
      13'd279: x = 8'he8;
      13'd280: x = 8'h20;
      13'd281: x = 8'h34;
      13'd282: x = 8'hee;
      13'd283: x = 8'hf0;
      13'd284: x = 8'he7;
      13'd285: x = 8'h38;
      13'd286: x = 8'he9;
      13'd287: x = 8'h01;
      13'd288: x = 8'h60;
      13'd289: x = 8'h20;
      13'd290: x = 8'h18;
      13'd291: x = 8'he1;
      13'd292: x = 8'h95;
      13'd293: x = 8'h50;
      13'd294: x = 8'h18;
      13'd295: x = 8'hf5;
      13'd296: x = 8'h78;
      13'd297: x = 8'h4c;
      13'd298: x = 8'h02;
      13'd299: x = 8'he1;
      13'd300: x = 8'ha0;
      13'd301: x = 8'h14;
      13'd302: x = 8'hd0;
      13'd303: x = 8'hd6;
      13'd304: x = 8'h20;
      13'd305: x = 8'h18;
      13'd306: x = 8'he1;
      13'd307: x = 8'he8;
      13'd308: x = 8'hb5;
      13'd309: x = 8'h50;
      13'd310: x = 8'h85;
      13'd311: x = 8'hda;
      13'd312: x = 8'h65;
      13'd313: x = 8'hce;
      13'd314: x = 8'h48;
      13'd315: x = 8'ha8;
      13'd316: x = 8'hb5;
      13'd317: x = 8'h78;
      13'd318: x = 8'h85;
      13'd319: x = 8'hdb;
      13'd320: x = 8'h65;
      13'd321: x = 8'hcf;
      13'd322: x = 8'h48;
      13'd323: x = 8'hc4;
      13'd324: x = 8'hca;
      13'd325: x = 8'he5;
      13'd326: x = 8'hcb;
      13'd327: x = 8'hb0;
      13'd328: x = 8'he3;
      13'd329: x = 8'ha5;
      13'd330: x = 8'hda;
      13'd331: x = 8'h69;
      13'd332: x = 8'hfe;
      13'd333: x = 8'h85;
      13'd334: x = 8'hda;
      13'd335: x = 8'ha9;
      13'd336: x = 8'hff;
      13'd337: x = 8'ha8;
      13'd338: x = 8'h65;
      13'd339: x = 8'hdb;
      13'd340: x = 8'h85;
      13'd341: x = 8'hdb;
      13'd342: x = 8'hc8;
      13'd343: x = 8'hb1;
      13'd344: x = 8'hda;
      13'd345: x = 8'hd9;
      13'd346: x = 8'hcc;
      13'd347: x = 8'h00;
      13'd348: x = 8'hd0;
      13'd349: x = 8'h0f;
      13'd350: x = 8'h98;
      13'd351: x = 8'hf0;
      13'd352: x = 8'hf5;
      13'd353: x = 8'h68;
      13'd354: x = 8'h91;
      13'd355: x = 8'hda;
      13'd356: x = 8'h99;
      13'd357: x = 8'hcc;
      13'd358: x = 8'h00;
      13'd359: x = 8'h88;
      13'd360: x = 8'h10;
      13'd361: x = 8'hf7;
      13'd362: x = 8'he8;
      13'd363: x = 8'h60;
      13'd364: x = 8'hea;
      13'd365: x = 8'ha0;
      13'd366: x = 8'h80;
      13'd367: x = 8'hd0;
      13'd368: x = 8'h95;
      13'd369: x = 8'ha9;
      13'd370: x = 8'h00;
      13'd371: x = 8'h20;
      13'd372: x = 8'h0a;
      13'd373: x = 8'he7;
      13'd374: x = 8'ha0;
      13'd375: x = 8'h02;
      13'd376: x = 8'h94;
      13'd377: x = 8'h78;
      13'd378: x = 8'h20;
      13'd379: x = 8'h0a;
      13'd380: x = 8'he7;
      13'd381: x = 8'ha9;
      13'd382: x = 8'hbf;
      13'd383: x = 8'h20;
      13'd384: x = 8'hc9;
      13'd385: x = 8'he3;
      13'd386: x = 8'ha0;
      13'd387: x = 8'h00;
      13'd388: x = 8'h20;
      13'd389: x = 8'h9e;
      13'd390: x = 8'he2;
      13'd391: x = 8'h94;
      13'd392: x = 8'h78;
      13'd393: x = 8'hea;
      13'd394: x = 8'hea;
      13'd395: x = 8'hea;
      13'd396: x = 8'hb5;
      13'd397: x = 8'h51;
      13'd398: x = 8'h85;
      13'd399: x = 8'hce;
      13'd400: x = 8'hb5;
      13'd401: x = 8'h79;
      13'd402: x = 8'h85;
      13'd403: x = 8'hcf;
      13'd404: x = 8'he8;
      13'd405: x = 8'he8;
      13'd406: x = 8'h20;
      13'd407: x = 8'hbc;
      13'd408: x = 8'he1;
      13'd409: x = 8'hb5;
      13'd410: x = 8'h4e;
      13'd411: x = 8'hd5;
      13'd412: x = 8'h76;
      13'd413: x = 8'hb0;
      13'd414: x = 8'h15;
      13'd415: x = 8'hf6;
      13'd416: x = 8'h4e;
      13'd417: x = 8'ha8;
      13'd418: x = 8'hb1;
      13'd419: x = 8'hce;
      13'd420: x = 8'hb4;
      13'd421: x = 8'h50;
      13'd422: x = 8'hc4;
      13'd423: x = 8'he4;
      13'd424: x = 8'h90;
      13'd425: x = 8'h04;
      13'd426: x = 8'ha0;
      13'd427: x = 8'h83;
      13'd428: x = 8'hd0;
      13'd429: x = 8'hc1;
      13'd430: x = 8'h91;
      13'd431: x = 8'hda;
      13'd432: x = 8'hf6;
      13'd433: x = 8'h50;
      13'd434: x = 8'h90;
      13'd435: x = 8'he5;
      13'd436: x = 8'hb4;
      13'd437: x = 8'h50;
      13'd438: x = 8'h8a;
      13'd439: x = 8'h91;
      13'd440: x = 8'hda;
      13'd441: x = 8'he8;
      13'd442: x = 8'he8;
      13'd443: x = 8'h60;
      13'd444: x = 8'hb5;
      13'd445: x = 8'h51;
      13'd446: x = 8'h85;
      13'd447: x = 8'hda;
      13'd448: x = 8'h38;
      13'd449: x = 8'he9;
      13'd450: x = 8'h02;
      13'd451: x = 8'h85;
      13'd452: x = 8'he4;
      13'd453: x = 8'hb5;
      13'd454: x = 8'h79;
      13'd455: x = 8'h85;
      13'd456: x = 8'hdb;
      13'd457: x = 8'he9;
      13'd458: x = 8'h00;
      13'd459: x = 8'h85;
      13'd460: x = 8'he5;
      13'd461: x = 8'ha0;
      13'd462: x = 8'h00;
      13'd463: x = 8'hb1;
      13'd464: x = 8'he4;
      13'd465: x = 8'h18;
      13'd466: x = 8'he5;
      13'd467: x = 8'hda;
      13'd468: x = 8'h85;
      13'd469: x = 8'he4;
      13'd470: x = 8'h60;
      13'd471: x = 8'hb5;
      13'd472: x = 8'h53;
      13'd473: x = 8'h85;
      13'd474: x = 8'hce;
      13'd475: x = 8'hb5;
      13'd476: x = 8'h7b;
      13'd477: x = 8'h85;
      13'd478: x = 8'hcf;
      13'd479: x = 8'hb5;
      13'd480: x = 8'h51;
      13'd481: x = 8'h85;
      13'd482: x = 8'hda;
      13'd483: x = 8'hb5;
      13'd484: x = 8'h79;
      13'd485: x = 8'h85;
      13'd486: x = 8'hdb;
      13'd487: x = 8'he8;
      13'd488: x = 8'he8;
      13'd489: x = 8'he8;
      13'd490: x = 8'ha0;
      13'd491: x = 8'h00;
      13'd492: x = 8'h94;
      13'd493: x = 8'h78;
      13'd494: x = 8'h94;
      13'd495: x = 8'ha0;
      13'd496: x = 8'hc8;
      13'd497: x = 8'h94;
      13'd498: x = 8'h50;
      13'd499: x = 8'hb5;
      13'd500: x = 8'h4d;
      13'd501: x = 8'hd5;
      13'd502: x = 8'h75;
      13'd503: x = 8'h08;
      13'd504: x = 8'h48;
      13'd505: x = 8'hb5;
      13'd506: x = 8'h4f;
      13'd507: x = 8'hd5;
      13'd508: x = 8'h77;
      13'd509: x = 8'h90;
      13'd510: x = 8'h07;
      13'd511: x = 8'h68;
      13'd512: x = 8'h28;
      13'd513: x = 8'hb0;
      13'd514: x = 8'h02;
      13'd515: x = 8'h56;
      13'd516: x = 8'h50;
      13'd517: x = 8'h60;
      13'd518: x = 8'ha8;
      13'd519: x = 8'hb1;
      13'd520: x = 8'hce;
      13'd521: x = 8'h85;
      13'd522: x = 8'he4;
      13'd523: x = 8'h68;
      13'd524: x = 8'ha8;
      13'd525: x = 8'h28;
      13'd526: x = 8'hb0;
      13'd527: x = 8'hf3;
      13'd528: x = 8'hb1;
      13'd529: x = 8'hda;
      13'd530: x = 8'hc5;
      13'd531: x = 8'he4;
      13'd532: x = 8'hd0;
      13'd533: x = 8'hed;
      13'd534: x = 8'hf6;
      13'd535: x = 8'h4f;
      13'd536: x = 8'hf6;
      13'd537: x = 8'h4d;
      13'd538: x = 8'hb0;
      13'd539: x = 8'hd7;
      13'd540: x = 8'h20;
      13'd541: x = 8'hd7;
      13'd542: x = 8'he1;
      13'd543: x = 8'h4c;
      13'd544: x = 8'h36;
      13'd545: x = 8'he7;
      13'd546: x = 8'h20;
      13'd547: x = 8'h54;
      13'd548: x = 8'he2;
      13'd549: x = 8'h06;
      13'd550: x = 8'hce;
      13'd551: x = 8'h26;
      13'd552: x = 8'hcf;
      13'd553: x = 8'h90;
      13'd554: x = 8'h0d;
      13'd555: x = 8'h18;
      13'd556: x = 8'ha5;
      13'd557: x = 8'he6;
      13'd558: x = 8'h65;
      13'd559: x = 8'hda;
      13'd560: x = 8'h85;
      13'd561: x = 8'he6;
      13'd562: x = 8'ha5;
      13'd563: x = 8'he7;
      13'd564: x = 8'h65;
      13'd565: x = 8'hdb;
      13'd566: x = 8'h85;
      13'd567: x = 8'he7;
      13'd568: x = 8'h88;
      13'd569: x = 8'hf0;
      13'd570: x = 8'h09;
      13'd571: x = 8'h06;
      13'd572: x = 8'he6;
      13'd573: x = 8'h26;
      13'd574: x = 8'he7;
      13'd575: x = 8'h10;
      13'd576: x = 8'he4;
      13'd577: x = 8'h4c;
      13'd578: x = 8'h7e;
      13'd579: x = 8'he7;
      13'd580: x = 8'ha5;
      13'd581: x = 8'he6;
      13'd582: x = 8'h20;
      13'd583: x = 8'h08;
      13'd584: x = 8'he7;
      13'd585: x = 8'ha5;
      13'd586: x = 8'he7;
      13'd587: x = 8'h95;
      13'd588: x = 8'ha0;
      13'd589: x = 8'h06;
      13'd590: x = 8'he5;
      13'd591: x = 8'h90;
      13'd592: x = 8'h28;
      13'd593: x = 8'h4c;
      13'd594: x = 8'h6f;
      13'd595: x = 8'he7;
      13'd596: x = 8'ha9;
      13'd597: x = 8'h55;
      13'd598: x = 8'h85;
      13'd599: x = 8'he5;
      13'd600: x = 8'h20;
      13'd601: x = 8'h5b;
      13'd602: x = 8'he2;
      13'd603: x = 8'ha5;
      13'd604: x = 8'hce;
      13'd605: x = 8'h85;
      13'd606: x = 8'hda;
      13'd607: x = 8'ha5;
      13'd608: x = 8'hcf;
      13'd609: x = 8'h85;
      13'd610: x = 8'hdb;
      13'd611: x = 8'h20;
      13'd612: x = 8'h15;
      13'd613: x = 8'he7;
      13'd614: x = 8'h84;
      13'd615: x = 8'he6;
      13'd616: x = 8'h84;
      13'd617: x = 8'he7;
      13'd618: x = 8'ha5;
      13'd619: x = 8'hcf;
      13'd620: x = 8'h10;
      13'd621: x = 8'h09;
      13'd622: x = 8'hca;
      13'd623: x = 8'h06;
      13'd624: x = 8'he5;
      13'd625: x = 8'h20;
      13'd626: x = 8'h6f;
      13'd627: x = 8'he7;
      13'd628: x = 8'h20;
      13'd629: x = 8'h15;
      13'd630: x = 8'he7;
      13'd631: x = 8'ha0;
      13'd632: x = 8'h10;
      13'd633: x = 8'h60;
      13'd634: x = 8'h20;
      13'd635: x = 8'h6c;
      13'd636: x = 8'hee;
      13'd637: x = 8'hf0;
      13'd638: x = 8'hc5;
      13'd639: x = 8'hff;
      13'd640: x = 8'hc9;
      13'd641: x = 8'h84;
      13'd642: x = 8'hd0;
      13'd643: x = 8'h02;
      13'd644: x = 8'h46;
      13'd645: x = 8'hf8;
      13'd646: x = 8'hc9;
      13'd647: x = 8'hdf;
      13'd648: x = 8'hf0;
      13'd649: x = 8'h11;
      13'd650: x = 8'hc9;
      13'd651: x = 8'h9b;
      13'd652: x = 8'hf0;
      13'd653: x = 8'h06;
      13'd654: x = 8'h99;
      13'd655: x = 8'h00;
      13'd656: x = 8'h02;
      13'd657: x = 8'hc8;
      13'd658: x = 8'h10;
      13'd659: x = 8'h0a;
      13'd660: x = 8'ha0;
      13'd661: x = 8'h8b;
      13'd662: x = 8'h20;
      13'd663: x = 8'hc4;
      13'd664: x = 8'he3;
      13'd665: x = 8'ha0;
      13'd666: x = 8'h01;
      13'd667: x = 8'h88;
      13'd668: x = 8'h30;
      13'd669: x = 8'hf6;
      13'd670: x = 8'h20;
      13'd671: x = 8'h03;
      13'd672: x = 8'he0;
      13'd673: x = 8'hea;
      13'd674: x = 8'hea;
      13'd675: x = 8'h20;
      13'd676: x = 8'hc9;
      13'd677: x = 8'he3;
      13'd678: x = 8'hc9;
      13'd679: x = 8'h8d;
      13'd680: x = 8'hd0;
      13'd681: x = 8'hd6;
      13'd682: x = 8'ha9;
      13'd683: x = 8'hdf;
      13'd684: x = 8'h99;
      13'd685: x = 8'h00;
      13'd686: x = 8'h02;
      13'd687: x = 8'h60;
      13'd688: x = 8'h20;
      13'd689: x = 8'hd3;
      13'd690: x = 8'hef;
      13'd691: x = 8'h20;
      13'd692: x = 8'hcd;
      13'd693: x = 8'he3;
      13'd694: x = 8'h46;
      13'd695: x = 8'hd9;
      13'd696: x = 8'ha9;
      13'd697: x = 8'hbe;
      13'd698: x = 8'h20;
      13'd699: x = 8'hc9;
      13'd700: x = 8'he3;
      13'd701: x = 8'ha0;
      13'd702: x = 8'h00;
      13'd703: x = 8'h84;
      13'd704: x = 8'hfa;
      13'd705: x = 8'h24;
      13'd706: x = 8'hf8;
      13'd707: x = 8'h10;
      13'd708: x = 8'h0c;
      13'd709: x = 8'ha6;
      13'd710: x = 8'hf6;
      13'd711: x = 8'ha5;
      13'd712: x = 8'hf7;
      13'd713: x = 8'h20;
      13'd714: x = 8'h1b;
      13'd715: x = 8'he5;
      13'd716: x = 8'ha9;
      13'd717: x = 8'ha0;
      13'd718: x = 8'h20;
      13'd719: x = 8'hc9;
      13'd720: x = 8'he3;
      13'd721: x = 8'ha2;
      13'd722: x = 8'hff;
      13'd723: x = 8'h9a;
      13'd724: x = 8'h20;
      13'd725: x = 8'h9e;
      13'd726: x = 8'he2;
      13'd727: x = 8'h84;
      13'd728: x = 8'hf1;
      13'd729: x = 8'h8a;
      13'd730: x = 8'h85;
      13'd731: x = 8'hc8;
      13'd732: x = 8'ha2;
      13'd733: x = 8'h20;
      13'd734: x = 8'h20;
      13'd735: x = 8'h91;
      13'd736: x = 8'he4;
      13'd737: x = 8'ha5;
      13'd738: x = 8'hc8;
      13'd739: x = 8'h69;
      13'd740: x = 8'h00;
      13'd741: x = 8'h85;
      13'd742: x = 8'he0;
      13'd743: x = 8'ha9;
      13'd744: x = 8'h00;
      13'd745: x = 8'haa;
      13'd746: x = 8'h69;
      13'd747: x = 8'h02;
      13'd748: x = 8'h85;
      13'd749: x = 8'he1;
      13'd750: x = 8'ha1;
      13'd751: x = 8'he0;
      13'd752: x = 8'h29;
      13'd753: x = 8'hf0;
      13'd754: x = 8'hc9;
      13'd755: x = 8'hb0;
      13'd756: x = 8'hf0;
      13'd757: x = 8'h03;
      13'd758: x = 8'h4c;
      13'd759: x = 8'h83;
      13'd760: x = 8'he8;
      13'd761: x = 8'ha0;
      13'd762: x = 8'h02;
      13'd763: x = 8'hb1;
      13'd764: x = 8'he0;
      13'd765: x = 8'h99;
      13'd766: x = 8'hcd;
      13'd767: x = 8'h00;
      13'd768: x = 8'h88;
      13'd769: x = 8'hd0;
      13'd770: x = 8'hf8;
      13'd771: x = 8'h20;
      13'd772: x = 8'h8a;
      13'd773: x = 8'he3;
      13'd774: x = 8'ha5;
      13'd775: x = 8'hf1;
      13'd776: x = 8'he5;
      13'd777: x = 8'hc8;
      13'd778: x = 8'hc9;
      13'd779: x = 8'h04;
      13'd780: x = 8'hf0;
      13'd781: x = 8'ha8;
      13'd782: x = 8'h91;
      13'd783: x = 8'he0;
      13'd784: x = 8'ha5;
      13'd785: x = 8'hca;
      13'd786: x = 8'hf1;
      13'd787: x = 8'he0;
      13'd788: x = 8'h85;
      13'd789: x = 8'he4;
      13'd790: x = 8'ha5;
      13'd791: x = 8'hcb;
      13'd792: x = 8'he9;
      13'd793: x = 8'h00;
      13'd794: x = 8'h85;
      13'd795: x = 8'he5;
      13'd796: x = 8'ha5;
      13'd797: x = 8'he4;
      13'd798: x = 8'hc5;
      13'd799: x = 8'hcc;
      13'd800: x = 8'ha5;
      13'd801: x = 8'he5;
      13'd802: x = 8'he5;
      13'd803: x = 8'hcd;
      13'd804: x = 8'h90;
      13'd805: x = 8'h45;
      13'd806: x = 8'ha5;
      13'd807: x = 8'hca;
      13'd808: x = 8'hf1;
      13'd809: x = 8'he0;
      13'd810: x = 8'h85;
      13'd811: x = 8'he6;
      13'd812: x = 8'ha5;
      13'd813: x = 8'hcb;
      13'd814: x = 8'he9;
      13'd815: x = 8'h00;
      13'd816: x = 8'h85;
      13'd817: x = 8'he7;
      13'd818: x = 8'hb1;
      13'd819: x = 8'hca;
      13'd820: x = 8'h91;
      13'd821: x = 8'he6;
      13'd822: x = 8'he6;
      13'd823: x = 8'hca;
      13'd824: x = 8'hd0;
      13'd825: x = 8'h02;
      13'd826: x = 8'he6;
      13'd827: x = 8'hcb;
      13'd828: x = 8'ha5;
      13'd829: x = 8'he2;
      13'd830: x = 8'hc5;
      13'd831: x = 8'hca;
      13'd832: x = 8'ha5;
      13'd833: x = 8'he3;
      13'd834: x = 8'he5;
      13'd835: x = 8'hcb;
      13'd836: x = 8'hb0;
      13'd837: x = 8'he0;
      13'd838: x = 8'hb5;
      13'd839: x = 8'he4;
      13'd840: x = 8'h95;
      13'd841: x = 8'hca;
      13'd842: x = 8'hca;
      13'd843: x = 8'h10;
      13'd844: x = 8'hf9;
      13'd845: x = 8'hb1;
      13'd846: x = 8'he0;
      13'd847: x = 8'ha8;
      13'd848: x = 8'h88;
      13'd849: x = 8'hb1;
      13'd850: x = 8'he0;
      13'd851: x = 8'h91;
      13'd852: x = 8'he6;
      13'd853: x = 8'h98;
      13'd854: x = 8'hd0;
      13'd855: x = 8'hf8;
      13'd856: x = 8'h24;
      13'd857: x = 8'hf8;
      13'd858: x = 8'h10;
      13'd859: x = 8'h09;
      13'd860: x = 8'hb5;
      13'd861: x = 8'hf7;
      13'd862: x = 8'h75;
      13'd863: x = 8'hf5;
      13'd864: x = 8'h95;
      13'd865: x = 8'hf7;
      13'd866: x = 8'he8;
      13'd867: x = 8'hf0;
      13'd868: x = 8'hf7;
      13'd869: x = 8'h10;
      13'd870: x = 8'h7e;
      13'd871: x = 8'h00;
      13'd872: x = 8'h00;
      13'd873: x = 8'h00;
      13'd874: x = 8'h00;
      13'd875: x = 8'ha0;
      13'd876: x = 8'h14;
      13'd877: x = 8'hd0;
      13'd878: x = 8'h71;
      13'd879: x = 8'h20;
      13'd880: x = 8'h15;
      13'd881: x = 8'he7;
      13'd882: x = 8'ha5;
      13'd883: x = 8'he2;
      13'd884: x = 8'h85;
      13'd885: x = 8'he6;
      13'd886: x = 8'ha5;
      13'd887: x = 8'he3;
      13'd888: x = 8'h85;
      13'd889: x = 8'he7;
      13'd890: x = 8'h20;
      13'd891: x = 8'h75;
      13'd892: x = 8'he5;
      13'd893: x = 8'ha5;
      13'd894: x = 8'he2;
      13'd895: x = 8'h85;
      13'd896: x = 8'he4;
      13'd897: x = 8'ha5;
      13'd898: x = 8'he3;
      13'd899: x = 8'h85;
      13'd900: x = 8'he5;
      13'd901: x = 8'hd0;
      13'd902: x = 8'h0e;
      13'd903: x = 8'h20;
      13'd904: x = 8'h15;
      13'd905: x = 8'he7;
      13'd906: x = 8'h20;
      13'd907: x = 8'h6d;
      13'd908: x = 8'he5;
      13'd909: x = 8'ha5;
      13'd910: x = 8'he6;
      13'd911: x = 8'h85;
      13'd912: x = 8'he2;
      13'd913: x = 8'ha5;
      13'd914: x = 8'he7;
      13'd915: x = 8'h85;
      13'd916: x = 8'he3;
      13'd917: x = 8'ha0;
      13'd918: x = 8'h00;
      13'd919: x = 8'ha5;
      13'd920: x = 8'hca;
      13'd921: x = 8'hc5;
      13'd922: x = 8'he4;
      13'd923: x = 8'ha5;
      13'd924: x = 8'hcb;
      13'd925: x = 8'he5;
      13'd926: x = 8'he5;
      13'd927: x = 8'hb0;
      13'd928: x = 8'h16;
      13'd929: x = 8'ha5;
      13'd930: x = 8'he4;
      13'd931: x = 8'hd0;
      13'd932: x = 8'h02;
      13'd933: x = 8'hc6;
      13'd934: x = 8'he5;
      13'd935: x = 8'hc6;
      13'd936: x = 8'he4;
      13'd937: x = 8'ha5;
      13'd938: x = 8'he6;
      13'd939: x = 8'hd0;
      13'd940: x = 8'h02;
      13'd941: x = 8'hc6;
      13'd942: x = 8'he7;
      13'd943: x = 8'hc6;
      13'd944: x = 8'he6;
      13'd945: x = 8'hb1;
      13'd946: x = 8'he4;
      13'd947: x = 8'h91;
      13'd948: x = 8'he6;
      13'd949: x = 8'h90;
      13'd950: x = 8'he0;
      13'd951: x = 8'ha5;
      13'd952: x = 8'he6;
      13'd953: x = 8'h85;
      13'd954: x = 8'hca;
      13'd955: x = 8'ha5;
      13'd956: x = 8'he7;
      13'd957: x = 8'h85;
      13'd958: x = 8'hcb;
      13'd959: x = 8'h60;
      13'd960: x = 8'h20;
      13'd961: x = 8'hc9;
      13'd962: x = 8'he3;
      13'd963: x = 8'hc8;
      13'd964: x = 8'hb9;
      13'd965: x = 8'h00;
      13'd966: x = 8'heb;
      13'd967: x = 8'h30;
      13'd968: x = 8'hf7;
      13'd969: x = 8'hc9;
      13'd970: x = 8'h8d;
      13'd971: x = 8'hd0;
      13'd972: x = 8'h06;
      13'd973: x = 8'ha9;
      13'd974: x = 8'h00;
      13'd975: x = 8'h85;
      13'd976: x = 8'h24;
      13'd977: x = 8'ha9;
      13'd978: x = 8'h8d;
      13'd979: x = 8'he6;
      13'd980: x = 8'h24;
      13'd981: x = 8'h2c;
      13'd982: x = 8'h12;
      13'd983: x = 8'hd0;
      13'd984: x = 8'h30;
      13'd985: x = 8'hfb;
      13'd986: x = 8'h8d;
      13'd987: x = 8'h12;
      13'd988: x = 8'hd0;
      13'd989: x = 8'h60;
      13'd990: x = 8'ha0;
      13'd991: x = 8'h06;
      13'd992: x = 8'h20;
      13'd993: x = 8'hd3;
      13'd994: x = 8'hee;
      13'd995: x = 8'h24;
      13'd996: x = 8'hd9;
      13'd997: x = 8'h30;
      13'd998: x = 8'h03;
      13'd999: x = 8'h4c;
      13'd1000: x = 8'hb6;
      13'd1001: x = 8'he2;
      13'd1002: x = 8'h4c;
      13'd1003: x = 8'h9a;
      13'd1004: x = 8'heb;
      13'd1005: x = 8'h2a;
      13'd1006: x = 8'h69;
      13'd1007: x = 8'ha0;
      13'd1008: x = 8'hdd;
      13'd1009: x = 8'h00;
      13'd1010: x = 8'h02;
      13'd1011: x = 8'hd0;
      13'd1012: x = 8'h53;
      13'd1013: x = 8'hb1;
      13'd1014: x = 8'hfe;
      13'd1015: x = 8'h0a;
      13'd1016: x = 8'h30;
      13'd1017: x = 8'h06;
      13'd1018: x = 8'h88;
      13'd1019: x = 8'hb1;
      13'd1020: x = 8'hfe;
      13'd1021: x = 8'h30;
      13'd1022: x = 8'h29;
      13'd1023: x = 8'hc8;
      13'd1024: x = 8'h86;
      13'd1025: x = 8'hc8;
      13'd1026: x = 8'h98;
      13'd1027: x = 8'h48;
      13'd1028: x = 8'ha2;
      13'd1029: x = 8'h00;
      13'd1030: x = 8'ha1;
      13'd1031: x = 8'hfe;
      13'd1032: x = 8'haa;
      13'd1033: x = 8'h4a;
      13'd1034: x = 8'h49;
      13'd1035: x = 8'h48;
      13'd1036: x = 8'h11;
      13'd1037: x = 8'hfe;
      13'd1038: x = 8'hc9;
      13'd1039: x = 8'hc0;
      13'd1040: x = 8'h90;
      13'd1041: x = 8'h01;
      13'd1042: x = 8'he8;
      13'd1043: x = 8'hc8;
      13'd1044: x = 8'hd0;
      13'd1045: x = 8'hf3;
      13'd1046: x = 8'h68;
      13'd1047: x = 8'ha8;
      13'd1048: x = 8'h8a;
      13'd1049: x = 8'h4c;
      13'd1050: x = 8'hc0;
      13'd1051: x = 8'he4;
      13'd1052: x = 8'he6;
      13'd1053: x = 8'hf1;
      13'd1054: x = 8'ha6;
      13'd1055: x = 8'hf1;
      13'd1056: x = 8'hf0;
      13'd1057: x = 8'hbc;
      13'd1058: x = 8'h9d;
      13'd1059: x = 8'h00;
      13'd1060: x = 8'h02;
      13'd1061: x = 8'h60;
      13'd1062: x = 8'ha6;
      13'd1063: x = 8'hc8;
      13'd1064: x = 8'ha9;
      13'd1065: x = 8'ha0;
      13'd1066: x = 8'he8;
      13'd1067: x = 8'hdd;
      13'd1068: x = 8'h00;
      13'd1069: x = 8'h02;
      13'd1070: x = 8'hb0;
      13'd1071: x = 8'hfa;
      13'd1072: x = 8'hb1;
      13'd1073: x = 8'hfe;
      13'd1074: x = 8'h29;
      13'd1075: x = 8'h3f;
      13'd1076: x = 8'h4a;
      13'd1077: x = 8'hd0;
      13'd1078: x = 8'hb6;
      13'd1079: x = 8'hbd;
      13'd1080: x = 8'h00;
      13'd1081: x = 8'h02;
      13'd1082: x = 8'hb0;
      13'd1083: x = 8'h06;
      13'd1084: x = 8'h69;
      13'd1085: x = 8'h3f;
      13'd1086: x = 8'hc9;
      13'd1087: x = 8'h1a;
      13'd1088: x = 8'h90;
      13'd1089: x = 8'h6f;
      13'd1090: x = 8'h69;
      13'd1091: x = 8'h4f;
      13'd1092: x = 8'hc9;
      13'd1093: x = 8'h0a;
      13'd1094: x = 8'h90;
      13'd1095: x = 8'h69;
      13'd1096: x = 8'ha6;
      13'd1097: x = 8'hfd;
      13'd1098: x = 8'hc8;
      13'd1099: x = 8'hb1;
      13'd1100: x = 8'hfe;
      13'd1101: x = 8'h29;
      13'd1102: x = 8'he0;
      13'd1103: x = 8'hc9;
      13'd1104: x = 8'h20;
      13'd1105: x = 8'hf0;
      13'd1106: x = 8'h7a;
      13'd1107: x = 8'hb5;
      13'd1108: x = 8'ha8;
      13'd1109: x = 8'h85;
      13'd1110: x = 8'hc8;
      13'd1111: x = 8'hb5;
      13'd1112: x = 8'hd1;
      13'd1113: x = 8'h85;
      13'd1114: x = 8'hf1;
      13'd1115: x = 8'h88;
      13'd1116: x = 8'hb1;
      13'd1117: x = 8'hfe;
      13'd1118: x = 8'h0a;
      13'd1119: x = 8'h10;
      13'd1120: x = 8'hfa;
      13'd1121: x = 8'h88;
      13'd1122: x = 8'hb0;
      13'd1123: x = 8'h38;
      13'd1124: x = 8'h0a;
      13'd1125: x = 8'h30;
      13'd1126: x = 8'h35;
      13'd1127: x = 8'hb4;
      13'd1128: x = 8'h58;
      13'd1129: x = 8'h84;
      13'd1130: x = 8'hff;
      13'd1131: x = 8'hb4;
      13'd1132: x = 8'h80;
      13'd1133: x = 8'he8;
      13'd1134: x = 8'h10;
      13'd1135: x = 8'hda;
      13'd1136: x = 8'hf0;
      13'd1137: x = 8'hb3;
      13'd1138: x = 8'hc9;
      13'd1139: x = 8'h7e;
      13'd1140: x = 8'hb0;
      13'd1141: x = 8'h22;
      13'd1142: x = 8'hca;
      13'd1143: x = 8'h10;
      13'd1144: x = 8'h04;
      13'd1145: x = 8'ha0;
      13'd1146: x = 8'h06;
      13'd1147: x = 8'h10;
      13'd1148: x = 8'h29;
      13'd1149: x = 8'h94;
      13'd1150: x = 8'h80;
      13'd1151: x = 8'ha4;
      13'd1152: x = 8'hff;
      13'd1153: x = 8'h94;
      13'd1154: x = 8'h58;
      13'd1155: x = 8'ha4;
      13'd1156: x = 8'hc8;
      13'd1157: x = 8'h94;
      13'd1158: x = 8'ha8;
      13'd1159: x = 8'ha4;
      13'd1160: x = 8'hf1;
      13'd1161: x = 8'h94;
      13'd1162: x = 8'hd1;
      13'd1163: x = 8'h29;
      13'd1164: x = 8'h1f;
      13'd1165: x = 8'ha8;
      13'd1166: x = 8'hb9;
      13'd1167: x = 8'h20;
      13'd1168: x = 8'hec;
      13'd1169: x = 8'h0a;
      13'd1170: x = 8'ha8;
      13'd1171: x = 8'ha9;
      13'd1172: x = 8'h76;
      13'd1173: x = 8'h2a;
      13'd1174: x = 8'h85;
      13'd1175: x = 8'hff;
      13'd1176: x = 8'hd0;
      13'd1177: x = 8'h01;
      13'd1178: x = 8'hc8;
      13'd1179: x = 8'hc8;
      13'd1180: x = 8'h86;
      13'd1181: x = 8'hfd;
      13'd1182: x = 8'hb1;
      13'd1183: x = 8'hfe;
      13'd1184: x = 8'h30;
      13'd1185: x = 8'h84;
      13'd1186: x = 8'hd0;
      13'd1187: x = 8'h05;
      13'd1188: x = 8'ha0;
      13'd1189: x = 8'h0e;
      13'd1190: x = 8'h4c;
      13'd1191: x = 8'he0;
      13'd1192: x = 8'he3;
      13'd1193: x = 8'hc9;
      13'd1194: x = 8'h03;
      13'd1195: x = 8'hb0;
      13'd1196: x = 8'hc3;
      13'd1197: x = 8'h4a;
      13'd1198: x = 8'ha6;
      13'd1199: x = 8'hc8;
      13'd1200: x = 8'he8;
      13'd1201: x = 8'hbd;
      13'd1202: x = 8'h00;
      13'd1203: x = 8'h02;
      13'd1204: x = 8'h90;
      13'd1205: x = 8'h04;
      13'd1206: x = 8'hc9;
      13'd1207: x = 8'ha2;
      13'd1208: x = 8'hf0;
      13'd1209: x = 8'h0a;
      13'd1210: x = 8'hc9;
      13'd1211: x = 8'hdf;
      13'd1212: x = 8'hf0;
      13'd1213: x = 8'h06;
      13'd1214: x = 8'h86;
      13'd1215: x = 8'hc8;
      13'd1216: x = 8'h20;
      13'd1217: x = 8'h1c;
      13'd1218: x = 8'he4;
      13'd1219: x = 8'hc8;
      13'd1220: x = 8'h88;
      13'd1221: x = 8'ha6;
      13'd1222: x = 8'hfd;
      13'd1223: x = 8'hb1;
      13'd1224: x = 8'hfe;
      13'd1225: x = 8'h88;
      13'd1226: x = 8'h0a;
      13'd1227: x = 8'h10;
      13'd1228: x = 8'hcf;
      13'd1229: x = 8'hb4;
      13'd1230: x = 8'h58;
      13'd1231: x = 8'h84;
      13'd1232: x = 8'hff;
      13'd1233: x = 8'hb4;
      13'd1234: x = 8'h80;
      13'd1235: x = 8'he8;
      13'd1236: x = 8'hb1;
      13'd1237: x = 8'hfe;
      13'd1238: x = 8'h29;
      13'd1239: x = 8'h9f;
      13'd1240: x = 8'hd0;
      13'd1241: x = 8'hed;
      13'd1242: x = 8'h85;
      13'd1243: x = 8'hf2;
      13'd1244: x = 8'h85;
      13'd1245: x = 8'hf3;
      13'd1246: x = 8'h98;
      13'd1247: x = 8'h48;
      13'd1248: x = 8'h86;
      13'd1249: x = 8'hfd;
      13'd1250: x = 8'hb4;
      13'd1251: x = 8'hd0;
      13'd1252: x = 8'h84;
      13'd1253: x = 8'hc9;
      13'd1254: x = 8'h18;
      13'd1255: x = 8'ha9;
      13'd1256: x = 8'h0a;
      13'd1257: x = 8'h85;
      13'd1258: x = 8'hf9;
      13'd1259: x = 8'ha2;
      13'd1260: x = 8'h00;
      13'd1261: x = 8'hc8;
      13'd1262: x = 8'hb9;
      13'd1263: x = 8'h00;
      13'd1264: x = 8'h02;
      13'd1265: x = 8'h29;
      13'd1266: x = 8'h0f;
      13'd1267: x = 8'h65;
      13'd1268: x = 8'hf2;
      13'd1269: x = 8'h48;
      13'd1270: x = 8'h8a;
      13'd1271: x = 8'h65;
      13'd1272: x = 8'hf3;
      13'd1273: x = 8'h30;
      13'd1274: x = 8'h1c;
      13'd1275: x = 8'haa;
      13'd1276: x = 8'h68;
      13'd1277: x = 8'hc6;
      13'd1278: x = 8'hf9;
      13'd1279: x = 8'hd0;
      13'd1280: x = 8'hf2;
      13'd1281: x = 8'h85;
      13'd1282: x = 8'hf2;
      13'd1283: x = 8'h86;
      13'd1284: x = 8'hf3;
      13'd1285: x = 8'hc4;
      13'd1286: x = 8'hf1;
      13'd1287: x = 8'hd0;
      13'd1288: x = 8'hde;
      13'd1289: x = 8'ha4;
      13'd1290: x = 8'hc9;
      13'd1291: x = 8'hc8;
      13'd1292: x = 8'h84;
      13'd1293: x = 8'hf1;
      13'd1294: x = 8'h20;
      13'd1295: x = 8'h1c;
      13'd1296: x = 8'he4;
      13'd1297: x = 8'h68;
      13'd1298: x = 8'ha8;
      13'd1299: x = 8'ha5;
      13'd1300: x = 8'hf3;
      13'd1301: x = 8'hb0;
      13'd1302: x = 8'ha9;
      13'd1303: x = 8'ha0;
      13'd1304: x = 8'h00;
      13'd1305: x = 8'h10;
      13'd1306: x = 8'h8b;
      13'd1307: x = 8'h85;
      13'd1308: x = 8'hf3;
      13'd1309: x = 8'h86;
      13'd1310: x = 8'hf2;
      13'd1311: x = 8'ha2;
      13'd1312: x = 8'h04;
      13'd1313: x = 8'h86;
      13'd1314: x = 8'hc9;
      13'd1315: x = 8'ha9;
      13'd1316: x = 8'hb0;
      13'd1317: x = 8'h85;
      13'd1318: x = 8'hf9;
      13'd1319: x = 8'ha5;
      13'd1320: x = 8'hf2;
      13'd1321: x = 8'hdd;
      13'd1322: x = 8'h63;
      13'd1323: x = 8'he5;
      13'd1324: x = 8'ha5;
      13'd1325: x = 8'hf3;
      13'd1326: x = 8'hfd;
      13'd1327: x = 8'h68;
      13'd1328: x = 8'he5;
      13'd1329: x = 8'h90;
      13'd1330: x = 8'h0d;
      13'd1331: x = 8'h85;
      13'd1332: x = 8'hf3;
      13'd1333: x = 8'ha5;
      13'd1334: x = 8'hf2;
      13'd1335: x = 8'hfd;
      13'd1336: x = 8'h63;
      13'd1337: x = 8'he5;
      13'd1338: x = 8'h85;
      13'd1339: x = 8'hf2;
      13'd1340: x = 8'he6;
      13'd1341: x = 8'hf9;
      13'd1342: x = 8'hd0;
      13'd1343: x = 8'he7;
      13'd1344: x = 8'ha5;
      13'd1345: x = 8'hf9;
      13'd1346: x = 8'he8;
      13'd1347: x = 8'hca;
      13'd1348: x = 8'hf0;
      13'd1349: x = 8'h0e;
      13'd1350: x = 8'hc9;
      13'd1351: x = 8'hb0;
      13'd1352: x = 8'hf0;
      13'd1353: x = 8'h02;
      13'd1354: x = 8'h85;
      13'd1355: x = 8'hc9;
      13'd1356: x = 8'h24;
      13'd1357: x = 8'hc9;
      13'd1358: x = 8'h30;
      13'd1359: x = 8'h04;
      13'd1360: x = 8'ha5;
      13'd1361: x = 8'hfa;
      13'd1362: x = 8'hf0;
      13'd1363: x = 8'h0b;
      13'd1364: x = 8'h20;
      13'd1365: x = 8'hc9;
      13'd1366: x = 8'he3;
      13'd1367: x = 8'h24;
      13'd1368: x = 8'hf8;
      13'd1369: x = 8'h10;
      13'd1370: x = 8'h04;
      13'd1371: x = 8'h99;
      13'd1372: x = 8'h00;
      13'd1373: x = 8'h02;
      13'd1374: x = 8'hc8;
      13'd1375: x = 8'hca;
      13'd1376: x = 8'h10;
      13'd1377: x = 8'hc1;
      13'd1378: x = 8'h60;
      13'd1379: x = 8'h01;
      13'd1380: x = 8'h0a;
      13'd1381: x = 8'h64;
      13'd1382: x = 8'he8;
      13'd1383: x = 8'h10;
      13'd1384: x = 8'h00;
      13'd1385: x = 8'h00;
      13'd1386: x = 8'h00;
      13'd1387: x = 8'h03;
      13'd1388: x = 8'h27;
      13'd1389: x = 8'ha5;
      13'd1390: x = 8'hca;
      13'd1391: x = 8'h85;
      13'd1392: x = 8'he6;
      13'd1393: x = 8'ha5;
      13'd1394: x = 8'hcb;
      13'd1395: x = 8'h85;
      13'd1396: x = 8'he7;
      13'd1397: x = 8'he8;
      13'd1398: x = 8'ha5;
      13'd1399: x = 8'he7;
      13'd1400: x = 8'h85;
      13'd1401: x = 8'he5;
      13'd1402: x = 8'ha5;
      13'd1403: x = 8'he6;
      13'd1404: x = 8'h85;
      13'd1405: x = 8'he4;
      13'd1406: x = 8'hc5;
      13'd1407: x = 8'h4c;
      13'd1408: x = 8'ha5;
      13'd1409: x = 8'he5;
      13'd1410: x = 8'he5;
      13'd1411: x = 8'h4d;
      13'd1412: x = 8'hb0;
      13'd1413: x = 8'h26;
      13'd1414: x = 8'ha0;
      13'd1415: x = 8'h01;
      13'd1416: x = 8'hb1;
      13'd1417: x = 8'he4;
      13'd1418: x = 8'he5;
      13'd1419: x = 8'hce;
      13'd1420: x = 8'hc8;
      13'd1421: x = 8'hb1;
      13'd1422: x = 8'he4;
      13'd1423: x = 8'he5;
      13'd1424: x = 8'hcf;
      13'd1425: x = 8'hb0;
      13'd1426: x = 8'h19;
      13'd1427: x = 8'ha0;
      13'd1428: x = 8'h00;
      13'd1429: x = 8'ha5;
      13'd1430: x = 8'he6;
      13'd1431: x = 8'h71;
      13'd1432: x = 8'he4;
      13'd1433: x = 8'h85;
      13'd1434: x = 8'he6;
      13'd1435: x = 8'h90;
      13'd1436: x = 8'h03;
      13'd1437: x = 8'he6;
      13'd1438: x = 8'he7;
      13'd1439: x = 8'h18;
      13'd1440: x = 8'hc8;
      13'd1441: x = 8'ha5;
      13'd1442: x = 8'hce;
      13'd1443: x = 8'hf1;
      13'd1444: x = 8'he4;
      13'd1445: x = 8'hc8;
      13'd1446: x = 8'ha5;
      13'd1447: x = 8'hcf;
      13'd1448: x = 8'hf1;
      13'd1449: x = 8'he4;
      13'd1450: x = 8'hb0;
      13'd1451: x = 8'hca;
      13'd1452: x = 8'h60;
      13'd1453: x = 8'h46;
      13'd1454: x = 8'hf8;
      13'd1455: x = 8'ha5;
      13'd1456: x = 8'h4c;
      13'd1457: x = 8'h85;
      13'd1458: x = 8'hca;
      13'd1459: x = 8'ha5;
      13'd1460: x = 8'h4d;
      13'd1461: x = 8'h85;
      13'd1462: x = 8'hcb;
      13'd1463: x = 8'ha5;
      13'd1464: x = 8'h4a;
      13'd1465: x = 8'h85;
      13'd1466: x = 8'hcc;
      13'd1467: x = 8'ha5;
      13'd1468: x = 8'h4b;
      13'd1469: x = 8'h85;
      13'd1470: x = 8'hcd;
      13'd1471: x = 8'ha9;
      13'd1472: x = 8'h00;
      13'd1473: x = 8'h85;
      13'd1474: x = 8'hfb;
      13'd1475: x = 8'h85;
      13'd1476: x = 8'hfc;
      13'd1477: x = 8'h85;
      13'd1478: x = 8'hfe;
      13'd1479: x = 8'ha9;
      13'd1480: x = 8'h00;
      13'd1481: x = 8'h85;
      13'd1482: x = 8'h1d;
      13'd1483: x = 8'h60;
      13'd1484: x = 8'ha5;
      13'd1485: x = 8'hd0;
      13'd1486: x = 8'h69;
      13'd1487: x = 8'h05;
      13'd1488: x = 8'h85;
      13'd1489: x = 8'hd2;
      13'd1490: x = 8'ha5;
      13'd1491: x = 8'hd1;
      13'd1492: x = 8'h69;
      13'd1493: x = 8'h00;
      13'd1494: x = 8'h85;
      13'd1495: x = 8'hd3;
      13'd1496: x = 8'ha5;
      13'd1497: x = 8'hd2;
      13'd1498: x = 8'hc5;
      13'd1499: x = 8'hca;
      13'd1500: x = 8'ha5;
      13'd1501: x = 8'hd3;
      13'd1502: x = 8'he5;
      13'd1503: x = 8'hcb;
      13'd1504: x = 8'h90;
      13'd1505: x = 8'h03;
      13'd1506: x = 8'h4c;
      13'd1507: x = 8'h6b;
      13'd1508: x = 8'he3;
      13'd1509: x = 8'ha5;
      13'd1510: x = 8'hce;
      13'd1511: x = 8'h91;
      13'd1512: x = 8'hd0;
      13'd1513: x = 8'ha5;
      13'd1514: x = 8'hcf;
      13'd1515: x = 8'hc8;
      13'd1516: x = 8'h91;
      13'd1517: x = 8'hd0;
      13'd1518: x = 8'ha5;
      13'd1519: x = 8'hd2;
      13'd1520: x = 8'hc8;
      13'd1521: x = 8'h91;
      13'd1522: x = 8'hd0;
      13'd1523: x = 8'ha5;
      13'd1524: x = 8'hd3;
      13'd1525: x = 8'hc8;
      13'd1526: x = 8'h91;
      13'd1527: x = 8'hd0;
      13'd1528: x = 8'ha9;
      13'd1529: x = 8'h00;
      13'd1530: x = 8'hc8;
      13'd1531: x = 8'h91;
      13'd1532: x = 8'hd0;
      13'd1533: x = 8'hc8;
      13'd1534: x = 8'h91;
      13'd1535: x = 8'hd0;
      13'd1536: x = 8'ha5;
      13'd1537: x = 8'hd2;
      13'd1538: x = 8'h85;
      13'd1539: x = 8'hcc;
      13'd1540: x = 8'ha5;
      13'd1541: x = 8'hd3;
      13'd1542: x = 8'h85;
      13'd1543: x = 8'hcd;
      13'd1544: x = 8'ha5;
      13'd1545: x = 8'hd0;
      13'd1546: x = 8'h90;
      13'd1547: x = 8'h43;
      13'd1548: x = 8'h85;
      13'd1549: x = 8'hce;
      13'd1550: x = 8'h84;
      13'd1551: x = 8'hcf;
      13'd1552: x = 8'h20;
      13'd1553: x = 8'hff;
      13'd1554: x = 8'he6;
      13'd1555: x = 8'h30;
      13'd1556: x = 8'h0e;
      13'd1557: x = 8'hc9;
      13'd1558: x = 8'h40;
      13'd1559: x = 8'hf0;
      13'd1560: x = 8'h0a;
      13'd1561: x = 8'h4c;
      13'd1562: x = 8'h28;
      13'd1563: x = 8'he6;
      13'd1564: x = 8'h06;
      13'd1565: x = 8'hc9;
      13'd1566: x = 8'h49;
      13'd1567: x = 8'hd0;
      13'd1568: x = 8'h07;
      13'd1569: x = 8'ha9;
      13'd1570: x = 8'h49;
      13'd1571: x = 8'h85;
      13'd1572: x = 8'hcf;
      13'd1573: x = 8'h20;
      13'd1574: x = 8'hff;
      13'd1575: x = 8'he6;
      13'd1576: x = 8'ha5;
      13'd1577: x = 8'h4b;
      13'd1578: x = 8'h85;
      13'd1579: x = 8'hd1;
      13'd1580: x = 8'ha5;
      13'd1581: x = 8'h4a;
      13'd1582: x = 8'h85;
      13'd1583: x = 8'hd0;
      13'd1584: x = 8'hc5;
      13'd1585: x = 8'hcc;
      13'd1586: x = 8'ha5;
      13'd1587: x = 8'hd1;
      13'd1588: x = 8'he5;
      13'd1589: x = 8'hcd;
      13'd1590: x = 8'hb0;
      13'd1591: x = 8'h94;
      13'd1592: x = 8'hb1;
      13'd1593: x = 8'hd0;
      13'd1594: x = 8'hc8;
      13'd1595: x = 8'hc5;
      13'd1596: x = 8'hce;
      13'd1597: x = 8'hd0;
      13'd1598: x = 8'h06;
      13'd1599: x = 8'hb1;
      13'd1600: x = 8'hd0;
      13'd1601: x = 8'hc5;
      13'd1602: x = 8'hcf;
      13'd1603: x = 8'hf0;
      13'd1604: x = 8'h0e;
      13'd1605: x = 8'hc8;
      13'd1606: x = 8'hb1;
      13'd1607: x = 8'hd0;
      13'd1608: x = 8'h48;
      13'd1609: x = 8'hc8;
      13'd1610: x = 8'hb1;
      13'd1611: x = 8'hd0;
      13'd1612: x = 8'h85;
      13'd1613: x = 8'hd1;
      13'd1614: x = 8'h68;
      13'd1615: x = 8'ha0;
      13'd1616: x = 8'h00;
      13'd1617: x = 8'hf0;
      13'd1618: x = 8'hdb;
      13'd1619: x = 8'ha5;
      13'd1620: x = 8'hd0;
      13'd1621: x = 8'h69;
      13'd1622: x = 8'h03;
      13'd1623: x = 8'h20;
      13'd1624: x = 8'h0a;
      13'd1625: x = 8'he7;
      13'd1626: x = 8'ha5;
      13'd1627: x = 8'hd1;
      13'd1628: x = 8'h69;
      13'd1629: x = 8'h00;
      13'd1630: x = 8'h95;
      13'd1631: x = 8'h78;
      13'd1632: x = 8'ha5;
      13'd1633: x = 8'hcf;
      13'd1634: x = 8'hc9;
      13'd1635: x = 8'h40;
      13'd1636: x = 8'hd0;
      13'd1637: x = 8'h1c;
      13'd1638: x = 8'h88;
      13'd1639: x = 8'h98;
      13'd1640: x = 8'h20;
      13'd1641: x = 8'h0a;
      13'd1642: x = 8'he7;
      13'd1643: x = 8'h88;
      13'd1644: x = 8'h94;
      13'd1645: x = 8'h78;
      13'd1646: x = 8'ha0;
      13'd1647: x = 8'h03;
      13'd1648: x = 8'hf6;
      13'd1649: x = 8'h78;
      13'd1650: x = 8'hc8;
      13'd1651: x = 8'hb1;
      13'd1652: x = 8'hd0;
      13'd1653: x = 8'h30;
      13'd1654: x = 8'hf9;
      13'd1655: x = 8'h10;
      13'd1656: x = 8'h09;
      13'd1657: x = 8'ha9;
      13'd1658: x = 8'h00;
      13'd1659: x = 8'h85;
      13'd1660: x = 8'hd4;
      13'd1661: x = 8'h85;
      13'd1662: x = 8'hd5;
      13'd1663: x = 8'ha2;
      13'd1664: x = 8'h20;
      13'd1665: x = 8'h48;
      13'd1666: x = 8'ha0;
      13'd1667: x = 8'h00;
      13'd1668: x = 8'hb1;
      13'd1669: x = 8'he0;
      13'd1670: x = 8'h10;
      13'd1671: x = 8'h18;
      13'd1672: x = 8'h0a;
      13'd1673: x = 8'h30;
      13'd1674: x = 8'h81;
      13'd1675: x = 8'h20;
      13'd1676: x = 8'hff;
      13'd1677: x = 8'he6;
      13'd1678: x = 8'h20;
      13'd1679: x = 8'h08;
      13'd1680: x = 8'he7;
      13'd1681: x = 8'h20;
      13'd1682: x = 8'hff;
      13'd1683: x = 8'he6;
      13'd1684: x = 8'h95;
      13'd1685: x = 8'ha0;
      13'd1686: x = 8'h24;
      13'd1687: x = 8'hd4;
      13'd1688: x = 8'h10;
      13'd1689: x = 8'h01;
      13'd1690: x = 8'hca;
      13'd1691: x = 8'h20;
      13'd1692: x = 8'hff;
      13'd1693: x = 8'he6;
      13'd1694: x = 8'hb0;
      13'd1695: x = 8'he6;
      13'd1696: x = 8'hc9;
      13'd1697: x = 8'h28;
      13'd1698: x = 8'hd0;
      13'd1699: x = 8'h1f;
      13'd1700: x = 8'ha5;
      13'd1701: x = 8'he0;
      13'd1702: x = 8'h20;
      13'd1703: x = 8'h0a;
      13'd1704: x = 8'he7;
      13'd1705: x = 8'ha5;
      13'd1706: x = 8'he1;
      13'd1707: x = 8'h95;
      13'd1708: x = 8'h78;
      13'd1709: x = 8'h24;
      13'd1710: x = 8'hd4;
      13'd1711: x = 8'h30;
      13'd1712: x = 8'h0b;
      13'd1713: x = 8'ha9;
      13'd1714: x = 8'h01;
      13'd1715: x = 8'h20;
      13'd1716: x = 8'h0a;
      13'd1717: x = 8'he7;
      13'd1718: x = 8'ha9;
      13'd1719: x = 8'h00;
      13'd1720: x = 8'h95;
      13'd1721: x = 8'h78;
      13'd1722: x = 8'hf6;
      13'd1723: x = 8'h78;
      13'd1724: x = 8'h20;
      13'd1725: x = 8'hff;
      13'd1726: x = 8'he6;
      13'd1727: x = 8'h30;
      13'd1728: x = 8'hf9;
      13'd1729: x = 8'hb0;
      13'd1730: x = 8'hd3;
      13'd1731: x = 8'h24;
      13'd1732: x = 8'hd4;
      13'd1733: x = 8'h10;
      13'd1734: x = 8'h06;
      13'd1735: x = 8'hc9;
      13'd1736: x = 8'h04;
      13'd1737: x = 8'hb0;
      13'd1738: x = 8'hd0;
      13'd1739: x = 8'h46;
      13'd1740: x = 8'hd4;
      13'd1741: x = 8'ha8;
      13'd1742: x = 8'h85;
      13'd1743: x = 8'hd6;
      13'd1744: x = 8'hb9;
      13'd1745: x = 8'h98;
      13'd1746: x = 8'he9;
      13'd1747: x = 8'h29;
      13'd1748: x = 8'h55;
      13'd1749: x = 8'h0a;
      13'd1750: x = 8'h85;
      13'd1751: x = 8'hd7;
      13'd1752: x = 8'h68;
      13'd1753: x = 8'ha8;
      13'd1754: x = 8'hb9;
      13'd1755: x = 8'h98;
      13'd1756: x = 8'he9;
      13'd1757: x = 8'h29;
      13'd1758: x = 8'haa;
      13'd1759: x = 8'hc5;
      13'd1760: x = 8'hd7;
      13'd1761: x = 8'hb0;
      13'd1762: x = 8'h09;
      13'd1763: x = 8'h98;
      13'd1764: x = 8'h48;
      13'd1765: x = 8'h20;
      13'd1766: x = 8'hff;
      13'd1767: x = 8'he6;
      13'd1768: x = 8'ha5;
      13'd1769: x = 8'hd6;
      13'd1770: x = 8'h90;
      13'd1771: x = 8'h95;
      13'd1772: x = 8'hb9;
      13'd1773: x = 8'h10;
      13'd1774: x = 8'hea;
      13'd1775: x = 8'h85;
      13'd1776: x = 8'hce;
      13'd1777: x = 8'hb9;
      13'd1778: x = 8'h88;
      13'd1779: x = 8'hea;
      13'd1780: x = 8'h85;
      13'd1781: x = 8'hcf;
      13'd1782: x = 8'h20;
      13'd1783: x = 8'hfc;
      13'd1784: x = 8'he6;
      13'd1785: x = 8'h4c;
      13'd1786: x = 8'hd8;
      13'd1787: x = 8'he6;
      13'd1788: x = 8'h6c;
      13'd1789: x = 8'hce;
      13'd1790: x = 8'h00;
      13'd1791: x = 8'he6;
      13'd1792: x = 8'he0;
      13'd1793: x = 8'hd0;
      13'd1794: x = 8'h02;
      13'd1795: x = 8'he6;
      13'd1796: x = 8'he1;
      13'd1797: x = 8'hb1;
      13'd1798: x = 8'he0;
      13'd1799: x = 8'h60;
      13'd1800: x = 8'h94;
      13'd1801: x = 8'h77;
      13'd1802: x = 8'hca;
      13'd1803: x = 8'h30;
      13'd1804: x = 8'h03;
      13'd1805: x = 8'h95;
      13'd1806: x = 8'h50;
      13'd1807: x = 8'h60;
      13'd1808: x = 8'ha0;
      13'd1809: x = 8'h66;
      13'd1810: x = 8'h4c;
      13'd1811: x = 8'he0;
      13'd1812: x = 8'he3;
      13'd1813: x = 8'ha0;
      13'd1814: x = 8'h00;
      13'd1815: x = 8'hb5;
      13'd1816: x = 8'h50;
      13'd1817: x = 8'h85;
      13'd1818: x = 8'hce;
      13'd1819: x = 8'hb5;
      13'd1820: x = 8'ha0;
      13'd1821: x = 8'h85;
      13'd1822: x = 8'hcf;
      13'd1823: x = 8'hb5;
      13'd1824: x = 8'h78;
      13'd1825: x = 8'hf0;
      13'd1826: x = 8'h0e;
      13'd1827: x = 8'h85;
      13'd1828: x = 8'hcf;
      13'd1829: x = 8'hb1;
      13'd1830: x = 8'hce;
      13'd1831: x = 8'h48;
      13'd1832: x = 8'hc8;
      13'd1833: x = 8'hb1;
      13'd1834: x = 8'hce;
      13'd1835: x = 8'h85;
      13'd1836: x = 8'hcf;
      13'd1837: x = 8'h68;
      13'd1838: x = 8'h85;
      13'd1839: x = 8'hce;
      13'd1840: x = 8'h88;
      13'd1841: x = 8'he8;
      13'd1842: x = 8'h60;
      13'd1843: x = 8'h20;
      13'd1844: x = 8'h4a;
      13'd1845: x = 8'he7;
      13'd1846: x = 8'h20;
      13'd1847: x = 8'h15;
      13'd1848: x = 8'he7;
      13'd1849: x = 8'h98;
      13'd1850: x = 8'h20;
      13'd1851: x = 8'h08;
      13'd1852: x = 8'he7;
      13'd1853: x = 8'h95;
      13'd1854: x = 8'ha0;
      13'd1855: x = 8'hc5;
      13'd1856: x = 8'hce;
      13'd1857: x = 8'hd0;
      13'd1858: x = 8'h06;
      13'd1859: x = 8'hc5;
      13'd1860: x = 8'hcf;
      13'd1861: x = 8'hd0;
      13'd1862: x = 8'h02;
      13'd1863: x = 8'hf6;
      13'd1864: x = 8'h50;
      13'd1865: x = 8'h60;
      13'd1866: x = 8'h20;
      13'd1867: x = 8'h82;
      13'd1868: x = 8'he7;
      13'd1869: x = 8'h20;
      13'd1870: x = 8'h59;
      13'd1871: x = 8'he7;
      13'd1872: x = 8'h20;
      13'd1873: x = 8'h15;
      13'd1874: x = 8'he7;
      13'd1875: x = 8'h24;
      13'd1876: x = 8'hcf;
      13'd1877: x = 8'h30;
      13'd1878: x = 8'h1b;
      13'd1879: x = 8'hca;
      13'd1880: x = 8'h60;
      13'd1881: x = 8'h20;
      13'd1882: x = 8'h15;
      13'd1883: x = 8'he7;
      13'd1884: x = 8'ha5;
      13'd1885: x = 8'hcf;
      13'd1886: x = 8'hd0;
      13'd1887: x = 8'h04;
      13'd1888: x = 8'ha5;
      13'd1889: x = 8'hce;
      13'd1890: x = 8'hf0;
      13'd1891: x = 8'hf3;
      13'd1892: x = 8'ha9;
      13'd1893: x = 8'hff;
      13'd1894: x = 8'h20;
      13'd1895: x = 8'h08;
      13'd1896: x = 8'he7;
      13'd1897: x = 8'h95;
      13'd1898: x = 8'ha0;
      13'd1899: x = 8'h24;
      13'd1900: x = 8'hcf;
      13'd1901: x = 8'h30;
      13'd1902: x = 8'he9;
      13'd1903: x = 8'h20;
      13'd1904: x = 8'h15;
      13'd1905: x = 8'he7;
      13'd1906: x = 8'h98;
      13'd1907: x = 8'h38;
      13'd1908: x = 8'he5;
      13'd1909: x = 8'hce;
      13'd1910: x = 8'h20;
      13'd1911: x = 8'h08;
      13'd1912: x = 8'he7;
      13'd1913: x = 8'h98;
      13'd1914: x = 8'he5;
      13'd1915: x = 8'hcf;
      13'd1916: x = 8'h50;
      13'd1917: x = 8'h23;
      13'd1918: x = 8'ha0;
      13'd1919: x = 8'h00;
      13'd1920: x = 8'h10;
      13'd1921: x = 8'h90;
      13'd1922: x = 8'h20;
      13'd1923: x = 8'h6f;
      13'd1924: x = 8'he7;
      13'd1925: x = 8'h20;
      13'd1926: x = 8'h15;
      13'd1927: x = 8'he7;
      13'd1928: x = 8'ha5;
      13'd1929: x = 8'hce;
      13'd1930: x = 8'h85;
      13'd1931: x = 8'hda;
      13'd1932: x = 8'ha5;
      13'd1933: x = 8'hcf;
      13'd1934: x = 8'h85;
      13'd1935: x = 8'hdb;
      13'd1936: x = 8'h20;
      13'd1937: x = 8'h15;
      13'd1938: x = 8'he7;
      13'd1939: x = 8'h18;
      13'd1940: x = 8'ha5;
      13'd1941: x = 8'hce;
      13'd1942: x = 8'h65;
      13'd1943: x = 8'hda;
      13'd1944: x = 8'h20;
      13'd1945: x = 8'h08;
      13'd1946: x = 8'he7;
      13'd1947: x = 8'ha5;
      13'd1948: x = 8'hcf;
      13'd1949: x = 8'h65;
      13'd1950: x = 8'hdb;
      13'd1951: x = 8'h70;
      13'd1952: x = 8'hdd;
      13'd1953: x = 8'h95;
      13'd1954: x = 8'ha0;
      13'd1955: x = 8'h60;
      13'd1956: x = 8'h20;
      13'd1957: x = 8'h15;
      13'd1958: x = 8'he7;
      13'd1959: x = 8'ha4;
      13'd1960: x = 8'hce;
      13'd1961: x = 8'hf0;
      13'd1962: x = 8'h05;
      13'd1963: x = 8'h88;
      13'd1964: x = 8'ha5;
      13'd1965: x = 8'hcf;
      13'd1966: x = 8'hf0;
      13'd1967: x = 8'h0c;
      13'd1968: x = 8'h60;
      13'd1969: x = 8'ha5;
      13'd1970: x = 8'h24;
      13'd1971: x = 8'h09;
      13'd1972: x = 8'h07;
      13'd1973: x = 8'ha8;
      13'd1974: x = 8'hc8;
      13'd1975: x = 8'ha9;
      13'd1976: x = 8'ha0;
      13'd1977: x = 8'h20;
      13'd1978: x = 8'hc9;
      13'd1979: x = 8'he3;
      13'd1980: x = 8'hc4;
      13'd1981: x = 8'h24;
      13'd1982: x = 8'hb0;
      13'd1983: x = 8'hf7;
      13'd1984: x = 8'h60;
      13'd1985: x = 8'h20;
      13'd1986: x = 8'hb1;
      13'd1987: x = 8'he7;
      13'd1988: x = 8'h20;
      13'd1989: x = 8'h15;
      13'd1990: x = 8'he7;
      13'd1991: x = 8'ha5;
      13'd1992: x = 8'hcf;
      13'd1993: x = 8'h10;
      13'd1994: x = 8'h0a;
      13'd1995: x = 8'ha9;
      13'd1996: x = 8'had;
      13'd1997: x = 8'h20;
      13'd1998: x = 8'hc9;
      13'd1999: x = 8'he3;
      13'd2000: x = 8'h20;
      13'd2001: x = 8'h72;
      13'd2002: x = 8'he7;
      13'd2003: x = 8'h50;
      13'd2004: x = 8'hef;
      13'd2005: x = 8'h88;
      13'd2006: x = 8'h84;
      13'd2007: x = 8'hd5;
      13'd2008: x = 8'h86;
      13'd2009: x = 8'hcf;
      13'd2010: x = 8'ha6;
      13'd2011: x = 8'hce;
      13'd2012: x = 8'h20;
      13'd2013: x = 8'h1b;
      13'd2014: x = 8'he5;
      13'd2015: x = 8'ha6;
      13'd2016: x = 8'hcf;
      13'd2017: x = 8'h60;
      13'd2018: x = 8'h20;
      13'd2019: x = 8'h15;
      13'd2020: x = 8'he7;
      13'd2021: x = 8'ha5;
      13'd2022: x = 8'hce;
      13'd2023: x = 8'h85;
      13'd2024: x = 8'hf6;
      13'd2025: x = 8'ha5;
      13'd2026: x = 8'hcf;
      13'd2027: x = 8'h85;
      13'd2028: x = 8'hf7;
      13'd2029: x = 8'h88;
      13'd2030: x = 8'h84;
      13'd2031: x = 8'hf8;
      13'd2032: x = 8'hc8;
      13'd2033: x = 8'ha9;
      13'd2034: x = 8'h0a;
      13'd2035: x = 8'h85;
      13'd2036: x = 8'hf4;
      13'd2037: x = 8'h84;
      13'd2038: x = 8'hf5;
      13'd2039: x = 8'h60;
      13'd2040: x = 8'h20;
      13'd2041: x = 8'h15;
      13'd2042: x = 8'he7;
      13'd2043: x = 8'ha5;
      13'd2044: x = 8'hce;
      13'd2045: x = 8'ha4;
      13'd2046: x = 8'hcf;
      13'd2047: x = 8'h10;
      13'd2048: x = 8'hf2;
      13'd2049: x = 8'h20;
      13'd2050: x = 8'h15;
      13'd2051: x = 8'he7;
      13'd2052: x = 8'hb5;
      13'd2053: x = 8'h50;
      13'd2054: x = 8'h85;
      13'd2055: x = 8'hda;
      13'd2056: x = 8'hb5;
      13'd2057: x = 8'h78;
      13'd2058: x = 8'h85;
      13'd2059: x = 8'hdb;
      13'd2060: x = 8'ha5;
      13'd2061: x = 8'hce;
      13'd2062: x = 8'h91;
      13'd2063: x = 8'hda;
      13'd2064: x = 8'hc8;
      13'd2065: x = 8'ha5;
      13'd2066: x = 8'hcf;
      13'd2067: x = 8'h91;
      13'd2068: x = 8'hda;
      13'd2069: x = 8'he8;
      13'd2070: x = 8'h60;
      13'd2071: x = 8'h68;
      13'd2072: x = 8'h68;
      13'd2073: x = 8'h24;
      13'd2074: x = 8'hd5;
      13'd2075: x = 8'h10;
      13'd2076: x = 8'h05;
      13'd2077: x = 8'h20;
      13'd2078: x = 8'hcd;
      13'd2079: x = 8'he3;
      13'd2080: x = 8'h46;
      13'd2081: x = 8'hd5;
      13'd2082: x = 8'h60;
      13'd2083: x = 8'ha0;
      13'd2084: x = 8'hff;
      13'd2085: x = 8'h84;
      13'd2086: x = 8'hd7;
      13'd2087: x = 8'h60;
      13'd2088: x = 8'h20;
      13'd2089: x = 8'hcd;
      13'd2090: x = 8'hef;
      13'd2091: x = 8'hf0;
      13'd2092: x = 8'h07;
      13'd2093: x = 8'ha9;
      13'd2094: x = 8'h25;
      13'd2095: x = 8'h85;
      13'd2096: x = 8'hd6;
      13'd2097: x = 8'h88;
      13'd2098: x = 8'h84;
      13'd2099: x = 8'hd4;
      13'd2100: x = 8'he8;
      13'd2101: x = 8'h60;
      13'd2102: x = 8'ha5;
      13'd2103: x = 8'hca;
      13'd2104: x = 8'ha4;
      13'd2105: x = 8'hcb;
      13'd2106: x = 8'hd0;
      13'd2107: x = 8'h5a;
      13'd2108: x = 8'ha0;
      13'd2109: x = 8'h41;
      13'd2110: x = 8'ha5;
      13'd2111: x = 8'hfc;
      13'd2112: x = 8'hc9;
      13'd2113: x = 8'h08;
      13'd2114: x = 8'hb0;
      13'd2115: x = 8'h5e;
      13'd2116: x = 8'ha8;
      13'd2117: x = 8'he6;
      13'd2118: x = 8'hfc;
      13'd2119: x = 8'ha5;
      13'd2120: x = 8'he0;
      13'd2121: x = 8'h99;
      13'd2122: x = 8'h00;
      13'd2123: x = 8'h01;
      13'd2124: x = 8'ha5;
      13'd2125: x = 8'he1;
      13'd2126: x = 8'h99;
      13'd2127: x = 8'h08;
      13'd2128: x = 8'h01;
      13'd2129: x = 8'ha5;
      13'd2130: x = 8'hdc;
      13'd2131: x = 8'h99;
      13'd2132: x = 8'h10;
      13'd2133: x = 8'h01;
      13'd2134: x = 8'ha5;
      13'd2135: x = 8'hdd;
      13'd2136: x = 8'h99;
      13'd2137: x = 8'h18;
      13'd2138: x = 8'h01;
      13'd2139: x = 8'h20;
      13'd2140: x = 8'h15;
      13'd2141: x = 8'he7;
      13'd2142: x = 8'h20;
      13'd2143: x = 8'h6d;
      13'd2144: x = 8'he5;
      13'd2145: x = 8'h90;
      13'd2146: x = 8'h04;
      13'd2147: x = 8'ha0;
      13'd2148: x = 8'h37;
      13'd2149: x = 8'hd0;
      13'd2150: x = 8'h3b;
      13'd2151: x = 8'ha5;
      13'd2152: x = 8'he4;
      13'd2153: x = 8'ha4;
      13'd2154: x = 8'he5;
      13'd2155: x = 8'h85;
      13'd2156: x = 8'hdc;
      13'd2157: x = 8'h84;
      13'd2158: x = 8'hdd;
      13'd2159: x = 8'h2c;
      13'd2160: x = 8'h11;
      13'd2161: x = 8'hd0;
      13'd2162: x = 8'h30;
      13'd2163: x = 8'h4f;
      13'd2164: x = 8'h18;
      13'd2165: x = 8'h69;
      13'd2166: x = 8'h03;
      13'd2167: x = 8'h90;
      13'd2168: x = 8'h01;
      13'd2169: x = 8'hc8;
      13'd2170: x = 8'ha2;
      13'd2171: x = 8'hff;
      13'd2172: x = 8'h86;
      13'd2173: x = 8'hd9;
      13'd2174: x = 8'h9a;
      13'd2175: x = 8'h85;
      13'd2176: x = 8'he0;
      13'd2177: x = 8'h84;
      13'd2178: x = 8'he1;
      13'd2179: x = 8'h20;
      13'd2180: x = 8'h79;
      13'd2181: x = 8'he6;
      13'd2182: x = 8'h24;
      13'd2183: x = 8'hd9;
      13'd2184: x = 8'h10;
      13'd2185: x = 8'h49;
      13'd2186: x = 8'h18;
      13'd2187: x = 8'ha0;
      13'd2188: x = 8'h00;
      13'd2189: x = 8'ha5;
      13'd2190: x = 8'hdc;
      13'd2191: x = 8'h71;
      13'd2192: x = 8'hdc;
      13'd2193: x = 8'ha4;
      13'd2194: x = 8'hdd;
      13'd2195: x = 8'h90;
      13'd2196: x = 8'h01;
      13'd2197: x = 8'hc8;
      13'd2198: x = 8'hc5;
      13'd2199: x = 8'h4c;
      13'd2200: x = 8'hd0;
      13'd2201: x = 8'hd1;
      13'd2202: x = 8'hc4;
      13'd2203: x = 8'h4d;
      13'd2204: x = 8'hd0;
      13'd2205: x = 8'hcd;
      13'd2206: x = 8'ha0;
      13'd2207: x = 8'h34;
      13'd2208: x = 8'h46;
      13'd2209: x = 8'hd9;
      13'd2210: x = 8'h4c;
      13'd2211: x = 8'he0;
      13'd2212: x = 8'he3;
      13'd2213: x = 8'ha0;
      13'd2214: x = 8'h4a;
      13'd2215: x = 8'ha5;
      13'd2216: x = 8'hfc;
      13'd2217: x = 8'hf0;
      13'd2218: x = 8'hf7;
      13'd2219: x = 8'hc6;
      13'd2220: x = 8'hfc;
      13'd2221: x = 8'ha8;
      13'd2222: x = 8'hb9;
      13'd2223: x = 8'h0f;
      13'd2224: x = 8'h01;
      13'd2225: x = 8'h85;
      13'd2226: x = 8'hdc;
      13'd2227: x = 8'hb9;
      13'd2228: x = 8'h17;
      13'd2229: x = 8'h01;
      13'd2230: x = 8'h85;
      13'd2231: x = 8'hdd;
      13'd2232: x = 8'hbe;
      13'd2233: x = 8'hff;
      13'd2234: x = 8'h00;
      13'd2235: x = 8'hb9;
      13'd2236: x = 8'h07;
      13'd2237: x = 8'h01;
      13'd2238: x = 8'ha8;
      13'd2239: x = 8'h8a;
      13'd2240: x = 8'h4c;
      13'd2241: x = 8'h7a;
      13'd2242: x = 8'he8;
      13'd2243: x = 8'ha0;
      13'd2244: x = 8'h63;
      13'd2245: x = 8'h20;
      13'd2246: x = 8'hc4;
      13'd2247: x = 8'he3;
      13'd2248: x = 8'ha0;
      13'd2249: x = 8'h01;
      13'd2250: x = 8'hb1;
      13'd2251: x = 8'hdc;
      13'd2252: x = 8'haa;
      13'd2253: x = 8'hc8;
      13'd2254: x = 8'hb1;
      13'd2255: x = 8'hdc;
      13'd2256: x = 8'h20;
      13'd2257: x = 8'h1b;
      13'd2258: x = 8'he5;
      13'd2259: x = 8'h4c;
      13'd2260: x = 8'hb3;
      13'd2261: x = 8'he2;
      13'd2262: x = 8'hc6;
      13'd2263: x = 8'hfb;
      13'd2264: x = 8'ha0;
      13'd2265: x = 8'h5b;
      13'd2266: x = 8'ha5;
      13'd2267: x = 8'hfb;
      13'd2268: x = 8'hf0;
      13'd2269: x = 8'hc4;
      13'd2270: x = 8'ha8;
      13'd2271: x = 8'hb5;
      13'd2272: x = 8'h50;
      13'd2273: x = 8'hd9;
      13'd2274: x = 8'h1f;
      13'd2275: x = 8'h01;
      13'd2276: x = 8'hd0;
      13'd2277: x = 8'hf0;
      13'd2278: x = 8'hb5;
      13'd2279: x = 8'h78;
      13'd2280: x = 8'hd9;
      13'd2281: x = 8'h27;
      13'd2282: x = 8'h01;
      13'd2283: x = 8'hd0;
      13'd2284: x = 8'he9;
      13'd2285: x = 8'hb9;
      13'd2286: x = 8'h2f;
      13'd2287: x = 8'h01;
      13'd2288: x = 8'h85;
      13'd2289: x = 8'hda;
      13'd2290: x = 8'hb9;
      13'd2291: x = 8'h37;
      13'd2292: x = 8'h01;
      13'd2293: x = 8'h85;
      13'd2294: x = 8'hdb;
      13'd2295: x = 8'h20;
      13'd2296: x = 8'h15;
      13'd2297: x = 8'he7;
      13'd2298: x = 8'hca;
      13'd2299: x = 8'h20;
      13'd2300: x = 8'h93;
      13'd2301: x = 8'he7;
      13'd2302: x = 8'h20;
      13'd2303: x = 8'h01;
      13'd2304: x = 8'he8;
      13'd2305: x = 8'hca;
      13'd2306: x = 8'ha4;
      13'd2307: x = 8'hfb;
      13'd2308: x = 8'hb9;
      13'd2309: x = 8'h67;
      13'd2310: x = 8'h01;
      13'd2311: x = 8'h95;
      13'd2312: x = 8'h9f;
      13'd2313: x = 8'hb9;
      13'd2314: x = 8'h5f;
      13'd2315: x = 8'h01;
      13'd2316: x = 8'ha0;
      13'd2317: x = 8'h00;
      13'd2318: x = 8'h20;
      13'd2319: x = 8'h08;
      13'd2320: x = 8'he7;
      13'd2321: x = 8'h20;
      13'd2322: x = 8'h82;
      13'd2323: x = 8'he7;
      13'd2324: x = 8'h20;
      13'd2325: x = 8'h59;
      13'd2326: x = 8'he7;
      13'd2327: x = 8'h20;
      13'd2328: x = 8'h15;
      13'd2329: x = 8'he7;
      13'd2330: x = 8'ha4;
      13'd2331: x = 8'hfb;
      13'd2332: x = 8'ha5;
      13'd2333: x = 8'hce;
      13'd2334: x = 8'hf0;
      13'd2335: x = 8'h05;
      13'd2336: x = 8'h59;
      13'd2337: x = 8'h37;
      13'd2338: x = 8'h01;
      13'd2339: x = 8'h10;
      13'd2340: x = 8'h12;
      13'd2341: x = 8'hb9;
      13'd2342: x = 8'h3f;
      13'd2343: x = 8'h01;
      13'd2344: x = 8'h85;
      13'd2345: x = 8'hdc;
      13'd2346: x = 8'hb9;
      13'd2347: x = 8'h47;
      13'd2348: x = 8'h01;
      13'd2349: x = 8'h85;
      13'd2350: x = 8'hdd;
      13'd2351: x = 8'hbe;
      13'd2352: x = 8'h4f;
      13'd2353: x = 8'h01;
      13'd2354: x = 8'hb9;
      13'd2355: x = 8'h57;
      13'd2356: x = 8'h01;
      13'd2357: x = 8'hd0;
      13'd2358: x = 8'h87;
      13'd2359: x = 8'hc6;
      13'd2360: x = 8'hfb;
      13'd2361: x = 8'h60;
      13'd2362: x = 8'ha0;
      13'd2363: x = 8'h54;
      13'd2364: x = 8'ha5;
      13'd2365: x = 8'hfb;
      13'd2366: x = 8'hc9;
      13'd2367: x = 8'h08;
      13'd2368: x = 8'hf0;
      13'd2369: x = 8'h9a;
      13'd2370: x = 8'he6;
      13'd2371: x = 8'hfb;
      13'd2372: x = 8'ha8;
      13'd2373: x = 8'hb5;
      13'd2374: x = 8'h50;
      13'd2375: x = 8'h99;
      13'd2376: x = 8'h20;
      13'd2377: x = 8'h01;
      13'd2378: x = 8'hb5;
      13'd2379: x = 8'h78;
      13'd2380: x = 8'h99;
      13'd2381: x = 8'h28;
      13'd2382: x = 8'h01;
      13'd2383: x = 8'h60;
      13'd2384: x = 8'h20;
      13'd2385: x = 8'h15;
      13'd2386: x = 8'he7;
      13'd2387: x = 8'ha4;
      13'd2388: x = 8'hfb;
      13'd2389: x = 8'ha5;
      13'd2390: x = 8'hce;
      13'd2391: x = 8'h99;
      13'd2392: x = 8'h5f;
      13'd2393: x = 8'h01;
      13'd2394: x = 8'ha5;
      13'd2395: x = 8'hcf;
      13'd2396: x = 8'h99;
      13'd2397: x = 8'h67;
      13'd2398: x = 8'h01;
      13'd2399: x = 8'ha9;
      13'd2400: x = 8'h01;
      13'd2401: x = 8'h99;
      13'd2402: x = 8'h2f;
      13'd2403: x = 8'h01;
      13'd2404: x = 8'ha9;
      13'd2405: x = 8'h00;
      13'd2406: x = 8'h99;
      13'd2407: x = 8'h37;
      13'd2408: x = 8'h01;
      13'd2409: x = 8'ha5;
      13'd2410: x = 8'hdc;
      13'd2411: x = 8'h99;
      13'd2412: x = 8'h3f;
      13'd2413: x = 8'h01;
      13'd2414: x = 8'ha5;
      13'd2415: x = 8'hdd;
      13'd2416: x = 8'h99;
      13'd2417: x = 8'h47;
      13'd2418: x = 8'h01;
      13'd2419: x = 8'ha5;
      13'd2420: x = 8'he0;
      13'd2421: x = 8'h99;
      13'd2422: x = 8'h4f;
      13'd2423: x = 8'h01;
      13'd2424: x = 8'ha5;
      13'd2425: x = 8'he1;
      13'd2426: x = 8'h99;
      13'd2427: x = 8'h57;
      13'd2428: x = 8'h01;
      13'd2429: x = 8'h60;
      13'd2430: x = 8'h20;
      13'd2431: x = 8'h15;
      13'd2432: x = 8'he7;
      13'd2433: x = 8'ha4;
      13'd2434: x = 8'hfb;
      13'd2435: x = 8'ha5;
      13'd2436: x = 8'hce;
      13'd2437: x = 8'h99;
      13'd2438: x = 8'h2f;
      13'd2439: x = 8'h01;
      13'd2440: x = 8'ha5;
      13'd2441: x = 8'hcf;
      13'd2442: x = 8'h4c;
      13'd2443: x = 8'h66;
      13'd2444: x = 8'he9;
      13'd2445: x = 8'h00;
      13'd2446: x = 8'h00;
      13'd2447: x = 8'h00;
      13'd2448: x = 8'h00;
      13'd2449: x = 8'h00;
      13'd2450: x = 8'h00;
      13'd2451: x = 8'h00;
      13'd2452: x = 8'h00;
      13'd2453: x = 8'h00;
      13'd2454: x = 8'h00;
      13'd2455: x = 8'h00;
      13'd2456: x = 8'h00;
      13'd2457: x = 8'h00;
      13'd2458: x = 8'h00;
      13'd2459: x = 8'hab;
      13'd2460: x = 8'h03;
      13'd2461: x = 8'h03;
      13'd2462: x = 8'h03;
      13'd2463: x = 8'h03;
      13'd2464: x = 8'h03;
      13'd2465: x = 8'h03;
      13'd2466: x = 8'h03;
      13'd2467: x = 8'h03;
      13'd2468: x = 8'h03;
      13'd2469: x = 8'h03;
      13'd2470: x = 8'h03;
      13'd2471: x = 8'h03;
      13'd2472: x = 8'h03;
      13'd2473: x = 8'h03;
      13'd2474: x = 8'h3f;
      13'd2475: x = 8'h3f;
      13'd2476: x = 8'hc0;
      13'd2477: x = 8'hc0;
      13'd2478: x = 8'h3c;
      13'd2479: x = 8'h3c;
      13'd2480: x = 8'h3c;
      13'd2481: x = 8'h3c;
      13'd2482: x = 8'h3c;
      13'd2483: x = 8'h3c;
      13'd2484: x = 8'h3c;
      13'd2485: x = 8'h30;
      13'd2486: x = 8'h0f;
      13'd2487: x = 8'hc0;
      13'd2488: x = 8'hcc;
      13'd2489: x = 8'hff;
      13'd2490: x = 8'h55;
      13'd2491: x = 8'h00;
      13'd2492: x = 8'hab;
      13'd2493: x = 8'hab;
      13'd2494: x = 8'h03;
      13'd2495: x = 8'h03;
      13'd2496: x = 8'hff;
      13'd2497: x = 8'hff;
      13'd2498: x = 8'h55;
      13'd2499: x = 8'hff;
      13'd2500: x = 8'hff;
      13'd2501: x = 8'h55;
      13'd2502: x = 8'hcf;
      13'd2503: x = 8'hcf;
      13'd2504: x = 8'hcf;
      13'd2505: x = 8'hcf;
      13'd2506: x = 8'hcf;
      13'd2507: x = 8'hff;
      13'd2508: x = 8'h55;
      13'd2509: x = 8'hc3;
      13'd2510: x = 8'hc3;
      13'd2511: x = 8'hc3;
      13'd2512: x = 8'h55;
      13'd2513: x = 8'hf0;
      13'd2514: x = 8'hf0;
      13'd2515: x = 8'hcf;
      13'd2516: x = 8'h56;
      13'd2517: x = 8'h56;
      13'd2518: x = 8'h56;
      13'd2519: x = 8'h55;
      13'd2520: x = 8'hff;
      13'd2521: x = 8'hff;
      13'd2522: x = 8'h55;
      13'd2523: x = 8'h03;
      13'd2524: x = 8'h03;
      13'd2525: x = 8'h03;
      13'd2526: x = 8'h03;
      13'd2527: x = 8'h03;
      13'd2528: x = 8'h03;
      13'd2529: x = 8'h03;
      13'd2530: x = 8'hff;
      13'd2531: x = 8'hff;
      13'd2532: x = 8'hff;
      13'd2533: x = 8'h03;
      13'd2534: x = 8'h03;
      13'd2535: x = 8'h03;
      13'd2536: x = 8'h03;
      13'd2537: x = 8'h03;
      13'd2538: x = 8'h03;
      13'd2539: x = 8'h03;
      13'd2540: x = 8'h03;
      13'd2541: x = 8'h03;
      13'd2542: x = 8'h03;
      13'd2543: x = 8'h03;
      13'd2544: x = 8'h03;
      13'd2545: x = 8'h03;
      13'd2546: x = 8'h03;
      13'd2547: x = 8'h03;
      13'd2548: x = 8'h03;
      13'd2549: x = 8'h00;
      13'd2550: x = 8'hab;
      13'd2551: x = 8'h03;
      13'd2552: x = 8'h57;
      13'd2553: x = 8'h03;
      13'd2554: x = 8'h03;
      13'd2555: x = 8'h03;
      13'd2556: x = 8'h03;
      13'd2557: x = 8'h07;
      13'd2558: x = 8'h03;
      13'd2559: x = 8'h03;
      13'd2560: x = 8'h03;
      13'd2561: x = 8'h03;
      13'd2562: x = 8'h03;
      13'd2563: x = 8'h03;
      13'd2564: x = 8'h03;
      13'd2565: x = 8'h03;
      13'd2566: x = 8'h03;
      13'd2567: x = 8'h03;
      13'd2568: x = 8'h03;
      13'd2569: x = 8'h03;
      13'd2570: x = 8'haa;
      13'd2571: x = 8'hff;
      13'd2572: x = 8'hff;
      13'd2573: x = 8'hff;
      13'd2574: x = 8'hff;
      13'd2575: x = 8'hff;
      13'd2576: x = 8'h17;
      13'd2577: x = 8'hff;
      13'd2578: x = 8'hff;
      13'd2579: x = 8'h19;
      13'd2580: x = 8'h5d;
      13'd2581: x = 8'h35;
      13'd2582: x = 8'h4b;
      13'd2583: x = 8'hf2;
      13'd2584: x = 8'hec;
      13'd2585: x = 8'h87;
      13'd2586: x = 8'h6f;
      13'd2587: x = 8'had;
      13'd2588: x = 8'hb7;
      13'd2589: x = 8'he2;
      13'd2590: x = 8'hf8;
      13'd2591: x = 8'h54;
      13'd2592: x = 8'h80;
      13'd2593: x = 8'h96;
      13'd2594: x = 8'h85;
      13'd2595: x = 8'h82;
      13'd2596: x = 8'h22;
      13'd2597: x = 8'h10;
      13'd2598: x = 8'h33;
      13'd2599: x = 8'h4a;
      13'd2600: x = 8'h13;
      13'd2601: x = 8'h06;
      13'd2602: x = 8'h0b;
      13'd2603: x = 8'h4a;
      13'd2604: x = 8'h01;
      13'd2605: x = 8'h40;
      13'd2606: x = 8'h47;
      13'd2607: x = 8'h7a;
      13'd2608: x = 8'h00;
      13'd2609: x = 8'hff;
      13'd2610: x = 8'h23;
      13'd2611: x = 8'h09;
      13'd2612: x = 8'h5b;
      13'd2613: x = 8'h16;
      13'd2614: x = 8'hb6;
      13'd2615: x = 8'hcb;
      13'd2616: x = 8'hff;
      13'd2617: x = 8'hff;
      13'd2618: x = 8'hfb;
      13'd2619: x = 8'hff;
      13'd2620: x = 8'hff;
      13'd2621: x = 8'h24;
      13'd2622: x = 8'hf6;
      13'd2623: x = 8'h4e;
      13'd2624: x = 8'h59;
      13'd2625: x = 8'h50;
      13'd2626: x = 8'h00;
      13'd2627: x = 8'hff;
      13'd2628: x = 8'h23;
      13'd2629: x = 8'ha3;
      13'd2630: x = 8'h6f;
      13'd2631: x = 8'h36;
      13'd2632: x = 8'h23;
      13'd2633: x = 8'hd7;
      13'd2634: x = 8'h1c;
      13'd2635: x = 8'h22;
      13'd2636: x = 8'hc2;
      13'd2637: x = 8'hae;
      13'd2638: x = 8'hba;
      13'd2639: x = 8'h23;
      13'd2640: x = 8'hff;
      13'd2641: x = 8'hff;
      13'd2642: x = 8'h21;
      13'd2643: x = 8'h30;
      13'd2644: x = 8'h1e;
      13'd2645: x = 8'h03;
      13'd2646: x = 8'hc4;
      13'd2647: x = 8'h20;
      13'd2648: x = 8'h00;
      13'd2649: x = 8'hc1;
      13'd2650: x = 8'hff;
      13'd2651: x = 8'hff;
      13'd2652: x = 8'hff;
      13'd2653: x = 8'ha0;
      13'd2654: x = 8'h30;
      13'd2655: x = 8'h1e;
      13'd2656: x = 8'ha4;
      13'd2657: x = 8'hd3;
      13'd2658: x = 8'hb6;
      13'd2659: x = 8'hbc;
      13'd2660: x = 8'haa;
      13'd2661: x = 8'h3a;
      13'd2662: x = 8'h01;
      13'd2663: x = 8'h50;
      13'd2664: x = 8'h7e;
      13'd2665: x = 8'hd8;
      13'd2666: x = 8'hd8;
      13'd2667: x = 8'ha5;
      13'd2668: x = 8'h3c;
      13'd2669: x = 8'hff;
      13'd2670: x = 8'h16;
      13'd2671: x = 8'h5b;
      13'd2672: x = 8'h28;
      13'd2673: x = 8'h03;
      13'd2674: x = 8'hc4;
      13'd2675: x = 8'h1d;
      13'd2676: x = 8'h00;
      13'd2677: x = 8'h0c;
      13'd2678: x = 8'h4e;
      13'd2679: x = 8'h00;
      13'd2680: x = 8'h3e;
      13'd2681: x = 8'h00;
      13'd2682: x = 8'ha6;
      13'd2683: x = 8'hb0;
      13'd2684: x = 8'h00;
      13'd2685: x = 8'hbc;
      13'd2686: x = 8'hc6;
      13'd2687: x = 8'h57;
      13'd2688: x = 8'h8c;
      13'd2689: x = 8'h01;
      13'd2690: x = 8'h27;
      13'd2691: x = 8'hff;
      13'd2692: x = 8'hff;
      13'd2693: x = 8'hff;
      13'd2694: x = 8'hff;
      13'd2695: x = 8'hff;
      13'd2696: x = 8'he8;
      13'd2697: x = 8'hff;
      13'd2698: x = 8'hff;
      13'd2699: x = 8'he8;
      13'd2700: x = 8'he0;
      13'd2701: x = 8'he0;
      13'd2702: x = 8'he0;
      13'd2703: x = 8'hef;
      13'd2704: x = 8'hef;
      13'd2705: x = 8'he3;
      13'd2706: x = 8'he3;
      13'd2707: x = 8'he5;
      13'd2708: x = 8'he5;
      13'd2709: x = 8'he7;
      13'd2710: x = 8'he7;
      13'd2711: x = 8'hee;
      13'd2712: x = 8'hef;
      13'd2713: x = 8'hef;
      13'd2714: x = 8'he7;
      13'd2715: x = 8'he7;
      13'd2716: x = 8'he2;
      13'd2717: x = 8'hef;
      13'd2718: x = 8'he7;
      13'd2719: x = 8'he7;
      13'd2720: x = 8'hec;
      13'd2721: x = 8'hec;
      13'd2722: x = 8'hec;
      13'd2723: x = 8'he7;
      13'd2724: x = 8'hec;
      13'd2725: x = 8'hec;
      13'd2726: x = 8'hec;
      13'd2727: x = 8'he2;
      13'd2728: x = 8'h00;
      13'd2729: x = 8'hff;
      13'd2730: x = 8'he8;
      13'd2731: x = 8'he1;
      13'd2732: x = 8'he8;
      13'd2733: x = 8'he8;
      13'd2734: x = 8'hef;
      13'd2735: x = 8'heb;
      13'd2736: x = 8'hff;
      13'd2737: x = 8'hff;
      13'd2738: x = 8'he0;
      13'd2739: x = 8'hff;
      13'd2740: x = 8'hff;
      13'd2741: x = 8'hef;
      13'd2742: x = 8'hee;
      13'd2743: x = 8'hef;
      13'd2744: x = 8'he7;
      13'd2745: x = 8'he7;
      13'd2746: x = 8'h00;
      13'd2747: x = 8'hff;
      13'd2748: x = 8'he8;
      13'd2749: x = 8'he7;
      13'd2750: x = 8'he7;
      13'd2751: x = 8'he7;
      13'd2752: x = 8'he8;
      13'd2753: x = 8'he1;
      13'd2754: x = 8'he2;
      13'd2755: x = 8'hee;
      13'd2756: x = 8'hee;
      13'd2757: x = 8'hee;
      13'd2758: x = 8'hee;
      13'd2759: x = 8'he8;
      13'd2760: x = 8'hff;
      13'd2761: x = 8'hff;
      13'd2762: x = 8'he1;
      13'd2763: x = 8'he1;
      13'd2764: x = 8'hef;
      13'd2765: x = 8'hee;
      13'd2766: x = 8'he7;
      13'd2767: x = 8'he8;
      13'd2768: x = 8'hee;
      13'd2769: x = 8'he7;
      13'd2770: x = 8'hff;
      13'd2771: x = 8'hff;
      13'd2772: x = 8'hff;
      13'd2773: x = 8'hee;
      13'd2774: x = 8'he1;
      13'd2775: x = 8'hef;
      13'd2776: x = 8'he7;
      13'd2777: x = 8'he8;
      13'd2778: x = 8'hef;
      13'd2779: x = 8'hef;
      13'd2780: x = 8'heb;
      13'd2781: x = 8'he9;
      13'd2782: x = 8'he8;
      13'd2783: x = 8'he9;
      13'd2784: x = 8'he9;
      13'd2785: x = 8'he8;
      13'd2786: x = 8'he8;
      13'd2787: x = 8'he8;
      13'd2788: x = 8'he8;
      13'd2789: x = 8'hff;
      13'd2790: x = 8'he8;
      13'd2791: x = 8'he8;
      13'd2792: x = 8'he8;
      13'd2793: x = 8'hee;
      13'd2794: x = 8'he7;
      13'd2795: x = 8'he8;
      13'd2796: x = 8'hef;
      13'd2797: x = 8'hef;
      13'd2798: x = 8'hee;
      13'd2799: x = 8'hef;
      13'd2800: x = 8'hee;
      13'd2801: x = 8'hef;
      13'd2802: x = 8'hee;
      13'd2803: x = 8'hee;
      13'd2804: x = 8'hef;
      13'd2805: x = 8'hee;
      13'd2806: x = 8'hee;
      13'd2807: x = 8'hee;
      13'd2808: x = 8'he1;
      13'd2809: x = 8'he8;
      13'd2810: x = 8'he8;
      13'd2811: x = 8'hff;
      13'd2812: x = 8'hff;
      13'd2813: x = 8'hff;
      13'd2814: x = 8'hff;
      13'd2815: x = 8'hff;
      13'd2816: x = 8'hbe;
      13'd2817: x = 8'hb3;
      13'd2818: x = 8'hb2;
      13'd2819: x = 8'hb7;
      13'd2820: x = 8'hb6;
      13'd2821: x = 8'h37;
      13'd2822: x = 8'hd4;
      13'd2823: x = 8'hcf;
      13'd2824: x = 8'hcf;
      13'd2825: x = 8'ha0;
      13'd2826: x = 8'hcc;
      13'd2827: x = 8'hcf;
      13'd2828: x = 8'hce;
      13'd2829: x = 8'h47;
      13'd2830: x = 8'hd3;
      13'd2831: x = 8'hd9;
      13'd2832: x = 8'hce;
      13'd2833: x = 8'hd4;
      13'd2834: x = 8'hc1;
      13'd2835: x = 8'h58;
      13'd2836: x = 8'hcd;
      13'd2837: x = 8'hc5;
      13'd2838: x = 8'hcd;
      13'd2839: x = 8'ha0;
      13'd2840: x = 8'hc6;
      13'd2841: x = 8'hd5;
      13'd2842: x = 8'hcc;
      13'd2843: x = 8'h4c;
      13'd2844: x = 8'hd4;
      13'd2845: x = 8'hcf;
      13'd2846: x = 8'hcf;
      13'd2847: x = 8'ha0;
      13'd2848: x = 8'hcd;
      13'd2849: x = 8'hc1;
      13'd2850: x = 8'hce;
      13'd2851: x = 8'hd9;
      13'd2852: x = 8'ha0;
      13'd2853: x = 8'hd0;
      13'd2854: x = 8'hc1;
      13'd2855: x = 8'hd2;
      13'd2856: x = 8'hc5;
      13'd2857: x = 8'hce;
      13'd2858: x = 8'h53;
      13'd2859: x = 8'hd3;
      13'd2860: x = 8'hd4;
      13'd2861: x = 8'hd2;
      13'd2862: x = 8'hc9;
      13'd2863: x = 8'hce;
      13'd2864: x = 8'h47;
      13'd2865: x = 8'hce;
      13'd2866: x = 8'hcf;
      13'd2867: x = 8'ha0;
      13'd2868: x = 8'hc5;
      13'd2869: x = 8'hce;
      13'd2870: x = 8'h44;
      13'd2871: x = 8'hc2;
      13'd2872: x = 8'hc1;
      13'd2873: x = 8'hc4;
      13'd2874: x = 8'ha0;
      13'd2875: x = 8'hc2;
      13'd2876: x = 8'hd2;
      13'd2877: x = 8'hc1;
      13'd2878: x = 8'hce;
      13'd2879: x = 8'hc3;
      13'd2880: x = 8'h48;
      13'd2881: x = 8'hbe;
      13'd2882: x = 8'hb8;
      13'd2883: x = 8'ha0;
      13'd2884: x = 8'hc7;
      13'd2885: x = 8'hcf;
      13'd2886: x = 8'hd3;
      13'd2887: x = 8'hd5;
      13'd2888: x = 8'hc2;
      13'd2889: x = 8'h53;
      13'd2890: x = 8'hc2;
      13'd2891: x = 8'hc1;
      13'd2892: x = 8'hc4;
      13'd2893: x = 8'ha0;
      13'd2894: x = 8'hd2;
      13'd2895: x = 8'hc5;
      13'd2896: x = 8'hd4;
      13'd2897: x = 8'hd5;
      13'd2898: x = 8'hd2;
      13'd2899: x = 8'h4e;
      13'd2900: x = 8'hbe;
      13'd2901: x = 8'hb8;
      13'd2902: x = 8'ha0;
      13'd2903: x = 8'hc6;
      13'd2904: x = 8'hcf;
      13'd2905: x = 8'hd2;
      13'd2906: x = 8'h53;
      13'd2907: x = 8'hc2;
      13'd2908: x = 8'hc1;
      13'd2909: x = 8'hc4;
      13'd2910: x = 8'ha0;
      13'd2911: x = 8'hce;
      13'd2912: x = 8'hc5;
      13'd2913: x = 8'hd8;
      13'd2914: x = 8'h54;
      13'd2915: x = 8'hd3;
      13'd2916: x = 8'hd4;
      13'd2917: x = 8'hcf;
      13'd2918: x = 8'hd0;
      13'd2919: x = 8'hd0;
      13'd2920: x = 8'hc5;
      13'd2921: x = 8'hc4;
      13'd2922: x = 8'ha0;
      13'd2923: x = 8'hc1;
      13'd2924: x = 8'hd4;
      13'd2925: x = 8'h20;
      13'd2926: x = 8'haa;
      13'd2927: x = 8'haa;
      13'd2928: x = 8'haa;
      13'd2929: x = 8'h20;
      13'd2930: x = 8'ha0;
      13'd2931: x = 8'hc5;
      13'd2932: x = 8'hd2;
      13'd2933: x = 8'hd2;
      13'd2934: x = 8'h0d;
      13'd2935: x = 8'hbe;
      13'd2936: x = 8'hb2;
      13'd2937: x = 8'hb5;
      13'd2938: x = 8'h35;
      13'd2939: x = 8'hd2;
      13'd2940: x = 8'hc1;
      13'd2941: x = 8'hce;
      13'd2942: x = 8'hc7;
      13'd2943: x = 8'h45;
      13'd2944: x = 8'hc4;
      13'd2945: x = 8'hc9;
      13'd2946: x = 8'h4d;
      13'd2947: x = 8'hd3;
      13'd2948: x = 8'hd4;
      13'd2949: x = 8'hd2;
      13'd2950: x = 8'ha0;
      13'd2951: x = 8'hcf;
      13'd2952: x = 8'hd6;
      13'd2953: x = 8'hc6;
      13'd2954: x = 8'h4c;
      13'd2955: x = 8'hdc;
      13'd2956: x = 8'h0d;
      13'd2957: x = 8'hd2;
      13'd2958: x = 8'hc5;
      13'd2959: x = 8'hd4;
      13'd2960: x = 8'hd9;
      13'd2961: x = 8'hd0;
      13'd2962: x = 8'hc5;
      13'd2963: x = 8'ha0;
      13'd2964: x = 8'hcc;
      13'd2965: x = 8'hc9;
      13'd2966: x = 8'hce;
      13'd2967: x = 8'hc5;
      13'd2968: x = 8'h8d;
      13'd2969: x = 8'h3f;
      13'd2970: x = 8'h46;
      13'd2971: x = 8'hd9;
      13'd2972: x = 8'h90;
      13'd2973: x = 8'h03;
      13'd2974: x = 8'h4c;
      13'd2975: x = 8'hc3;
      13'd2976: x = 8'he8;
      13'd2977: x = 8'ha6;
      13'd2978: x = 8'hcf;
      13'd2979: x = 8'h9a;
      13'd2980: x = 8'ha6;
      13'd2981: x = 8'hce;
      13'd2982: x = 8'ha0;
      13'd2983: x = 8'h8d;
      13'd2984: x = 8'hd0;
      13'd2985: x = 8'h02;
      13'd2986: x = 8'ha0;
      13'd2987: x = 8'h99;
      13'd2988: x = 8'h20;
      13'd2989: x = 8'hc4;
      13'd2990: x = 8'he3;
      13'd2991: x = 8'h86;
      13'd2992: x = 8'hce;
      13'd2993: x = 8'hba;
      13'd2994: x = 8'h86;
      13'd2995: x = 8'hcf;
      13'd2996: x = 8'ha0;
      13'd2997: x = 8'hfe;
      13'd2998: x = 8'h84;
      13'd2999: x = 8'hd9;
      13'd3000: x = 8'hc8;
      13'd3001: x = 8'h84;
      13'd3002: x = 8'hc8;
      13'd3003: x = 8'h20;
      13'd3004: x = 8'h99;
      13'd3005: x = 8'he2;
      13'd3006: x = 8'h84;
      13'd3007: x = 8'hf1;
      13'd3008: x = 8'ha2;
      13'd3009: x = 8'h20;
      13'd3010: x = 8'ha9;
      13'd3011: x = 8'h30;
      13'd3012: x = 8'h20;
      13'd3013: x = 8'h91;
      13'd3014: x = 8'he4;
      13'd3015: x = 8'he6;
      13'd3016: x = 8'hd9;
      13'd3017: x = 8'ha6;
      13'd3018: x = 8'hce;
      13'd3019: x = 8'ha4;
      13'd3020: x = 8'hc8;
      13'd3021: x = 8'h0a;
      13'd3022: x = 8'h85;
      13'd3023: x = 8'hce;
      13'd3024: x = 8'hc8;
      13'd3025: x = 8'hb9;
      13'd3026: x = 8'h00;
      13'd3027: x = 8'h02;
      13'd3028: x = 8'hc9;
      13'd3029: x = 8'h74;
      13'd3030: x = 8'hf0;
      13'd3031: x = 8'hd2;
      13'd3032: x = 8'h49;
      13'd3033: x = 8'hb0;
      13'd3034: x = 8'hc9;
      13'd3035: x = 8'h0a;
      13'd3036: x = 8'hb0;
      13'd3037: x = 8'hf0;
      13'd3038: x = 8'hc8;
      13'd3039: x = 8'hc8;
      13'd3040: x = 8'h84;
      13'd3041: x = 8'hc8;
      13'd3042: x = 8'hb9;
      13'd3043: x = 8'h00;
      13'd3044: x = 8'h02;
      13'd3045: x = 8'h48;
      13'd3046: x = 8'hb9;
      13'd3047: x = 8'hff;
      13'd3048: x = 8'h01;
      13'd3049: x = 8'ha0;
      13'd3050: x = 8'h00;
      13'd3051: x = 8'h20;
      13'd3052: x = 8'h08;
      13'd3053: x = 8'he7;
      13'd3054: x = 8'h68;
      13'd3055: x = 8'h95;
      13'd3056: x = 8'ha0;
      13'd3057: x = 8'ha5;
      13'd3058: x = 8'hce;
      13'd3059: x = 8'hc9;
      13'd3060: x = 8'hc7;
      13'd3061: x = 8'hd0;
      13'd3062: x = 8'h03;
      13'd3063: x = 8'h20;
      13'd3064: x = 8'h6f;
      13'd3065: x = 8'he7;
      13'd3066: x = 8'h4c;
      13'd3067: x = 8'h01;
      13'd3068: x = 8'he8;
      13'd3069: x = 8'hff;
      13'd3070: x = 8'hff;
      13'd3071: x = 8'hff;
      13'd3072: x = 8'h50;
      13'd3073: x = 8'h20;
      13'd3074: x = 8'h13;
      13'd3075: x = 8'hec;
      13'd3076: x = 8'hd0;
      13'd3077: x = 8'h15;
      13'd3078: x = 8'h20;
      13'd3079: x = 8'h0b;
      13'd3080: x = 8'hec;
      13'd3081: x = 8'hd0;
      13'd3082: x = 8'h10;
      13'd3083: x = 8'h20;
      13'd3084: x = 8'h82;
      13'd3085: x = 8'he7;
      13'd3086: x = 8'h20;
      13'd3087: x = 8'h6f;
      13'd3088: x = 8'he7;
      13'd3089: x = 8'h50;
      13'd3090: x = 8'h03;
      13'd3091: x = 8'h20;
      13'd3092: x = 8'h82;
      13'd3093: x = 8'he7;
      13'd3094: x = 8'h20;
      13'd3095: x = 8'h59;
      13'd3096: x = 8'he7;
      13'd3097: x = 8'h56;
      13'd3098: x = 8'h50;
      13'd3099: x = 8'h4c;
      13'd3100: x = 8'h36;
      13'd3101: x = 8'he7;
      13'd3102: x = 8'hff;
      13'd3103: x = 8'hff;
      13'd3104: x = 8'hc1;
      13'd3105: x = 8'hff;
      13'd3106: x = 8'h7f;
      13'd3107: x = 8'hd1;
      13'd3108: x = 8'hcc;
      13'd3109: x = 8'hc7;
      13'd3110: x = 8'hcf;
      13'd3111: x = 8'hce;
      13'd3112: x = 8'hc5;
      13'd3113: x = 8'h9a;
      13'd3114: x = 8'h98;
      13'd3115: x = 8'h8b;
      13'd3116: x = 8'h96;
      13'd3117: x = 8'h95;
      13'd3118: x = 8'h93;
      13'd3119: x = 8'hbf;
      13'd3120: x = 8'hb2;
      13'd3121: x = 8'h32;
      13'd3122: x = 8'h2d;
      13'd3123: x = 8'h2b;
      13'd3124: x = 8'hbc;
      13'd3125: x = 8'hb0;
      13'd3126: x = 8'hac;
      13'd3127: x = 8'hbe;
      13'd3128: x = 8'h35;
      13'd3129: x = 8'h8e;
      13'd3130: x = 8'h61;
      13'd3131: x = 8'hff;
      13'd3132: x = 8'hff;
      13'd3133: x = 8'hff;
      13'd3134: x = 8'hdd;
      13'd3135: x = 8'hfb;
      13'd3136: x = 8'h20;
      13'd3137: x = 8'hc9;
      13'd3138: x = 8'hef;
      13'd3139: x = 8'h15;
      13'd3140: x = 8'h4f;
      13'd3141: x = 8'h10;
      13'd3142: x = 8'h05;
      13'd3143: x = 8'h20;
      13'd3144: x = 8'hc9;
      13'd3145: x = 8'hef;
      13'd3146: x = 8'h35;
      13'd3147: x = 8'h4f;
      13'd3148: x = 8'h95;
      13'd3149: x = 8'h50;
      13'd3150: x = 8'h10;
      13'd3151: x = 8'hcb;
      13'd3152: x = 8'h4c;
      13'd3153: x = 8'hc9;
      13'd3154: x = 8'hef;
      13'd3155: x = 8'h40;
      13'd3156: x = 8'h60;
      13'd3157: x = 8'h8d;
      13'd3158: x = 8'h60;
      13'd3159: x = 8'h8b;
      13'd3160: x = 8'h00;
      13'd3161: x = 8'h7e;
      13'd3162: x = 8'h8c;
      13'd3163: x = 8'h33;
      13'd3164: x = 8'h00;
      13'd3165: x = 8'h00;
      13'd3166: x = 8'h60;
      13'd3167: x = 8'h03;
      13'd3168: x = 8'hbf;
      13'd3169: x = 8'h12;
      13'd3170: x = 8'h00;
      13'd3171: x = 8'h40;
      13'd3172: x = 8'h89;
      13'd3173: x = 8'hc9;
      13'd3174: x = 8'h47;
      13'd3175: x = 8'h9d;
      13'd3176: x = 8'h17;
      13'd3177: x = 8'h68;
      13'd3178: x = 8'h9d;
      13'd3179: x = 8'h0a;
      13'd3180: x = 8'h00;
      13'd3181: x = 8'h40;
      13'd3182: x = 8'h60;
      13'd3183: x = 8'h8d;
      13'd3184: x = 8'h60;
      13'd3185: x = 8'h8b;
      13'd3186: x = 8'h00;
      13'd3187: x = 8'h7e;
      13'd3188: x = 8'h8c;
      13'd3189: x = 8'h3c;
      13'd3190: x = 8'h00;
      13'd3191: x = 8'h00;
      13'd3192: x = 8'h60;
      13'd3193: x = 8'h03;
      13'd3194: x = 8'hbf;
      13'd3195: x = 8'h1b;
      13'd3196: x = 8'h4b;
      13'd3197: x = 8'h67;
      13'd3198: x = 8'hb4;
      13'd3199: x = 8'ha1;
      13'd3200: x = 8'h07;
      13'd3201: x = 8'h8c;
      13'd3202: x = 8'h07;
      13'd3203: x = 8'hae;
      13'd3204: x = 8'ha9;
      13'd3205: x = 8'hac;
      13'd3206: x = 8'ha8;
      13'd3207: x = 8'h67;
      13'd3208: x = 8'h8c;
      13'd3209: x = 8'h07;
      13'd3210: x = 8'hb4;
      13'd3211: x = 8'haf;
      13'd3212: x = 8'hac;
      13'd3213: x = 8'hb0;
      13'd3214: x = 8'h67;
      13'd3215: x = 8'h9d;
      13'd3216: x = 8'hb2;
      13'd3217: x = 8'haf;
      13'd3218: x = 8'hac;
      13'd3219: x = 8'haf;
      13'd3220: x = 8'ha3;
      13'd3221: x = 8'h67;
      13'd3222: x = 8'h8c;
      13'd3223: x = 8'h07;
      13'd3224: x = 8'ha5;
      13'd3225: x = 8'hab;
      13'd3226: x = 8'haf;
      13'd3227: x = 8'hb0;
      13'd3228: x = 8'hf4;
      13'd3229: x = 8'hae;
      13'd3230: x = 8'ha9;
      13'd3231: x = 8'hb2;
      13'd3232: x = 8'hb0;
      13'd3233: x = 8'h7f;
      13'd3234: x = 8'h0e;
      13'd3235: x = 8'h27;
      13'd3236: x = 8'hb4;
      13'd3237: x = 8'hae;
      13'd3238: x = 8'ha9;
      13'd3239: x = 8'hb2;
      13'd3240: x = 8'hb0;
      13'd3241: x = 8'h7f;
      13'd3242: x = 8'h0e;
      13'd3243: x = 8'h28;
      13'd3244: x = 8'hb4;
      13'd3245: x = 8'hae;
      13'd3246: x = 8'ha9;
      13'd3247: x = 8'hb2;
      13'd3248: x = 8'hb0;
      13'd3249: x = 8'h64;
      13'd3250: x = 8'h07;
      13'd3251: x = 8'ha6;
      13'd3252: x = 8'ha9;
      13'd3253: x = 8'h67;
      13'd3254: x = 8'haf;
      13'd3255: x = 8'hb4;
      13'd3256: x = 8'haf;
      13'd3257: x = 8'ha7;
      13'd3258: x = 8'h78;
      13'd3259: x = 8'hb4;
      13'd3260: x = 8'ha5;
      13'd3261: x = 8'hac;
      13'd3262: x = 8'h78;
      13'd3263: x = 8'h7f;
      13'd3264: x = 8'h02;
      13'd3265: x = 8'had;
      13'd3266: x = 8'ha5;
      13'd3267: x = 8'hb2;
      13'd3268: x = 8'h67;
      13'd3269: x = 8'ha2;
      13'd3270: x = 8'hb5;
      13'd3271: x = 8'hb3;
      13'd3272: x = 8'haf;
      13'd3273: x = 8'ha7;
      13'd3274: x = 8'hee;
      13'd3275: x = 8'hb2;
      13'd3276: x = 8'hb5;
      13'd3277: x = 8'hb4;
      13'd3278: x = 8'ha5;
      13'd3279: x = 8'hb2;
      13'd3280: x = 8'h7e;
      13'd3281: x = 8'h8c;
      13'd3282: x = 8'h39;
      13'd3283: x = 8'hb4;
      13'd3284: x = 8'hb8;
      13'd3285: x = 8'ha5;
      13'd3286: x = 8'hae;
      13'd3287: x = 8'h67;
      13'd3288: x = 8'hb0;
      13'd3289: x = 8'ha5;
      13'd3290: x = 8'hb4;
      13'd3291: x = 8'hb3;
      13'd3292: x = 8'h27;
      13'd3293: x = 8'haf;
      13'd3294: x = 8'hb4;
      13'd3295: x = 8'h07;
      13'd3296: x = 8'h9d;
      13'd3297: x = 8'h19;
      13'd3298: x = 8'hb2;
      13'd3299: x = 8'haf;
      13'd3300: x = 8'ha6;
      13'd3301: x = 8'h7f;
      13'd3302: x = 8'h05;
      13'd3303: x = 8'h37;
      13'd3304: x = 8'hb4;
      13'd3305: x = 8'hb5;
      13'd3306: x = 8'hb0;
      13'd3307: x = 8'hae;
      13'd3308: x = 8'ha9;
      13'd3309: x = 8'h7f;
      13'd3310: x = 8'h05;
      13'd3311: x = 8'h28;
      13'd3312: x = 8'hb4;
      13'd3313: x = 8'hb5;
      13'd3314: x = 8'hb0;
      13'd3315: x = 8'hae;
      13'd3316: x = 8'ha9;
      13'd3317: x = 8'h7f;
      13'd3318: x = 8'h05;
      13'd3319: x = 8'h2a;
      13'd3320: x = 8'hb4;
      13'd3321: x = 8'hb5;
      13'd3322: x = 8'hb0;
      13'd3323: x = 8'hae;
      13'd3324: x = 8'ha9;
      13'd3325: x = 8'he4;
      13'd3326: x = 8'hae;
      13'd3327: x = 8'ha5;
      13'd3328: x = 8'h00;
      13'd3329: x = 8'hff;
      13'd3330: x = 8'hff;
      13'd3331: x = 8'h47;
      13'd3332: x = 8'ha2;
      13'd3333: x = 8'ha1;
      13'd3334: x = 8'hb4;
      13'd3335: x = 8'h7f;
      13'd3336: x = 8'h0d;
      13'd3337: x = 8'h30;
      13'd3338: x = 8'had;
      13'd3339: x = 8'ha9;
      13'd3340: x = 8'ha4;
      13'd3341: x = 8'h7f;
      13'd3342: x = 8'h0d;
      13'd3343: x = 8'h23;
      13'd3344: x = 8'had;
      13'd3345: x = 8'ha9;
      13'd3346: x = 8'ha4;
      13'd3347: x = 8'h67;
      13'd3348: x = 8'hac;
      13'd3349: x = 8'hac;
      13'd3350: x = 8'ha1;
      13'd3351: x = 8'ha3;
      13'd3352: x = 8'h00;
      13'd3353: x = 8'h40;
      13'd3354: x = 8'h80;
      13'd3355: x = 8'hc0;
      13'd3356: x = 8'hc1;
      13'd3357: x = 8'h80;
      13'd3358: x = 8'h00;
      13'd3359: x = 8'h47;
      13'd3360: x = 8'h8c;
      13'd3361: x = 8'h68;
      13'd3362: x = 8'h8c;
      13'd3363: x = 8'hdb;
      13'd3364: x = 8'h67;
      13'd3365: x = 8'h9b;
      13'd3366: x = 8'h68;
      13'd3367: x = 8'h9b;
      13'd3368: x = 8'h50;
      13'd3369: x = 8'h8c;
      13'd3370: x = 8'h63;
      13'd3371: x = 8'h8c;
      13'd3372: x = 8'h7f;
      13'd3373: x = 8'h01;
      13'd3374: x = 8'h51;
      13'd3375: x = 8'h07;
      13'd3376: x = 8'h88;
      13'd3377: x = 8'h29;
      13'd3378: x = 8'h84;
      13'd3379: x = 8'h80;
      13'd3380: x = 8'hc4;
      13'd3381: x = 8'h80;
      13'd3382: x = 8'h57;
      13'd3383: x = 8'h71;
      13'd3384: x = 8'h07;
      13'd3385: x = 8'h88;
      13'd3386: x = 8'h14;
      13'd3387: x = 8'hed;
      13'd3388: x = 8'ha5;
      13'd3389: x = 8'had;
      13'd3390: x = 8'haf;
      13'd3391: x = 8'hac;
      13'd3392: x = 8'hed;
      13'd3393: x = 8'ha5;
      13'd3394: x = 8'had;
      13'd3395: x = 8'ha9;
      13'd3396: x = 8'ha8;
      13'd3397: x = 8'hf2;
      13'd3398: x = 8'haf;
      13'd3399: x = 8'hac;
      13'd3400: x = 8'haf;
      13'd3401: x = 8'ha3;
      13'd3402: x = 8'h71;
      13'd3403: x = 8'h08;
      13'd3404: x = 8'h88;
      13'd3405: x = 8'hae;
      13'd3406: x = 8'ha5;
      13'd3407: x = 8'hac;
      13'd3408: x = 8'h68;
      13'd3409: x = 8'h83;
      13'd3410: x = 8'h08;
      13'd3411: x = 8'h68;
      13'd3412: x = 8'h9d;
      13'd3413: x = 8'h08;
      13'd3414: x = 8'h71;
      13'd3415: x = 8'h07;
      13'd3416: x = 8'h88;
      13'd3417: x = 8'h60;
      13'd3418: x = 8'h76;
      13'd3419: x = 8'hb4;
      13'd3420: x = 8'haf;
      13'd3421: x = 8'hae;
      13'd3422: x = 8'h76;
      13'd3423: x = 8'h8d;
      13'd3424: x = 8'h76;
      13'd3425: x = 8'h8b;
      13'd3426: x = 8'h51;
      13'd3427: x = 8'h07;
      13'd3428: x = 8'h88;
      13'd3429: x = 8'h19;
      13'd3430: x = 8'hb8;
      13'd3431: x = 8'ha4;
      13'd3432: x = 8'hae;
      13'd3433: x = 8'hb2;
      13'd3434: x = 8'hf2;
      13'd3435: x = 8'hb3;
      13'd3436: x = 8'hb5;
      13'd3437: x = 8'hf3;
      13'd3438: x = 8'ha2;
      13'd3439: x = 8'ha1;
      13'd3440: x = 8'hee;
      13'd3441: x = 8'ha7;
      13'd3442: x = 8'hb3;
      13'd3443: x = 8'he4;
      13'd3444: x = 8'hae;
      13'd3445: x = 8'hb2;
      13'd3446: x = 8'heb;
      13'd3447: x = 8'ha5;
      13'd3448: x = 8'ha5;
      13'd3449: x = 8'hb0;
      13'd3450: x = 8'h51;
      13'd3451: x = 8'h07;
      13'd3452: x = 8'h88;
      13'd3453: x = 8'h39;
      13'd3454: x = 8'h81;
      13'd3455: x = 8'hc1;
      13'd3456: x = 8'h4f;
      13'd3457: x = 8'h7f;
      13'd3458: x = 8'h0f;
      13'd3459: x = 8'h2f;
      13'd3460: x = 8'h00;
      13'd3461: x = 8'h51;
      13'd3462: x = 8'h06;
      13'd3463: x = 8'h88;
      13'd3464: x = 8'h29;
      13'd3465: x = 8'hc2;
      13'd3466: x = 8'h0c;
      13'd3467: x = 8'h82;
      13'd3468: x = 8'h57;
      13'd3469: x = 8'h8c;
      13'd3470: x = 8'h6a;
      13'd3471: x = 8'h8c;
      13'd3472: x = 8'h42;
      13'd3473: x = 8'hae;
      13'd3474: x = 8'ha5;
      13'd3475: x = 8'ha8;
      13'd3476: x = 8'hb4;
      13'd3477: x = 8'h60;
      13'd3478: x = 8'hae;
      13'd3479: x = 8'ha5;
      13'd3480: x = 8'ha8;
      13'd3481: x = 8'hb4;
      13'd3482: x = 8'h4f;
      13'd3483: x = 8'h7e;
      13'd3484: x = 8'h1e;
      13'd3485: x = 8'h35;
      13'd3486: x = 8'h8c;
      13'd3487: x = 8'h27;
      13'd3488: x = 8'h51;
      13'd3489: x = 8'h07;
      13'd3490: x = 8'h88;
      13'd3491: x = 8'h09;
      13'd3492: x = 8'h8b;
      13'd3493: x = 8'hfe;
      13'd3494: x = 8'he4;
      13'd3495: x = 8'haf;
      13'd3496: x = 8'had;
      13'd3497: x = 8'hf2;
      13'd3498: x = 8'haf;
      13'd3499: x = 8'he4;
      13'd3500: x = 8'hae;
      13'd3501: x = 8'ha1;
      13'd3502: x = 8'hdc;
      13'd3503: x = 8'hde;
      13'd3504: x = 8'h9c;
      13'd3505: x = 8'hdd;
      13'd3506: x = 8'h9c;
      13'd3507: x = 8'hde;
      13'd3508: x = 8'hdd;
      13'd3509: x = 8'h9e;
      13'd3510: x = 8'hc3;
      13'd3511: x = 8'hdd;
      13'd3512: x = 8'hcf;
      13'd3513: x = 8'hca;
      13'd3514: x = 8'hcd;
      13'd3515: x = 8'hcb;
      13'd3516: x = 8'h00;
      13'd3517: x = 8'h47;
      13'd3518: x = 8'h9d;
      13'd3519: x = 8'had;
      13'd3520: x = 8'ha5;
      13'd3521: x = 8'had;
      13'd3522: x = 8'haf;
      13'd3523: x = 8'hac;
      13'd3524: x = 8'h76;
      13'd3525: x = 8'h9d;
      13'd3526: x = 8'had;
      13'd3527: x = 8'ha5;
      13'd3528: x = 8'had;
      13'd3529: x = 8'ha9;
      13'd3530: x = 8'ha8;
      13'd3531: x = 8'he6;
      13'd3532: x = 8'ha6;
      13'd3533: x = 8'haf;
      13'd3534: x = 8'h60;
      13'd3535: x = 8'h8c;
      13'd3536: x = 8'h20;
      13'd3537: x = 8'haf;
      13'd3538: x = 8'hb4;
      13'd3539: x = 8'hb5;
      13'd3540: x = 8'ha1;
      13'd3541: x = 8'hf2;
      13'd3542: x = 8'hac;
      13'd3543: x = 8'ha3;
      13'd3544: x = 8'hf2;
      13'd3545: x = 8'ha3;
      13'd3546: x = 8'hb3;
      13'd3547: x = 8'h60;
      13'd3548: x = 8'h8c;
      13'd3549: x = 8'h20;
      13'd3550: x = 8'hac;
      13'd3551: x = 8'ha5;
      13'd3552: x = 8'ha4;
      13'd3553: x = 8'hee;
      13'd3554: x = 8'hb5;
      13'd3555: x = 8'hb2;
      13'd3556: x = 8'h60;
      13'd3557: x = 8'hae;
      13'd3558: x = 8'hb5;
      13'd3559: x = 8'hb2;
      13'd3560: x = 8'hf4;
      13'd3561: x = 8'hb3;
      13'd3562: x = 8'ha9;
      13'd3563: x = 8'hac;
      13'd3564: x = 8'h60;
      13'd3565: x = 8'h8c;
      13'd3566: x = 8'h20;
      13'd3567: x = 8'hb4;
      13'd3568: x = 8'hb3;
      13'd3569: x = 8'ha9;
      13'd3570: x = 8'hac;
      13'd3571: x = 8'h7a;
      13'd3572: x = 8'h7e;
      13'd3573: x = 8'h9a;
      13'd3574: x = 8'h22;
      13'd3575: x = 8'h20;
      13'd3576: x = 8'h00;
      13'd3577: x = 8'h60;
      13'd3578: x = 8'h03;
      13'd3579: x = 8'hbf;
      13'd3580: x = 8'h60;
      13'd3581: x = 8'h03;
      13'd3582: x = 8'hbf;
      13'd3583: x = 8'h1f;
      13'd3584: x = 8'h20;
      13'd3585: x = 8'hb1;
      13'd3586: x = 8'he7;
      13'd3587: x = 8'he8;
      13'd3588: x = 8'he8;
      13'd3589: x = 8'hb5;
      13'd3590: x = 8'h4f;
      13'd3591: x = 8'h85;
      13'd3592: x = 8'hda;
      13'd3593: x = 8'hb5;
      13'd3594: x = 8'h77;
      13'd3595: x = 8'h85;
      13'd3596: x = 8'hdb;
      13'd3597: x = 8'hb4;
      13'd3598: x = 8'h4e;
      13'd3599: x = 8'h98;
      13'd3600: x = 8'hd5;
      13'd3601: x = 8'h76;
      13'd3602: x = 8'hb0;
      13'd3603: x = 8'h09;
      13'd3604: x = 8'hb1;
      13'd3605: x = 8'hda;
      13'd3606: x = 8'h20;
      13'd3607: x = 8'hc9;
      13'd3608: x = 8'he3;
      13'd3609: x = 8'hc8;
      13'd3610: x = 8'h4c;
      13'd3611: x = 8'h0f;
      13'd3612: x = 8'hee;
      13'd3613: x = 8'ha9;
      13'd3614: x = 8'hff;
      13'd3615: x = 8'h85;
      13'd3616: x = 8'hd5;
      13'd3617: x = 8'h60;
      13'd3618: x = 8'he8;
      13'd3619: x = 8'ha9;
      13'd3620: x = 8'h00;
      13'd3621: x = 8'h95;
      13'd3622: x = 8'h78;
      13'd3623: x = 8'h95;
      13'd3624: x = 8'ha0;
      13'd3625: x = 8'hb5;
      13'd3626: x = 8'h77;
      13'd3627: x = 8'h38;
      13'd3628: x = 8'hf5;
      13'd3629: x = 8'h4f;
      13'd3630: x = 8'h95;
      13'd3631: x = 8'h50;
      13'd3632: x = 8'h4c;
      13'd3633: x = 8'h23;
      13'd3634: x = 8'he8;
      13'd3635: x = 8'hff;
      13'd3636: x = 8'h20;
      13'd3637: x = 8'h15;
      13'd3638: x = 8'he7;
      13'd3639: x = 8'ha5;
      13'd3640: x = 8'hcf;
      13'd3641: x = 8'hd0;
      13'd3642: x = 8'h28;
      13'd3643: x = 8'ha5;
      13'd3644: x = 8'hce;
      13'd3645: x = 8'h60;
      13'd3646: x = 8'h20;
      13'd3647: x = 8'h34;
      13'd3648: x = 8'hee;
      13'd3649: x = 8'ha4;
      13'd3650: x = 8'hc8;
      13'd3651: x = 8'hc9;
      13'd3652: x = 8'h30;
      13'd3653: x = 8'hb0;
      13'd3654: x = 8'h21;
      13'd3655: x = 8'hc0;
      13'd3656: x = 8'h28;
      13'd3657: x = 8'hb0;
      13'd3658: x = 8'h1d;
      13'd3659: x = 8'h60;
      13'd3660: x = 8'hea;
      13'd3661: x = 8'hea;
      13'd3662: x = 8'h20;
      13'd3663: x = 8'h34;
      13'd3664: x = 8'hee;
      13'd3665: x = 8'h60;
      13'd3666: x = 8'hea;
      13'd3667: x = 8'h8a;
      13'd3668: x = 8'ha2;
      13'd3669: x = 8'h01;
      13'd3670: x = 8'hb4;
      13'd3671: x = 8'hce;
      13'd3672: x = 8'h94;
      13'd3673: x = 8'h4c;
      13'd3674: x = 8'hb4;
      13'd3675: x = 8'h48;
      13'd3676: x = 8'h94;
      13'd3677: x = 8'hca;
      13'd3678: x = 8'hca;
      13'd3679: x = 8'hf0;
      13'd3680: x = 8'hf5;
      13'd3681: x = 8'haa;
      13'd3682: x = 8'h60;
      13'd3683: x = 8'ha0;
      13'd3684: x = 8'h77;
      13'd3685: x = 8'h4c;
      13'd3686: x = 8'he0;
      13'd3687: x = 8'he3;
      13'd3688: x = 8'ha0;
      13'd3689: x = 8'h7b;
      13'd3690: x = 8'hd0;
      13'd3691: x = 8'hf9;
      13'd3692: x = 8'h20;
      13'd3693: x = 8'h54;
      13'd3694: x = 8'he2;
      13'd3695: x = 8'ha5;
      13'd3696: x = 8'hda;
      13'd3697: x = 8'hd0;
      13'd3698: x = 8'h07;
      13'd3699: x = 8'ha5;
      13'd3700: x = 8'hdb;
      13'd3701: x = 8'hd0;
      13'd3702: x = 8'h03;
      13'd3703: x = 8'h4c;
      13'd3704: x = 8'h7e;
      13'd3705: x = 8'he7;
      13'd3706: x = 8'h06;
      13'd3707: x = 8'hce;
      13'd3708: x = 8'h26;
      13'd3709: x = 8'hcf;
      13'd3710: x = 8'h26;
      13'd3711: x = 8'he6;
      13'd3712: x = 8'h26;
      13'd3713: x = 8'he7;
      13'd3714: x = 8'ha5;
      13'd3715: x = 8'he6;
      13'd3716: x = 8'hc5;
      13'd3717: x = 8'hda;
      13'd3718: x = 8'ha5;
      13'd3719: x = 8'he7;
      13'd3720: x = 8'he5;
      13'd3721: x = 8'hdb;
      13'd3722: x = 8'h90;
      13'd3723: x = 8'h0a;
      13'd3724: x = 8'h85;
      13'd3725: x = 8'he7;
      13'd3726: x = 8'ha5;
      13'd3727: x = 8'he6;
      13'd3728: x = 8'he5;
      13'd3729: x = 8'hda;
      13'd3730: x = 8'h85;
      13'd3731: x = 8'he6;
      13'd3732: x = 8'he6;
      13'd3733: x = 8'hce;
      13'd3734: x = 8'h88;
      13'd3735: x = 8'hd0;
      13'd3736: x = 8'he1;
      13'd3737: x = 8'h60;
      13'd3738: x = 8'hff;
      13'd3739: x = 8'hff;
      13'd3740: x = 8'hff;
      13'd3741: x = 8'hff;
      13'd3742: x = 8'hff;
      13'd3743: x = 8'hff;
      13'd3744: x = 8'h20;
      13'd3745: x = 8'h15;
      13'd3746: x = 8'he7;
      13'd3747: x = 8'h6c;
      13'd3748: x = 8'hce;
      13'd3749: x = 8'h00;
      13'd3750: x = 8'ha5;
      13'd3751: x = 8'h4c;
      13'd3752: x = 8'hd0;
      13'd3753: x = 8'h02;
      13'd3754: x = 8'hc6;
      13'd3755: x = 8'h4d;
      13'd3756: x = 8'hc6;
      13'd3757: x = 8'h4c;
      13'd3758: x = 8'ha5;
      13'd3759: x = 8'h48;
      13'd3760: x = 8'hd0;
      13'd3761: x = 8'h02;
      13'd3762: x = 8'hc6;
      13'd3763: x = 8'h49;
      13'd3764: x = 8'hc6;
      13'd3765: x = 8'h48;
      13'd3766: x = 8'ha0;
      13'd3767: x = 8'h00;
      13'd3768: x = 8'hb1;
      13'd3769: x = 8'h4c;
      13'd3770: x = 8'h91;
      13'd3771: x = 8'h48;
      13'd3772: x = 8'ha5;
      13'd3773: x = 8'hca;
      13'd3774: x = 8'hc5;
      13'd3775: x = 8'h4c;
      13'd3776: x = 8'ha5;
      13'd3777: x = 8'hcb;
      13'd3778: x = 8'he5;
      13'd3779: x = 8'h4d;
      13'd3780: x = 8'h90;
      13'd3781: x = 8'he0;
      13'd3782: x = 8'h4c;
      13'd3783: x = 8'h53;
      13'd3784: x = 8'hee;
      13'd3785: x = 8'hc9;
      13'd3786: x = 8'h28;
      13'd3787: x = 8'hb0;
      13'd3788: x = 8'h9b;
      13'd3789: x = 8'ha8;
      13'd3790: x = 8'ha5;
      13'd3791: x = 8'hc8;
      13'd3792: x = 8'h60;
      13'd3793: x = 8'hea;
      13'd3794: x = 8'hea;
      13'd3795: x = 8'h98;
      13'd3796: x = 8'haa;
      13'd3797: x = 8'ha0;
      13'd3798: x = 8'h6e;
      13'd3799: x = 8'h20;
      13'd3800: x = 8'hc4;
      13'd3801: x = 8'he3;
      13'd3802: x = 8'h8a;
      13'd3803: x = 8'ha8;
      13'd3804: x = 8'h20;
      13'd3805: x = 8'hc4;
      13'd3806: x = 8'he3;
      13'd3807: x = 8'ha0;
      13'd3808: x = 8'h72;
      13'd3809: x = 8'h4c;
      13'd3810: x = 8'hc4;
      13'd3811: x = 8'he3;
      13'd3812: x = 8'h20;
      13'd3813: x = 8'h15;
      13'd3814: x = 8'he7;
      13'd3815: x = 8'h06;
      13'd3816: x = 8'hce;
      13'd3817: x = 8'h26;
      13'd3818: x = 8'hcf;
      13'd3819: x = 8'h30;
      13'd3820: x = 8'hfa;
      13'd3821: x = 8'hb0;
      13'd3822: x = 8'hdc;
      13'd3823: x = 8'hd0;
      13'd3824: x = 8'h04;
      13'd3825: x = 8'hc5;
      13'd3826: x = 8'hce;
      13'd3827: x = 8'hb0;
      13'd3828: x = 8'hd6;
      13'd3829: x = 8'h60;
      13'd3830: x = 8'h20;
      13'd3831: x = 8'h15;
      13'd3832: x = 8'he7;
      13'd3833: x = 8'hb1;
      13'd3834: x = 8'hce;
      13'd3835: x = 8'h94;
      13'd3836: x = 8'h9f;
      13'd3837: x = 8'h4c;
      13'd3838: x = 8'h08;
      13'd3839: x = 8'he7;
      13'd3840: x = 8'h20;
      13'd3841: x = 8'h34;
      13'd3842: x = 8'hee;
      13'd3843: x = 8'ha5;
      13'd3844: x = 8'hce;
      13'd3845: x = 8'h48;
      13'd3846: x = 8'h20;
      13'd3847: x = 8'h15;
      13'd3848: x = 8'he7;
      13'd3849: x = 8'h68;
      13'd3850: x = 8'h91;
      13'd3851: x = 8'hce;
      13'd3852: x = 8'h60;
      13'd3853: x = 8'hff;
      13'd3854: x = 8'hff;
      13'd3855: x = 8'hff;
      13'd3856: x = 8'h20;
      13'd3857: x = 8'h6c;
      13'd3858: x = 8'hee;
      13'd3859: x = 8'ha5;
      13'd3860: x = 8'hce;
      13'd3861: x = 8'h85;
      13'd3862: x = 8'he6;
      13'd3863: x = 8'ha5;
      13'd3864: x = 8'hcf;
      13'd3865: x = 8'h85;
      13'd3866: x = 8'he7;
      13'd3867: x = 8'h4c;
      13'd3868: x = 8'h44;
      13'd3869: x = 8'he2;
      13'd3870: x = 8'h20;
      13'd3871: x = 8'he4;
      13'd3872: x = 8'hee;
      13'd3873: x = 8'h4c;
      13'd3874: x = 8'h34;
      13'd3875: x = 8'he1;
      13'd3876: x = 8'h20;
      13'd3877: x = 8'he4;
      13'd3878: x = 8'hee;
      13'd3879: x = 8'hb4;
      13'd3880: x = 8'h78;
      13'd3881: x = 8'hb5;
      13'd3882: x = 8'h50;
      13'd3883: x = 8'h69;
      13'd3884: x = 8'hfe;
      13'd3885: x = 8'hb0;
      13'd3886: x = 8'h01;
      13'd3887: x = 8'h88;
      13'd3888: x = 8'h85;
      13'd3889: x = 8'hda;
      13'd3890: x = 8'h84;
      13'd3891: x = 8'hdb;
      13'd3892: x = 8'h18;
      13'd3893: x = 8'h65;
      13'd3894: x = 8'hce;
      13'd3895: x = 8'h95;
      13'd3896: x = 8'h50;
      13'd3897: x = 8'h98;
      13'd3898: x = 8'h65;
      13'd3899: x = 8'hcf;
      13'd3900: x = 8'h95;
      13'd3901: x = 8'h78;
      13'd3902: x = 8'ha0;
      13'd3903: x = 8'h00;
      13'd3904: x = 8'hb5;
      13'd3905: x = 8'h50;
      13'd3906: x = 8'hd1;
      13'd3907: x = 8'hda;
      13'd3908: x = 8'hc8;
      13'd3909: x = 8'hb5;
      13'd3910: x = 8'h78;
      13'd3911: x = 8'hf1;
      13'd3912: x = 8'hda;
      13'd3913: x = 8'hb0;
      13'd3914: x = 8'h80;
      13'd3915: x = 8'h4c;
      13'd3916: x = 8'h23;
      13'd3917: x = 8'he8;
      13'd3918: x = 8'h20;
      13'd3919: x = 8'h15;
      13'd3920: x = 8'he7;
      13'd3921: x = 8'ha5;
      13'd3922: x = 8'h4e;
      13'd3923: x = 8'h20;
      13'd3924: x = 8'h08;
      13'd3925: x = 8'he7;
      13'd3926: x = 8'ha5;
      13'd3927: x = 8'h4f;
      13'd3928: x = 8'hd0;
      13'd3929: x = 8'h04;
      13'd3930: x = 8'hc5;
      13'd3931: x = 8'h4e;
      13'd3932: x = 8'h69;
      13'd3933: x = 8'h00;
      13'd3934: x = 8'h29;
      13'd3935: x = 8'h7f;
      13'd3936: x = 8'h85;
      13'd3937: x = 8'h4f;
      13'd3938: x = 8'h95;
      13'd3939: x = 8'ha0;
      13'd3940: x = 8'ha0;
      13'd3941: x = 8'h11;
      13'd3942: x = 8'ha5;
      13'd3943: x = 8'h4f;
      13'd3944: x = 8'h0a;
      13'd3945: x = 8'h18;
      13'd3946: x = 8'h69;
      13'd3947: x = 8'h40;
      13'd3948: x = 8'h0a;
      13'd3949: x = 8'h26;
      13'd3950: x = 8'h4e;
      13'd3951: x = 8'h26;
      13'd3952: x = 8'h4f;
      13'd3953: x = 8'h88;
      13'd3954: x = 8'hd0;
      13'd3955: x = 8'hf2;
      13'd3956: x = 8'ha5;
      13'd3957: x = 8'hce;
      13'd3958: x = 8'h20;
      13'd3959: x = 8'h08;
      13'd3960: x = 8'he7;
      13'd3961: x = 8'ha5;
      13'd3962: x = 8'hcf;
      13'd3963: x = 8'h95;
      13'd3964: x = 8'ha0;
      13'd3965: x = 8'h4c;
      13'd3966: x = 8'h7a;
      13'd3967: x = 8'he2;
      13'd3968: x = 8'h20;
      13'd3969: x = 8'h15;
      13'd3970: x = 8'he7;
      13'd3971: x = 8'ha4;
      13'd3972: x = 8'hce;
      13'd3973: x = 8'hc4;
      13'd3974: x = 8'h4c;
      13'd3975: x = 8'ha5;
      13'd3976: x = 8'hcf;
      13'd3977: x = 8'he5;
      13'd3978: x = 8'h4d;
      13'd3979: x = 8'h90;
      13'd3980: x = 8'h1f;
      13'd3981: x = 8'h84;
      13'd3982: x = 8'h48;
      13'd3983: x = 8'ha5;
      13'd3984: x = 8'hcf;
      13'd3985: x = 8'h85;
      13'd3986: x = 8'h49;
      13'd3987: x = 8'h4c;
      13'd3988: x = 8'hb6;
      13'd3989: x = 8'hee;
      13'd3990: x = 8'h20;
      13'd3991: x = 8'h15;
      13'd3992: x = 8'he7;
      13'd3993: x = 8'ha4;
      13'd3994: x = 8'hce;
      13'd3995: x = 8'hc4;
      13'd3996: x = 8'hca;
      13'd3997: x = 8'ha5;
      13'd3998: x = 8'hcf;
      13'd3999: x = 8'he5;
      13'd4000: x = 8'hcb;
      13'd4001: x = 8'hb0;
      13'd4002: x = 8'h09;
      13'd4003: x = 8'h84;
      13'd4004: x = 8'h4a;
      13'd4005: x = 8'ha5;
      13'd4006: x = 8'hcf;
      13'd4007: x = 8'h85;
      13'd4008: x = 8'h4b;
      13'd4009: x = 8'h4c;
      13'd4010: x = 8'hb7;
      13'd4011: x = 8'he5;
      13'd4012: x = 8'h4c;
      13'd4013: x = 8'hcb;
      13'd4014: x = 8'hee;
      13'd4015: x = 8'hea;
      13'd4016: x = 8'hea;
      13'd4017: x = 8'hea;
      13'd4018: x = 8'hea;
      13'd4019: x = 8'h20;
      13'd4020: x = 8'hc9;
      13'd4021: x = 8'hef;
      13'd4022: x = 8'h20;
      13'd4023: x = 8'h71;
      13'd4024: x = 8'he1;
      13'd4025: x = 8'h4c;
      13'd4026: x = 8'hbf;
      13'd4027: x = 8'hef;
      13'd4028: x = 8'h20;
      13'd4029: x = 8'h03;
      13'd4030: x = 8'hee;
      13'd4031: x = 8'ha9;
      13'd4032: x = 8'hff;
      13'd4033: x = 8'h85;
      13'd4034: x = 8'hc8;
      13'd4035: x = 8'ha9;
      13'd4036: x = 8'h74;
      13'd4037: x = 8'h8d;
      13'd4038: x = 8'h00;
      13'd4039: x = 8'h02;
      13'd4040: x = 8'h60;
      13'd4041: x = 8'h20;
      13'd4042: x = 8'h36;
      13'd4043: x = 8'he7;
      13'd4044: x = 8'he8;
      13'd4045: x = 8'h20;
      13'd4046: x = 8'h36;
      13'd4047: x = 8'he7;
      13'd4048: x = 8'hb5;
      13'd4049: x = 8'h50;
      13'd4050: x = 8'h60;
      13'd4051: x = 8'ha9;
      13'd4052: x = 8'h00;
      13'd4053: x = 8'h85;
      13'd4054: x = 8'h4a;
      13'd4055: x = 8'h85;
      13'd4056: x = 8'h4c;
      13'd4057: x = 8'ha9;
      13'd4058: x = 8'h08;
      13'd4059: x = 8'h85;
      13'd4060: x = 8'h4b;
      13'd4061: x = 8'ha9;
      13'd4062: x = 8'h10;
      13'd4063: x = 8'h85;
      13'd4064: x = 8'h4d;
      13'd4065: x = 8'h4c;
      13'd4066: x = 8'had;
      13'd4067: x = 8'he5;
      13'd4068: x = 8'hd5;
      13'd4069: x = 8'h78;
      13'd4070: x = 8'hd0;
      13'd4071: x = 8'h01;
      13'd4072: x = 8'h18;
      13'd4073: x = 8'h4c;
      13'd4074: x = 8'h02;
      13'd4075: x = 8'he1;
      13'd4076: x = 8'h20;
      13'd4077: x = 8'hb7;
      13'd4078: x = 8'he5;
      13'd4079: x = 8'h4c;
      13'd4080: x = 8'h36;
      13'd4081: x = 8'he8;
      13'd4082: x = 8'h20;
      13'd4083: x = 8'hb7;
      13'd4084: x = 8'he5;
      13'd4085: x = 8'h4c;
      13'd4086: x = 8'h5b;
      13'd4087: x = 8'he8;
      13'd4088: x = 8'he0;
      13'd4089: x = 8'h80;
      13'd4090: x = 8'hd0;
      13'd4091: x = 8'h01;
      13'd4092: x = 8'h88;
      13'd4093: x = 8'h4c;
      13'd4094: x = 8'h0c;
      13'd4095: x = 8'he0;
      13'd4096: x = 8'h00;
      13'd4097: x = 8'h00;
      13'd4098: x = 8'h00;
      13'd4099: x = 8'h00;
      13'd4100: x = 8'h00;
      13'd4101: x = 8'h00;
      13'd4102: x = 8'h00;
      13'd4103: x = 8'h00;
      13'd4104: x = 8'h00;
      13'd4105: x = 8'h00;
      13'd4106: x = 8'h00;
      13'd4107: x = 8'h00;
      13'd4108: x = 8'h00;
      13'd4109: x = 8'h00;
      13'd4110: x = 8'h00;
      13'd4111: x = 8'h00;
      13'd4112: x = 8'h00;
      13'd4113: x = 8'h00;
      13'd4114: x = 8'h00;
      13'd4115: x = 8'h00;
      13'd4116: x = 8'h00;
      13'd4117: x = 8'h00;
      13'd4118: x = 8'h00;
      13'd4119: x = 8'h00;
      13'd4120: x = 8'h00;
      13'd4121: x = 8'h00;
      13'd4122: x = 8'h00;
      13'd4123: x = 8'h00;
      13'd4124: x = 8'h00;
      13'd4125: x = 8'h00;
      13'd4126: x = 8'h00;
      13'd4127: x = 8'h00;
      13'd4128: x = 8'h00;
      13'd4129: x = 8'h00;
      13'd4130: x = 8'h00;
      13'd4131: x = 8'h00;
      13'd4132: x = 8'h00;
      13'd4133: x = 8'h00;
      13'd4134: x = 8'h00;
      13'd4135: x = 8'h00;
      13'd4136: x = 8'h00;
      13'd4137: x = 8'h00;
      13'd4138: x = 8'h00;
      13'd4139: x = 8'h00;
      13'd4140: x = 8'h00;
      13'd4141: x = 8'h00;
      13'd4142: x = 8'h00;
      13'd4143: x = 8'h00;
      13'd4144: x = 8'h00;
      13'd4145: x = 8'h00;
      13'd4146: x = 8'h00;
      13'd4147: x = 8'h00;
      13'd4148: x = 8'h00;
      13'd4149: x = 8'h00;
      13'd4150: x = 8'h00;
      13'd4151: x = 8'h00;
      13'd4152: x = 8'h00;
      13'd4153: x = 8'h00;
      13'd4154: x = 8'h00;
      13'd4155: x = 8'h00;
      13'd4156: x = 8'h00;
      13'd4157: x = 8'h00;
      13'd4158: x = 8'h00;
      13'd4159: x = 8'h00;
      13'd4160: x = 8'h00;
      13'd4161: x = 8'h00;
      13'd4162: x = 8'h00;
      13'd4163: x = 8'h00;
      13'd4164: x = 8'h00;
      13'd4165: x = 8'h00;
      13'd4166: x = 8'h00;
      13'd4167: x = 8'h00;
      13'd4168: x = 8'h00;
      13'd4169: x = 8'h00;
      13'd4170: x = 8'h00;
      13'd4171: x = 8'h00;
      13'd4172: x = 8'h00;
      13'd4173: x = 8'h00;
      13'd4174: x = 8'h00;
      13'd4175: x = 8'h00;
      13'd4176: x = 8'h00;
      13'd4177: x = 8'h00;
      13'd4178: x = 8'h00;
      13'd4179: x = 8'h00;
      13'd4180: x = 8'h00;
      13'd4181: x = 8'h00;
      13'd4182: x = 8'h00;
      13'd4183: x = 8'h00;
      13'd4184: x = 8'h00;
      13'd4185: x = 8'h00;
      13'd4186: x = 8'h00;
      13'd4187: x = 8'h00;
      13'd4188: x = 8'h00;
      13'd4189: x = 8'h00;
      13'd4190: x = 8'h00;
      13'd4191: x = 8'h00;
      13'd4192: x = 8'h00;
      13'd4193: x = 8'h00;
      13'd4194: x = 8'h00;
      13'd4195: x = 8'h00;
      13'd4196: x = 8'h00;
      13'd4197: x = 8'h00;
      13'd4198: x = 8'h00;
      13'd4199: x = 8'h00;
      13'd4200: x = 8'h00;
      13'd4201: x = 8'h00;
      13'd4202: x = 8'h00;
      13'd4203: x = 8'h00;
      13'd4204: x = 8'h00;
      13'd4205: x = 8'h00;
      13'd4206: x = 8'h00;
      13'd4207: x = 8'h00;
      13'd4208: x = 8'h00;
      13'd4209: x = 8'h00;
      13'd4210: x = 8'h00;
      13'd4211: x = 8'h00;
      13'd4212: x = 8'h00;
      13'd4213: x = 8'h00;
      13'd4214: x = 8'h00;
      13'd4215: x = 8'h00;
      13'd4216: x = 8'h00;
      13'd4217: x = 8'h00;
      13'd4218: x = 8'h00;
      13'd4219: x = 8'h00;
      13'd4220: x = 8'h00;
      13'd4221: x = 8'h00;
      13'd4222: x = 8'h00;
      13'd4223: x = 8'h00;
      13'd4224: x = 8'h00;
      13'd4225: x = 8'h00;
      13'd4226: x = 8'h00;
      13'd4227: x = 8'h00;
      13'd4228: x = 8'h00;
      13'd4229: x = 8'h00;
      13'd4230: x = 8'h00;
      13'd4231: x = 8'h00;
      13'd4232: x = 8'h00;
      13'd4233: x = 8'h00;
      13'd4234: x = 8'h00;
      13'd4235: x = 8'h00;
      13'd4236: x = 8'h00;
      13'd4237: x = 8'h00;
      13'd4238: x = 8'h00;
      13'd4239: x = 8'h00;
      13'd4240: x = 8'h00;
      13'd4241: x = 8'h00;
      13'd4242: x = 8'h00;
      13'd4243: x = 8'h00;
      13'd4244: x = 8'h00;
      13'd4245: x = 8'h00;
      13'd4246: x = 8'h00;
      13'd4247: x = 8'h00;
      13'd4248: x = 8'h00;
      13'd4249: x = 8'h00;
      13'd4250: x = 8'h00;
      13'd4251: x = 8'h00;
      13'd4252: x = 8'h00;
      13'd4253: x = 8'h00;
      13'd4254: x = 8'h00;
      13'd4255: x = 8'h00;
      13'd4256: x = 8'h00;
      13'd4257: x = 8'h00;
      13'd4258: x = 8'h00;
      13'd4259: x = 8'h00;
      13'd4260: x = 8'h00;
      13'd4261: x = 8'h00;
      13'd4262: x = 8'h00;
      13'd4263: x = 8'h00;
      13'd4264: x = 8'h00;
      13'd4265: x = 8'h00;
      13'd4266: x = 8'h00;
      13'd4267: x = 8'h00;
      13'd4268: x = 8'h00;
      13'd4269: x = 8'h00;
      13'd4270: x = 8'h00;
      13'd4271: x = 8'h00;
      13'd4272: x = 8'h00;
      13'd4273: x = 8'h00;
      13'd4274: x = 8'h00;
      13'd4275: x = 8'h00;
      13'd4276: x = 8'h00;
      13'd4277: x = 8'h00;
      13'd4278: x = 8'h00;
      13'd4279: x = 8'h00;
      13'd4280: x = 8'h00;
      13'd4281: x = 8'h00;
      13'd4282: x = 8'h00;
      13'd4283: x = 8'h00;
      13'd4284: x = 8'h00;
      13'd4285: x = 8'h00;
      13'd4286: x = 8'h00;
      13'd4287: x = 8'h00;
      13'd4288: x = 8'h00;
      13'd4289: x = 8'h00;
      13'd4290: x = 8'h00;
      13'd4291: x = 8'h00;
      13'd4292: x = 8'h00;
      13'd4293: x = 8'h00;
      13'd4294: x = 8'h00;
      13'd4295: x = 8'h00;
      13'd4296: x = 8'h00;
      13'd4297: x = 8'h00;
      13'd4298: x = 8'h00;
      13'd4299: x = 8'h00;
      13'd4300: x = 8'h00;
      13'd4301: x = 8'h00;
      13'd4302: x = 8'h00;
      13'd4303: x = 8'h00;
      13'd4304: x = 8'h00;
      13'd4305: x = 8'h00;
      13'd4306: x = 8'h00;
      13'd4307: x = 8'h00;
      13'd4308: x = 8'h00;
      13'd4309: x = 8'h00;
      13'd4310: x = 8'h00;
      13'd4311: x = 8'h00;
      13'd4312: x = 8'h00;
      13'd4313: x = 8'h00;
      13'd4314: x = 8'h00;
      13'd4315: x = 8'h00;
      13'd4316: x = 8'h00;
      13'd4317: x = 8'h00;
      13'd4318: x = 8'h00;
      13'd4319: x = 8'h00;
      13'd4320: x = 8'h00;
      13'd4321: x = 8'h00;
      13'd4322: x = 8'h00;
      13'd4323: x = 8'h00;
      13'd4324: x = 8'h00;
      13'd4325: x = 8'h00;
      13'd4326: x = 8'h00;
      13'd4327: x = 8'h00;
      13'd4328: x = 8'h00;
      13'd4329: x = 8'h00;
      13'd4330: x = 8'h00;
      13'd4331: x = 8'h00;
      13'd4332: x = 8'h00;
      13'd4333: x = 8'h00;
      13'd4334: x = 8'h00;
      13'd4335: x = 8'h00;
      13'd4336: x = 8'h00;
      13'd4337: x = 8'h00;
      13'd4338: x = 8'h00;
      13'd4339: x = 8'h00;
      13'd4340: x = 8'h00;
      13'd4341: x = 8'h00;
      13'd4342: x = 8'h00;
      13'd4343: x = 8'h00;
      13'd4344: x = 8'h00;
      13'd4345: x = 8'h00;
      13'd4346: x = 8'h00;
      13'd4347: x = 8'h00;
      13'd4348: x = 8'h00;
      13'd4349: x = 8'h00;
      13'd4350: x = 8'h00;
      13'd4351: x = 8'h00;
      13'd4352: x = 8'h00;
      13'd4353: x = 8'h00;
      13'd4354: x = 8'h00;
      13'd4355: x = 8'h00;
      13'd4356: x = 8'h00;
      13'd4357: x = 8'h00;
      13'd4358: x = 8'h00;
      13'd4359: x = 8'h00;
      13'd4360: x = 8'h00;
      13'd4361: x = 8'h00;
      13'd4362: x = 8'h00;
      13'd4363: x = 8'h00;
      13'd4364: x = 8'h00;
      13'd4365: x = 8'h00;
      13'd4366: x = 8'h00;
      13'd4367: x = 8'h00;
      13'd4368: x = 8'h00;
      13'd4369: x = 8'h00;
      13'd4370: x = 8'h00;
      13'd4371: x = 8'h00;
      13'd4372: x = 8'h00;
      13'd4373: x = 8'h00;
      13'd4374: x = 8'h00;
      13'd4375: x = 8'h00;
      13'd4376: x = 8'h00;
      13'd4377: x = 8'h00;
      13'd4378: x = 8'h00;
      13'd4379: x = 8'h00;
      13'd4380: x = 8'h00;
      13'd4381: x = 8'h00;
      13'd4382: x = 8'h00;
      13'd4383: x = 8'h00;
      13'd4384: x = 8'h00;
      13'd4385: x = 8'h00;
      13'd4386: x = 8'h00;
      13'd4387: x = 8'h00;
      13'd4388: x = 8'h00;
      13'd4389: x = 8'h00;
      13'd4390: x = 8'h00;
      13'd4391: x = 8'h00;
      13'd4392: x = 8'h00;
      13'd4393: x = 8'h00;
      13'd4394: x = 8'h00;
      13'd4395: x = 8'h00;
      13'd4396: x = 8'h00;
      13'd4397: x = 8'h00;
      13'd4398: x = 8'h00;
      13'd4399: x = 8'h00;
      13'd4400: x = 8'h00;
      13'd4401: x = 8'h00;
      13'd4402: x = 8'h00;
      13'd4403: x = 8'h00;
      13'd4404: x = 8'h00;
      13'd4405: x = 8'h00;
      13'd4406: x = 8'h00;
      13'd4407: x = 8'h00;
      13'd4408: x = 8'h00;
      13'd4409: x = 8'h00;
      13'd4410: x = 8'h00;
      13'd4411: x = 8'h00;
      13'd4412: x = 8'h00;
      13'd4413: x = 8'h00;
      13'd4414: x = 8'h00;
      13'd4415: x = 8'h00;
      13'd4416: x = 8'h00;
      13'd4417: x = 8'h00;
      13'd4418: x = 8'h00;
      13'd4419: x = 8'h00;
      13'd4420: x = 8'h00;
      13'd4421: x = 8'h00;
      13'd4422: x = 8'h00;
      13'd4423: x = 8'h00;
      13'd4424: x = 8'h00;
      13'd4425: x = 8'h00;
      13'd4426: x = 8'h00;
      13'd4427: x = 8'h00;
      13'd4428: x = 8'h00;
      13'd4429: x = 8'h00;
      13'd4430: x = 8'h00;
      13'd4431: x = 8'h00;
      13'd4432: x = 8'h00;
      13'd4433: x = 8'h00;
      13'd4434: x = 8'h00;
      13'd4435: x = 8'h00;
      13'd4436: x = 8'h00;
      13'd4437: x = 8'h00;
      13'd4438: x = 8'h00;
      13'd4439: x = 8'h00;
      13'd4440: x = 8'h00;
      13'd4441: x = 8'h00;
      13'd4442: x = 8'h00;
      13'd4443: x = 8'h00;
      13'd4444: x = 8'h00;
      13'd4445: x = 8'h00;
      13'd4446: x = 8'h00;
      13'd4447: x = 8'h00;
      13'd4448: x = 8'h00;
      13'd4449: x = 8'h00;
      13'd4450: x = 8'h00;
      13'd4451: x = 8'h00;
      13'd4452: x = 8'h00;
      13'd4453: x = 8'h00;
      13'd4454: x = 8'h00;
      13'd4455: x = 8'h00;
      13'd4456: x = 8'h00;
      13'd4457: x = 8'h00;
      13'd4458: x = 8'h00;
      13'd4459: x = 8'h00;
      13'd4460: x = 8'h00;
      13'd4461: x = 8'h00;
      13'd4462: x = 8'h00;
      13'd4463: x = 8'h00;
      13'd4464: x = 8'h00;
      13'd4465: x = 8'h00;
      13'd4466: x = 8'h00;
      13'd4467: x = 8'h00;
      13'd4468: x = 8'h00;
      13'd4469: x = 8'h00;
      13'd4470: x = 8'h00;
      13'd4471: x = 8'h00;
      13'd4472: x = 8'h00;
      13'd4473: x = 8'h00;
      13'd4474: x = 8'h00;
      13'd4475: x = 8'h00;
      13'd4476: x = 8'h00;
      13'd4477: x = 8'h00;
      13'd4478: x = 8'h00;
      13'd4479: x = 8'h00;
      13'd4480: x = 8'h00;
      13'd4481: x = 8'h00;
      13'd4482: x = 8'h00;
      13'd4483: x = 8'h00;
      13'd4484: x = 8'h00;
      13'd4485: x = 8'h00;
      13'd4486: x = 8'h00;
      13'd4487: x = 8'h00;
      13'd4488: x = 8'h00;
      13'd4489: x = 8'h00;
      13'd4490: x = 8'h00;
      13'd4491: x = 8'h00;
      13'd4492: x = 8'h00;
      13'd4493: x = 8'h00;
      13'd4494: x = 8'h00;
      13'd4495: x = 8'h00;
      13'd4496: x = 8'h00;
      13'd4497: x = 8'h00;
      13'd4498: x = 8'h00;
      13'd4499: x = 8'h00;
      13'd4500: x = 8'h00;
      13'd4501: x = 8'h00;
      13'd4502: x = 8'h00;
      13'd4503: x = 8'h00;
      13'd4504: x = 8'h00;
      13'd4505: x = 8'h00;
      13'd4506: x = 8'h00;
      13'd4507: x = 8'h00;
      13'd4508: x = 8'h00;
      13'd4509: x = 8'h00;
      13'd4510: x = 8'h00;
      13'd4511: x = 8'h00;
      13'd4512: x = 8'h00;
      13'd4513: x = 8'h00;
      13'd4514: x = 8'h00;
      13'd4515: x = 8'h00;
      13'd4516: x = 8'h00;
      13'd4517: x = 8'h00;
      13'd4518: x = 8'h00;
      13'd4519: x = 8'h00;
      13'd4520: x = 8'h00;
      13'd4521: x = 8'h00;
      13'd4522: x = 8'h00;
      13'd4523: x = 8'h00;
      13'd4524: x = 8'h00;
      13'd4525: x = 8'h00;
      13'd4526: x = 8'h00;
      13'd4527: x = 8'h00;
      13'd4528: x = 8'h00;
      13'd4529: x = 8'h00;
      13'd4530: x = 8'h00;
      13'd4531: x = 8'h00;
      13'd4532: x = 8'h00;
      13'd4533: x = 8'h00;
      13'd4534: x = 8'h00;
      13'd4535: x = 8'h00;
      13'd4536: x = 8'h00;
      13'd4537: x = 8'h00;
      13'd4538: x = 8'h00;
      13'd4539: x = 8'h00;
      13'd4540: x = 8'h00;
      13'd4541: x = 8'h00;
      13'd4542: x = 8'h00;
      13'd4543: x = 8'h00;
      13'd4544: x = 8'h00;
      13'd4545: x = 8'h00;
      13'd4546: x = 8'h00;
      13'd4547: x = 8'h00;
      13'd4548: x = 8'h00;
      13'd4549: x = 8'h00;
      13'd4550: x = 8'h00;
      13'd4551: x = 8'h00;
      13'd4552: x = 8'h00;
      13'd4553: x = 8'h00;
      13'd4554: x = 8'h00;
      13'd4555: x = 8'h00;
      13'd4556: x = 8'h00;
      13'd4557: x = 8'h00;
      13'd4558: x = 8'h00;
      13'd4559: x = 8'h00;
      13'd4560: x = 8'h00;
      13'd4561: x = 8'h00;
      13'd4562: x = 8'h00;
      13'd4563: x = 8'h00;
      13'd4564: x = 8'h00;
      13'd4565: x = 8'h00;
      13'd4566: x = 8'h00;
      13'd4567: x = 8'h00;
      13'd4568: x = 8'h00;
      13'd4569: x = 8'h00;
      13'd4570: x = 8'h00;
      13'd4571: x = 8'h00;
      13'd4572: x = 8'h00;
      13'd4573: x = 8'h00;
      13'd4574: x = 8'h00;
      13'd4575: x = 8'h00;
      13'd4576: x = 8'h00;
      13'd4577: x = 8'h00;
      13'd4578: x = 8'h00;
      13'd4579: x = 8'h00;
      13'd4580: x = 8'h00;
      13'd4581: x = 8'h00;
      13'd4582: x = 8'h00;
      13'd4583: x = 8'h00;
      13'd4584: x = 8'h00;
      13'd4585: x = 8'h00;
      13'd4586: x = 8'h00;
      13'd4587: x = 8'h00;
      13'd4588: x = 8'h00;
      13'd4589: x = 8'h00;
      13'd4590: x = 8'h00;
      13'd4591: x = 8'h00;
      13'd4592: x = 8'h00;
      13'd4593: x = 8'h00;
      13'd4594: x = 8'h00;
      13'd4595: x = 8'h00;
      13'd4596: x = 8'h00;
      13'd4597: x = 8'h00;
      13'd4598: x = 8'h00;
      13'd4599: x = 8'h00;
      13'd4600: x = 8'h00;
      13'd4601: x = 8'h00;
      13'd4602: x = 8'h00;
      13'd4603: x = 8'h00;
      13'd4604: x = 8'h00;
      13'd4605: x = 8'h00;
      13'd4606: x = 8'h00;
      13'd4607: x = 8'h00;
      13'd4608: x = 8'h00;
      13'd4609: x = 8'h00;
      13'd4610: x = 8'h00;
      13'd4611: x = 8'h00;
      13'd4612: x = 8'h00;
      13'd4613: x = 8'h00;
      13'd4614: x = 8'h00;
      13'd4615: x = 8'h00;
      13'd4616: x = 8'h00;
      13'd4617: x = 8'h00;
      13'd4618: x = 8'h00;
      13'd4619: x = 8'h00;
      13'd4620: x = 8'h00;
      13'd4621: x = 8'h00;
      13'd4622: x = 8'h00;
      13'd4623: x = 8'h00;
      13'd4624: x = 8'h00;
      13'd4625: x = 8'h00;
      13'd4626: x = 8'h00;
      13'd4627: x = 8'h00;
      13'd4628: x = 8'h00;
      13'd4629: x = 8'h00;
      13'd4630: x = 8'h00;
      13'd4631: x = 8'h00;
      13'd4632: x = 8'h00;
      13'd4633: x = 8'h00;
      13'd4634: x = 8'h00;
      13'd4635: x = 8'h00;
      13'd4636: x = 8'h00;
      13'd4637: x = 8'h00;
      13'd4638: x = 8'h00;
      13'd4639: x = 8'h00;
      13'd4640: x = 8'h00;
      13'd4641: x = 8'h00;
      13'd4642: x = 8'h00;
      13'd4643: x = 8'h00;
      13'd4644: x = 8'h00;
      13'd4645: x = 8'h00;
      13'd4646: x = 8'h00;
      13'd4647: x = 8'h00;
      13'd4648: x = 8'h00;
      13'd4649: x = 8'h00;
      13'd4650: x = 8'h00;
      13'd4651: x = 8'h00;
      13'd4652: x = 8'h00;
      13'd4653: x = 8'h00;
      13'd4654: x = 8'h00;
      13'd4655: x = 8'h00;
      13'd4656: x = 8'h00;
      13'd4657: x = 8'h00;
      13'd4658: x = 8'h00;
      13'd4659: x = 8'h00;
      13'd4660: x = 8'h00;
      13'd4661: x = 8'h00;
      13'd4662: x = 8'h00;
      13'd4663: x = 8'h00;
      13'd4664: x = 8'h00;
      13'd4665: x = 8'h00;
      13'd4666: x = 8'h00;
      13'd4667: x = 8'h00;
      13'd4668: x = 8'h00;
      13'd4669: x = 8'h00;
      13'd4670: x = 8'h00;
      13'd4671: x = 8'h00;
      13'd4672: x = 8'h00;
      13'd4673: x = 8'h00;
      13'd4674: x = 8'h00;
      13'd4675: x = 8'h00;
      13'd4676: x = 8'h00;
      13'd4677: x = 8'h00;
      13'd4678: x = 8'h00;
      13'd4679: x = 8'h00;
      13'd4680: x = 8'h00;
      13'd4681: x = 8'h00;
      13'd4682: x = 8'h00;
      13'd4683: x = 8'h00;
      13'd4684: x = 8'h00;
      13'd4685: x = 8'h00;
      13'd4686: x = 8'h00;
      13'd4687: x = 8'h00;
      13'd4688: x = 8'h00;
      13'd4689: x = 8'h00;
      13'd4690: x = 8'h00;
      13'd4691: x = 8'h00;
      13'd4692: x = 8'h00;
      13'd4693: x = 8'h00;
      13'd4694: x = 8'h00;
      13'd4695: x = 8'h00;
      13'd4696: x = 8'h00;
      13'd4697: x = 8'h00;
      13'd4698: x = 8'h00;
      13'd4699: x = 8'h00;
      13'd4700: x = 8'h00;
      13'd4701: x = 8'h00;
      13'd4702: x = 8'h00;
      13'd4703: x = 8'h00;
      13'd4704: x = 8'h00;
      13'd4705: x = 8'h00;
      13'd4706: x = 8'h00;
      13'd4707: x = 8'h00;
      13'd4708: x = 8'h00;
      13'd4709: x = 8'h00;
      13'd4710: x = 8'h00;
      13'd4711: x = 8'h00;
      13'd4712: x = 8'h00;
      13'd4713: x = 8'h00;
      13'd4714: x = 8'h00;
      13'd4715: x = 8'h00;
      13'd4716: x = 8'h00;
      13'd4717: x = 8'h00;
      13'd4718: x = 8'h00;
      13'd4719: x = 8'h00;
      13'd4720: x = 8'h00;
      13'd4721: x = 8'h00;
      13'd4722: x = 8'h00;
      13'd4723: x = 8'h00;
      13'd4724: x = 8'h00;
      13'd4725: x = 8'h00;
      13'd4726: x = 8'h00;
      13'd4727: x = 8'h00;
      13'd4728: x = 8'h00;
      13'd4729: x = 8'h00;
      13'd4730: x = 8'h00;
      13'd4731: x = 8'h00;
      13'd4732: x = 8'h00;
      13'd4733: x = 8'h00;
      13'd4734: x = 8'h00;
      13'd4735: x = 8'h00;
      13'd4736: x = 8'h00;
      13'd4737: x = 8'h00;
      13'd4738: x = 8'h00;
      13'd4739: x = 8'h00;
      13'd4740: x = 8'h00;
      13'd4741: x = 8'h00;
      13'd4742: x = 8'h00;
      13'd4743: x = 8'h00;
      13'd4744: x = 8'h00;
      13'd4745: x = 8'h00;
      13'd4746: x = 8'h00;
      13'd4747: x = 8'h00;
      13'd4748: x = 8'h00;
      13'd4749: x = 8'h00;
      13'd4750: x = 8'h00;
      13'd4751: x = 8'h00;
      13'd4752: x = 8'h00;
      13'd4753: x = 8'h00;
      13'd4754: x = 8'h00;
      13'd4755: x = 8'h00;
      13'd4756: x = 8'h00;
      13'd4757: x = 8'h00;
      13'd4758: x = 8'h00;
      13'd4759: x = 8'h00;
      13'd4760: x = 8'h00;
      13'd4761: x = 8'h00;
      13'd4762: x = 8'h00;
      13'd4763: x = 8'h00;
      13'd4764: x = 8'h00;
      13'd4765: x = 8'h00;
      13'd4766: x = 8'h00;
      13'd4767: x = 8'h00;
      13'd4768: x = 8'h00;
      13'd4769: x = 8'h00;
      13'd4770: x = 8'h00;
      13'd4771: x = 8'h00;
      13'd4772: x = 8'h00;
      13'd4773: x = 8'h00;
      13'd4774: x = 8'h00;
      13'd4775: x = 8'h00;
      13'd4776: x = 8'h00;
      13'd4777: x = 8'h00;
      13'd4778: x = 8'h00;
      13'd4779: x = 8'h00;
      13'd4780: x = 8'h00;
      13'd4781: x = 8'h00;
      13'd4782: x = 8'h00;
      13'd4783: x = 8'h00;
      13'd4784: x = 8'h00;
      13'd4785: x = 8'h00;
      13'd4786: x = 8'h00;
      13'd4787: x = 8'h00;
      13'd4788: x = 8'h00;
      13'd4789: x = 8'h00;
      13'd4790: x = 8'h00;
      13'd4791: x = 8'h00;
      13'd4792: x = 8'h00;
      13'd4793: x = 8'h00;
      13'd4794: x = 8'h00;
      13'd4795: x = 8'h00;
      13'd4796: x = 8'h00;
      13'd4797: x = 8'h00;
      13'd4798: x = 8'h00;
      13'd4799: x = 8'h00;
      13'd4800: x = 8'h00;
      13'd4801: x = 8'h00;
      13'd4802: x = 8'h00;
      13'd4803: x = 8'h00;
      13'd4804: x = 8'h00;
      13'd4805: x = 8'h00;
      13'd4806: x = 8'h00;
      13'd4807: x = 8'h00;
      13'd4808: x = 8'h00;
      13'd4809: x = 8'h00;
      13'd4810: x = 8'h00;
      13'd4811: x = 8'h00;
      13'd4812: x = 8'h00;
      13'd4813: x = 8'h00;
      13'd4814: x = 8'h00;
      13'd4815: x = 8'h00;
      13'd4816: x = 8'h00;
      13'd4817: x = 8'h00;
      13'd4818: x = 8'h00;
      13'd4819: x = 8'h00;
      13'd4820: x = 8'h00;
      13'd4821: x = 8'h00;
      13'd4822: x = 8'h00;
      13'd4823: x = 8'h00;
      13'd4824: x = 8'h00;
      13'd4825: x = 8'h00;
      13'd4826: x = 8'h00;
      13'd4827: x = 8'h00;
      13'd4828: x = 8'h00;
      13'd4829: x = 8'h00;
      13'd4830: x = 8'h00;
      13'd4831: x = 8'h00;
      13'd4832: x = 8'h00;
      13'd4833: x = 8'h00;
      13'd4834: x = 8'h00;
      13'd4835: x = 8'h00;
      13'd4836: x = 8'h00;
      13'd4837: x = 8'h00;
      13'd4838: x = 8'h00;
      13'd4839: x = 8'h00;
      13'd4840: x = 8'h00;
      13'd4841: x = 8'h00;
      13'd4842: x = 8'h00;
      13'd4843: x = 8'h00;
      13'd4844: x = 8'h00;
      13'd4845: x = 8'h00;
      13'd4846: x = 8'h00;
      13'd4847: x = 8'h00;
      13'd4848: x = 8'h00;
      13'd4849: x = 8'h00;
      13'd4850: x = 8'h00;
      13'd4851: x = 8'h00;
      13'd4852: x = 8'h00;
      13'd4853: x = 8'h00;
      13'd4854: x = 8'h00;
      13'd4855: x = 8'h00;
      13'd4856: x = 8'h00;
      13'd4857: x = 8'h00;
      13'd4858: x = 8'h00;
      13'd4859: x = 8'h00;
      13'd4860: x = 8'h00;
      13'd4861: x = 8'h00;
      13'd4862: x = 8'h00;
      13'd4863: x = 8'h00;
      13'd4864: x = 8'h00;
      13'd4865: x = 8'h00;
      13'd4866: x = 8'h00;
      13'd4867: x = 8'h00;
      13'd4868: x = 8'h00;
      13'd4869: x = 8'h00;
      13'd4870: x = 8'h00;
      13'd4871: x = 8'h00;
      13'd4872: x = 8'h00;
      13'd4873: x = 8'h00;
      13'd4874: x = 8'h00;
      13'd4875: x = 8'h00;
      13'd4876: x = 8'h00;
      13'd4877: x = 8'h00;
      13'd4878: x = 8'h00;
      13'd4879: x = 8'h00;
      13'd4880: x = 8'h00;
      13'd4881: x = 8'h00;
      13'd4882: x = 8'h00;
      13'd4883: x = 8'h00;
      13'd4884: x = 8'h00;
      13'd4885: x = 8'h00;
      13'd4886: x = 8'h00;
      13'd4887: x = 8'h00;
      13'd4888: x = 8'h00;
      13'd4889: x = 8'h00;
      13'd4890: x = 8'h00;
      13'd4891: x = 8'h00;
      13'd4892: x = 8'h00;
      13'd4893: x = 8'h00;
      13'd4894: x = 8'h00;
      13'd4895: x = 8'h00;
      13'd4896: x = 8'h00;
      13'd4897: x = 8'h00;
      13'd4898: x = 8'h00;
      13'd4899: x = 8'h00;
      13'd4900: x = 8'h00;
      13'd4901: x = 8'h00;
      13'd4902: x = 8'h00;
      13'd4903: x = 8'h00;
      13'd4904: x = 8'h00;
      13'd4905: x = 8'h00;
      13'd4906: x = 8'h00;
      13'd4907: x = 8'h00;
      13'd4908: x = 8'h00;
      13'd4909: x = 8'h00;
      13'd4910: x = 8'h00;
      13'd4911: x = 8'h00;
      13'd4912: x = 8'h00;
      13'd4913: x = 8'h00;
      13'd4914: x = 8'h00;
      13'd4915: x = 8'h00;
      13'd4916: x = 8'h00;
      13'd4917: x = 8'h00;
      13'd4918: x = 8'h00;
      13'd4919: x = 8'h00;
      13'd4920: x = 8'h00;
      13'd4921: x = 8'h00;
      13'd4922: x = 8'h00;
      13'd4923: x = 8'h00;
      13'd4924: x = 8'h00;
      13'd4925: x = 8'h00;
      13'd4926: x = 8'h00;
      13'd4927: x = 8'h00;
      13'd4928: x = 8'h00;
      13'd4929: x = 8'h00;
      13'd4930: x = 8'h00;
      13'd4931: x = 8'h00;
      13'd4932: x = 8'h00;
      13'd4933: x = 8'h00;
      13'd4934: x = 8'h00;
      13'd4935: x = 8'h00;
      13'd4936: x = 8'h00;
      13'd4937: x = 8'h00;
      13'd4938: x = 8'h00;
      13'd4939: x = 8'h00;
      13'd4940: x = 8'h00;
      13'd4941: x = 8'h00;
      13'd4942: x = 8'h00;
      13'd4943: x = 8'h00;
      13'd4944: x = 8'h00;
      13'd4945: x = 8'h00;
      13'd4946: x = 8'h00;
      13'd4947: x = 8'h00;
      13'd4948: x = 8'h00;
      13'd4949: x = 8'h00;
      13'd4950: x = 8'h00;
      13'd4951: x = 8'h00;
      13'd4952: x = 8'h00;
      13'd4953: x = 8'h00;
      13'd4954: x = 8'h00;
      13'd4955: x = 8'h00;
      13'd4956: x = 8'h00;
      13'd4957: x = 8'h00;
      13'd4958: x = 8'h00;
      13'd4959: x = 8'h00;
      13'd4960: x = 8'h00;
      13'd4961: x = 8'h00;
      13'd4962: x = 8'h00;
      13'd4963: x = 8'h00;
      13'd4964: x = 8'h00;
      13'd4965: x = 8'h00;
      13'd4966: x = 8'h00;
      13'd4967: x = 8'h00;
      13'd4968: x = 8'h00;
      13'd4969: x = 8'h00;
      13'd4970: x = 8'h00;
      13'd4971: x = 8'h00;
      13'd4972: x = 8'h00;
      13'd4973: x = 8'h00;
      13'd4974: x = 8'h00;
      13'd4975: x = 8'h00;
      13'd4976: x = 8'h00;
      13'd4977: x = 8'h00;
      13'd4978: x = 8'h00;
      13'd4979: x = 8'h00;
      13'd4980: x = 8'h00;
      13'd4981: x = 8'h00;
      13'd4982: x = 8'h00;
      13'd4983: x = 8'h00;
      13'd4984: x = 8'h00;
      13'd4985: x = 8'h00;
      13'd4986: x = 8'h00;
      13'd4987: x = 8'h00;
      13'd4988: x = 8'h00;
      13'd4989: x = 8'h00;
      13'd4990: x = 8'h00;
      13'd4991: x = 8'h00;
      13'd4992: x = 8'h00;
      13'd4993: x = 8'h00;
      13'd4994: x = 8'h00;
      13'd4995: x = 8'h00;
      13'd4996: x = 8'h00;
      13'd4997: x = 8'h00;
      13'd4998: x = 8'h00;
      13'd4999: x = 8'h00;
      13'd5000: x = 8'h00;
      13'd5001: x = 8'h00;
      13'd5002: x = 8'h00;
      13'd5003: x = 8'h00;
      13'd5004: x = 8'h00;
      13'd5005: x = 8'h00;
      13'd5006: x = 8'h00;
      13'd5007: x = 8'h00;
      13'd5008: x = 8'h00;
      13'd5009: x = 8'h00;
      13'd5010: x = 8'h00;
      13'd5011: x = 8'h00;
      13'd5012: x = 8'h00;
      13'd5013: x = 8'h00;
      13'd5014: x = 8'h00;
      13'd5015: x = 8'h00;
      13'd5016: x = 8'h00;
      13'd5017: x = 8'h00;
      13'd5018: x = 8'h00;
      13'd5019: x = 8'h00;
      13'd5020: x = 8'h00;
      13'd5021: x = 8'h00;
      13'd5022: x = 8'h00;
      13'd5023: x = 8'h00;
      13'd5024: x = 8'h00;
      13'd5025: x = 8'h00;
      13'd5026: x = 8'h00;
      13'd5027: x = 8'h00;
      13'd5028: x = 8'h00;
      13'd5029: x = 8'h00;
      13'd5030: x = 8'h00;
      13'd5031: x = 8'h00;
      13'd5032: x = 8'h00;
      13'd5033: x = 8'h00;
      13'd5034: x = 8'h00;
      13'd5035: x = 8'h00;
      13'd5036: x = 8'h00;
      13'd5037: x = 8'h00;
      13'd5038: x = 8'h00;
      13'd5039: x = 8'h00;
      13'd5040: x = 8'h00;
      13'd5041: x = 8'h00;
      13'd5042: x = 8'h00;
      13'd5043: x = 8'h00;
      13'd5044: x = 8'h00;
      13'd5045: x = 8'h00;
      13'd5046: x = 8'h00;
      13'd5047: x = 8'h00;
      13'd5048: x = 8'h00;
      13'd5049: x = 8'h00;
      13'd5050: x = 8'h00;
      13'd5051: x = 8'h00;
      13'd5052: x = 8'h00;
      13'd5053: x = 8'h00;
      13'd5054: x = 8'h00;
      13'd5055: x = 8'h00;
      13'd5056: x = 8'h00;
      13'd5057: x = 8'h00;
      13'd5058: x = 8'h00;
      13'd5059: x = 8'h00;
      13'd5060: x = 8'h00;
      13'd5061: x = 8'h00;
      13'd5062: x = 8'h00;
      13'd5063: x = 8'h00;
      13'd5064: x = 8'h00;
      13'd5065: x = 8'h00;
      13'd5066: x = 8'h00;
      13'd5067: x = 8'h00;
      13'd5068: x = 8'h00;
      13'd5069: x = 8'h00;
      13'd5070: x = 8'h00;
      13'd5071: x = 8'h00;
      13'd5072: x = 8'h00;
      13'd5073: x = 8'h00;
      13'd5074: x = 8'h00;
      13'd5075: x = 8'h00;
      13'd5076: x = 8'h00;
      13'd5077: x = 8'h00;
      13'd5078: x = 8'h00;
      13'd5079: x = 8'h00;
      13'd5080: x = 8'h00;
      13'd5081: x = 8'h00;
      13'd5082: x = 8'h00;
      13'd5083: x = 8'h00;
      13'd5084: x = 8'h00;
      13'd5085: x = 8'h00;
      13'd5086: x = 8'h00;
      13'd5087: x = 8'h00;
      13'd5088: x = 8'h00;
      13'd5089: x = 8'h00;
      13'd5090: x = 8'h00;
      13'd5091: x = 8'h00;
      13'd5092: x = 8'h00;
      13'd5093: x = 8'h00;
      13'd5094: x = 8'h00;
      13'd5095: x = 8'h00;
      13'd5096: x = 8'h00;
      13'd5097: x = 8'h00;
      13'd5098: x = 8'h00;
      13'd5099: x = 8'h00;
      13'd5100: x = 8'h00;
      13'd5101: x = 8'h00;
      13'd5102: x = 8'h00;
      13'd5103: x = 8'h00;
      13'd5104: x = 8'h00;
      13'd5105: x = 8'h00;
      13'd5106: x = 8'h00;
      13'd5107: x = 8'h00;
      13'd5108: x = 8'h00;
      13'd5109: x = 8'h00;
      13'd5110: x = 8'h00;
      13'd5111: x = 8'h00;
      13'd5112: x = 8'h00;
      13'd5113: x = 8'h00;
      13'd5114: x = 8'h00;
      13'd5115: x = 8'h00;
      13'd5116: x = 8'h00;
      13'd5117: x = 8'h00;
      13'd5118: x = 8'h00;
      13'd5119: x = 8'h00;
      13'd5120: x = 8'h00;
      13'd5121: x = 8'h00;
      13'd5122: x = 8'h00;
      13'd5123: x = 8'h00;
      13'd5124: x = 8'h00;
      13'd5125: x = 8'h00;
      13'd5126: x = 8'h00;
      13'd5127: x = 8'h00;
      13'd5128: x = 8'h00;
      13'd5129: x = 8'h00;
      13'd5130: x = 8'h00;
      13'd5131: x = 8'h00;
      13'd5132: x = 8'h00;
      13'd5133: x = 8'h00;
      13'd5134: x = 8'h00;
      13'd5135: x = 8'h00;
      13'd5136: x = 8'h00;
      13'd5137: x = 8'h00;
      13'd5138: x = 8'h00;
      13'd5139: x = 8'h00;
      13'd5140: x = 8'h00;
      13'd5141: x = 8'h00;
      13'd5142: x = 8'h00;
      13'd5143: x = 8'h00;
      13'd5144: x = 8'h00;
      13'd5145: x = 8'h00;
      13'd5146: x = 8'h00;
      13'd5147: x = 8'h00;
      13'd5148: x = 8'h00;
      13'd5149: x = 8'h00;
      13'd5150: x = 8'h00;
      13'd5151: x = 8'h00;
      13'd5152: x = 8'h00;
      13'd5153: x = 8'h00;
      13'd5154: x = 8'h00;
      13'd5155: x = 8'h00;
      13'd5156: x = 8'h00;
      13'd5157: x = 8'h00;
      13'd5158: x = 8'h00;
      13'd5159: x = 8'h00;
      13'd5160: x = 8'h00;
      13'd5161: x = 8'h00;
      13'd5162: x = 8'h00;
      13'd5163: x = 8'h00;
      13'd5164: x = 8'h00;
      13'd5165: x = 8'h00;
      13'd5166: x = 8'h00;
      13'd5167: x = 8'h00;
      13'd5168: x = 8'h00;
      13'd5169: x = 8'h00;
      13'd5170: x = 8'h00;
      13'd5171: x = 8'h00;
      13'd5172: x = 8'h00;
      13'd5173: x = 8'h00;
      13'd5174: x = 8'h00;
      13'd5175: x = 8'h00;
      13'd5176: x = 8'h00;
      13'd5177: x = 8'h00;
      13'd5178: x = 8'h00;
      13'd5179: x = 8'h00;
      13'd5180: x = 8'h00;
      13'd5181: x = 8'h00;
      13'd5182: x = 8'h00;
      13'd5183: x = 8'h00;
      13'd5184: x = 8'h00;
      13'd5185: x = 8'h00;
      13'd5186: x = 8'h00;
      13'd5187: x = 8'h00;
      13'd5188: x = 8'h00;
      13'd5189: x = 8'h00;
      13'd5190: x = 8'h00;
      13'd5191: x = 8'h00;
      13'd5192: x = 8'h00;
      13'd5193: x = 8'h00;
      13'd5194: x = 8'h00;
      13'd5195: x = 8'h00;
      13'd5196: x = 8'h00;
      13'd5197: x = 8'h00;
      13'd5198: x = 8'h00;
      13'd5199: x = 8'h00;
      13'd5200: x = 8'h00;
      13'd5201: x = 8'h00;
      13'd5202: x = 8'h00;
      13'd5203: x = 8'h00;
      13'd5204: x = 8'h00;
      13'd5205: x = 8'h00;
      13'd5206: x = 8'h00;
      13'd5207: x = 8'h00;
      13'd5208: x = 8'h00;
      13'd5209: x = 8'h00;
      13'd5210: x = 8'h00;
      13'd5211: x = 8'h00;
      13'd5212: x = 8'h00;
      13'd5213: x = 8'h00;
      13'd5214: x = 8'h00;
      13'd5215: x = 8'h00;
      13'd5216: x = 8'h00;
      13'd5217: x = 8'h00;
      13'd5218: x = 8'h00;
      13'd5219: x = 8'h00;
      13'd5220: x = 8'h00;
      13'd5221: x = 8'h00;
      13'd5222: x = 8'h00;
      13'd5223: x = 8'h00;
      13'd5224: x = 8'h00;
      13'd5225: x = 8'h00;
      13'd5226: x = 8'h00;
      13'd5227: x = 8'h00;
      13'd5228: x = 8'h00;
      13'd5229: x = 8'h00;
      13'd5230: x = 8'h00;
      13'd5231: x = 8'h00;
      13'd5232: x = 8'h00;
      13'd5233: x = 8'h00;
      13'd5234: x = 8'h00;
      13'd5235: x = 8'h00;
      13'd5236: x = 8'h00;
      13'd5237: x = 8'h00;
      13'd5238: x = 8'h00;
      13'd5239: x = 8'h00;
      13'd5240: x = 8'h00;
      13'd5241: x = 8'h00;
      13'd5242: x = 8'h00;
      13'd5243: x = 8'h00;
      13'd5244: x = 8'h00;
      13'd5245: x = 8'h00;
      13'd5246: x = 8'h00;
      13'd5247: x = 8'h00;
      13'd5248: x = 8'h00;
      13'd5249: x = 8'h00;
      13'd5250: x = 8'h00;
      13'd5251: x = 8'h00;
      13'd5252: x = 8'h00;
      13'd5253: x = 8'h00;
      13'd5254: x = 8'h00;
      13'd5255: x = 8'h00;
      13'd5256: x = 8'h00;
      13'd5257: x = 8'h00;
      13'd5258: x = 8'h00;
      13'd5259: x = 8'h00;
      13'd5260: x = 8'h00;
      13'd5261: x = 8'h00;
      13'd5262: x = 8'h00;
      13'd5263: x = 8'h00;
      13'd5264: x = 8'h00;
      13'd5265: x = 8'h00;
      13'd5266: x = 8'h00;
      13'd5267: x = 8'h00;
      13'd5268: x = 8'h00;
      13'd5269: x = 8'h00;
      13'd5270: x = 8'h00;
      13'd5271: x = 8'h00;
      13'd5272: x = 8'h00;
      13'd5273: x = 8'h00;
      13'd5274: x = 8'h00;
      13'd5275: x = 8'h00;
      13'd5276: x = 8'h00;
      13'd5277: x = 8'h00;
      13'd5278: x = 8'h00;
      13'd5279: x = 8'h00;
      13'd5280: x = 8'h00;
      13'd5281: x = 8'h00;
      13'd5282: x = 8'h00;
      13'd5283: x = 8'h00;
      13'd5284: x = 8'h00;
      13'd5285: x = 8'h00;
      13'd5286: x = 8'h00;
      13'd5287: x = 8'h00;
      13'd5288: x = 8'h00;
      13'd5289: x = 8'h00;
      13'd5290: x = 8'h00;
      13'd5291: x = 8'h00;
      13'd5292: x = 8'h00;
      13'd5293: x = 8'h00;
      13'd5294: x = 8'h00;
      13'd5295: x = 8'h00;
      13'd5296: x = 8'h00;
      13'd5297: x = 8'h00;
      13'd5298: x = 8'h00;
      13'd5299: x = 8'h00;
      13'd5300: x = 8'h00;
      13'd5301: x = 8'h00;
      13'd5302: x = 8'h00;
      13'd5303: x = 8'h00;
      13'd5304: x = 8'h00;
      13'd5305: x = 8'h00;
      13'd5306: x = 8'h00;
      13'd5307: x = 8'h00;
      13'd5308: x = 8'h00;
      13'd5309: x = 8'h00;
      13'd5310: x = 8'h00;
      13'd5311: x = 8'h00;
      13'd5312: x = 8'h00;
      13'd5313: x = 8'h00;
      13'd5314: x = 8'h00;
      13'd5315: x = 8'h00;
      13'd5316: x = 8'h00;
      13'd5317: x = 8'h00;
      13'd5318: x = 8'h00;
      13'd5319: x = 8'h00;
      13'd5320: x = 8'h00;
      13'd5321: x = 8'h00;
      13'd5322: x = 8'h00;
      13'd5323: x = 8'h00;
      13'd5324: x = 8'h00;
      13'd5325: x = 8'h00;
      13'd5326: x = 8'h00;
      13'd5327: x = 8'h00;
      13'd5328: x = 8'h00;
      13'd5329: x = 8'h00;
      13'd5330: x = 8'h00;
      13'd5331: x = 8'h00;
      13'd5332: x = 8'h00;
      13'd5333: x = 8'h00;
      13'd5334: x = 8'h00;
      13'd5335: x = 8'h00;
      13'd5336: x = 8'h00;
      13'd5337: x = 8'h00;
      13'd5338: x = 8'h00;
      13'd5339: x = 8'h00;
      13'd5340: x = 8'h00;
      13'd5341: x = 8'h00;
      13'd5342: x = 8'h00;
      13'd5343: x = 8'h00;
      13'd5344: x = 8'h00;
      13'd5345: x = 8'h00;
      13'd5346: x = 8'h00;
      13'd5347: x = 8'h00;
      13'd5348: x = 8'h00;
      13'd5349: x = 8'h00;
      13'd5350: x = 8'h00;
      13'd5351: x = 8'h00;
      13'd5352: x = 8'h00;
      13'd5353: x = 8'h00;
      13'd5354: x = 8'h00;
      13'd5355: x = 8'h00;
      13'd5356: x = 8'h00;
      13'd5357: x = 8'h00;
      13'd5358: x = 8'h00;
      13'd5359: x = 8'h00;
      13'd5360: x = 8'h00;
      13'd5361: x = 8'h00;
      13'd5362: x = 8'h00;
      13'd5363: x = 8'h00;
      13'd5364: x = 8'h00;
      13'd5365: x = 8'h00;
      13'd5366: x = 8'h00;
      13'd5367: x = 8'h00;
      13'd5368: x = 8'h00;
      13'd5369: x = 8'h00;
      13'd5370: x = 8'h00;
      13'd5371: x = 8'h00;
      13'd5372: x = 8'h00;
      13'd5373: x = 8'h00;
      13'd5374: x = 8'h00;
      13'd5375: x = 8'h00;
      13'd5376: x = 8'h00;
      13'd5377: x = 8'h00;
      13'd5378: x = 8'h00;
      13'd5379: x = 8'h00;
      13'd5380: x = 8'h00;
      13'd5381: x = 8'h00;
      13'd5382: x = 8'h00;
      13'd5383: x = 8'h00;
      13'd5384: x = 8'h00;
      13'd5385: x = 8'h00;
      13'd5386: x = 8'h00;
      13'd5387: x = 8'h00;
      13'd5388: x = 8'h00;
      13'd5389: x = 8'h00;
      13'd5390: x = 8'h00;
      13'd5391: x = 8'h00;
      13'd5392: x = 8'h00;
      13'd5393: x = 8'h00;
      13'd5394: x = 8'h00;
      13'd5395: x = 8'h00;
      13'd5396: x = 8'h00;
      13'd5397: x = 8'h00;
      13'd5398: x = 8'h00;
      13'd5399: x = 8'h00;
      13'd5400: x = 8'h00;
      13'd5401: x = 8'h00;
      13'd5402: x = 8'h00;
      13'd5403: x = 8'h00;
      13'd5404: x = 8'h00;
      13'd5405: x = 8'h00;
      13'd5406: x = 8'h00;
      13'd5407: x = 8'h00;
      13'd5408: x = 8'h00;
      13'd5409: x = 8'h00;
      13'd5410: x = 8'h00;
      13'd5411: x = 8'h00;
      13'd5412: x = 8'h00;
      13'd5413: x = 8'h00;
      13'd5414: x = 8'h00;
      13'd5415: x = 8'h00;
      13'd5416: x = 8'h00;
      13'd5417: x = 8'h00;
      13'd5418: x = 8'h00;
      13'd5419: x = 8'h00;
      13'd5420: x = 8'h00;
      13'd5421: x = 8'h00;
      13'd5422: x = 8'h00;
      13'd5423: x = 8'h00;
      13'd5424: x = 8'h00;
      13'd5425: x = 8'h00;
      13'd5426: x = 8'h00;
      13'd5427: x = 8'h00;
      13'd5428: x = 8'h00;
      13'd5429: x = 8'h00;
      13'd5430: x = 8'h00;
      13'd5431: x = 8'h00;
      13'd5432: x = 8'h00;
      13'd5433: x = 8'h00;
      13'd5434: x = 8'h00;
      13'd5435: x = 8'h00;
      13'd5436: x = 8'h00;
      13'd5437: x = 8'h00;
      13'd5438: x = 8'h00;
      13'd5439: x = 8'h00;
      13'd5440: x = 8'h00;
      13'd5441: x = 8'h00;
      13'd5442: x = 8'h00;
      13'd5443: x = 8'h00;
      13'd5444: x = 8'h00;
      13'd5445: x = 8'h00;
      13'd5446: x = 8'h00;
      13'd5447: x = 8'h00;
      13'd5448: x = 8'h00;
      13'd5449: x = 8'h00;
      13'd5450: x = 8'h00;
      13'd5451: x = 8'h00;
      13'd5452: x = 8'h00;
      13'd5453: x = 8'h00;
      13'd5454: x = 8'h00;
      13'd5455: x = 8'h00;
      13'd5456: x = 8'h00;
      13'd5457: x = 8'h00;
      13'd5458: x = 8'h00;
      13'd5459: x = 8'h00;
      13'd5460: x = 8'h00;
      13'd5461: x = 8'h00;
      13'd5462: x = 8'h00;
      13'd5463: x = 8'h00;
      13'd5464: x = 8'h00;
      13'd5465: x = 8'h00;
      13'd5466: x = 8'h00;
      13'd5467: x = 8'h00;
      13'd5468: x = 8'h00;
      13'd5469: x = 8'h00;
      13'd5470: x = 8'h00;
      13'd5471: x = 8'h00;
      13'd5472: x = 8'h00;
      13'd5473: x = 8'h00;
      13'd5474: x = 8'h00;
      13'd5475: x = 8'h00;
      13'd5476: x = 8'h00;
      13'd5477: x = 8'h00;
      13'd5478: x = 8'h00;
      13'd5479: x = 8'h00;
      13'd5480: x = 8'h00;
      13'd5481: x = 8'h00;
      13'd5482: x = 8'h00;
      13'd5483: x = 8'h00;
      13'd5484: x = 8'h00;
      13'd5485: x = 8'h00;
      13'd5486: x = 8'h00;
      13'd5487: x = 8'h00;
      13'd5488: x = 8'h00;
      13'd5489: x = 8'h00;
      13'd5490: x = 8'h00;
      13'd5491: x = 8'h00;
      13'd5492: x = 8'h00;
      13'd5493: x = 8'h00;
      13'd5494: x = 8'h00;
      13'd5495: x = 8'h00;
      13'd5496: x = 8'h00;
      13'd5497: x = 8'h00;
      13'd5498: x = 8'h00;
      13'd5499: x = 8'h00;
      13'd5500: x = 8'h00;
      13'd5501: x = 8'h00;
      13'd5502: x = 8'h00;
      13'd5503: x = 8'h00;
      13'd5504: x = 8'h00;
      13'd5505: x = 8'h00;
      13'd5506: x = 8'h00;
      13'd5507: x = 8'h00;
      13'd5508: x = 8'h00;
      13'd5509: x = 8'h00;
      13'd5510: x = 8'h00;
      13'd5511: x = 8'h00;
      13'd5512: x = 8'h00;
      13'd5513: x = 8'h00;
      13'd5514: x = 8'h00;
      13'd5515: x = 8'h00;
      13'd5516: x = 8'h00;
      13'd5517: x = 8'h00;
      13'd5518: x = 8'h00;
      13'd5519: x = 8'h00;
      13'd5520: x = 8'h00;
      13'd5521: x = 8'h00;
      13'd5522: x = 8'h00;
      13'd5523: x = 8'h00;
      13'd5524: x = 8'h00;
      13'd5525: x = 8'h00;
      13'd5526: x = 8'h00;
      13'd5527: x = 8'h00;
      13'd5528: x = 8'h00;
      13'd5529: x = 8'h00;
      13'd5530: x = 8'h00;
      13'd5531: x = 8'h00;
      13'd5532: x = 8'h00;
      13'd5533: x = 8'h00;
      13'd5534: x = 8'h00;
      13'd5535: x = 8'h00;
      13'd5536: x = 8'h00;
      13'd5537: x = 8'h00;
      13'd5538: x = 8'h00;
      13'd5539: x = 8'h00;
      13'd5540: x = 8'h00;
      13'd5541: x = 8'h00;
      13'd5542: x = 8'h00;
      13'd5543: x = 8'h00;
      13'd5544: x = 8'h00;
      13'd5545: x = 8'h00;
      13'd5546: x = 8'h00;
      13'd5547: x = 8'h00;
      13'd5548: x = 8'h00;
      13'd5549: x = 8'h00;
      13'd5550: x = 8'h00;
      13'd5551: x = 8'h00;
      13'd5552: x = 8'h00;
      13'd5553: x = 8'h00;
      13'd5554: x = 8'h00;
      13'd5555: x = 8'h00;
      13'd5556: x = 8'h00;
      13'd5557: x = 8'h00;
      13'd5558: x = 8'h00;
      13'd5559: x = 8'h00;
      13'd5560: x = 8'h00;
      13'd5561: x = 8'h00;
      13'd5562: x = 8'h00;
      13'd5563: x = 8'h00;
      13'd5564: x = 8'h00;
      13'd5565: x = 8'h00;
      13'd5566: x = 8'h00;
      13'd5567: x = 8'h00;
      13'd5568: x = 8'h00;
      13'd5569: x = 8'h00;
      13'd5570: x = 8'h00;
      13'd5571: x = 8'h00;
      13'd5572: x = 8'h00;
      13'd5573: x = 8'h00;
      13'd5574: x = 8'h00;
      13'd5575: x = 8'h00;
      13'd5576: x = 8'h00;
      13'd5577: x = 8'h00;
      13'd5578: x = 8'h00;
      13'd5579: x = 8'h00;
      13'd5580: x = 8'h00;
      13'd5581: x = 8'h00;
      13'd5582: x = 8'h00;
      13'd5583: x = 8'h00;
      13'd5584: x = 8'h00;
      13'd5585: x = 8'h00;
      13'd5586: x = 8'h00;
      13'd5587: x = 8'h00;
      13'd5588: x = 8'h00;
      13'd5589: x = 8'h00;
      13'd5590: x = 8'h00;
      13'd5591: x = 8'h00;
      13'd5592: x = 8'h00;
      13'd5593: x = 8'h00;
      13'd5594: x = 8'h00;
      13'd5595: x = 8'h00;
      13'd5596: x = 8'h00;
      13'd5597: x = 8'h00;
      13'd5598: x = 8'h00;
      13'd5599: x = 8'h00;
      13'd5600: x = 8'h00;
      13'd5601: x = 8'h00;
      13'd5602: x = 8'h00;
      13'd5603: x = 8'h00;
      13'd5604: x = 8'h00;
      13'd5605: x = 8'h00;
      13'd5606: x = 8'h00;
      13'd5607: x = 8'h00;
      13'd5608: x = 8'h00;
      13'd5609: x = 8'h00;
      13'd5610: x = 8'h00;
      13'd5611: x = 8'h00;
      13'd5612: x = 8'h00;
      13'd5613: x = 8'h00;
      13'd5614: x = 8'h00;
      13'd5615: x = 8'h00;
      13'd5616: x = 8'h00;
      13'd5617: x = 8'h00;
      13'd5618: x = 8'h00;
      13'd5619: x = 8'h00;
      13'd5620: x = 8'h00;
      13'd5621: x = 8'h00;
      13'd5622: x = 8'h00;
      13'd5623: x = 8'h00;
      13'd5624: x = 8'h00;
      13'd5625: x = 8'h00;
      13'd5626: x = 8'h00;
      13'd5627: x = 8'h00;
      13'd5628: x = 8'h00;
      13'd5629: x = 8'h00;
      13'd5630: x = 8'h00;
      13'd5631: x = 8'h00;
      13'd5632: x = 8'h00;
      13'd5633: x = 8'h00;
      13'd5634: x = 8'h00;
      13'd5635: x = 8'h00;
      13'd5636: x = 8'h00;
      13'd5637: x = 8'h00;
      13'd5638: x = 8'h00;
      13'd5639: x = 8'h00;
      13'd5640: x = 8'h00;
      13'd5641: x = 8'h00;
      13'd5642: x = 8'h00;
      13'd5643: x = 8'h00;
      13'd5644: x = 8'h00;
      13'd5645: x = 8'h00;
      13'd5646: x = 8'h00;
      13'd5647: x = 8'h00;
      13'd5648: x = 8'h00;
      13'd5649: x = 8'h00;
      13'd5650: x = 8'h00;
      13'd5651: x = 8'h00;
      13'd5652: x = 8'h00;
      13'd5653: x = 8'h00;
      13'd5654: x = 8'h00;
      13'd5655: x = 8'h00;
      13'd5656: x = 8'h00;
      13'd5657: x = 8'h00;
      13'd5658: x = 8'h00;
      13'd5659: x = 8'h00;
      13'd5660: x = 8'h00;
      13'd5661: x = 8'h00;
      13'd5662: x = 8'h00;
      13'd5663: x = 8'h00;
      13'd5664: x = 8'h00;
      13'd5665: x = 8'h00;
      13'd5666: x = 8'h00;
      13'd5667: x = 8'h00;
      13'd5668: x = 8'h00;
      13'd5669: x = 8'h00;
      13'd5670: x = 8'h00;
      13'd5671: x = 8'h00;
      13'd5672: x = 8'h00;
      13'd5673: x = 8'h00;
      13'd5674: x = 8'h00;
      13'd5675: x = 8'h00;
      13'd5676: x = 8'h00;
      13'd5677: x = 8'h00;
      13'd5678: x = 8'h00;
      13'd5679: x = 8'h00;
      13'd5680: x = 8'h00;
      13'd5681: x = 8'h00;
      13'd5682: x = 8'h00;
      13'd5683: x = 8'h00;
      13'd5684: x = 8'h00;
      13'd5685: x = 8'h00;
      13'd5686: x = 8'h00;
      13'd5687: x = 8'h00;
      13'd5688: x = 8'h00;
      13'd5689: x = 8'h00;
      13'd5690: x = 8'h00;
      13'd5691: x = 8'h00;
      13'd5692: x = 8'h00;
      13'd5693: x = 8'h00;
      13'd5694: x = 8'h00;
      13'd5695: x = 8'h00;
      13'd5696: x = 8'h00;
      13'd5697: x = 8'h00;
      13'd5698: x = 8'h00;
      13'd5699: x = 8'h00;
      13'd5700: x = 8'h00;
      13'd5701: x = 8'h00;
      13'd5702: x = 8'h00;
      13'd5703: x = 8'h00;
      13'd5704: x = 8'h00;
      13'd5705: x = 8'h00;
      13'd5706: x = 8'h00;
      13'd5707: x = 8'h00;
      13'd5708: x = 8'h00;
      13'd5709: x = 8'h00;
      13'd5710: x = 8'h00;
      13'd5711: x = 8'h00;
      13'd5712: x = 8'h00;
      13'd5713: x = 8'h00;
      13'd5714: x = 8'h00;
      13'd5715: x = 8'h00;
      13'd5716: x = 8'h00;
      13'd5717: x = 8'h00;
      13'd5718: x = 8'h00;
      13'd5719: x = 8'h00;
      13'd5720: x = 8'h00;
      13'd5721: x = 8'h00;
      13'd5722: x = 8'h00;
      13'd5723: x = 8'h00;
      13'd5724: x = 8'h00;
      13'd5725: x = 8'h00;
      13'd5726: x = 8'h00;
      13'd5727: x = 8'h00;
      13'd5728: x = 8'h00;
      13'd5729: x = 8'h00;
      13'd5730: x = 8'h00;
      13'd5731: x = 8'h00;
      13'd5732: x = 8'h00;
      13'd5733: x = 8'h00;
      13'd5734: x = 8'h00;
      13'd5735: x = 8'h00;
      13'd5736: x = 8'h00;
      13'd5737: x = 8'h00;
      13'd5738: x = 8'h00;
      13'd5739: x = 8'h00;
      13'd5740: x = 8'h00;
      13'd5741: x = 8'h00;
      13'd5742: x = 8'h00;
      13'd5743: x = 8'h00;
      13'd5744: x = 8'h00;
      13'd5745: x = 8'h00;
      13'd5746: x = 8'h00;
      13'd5747: x = 8'h00;
      13'd5748: x = 8'h00;
      13'd5749: x = 8'h00;
      13'd5750: x = 8'h00;
      13'd5751: x = 8'h00;
      13'd5752: x = 8'h00;
      13'd5753: x = 8'h00;
      13'd5754: x = 8'h00;
      13'd5755: x = 8'h00;
      13'd5756: x = 8'h00;
      13'd5757: x = 8'h00;
      13'd5758: x = 8'h00;
      13'd5759: x = 8'h00;
      13'd5760: x = 8'h00;
      13'd5761: x = 8'h00;
      13'd5762: x = 8'h00;
      13'd5763: x = 8'h00;
      13'd5764: x = 8'h00;
      13'd5765: x = 8'h00;
      13'd5766: x = 8'h00;
      13'd5767: x = 8'h00;
      13'd5768: x = 8'h00;
      13'd5769: x = 8'h00;
      13'd5770: x = 8'h00;
      13'd5771: x = 8'h00;
      13'd5772: x = 8'h00;
      13'd5773: x = 8'h00;
      13'd5774: x = 8'h00;
      13'd5775: x = 8'h00;
      13'd5776: x = 8'h00;
      13'd5777: x = 8'h00;
      13'd5778: x = 8'h00;
      13'd5779: x = 8'h00;
      13'd5780: x = 8'h00;
      13'd5781: x = 8'h00;
      13'd5782: x = 8'h00;
      13'd5783: x = 8'h00;
      13'd5784: x = 8'h00;
      13'd5785: x = 8'h00;
      13'd5786: x = 8'h00;
      13'd5787: x = 8'h00;
      13'd5788: x = 8'h00;
      13'd5789: x = 8'h00;
      13'd5790: x = 8'h00;
      13'd5791: x = 8'h00;
      13'd5792: x = 8'h00;
      13'd5793: x = 8'h00;
      13'd5794: x = 8'h00;
      13'd5795: x = 8'h00;
      13'd5796: x = 8'h00;
      13'd5797: x = 8'h00;
      13'd5798: x = 8'h00;
      13'd5799: x = 8'h00;
      13'd5800: x = 8'h00;
      13'd5801: x = 8'h00;
      13'd5802: x = 8'h00;
      13'd5803: x = 8'h00;
      13'd5804: x = 8'h00;
      13'd5805: x = 8'h00;
      13'd5806: x = 8'h00;
      13'd5807: x = 8'h00;
      13'd5808: x = 8'h00;
      13'd5809: x = 8'h00;
      13'd5810: x = 8'h00;
      13'd5811: x = 8'h00;
      13'd5812: x = 8'h00;
      13'd5813: x = 8'h00;
      13'd5814: x = 8'h00;
      13'd5815: x = 8'h00;
      13'd5816: x = 8'h00;
      13'd5817: x = 8'h00;
      13'd5818: x = 8'h00;
      13'd5819: x = 8'h00;
      13'd5820: x = 8'h00;
      13'd5821: x = 8'h00;
      13'd5822: x = 8'h00;
      13'd5823: x = 8'h00;
      13'd5824: x = 8'h00;
      13'd5825: x = 8'h00;
      13'd5826: x = 8'h00;
      13'd5827: x = 8'h00;
      13'd5828: x = 8'h00;
      13'd5829: x = 8'h00;
      13'd5830: x = 8'h00;
      13'd5831: x = 8'h00;
      13'd5832: x = 8'h00;
      13'd5833: x = 8'h00;
      13'd5834: x = 8'h00;
      13'd5835: x = 8'h00;
      13'd5836: x = 8'h00;
      13'd5837: x = 8'h00;
      13'd5838: x = 8'h00;
      13'd5839: x = 8'h00;
      13'd5840: x = 8'h00;
      13'd5841: x = 8'h00;
      13'd5842: x = 8'h00;
      13'd5843: x = 8'h00;
      13'd5844: x = 8'h00;
      13'd5845: x = 8'h00;
      13'd5846: x = 8'h00;
      13'd5847: x = 8'h00;
      13'd5848: x = 8'h00;
      13'd5849: x = 8'h00;
      13'd5850: x = 8'h00;
      13'd5851: x = 8'h00;
      13'd5852: x = 8'h00;
      13'd5853: x = 8'h00;
      13'd5854: x = 8'h00;
      13'd5855: x = 8'h00;
      13'd5856: x = 8'h00;
      13'd5857: x = 8'h00;
      13'd5858: x = 8'h00;
      13'd5859: x = 8'h00;
      13'd5860: x = 8'h00;
      13'd5861: x = 8'h00;
      13'd5862: x = 8'h00;
      13'd5863: x = 8'h00;
      13'd5864: x = 8'h00;
      13'd5865: x = 8'h00;
      13'd5866: x = 8'h00;
      13'd5867: x = 8'h00;
      13'd5868: x = 8'h00;
      13'd5869: x = 8'h00;
      13'd5870: x = 8'h00;
      13'd5871: x = 8'h00;
      13'd5872: x = 8'h00;
      13'd5873: x = 8'h00;
      13'd5874: x = 8'h00;
      13'd5875: x = 8'h00;
      13'd5876: x = 8'h00;
      13'd5877: x = 8'h00;
      13'd5878: x = 8'h00;
      13'd5879: x = 8'h00;
      13'd5880: x = 8'h00;
      13'd5881: x = 8'h00;
      13'd5882: x = 8'h00;
      13'd5883: x = 8'h00;
      13'd5884: x = 8'h00;
      13'd5885: x = 8'h00;
      13'd5886: x = 8'h00;
      13'd5887: x = 8'h00;
      13'd5888: x = 8'h00;
      13'd5889: x = 8'h00;
      13'd5890: x = 8'h00;
      13'd5891: x = 8'h00;
      13'd5892: x = 8'h00;
      13'd5893: x = 8'h00;
      13'd5894: x = 8'h00;
      13'd5895: x = 8'h00;
      13'd5896: x = 8'h00;
      13'd5897: x = 8'h00;
      13'd5898: x = 8'h00;
      13'd5899: x = 8'h00;
      13'd5900: x = 8'h00;
      13'd5901: x = 8'h00;
      13'd5902: x = 8'h00;
      13'd5903: x = 8'h00;
      13'd5904: x = 8'h00;
      13'd5905: x = 8'h00;
      13'd5906: x = 8'h00;
      13'd5907: x = 8'h00;
      13'd5908: x = 8'h00;
      13'd5909: x = 8'h00;
      13'd5910: x = 8'h00;
      13'd5911: x = 8'h00;
      13'd5912: x = 8'h00;
      13'd5913: x = 8'h00;
      13'd5914: x = 8'h00;
      13'd5915: x = 8'h00;
      13'd5916: x = 8'h00;
      13'd5917: x = 8'h00;
      13'd5918: x = 8'h00;
      13'd5919: x = 8'h00;
      13'd5920: x = 8'h00;
      13'd5921: x = 8'h00;
      13'd5922: x = 8'h00;
      13'd5923: x = 8'h00;
      13'd5924: x = 8'h00;
      13'd5925: x = 8'h00;
      13'd5926: x = 8'h00;
      13'd5927: x = 8'h00;
      13'd5928: x = 8'h00;
      13'd5929: x = 8'h00;
      13'd5930: x = 8'h00;
      13'd5931: x = 8'h00;
      13'd5932: x = 8'h00;
      13'd5933: x = 8'h00;
      13'd5934: x = 8'h00;
      13'd5935: x = 8'h00;
      13'd5936: x = 8'h00;
      13'd5937: x = 8'h00;
      13'd5938: x = 8'h00;
      13'd5939: x = 8'h00;
      13'd5940: x = 8'h00;
      13'd5941: x = 8'h00;
      13'd5942: x = 8'h00;
      13'd5943: x = 8'h00;
      13'd5944: x = 8'h00;
      13'd5945: x = 8'h00;
      13'd5946: x = 8'h00;
      13'd5947: x = 8'h00;
      13'd5948: x = 8'h00;
      13'd5949: x = 8'h00;
      13'd5950: x = 8'h00;
      13'd5951: x = 8'h00;
      13'd5952: x = 8'h00;
      13'd5953: x = 8'h00;
      13'd5954: x = 8'h00;
      13'd5955: x = 8'h00;
      13'd5956: x = 8'h00;
      13'd5957: x = 8'h00;
      13'd5958: x = 8'h00;
      13'd5959: x = 8'h00;
      13'd5960: x = 8'h00;
      13'd5961: x = 8'h00;
      13'd5962: x = 8'h00;
      13'd5963: x = 8'h00;
      13'd5964: x = 8'h00;
      13'd5965: x = 8'h00;
      13'd5966: x = 8'h00;
      13'd5967: x = 8'h00;
      13'd5968: x = 8'h00;
      13'd5969: x = 8'h00;
      13'd5970: x = 8'h00;
      13'd5971: x = 8'h00;
      13'd5972: x = 8'h00;
      13'd5973: x = 8'h00;
      13'd5974: x = 8'h00;
      13'd5975: x = 8'h00;
      13'd5976: x = 8'h00;
      13'd5977: x = 8'h00;
      13'd5978: x = 8'h00;
      13'd5979: x = 8'h00;
      13'd5980: x = 8'h00;
      13'd5981: x = 8'h00;
      13'd5982: x = 8'h00;
      13'd5983: x = 8'h00;
      13'd5984: x = 8'h00;
      13'd5985: x = 8'h00;
      13'd5986: x = 8'h00;
      13'd5987: x = 8'h00;
      13'd5988: x = 8'h00;
      13'd5989: x = 8'h00;
      13'd5990: x = 8'h00;
      13'd5991: x = 8'h00;
      13'd5992: x = 8'h00;
      13'd5993: x = 8'h00;
      13'd5994: x = 8'h00;
      13'd5995: x = 8'h00;
      13'd5996: x = 8'h00;
      13'd5997: x = 8'h00;
      13'd5998: x = 8'h00;
      13'd5999: x = 8'h00;
      13'd6000: x = 8'h00;
      13'd6001: x = 8'h00;
      13'd6002: x = 8'h00;
      13'd6003: x = 8'h00;
      13'd6004: x = 8'h00;
      13'd6005: x = 8'h00;
      13'd6006: x = 8'h00;
      13'd6007: x = 8'h00;
      13'd6008: x = 8'h00;
      13'd6009: x = 8'h00;
      13'd6010: x = 8'h00;
      13'd6011: x = 8'h00;
      13'd6012: x = 8'h00;
      13'd6013: x = 8'h00;
      13'd6014: x = 8'h00;
      13'd6015: x = 8'h00;
      13'd6016: x = 8'h00;
      13'd6017: x = 8'h00;
      13'd6018: x = 8'h00;
      13'd6019: x = 8'h00;
      13'd6020: x = 8'h00;
      13'd6021: x = 8'h00;
      13'd6022: x = 8'h00;
      13'd6023: x = 8'h00;
      13'd6024: x = 8'h00;
      13'd6025: x = 8'h00;
      13'd6026: x = 8'h00;
      13'd6027: x = 8'h00;
      13'd6028: x = 8'h00;
      13'd6029: x = 8'h00;
      13'd6030: x = 8'h00;
      13'd6031: x = 8'h00;
      13'd6032: x = 8'h00;
      13'd6033: x = 8'h00;
      13'd6034: x = 8'h00;
      13'd6035: x = 8'h00;
      13'd6036: x = 8'h00;
      13'd6037: x = 8'h00;
      13'd6038: x = 8'h00;
      13'd6039: x = 8'h00;
      13'd6040: x = 8'h00;
      13'd6041: x = 8'h00;
      13'd6042: x = 8'h00;
      13'd6043: x = 8'h00;
      13'd6044: x = 8'h00;
      13'd6045: x = 8'h00;
      13'd6046: x = 8'h00;
      13'd6047: x = 8'h00;
      13'd6048: x = 8'h00;
      13'd6049: x = 8'h00;
      13'd6050: x = 8'h00;
      13'd6051: x = 8'h00;
      13'd6052: x = 8'h00;
      13'd6053: x = 8'h00;
      13'd6054: x = 8'h00;
      13'd6055: x = 8'h00;
      13'd6056: x = 8'h00;
      13'd6057: x = 8'h00;
      13'd6058: x = 8'h00;
      13'd6059: x = 8'h00;
      13'd6060: x = 8'h00;
      13'd6061: x = 8'h00;
      13'd6062: x = 8'h00;
      13'd6063: x = 8'h00;
      13'd6064: x = 8'h00;
      13'd6065: x = 8'h00;
      13'd6066: x = 8'h00;
      13'd6067: x = 8'h00;
      13'd6068: x = 8'h00;
      13'd6069: x = 8'h00;
      13'd6070: x = 8'h00;
      13'd6071: x = 8'h00;
      13'd6072: x = 8'h00;
      13'd6073: x = 8'h00;
      13'd6074: x = 8'h00;
      13'd6075: x = 8'h00;
      13'd6076: x = 8'h00;
      13'd6077: x = 8'h00;
      13'd6078: x = 8'h00;
      13'd6079: x = 8'h00;
      13'd6080: x = 8'h00;
      13'd6081: x = 8'h00;
      13'd6082: x = 8'h00;
      13'd6083: x = 8'h00;
      13'd6084: x = 8'h00;
      13'd6085: x = 8'h00;
      13'd6086: x = 8'h00;
      13'd6087: x = 8'h00;
      13'd6088: x = 8'h00;
      13'd6089: x = 8'h00;
      13'd6090: x = 8'h00;
      13'd6091: x = 8'h00;
      13'd6092: x = 8'h00;
      13'd6093: x = 8'h00;
      13'd6094: x = 8'h00;
      13'd6095: x = 8'h00;
      13'd6096: x = 8'h00;
      13'd6097: x = 8'h00;
      13'd6098: x = 8'h00;
      13'd6099: x = 8'h00;
      13'd6100: x = 8'h00;
      13'd6101: x = 8'h00;
      13'd6102: x = 8'h00;
      13'd6103: x = 8'h00;
      13'd6104: x = 8'h00;
      13'd6105: x = 8'h00;
      13'd6106: x = 8'h00;
      13'd6107: x = 8'h00;
      13'd6108: x = 8'h00;
      13'd6109: x = 8'h00;
      13'd6110: x = 8'h00;
      13'd6111: x = 8'h00;
      13'd6112: x = 8'h00;
      13'd6113: x = 8'h00;
      13'd6114: x = 8'h00;
      13'd6115: x = 8'h00;
      13'd6116: x = 8'h00;
      13'd6117: x = 8'h00;
      13'd6118: x = 8'h00;
      13'd6119: x = 8'h00;
      13'd6120: x = 8'h00;
      13'd6121: x = 8'h00;
      13'd6122: x = 8'h00;
      13'd6123: x = 8'h00;
      13'd6124: x = 8'h00;
      13'd6125: x = 8'h00;
      13'd6126: x = 8'h00;
      13'd6127: x = 8'h00;
      13'd6128: x = 8'h00;
      13'd6129: x = 8'h00;
      13'd6130: x = 8'h00;
      13'd6131: x = 8'h00;
      13'd6132: x = 8'h00;
      13'd6133: x = 8'h00;
      13'd6134: x = 8'h00;
      13'd6135: x = 8'h00;
      13'd6136: x = 8'h00;
      13'd6137: x = 8'h00;
      13'd6138: x = 8'h00;
      13'd6139: x = 8'h00;
      13'd6140: x = 8'h00;
      13'd6141: x = 8'h00;
      13'd6142: x = 8'h00;
      13'd6143: x = 8'h00;
      13'd6144: x = 8'h00;
      13'd6145: x = 8'h00;
      13'd6146: x = 8'h00;
      13'd6147: x = 8'h00;
      13'd6148: x = 8'h00;
      13'd6149: x = 8'h00;
      13'd6150: x = 8'h00;
      13'd6151: x = 8'h00;
      13'd6152: x = 8'h00;
      13'd6153: x = 8'h00;
      13'd6154: x = 8'h00;
      13'd6155: x = 8'h00;
      13'd6156: x = 8'h00;
      13'd6157: x = 8'h00;
      13'd6158: x = 8'h00;
      13'd6159: x = 8'h00;
      13'd6160: x = 8'h00;
      13'd6161: x = 8'h00;
      13'd6162: x = 8'h00;
      13'd6163: x = 8'h00;
      13'd6164: x = 8'h00;
      13'd6165: x = 8'h00;
      13'd6166: x = 8'h00;
      13'd6167: x = 8'h00;
      13'd6168: x = 8'h00;
      13'd6169: x = 8'h00;
      13'd6170: x = 8'h00;
      13'd6171: x = 8'h00;
      13'd6172: x = 8'h00;
      13'd6173: x = 8'h00;
      13'd6174: x = 8'h00;
      13'd6175: x = 8'h00;
      13'd6176: x = 8'h00;
      13'd6177: x = 8'h00;
      13'd6178: x = 8'h00;
      13'd6179: x = 8'h00;
      13'd6180: x = 8'h00;
      13'd6181: x = 8'h00;
      13'd6182: x = 8'h00;
      13'd6183: x = 8'h00;
      13'd6184: x = 8'h00;
      13'd6185: x = 8'h00;
      13'd6186: x = 8'h00;
      13'd6187: x = 8'h00;
      13'd6188: x = 8'h00;
      13'd6189: x = 8'h00;
      13'd6190: x = 8'h00;
      13'd6191: x = 8'h00;
      13'd6192: x = 8'h00;
      13'd6193: x = 8'h00;
      13'd6194: x = 8'h00;
      13'd6195: x = 8'h00;
      13'd6196: x = 8'h00;
      13'd6197: x = 8'h00;
      13'd6198: x = 8'h00;
      13'd6199: x = 8'h00;
      13'd6200: x = 8'h00;
      13'd6201: x = 8'h00;
      13'd6202: x = 8'h00;
      13'd6203: x = 8'h00;
      13'd6204: x = 8'h00;
      13'd6205: x = 8'h00;
      13'd6206: x = 8'h00;
      13'd6207: x = 8'h00;
      13'd6208: x = 8'h00;
      13'd6209: x = 8'h00;
      13'd6210: x = 8'h00;
      13'd6211: x = 8'h00;
      13'd6212: x = 8'h00;
      13'd6213: x = 8'h00;
      13'd6214: x = 8'h00;
      13'd6215: x = 8'h00;
      13'd6216: x = 8'h00;
      13'd6217: x = 8'h00;
      13'd6218: x = 8'h00;
      13'd6219: x = 8'h00;
      13'd6220: x = 8'h00;
      13'd6221: x = 8'h00;
      13'd6222: x = 8'h00;
      13'd6223: x = 8'h00;
      13'd6224: x = 8'h00;
      13'd6225: x = 8'h00;
      13'd6226: x = 8'h00;
      13'd6227: x = 8'h00;
      13'd6228: x = 8'h00;
      13'd6229: x = 8'h00;
      13'd6230: x = 8'h00;
      13'd6231: x = 8'h00;
      13'd6232: x = 8'h00;
      13'd6233: x = 8'h00;
      13'd6234: x = 8'h00;
      13'd6235: x = 8'h00;
      13'd6236: x = 8'h00;
      13'd6237: x = 8'h00;
      13'd6238: x = 8'h00;
      13'd6239: x = 8'h00;
      13'd6240: x = 8'h00;
      13'd6241: x = 8'h00;
      13'd6242: x = 8'h00;
      13'd6243: x = 8'h00;
      13'd6244: x = 8'h00;
      13'd6245: x = 8'h00;
      13'd6246: x = 8'h00;
      13'd6247: x = 8'h00;
      13'd6248: x = 8'h00;
      13'd6249: x = 8'h00;
      13'd6250: x = 8'h00;
      13'd6251: x = 8'h00;
      13'd6252: x = 8'h00;
      13'd6253: x = 8'h00;
      13'd6254: x = 8'h00;
      13'd6255: x = 8'h00;
      13'd6256: x = 8'h00;
      13'd6257: x = 8'h00;
      13'd6258: x = 8'h00;
      13'd6259: x = 8'h00;
      13'd6260: x = 8'h00;
      13'd6261: x = 8'h00;
      13'd6262: x = 8'h00;
      13'd6263: x = 8'h00;
      13'd6264: x = 8'h00;
      13'd6265: x = 8'h00;
      13'd6266: x = 8'h00;
      13'd6267: x = 8'h00;
      13'd6268: x = 8'h00;
      13'd6269: x = 8'h00;
      13'd6270: x = 8'h00;
      13'd6271: x = 8'h00;
      13'd6272: x = 8'h00;
      13'd6273: x = 8'h00;
      13'd6274: x = 8'h00;
      13'd6275: x = 8'h00;
      13'd6276: x = 8'h00;
      13'd6277: x = 8'h00;
      13'd6278: x = 8'h00;
      13'd6279: x = 8'h00;
      13'd6280: x = 8'h00;
      13'd6281: x = 8'h00;
      13'd6282: x = 8'h00;
      13'd6283: x = 8'h00;
      13'd6284: x = 8'h00;
      13'd6285: x = 8'h00;
      13'd6286: x = 8'h00;
      13'd6287: x = 8'h00;
      13'd6288: x = 8'h00;
      13'd6289: x = 8'h00;
      13'd6290: x = 8'h00;
      13'd6291: x = 8'h00;
      13'd6292: x = 8'h00;
      13'd6293: x = 8'h00;
      13'd6294: x = 8'h00;
      13'd6295: x = 8'h00;
      13'd6296: x = 8'h00;
      13'd6297: x = 8'h00;
      13'd6298: x = 8'h00;
      13'd6299: x = 8'h00;
      13'd6300: x = 8'h00;
      13'd6301: x = 8'h00;
      13'd6302: x = 8'h00;
      13'd6303: x = 8'h00;
      13'd6304: x = 8'h00;
      13'd6305: x = 8'h00;
      13'd6306: x = 8'h00;
      13'd6307: x = 8'h00;
      13'd6308: x = 8'h00;
      13'd6309: x = 8'h00;
      13'd6310: x = 8'h00;
      13'd6311: x = 8'h00;
      13'd6312: x = 8'h00;
      13'd6313: x = 8'h00;
      13'd6314: x = 8'h00;
      13'd6315: x = 8'h00;
      13'd6316: x = 8'h00;
      13'd6317: x = 8'h00;
      13'd6318: x = 8'h00;
      13'd6319: x = 8'h00;
      13'd6320: x = 8'h00;
      13'd6321: x = 8'h00;
      13'd6322: x = 8'h00;
      13'd6323: x = 8'h00;
      13'd6324: x = 8'h00;
      13'd6325: x = 8'h00;
      13'd6326: x = 8'h00;
      13'd6327: x = 8'h00;
      13'd6328: x = 8'h00;
      13'd6329: x = 8'h00;
      13'd6330: x = 8'h00;
      13'd6331: x = 8'h00;
      13'd6332: x = 8'h00;
      13'd6333: x = 8'h00;
      13'd6334: x = 8'h00;
      13'd6335: x = 8'h00;
      13'd6336: x = 8'h00;
      13'd6337: x = 8'h00;
      13'd6338: x = 8'h00;
      13'd6339: x = 8'h00;
      13'd6340: x = 8'h00;
      13'd6341: x = 8'h00;
      13'd6342: x = 8'h00;
      13'd6343: x = 8'h00;
      13'd6344: x = 8'h00;
      13'd6345: x = 8'h00;
      13'd6346: x = 8'h00;
      13'd6347: x = 8'h00;
      13'd6348: x = 8'h00;
      13'd6349: x = 8'h00;
      13'd6350: x = 8'h00;
      13'd6351: x = 8'h00;
      13'd6352: x = 8'h00;
      13'd6353: x = 8'h00;
      13'd6354: x = 8'h00;
      13'd6355: x = 8'h00;
      13'd6356: x = 8'h00;
      13'd6357: x = 8'h00;
      13'd6358: x = 8'h00;
      13'd6359: x = 8'h00;
      13'd6360: x = 8'h00;
      13'd6361: x = 8'h00;
      13'd6362: x = 8'h00;
      13'd6363: x = 8'h00;
      13'd6364: x = 8'h00;
      13'd6365: x = 8'h00;
      13'd6366: x = 8'h00;
      13'd6367: x = 8'h00;
      13'd6368: x = 8'h00;
      13'd6369: x = 8'h00;
      13'd6370: x = 8'h00;
      13'd6371: x = 8'h00;
      13'd6372: x = 8'h00;
      13'd6373: x = 8'h00;
      13'd6374: x = 8'h00;
      13'd6375: x = 8'h00;
      13'd6376: x = 8'h00;
      13'd6377: x = 8'h00;
      13'd6378: x = 8'h00;
      13'd6379: x = 8'h00;
      13'd6380: x = 8'h00;
      13'd6381: x = 8'h00;
      13'd6382: x = 8'h00;
      13'd6383: x = 8'h00;
      13'd6384: x = 8'h00;
      13'd6385: x = 8'h00;
      13'd6386: x = 8'h00;
      13'd6387: x = 8'h00;
      13'd6388: x = 8'h00;
      13'd6389: x = 8'h00;
      13'd6390: x = 8'h00;
      13'd6391: x = 8'h00;
      13'd6392: x = 8'h00;
      13'd6393: x = 8'h00;
      13'd6394: x = 8'h00;
      13'd6395: x = 8'h00;
      13'd6396: x = 8'h00;
      13'd6397: x = 8'h00;
      13'd6398: x = 8'h00;
      13'd6399: x = 8'h00;
      13'd6400: x = 8'h00;
      13'd6401: x = 8'h00;
      13'd6402: x = 8'h00;
      13'd6403: x = 8'h00;
      13'd6404: x = 8'h00;
      13'd6405: x = 8'h00;
      13'd6406: x = 8'h00;
      13'd6407: x = 8'h00;
      13'd6408: x = 8'h00;
      13'd6409: x = 8'h00;
      13'd6410: x = 8'h00;
      13'd6411: x = 8'h00;
      13'd6412: x = 8'h00;
      13'd6413: x = 8'h00;
      13'd6414: x = 8'h00;
      13'd6415: x = 8'h00;
      13'd6416: x = 8'h00;
      13'd6417: x = 8'h00;
      13'd6418: x = 8'h00;
      13'd6419: x = 8'h00;
      13'd6420: x = 8'h00;
      13'd6421: x = 8'h00;
      13'd6422: x = 8'h00;
      13'd6423: x = 8'h00;
      13'd6424: x = 8'h00;
      13'd6425: x = 8'h00;
      13'd6426: x = 8'h00;
      13'd6427: x = 8'h00;
      13'd6428: x = 8'h00;
      13'd6429: x = 8'h00;
      13'd6430: x = 8'h00;
      13'd6431: x = 8'h00;
      13'd6432: x = 8'h00;
      13'd6433: x = 8'h00;
      13'd6434: x = 8'h00;
      13'd6435: x = 8'h00;
      13'd6436: x = 8'h00;
      13'd6437: x = 8'h00;
      13'd6438: x = 8'h00;
      13'd6439: x = 8'h00;
      13'd6440: x = 8'h00;
      13'd6441: x = 8'h00;
      13'd6442: x = 8'h00;
      13'd6443: x = 8'h00;
      13'd6444: x = 8'h00;
      13'd6445: x = 8'h00;
      13'd6446: x = 8'h00;
      13'd6447: x = 8'h00;
      13'd6448: x = 8'h00;
      13'd6449: x = 8'h00;
      13'd6450: x = 8'h00;
      13'd6451: x = 8'h00;
      13'd6452: x = 8'h00;
      13'd6453: x = 8'h00;
      13'd6454: x = 8'h00;
      13'd6455: x = 8'h00;
      13'd6456: x = 8'h00;
      13'd6457: x = 8'h00;
      13'd6458: x = 8'h00;
      13'd6459: x = 8'h00;
      13'd6460: x = 8'h00;
      13'd6461: x = 8'h00;
      13'd6462: x = 8'h00;
      13'd6463: x = 8'h00;
      13'd6464: x = 8'h00;
      13'd6465: x = 8'h00;
      13'd6466: x = 8'h00;
      13'd6467: x = 8'h00;
      13'd6468: x = 8'h00;
      13'd6469: x = 8'h00;
      13'd6470: x = 8'h00;
      13'd6471: x = 8'h00;
      13'd6472: x = 8'h00;
      13'd6473: x = 8'h00;
      13'd6474: x = 8'h00;
      13'd6475: x = 8'h00;
      13'd6476: x = 8'h00;
      13'd6477: x = 8'h00;
      13'd6478: x = 8'h00;
      13'd6479: x = 8'h00;
      13'd6480: x = 8'h00;
      13'd6481: x = 8'h00;
      13'd6482: x = 8'h00;
      13'd6483: x = 8'h00;
      13'd6484: x = 8'h00;
      13'd6485: x = 8'h00;
      13'd6486: x = 8'h00;
      13'd6487: x = 8'h00;
      13'd6488: x = 8'h00;
      13'd6489: x = 8'h00;
      13'd6490: x = 8'h00;
      13'd6491: x = 8'h00;
      13'd6492: x = 8'h00;
      13'd6493: x = 8'h00;
      13'd6494: x = 8'h00;
      13'd6495: x = 8'h00;
      13'd6496: x = 8'h00;
      13'd6497: x = 8'h00;
      13'd6498: x = 8'h00;
      13'd6499: x = 8'h00;
      13'd6500: x = 8'h00;
      13'd6501: x = 8'h00;
      13'd6502: x = 8'h00;
      13'd6503: x = 8'h00;
      13'd6504: x = 8'h00;
      13'd6505: x = 8'h00;
      13'd6506: x = 8'h00;
      13'd6507: x = 8'h00;
      13'd6508: x = 8'h00;
      13'd6509: x = 8'h00;
      13'd6510: x = 8'h00;
      13'd6511: x = 8'h00;
      13'd6512: x = 8'h00;
      13'd6513: x = 8'h00;
      13'd6514: x = 8'h00;
      13'd6515: x = 8'h00;
      13'd6516: x = 8'h00;
      13'd6517: x = 8'h00;
      13'd6518: x = 8'h00;
      13'd6519: x = 8'h00;
      13'd6520: x = 8'h00;
      13'd6521: x = 8'h00;
      13'd6522: x = 8'h00;
      13'd6523: x = 8'h00;
      13'd6524: x = 8'h00;
      13'd6525: x = 8'h00;
      13'd6526: x = 8'h00;
      13'd6527: x = 8'h00;
      13'd6528: x = 8'h00;
      13'd6529: x = 8'h00;
      13'd6530: x = 8'h00;
      13'd6531: x = 8'h00;
      13'd6532: x = 8'h00;
      13'd6533: x = 8'h00;
      13'd6534: x = 8'h00;
      13'd6535: x = 8'h00;
      13'd6536: x = 8'h00;
      13'd6537: x = 8'h00;
      13'd6538: x = 8'h00;
      13'd6539: x = 8'h00;
      13'd6540: x = 8'h00;
      13'd6541: x = 8'h00;
      13'd6542: x = 8'h00;
      13'd6543: x = 8'h00;
      13'd6544: x = 8'h00;
      13'd6545: x = 8'h00;
      13'd6546: x = 8'h00;
      13'd6547: x = 8'h00;
      13'd6548: x = 8'h00;
      13'd6549: x = 8'h00;
      13'd6550: x = 8'h00;
      13'd6551: x = 8'h00;
      13'd6552: x = 8'h00;
      13'd6553: x = 8'h00;
      13'd6554: x = 8'h00;
      13'd6555: x = 8'h00;
      13'd6556: x = 8'h00;
      13'd6557: x = 8'h00;
      13'd6558: x = 8'h00;
      13'd6559: x = 8'h00;
      13'd6560: x = 8'h00;
      13'd6561: x = 8'h00;
      13'd6562: x = 8'h00;
      13'd6563: x = 8'h00;
      13'd6564: x = 8'h00;
      13'd6565: x = 8'h00;
      13'd6566: x = 8'h00;
      13'd6567: x = 8'h00;
      13'd6568: x = 8'h00;
      13'd6569: x = 8'h00;
      13'd6570: x = 8'h00;
      13'd6571: x = 8'h00;
      13'd6572: x = 8'h00;
      13'd6573: x = 8'h00;
      13'd6574: x = 8'h00;
      13'd6575: x = 8'h00;
      13'd6576: x = 8'h00;
      13'd6577: x = 8'h00;
      13'd6578: x = 8'h00;
      13'd6579: x = 8'h00;
      13'd6580: x = 8'h00;
      13'd6581: x = 8'h00;
      13'd6582: x = 8'h00;
      13'd6583: x = 8'h00;
      13'd6584: x = 8'h00;
      13'd6585: x = 8'h00;
      13'd6586: x = 8'h00;
      13'd6587: x = 8'h00;
      13'd6588: x = 8'h00;
      13'd6589: x = 8'h00;
      13'd6590: x = 8'h00;
      13'd6591: x = 8'h00;
      13'd6592: x = 8'h00;
      13'd6593: x = 8'h00;
      13'd6594: x = 8'h00;
      13'd6595: x = 8'h00;
      13'd6596: x = 8'h00;
      13'd6597: x = 8'h00;
      13'd6598: x = 8'h00;
      13'd6599: x = 8'h00;
      13'd6600: x = 8'h00;
      13'd6601: x = 8'h00;
      13'd6602: x = 8'h00;
      13'd6603: x = 8'h00;
      13'd6604: x = 8'h00;
      13'd6605: x = 8'h00;
      13'd6606: x = 8'h00;
      13'd6607: x = 8'h00;
      13'd6608: x = 8'h00;
      13'd6609: x = 8'h00;
      13'd6610: x = 8'h00;
      13'd6611: x = 8'h00;
      13'd6612: x = 8'h00;
      13'd6613: x = 8'h00;
      13'd6614: x = 8'h00;
      13'd6615: x = 8'h00;
      13'd6616: x = 8'h00;
      13'd6617: x = 8'h00;
      13'd6618: x = 8'h00;
      13'd6619: x = 8'h00;
      13'd6620: x = 8'h00;
      13'd6621: x = 8'h00;
      13'd6622: x = 8'h00;
      13'd6623: x = 8'h00;
      13'd6624: x = 8'h00;
      13'd6625: x = 8'h00;
      13'd6626: x = 8'h00;
      13'd6627: x = 8'h00;
      13'd6628: x = 8'h00;
      13'd6629: x = 8'h00;
      13'd6630: x = 8'h00;
      13'd6631: x = 8'h00;
      13'd6632: x = 8'h00;
      13'd6633: x = 8'h00;
      13'd6634: x = 8'h00;
      13'd6635: x = 8'h00;
      13'd6636: x = 8'h00;
      13'd6637: x = 8'h00;
      13'd6638: x = 8'h00;
      13'd6639: x = 8'h00;
      13'd6640: x = 8'h00;
      13'd6641: x = 8'h00;
      13'd6642: x = 8'h00;
      13'd6643: x = 8'h00;
      13'd6644: x = 8'h00;
      13'd6645: x = 8'h00;
      13'd6646: x = 8'h00;
      13'd6647: x = 8'h00;
      13'd6648: x = 8'h00;
      13'd6649: x = 8'h00;
      13'd6650: x = 8'h00;
      13'd6651: x = 8'h00;
      13'd6652: x = 8'h00;
      13'd6653: x = 8'h00;
      13'd6654: x = 8'h00;
      13'd6655: x = 8'h00;
      13'd6656: x = 8'h00;
      13'd6657: x = 8'h00;
      13'd6658: x = 8'h00;
      13'd6659: x = 8'h00;
      13'd6660: x = 8'h00;
      13'd6661: x = 8'h00;
      13'd6662: x = 8'h00;
      13'd6663: x = 8'h00;
      13'd6664: x = 8'h00;
      13'd6665: x = 8'h00;
      13'd6666: x = 8'h00;
      13'd6667: x = 8'h00;
      13'd6668: x = 8'h00;
      13'd6669: x = 8'h00;
      13'd6670: x = 8'h00;
      13'd6671: x = 8'h00;
      13'd6672: x = 8'h00;
      13'd6673: x = 8'h00;
      13'd6674: x = 8'h00;
      13'd6675: x = 8'h00;
      13'd6676: x = 8'h00;
      13'd6677: x = 8'h00;
      13'd6678: x = 8'h00;
      13'd6679: x = 8'h00;
      13'd6680: x = 8'h00;
      13'd6681: x = 8'h00;
      13'd6682: x = 8'h00;
      13'd6683: x = 8'h00;
      13'd6684: x = 8'h00;
      13'd6685: x = 8'h00;
      13'd6686: x = 8'h00;
      13'd6687: x = 8'h00;
      13'd6688: x = 8'h00;
      13'd6689: x = 8'h00;
      13'd6690: x = 8'h00;
      13'd6691: x = 8'h00;
      13'd6692: x = 8'h00;
      13'd6693: x = 8'h00;
      13'd6694: x = 8'h00;
      13'd6695: x = 8'h00;
      13'd6696: x = 8'h00;
      13'd6697: x = 8'h00;
      13'd6698: x = 8'h00;
      13'd6699: x = 8'h00;
      13'd6700: x = 8'h00;
      13'd6701: x = 8'h00;
      13'd6702: x = 8'h00;
      13'd6703: x = 8'h00;
      13'd6704: x = 8'h00;
      13'd6705: x = 8'h00;
      13'd6706: x = 8'h00;
      13'd6707: x = 8'h00;
      13'd6708: x = 8'h00;
      13'd6709: x = 8'h00;
      13'd6710: x = 8'h00;
      13'd6711: x = 8'h00;
      13'd6712: x = 8'h00;
      13'd6713: x = 8'h00;
      13'd6714: x = 8'h00;
      13'd6715: x = 8'h00;
      13'd6716: x = 8'h00;
      13'd6717: x = 8'h00;
      13'd6718: x = 8'h00;
      13'd6719: x = 8'h00;
      13'd6720: x = 8'h00;
      13'd6721: x = 8'h00;
      13'd6722: x = 8'h00;
      13'd6723: x = 8'h00;
      13'd6724: x = 8'h00;
      13'd6725: x = 8'h00;
      13'd6726: x = 8'h00;
      13'd6727: x = 8'h00;
      13'd6728: x = 8'h00;
      13'd6729: x = 8'h00;
      13'd6730: x = 8'h00;
      13'd6731: x = 8'h00;
      13'd6732: x = 8'h00;
      13'd6733: x = 8'h00;
      13'd6734: x = 8'h00;
      13'd6735: x = 8'h00;
      13'd6736: x = 8'h00;
      13'd6737: x = 8'h00;
      13'd6738: x = 8'h00;
      13'd6739: x = 8'h00;
      13'd6740: x = 8'h00;
      13'd6741: x = 8'h00;
      13'd6742: x = 8'h00;
      13'd6743: x = 8'h00;
      13'd6744: x = 8'h00;
      13'd6745: x = 8'h00;
      13'd6746: x = 8'h00;
      13'd6747: x = 8'h00;
      13'd6748: x = 8'h00;
      13'd6749: x = 8'h00;
      13'd6750: x = 8'h00;
      13'd6751: x = 8'h00;
      13'd6752: x = 8'h00;
      13'd6753: x = 8'h00;
      13'd6754: x = 8'h00;
      13'd6755: x = 8'h00;
      13'd6756: x = 8'h00;
      13'd6757: x = 8'h00;
      13'd6758: x = 8'h00;
      13'd6759: x = 8'h00;
      13'd6760: x = 8'h00;
      13'd6761: x = 8'h00;
      13'd6762: x = 8'h00;
      13'd6763: x = 8'h00;
      13'd6764: x = 8'h00;
      13'd6765: x = 8'h00;
      13'd6766: x = 8'h00;
      13'd6767: x = 8'h00;
      13'd6768: x = 8'h00;
      13'd6769: x = 8'h00;
      13'd6770: x = 8'h00;
      13'd6771: x = 8'h00;
      13'd6772: x = 8'h00;
      13'd6773: x = 8'h00;
      13'd6774: x = 8'h00;
      13'd6775: x = 8'h00;
      13'd6776: x = 8'h00;
      13'd6777: x = 8'h00;
      13'd6778: x = 8'h00;
      13'd6779: x = 8'h00;
      13'd6780: x = 8'h00;
      13'd6781: x = 8'h00;
      13'd6782: x = 8'h00;
      13'd6783: x = 8'h00;
      13'd6784: x = 8'h00;
      13'd6785: x = 8'h00;
      13'd6786: x = 8'h00;
      13'd6787: x = 8'h00;
      13'd6788: x = 8'h00;
      13'd6789: x = 8'h00;
      13'd6790: x = 8'h00;
      13'd6791: x = 8'h00;
      13'd6792: x = 8'h00;
      13'd6793: x = 8'h00;
      13'd6794: x = 8'h00;
      13'd6795: x = 8'h00;
      13'd6796: x = 8'h00;
      13'd6797: x = 8'h00;
      13'd6798: x = 8'h00;
      13'd6799: x = 8'h00;
      13'd6800: x = 8'h00;
      13'd6801: x = 8'h00;
      13'd6802: x = 8'h00;
      13'd6803: x = 8'h00;
      13'd6804: x = 8'h00;
      13'd6805: x = 8'h00;
      13'd6806: x = 8'h00;
      13'd6807: x = 8'h00;
      13'd6808: x = 8'h00;
      13'd6809: x = 8'h00;
      13'd6810: x = 8'h00;
      13'd6811: x = 8'h00;
      13'd6812: x = 8'h00;
      13'd6813: x = 8'h00;
      13'd6814: x = 8'h00;
      13'd6815: x = 8'h00;
      13'd6816: x = 8'h00;
      13'd6817: x = 8'h00;
      13'd6818: x = 8'h00;
      13'd6819: x = 8'h00;
      13'd6820: x = 8'h00;
      13'd6821: x = 8'h00;
      13'd6822: x = 8'h00;
      13'd6823: x = 8'h00;
      13'd6824: x = 8'h00;
      13'd6825: x = 8'h00;
      13'd6826: x = 8'h00;
      13'd6827: x = 8'h00;
      13'd6828: x = 8'h00;
      13'd6829: x = 8'h00;
      13'd6830: x = 8'h00;
      13'd6831: x = 8'h00;
      13'd6832: x = 8'h00;
      13'd6833: x = 8'h00;
      13'd6834: x = 8'h00;
      13'd6835: x = 8'h00;
      13'd6836: x = 8'h00;
      13'd6837: x = 8'h00;
      13'd6838: x = 8'h00;
      13'd6839: x = 8'h00;
      13'd6840: x = 8'h00;
      13'd6841: x = 8'h00;
      13'd6842: x = 8'h00;
      13'd6843: x = 8'h00;
      13'd6844: x = 8'h00;
      13'd6845: x = 8'h00;
      13'd6846: x = 8'h00;
      13'd6847: x = 8'h00;
      13'd6848: x = 8'h00;
      13'd6849: x = 8'h00;
      13'd6850: x = 8'h00;
      13'd6851: x = 8'h00;
      13'd6852: x = 8'h00;
      13'd6853: x = 8'h00;
      13'd6854: x = 8'h00;
      13'd6855: x = 8'h00;
      13'd6856: x = 8'h00;
      13'd6857: x = 8'h00;
      13'd6858: x = 8'h00;
      13'd6859: x = 8'h00;
      13'd6860: x = 8'h00;
      13'd6861: x = 8'h00;
      13'd6862: x = 8'h00;
      13'd6863: x = 8'h00;
      13'd6864: x = 8'h00;
      13'd6865: x = 8'h00;
      13'd6866: x = 8'h00;
      13'd6867: x = 8'h00;
      13'd6868: x = 8'h00;
      13'd6869: x = 8'h00;
      13'd6870: x = 8'h00;
      13'd6871: x = 8'h00;
      13'd6872: x = 8'h00;
      13'd6873: x = 8'h00;
      13'd6874: x = 8'h00;
      13'd6875: x = 8'h00;
      13'd6876: x = 8'h00;
      13'd6877: x = 8'h00;
      13'd6878: x = 8'h00;
      13'd6879: x = 8'h00;
      13'd6880: x = 8'h00;
      13'd6881: x = 8'h00;
      13'd6882: x = 8'h00;
      13'd6883: x = 8'h00;
      13'd6884: x = 8'h00;
      13'd6885: x = 8'h00;
      13'd6886: x = 8'h00;
      13'd6887: x = 8'h00;
      13'd6888: x = 8'h00;
      13'd6889: x = 8'h00;
      13'd6890: x = 8'h00;
      13'd6891: x = 8'h00;
      13'd6892: x = 8'h00;
      13'd6893: x = 8'h00;
      13'd6894: x = 8'h00;
      13'd6895: x = 8'h00;
      13'd6896: x = 8'h00;
      13'd6897: x = 8'h00;
      13'd6898: x = 8'h00;
      13'd6899: x = 8'h00;
      13'd6900: x = 8'h00;
      13'd6901: x = 8'h00;
      13'd6902: x = 8'h00;
      13'd6903: x = 8'h00;
      13'd6904: x = 8'h00;
      13'd6905: x = 8'h00;
      13'd6906: x = 8'h00;
      13'd6907: x = 8'h00;
      13'd6908: x = 8'h00;
      13'd6909: x = 8'h00;
      13'd6910: x = 8'h00;
      13'd6911: x = 8'h00;
      13'd6912: x = 8'h00;
      13'd6913: x = 8'h00;
      13'd6914: x = 8'h00;
      13'd6915: x = 8'h00;
      13'd6916: x = 8'h00;
      13'd6917: x = 8'h00;
      13'd6918: x = 8'h00;
      13'd6919: x = 8'h00;
      13'd6920: x = 8'h00;
      13'd6921: x = 8'h00;
      13'd6922: x = 8'h00;
      13'd6923: x = 8'h00;
      13'd6924: x = 8'h00;
      13'd6925: x = 8'h00;
      13'd6926: x = 8'h00;
      13'd6927: x = 8'h00;
      13'd6928: x = 8'h00;
      13'd6929: x = 8'h00;
      13'd6930: x = 8'h00;
      13'd6931: x = 8'h00;
      13'd6932: x = 8'h00;
      13'd6933: x = 8'h00;
      13'd6934: x = 8'h00;
      13'd6935: x = 8'h00;
      13'd6936: x = 8'h00;
      13'd6937: x = 8'h00;
      13'd6938: x = 8'h00;
      13'd6939: x = 8'h00;
      13'd6940: x = 8'h00;
      13'd6941: x = 8'h00;
      13'd6942: x = 8'h00;
      13'd6943: x = 8'h00;
      13'd6944: x = 8'h00;
      13'd6945: x = 8'h00;
      13'd6946: x = 8'h00;
      13'd6947: x = 8'h00;
      13'd6948: x = 8'h00;
      13'd6949: x = 8'h00;
      13'd6950: x = 8'h00;
      13'd6951: x = 8'h00;
      13'd6952: x = 8'h00;
      13'd6953: x = 8'h00;
      13'd6954: x = 8'h00;
      13'd6955: x = 8'h00;
      13'd6956: x = 8'h00;
      13'd6957: x = 8'h00;
      13'd6958: x = 8'h00;
      13'd6959: x = 8'h00;
      13'd6960: x = 8'h00;
      13'd6961: x = 8'h00;
      13'd6962: x = 8'h00;
      13'd6963: x = 8'h00;
      13'd6964: x = 8'h00;
      13'd6965: x = 8'h00;
      13'd6966: x = 8'h00;
      13'd6967: x = 8'h00;
      13'd6968: x = 8'h00;
      13'd6969: x = 8'h00;
      13'd6970: x = 8'h00;
      13'd6971: x = 8'h00;
      13'd6972: x = 8'h00;
      13'd6973: x = 8'h00;
      13'd6974: x = 8'h00;
      13'd6975: x = 8'h00;
      13'd6976: x = 8'h00;
      13'd6977: x = 8'h00;
      13'd6978: x = 8'h00;
      13'd6979: x = 8'h00;
      13'd6980: x = 8'h00;
      13'd6981: x = 8'h00;
      13'd6982: x = 8'h00;
      13'd6983: x = 8'h00;
      13'd6984: x = 8'h00;
      13'd6985: x = 8'h00;
      13'd6986: x = 8'h00;
      13'd6987: x = 8'h00;
      13'd6988: x = 8'h00;
      13'd6989: x = 8'h00;
      13'd6990: x = 8'h00;
      13'd6991: x = 8'h00;
      13'd6992: x = 8'h00;
      13'd6993: x = 8'h00;
      13'd6994: x = 8'h00;
      13'd6995: x = 8'h00;
      13'd6996: x = 8'h00;
      13'd6997: x = 8'h00;
      13'd6998: x = 8'h00;
      13'd6999: x = 8'h00;
      13'd7000: x = 8'h00;
      13'd7001: x = 8'h00;
      13'd7002: x = 8'h00;
      13'd7003: x = 8'h00;
      13'd7004: x = 8'h00;
      13'd7005: x = 8'h00;
      13'd7006: x = 8'h00;
      13'd7007: x = 8'h00;
      13'd7008: x = 8'h00;
      13'd7009: x = 8'h00;
      13'd7010: x = 8'h00;
      13'd7011: x = 8'h00;
      13'd7012: x = 8'h00;
      13'd7013: x = 8'h00;
      13'd7014: x = 8'h00;
      13'd7015: x = 8'h00;
      13'd7016: x = 8'h00;
      13'd7017: x = 8'h00;
      13'd7018: x = 8'h00;
      13'd7019: x = 8'h00;
      13'd7020: x = 8'h00;
      13'd7021: x = 8'h00;
      13'd7022: x = 8'h00;
      13'd7023: x = 8'h00;
      13'd7024: x = 8'h00;
      13'd7025: x = 8'h00;
      13'd7026: x = 8'h00;
      13'd7027: x = 8'h00;
      13'd7028: x = 8'h00;
      13'd7029: x = 8'h00;
      13'd7030: x = 8'h00;
      13'd7031: x = 8'h00;
      13'd7032: x = 8'h00;
      13'd7033: x = 8'h00;
      13'd7034: x = 8'h00;
      13'd7035: x = 8'h00;
      13'd7036: x = 8'h00;
      13'd7037: x = 8'h00;
      13'd7038: x = 8'h00;
      13'd7039: x = 8'h00;
      13'd7040: x = 8'h00;
      13'd7041: x = 8'h00;
      13'd7042: x = 8'h00;
      13'd7043: x = 8'h00;
      13'd7044: x = 8'h00;
      13'd7045: x = 8'h00;
      13'd7046: x = 8'h00;
      13'd7047: x = 8'h00;
      13'd7048: x = 8'h00;
      13'd7049: x = 8'h00;
      13'd7050: x = 8'h00;
      13'd7051: x = 8'h00;
      13'd7052: x = 8'h00;
      13'd7053: x = 8'h00;
      13'd7054: x = 8'h00;
      13'd7055: x = 8'h00;
      13'd7056: x = 8'h00;
      13'd7057: x = 8'h00;
      13'd7058: x = 8'h00;
      13'd7059: x = 8'h00;
      13'd7060: x = 8'h00;
      13'd7061: x = 8'h00;
      13'd7062: x = 8'h00;
      13'd7063: x = 8'h00;
      13'd7064: x = 8'h00;
      13'd7065: x = 8'h00;
      13'd7066: x = 8'h00;
      13'd7067: x = 8'h00;
      13'd7068: x = 8'h00;
      13'd7069: x = 8'h00;
      13'd7070: x = 8'h00;
      13'd7071: x = 8'h00;
      13'd7072: x = 8'h00;
      13'd7073: x = 8'h00;
      13'd7074: x = 8'h00;
      13'd7075: x = 8'h00;
      13'd7076: x = 8'h00;
      13'd7077: x = 8'h00;
      13'd7078: x = 8'h00;
      13'd7079: x = 8'h00;
      13'd7080: x = 8'h00;
      13'd7081: x = 8'h00;
      13'd7082: x = 8'h00;
      13'd7083: x = 8'h00;
      13'd7084: x = 8'h00;
      13'd7085: x = 8'h00;
      13'd7086: x = 8'h00;
      13'd7087: x = 8'h00;
      13'd7088: x = 8'h00;
      13'd7089: x = 8'h00;
      13'd7090: x = 8'h00;
      13'd7091: x = 8'h00;
      13'd7092: x = 8'h00;
      13'd7093: x = 8'h00;
      13'd7094: x = 8'h00;
      13'd7095: x = 8'h00;
      13'd7096: x = 8'h00;
      13'd7097: x = 8'h00;
      13'd7098: x = 8'h00;
      13'd7099: x = 8'h00;
      13'd7100: x = 8'h00;
      13'd7101: x = 8'h00;
      13'd7102: x = 8'h00;
      13'd7103: x = 8'h00;
      13'd7104: x = 8'h00;
      13'd7105: x = 8'h00;
      13'd7106: x = 8'h00;
      13'd7107: x = 8'h00;
      13'd7108: x = 8'h00;
      13'd7109: x = 8'h00;
      13'd7110: x = 8'h00;
      13'd7111: x = 8'h00;
      13'd7112: x = 8'h00;
      13'd7113: x = 8'h00;
      13'd7114: x = 8'h00;
      13'd7115: x = 8'h00;
      13'd7116: x = 8'h00;
      13'd7117: x = 8'h00;
      13'd7118: x = 8'h00;
      13'd7119: x = 8'h00;
      13'd7120: x = 8'h00;
      13'd7121: x = 8'h00;
      13'd7122: x = 8'h00;
      13'd7123: x = 8'h00;
      13'd7124: x = 8'h00;
      13'd7125: x = 8'h00;
      13'd7126: x = 8'h00;
      13'd7127: x = 8'h00;
      13'd7128: x = 8'h00;
      13'd7129: x = 8'h00;
      13'd7130: x = 8'h00;
      13'd7131: x = 8'h00;
      13'd7132: x = 8'h00;
      13'd7133: x = 8'h00;
      13'd7134: x = 8'h00;
      13'd7135: x = 8'h00;
      13'd7136: x = 8'h00;
      13'd7137: x = 8'h00;
      13'd7138: x = 8'h00;
      13'd7139: x = 8'h00;
      13'd7140: x = 8'h00;
      13'd7141: x = 8'h00;
      13'd7142: x = 8'h00;
      13'd7143: x = 8'h00;
      13'd7144: x = 8'h00;
      13'd7145: x = 8'h00;
      13'd7146: x = 8'h00;
      13'd7147: x = 8'h00;
      13'd7148: x = 8'h00;
      13'd7149: x = 8'h00;
      13'd7150: x = 8'h00;
      13'd7151: x = 8'h00;
      13'd7152: x = 8'h00;
      13'd7153: x = 8'h00;
      13'd7154: x = 8'h00;
      13'd7155: x = 8'h00;
      13'd7156: x = 8'h00;
      13'd7157: x = 8'h00;
      13'd7158: x = 8'h00;
      13'd7159: x = 8'h00;
      13'd7160: x = 8'h00;
      13'd7161: x = 8'h00;
      13'd7162: x = 8'h00;
      13'd7163: x = 8'h00;
      13'd7164: x = 8'h00;
      13'd7165: x = 8'h00;
      13'd7166: x = 8'h00;
      13'd7167: x = 8'h00;
      13'd7168: x = 8'h00;
      13'd7169: x = 8'h00;
      13'd7170: x = 8'h00;
      13'd7171: x = 8'h00;
      13'd7172: x = 8'h00;
      13'd7173: x = 8'h00;
      13'd7174: x = 8'h00;
      13'd7175: x = 8'h00;
      13'd7176: x = 8'h00;
      13'd7177: x = 8'h00;
      13'd7178: x = 8'h00;
      13'd7179: x = 8'h00;
      13'd7180: x = 8'h00;
      13'd7181: x = 8'h00;
      13'd7182: x = 8'h00;
      13'd7183: x = 8'h00;
      13'd7184: x = 8'h00;
      13'd7185: x = 8'h00;
      13'd7186: x = 8'h00;
      13'd7187: x = 8'h00;
      13'd7188: x = 8'h00;
      13'd7189: x = 8'h00;
      13'd7190: x = 8'h00;
      13'd7191: x = 8'h00;
      13'd7192: x = 8'h00;
      13'd7193: x = 8'h00;
      13'd7194: x = 8'h00;
      13'd7195: x = 8'h00;
      13'd7196: x = 8'h00;
      13'd7197: x = 8'h00;
      13'd7198: x = 8'h00;
      13'd7199: x = 8'h00;
      13'd7200: x = 8'h00;
      13'd7201: x = 8'h00;
      13'd7202: x = 8'h00;
      13'd7203: x = 8'h00;
      13'd7204: x = 8'h00;
      13'd7205: x = 8'h00;
      13'd7206: x = 8'h00;
      13'd7207: x = 8'h00;
      13'd7208: x = 8'h00;
      13'd7209: x = 8'h00;
      13'd7210: x = 8'h00;
      13'd7211: x = 8'h00;
      13'd7212: x = 8'h00;
      13'd7213: x = 8'h00;
      13'd7214: x = 8'h00;
      13'd7215: x = 8'h00;
      13'd7216: x = 8'h00;
      13'd7217: x = 8'h00;
      13'd7218: x = 8'h00;
      13'd7219: x = 8'h00;
      13'd7220: x = 8'h00;
      13'd7221: x = 8'h00;
      13'd7222: x = 8'h00;
      13'd7223: x = 8'h00;
      13'd7224: x = 8'h00;
      13'd7225: x = 8'h00;
      13'd7226: x = 8'h00;
      13'd7227: x = 8'h00;
      13'd7228: x = 8'h00;
      13'd7229: x = 8'h00;
      13'd7230: x = 8'h00;
      13'd7231: x = 8'h00;
      13'd7232: x = 8'h00;
      13'd7233: x = 8'h00;
      13'd7234: x = 8'h00;
      13'd7235: x = 8'h00;
      13'd7236: x = 8'h00;
      13'd7237: x = 8'h00;
      13'd7238: x = 8'h00;
      13'd7239: x = 8'h00;
      13'd7240: x = 8'h00;
      13'd7241: x = 8'h00;
      13'd7242: x = 8'h00;
      13'd7243: x = 8'h00;
      13'd7244: x = 8'h00;
      13'd7245: x = 8'h00;
      13'd7246: x = 8'h00;
      13'd7247: x = 8'h00;
      13'd7248: x = 8'h00;
      13'd7249: x = 8'h00;
      13'd7250: x = 8'h00;
      13'd7251: x = 8'h00;
      13'd7252: x = 8'h00;
      13'd7253: x = 8'h00;
      13'd7254: x = 8'h00;
      13'd7255: x = 8'h00;
      13'd7256: x = 8'h00;
      13'd7257: x = 8'h00;
      13'd7258: x = 8'h00;
      13'd7259: x = 8'h00;
      13'd7260: x = 8'h00;
      13'd7261: x = 8'h00;
      13'd7262: x = 8'h00;
      13'd7263: x = 8'h00;
      13'd7264: x = 8'h00;
      13'd7265: x = 8'h00;
      13'd7266: x = 8'h00;
      13'd7267: x = 8'h00;
      13'd7268: x = 8'h00;
      13'd7269: x = 8'h00;
      13'd7270: x = 8'h00;
      13'd7271: x = 8'h00;
      13'd7272: x = 8'h00;
      13'd7273: x = 8'h00;
      13'd7274: x = 8'h00;
      13'd7275: x = 8'h00;
      13'd7276: x = 8'h00;
      13'd7277: x = 8'h00;
      13'd7278: x = 8'h00;
      13'd7279: x = 8'h00;
      13'd7280: x = 8'h00;
      13'd7281: x = 8'h00;
      13'd7282: x = 8'h00;
      13'd7283: x = 8'h00;
      13'd7284: x = 8'h00;
      13'd7285: x = 8'h00;
      13'd7286: x = 8'h00;
      13'd7287: x = 8'h00;
      13'd7288: x = 8'h00;
      13'd7289: x = 8'h00;
      13'd7290: x = 8'h00;
      13'd7291: x = 8'h00;
      13'd7292: x = 8'h00;
      13'd7293: x = 8'h00;
      13'd7294: x = 8'h00;
      13'd7295: x = 8'h00;
      13'd7296: x = 8'h00;
      13'd7297: x = 8'h00;
      13'd7298: x = 8'h00;
      13'd7299: x = 8'h00;
      13'd7300: x = 8'h00;
      13'd7301: x = 8'h00;
      13'd7302: x = 8'h00;
      13'd7303: x = 8'h00;
      13'd7304: x = 8'h00;
      13'd7305: x = 8'h00;
      13'd7306: x = 8'h00;
      13'd7307: x = 8'h00;
      13'd7308: x = 8'h00;
      13'd7309: x = 8'h00;
      13'd7310: x = 8'h00;
      13'd7311: x = 8'h00;
      13'd7312: x = 8'h00;
      13'd7313: x = 8'h00;
      13'd7314: x = 8'h00;
      13'd7315: x = 8'h00;
      13'd7316: x = 8'h00;
      13'd7317: x = 8'h00;
      13'd7318: x = 8'h00;
      13'd7319: x = 8'h00;
      13'd7320: x = 8'h00;
      13'd7321: x = 8'h00;
      13'd7322: x = 8'h00;
      13'd7323: x = 8'h00;
      13'd7324: x = 8'h00;
      13'd7325: x = 8'h00;
      13'd7326: x = 8'h00;
      13'd7327: x = 8'h00;
      13'd7328: x = 8'h00;
      13'd7329: x = 8'h00;
      13'd7330: x = 8'h00;
      13'd7331: x = 8'h00;
      13'd7332: x = 8'h00;
      13'd7333: x = 8'h00;
      13'd7334: x = 8'h00;
      13'd7335: x = 8'h00;
      13'd7336: x = 8'h00;
      13'd7337: x = 8'h00;
      13'd7338: x = 8'h00;
      13'd7339: x = 8'h00;
      13'd7340: x = 8'h00;
      13'd7341: x = 8'h00;
      13'd7342: x = 8'h00;
      13'd7343: x = 8'h00;
      13'd7344: x = 8'h00;
      13'd7345: x = 8'h00;
      13'd7346: x = 8'h00;
      13'd7347: x = 8'h00;
      13'd7348: x = 8'h00;
      13'd7349: x = 8'h00;
      13'd7350: x = 8'h00;
      13'd7351: x = 8'h00;
      13'd7352: x = 8'h00;
      13'd7353: x = 8'h00;
      13'd7354: x = 8'h00;
      13'd7355: x = 8'h00;
      13'd7356: x = 8'h00;
      13'd7357: x = 8'h00;
      13'd7358: x = 8'h00;
      13'd7359: x = 8'h00;
      13'd7360: x = 8'h00;
      13'd7361: x = 8'h00;
      13'd7362: x = 8'h00;
      13'd7363: x = 8'h00;
      13'd7364: x = 8'h00;
      13'd7365: x = 8'h00;
      13'd7366: x = 8'h00;
      13'd7367: x = 8'h00;
      13'd7368: x = 8'h00;
      13'd7369: x = 8'h00;
      13'd7370: x = 8'h00;
      13'd7371: x = 8'h00;
      13'd7372: x = 8'h00;
      13'd7373: x = 8'h00;
      13'd7374: x = 8'h00;
      13'd7375: x = 8'h00;
      13'd7376: x = 8'h00;
      13'd7377: x = 8'h00;
      13'd7378: x = 8'h00;
      13'd7379: x = 8'h00;
      13'd7380: x = 8'h00;
      13'd7381: x = 8'h00;
      13'd7382: x = 8'h00;
      13'd7383: x = 8'h00;
      13'd7384: x = 8'h00;
      13'd7385: x = 8'h00;
      13'd7386: x = 8'h00;
      13'd7387: x = 8'h00;
      13'd7388: x = 8'h00;
      13'd7389: x = 8'h00;
      13'd7390: x = 8'h00;
      13'd7391: x = 8'h00;
      13'd7392: x = 8'h00;
      13'd7393: x = 8'h00;
      13'd7394: x = 8'h00;
      13'd7395: x = 8'h00;
      13'd7396: x = 8'h00;
      13'd7397: x = 8'h00;
      13'd7398: x = 8'h00;
      13'd7399: x = 8'h00;
      13'd7400: x = 8'h00;
      13'd7401: x = 8'h00;
      13'd7402: x = 8'h00;
      13'd7403: x = 8'h00;
      13'd7404: x = 8'h00;
      13'd7405: x = 8'h00;
      13'd7406: x = 8'h00;
      13'd7407: x = 8'h00;
      13'd7408: x = 8'h00;
      13'd7409: x = 8'h00;
      13'd7410: x = 8'h00;
      13'd7411: x = 8'h00;
      13'd7412: x = 8'h00;
      13'd7413: x = 8'h00;
      13'd7414: x = 8'h00;
      13'd7415: x = 8'h00;
      13'd7416: x = 8'h00;
      13'd7417: x = 8'h00;
      13'd7418: x = 8'h00;
      13'd7419: x = 8'h00;
      13'd7420: x = 8'h00;
      13'd7421: x = 8'h00;
      13'd7422: x = 8'h00;
      13'd7423: x = 8'h00;
      13'd7424: x = 8'h00;
      13'd7425: x = 8'h00;
      13'd7426: x = 8'h00;
      13'd7427: x = 8'h00;
      13'd7428: x = 8'h00;
      13'd7429: x = 8'h00;
      13'd7430: x = 8'h00;
      13'd7431: x = 8'h00;
      13'd7432: x = 8'h00;
      13'd7433: x = 8'h00;
      13'd7434: x = 8'h00;
      13'd7435: x = 8'h00;
      13'd7436: x = 8'h00;
      13'd7437: x = 8'h00;
      13'd7438: x = 8'h00;
      13'd7439: x = 8'h00;
      13'd7440: x = 8'h00;
      13'd7441: x = 8'h00;
      13'd7442: x = 8'h00;
      13'd7443: x = 8'h00;
      13'd7444: x = 8'h00;
      13'd7445: x = 8'h00;
      13'd7446: x = 8'h00;
      13'd7447: x = 8'h00;
      13'd7448: x = 8'h00;
      13'd7449: x = 8'h00;
      13'd7450: x = 8'h00;
      13'd7451: x = 8'h00;
      13'd7452: x = 8'h00;
      13'd7453: x = 8'h00;
      13'd7454: x = 8'h00;
      13'd7455: x = 8'h00;
      13'd7456: x = 8'h00;
      13'd7457: x = 8'h00;
      13'd7458: x = 8'h00;
      13'd7459: x = 8'h00;
      13'd7460: x = 8'h00;
      13'd7461: x = 8'h00;
      13'd7462: x = 8'h00;
      13'd7463: x = 8'h00;
      13'd7464: x = 8'h00;
      13'd7465: x = 8'h00;
      13'd7466: x = 8'h00;
      13'd7467: x = 8'h00;
      13'd7468: x = 8'h00;
      13'd7469: x = 8'h00;
      13'd7470: x = 8'h00;
      13'd7471: x = 8'h00;
      13'd7472: x = 8'h00;
      13'd7473: x = 8'h00;
      13'd7474: x = 8'h00;
      13'd7475: x = 8'h00;
      13'd7476: x = 8'h00;
      13'd7477: x = 8'h00;
      13'd7478: x = 8'h00;
      13'd7479: x = 8'h00;
      13'd7480: x = 8'h00;
      13'd7481: x = 8'h00;
      13'd7482: x = 8'h00;
      13'd7483: x = 8'h00;
      13'd7484: x = 8'h00;
      13'd7485: x = 8'h00;
      13'd7486: x = 8'h00;
      13'd7487: x = 8'h00;
      13'd7488: x = 8'h00;
      13'd7489: x = 8'h00;
      13'd7490: x = 8'h00;
      13'd7491: x = 8'h00;
      13'd7492: x = 8'h00;
      13'd7493: x = 8'h00;
      13'd7494: x = 8'h00;
      13'd7495: x = 8'h00;
      13'd7496: x = 8'h00;
      13'd7497: x = 8'h00;
      13'd7498: x = 8'h00;
      13'd7499: x = 8'h00;
      13'd7500: x = 8'h00;
      13'd7501: x = 8'h00;
      13'd7502: x = 8'h00;
      13'd7503: x = 8'h00;
      13'd7504: x = 8'h00;
      13'd7505: x = 8'h00;
      13'd7506: x = 8'h00;
      13'd7507: x = 8'h00;
      13'd7508: x = 8'h00;
      13'd7509: x = 8'h00;
      13'd7510: x = 8'h00;
      13'd7511: x = 8'h00;
      13'd7512: x = 8'h00;
      13'd7513: x = 8'h00;
      13'd7514: x = 8'h00;
      13'd7515: x = 8'h00;
      13'd7516: x = 8'h00;
      13'd7517: x = 8'h00;
      13'd7518: x = 8'h00;
      13'd7519: x = 8'h00;
      13'd7520: x = 8'h00;
      13'd7521: x = 8'h00;
      13'd7522: x = 8'h00;
      13'd7523: x = 8'h00;
      13'd7524: x = 8'h00;
      13'd7525: x = 8'h00;
      13'd7526: x = 8'h00;
      13'd7527: x = 8'h00;
      13'd7528: x = 8'h00;
      13'd7529: x = 8'h00;
      13'd7530: x = 8'h00;
      13'd7531: x = 8'h00;
      13'd7532: x = 8'h00;
      13'd7533: x = 8'h00;
      13'd7534: x = 8'h00;
      13'd7535: x = 8'h00;
      13'd7536: x = 8'h00;
      13'd7537: x = 8'h00;
      13'd7538: x = 8'h00;
      13'd7539: x = 8'h00;
      13'd7540: x = 8'h00;
      13'd7541: x = 8'h00;
      13'd7542: x = 8'h00;
      13'd7543: x = 8'h00;
      13'd7544: x = 8'h00;
      13'd7545: x = 8'h00;
      13'd7546: x = 8'h00;
      13'd7547: x = 8'h00;
      13'd7548: x = 8'h00;
      13'd7549: x = 8'h00;
      13'd7550: x = 8'h00;
      13'd7551: x = 8'h00;
      13'd7552: x = 8'h00;
      13'd7553: x = 8'h00;
      13'd7554: x = 8'h00;
      13'd7555: x = 8'h00;
      13'd7556: x = 8'h00;
      13'd7557: x = 8'h00;
      13'd7558: x = 8'h00;
      13'd7559: x = 8'h00;
      13'd7560: x = 8'h00;
      13'd7561: x = 8'h00;
      13'd7562: x = 8'h00;
      13'd7563: x = 8'h00;
      13'd7564: x = 8'h00;
      13'd7565: x = 8'h00;
      13'd7566: x = 8'h00;
      13'd7567: x = 8'h00;
      13'd7568: x = 8'h00;
      13'd7569: x = 8'h00;
      13'd7570: x = 8'h00;
      13'd7571: x = 8'h00;
      13'd7572: x = 8'h00;
      13'd7573: x = 8'h00;
      13'd7574: x = 8'h00;
      13'd7575: x = 8'h00;
      13'd7576: x = 8'h00;
      13'd7577: x = 8'h00;
      13'd7578: x = 8'h00;
      13'd7579: x = 8'h00;
      13'd7580: x = 8'h00;
      13'd7581: x = 8'h00;
      13'd7582: x = 8'h00;
      13'd7583: x = 8'h00;
      13'd7584: x = 8'h00;
      13'd7585: x = 8'h00;
      13'd7586: x = 8'h00;
      13'd7587: x = 8'h00;
      13'd7588: x = 8'h00;
      13'd7589: x = 8'h00;
      13'd7590: x = 8'h00;
      13'd7591: x = 8'h00;
      13'd7592: x = 8'h00;
      13'd7593: x = 8'h00;
      13'd7594: x = 8'h00;
      13'd7595: x = 8'h00;
      13'd7596: x = 8'h00;
      13'd7597: x = 8'h00;
      13'd7598: x = 8'h00;
      13'd7599: x = 8'h00;
      13'd7600: x = 8'h00;
      13'd7601: x = 8'h00;
      13'd7602: x = 8'h00;
      13'd7603: x = 8'h00;
      13'd7604: x = 8'h00;
      13'd7605: x = 8'h00;
      13'd7606: x = 8'h00;
      13'd7607: x = 8'h00;
      13'd7608: x = 8'h00;
      13'd7609: x = 8'h00;
      13'd7610: x = 8'h00;
      13'd7611: x = 8'h00;
      13'd7612: x = 8'h00;
      13'd7613: x = 8'h00;
      13'd7614: x = 8'h00;
      13'd7615: x = 8'h00;
      13'd7616: x = 8'h00;
      13'd7617: x = 8'h00;
      13'd7618: x = 8'h00;
      13'd7619: x = 8'h00;
      13'd7620: x = 8'h00;
      13'd7621: x = 8'h00;
      13'd7622: x = 8'h00;
      13'd7623: x = 8'h00;
      13'd7624: x = 8'h00;
      13'd7625: x = 8'h00;
      13'd7626: x = 8'h00;
      13'd7627: x = 8'h00;
      13'd7628: x = 8'h00;
      13'd7629: x = 8'h00;
      13'd7630: x = 8'h00;
      13'd7631: x = 8'h00;
      13'd7632: x = 8'h00;
      13'd7633: x = 8'h00;
      13'd7634: x = 8'h00;
      13'd7635: x = 8'h00;
      13'd7636: x = 8'h00;
      13'd7637: x = 8'h00;
      13'd7638: x = 8'h00;
      13'd7639: x = 8'h00;
      13'd7640: x = 8'h00;
      13'd7641: x = 8'h00;
      13'd7642: x = 8'h00;
      13'd7643: x = 8'h00;
      13'd7644: x = 8'h00;
      13'd7645: x = 8'h00;
      13'd7646: x = 8'h00;
      13'd7647: x = 8'h00;
      13'd7648: x = 8'h00;
      13'd7649: x = 8'h00;
      13'd7650: x = 8'h00;
      13'd7651: x = 8'h00;
      13'd7652: x = 8'h00;
      13'd7653: x = 8'h00;
      13'd7654: x = 8'h00;
      13'd7655: x = 8'h00;
      13'd7656: x = 8'h00;
      13'd7657: x = 8'h00;
      13'd7658: x = 8'h00;
      13'd7659: x = 8'h00;
      13'd7660: x = 8'h00;
      13'd7661: x = 8'h00;
      13'd7662: x = 8'h00;
      13'd7663: x = 8'h00;
      13'd7664: x = 8'h00;
      13'd7665: x = 8'h00;
      13'd7666: x = 8'h00;
      13'd7667: x = 8'h00;
      13'd7668: x = 8'h00;
      13'd7669: x = 8'h00;
      13'd7670: x = 8'h00;
      13'd7671: x = 8'h00;
      13'd7672: x = 8'h00;
      13'd7673: x = 8'h00;
      13'd7674: x = 8'h00;
      13'd7675: x = 8'h00;
      13'd7676: x = 8'h00;
      13'd7677: x = 8'h00;
      13'd7678: x = 8'h00;
      13'd7679: x = 8'h00;
      13'd7680: x = 8'h00;
      13'd7681: x = 8'h00;
      13'd7682: x = 8'h00;
      13'd7683: x = 8'h00;
      13'd7684: x = 8'h00;
      13'd7685: x = 8'h00;
      13'd7686: x = 8'h00;
      13'd7687: x = 8'h00;
      13'd7688: x = 8'h00;
      13'd7689: x = 8'h00;
      13'd7690: x = 8'h00;
      13'd7691: x = 8'h00;
      13'd7692: x = 8'h00;
      13'd7693: x = 8'h00;
      13'd7694: x = 8'h00;
      13'd7695: x = 8'h00;
      13'd7696: x = 8'h00;
      13'd7697: x = 8'h00;
      13'd7698: x = 8'h00;
      13'd7699: x = 8'h00;
      13'd7700: x = 8'h00;
      13'd7701: x = 8'h00;
      13'd7702: x = 8'h00;
      13'd7703: x = 8'h00;
      13'd7704: x = 8'h00;
      13'd7705: x = 8'h00;
      13'd7706: x = 8'h00;
      13'd7707: x = 8'h00;
      13'd7708: x = 8'h00;
      13'd7709: x = 8'h00;
      13'd7710: x = 8'h00;
      13'd7711: x = 8'h00;
      13'd7712: x = 8'h00;
      13'd7713: x = 8'h00;
      13'd7714: x = 8'h00;
      13'd7715: x = 8'h00;
      13'd7716: x = 8'h00;
      13'd7717: x = 8'h00;
      13'd7718: x = 8'h00;
      13'd7719: x = 8'h00;
      13'd7720: x = 8'h00;
      13'd7721: x = 8'h00;
      13'd7722: x = 8'h00;
      13'd7723: x = 8'h00;
      13'd7724: x = 8'h00;
      13'd7725: x = 8'h00;
      13'd7726: x = 8'h00;
      13'd7727: x = 8'h00;
      13'd7728: x = 8'h00;
      13'd7729: x = 8'h00;
      13'd7730: x = 8'h00;
      13'd7731: x = 8'h00;
      13'd7732: x = 8'h00;
      13'd7733: x = 8'h00;
      13'd7734: x = 8'h00;
      13'd7735: x = 8'h00;
      13'd7736: x = 8'h00;
      13'd7737: x = 8'h00;
      13'd7738: x = 8'h00;
      13'd7739: x = 8'h00;
      13'd7740: x = 8'h00;
      13'd7741: x = 8'h00;
      13'd7742: x = 8'h00;
      13'd7743: x = 8'h00;
      13'd7744: x = 8'h00;
      13'd7745: x = 8'h00;
      13'd7746: x = 8'h00;
      13'd7747: x = 8'h00;
      13'd7748: x = 8'h00;
      13'd7749: x = 8'h00;
      13'd7750: x = 8'h00;
      13'd7751: x = 8'h00;
      13'd7752: x = 8'h00;
      13'd7753: x = 8'h00;
      13'd7754: x = 8'h00;
      13'd7755: x = 8'h00;
      13'd7756: x = 8'h00;
      13'd7757: x = 8'h00;
      13'd7758: x = 8'h00;
      13'd7759: x = 8'h00;
      13'd7760: x = 8'h00;
      13'd7761: x = 8'h00;
      13'd7762: x = 8'h00;
      13'd7763: x = 8'h00;
      13'd7764: x = 8'h00;
      13'd7765: x = 8'h00;
      13'd7766: x = 8'h00;
      13'd7767: x = 8'h00;
      13'd7768: x = 8'h00;
      13'd7769: x = 8'h00;
      13'd7770: x = 8'h00;
      13'd7771: x = 8'h00;
      13'd7772: x = 8'h00;
      13'd7773: x = 8'h00;
      13'd7774: x = 8'h00;
      13'd7775: x = 8'h00;
      13'd7776: x = 8'h00;
      13'd7777: x = 8'h00;
      13'd7778: x = 8'h00;
      13'd7779: x = 8'h00;
      13'd7780: x = 8'h00;
      13'd7781: x = 8'h00;
      13'd7782: x = 8'h00;
      13'd7783: x = 8'h00;
      13'd7784: x = 8'h00;
      13'd7785: x = 8'h00;
      13'd7786: x = 8'h00;
      13'd7787: x = 8'h00;
      13'd7788: x = 8'h00;
      13'd7789: x = 8'h00;
      13'd7790: x = 8'h00;
      13'd7791: x = 8'h00;
      13'd7792: x = 8'h00;
      13'd7793: x = 8'h00;
      13'd7794: x = 8'h00;
      13'd7795: x = 8'h00;
      13'd7796: x = 8'h00;
      13'd7797: x = 8'h00;
      13'd7798: x = 8'h00;
      13'd7799: x = 8'h00;
      13'd7800: x = 8'h00;
      13'd7801: x = 8'h00;
      13'd7802: x = 8'h00;
      13'd7803: x = 8'h00;
      13'd7804: x = 8'h00;
      13'd7805: x = 8'h00;
      13'd7806: x = 8'h00;
      13'd7807: x = 8'h00;
      13'd7808: x = 8'h00;
      13'd7809: x = 8'h00;
      13'd7810: x = 8'h00;
      13'd7811: x = 8'h00;
      13'd7812: x = 8'h00;
      13'd7813: x = 8'h00;
      13'd7814: x = 8'h00;
      13'd7815: x = 8'h00;
      13'd7816: x = 8'h00;
      13'd7817: x = 8'h00;
      13'd7818: x = 8'h00;
      13'd7819: x = 8'h00;
      13'd7820: x = 8'h00;
      13'd7821: x = 8'h00;
      13'd7822: x = 8'h00;
      13'd7823: x = 8'h00;
      13'd7824: x = 8'h00;
      13'd7825: x = 8'h00;
      13'd7826: x = 8'h00;
      13'd7827: x = 8'h00;
      13'd7828: x = 8'h00;
      13'd7829: x = 8'h00;
      13'd7830: x = 8'h00;
      13'd7831: x = 8'h00;
      13'd7832: x = 8'h00;
      13'd7833: x = 8'h00;
      13'd7834: x = 8'h00;
      13'd7835: x = 8'h00;
      13'd7836: x = 8'h00;
      13'd7837: x = 8'h00;
      13'd7838: x = 8'h00;
      13'd7839: x = 8'h00;
      13'd7840: x = 8'h00;
      13'd7841: x = 8'h00;
      13'd7842: x = 8'h00;
      13'd7843: x = 8'h00;
      13'd7844: x = 8'h00;
      13'd7845: x = 8'h00;
      13'd7846: x = 8'h00;
      13'd7847: x = 8'h00;
      13'd7848: x = 8'h00;
      13'd7849: x = 8'h00;
      13'd7850: x = 8'h00;
      13'd7851: x = 8'h00;
      13'd7852: x = 8'h00;
      13'd7853: x = 8'h00;
      13'd7854: x = 8'h00;
      13'd7855: x = 8'h00;
      13'd7856: x = 8'h00;
      13'd7857: x = 8'h00;
      13'd7858: x = 8'h00;
      13'd7859: x = 8'h00;
      13'd7860: x = 8'h00;
      13'd7861: x = 8'h00;
      13'd7862: x = 8'h00;
      13'd7863: x = 8'h00;
      13'd7864: x = 8'h00;
      13'd7865: x = 8'h00;
      13'd7866: x = 8'h00;
      13'd7867: x = 8'h00;
      13'd7868: x = 8'h00;
      13'd7869: x = 8'h00;
      13'd7870: x = 8'h00;
      13'd7871: x = 8'h00;
      13'd7872: x = 8'h00;
      13'd7873: x = 8'h00;
      13'd7874: x = 8'h00;
      13'd7875: x = 8'h00;
      13'd7876: x = 8'h00;
      13'd7877: x = 8'h00;
      13'd7878: x = 8'h00;
      13'd7879: x = 8'h00;
      13'd7880: x = 8'h00;
      13'd7881: x = 8'h00;
      13'd7882: x = 8'h00;
      13'd7883: x = 8'h00;
      13'd7884: x = 8'h00;
      13'd7885: x = 8'h00;
      13'd7886: x = 8'h00;
      13'd7887: x = 8'h00;
      13'd7888: x = 8'h00;
      13'd7889: x = 8'h00;
      13'd7890: x = 8'h00;
      13'd7891: x = 8'h00;
      13'd7892: x = 8'h00;
      13'd7893: x = 8'h00;
      13'd7894: x = 8'h00;
      13'd7895: x = 8'h00;
      13'd7896: x = 8'h00;
      13'd7897: x = 8'h00;
      13'd7898: x = 8'h00;
      13'd7899: x = 8'h00;
      13'd7900: x = 8'h00;
      13'd7901: x = 8'h00;
      13'd7902: x = 8'h00;
      13'd7903: x = 8'h00;
      13'd7904: x = 8'h00;
      13'd7905: x = 8'h00;
      13'd7906: x = 8'h00;
      13'd7907: x = 8'h00;
      13'd7908: x = 8'h00;
      13'd7909: x = 8'h00;
      13'd7910: x = 8'h00;
      13'd7911: x = 8'h00;
      13'd7912: x = 8'h00;
      13'd7913: x = 8'h00;
      13'd7914: x = 8'h00;
      13'd7915: x = 8'h00;
      13'd7916: x = 8'h00;
      13'd7917: x = 8'h00;
      13'd7918: x = 8'h00;
      13'd7919: x = 8'h00;
      13'd7920: x = 8'h00;
      13'd7921: x = 8'h00;
      13'd7922: x = 8'h00;
      13'd7923: x = 8'h00;
      13'd7924: x = 8'h00;
      13'd7925: x = 8'h00;
      13'd7926: x = 8'h00;
      13'd7927: x = 8'h00;
      13'd7928: x = 8'h00;
      13'd7929: x = 8'h00;
      13'd7930: x = 8'h00;
      13'd7931: x = 8'h00;
      13'd7932: x = 8'h00;
      13'd7933: x = 8'h00;
      13'd7934: x = 8'h00;
      13'd7935: x = 8'h00;
      13'd7936: x = 8'hd8;
      13'd7937: x = 8'h58;
      13'd7938: x = 8'ha0;
      13'd7939: x = 8'h7f;
      13'd7940: x = 8'h8c;
      13'd7941: x = 8'h12;
      13'd7942: x = 8'hd0;
      13'd7943: x = 8'ha9;
      13'd7944: x = 8'ha7;
      13'd7945: x = 8'h8d;
      13'd7946: x = 8'h11;
      13'd7947: x = 8'hd0;
      13'd7948: x = 8'h8d;
      13'd7949: x = 8'h13;
      13'd7950: x = 8'hd0;
      13'd7951: x = 8'hc9;
      13'd7952: x = 8'hdf;
      13'd7953: x = 8'hf0;
      13'd7954: x = 8'h13;
      13'd7955: x = 8'hc9;
      13'd7956: x = 8'h9b;
      13'd7957: x = 8'hf0;
      13'd7958: x = 8'h03;
      13'd7959: x = 8'hc8;
      13'd7960: x = 8'h10;
      13'd7961: x = 8'h0f;
      13'd7962: x = 8'ha9;
      13'd7963: x = 8'hdc;
      13'd7964: x = 8'h20;
      13'd7965: x = 8'hef;
      13'd7966: x = 8'hff;
      13'd7967: x = 8'ha9;
      13'd7968: x = 8'h8d;
      13'd7969: x = 8'h20;
      13'd7970: x = 8'hef;
      13'd7971: x = 8'hff;
      13'd7972: x = 8'ha0;
      13'd7973: x = 8'h01;
      13'd7974: x = 8'h88;
      13'd7975: x = 8'h30;
      13'd7976: x = 8'hf6;
      13'd7977: x = 8'had;
      13'd7978: x = 8'h11;
      13'd7979: x = 8'hd0;
      13'd7980: x = 8'h10;
      13'd7981: x = 8'hfb;
      13'd7982: x = 8'had;
      13'd7983: x = 8'h10;
      13'd7984: x = 8'hd0;
      13'd7985: x = 8'h99;
      13'd7986: x = 8'h00;
      13'd7987: x = 8'h02;
      13'd7988: x = 8'h20;
      13'd7989: x = 8'hef;
      13'd7990: x = 8'hff;
      13'd7991: x = 8'hc9;
      13'd7992: x = 8'h8d;
      13'd7993: x = 8'hd0;
      13'd7994: x = 8'hd4;
      13'd7995: x = 8'ha0;
      13'd7996: x = 8'hff;
      13'd7997: x = 8'ha9;
      13'd7998: x = 8'h00;
      13'd7999: x = 8'haa;
      13'd8000: x = 8'h0a;
      13'd8001: x = 8'h85;
      13'd8002: x = 8'h2b;
      13'd8003: x = 8'hc8;
      13'd8004: x = 8'hb9;
      13'd8005: x = 8'h00;
      13'd8006: x = 8'h02;
      13'd8007: x = 8'hc9;
      13'd8008: x = 8'h8d;
      13'd8009: x = 8'hf0;
      13'd8010: x = 8'hd4;
      13'd8011: x = 8'hc9;
      13'd8012: x = 8'hae;
      13'd8013: x = 8'h90;
      13'd8014: x = 8'hf4;
      13'd8015: x = 8'hf0;
      13'd8016: x = 8'hf0;
      13'd8017: x = 8'hc9;
      13'd8018: x = 8'hba;
      13'd8019: x = 8'hf0;
      13'd8020: x = 8'heb;
      13'd8021: x = 8'hc9;
      13'd8022: x = 8'hd2;
      13'd8023: x = 8'hf0;
      13'd8024: x = 8'h3b;
      13'd8025: x = 8'h86;
      13'd8026: x = 8'h28;
      13'd8027: x = 8'h86;
      13'd8028: x = 8'h29;
      13'd8029: x = 8'h84;
      13'd8030: x = 8'h2a;
      13'd8031: x = 8'hb9;
      13'd8032: x = 8'h00;
      13'd8033: x = 8'h02;
      13'd8034: x = 8'h49;
      13'd8035: x = 8'hb0;
      13'd8036: x = 8'hc9;
      13'd8037: x = 8'h0a;
      13'd8038: x = 8'h90;
      13'd8039: x = 8'h06;
      13'd8040: x = 8'h69;
      13'd8041: x = 8'h88;
      13'd8042: x = 8'hc9;
      13'd8043: x = 8'hfa;
      13'd8044: x = 8'h90;
      13'd8045: x = 8'h11;
      13'd8046: x = 8'h0a;
      13'd8047: x = 8'h0a;
      13'd8048: x = 8'h0a;
      13'd8049: x = 8'h0a;
      13'd8050: x = 8'ha2;
      13'd8051: x = 8'h04;
      13'd8052: x = 8'h0a;
      13'd8053: x = 8'h26;
      13'd8054: x = 8'h28;
      13'd8055: x = 8'h26;
      13'd8056: x = 8'h29;
      13'd8057: x = 8'hca;
      13'd8058: x = 8'hd0;
      13'd8059: x = 8'hf8;
      13'd8060: x = 8'hc8;
      13'd8061: x = 8'hd0;
      13'd8062: x = 8'he0;
      13'd8063: x = 8'hc4;
      13'd8064: x = 8'h2a;
      13'd8065: x = 8'hf0;
      13'd8066: x = 8'h97;
      13'd8067: x = 8'h24;
      13'd8068: x = 8'h2b;
      13'd8069: x = 8'h50;
      13'd8070: x = 8'h10;
      13'd8071: x = 8'ha5;
      13'd8072: x = 8'h28;
      13'd8073: x = 8'h81;
      13'd8074: x = 8'h26;
      13'd8075: x = 8'he6;
      13'd8076: x = 8'h26;
      13'd8077: x = 8'hd0;
      13'd8078: x = 8'hb5;
      13'd8079: x = 8'he6;
      13'd8080: x = 8'h27;
      13'd8081: x = 8'h4c;
      13'd8082: x = 8'h44;
      13'd8083: x = 8'hff;
      13'd8084: x = 8'h6c;
      13'd8085: x = 8'h24;
      13'd8086: x = 8'h00;
      13'd8087: x = 8'h30;
      13'd8088: x = 8'h2b;
      13'd8089: x = 8'ha2;
      13'd8090: x = 8'h02;
      13'd8091: x = 8'hb5;
      13'd8092: x = 8'h27;
      13'd8093: x = 8'h95;
      13'd8094: x = 8'h25;
      13'd8095: x = 8'h95;
      13'd8096: x = 8'h23;
      13'd8097: x = 8'hca;
      13'd8098: x = 8'hd0;
      13'd8099: x = 8'hf7;
      13'd8100: x = 8'hd0;
      13'd8101: x = 8'h14;
      13'd8102: x = 8'ha9;
      13'd8103: x = 8'h8d;
      13'd8104: x = 8'h20;
      13'd8105: x = 8'hef;
      13'd8106: x = 8'hff;
      13'd8107: x = 8'ha5;
      13'd8108: x = 8'h25;
      13'd8109: x = 8'h20;
      13'd8110: x = 8'hdc;
      13'd8111: x = 8'hff;
      13'd8112: x = 8'ha5;
      13'd8113: x = 8'h24;
      13'd8114: x = 8'h20;
      13'd8115: x = 8'hdc;
      13'd8116: x = 8'hff;
      13'd8117: x = 8'ha9;
      13'd8118: x = 8'hba;
      13'd8119: x = 8'h20;
      13'd8120: x = 8'hef;
      13'd8121: x = 8'hff;
      13'd8122: x = 8'ha9;
      13'd8123: x = 8'ha0;
      13'd8124: x = 8'h20;
      13'd8125: x = 8'hef;
      13'd8126: x = 8'hff;
      13'd8127: x = 8'ha1;
      13'd8128: x = 8'h24;
      13'd8129: x = 8'h20;
      13'd8130: x = 8'hdc;
      13'd8131: x = 8'hff;
      13'd8132: x = 8'h86;
      13'd8133: x = 8'h2b;
      13'd8134: x = 8'ha5;
      13'd8135: x = 8'h24;
      13'd8136: x = 8'hc5;
      13'd8137: x = 8'h28;
      13'd8138: x = 8'ha5;
      13'd8139: x = 8'h25;
      13'd8140: x = 8'he5;
      13'd8141: x = 8'h29;
      13'd8142: x = 8'hb0;
      13'd8143: x = 8'hc1;
      13'd8144: x = 8'he6;
      13'd8145: x = 8'h24;
      13'd8146: x = 8'hd0;
      13'd8147: x = 8'h02;
      13'd8148: x = 8'he6;
      13'd8149: x = 8'h25;
      13'd8150: x = 8'ha5;
      13'd8151: x = 8'h24;
      13'd8152: x = 8'h29;
      13'd8153: x = 8'h07;
      13'd8154: x = 8'h10;
      13'd8155: x = 8'hc8;
      13'd8156: x = 8'h48;
      13'd8157: x = 8'h4a;
      13'd8158: x = 8'h4a;
      13'd8159: x = 8'h4a;
      13'd8160: x = 8'h4a;
      13'd8161: x = 8'h20;
      13'd8162: x = 8'he5;
      13'd8163: x = 8'hff;
      13'd8164: x = 8'h68;
      13'd8165: x = 8'h29;
      13'd8166: x = 8'h0f;
      13'd8167: x = 8'h09;
      13'd8168: x = 8'hb0;
      13'd8169: x = 8'hc9;
      13'd8170: x = 8'hba;
      13'd8171: x = 8'h90;
      13'd8172: x = 8'h02;
      13'd8173: x = 8'h69;
      13'd8174: x = 8'h06;
      13'd8175: x = 8'h2c;
      13'd8176: x = 8'h12;
      13'd8177: x = 8'hd0;
      13'd8178: x = 8'h30;
      13'd8179: x = 8'hfb;
      13'd8180: x = 8'h8d;
      13'd8181: x = 8'h12;
      13'd8182: x = 8'hd0;
      13'd8183: x = 8'h60;
      13'd8184: x = 8'h00;
      13'd8185: x = 8'h00;
      13'd8186: x = 8'h00;
      13'd8187: x = 8'h0f;
      13'd8188: x = 8'h00;
      13'd8189: x = 8'hff;
      13'd8190: x = 8'h00;
      13'd8191: x = 8'h00;
    endcase

endmodule
