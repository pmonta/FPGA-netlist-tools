* SPICE3 file created from 4004.ext - technology: 4004-nmos-buried-stacked

.option scale=0.001u

M1000 vss N0770 N0385 vss efet w=89900 l=11600
M1001 vss vss test vss efet w=119625 l=15225
M1002 reset vss vss vss efet w=118175 l=15225
M1003 vss N0754 N0761 vss efet w=26100 l=13050
M1004 vss PC0_11 N0785 vss efet w=30450 l=12325
M1005 N0785 N0406 N0770 vss efet w=26100 l=13050
M1006 vss N0301 N0754 vss efet w=21750 l=11600
M1007 N0761 N0301 N0753 vss efet w=78300 l=11600
M1008 N0754 vcc vcc vss efet w=7250 l=69600
M1009 N0754 N0289 vss vss efet w=23925 l=13775
M1010 vcc vcc N0761 vss efet w=8700 l=30450
M1011 N0753 N0289 vss vss efet w=136300 l=20300
M1012 D3 RADB1 N0386 vss efet w=44225 l=13775
M1013 N0385 RADB2 D3 vss efet w=49300 l=12325
M1014 N0770 WADB2 N0761 vss efet w=14500 l=13050
M1015 vss N0289 N0311 vss efet w=15225 l=12325
M1016 vcc N0325 N0301 vss efet w=9425 l=13775
M1017 N0289 M12_M22_CLK1__M11_M12_ D3 vss efet w=21025 l=12325
M1018 N0387 RADB0 D3 vss efet w=44950 l=10875
M1019 N0290 M12_M22_CLK1__M11_M12_ D2 vss efet w=20300 l=11600
M1020 N0311 N0290 N0312 vss efet w=14500 l=12325
M1021 N0301 N0290 N0302 vss efet w=26100 l=11600
M1022 vss N0290 N0755 vss efet w=123250 l=11600
M1023 vss N0740 sync vss efet w=1224525 l=10875
M1025 vcc vcc S00531 vss efet w=5800 l=13050
M1026 vcc S00531 N0740 vss efet w=10150 l=13050
M1028 vcc S00536 N0738 vss efet w=11600 l=11600
M1029 vcc vcc S00536 vss efet w=6525 l=13775
M1030 sync N0738 vcc vss efet w=679325 l=13050
M1031 N0388 RADB0 D2 vss efet w=42050 l=11600
M1032 vcc N0325 N0298 vss efet w=13050 l=14500
M1033 N0762 N0298 N0755 vss efet w=68150 l=11600
M1034 vss N0290 N0756 vss efet w=23200 l=10150
M1035 N0756 vcc vcc vss efet w=7250 l=68150
M1036 vcc vcc N0762 vss efet w=7250 l=27550
M1037 N0756 N0298 vss vss efet w=23925 l=12325
M1038 N0762 N0756 vss vss efet w=26100 l=11600
M1039 vss N0758 N0763 vss efet w=26100 l=11600
M1040 vss N0293 N0758 vss efet w=23925 l=11600
M1041 N0763 N0293 N0757 vss efet w=70325 l=12325
M1042 N0758 vcc vcc vss efet w=7975 l=67425
M1043 N0758 N0291 vss vss efet w=23200 l=11600
M1044 vcc vcc N0763 vss efet w=7975 l=29725
M1045 N0757 N0291 vss vss efet w=125425 l=12325
M1046 N0298 N0291 N0299 vss efet w=23200 l=18850
M1047 N0312 N0291 N0313 vss efet w=13050 l=11600
M1048 N0302 N0291 N0303 vss efet w=23200 l=11600
M1049 vcc N0325 N0293 vss efet w=9425 l=13775
M1050 N0291 M12_M22_CLK1__M11_M12_ D1 vss efet w=20300 l=11600
M1051 N0761 WADB1 N0774 vss efet w=14500 l=13775
M1052 N0778 WADB0 N0761 vss efet w=14500 l=11600
M1053 N0779 WADB0 N0762 vss efet w=17400 l=10150
M1054 N0762 WADB1 N0775 vss efet w=15950 l=13050
M1055 D2 RADB1 N0389 vss efet w=44225 l=12325
M1056 N0390 RADB2 D2 vss efet w=47125 l=10875
M1057 D1 RADB1 N0392 vss efet w=44225 l=14500
M1058 N0391 RADB2 D1 vss efet w=53650 l=10150
M1059 N0393 RADB0 D1 vss efet w=43500 l=11600
M1060 N0313 N0292 N0305 vss efet w=13050 l=11600
M1061 N0303 N0292 N0294 vss efet w=23200 l=11600
M1062 N0299 N0292 N0294 vss efet w=17400 l=11600
M1063 N0293 N0292 N0294 vss efet w=8700 l=11600
M1064 N0292 M12_M22_CLK1__M11_M12_ D0 vss efet w=23200 l=12325
M1065 vss N0292 N0759 vss efet w=125425 l=12325
M1066 N0305 N0325 vcc vss efet w=7975 l=12325
M1067 N0394 RADB0 D0 vss efet w=43500 l=13775
M1068 vcc N0325 N0752 vss efet w=10875 l=14500
M1069 N0764 N0752 N0759 vss efet w=69600 l=11600
M1070 vss N0292 N0760 vss efet w=29000 l=11600
M1071 N0760 vcc vcc vss efet w=7975 l=67425
M1072 vcc vcc N0764 vss efet w=7250 l=27550
M1073 vss N0307 N0294 vss efet w=31900 l=13050
M1074 N0760 N0752 vss vss efet w=21750 l=10150
M1075 N0752 N0307 vss vss efet w=14500 l=11600
M1076 N0764 N0760 vss vss efet w=27550 l=10150
M1077 vss N0738 N0740 vss efet w=101500 l=13050
M1078 N0305 N0307 N0306 vss efet w=14500 l=11600
M1079 vss N0295 N0738 vss efet w=112375 l=13775
M1080 vss PC2_11 N0821 vss efet w=26100 l=14500
M1081 N0806 PC1_11 vss vss efet w=19575 l=10875
M1082 N0770 N0424 N0806 vss efet w=26825 l=12325
M1083 N0821 N0434 N0770 vss efet w=26100 l=12325
M1084 N0770 N0444 N0834 vss efet w=28275 l=12325
M1085 N0834 PC3_11 vss vss efet w=23200 l=11600
M1086 N0386 N0774 vss vss efet w=72500 l=16675
M1087 N0385 N0381 PC0_11 vss efet w=6525 l=12325
M1088 PC1_11 N0410 N0385 vss efet w=7975 l=10875
M1089 N0386 N0381 PC0_7 vss efet w=6525 l=12325
M1090 PC1_7 N0410 N0386 vss efet w=5800 l=10150
M1091 N0786 N0406 N0774 vss efet w=27550 l=11600
M1092 vss PC0_7 N0786 vss efet w=25375 l=15225
M1093 N0385 N0426 PC2_11 vss efet w=6525 l=12325
M1094 PC3_11 N0439 N0385 vss efet w=5800 l=11600
M1095 N0386 N0426 PC2_7 vss efet w=6525 l=12325
M1096 vss N0778 N0387 vss efet w=72500 l=13775
M1097 N0787 N0406 N0778 vss efet w=24650 l=10875
M1098 vss PC0_3 N0787 vss efet w=24650 l=15225
M1099 N0807 PC1_7 vss vss efet w=22475 l=13775
M1100 N0774 N0424 N0807 vss efet w=27550 l=11600
M1101 N0822 N0434 N0774 vss efet w=26825 l=10875
M1102 vss PC2_7 N0822 vss efet w=23925 l=12325
M1103 N0388 N0779 vss vss efet w=71050 l=13775
M1104 N0387 N0381 PC0_3 vss efet w=7975 l=12325
M1105 N0808 PC1_3 vss vss efet w=23925 l=15225
M1106 PC3_7 N0439 N0386 vss efet w=5800 l=13050
M1107 vcc __INH__X11_X31_CLK1 N0770 vss efet w=8700 l=11600
M1108 D0 M12_M22_CLK1__M11_M12_ N0497 vss efet w=14500 l=13050
M1109 N0862 WRAB1 N0866 vss efet w=17400 l=13050
M1110 vss N0866 N0531 vss efet w=63800 l=11600
M1111 vcc vcc N0385 vss efet w=6525 l=31175
M1112 vss N0497 N0862 vss efet w=109475 l=12325
M1113 vcc vcc N0386 vss efet w=7250 l=30450
M1114 vss PC2_3 N0823 vss efet w=25375 l=12325
M1115 N0778 N0424 N0808 vss efet w=25375 l=11600
M1116 N0823 N0434 N0778 vss efet w=26825 l=10875
M1117 N0835 PC3_7 vss vss efet w=23925 l=13775
M1118 N0774 N0444 N0835 vss efet w=26825 l=10875
M1119 vcc __INH__X11_X31_CLK1 N0774 vss efet w=9425 l=13050
M1120 D0 RRAB1 N0531 vss efet w=46400 l=11600
M1121 N0532 RRAB0 D0 vss efet w=45675 l=13050
M1122 N0862 vcc vcc vss efet w=7975 l=22475
M1123 N0836 PC3_3 vss vss efet w=23925 l=13775
M1124 N0778 N0444 N0836 vss efet w=28275 l=10875
M1125 PC1_3 N0410 N0387 vss efet w=6525 l=10150
M1126 N0388 N0381 PC0_2 vss efet w=5800 l=10150
M1127 PC1_2 N0410 N0388 vss efet w=5800 l=10150
M1128 N0788 N0406 N0779 vss efet w=28275 l=10875
M1129 vss PC0_2 N0788 vss efet w=24650 l=13050
M1130 N0387 N0426 PC2_3 vss efet w=6525 l=12325
M1131 vcc __INH__X11_X31_CLK1 N0778 vss efet w=9425 l=13775
M1132 N0863 vcc vcc vss efet w=7975 l=21025
M1133 PC3_3 N0439 N0387 vss efet w=5800 l=11600
M1134 N0388 N0426 PC2_2 vss efet w=6525 l=10150
M1135 PC3_2 N0439 N0388 vss efet w=5800 l=11600
M1136 vss N0775 N0389 vss efet w=63800 l=11600
M1137 vss N0771 N0390 vss efet w=68875 l=13775
M1138 N0771 WADB2 N0762 vss efet w=13050 l=11600
M1139 N0789 N0406 N0775 vss efet w=24650 l=10875
M1140 vss PC0_6 N0789 vss efet w=24650 l=14500
M1141 N0809 PC1_2 vss vss efet w=23925 l=13775
M1142 N0779 N0424 N0809 vss efet w=26100 l=11600
M1143 N0824 N0434 N0779 vss efet w=26825 l=10875
M1144 vss PC2_2 N0824 vss efet w=24650 l=11600
M1145 vss N0498 N0863 vss efet w=114550 l=11600
M1146 vcc vcc N0387 vss efet w=7250 l=31900
M1147 vcc vcc N0388 vss efet w=7975 l=29725
M1148 N0837 PC3_2 vss vss efet w=23925 l=18125
M1149 N0810 PC1_6 vss vss efet w=22475 l=15225
M1150 vss PC2_6 N0825 vss efet w=23925 l=12325
M1151 N0775 N0424 N0810 vss efet w=26825 l=10875
M1152 N0825 N0434 N0775 vss efet w=25375 l=10875
M1153 N0779 N0444 N0837 vss efet w=26100 l=11600
M1154 vcc __INH__X11_X31_CLK1 N0779 vss efet w=8700 l=13050
M1155 D1 RRAB1 N0534 vss efet w=44950 l=11600
M1156 N0533 RRAB0 D1 vss efet w=46400 l=11600
M1157 N0880 WRAB0 N0862 vss efet w=13775 l=13050
M1158 N0532 N0880 vss vss efet w=59450 l=11600
M1159 N0903 N0543 N0866 vss efet w=24650 l=13050
M1160 vss R1_0 N0903 vss efet w=26100 l=14500
M1161 N0920 R3_0 vss vss efet w=24650 l=14500
M1162 N0866 N0565 N0920 vss efet w=24650 l=13050
M1163 N0929 N0581 N0866 vss efet w=26100 l=13050
M1164 vss R5_0 N0929 vss efet w=23925 l=13775
M1165 N0947 R7_0 vss vss efet w=25375 l=16675
M1166 N0866 N0591 N0947 vss efet w=24650 l=13775
M1167 N0956 N0616 N0866 vss efet w=26100 l=14500
M1168 vss R9_0 N0956 vss efet w=26825 l=19575
M1169 N0966 R11_0 vss vss efet w=25375 l=13775
M1170 N0531 N0529 R1_0 vss efet w=5800 l=11600
M1171 R3_0 N0544 N0531 vss efet w=5800 l=11600
M1172 N0531 N0569 R5_0 vss efet w=6525 l=12325
M1173 N0532 N0529 R0_0 vss efet w=5800 l=11600
M1174 R2_0 N0544 N0532 vss efet w=5800 l=11600
M1175 N0904 N0543 N0880 vss efet w=27550 l=13050
M1176 vss R0_0 N0904 vss efet w=24650 l=12325
M1177 R7_0 N0583 N0531 vss efet w=5800 l=11600
M1178 vss R0_1 N0905 vss efet w=23925 l=13775
M1179 N0498 M12_M22_CLK1__M11_M12_ D1 vss efet w=13050 l=11600
M1180 N0838 PC3_6 vss vss efet w=24650 l=16675
M1181 N0775 N0444 N0838 vss efet w=25375 l=10875
M1182 N0389 N0381 PC0_6 vss efet w=7975 l=12325
M1183 PC1_6 N0410 N0389 vss efet w=5800 l=12325
M1184 N0390 N0381 PC0_10 vss efet w=5800 l=10150
M1185 PC1_10 N0410 N0390 vss efet w=5800 l=10150
M1186 N0790 N0406 N0771 vss efet w=27550 l=10875
M1187 vss PC0_10 N0790 vss efet w=23925 l=12325
M1188 N0389 N0426 PC2_6 vss efet w=6525 l=10875
M1189 PC3_6 N0439 N0389 vss efet w=5800 l=10150
M1190 N0390 N0426 PC2_10 vss efet w=5800 l=10150
M1191 PC3_10 N0439 N0390 vss efet w=5800 l=10150
M1192 vss N0772 N0391 vss efet w=73225 l=12325
M1193 N0772 WADB2 N0763 vss efet w=14500 l=10875
M1194 N0763 WADB1 N0776 vss efet w=14500 l=13050
M1195 N0791 N0406 N0772 vss efet w=26825 l=10875
M1196 vss PC0_9 N0791 vss efet w=24650 l=13050
M1197 N0811 PC1_10 vss vss efet w=23200 l=14500
M1198 N0771 N0424 N0811 vss efet w=27550 l=11600
M1199 N0826 N0434 N0771 vss efet w=27550 l=11600
M1200 vss PC2_10 N0826 vss efet w=24650 l=11600
M1201 vcc __INH__X11_X31_CLK1 N0775 vss efet w=8700 l=11600
M1202 N0499 M12_M22_CLK1__M11_M12_ D2 vss efet w=14500 l=13050
M1203 N0780 WADB0 N0763 vss efet w=14500 l=13050
M1204 N0781 WADB0 N0764 vss efet w=15225 l=12325
M1205 N0392 N0776 vss vss efet w=65975 l=10875
M1206 N0391 N0381 PC0_9 vss efet w=6525 l=13050
M1207 N0812 PC1_9 vss vss efet w=23200 l=14500
M1208 vss PC2_9 N0827 vss efet w=26100 l=13050
M1209 N0772 N0424 N0812 vss efet w=25375 l=12325
M1210 N0827 N0434 N0772 vss efet w=26100 l=11600
M1211 N0839 PC3_10 vss vss efet w=24650 l=13050
M1212 N0771 N0444 N0839 vss efet w=26100 l=11600
M1213 vcc vcc N0389 vss efet w=6525 l=29725
M1214 D2 RRAB1 N0535 vss efet w=44225 l=12325
M1215 vss N0499 N0864 vss efet w=109475 l=10875
M1216 vcc vcc N0390 vss efet w=7975 l=28275
M1217 vcc __INH__X11_X31_CLK1 N0771 vss efet w=10150 l=11600
M1218 N0881 WRAB0 N0863 vss efet w=13050 l=13050
M1219 N0863 WRAB1 N0867 vss efet w=13050 l=11600
M1220 N0864 WRAB1 N0868 vss efet w=13050 l=11600
M1221 N0840 PC3_9 vss vss efet w=25375 l=13775
M1222 PC1_9 N0410 N0391 vss efet w=5800 l=11600
M1223 PC1_5 N0410 N0392 vss efet w=5800 l=13050
M1224 N0392 N0381 PC0_5 vss efet w=5800 l=11600
M1225 N0792 N0406 N0776 vss efet w=28275 l=10875
M1226 vss PC0_5 N0792 vss efet w=23925 l=12325
M1227 N0391 N0426 PC2_9 vss efet w=5800 l=10150
M1228 N0772 N0444 N0840 vss efet w=25375 l=12325
M1229 PC3_9 N0439 N0391 vss efet w=5800 l=10150
M1230 N0392 N0426 PC2_5 vss efet w=5800 l=10150
M1231 N0813 PC1_5 vss vss efet w=23925 l=12325
M1232 vss PC0_1 N0793 vss efet w=25375 l=13775
M1233 vss N0780 N0393 vss efet w=69600 l=11600
M1234 N0793 N0406 N0780 vss efet w=25375 l=10875
M1235 N0776 N0424 N0813 vss efet w=26825 l=10875
M1236 N0828 N0434 N0776 vss efet w=26100 l=11600
M1237 vss PC2_5 N0828 vss efet w=26100 l=11600
M1238 PC3_5 N0439 N0392 vss efet w=5800 l=11600
M1239 N0841 PC3_5 vss vss efet w=23925 l=13775
M1240 N0776 N0444 N0841 vss efet w=24650 l=11600
M1241 N0394 N0781 vss vss efet w=68150 l=13050
M1242 N0393 N0381 PC0_1 vss efet w=5800 l=11600
M1243 N0814 PC1_1 vss vss efet w=24650 l=13050
M1244 vss PC2_1 N0829 vss efet w=23925 l=12325
M1245 N0780 N0424 N0814 vss efet w=26100 l=11600
M1246 N0829 N0434 N0780 vss efet w=26100 l=11600
M1247 N0864 vcc vcc vss efet w=7250 l=20300
M1248 vcc __INH__X11_X31_CLK1 N0772 vss efet w=9425 l=13775
M1249 vcc vcc N0391 vss efet w=7975 l=28275
M1250 N0865 vcc vcc vss efet w=7975 l=20300
M1251 vss N0500 N0865 vss efet w=114550 l=13050
M1252 N0536 RRAB0 D2 vss efet w=44950 l=11600
M1253 vss N0881 N0533 vss efet w=59450 l=11600
M1254 N0534 N0867 vss vss efet w=60175 l=10875
M1255 N0905 N0543 N0881 vss efet w=26100 l=11600
M1256 N0921 R2_0 vss vss efet w=29000 l=14500
M1257 N0880 N0565 N0921 vss efet w=27550 l=11600
M1258 N0930 N0581 N0880 vss efet w=26100 l=13050
M1259 N0532 N0569 R4_0 vss efet w=5800 l=11600
M1260 vss R4_0 N0930 vss efet w=21750 l=13050
M1261 N0922 R2_1 vss vss efet w=26825 l=15225
M1262 N0533 N0529 R0_1 vss efet w=5800 l=11600
M1263 R6_0 N0583 N0532 vss efet w=5800 l=11600
M1264 N0948 R6_0 vss vss efet w=24650 l=15950
M1265 N0866 N0632 N0966 vss efet w=30450 l=13050
M1266 N0975 N0645 N0866 vss efet w=27550 l=13050
M1267 vss R13_0 N0975 vss efet w=26825 l=18850
M1268 N0984 R15_0 vss vss efet w=27550 l=13050
M1269 N0866 N0657 N0984 vss efet w=29000 l=13775
M1270 N0880 N0591 N0948 vss efet w=26825 l=13775
M1271 N0531 N0598 R9_0 vss efet w=5800 l=13050
M1272 R11_0 N0619 N0531 vss efet w=7975 l=12325
M1273 N0532 N0598 R8_0 vss efet w=7250 l=13050
M1274 vss R8_0 N0957 vss efet w=21750 l=14500
M1275 R10_0 N0619 N0532 vss efet w=6525 l=12325
M1276 N0957 N0616 N0880 vss efet w=24650 l=11600
M1277 vss R4_1 N0931 vss efet w=23200 l=15225
M1278 N0881 N0565 N0922 vss efet w=28275 l=10875
M1279 N0931 N0581 N0881 vss efet w=25375 l=10875
M1280 N0531 N0634 R13_0 vss efet w=5800 l=13050
M1281 R15_0 N0647 N0531 vss efet w=5800 l=14500
M1282 N0532 N0634 R12_0 vss efet w=7250 l=13775
M1283 N0949 R6_1 vss vss efet w=25375 l=16675
M1284 N0881 N0591 N0949 vss efet w=27550 l=13050
M1285 R2_1 N0544 N0533 vss efet w=5800 l=11600
M1286 N0534 N0529 R1_1 vss efet w=5800 l=11600
M1287 R3_1 N0544 N0534 vss efet w=5800 l=11600
M1288 N0906 N0543 N0867 vss efet w=27550 l=11600
M1289 vss R1_1 N0906 vss efet w=23200 l=13050
M1290 N0533 N0569 R4_1 vss efet w=6525 l=10875
M1291 N0958 N0616 N0881 vss efet w=25375 l=13050
M1292 vss R8_1 N0958 vss efet w=22475 l=13775
M1293 N0967 R10_0 vss vss efet w=26825 l=13775
M1294 N0880 N0632 N0967 vss efet w=25375 l=12325
M1295 N0976 N0645 N0880 vss efet w=25375 l=12325
M1296 vss R12_0 N0976 vss efet w=20300 l=13050
M1297 R14_0 N0647 N0532 vss efet w=7975 l=15225
M1298 N0968 R10_1 vss vss efet w=26100 l=13050
M1299 N0881 N0632 N0968 vss efet w=26100 l=12325
M1300 N0985 R14_0 vss vss efet w=26100 l=13050
M1301 N0880 N0657 N0985 vss efet w=26100 l=14500
M1302 R6_1 N0583 N0533 vss efet w=5800 l=11600
M1303 N0534 N0569 R5_1 vss efet w=5800 l=10875
M1304 R7_1 N0583 N0534 vss efet w=5800 l=11600
M1305 N0923 R3_1 vss vss efet w=24650 l=13050
M1306 vss R1_2 N0907 vss efet w=23925 l=13775
M1307 vss N0868 N0535 vss efet w=58725 l=12325
M1308 N0907 N0543 N0868 vss efet w=25375 l=12325
M1309 N0867 N0565 N0923 vss efet w=29000 l=10875
M1310 N0932 N0581 N0867 vss efet w=26100 l=11600
M1311 vss R5_1 N0932 vss efet w=23200 l=13050
M1312 N0533 N0598 R8_1 vss efet w=5800 l=13050
M1313 N0977 N0645 N0881 vss efet w=24650 l=11600
M1314 vss R12_1 N0977 vss efet w=21025 l=13775
M1315 vcc SC_A22_M22_CLK2 N0866 vss efet w=11600 l=14500
M1316 vcc vcc N0531 vss efet w=8700 l=33350
M1317 vcc vcc N0532 vss efet w=8700 l=33350
M1318 vcc SC_A22_M22_CLK2 N0880 vss efet w=13050 l=11600
M1319 N0986 R14_1 vss vss efet w=26100 l=13050
M1320 R10_1 N0619 N0533 vss efet w=5800 l=11600
M1321 N0534 N0598 R9_1 vss efet w=5800 l=14500
M1322 N0536 N0882 vss vss efet w=62350 l=11600
M1323 N0882 WRAB0 N0864 vss efet w=13050 l=11600
M1324 N0924 R3_2 vss vss efet w=23200 l=13050
M1325 N0868 N0565 N0924 vss efet w=27550 l=11600
M1326 N0933 N0581 N0868 vss efet w=24650 l=11600
M1327 vss R5_2 N0933 vss efet w=23200 l=13050
M1328 N0950 R7_1 vss vss efet w=23925 l=13775
M1329 N0867 N0591 N0950 vss efet w=27550 l=11600
M1330 N0959 N0616 N0867 vss efet w=26100 l=11600
M1331 vss R9_1 N0959 vss efet w=23200 l=14500
M1332 R11_1 N0619 N0534 vss efet w=7250 l=13050
M1333 N0533 N0634 R12_1 vss efet w=5800 l=13050
M1334 N0881 N0657 N0986 vss efet w=26100 l=14500
M1335 R14_1 N0647 N0533 vss efet w=6525 l=13775
M1336 N0534 N0634 R13_1 vss efet w=7250 l=13050
M1337 N0969 R11_1 vss vss efet w=23200 l=13775
M1338 N0867 N0632 N0969 vss efet w=25375 l=13775
M1339 N0978 N0645 N0867 vss efet w=24650 l=12325
M1340 vss R13_1 N0978 vss efet w=20300 l=11600
M1341 N0951 R7_2 vss vss efet w=23200 l=14500
M1342 N0535 N0529 R1_2 vss efet w=5800 l=12325
M1343 R3_2 N0544 N0535 vss efet w=6525 l=12325
M1344 N0536 N0529 R0_2 vss efet w=7975 l=10875
M1345 R2_2 N0544 N0536 vss efet w=5800 l=11600
M1346 N0908 N0543 N0882 vss efet w=24650 l=11600
M1347 vss R0_2 N0908 vss efet w=23200 l=13050
M1348 N0868 N0591 N0951 vss efet w=24650 l=11600
M1349 N0960 N0616 N0868 vss efet w=24650 l=11600
M1350 vss R9_2 N0960 vss efet w=23925 l=16675
M1351 R15_1 N0647 N0534 vss efet w=7975 l=15225
M1352 N0987 R15_1 vss vss efet w=27550 l=14500
M1353 N0970 R11_2 vss vss efet w=23200 l=14500
M1354 N0535 N0569 R5_2 vss efet w=5800 l=13050
M1355 R7_2 N0583 N0535 vss efet w=7250 l=10875
M1356 N0536 N0569 R4_2 vss efet w=5800 l=11600
M1357 vss R0_3 N0909 vss efet w=23925 l=13775
M1358 vcc vcc N0392 vss efet w=7250 l=29000
M1359 vcc __INH__X11_X31_CLK1 N0776 vss efet w=10875 l=11600
M1360 N0500 M12_M22_CLK1__M11_M12_ D3 vss efet w=13050 l=11600
M1361 D3 RRAB1 N0538 vss efet w=46400 l=11600
M1362 N0537 RRAB0 D3 vss efet w=44950 l=11600
M1363 N0842 PC3_1 vss vss efet w=23925 l=15225
M1364 PC1_1 N0410 N0393 vss efet w=5800 l=11600
M1365 N0780 N0444 N0842 vss efet w=25375 l=11600
M1366 N0393 N0426 PC2_1 vss efet w=5800 l=10150
M1367 PC3_1 N0439 N0393 vss efet w=5800 l=10150
M1368 N0394 N0381 PC0_0 vss efet w=5800 l=11600
M1369 N0794 N0406 N0781 vss efet w=27550 l=10875
M1370 vss PC0_0 N0794 vss efet w=23925 l=12325
M1371 PC1_0 N0410 N0394 vss efet w=5800 l=11600
M1372 N0815 PC1_0 vss vss efet w=23925 l=13775
M1373 N0394 N0426 PC2_0 vss efet w=5800 l=10150
M1374 vss N0777 N0395 vss efet w=68150 l=11600
M1375 vss PC0_4 N0795 vss efet w=24650 l=14500
M1376 N0764 WADB1 N0777 vss efet w=14500 l=11600
M1377 D0 RADB1 N0395 vss efet w=43500 l=11600
M1378 N0396 RADB2 D0 vss efet w=48575 l=10875
M1379 vcc N0325 N0306 vss efet w=7250 l=11600
M1380 N0314 N0306 vss vss efet w=29000 l=11600
M1381 N0795 N0406 N0777 vss efet w=26100 l=11600
M1382 N0781 N0424 N0815 vss efet w=25375 l=10875
M1383 N0830 N0434 N0781 vss efet w=26100 l=11600
M1384 vss PC2_0 N0830 vss efet w=23925 l=13050
M1385 PC3_0 N0439 N0394 vss efet w=5800 l=10875
M1386 N0843 PC3_0 vss vss efet w=22475 l=15225
M1387 N0816 PC1_4 vss vss efet w=21750 l=14500
M1388 N0777 N0424 N0816 vss efet w=25375 l=10875
M1389 vss N0773 N0396 vss efet w=68875 l=13775
M1390 N0773 WADB2 N0764 vss efet w=13050 l=11600
M1391 N0395 N0381 PC0_4 vss efet w=6525 l=13775
M1392 N0831 N0434 N0777 vss efet w=24650 l=11600
M1393 vss PC2_4 N0831 vss efet w=23200 l=14500
M1394 N0781 N0444 N0843 vss efet w=24650 l=11600
M1395 vcc __INH__X11_X31_CLK1 N0780 vss efet w=8700 l=13050
M1396 N0883 WRAB0 N0865 vss efet w=13050 l=11600
M1397 N0865 WRAB1 N0869 vss efet w=15225 l=10150
M1398 vss N0883 N0537 vss efet w=59450 l=11600
M1399 N0909 N0543 N0883 vss efet w=24650 l=11600
M1400 N0925 R2_2 vss vss efet w=23925 l=13775
M1401 N0882 N0565 N0925 vss efet w=24650 l=11600
M1402 N0934 N0581 N0882 vss efet w=24650 l=13050
M1403 vss R4_2 N0934 vss efet w=25375 l=12325
M1404 N0926 R2_3 vss vss efet w=23200 l=13050
M1405 R6_2 N0583 N0536 vss efet w=5800 l=11600
M1406 N0868 N0632 N0970 vss efet w=25375 l=12325
M1407 N0979 N0645 N0868 vss efet w=27550 l=11600
M1408 vss R13_2 N0979 vss efet w=20300 l=11600
M1409 N0535 N0598 R9_2 vss efet w=5800 l=11600
M1410 R11_2 N0619 N0535 vss efet w=6525 l=13050
M1411 N0867 N0657 N0987 vss efet w=25375 l=12325
M1412 vcc SC_A22_M22_CLK2 N0881 vss efet w=11600 l=14500
M1413 vcc vcc N0533 vss efet w=7250 l=37700
M1414 vcc vcc N0534 vss efet w=7975 l=35525
M1415 vcc SC_A22_M22_CLK2 N0867 vss efet w=12325 l=13775
M1416 N0988 R15_2 vss vss efet w=27550 l=14500
M1417 N0868 N0657 N0988 vss efet w=26100 l=12325
M1418 N0536 N0598 R8_2 vss efet w=5800 l=11600
M1419 N0538 N0869 vss vss efet w=59450 l=11600
M1420 N0883 N0565 N0926 vss efet w=24650 l=11600
M1421 N0935 N0581 N0883 vss efet w=24650 l=11600
M1422 vss R4_3 N0935 vss efet w=26825 l=13050
M1423 N0952 R6_2 vss vss efet w=23925 l=15225
M1424 N0882 N0591 N0952 vss efet w=28275 l=10875
M1425 N0961 N0616 N0882 vss efet w=29725 l=10875
M1426 vss R8_2 N0961 vss efet w=25375 l=13775
M1427 R10_2 N0619 N0536 vss efet w=5800 l=11600
M1428 N0535 N0634 R13_2 vss efet w=5800 l=12325
M1429 R15_2 N0647 N0535 vss efet w=6525 l=13775
M1430 N0536 N0634 R12_2 vss efet w=6525 l=13775
M1431 R14_2 N0647 N0536 vss efet w=6525 l=15225
M1432 N0971 R10_2 vss vss efet w=24650 l=13050
M1433 N0882 N0632 N0971 vss efet w=26825 l=12325
M1434 N0980 N0645 N0882 vss efet w=29000 l=11600
M1435 N0953 R6_3 vss vss efet w=23200 l=13775
M1436 N0537 N0529 R0_3 vss efet w=6525 l=13775
M1437 R2_3 N0544 N0537 vss efet w=4350 l=12325
M1438 N0538 N0529 R1_3 vss efet w=7250 l=11600
M1439 R3_3 N0544 N0538 vss efet w=5800 l=11600
M1440 N0910 N0543 N0869 vss efet w=24650 l=13775
M1441 vss R1_3 N0910 vss efet w=23200 l=13050
M1442 N0537 N0569 R4_3 vss efet w=7250 l=11600
M1443 N0883 N0591 N0953 vss efet w=26825 l=11600
M1444 N0962 N0616 N0883 vss efet w=26825 l=12325
M1445 vss R8_3 N0962 vss efet w=26100 l=15950
M1446 vss R12_2 N0980 vss efet w=21025 l=15225
M1447 N0972 R10_3 vss vss efet w=24650 l=14500
M1448 R6_3 N0583 N0537 vss efet w=6525 l=13775
M1449 N0538 N0569 R5_3 vss efet w=5800 l=11600
M1450 vcc vcc N0393 vss efet w=5800 l=30450
M1451 vss N0461 N0469 vss efet w=13050 l=13050
M1452 N0469 vcc vcc vss efet w=8700 l=65250
M1453 N0461 N0469 vss vss efet w=11600 l=11600
M1454 N0927 R3_3 vss vss efet w=23925 l=13775
M1455 N0869 N0565 N0927 vss efet w=27550 l=11600
M1456 N0936 N0581 N0869 vss efet w=27550 l=13050
M1457 vss R5_3 N0936 vss efet w=27550 l=13050
M1458 R7_3 N0583 N0538 vss efet w=5800 l=11600
M1459 N0883 N0632 N0972 vss efet w=26100 l=13050
M1460 N0981 N0645 N0883 vss efet w=31175 l=13775
M1461 vss R12_3 N0981 vss efet w=22475 l=17400
M1462 N0989 R14_2 vss vss efet w=29725 l=15225
M1463 N0882 N0657 N0989 vss efet w=27550 l=13050
M1464 vcc SC_A22_M22_CLK2 N0868 vss efet w=14500 l=14500
M1465 vcc vcc N0535 vss efet w=8700 l=34075
M1466 vcc vcc N0536 vss efet w=7975 l=32625
M1467 vcc SC_A22_M22_CLK2 N0882 vss efet w=11600 l=13050
M1468 N0990 R14_3 vss vss efet w=29000 l=13050
M1469 N0883 N0657 N0990 vss efet w=29000 l=11600
M1470 N0537 N0598 R8_3 vss efet w=5800 l=11600
M1471 R10_3 N0619 N0537 vss efet w=5800 l=13775
M1472 N0538 N0598 R9_3 vss efet w=5800 l=11600
M1473 N0954 R7_3 vss vss efet w=23925 l=13775
M1474 N0869 N0591 N0954 vss efet w=27550 l=11600
M1475 N0963 N0616 N0869 vss efet w=27550 l=11600
M1476 vss R9_3 N0963 vss efet w=25375 l=13775
M1477 R11_3 N0619 N0538 vss efet w=5800 l=11600
M1478 N0973 R11_3 vss vss efet w=26825 l=14500
M1479 N0537 N0634 R12_3 vss efet w=5800 l=11600
M1480 vcc SC_A22_M22_CLK2 N0883 vss efet w=11600 l=13050
M1481 R14_3 N0647 N0537 vss efet w=5800 l=13050
M1482 N0538 N0634 R13_3 vss efet w=5800 l=13050
M1483 R15_3 N0647 N0538 vss efet w=7250 l=14500
M1484 N0869 N0632 N0973 vss efet w=26100 l=12325
M1485 N0982 N0645 N0869 vss efet w=26100 l=13050
M1486 vss R13_3 N0982 vss efet w=27550 l=15950
M1487 vcc vcc N0537 vss efet w=8700 l=34075
M1488 vss vss clk2 vss efet w=118175 l=13775
M1489 vss vss clk1 vss efet w=113100 l=13050
M1490 vcc vcc N0538 vss efet w=8700 l=34075
M1491 N0991 R15_3 vss vss efet w=26100 l=15950
M1492 N0869 N0657 N0991 vss efet w=26825 l=12325
M1493 vcc SC_A22_M22_CLK2 N0869 vss efet w=11600 l=14500
M1494 vcc vcc N0394 vss efet w=5800 l=29000
M1495 vcc vcc N0461 vss efet w=5800 l=65250
M1496 ADDR_RFSH_1 vcc vcc vss efet w=8700 l=66700
M1497 vss N0461 ADDR_RFSH_1 vss efet w=15225 l=10875
M1498 N0453 N0469 vss vss efet w=14500 l=11600
M1499 vss N0902 N0543 vss efet w=14500 l=11600
M1500 vss N0902 N0529 vss efet w=11600 l=11600
M1501 vss N0919 N0544 vss efet w=11600 l=11600
M1502 vss N0919 N0565 vss efet w=14500 l=11600
M1503 vcc vcc N0453 vss efet w=9425 l=65975
M1504 vcc __INH__X11_X31_CLK1 N0781 vss efet w=9425 l=10875
M1505 N0902 vcc vcc vss efet w=6525 l=61625
M1506 N0543 N0530 __POC__CLK2_SC_A32_X12_ vss efet w=16675 l=10875
M1507 N0529 N0530 CLK2_SC_A12_M12_ vss efet w=13775 l=13050
M1508 N0544 N0545 CLK2_SC_A12_M12_ vss efet w=12325 l=10875
M1509 N0565 N0545 __POC__CLK2_SC_A32_X12_ vss efet w=16675 l=12325
M1510 N0844 PC3_4 vss vss efet w=22475 l=18125
M1511 ADDR_RFSH_1 N0455 N0489 vss efet w=8700 l=10150
M1512 N0453 N0455 N0454 vss efet w=8700 l=13050
M1513 PC1_4 N0410 N0395 vss efet w=6525 l=12325
M1514 N0396 N0381 PC0_8 vss efet w=5800 l=11600
M1515 N0796 N0406 N0773 vss efet w=27550 l=13050
M1516 vcc vcc N0314 vss efet w=7250 l=65250
M1517 vss A32 N0712 vss efet w=24650 l=11600
M1518 N0314 clk2 N0315 vss efet w=13050 l=14500
M1519 cm_rom N0717 vcc vss efet w=417600 l=11600
M1520 vss N0737 cm_rom vss efet w=607550 l=10875
M1521 N0712 A22 vss vss efet w=26825 l=12325
M1522 N0325 vcc clk1 vss efet w=34800 l=11600
M1523 vcc vcc WADB1 vss efet w=5800 l=27550
M1524 vss A12 N0711 vss efet w=13050 l=12325
M1525 N0316 N0315 vss vss efet w=20300 l=11600
M1526 WADB0 vcc vcc vss efet w=7250 l=27550
M1527 vss N0300 WADB0 vss efet w=29000 l=13050
M1528 vcc vcc N0316 vss efet w=6525 l=51475
M1529 N0711 vcc vcc vss efet w=6525 l=67425
M1530 N0317 clk1 N0316 vss efet w=8700 l=11600
M1531 vss N0326 WADB0 vss efet w=36250 l=11600
M1532 vss PC0_8 N0796 vss efet w=23925 l=12325
M1533 PC1_8 N0410 N0396 vss efet w=5800 l=11600
M1534 N0777 N0444 N0844 vss efet w=24650 l=11600
M1535 N0395 N0426 PC2_4 vss efet w=6525 l=10875
M1536 PC3_4 N0439 N0395 vss efet w=5800 l=10150
M1537 N0396 N0426 PC2_8 vss efet w=5800 l=10150
M1538 PC3_8 N0439 N0396 vss efet w=5800 l=10150
M1539 N0817 PC1_8 vss vss efet w=26100 l=13050
M1540 N0773 N0424 N0817 vss efet w=27550 l=13050
M1541 N0832 N0434 N0773 vss efet w=25375 l=12325
M1542 WADB2 vcc vcc vss efet w=7975 l=31175
M1543 vss PC2_8 N0832 vss efet w=25375 l=13050
M1544 N0845 PC3_8 vss vss efet w=23925 l=15225
M1545 N0773 N0444 N0845 vss efet w=26825 l=13775
M1546 vcc __INH__X11_X31_CLK1 N0777 vss efet w=8700 l=11600
M1547 N0488 N0463 N0469 vss efet w=21750 l=12325
M1548 vcc vcc N0395 vss efet w=6525 l=32625
M1549 vss N0489 N0488 vss efet w=34075 l=11600
M1550 N0462 N0454 vss vss efet w=34800 l=11600
M1551 N0461 N0463 N0462 vss efet w=20300 l=11600
M1552 vcc vcc N0396 vss efet w=6525 l=31175
M1553 vss N0928 N0581 vss efet w=14500 l=10150
M1554 vss N0928 N0569 vss efet w=11600 l=10150
M1555 vss N0938 N0583 vss efet w=13050 l=10150
M1556 vss N0938 N0591 vss efet w=15950 l=10150
M1557 vss N0955 N0616 vss efet w=13775 l=10875
M1558 N0581 N0570 __POC__CLK2_SC_A32_X12_ vss efet w=14500 l=11600
M1559 N0569 N0570 CLK2_SC_A12_M12_ vss efet w=12325 l=12325
M1560 N0583 N0584 CLK2_SC_A12_M12_ vss efet w=13050 l=11600
M1561 N0591 N0584 __POC__CLK2_SC_A32_X12_ vss efet w=14500 l=13050
M1562 vss N0530 N0902 vss efet w=11600 l=13050
M1563 N0919 N0545 vss vss efet w=10150 l=11600
M1564 vss N0570 N0928 vss efet w=10875 l=12325
M1565 N0938 N0584 vss vss efet w=10150 l=13050
M1566 vss N0955 N0598 vss efet w=13050 l=10875
M1567 vss N0965 N0619 vss efet w=11600 l=11600
M1568 vss N0965 N0632 vss efet w=13050 l=12325
M1569 N0616 N0599 __POC__CLK2_SC_A32_X12_ vss efet w=14500 l=10875
M1570 CLK2_SC_A12_M12_ N0599 N0598 vss efet w=12325 l=10875
M1571 N0619 N0620 CLK2_SC_A12_M12_ vss efet w=12325 l=10875
M1572 N0632 N0620 __POC__CLK2_SC_A32_X12_ vss efet w=13050 l=10150
M1573 vss N0599 N0955 vss efet w=12325 l=12325
M1575 RRAB1 S00557 vcc vss efet w=10150 l=23200
M1576 S00557 vcc vcc vss efet w=6525 l=13775
M1577 vcc __INH__X11_X31_CLK1 N0773 vss efet w=10150 l=11600
M1578 N0463 vcc vcc vss efet w=6525 l=71775
M1579 vss N0455 N0463 vss efet w=11600 l=11600
M1580 N0455 N0463 vss vss efet w=13050 l=11600
M1581 N0919 vcc vcc vss efet w=6525 l=45675
M1582 vcc vcc N0928 vss efet w=7975 l=51475
M1583 N0965 N0620 vss vss efet w=11600 l=13050
M1584 vss N0974 N0645 vss efet w=14500 l=11600
M1585 vss N0974 N0634 vss efet w=11600 l=11600
M1586 vss N0983 N0647 vss efet w=11600 l=11600
M1587 vss N0983 N0657 vss efet w=14500 l=11600
M1588 N0645 N0635 __POC__CLK2_SC_A32_X12_ vss efet w=15225 l=10875
M1589 N0634 N0635 CLK2_SC_A12_M12_ vss efet w=12325 l=10875
M1590 N0647 N0648 CLK2_SC_A12_M12_ vss efet w=12325 l=10875
M1591 N0657 N0648 __POC__CLK2_SC_A32_X12_ vss efet w=14500 l=11600
M1592 N0938 vcc vcc vss efet w=5800 l=47850
M1593 vcc vcc N0955 vss efet w=6525 l=52925
M1594 vss N0635 N0974 vss efet w=10150 l=13050
M1595 N0983 N0648 vss vss efet w=10150 l=13050
M1596 vcc vcc N0613 vss efet w=13050 l=45675
M1597 N0965 vcc vcc vss efet w=6525 l=48575
M1598 vcc vcc N0974 vss efet w=5800 l=47850
M1599 N0983 vcc vcc vss efet w=5800 l=47850
M1600 N0539 N0540 vss vss efet w=27550 l=13050
M1601 vcc vcc N0540 vss efet w=7250 l=29000
M1602 vcc vcc N0455 vss efet w=6525 l=68875
M1603 ADDR_RFSH_0 vcc vcc vss efet w=9425 l=73950
M1604 vss N0455 ADDR_RFSH_0 vss efet w=13775 l=10875
M1605 N0503 N0463 vss vss efet w=13050 l=11600
M1606 vcc vcc N0503 vss efet w=8700 l=66700
M1607 S00564 vcc vcc vss efet w=6525 l=13775
M1609 RRAB0 S00564 vcc vss efet w=7250 l=21750
M1610 WADB1 N0318 vss vss efet w=27550 l=11600
M1611 vss N0304 WADB2 vss efet w=29000 l=13050
M1612 vss N0300 WADB1 vss efet w=27550 l=12325
M1613 WADB2 N0300 vss vss efet w=29725 l=10875
M1614 vss N0783 N0406 vss efet w=15950 l=10150
M1615 vss N0783 N0381 vss efet w=11600 l=10150
M1616 vss N0804 N0410 vss efet w=11600 l=11600
M1617 vss N0804 N0424 vss efet w=15950 l=10150
M1618 N0406 N0382 __POC_CLK2_X12_X32__INH vss efet w=15950 l=11600
M1619 N0381 N0382 ___SC__JIN_FIN__CLK1_M11_X21_INH_ vss efet w=10150 l=11600
M1620 N0410 N0411 ___SC__JIN_FIN__CLK1_M11_X21_INH_ vss efet w=12325 l=12325
M1621 N0424 N0411 __POC_CLK2_X12_X32__INH vss efet w=15950 l=11600
M1622 N0737 vcc vcc vss efet w=9425 l=13775
M1623 N0711 N0732 N0712 vss efet w=23200 l=10150
M1624 vss N0820 N0434 vss efet w=15950 l=10150
M1625 N0426 N0820 vss vss efet w=11600 l=11600
M1626 vss N0833 N0439 vss efet w=11600 l=11600
M1627 N0444 N0833 vss vss efet w=15950 l=13050
M1628 ADDR_RFSH_0 clk1 N0519 vss efet w=7250 l=11600
M1629 N0545 N0540 vss vss efet w=14500 l=10150
M1630 N0570 N0540 vss vss efet w=14500 l=11600
M1631 N0584 N0540 vss vss efet w=13775 l=14500
M1632 N0599 N0613 vss vss efet w=13775 l=13775
M1633 vss N0613 N0540 vss efet w=32625 l=10875
M1634 N0620 N0613 vss vss efet w=15225 l=12325
M1635 N0635 N0613 vss vss efet w=13775 l=13775
M1636 N0648 N0613 vss vss efet w=16675 l=13050
M1637 N0613 N0646 vss vss efet w=52925 l=15225
M1638 N0539 N0541 vss vss efet w=27550 l=10150
M1639 N0545 N0541 vss vss efet w=14500 l=10875
M1640 vss N0541 N0599 vss efet w=13775 l=12325
M1641 vss N0541 N0620 vss efet w=13775 l=10875
M1642 N0570 N0577 vss vss efet w=13775 l=13775
M1643 vss N0542 N0539 vss efet w=29000 l=11600
M1644 N0584 N0577 vss vss efet w=13775 l=13775
M1645 N0503 clk1 N0504 vss efet w=7250 l=13050
M1646 N0635 N0577 vss vss efet w=13050 l=10150
M1647 N0648 N0577 vss vss efet w=15950 l=15950
M1648 vcc vcc N0541 vss efet w=9425 l=38425
M1649 N0570 N0542 vss vss efet w=14500 l=15950
M1650 N0434 N0427 __POC_CLK2_X12_X32__INH vss efet w=15950 l=11600
M1651 N0426 N0427 ___SC__JIN_FIN__CLK1_M11_X21_INH_ vss efet w=10875 l=13775
M1652 N0439 N0440 ___SC__JIN_FIN__CLK1_M11_X21_INH_ vss efet w=11600 l=11600
M1653 N0444 N0440 __POC_CLK2_X12_X32__INH vss efet w=18125 l=12325
M1654 vss N0519 N0518 vss efet w=40600 l=11600
M1655 vss N0382 N0783 vss efet w=12325 l=12325
M1656 N0804 N0411 vss vss efet w=11600 l=11600
M1657 N0518 __INH__X32_CLK2 N0463 vss efet w=21750 l=13050
M1658 N0508 N0504 vss vss efet w=38425 l=12325
M1659 vss N0542 N0599 vss efet w=14500 l=13050
M1660 vss N0542 N0635 vss efet w=13050 l=10150
M1661 N0541 N0577 vss vss efet w=26100 l=11600
M1662 N0577 N0617 vss vss efet w=52200 l=13050
M1663 N0455 __INH__X32_CLK2 N0508 vss efet w=19575 l=13050
M1664 N0539 __FIN_X12_ N0530 vss efet w=41325 l=12325
M1665 N0561 vcc vcc vss efet w=8700 l=40600
M1666 vss __FIN_X12_ N0561 vss efet w=29000 l=11600
M1667 vcc vcc N0833 vss efet w=5800 l=60900
M1668 vss N0427 N0820 vss efet w=11600 l=10875
M1669 N0833 N0440 vss vss efet w=11600 l=11600
M1670 N0732 N0317 vss vss efet w=19575 l=12325
M1671 vcc vcc N0732 vss efet w=8700 l=65250
M1672 vss N0711 N0307 vss efet w=13775 l=11600
M1673 vss N0416 RADB0 vss efet w=43500 l=13050
M1674 RADB2 vcc vcc vss efet w=7975 l=23200
M1675 N0300 clk2 vss vss efet w=26100 l=13050
M1676 N0307 vcc vcc vss efet w=10150 l=50750
M1677 vss clk1 N0307 vss efet w=15950 l=10150
M1678 vcc vcc N0300 vss efet w=6525 l=29725
M1679 vss N0717 N0737 vss efet w=94250 l=13050
M1680 M12_M22_CLK1__M11_M12_ N0710 vcc vss efet w=23925 l=15225
M1681 vss N0708 M12_M22_CLK1__M11_M12_ vss efet w=20300 l=13775
M1683 S00609 vcc vcc vss efet w=7250 l=11600
M1684 vss N0708 N0710 vss efet w=14500 l=11600
M1685 N0402 vcc vcc vss efet w=7975 l=60900
M1686 vss X32 N0402 vss efet w=15950 l=10150
M1687 RADB1 vcc vcc vss efet w=7975 l=26825
M1688 RADB0 vcc vcc vss efet w=8700 l=21750
M1689 RADB1 clk2 vss vss efet w=50750 l=11600
M1690 vss N0384 RADB1 vss efet w=42775 l=13775
M1691 RADB2 clk2 vss vss efet w=53650 l=13050
M1692 vss N0374 RADB2 vss efet w=50025 l=11600
M1693 vcc vcc N0783 vss efet w=5800 l=62350
M1694 vcc vcc N0804 vss efet w=6525 l=50025
M1695 N0820 vcc vcc vss efet w=5800 l=52200
M1696 N0400 N0409 vss vss efet w=23925 l=10875
M1697 vss N0560 N0545 vss efet w=15225 l=10875
M1698 N0584 N0560 vss vss efet w=14500 l=11600
M1699 N0620 N0560 vss vss efet w=14500 l=10150
M1700 N0648 N0560 vss vss efet w=14500 l=12325
M1701 N0545 N0561 vss vss efet w=14500 l=13775
M1702 N0570 N0561 vss vss efet w=15225 l=13775
M1703 N0584 N0561 vss vss efet w=15225 l=12325
M1704 N0599 N0561 vss vss efet w=16675 l=11600
M1705 N0620 N0561 vss vss efet w=15225 l=10875
M1706 N0635 N0561 vss vss efet w=14500 l=11600
M1707 N0648 N0561 vss vss efet w=14500 l=13050
M1709 vcc vcc N0400 vss efet w=8700 l=65250
M1711 N0427 N0400 vss vss efet w=11600 l=13050
M1712 N0475 vcc vcc vss efet w=7250 l=65250
M1713 vss N0464 N0475 vss efet w=14500 l=13050
M1714 ADDR_PTR_1 vcc vcc vss efet w=8700 l=68150
M1715 vss N0464 ADDR_PTR_1 vss efet w=15225 l=13050
M1716 N0464 N0475 vss vss efet w=13050 l=11600
M1717 vcc vcc N0464 vss efet w=6525 l=67425
M1718 N0457 N0475 vss vss efet w=14500 l=13050
M1719 vcc vcc N0457 vss efet w=8700 l=66700
M1720 N0440 N0409 vss vss efet w=19575 l=12325
M1721 ADDR_PTR_1 N0459 N0492 vss efet w=8700 l=11600
M1722 N0457 N0459 N0458 vss efet w=9425 l=12325
M1723 N0402 clk2 N0416 vss efet w=7250 l=13050
M1724 N0384 clk2 N0379 vss efet w=7250 l=11600
M1725 N0374 clk2 N0365 vss efet w=7975 l=13775
M1726 N0710 S00609 vcc vss efet w=7975 l=37700
M1727 N0379 A12 vss vss efet w=14500 l=11600
M1728 vss A22 N0365 vss efet w=15950 l=10150
M1729 vcc vcc N0365 vss efet w=9425 l=55825
M1730 vcc vcc N0708 vss efet w=8700 l=34800
M1731 N0708 clk1 N0709 vss efet w=48575 l=15225
M1732 N0709 N0278 vss vss efet w=44225 l=12325
M1733 vcc vcc N0279 vss efet w=6525 l=41325
M1734 vss M12 N0708 vss efet w=22475 l=13050
M1735 N0708 M22 vss vss efet w=23200 l=8700
M1736 vcc vcc N0379 vss efet w=6525 l=52925
M1737 N0278 clk2 N0279 vss efet w=14500 l=11600
M1738 vss M12 N0279 vss efet w=21025 l=12325
M1739 RADB0 clk2 vss vss efet w=43500 l=11600
M1740 N0382 N0400 vss vss efet w=13050 l=10150
M1741 N0411 N0409 vss vss efet w=20300 l=10150
M1742 N0382 N0401 vss vss efet w=12325 l=10150
M1743 N0411 N0401 vss vss efet w=13050 l=11600
M1744 vss N0420 N0427 vss efet w=20300 l=10150
M1745 N0440 N0420 vss vss efet w=20300 l=13050
M1747 vss A32 N0279 vss efet w=23200 l=11600
M1748 vcc vcc N0304 vss efet w=7250 l=69600
M1749 N0382 S00598 vcc vss efet w=7250 l=56550
M1752 vss N0492 N0491 vss efet w=39150 l=11600
M1754 N0411 S00599 vcc vss efet w=7250 l=55100
M1755 N0427 S00600 vcc vss efet w=7250 l=56550
M1756 N0401 N0420 vss vss efet w=24650 l=11600
M1757 vcc vcc N0401 vss efet w=8700 l=66700
M1758 N0491 N0466 N0475 vss efet w=21750 l=14500
M1759 N0465 N0458 vss vss efet w=39150 l=13050
M1760 N0464 N0466 N0465 vss efet w=19575 l=13775
M1761 N0530 S00578 vcc vss efet w=10150 l=55825
M1763 N0545 S00579 vcc vss efet w=7975 l=60175
M1764 N0570 S00580 vcc vss efet w=7250 l=56550
M1769 N0584 S00581 vcc vss efet w=7250 l=56550
M1770 N0599 S00582 vcc vss efet w=8700 l=59450
M1771 N0620 S00583 vcc vss efet w=9425 l=54375
M1772 N0635 S00584 vcc vss efet w=9425 l=55825
M1773 vcc vcc N0577 vss efet w=8700 l=37700
M1774 vcc vcc N0542 vss efet w=11600 l=42775
M1776 N0542 N0560 vss vss efet w=26100 l=10150
M1777 N0560 N0582 vss vss efet w=48575 l=10875
M1778 vcc vcc N0560 vss efet w=10150 l=44225
M1779 N0648 S00585 vcc vss efet w=7250 l=53650
M1780 D1 SC_M22_CLK2 N0582 vss efet w=8700 l=13050
M1781 D2 SC_M22_CLK2 N0617 vss efet w=7250 l=13050
M1782 S00578 vcc vcc vss efet w=8700 l=11600
M1783 S00579 vcc vcc vss efet w=8700 l=12325
M1784 S00580 vcc vcc vss efet w=10150 l=10150
M1785 S00581 vcc vcc vss efet w=10150 l=10150
M1786 S00582 vcc vcc vss efet w=8700 l=10150
M1787 S00583 vcc vcc vss efet w=9425 l=10875
M1788 S00584 vcc vcc vss efet w=10875 l=14500
M1789 S00585 vcc vcc vss efet w=10150 l=11600
M1790 vcc vcc N0571 vss efet w=5800 l=68875
M1791 vcc vcc N0574 vss efet w=6525 l=65975
M1792 vcc vcc N0573 vss efet w=5800 l=66700
M1793 vcc vcc N0600 vss efet w=5800 l=63800
M1794 N0582 SC_A22 REG_RFSH_0 vss efet w=8700 l=11600
M1795 vcc vcc REG_RFSH_0 vss efet w=5800 l=33350
M1796 vcc vcc N0610 vss efet w=5800 l=72500
M1797 vcc vcc N0609 vss efet w=5800 l=63800
M1798 vcc vcc REG_RFSH_1 vss efet w=6525 l=41325
M1799 N0617 SC_A22 REG_RFSH_1 vss efet w=10875 l=10875
M1800 N0440 S00601 vcc vss efet w=7250 l=53650
M1801 N0409 X12 ADDR_RFSH_1 vss efet w=8700 l=11600
M1802 ADDR_PTR_1 X32 N0409 vss efet w=8700 l=11600
M1803 N0420 X12 ADDR_RFSH_0 vss efet w=8700 l=11600
M1804 ADDR_PTR_0 X32 N0420 vss efet w=7975 l=13050
M1806 vcc vcc N0450 vss efet w=7250 l=59450
M1807 S00598 vcc vcc vss efet w=10150 l=11600
M1808 S00599 vcc vcc vss efet w=11600 l=10150
M1809 S00600 vcc vcc vss efet w=10875 l=10150
M1810 S00601 vcc vcc vss efet w=11600 l=11600
M1811 __POC_CLK2_X12_X32__INH N0449 vcc vss efet w=41325 l=21025
M1812 vcc vcc S00613 vss efet w=7975 l=12325
M1813 vss JUN_JMS N0309 vss efet w=34075 l=13775
M1814 vcc S00613 N0449 vss efet w=5800 l=43500
M1815 vss N0450 __POC_CLK2_X12_X32__INH vss efet w=29725 l=12325
M1816 vcc vcc N0318 vss efet w=6525 l=68875
M1817 N0308 X22 N0304 vss efet w=30450 l=11600
M1818 N0309 N0310 N0308 vss efet w=30450 l=11600
M1819 N0323 M12 vss vss efet w=32625 l=12325
M1820 N0304 A32 vss vss efet w=13050 l=11600
M1821 N0323 JUN_JMS N0324 vss efet w=36975 l=20300
M1822 N0320 SC vss vss efet w=30450 l=13050
M1823 N0319 JIN_FIN N0320 vss efet w=29000 l=13050
M1824 N0318 X22 N0319 vss efet w=30450 l=11600
M1825 N0324 N0310 N0318 vss efet w=29000 l=11600
M1826 N0321 JCN_ISZ N0323 vss efet w=30450 l=11600
M1827 N0318 N0322 N0321 vss efet w=31175 l=12325
M1828 N0450 N0449 vss vss efet w=13050 l=14500
M1829 vcc vcc N0437 vss efet w=8700 l=51475
M1830 vss N0437 ___SC__JIN_FIN__CLK1_M11_X21_INH_ vss efet w=20300 l=10150
M1831 vcc S00612 N0436 vss efet w=7250 l=40600
M1832 vcc vcc S00612 vss efet w=5800 l=10150
M1833 S00628 vcc vcc vss efet w=5800 l=11600
M1834 vcc S00628 __INH__X11_X31_CLK1 vss efet w=7975 l=18125
M1836 vcc N0436 ___SC__JIN_FIN__CLK1_M11_X21_INH_ vss efet w=21025 l=12325
M1837 vss N0436 N0437 vss efet w=13775 l=13775
M1839 __INH__X11_X31_CLK1 N0517 vss vss efet w=35525 l=12325
M1840 vss INH __INH__X11_X31_CLK1 vss efet w=36250 l=11600
M1841 vss N0522 __INH__X11_X31_CLK1 vss efet w=34800 l=11600
M1842 vcc vcc N0451 vss efet w=5800 l=50750
M1843 N0449 INH vss vss efet w=13775 l=10875
M1844 N0436 N0443 vss vss efet w=13775 l=10875
M1845 N0436 N0435 N0441 vss efet w=29725 l=10875
M1846 N0449 POC vss vss efet w=15225 l=12325
M1847 vss N0447 N0449 vss efet w=14500 l=12325
M1848 N0449 N0451 vss vss efet w=14500 l=11600
M1849 N0441 JIN_FIN vss vss efet w=29725 l=10875
M1850 vss N0438 N0436 vss efet w=15225 l=10875
M1851 vss A22 N0318 vss efet w=18125 l=13775
M1852 N0451 clk2 vss vss efet w=14500 l=10150
M1853 vss _CN N0322 vss efet w=34075 l=13775
M1854 N0322 SC vss vss efet w=26825 l=13775
M1855 N0333 SC N0326 vss efet w=32625 l=10150
M1856 N0326 A12 vss vss efet w=12325 l=10875
M1857 N0334 JIN_FIN N0333 vss efet w=31900 l=10150
M1858 vss X32 N0334 vss efet w=30450 l=10150
M1859 vcc vcc N0326 vss efet w=7975 l=64525
M1860 N0341 N0310 N0339 vss efet w=36250 l=11600
M1861 N0326 JUN_JMS N0341 vss efet w=38425 l=10875
M1862 N0338 JCN_ISZ N0326 vss efet w=33350 l=11600
M1863 N0339 N0322 N0338 vss efet w=33350 l=11600
M1864 vss M22 N0339 vss efet w=34800 l=10150
M1865 vss SC N0310 vss efet w=27550 l=10875
M1866 N0310 vcc vcc vss efet w=5800 l=27550
M1867 N0322 vcc vcc vss efet w=6525 l=28275
M1868 N0344 S00654 vcc vss efet w=6525 l=28275
M1869 vcc N0344 SC vss efet w=37700 l=11600
M1870 vcc vcc S00654 vss efet w=6525 l=13050
M1871 vss X12 N0447 vss efet w=15225 l=12325
M1872 vss X32 N0447 vss efet w=12325 l=12325
M1873 vcc vcc N0443 vss efet w=6525 l=51475
M1874 N0447 vcc vcc vss efet w=5800 l=66700
M1875 N0443 clk1 vss vss efet w=14500 l=10150
M1876 vcc vcc _INH vss efet w=5800 l=27550
M1877 vcc vcc INH vss efet w=5800 l=29000
M1878 N0511 vcc vcc vss efet w=7975 l=54375
M1879 N0517 clk2 N0511 vss efet w=9425 l=15225
M1880 N0466 vcc vcc vss efet w=6525 l=73225
M1881 vss N0459 N0466 vss efet w=11600 l=11600
M1882 vss N0459 ADDR_PTR_0 vss efet w=18850 l=10150
M1883 ADDR_PTR_0 vcc vcc vss efet w=7975 l=68875
M1884 N0459 N0466 vss vss efet w=13050 l=11600
M1885 vcc vcc N0459 vss efet w=6525 l=65250
M1886 N0505 N0466 vss vss efet w=14500 l=11600
M1887 vcc vcc N0505 vss efet w=9425 l=76125
M1888 N0521 clk1 ADDR_PTR_0 vss efet w=8700 l=10875
M1889 N0505 clk1 N0506 vss efet w=7250 l=10150
M1890 REG_RFSH_0 clk1 N0566 vss efet w=7975 l=15225
M1891 N0571 SC_A12_CLK2 N0572 vss efet w=24650 l=12325
M1892 N0572 N0566 vss vss efet w=34075 l=12325
M1893 vss N0574 REG_RFSH_0 vss efet w=21750 l=11600
M1894 vss N0574 N0571 vss efet w=12325 l=12325
M1895 N0586 clk1 N0573 vss efet w=7975 l=13775
M1896 N0573 N0571 vss vss efet w=12325 l=12325
M1897 N0574 N0571 vss vss efet w=12325 l=12325
M1898 REG_RFSH_1 N0571 N0593 vss efet w=10150 l=12325
M1899 vss N0521 N0520 vss efet w=39150 l=13050
M1900 vcc vcc N0494 vss efet w=7250 l=65250
M1901 __INH__X32_CLK2 vcc vcc vss efet w=6525 l=28275
M1902 N0520 CLK2_JMS_DC_M22_BBL_M22_X12_X22__ N0466 vss efet w=19575 l=14500
M1903 N0509 N0506 vss vss efet w=39150 l=11600
M1904 N0459 CLK2_JMS_DC_M22_BBL_M22_X12_X22__ N0509 vss efet w=20300 l=13050
M1905 vss N0592 RRAB1 vss efet w=40600 l=12325
M1906 vss N0494 __INH__X32_CLK2 vss efet w=26100 l=11600
M1907 vcc vcc N0522 vss efet w=5800 l=36250
M1908 CLK2_JMS_DC_M22_BBL_M22_X12_X22__ N0467 vss vss efet w=26825 l=13050
M1909 vss DC RRAB1 vss efet w=31175 l=15225
M1910 N0574 SC_A12_CLK2 N0585 vss efet w=21025 l=12325
M1911 N0625 N0571 N0609 vss efet w=8700 l=13050
M1912 vss N0600 N0609 vss efet w=13050 l=12325
M1913 N0600 N0574 N0601 vss efet w=21750 l=13050
M1914 vss N0610 REG_RFSH_1 vss efet w=21750 l=10150
M1915 N0600 N0610 vss vss efet w=11600 l=10150
M1916 N0585 N0586 vss vss efet w=35525 l=13050
M1917 N0601 N0593 vss vss efet w=33350 l=11600
M1918 RRAB1 clk2 vss vss efet w=29000 l=13050
M1919 vcc vcc CLK2_JMS_DC_M22_BBL_M22_X12_X22__ vss efet w=9425 l=30450
M1920 vss clk2 N0496 vss efet w=29725 l=15225
M1921 N0496 X32 N0495 vss efet w=31175 l=12325
M1922 vss INH _INH vss efet w=26100 l=13775
M1923 vss N0524 INH vss efet w=26100 l=11600
M1924 vss M22 N0511 vss efet w=18850 l=11600
M1925 N0522 clk1 vss vss efet w=23200 l=11600
M1926 N0495 _INH N0494 vss efet w=29000 l=11600
M1927 N0429 X12 vss vss efet w=21750 l=13050
M1928 N0438 clk2 N0428 vss efet w=7975 l=12325
M1929 N0428 _INH N0429 vss efet w=21750 l=11600
M1930 N0435 SC vss vss efet w=14500 l=10875
M1931 vcc vcc N0528 vss efet w=5800 l=52200
M1932 N0428 vcc vcc vss efet w=5800 l=65250
M1933 N0428 A32 vss vss efet w=14500 l=10875
M1934 N0435 vcc vcc vss efet w=7250 l=47850
M1935 vss X22 N0511 vss efet w=15225 l=12325
M1936 vss DC N0526 vss efet w=29725 l=12325
M1937 vss _CN N0528 vss efet w=16675 l=11600
M1938 vss SC N0525 vss efet w=21750 l=11600
M1939 N0525 JIN_FIN N0524 vss efet w=25375 l=10875
M1940 N0526 N0528 N0527 vss efet w=29725 l=12325
M1941 vcc vcc N0467 vss efet w=5800 l=63800
M1942 N0485 JMS vss vss efet w=30450 l=11600
M1943 N0484 M22 N0485 vss efet w=31900 l=11600
M1944 N0467 DC N0484 vss efet w=30450 l=11600
M1945 vcc vcc N0460 vss efet w=5800 l=33350
M1946 vcc vcc N0588 vss efet w=5800 l=70325
M1947 N0592 clk2 N0588 vss efet w=13050 l=13050
M1948 vss clk2 N0460 vss efet w=21750 l=11600
M1949 N0610 N0600 vss vss efet w=12325 l=10875
M1950 N0610 N0574 N0624 vss efet w=21750 l=13050
M1951 N0624 N0625 vss vss efet w=36250 l=11600
M1952 D3 SC_M22_CLK2 N0646 vss efet w=10150 l=13050
M1953 vcc vcc N0637 vss efet w=5800 l=65250
M1954 vcc vcc N0642 vss efet w=6525 l=67425
M1955 vcc vcc N0641 vss efet w=7250 l=69600
M1956 N0646 SC_A22 REG_RFSH_2 vss efet w=7250 l=11600
M1957 vcc vcc REG_RFSH_2 vss efet w=5075 l=34075
M1958 REG_RFSH_2 N0600 N0633 vss efet w=7975 l=12325
M1959 N0637 N0610 N0638 vss efet w=21025 l=12325
M1960 vss N0642 REG_RFSH_2 vss efet w=21750 l=11600
M1961 N0637 N0642 vss vss efet w=13050 l=11600
M1962 N0638 N0633 vss vss efet w=36250 l=11600
M1963 N0653 N0600 N0641 vss efet w=10875 l=15225
M1964 N0641 N0637 vss vss efet w=11600 l=10150
M1965 N0642 N0637 vss vss efet w=13050 l=11600
M1966 vcc vcc __FIN_X12_ vss efet w=5800 l=51475
M1967 vss N0578 WRAB1 vss efet w=24650 l=11600
M1968 vss N0649 SC_A12_CLK2 vss efet w=21025 l=12325
M1970 RRAB0 DC vss vss efet w=39150 l=14500
M1971 vcc vcc N0608 vss efet w=5800 l=71050
M1972 vss N0615 RRAB0 vss efet w=36975 l=14500
M1973 vss N0460 CLK2_JMS_DC_M22_BBL_M22_X12_X22__ vss efet w=29725 l=12325
M1974 N0608 clk2 N0615 vss efet w=16675 l=10875
M1975 N0589 X22 vss vss efet w=22475 l=12325
M1976 N0594 N0580 N0588 vss efet w=32625 l=13775
M1977 N0588 FIN_FIM_SRC_JIN N0589 vss efet w=21750 l=12325
M1978 N0595 X12 N0594 vss efet w=29725 l=13775
M1979 N0468 BBL vss vss efet w=23925 l=12325
M1980 N0527 JCN_ISZ N0524 vss efet w=29000 l=11600
M1981 N0524 JUN_JMS N0526 vss efet w=21750 l=11600
M1982 N0468 M22 N0467 vss efet w=25375 l=13775
M1983 N0467 X22 N0468 vss efet w=23200 l=11600
M1984 N0467 X12 N0468 vss efet w=21750 l=13050
M1985 vss INC_ISZ_ADD_SUB_XCH_LD N0595 vss efet w=30450 l=13050
M1986 vss clk2 RRAB0 vss efet w=34800 l=15950
M1987 N0608 X12 N0602 vss efet w=31175 l=15225
M1988 __FIN_X12_ X12 N0639 vss efet w=42775 l=13775
M1989 vcc vcc DC vss efet w=8700 l=24650
M1990 WRAB1 vcc vcc vss efet w=5800 l=33350
M1991 N0547 vcc vcc vss efet w=5800 l=69600
M1992 vcc vcc WRAB0 vss efet w=7250 l=29000
M1993 SC_A12_CLK2 vcc vcc vss efet w=5800 l=36250
M1994 SC_A22_M22_CLK2 S00624 vcc vss efet w=10150 l=27550
M1995 SC_A22_M22_CLK2 N0655 vss vss efet w=37700 l=14500
M1996 N0642 N0610 N0652 vss efet w=24650 l=15950
M1997 N0652 N0653 vss vss efet w=33350 l=11600
M1998 vss N0622 N0621 vss efet w=12325 l=12325
M2000 vcc S00620 N0621 vss efet w=6525 l=54375
M2001 vss N0622 CLK2_SC_A12_M12_ vss efet w=20300 l=11600
M2002 vss N0626 N0627 vss efet w=11600 l=11600
M2004 CLK2_SC_A12_M12_ N0621 vcc vss efet w=18850 l=11600
M2005 __POC__CLK2_SC_A32_X12_ N0627 vss vss efet w=24650 l=11600
M2006 S00624 vcc vcc vss efet w=6525 l=10875
M2007 WRAB0 N0547 vss vss efet w=33350 l=13775
M2008 N0602 _OPA_0 N0614 vss efet w=52925 l=12325
M2009 N0640 _OPA_0 N0639 vss efet w=80475 l=13050
M2010 vss N0636 N0640 vss efet w=42775 l=13775
M2011 vss INC_ISZ_ADD_SUB_XCH_LD N0614 vss efet w=29725 l=12325
M2012 vss SC N0612 vss efet w=29725 l=13775
M2013 DC SC vss vss efet w=60175 l=13050
M2014 vss FIN_FIM_SRC_JIN N0602 vss efet w=21750 l=10150
M2015 N0580 _OPA_0 vss vss efet w=55100 l=11600
M2016 vss DC N0597 vss efet w=30450 l=11600
M2017 N0597 FIN_FIM_SRC_JIN N0596 vss efet w=31175 l=10875
M2018 N0649 vcc vcc vss efet w=5800 l=71050
M2019 vcc vcc N0655 vss efet w=5800 l=71050
M2020 S00620 vcc vcc vss efet w=7250 l=11600
M2021 N0655 clk2 N0656 vss efet w=30450 l=10150
M2022 N0649 clk2 N0650 vss efet w=30450 l=11600
M2023 N0626 S00627 vcc vss efet w=5800 l=52200
M2024 N0612 X32 N0611 vss efet w=36975 l=12325
M2025 N0564 N0590 vss vss efet w=29725 l=14500
M2026 N0524 vcc vcc vss efet w=5800 l=60900
M2027 vss _OPR_3 IO vss efet w=31900 l=12325
M2028 OPE _OPR_3 vss vss efet w=32625 l=10875
M2029 vss DC INC_ISZ vss efet w=24650 l=11600
M2030 N0580 vcc vcc vss efet w=5800 l=27550
M2031 vss N0603 N0568 vss efet w=28275 l=14500
M2032 N0596 _OPA_0 N0590 vss efet w=54375 l=12325
M2033 N0568 vcc vcc vss efet w=5800 l=27550
M2034 N0563 N0564 N0562 vss efet w=34075 l=15950
M2035 vss M12 N0563 vss efet w=34075 l=13050
M2036 N0576 M22 vss vss efet w=31175 l=13775
M2037 N0575 N0564 N0576 vss efet w=30450 l=13050
M2038 N0562 clk2 N0547 vss efet w=34075 l=12325
M2039 N0567 _OPA_0 N0562 vss efet w=53650 l=13775
M2040 N0603 INC_ISZ_XCH N0611 vss efet w=31175 l=12325
M2041 vcc vcc N0603 vss efet w=6525 l=64525
M2042 N0564 vcc vcc vss efet w=5800 l=27550
M2043 N0579 N0568 vss vss efet w=31175 l=13775
M2044 vss N0568 N0567 vss efet w=30450 l=13050
M2045 N0575 N0580 N0579 vss efet w=30450 l=13050
M2046 N0654 SC N0656 vss efet w=32625 l=15225
M2047 N0651 A12 N0650 vss efet w=32625 l=13775
M2048 vss SC N0651 vss efet w=30450 l=14500
M2049 vss M22 N0654 vss efet w=31175 l=15225
M2050 vcc vcc N0622 vss efet w=7250 l=68150
M2051 S00627 vcc vcc vss efet w=6525 l=10875
M2052 vcc vcc N0627 vss efet w=5800 l=52200
M2053 N0622 clk2 N0623 vss efet w=36975 l=10875
M2054 vss M12 N0618 vss efet w=30450 l=11600
M2055 N0682 X12 N0683 vss efet w=84825 l=16675
M2056 N0618 A12 vss vss efet w=36250 l=15225
M2057 vss A22 N0654 vss efet w=29725 l=13775
M2058 N0578 clk2 N0575 vss efet w=31900 l=13050
M2059 vcc vcc N0578 vss efet w=7975 l=67425
M2060 N0590 vcc vcc vss efet w=5800 l=65250
M2061 N0618 SC N0623 vss efet w=34075 l=15225
M2062 vss POC N0683 vss efet w=86275 l=12325
M2063 vcc vcc SC_A22 vss efet w=5800 l=34800
M2064 __POC__CLK2_SC_A32_X12_ N0626 vcc vss efet w=21750 l=10150
M2065 vcc vcc N0679 vss efet w=9425 l=65975
M2066 vcc vcc SC_M22_CLK2 vss efet w=7975 l=25375
M2067 SC_M22_CLK2 N0679 vss vss efet w=37700 l=14500
M2068 N0626 N0630 vss vss efet w=13775 l=10875
M2069 vss POC N0626 vss efet w=16675 l=12325
M2070 N0679 M22 N0680 vss efet w=32625 l=12325
M2071 vss N0643 SC_A22 vss efet w=25375 l=15225
M2072 N0703 clk2 N0682 vss efet w=14500 l=13050
M2073 N0681 clk2 N0680 vss efet w=30450 l=11600
M2074 N0681 SC vss vss efet w=30450 l=11600
M2075 N0629 X12 vss vss efet w=31175 l=12325
M2076 XCH _OPR_3 vss vss efet w=30450 l=15225
M2077 vss _OPR_3 BBL vss efet w=30450 l=13050
M2078 N0628 _OPR_3 vss vss efet w=53650 l=11600
M2079 INC_ISZ_XCH _OPR_3 N0587 vss efet w=47850 l=11600
M2080 LD _OPR_3 vss vss efet w=31175 l=11600
M2081 SUB _OPR_3 vss vss efet w=30450 l=10875
M2082 ADD _OPR_3 vss vss efet w=31175 l=13050
M2083 JCN_ISZ OPR_3 vss vss efet w=50025 l=11600
M2084 vss OPR_3 JCN vss efet w=25375 l=13050
M2085 FIN_FIM OPR_3 vss vss efet w=23925 l=13775
M2086 N0361 vcc vcc vss efet w=6525 l=35525
M2088 vss N0343 SC vss efet w=30450 l=11600
M2089 N0344 N0343 vss vss efet w=29000 l=11600
M2090 vss OPR_3 ISZ vss efet w=24650 l=11600
M2091 vss OPR_3 FIM_SRC vss efet w=23925 l=12325
M2092 vss OPR_3 JIN_FIN vss efet w=44950 l=11600
M2093 JUN_JMS OPR_3 vss vss efet w=44225 l=11600
M2094 vss OPR_3 INC_ISZ vss efet w=23200 l=13050
M2095 ISZ _OPR_2 vss vss efet w=31175 l=11600
M2096 IO _OPR_2 vss vss efet w=29725 l=12325
M2097 OPE _OPR_2 vss vss efet w=31175 l=11600
M2098 JUN_JMS _OPR_2 vss vss efet w=55825 l=13775
M2099 vss OPR_3 JMS vss efet w=24650 l=11600
M2100 vss OPR_3 N0636 vss efet w=23200 l=11600
M2101 LDM_BBL _OPR_3 vss vss efet w=31900 l=13050
M2102 vss A32 N0629 vss efet w=29725 l=13775
M2103 N0629 SC N0631 vss efet w=34075 l=13775
M2104 vss IOR N0683 vss efet w=81925 l=12325
M2105 vss A32 N0682 vss efet w=51475 l=15225
M2106 N0682 M12 vss vss efet w=36975 l=13775
M2107 vss N0703 L vss efet w=52925 l=13775
M2108 L N0703 vss vss efet w=60900 l=14500
M2109 N0631 clk2 N0630 vss efet w=30450 l=8700
M2110 vss M12 N0662 vss efet w=29725 l=10875
M2111 N0662 SC N0661 vss efet w=29725 l=10875
M2112 N0644 A22 N0643 vss efet w=23925 l=9425
M2113 vss SC N0644 vss efet w=23200 l=11600
M2114 N0661 clk2 N0660 vss efet w=30450 l=10150
M2115 N0682 vcc vcc vss efet w=9425 l=35525
M2116 vcc vcc N0630 vss efet w=6525 l=64525
M2117 INC_ISZ_ADD_SUB_XCH_LD OPR_3 N0628 vss efet w=47850 l=13050
M2118 N0587 OPR_3 vss vss efet w=39875 l=13775
M2119 vss _OPR_2 N0523 vss efet w=92075 l=10875
M2120 INC_ISZ _OPR_2 vss vss efet w=30450 l=12325
M2121 BBL _OPR_2 vss vss efet w=30450 l=12325
M2122 N0373 JCN_ISZ N0372 vss efet w=36250 l=15950
M2123 N0372 FIN_FIM N0373 vss efet w=33350 l=14500
M2124 JMS _OPR_2 vss vss efet w=31900 l=11600
M2125 vss OPR_3 FIN_FIM_SRC_JIN vss efet w=24650 l=11600
M2126 vss OPR_3 JUN2_JMS2 vss efet w=24650 l=11600
M2127 N0628 _OPR_2 INC_ISZ_ADD_SUB_XCH_LD vss efet w=56550 l=11600
M2128 N0587 _OPR_2 vss vss efet w=46400 l=13775
M2129 LDM_BBL _OPR_2 vss vss efet w=32625 l=12325
M2130 N0523 OPR_2 JCN_ISZ vss efet w=98600 l=11600
M2131 vss OPR_2 FIN_FIM vss efet w=23200 l=11600
M2132 vss OPR_2 JCN vss efet w=23925 l=13775
M2133 FIM_SRC OPR_2 vss vss efet w=23200 l=11600
M2134 JUN2_JMS2 _OPR_2 vss vss efet w=32625 l=12325
M2135 vss OPR_2 JIN_FIN vss efet w=44950 l=10150
M2136 FIN_FIM _OPR_1 vss vss efet w=31175 l=12325
M2137 ISZ _OPR_1 vss vss efet w=31900 l=13050
M2138 vss OPR_2 XCH vss efet w=23200 l=11600
M2139 vss OPR_2 N0636 vss efet w=23925 l=12325
M2140 N0628 OPR_2 vss vss efet w=46400 l=15950
M2141 OPR_2 N0995 vcc vss efet w=47850 l=20300
M2142 vcc N0994 _OPR_2 vss efet w=33350 l=15950
M2143 N0587 OPR_2 INC_ISZ_XCH vss efet w=40600 l=13050
M2144 vss OPR_2 FIN_FIM_SRC_JIN vss efet w=25375 l=12325
M2145 FIM_SRC _OPR_1 vss vss efet w=29725 l=11600
M2146 IO _OPR_1 vss vss efet w=29725 l=11600
M2147 OPE _OPR_1 vss vss efet w=30450 l=12325
M2148 JIN_FIN _OPR_1 vss vss efet w=53650 l=11600
M2149 INC_ISZ _OPR_1 vss vss efet w=29725 l=10875
M2150 N0523 _OPR_1 vss vss efet w=89175 l=13050
M2151 XCH _OPR_1 vss vss efet w=30450 l=12325
M2152 vss OPR_2 LD vss efet w=24650 l=11600
M2153 vss OPR_2 SUB vss efet w=23200 l=12325
M2154 vss OPR_2 ADD vss efet w=23200 l=11600
M2155 N0628 _OPR_1 INC_ISZ_ADD_SUB_XCH_LD vss efet w=57275 l=14500
M2156 vss _OPR_1 N0587 vss efet w=45675 l=11600
M2157 N0361 clk1 N0343 vss efet w=14500 l=13050
M2158 N0372 X32 vss vss efet w=37700 l=13050
M2159 N0352 vcc vcc vss efet w=7975 l=64525
M2160 vss N0362 N0361 vss efet w=22475 l=10875
M2161 N0373 JUN_JMS N0372 vss efet w=31900 l=13050
M2162 N0368 SC N0373 vss efet w=34800 l=11600
M2163 vss OPR_1 JCN vss efet w=23925 l=12325
M2164 vss OPR_1 JUN_JMS vss efet w=46400 l=13050
M2165 N0636 _OPR_1 vss vss efet w=23200 l=10150
M2166 N0523 OPR_1 JCN_ISZ vss efet w=96425 l=14500
M2167 vss OPR_1 BBL vss efet w=23200 l=11600
M2168 vss OPR_1 JMS vss efet w=26100 l=11600
M2169 INC_ISZ_XCH _OPR_1 N0587 vss efet w=46400 l=13050
M2170 FIN_FIM_SRC_JIN _OPR_1 vss vss efet w=30450 l=12325
M2171 LD _OPR_1 vss vss efet w=31900 l=11600
M2172 vss N0995 _OPR_2 vss efet w=32625 l=13775
M2173 OPR_2 N0994 vss vss efet w=29725 l=13775
M2174 L vcc vcc vss efet w=10150 l=14500
M2175 OPR_3 N0993 vcc vss efet w=39150 l=14500
M2176 vcc N0992 _OPR_3 vss efet w=20300 l=14500
M2177 vcc vcc N0643 vss efet w=7250 l=60900
M2178 N0660 vcc vcc vss efet w=6525 l=63075
M2179 vss N0660 SC_M12_CLK2 vss efet w=36975 l=9425
M2180 SC_M12_CLK2 vcc vcc vss efet w=6525 l=26100
M2181 D0 SC_M12_CLK2 N1011 vss efet w=11600 l=12325
M2182 D2 SC_M12_CLK2 N1009 vss efet w=10875 l=11600
M2183 OPR_3 N0992 vss vss efet w=29725 l=15225
M2184 vss N0993 _OPR_3 vss efet w=20300 l=11600
M2185 N0998 vcc vcc vss efet w=8700 l=30450
M2186 N0994 vcc vcc vss efet w=10150 l=32625
M2187 vss N1011 N0998 vss efet w=58725 l=13775
M2188 vss N1008 N0992 vss efet w=62350 l=11600
M2189 D1 SC_M12_CLK2 N1010 vss efet w=10875 l=12325
M2190 N0996 vcc vcc vss efet w=12325 l=29000
M2191 vss N1009 N0994 vss efet w=61625 l=12325
M2192 N0992 vcc vcc vss efet w=8700 l=33350
M2193 vss OPR_1 SUB vss efet w=23925 l=10875
M2194 vss OPR_1 ADD vss efet w=23925 l=10875
M2195 LDM_BBL OPR_1 vss vss efet w=23925 l=12325
M2196 ISZ _OPR_0 vss vss efet w=31900 l=13050
M2197 JCN _OPR_0 vss vss efet w=31175 l=12325
M2198 OPE _OPR_0 vss vss efet w=30450 l=12325
M2199 JIN_FIN _OPR_0 vss vss efet w=52200 l=10875
M2200 vss X32 N0352 vss efet w=12325 l=12325
M2201 N0367 N0352 vss vss efet w=21750 l=11600
M2202 N0368 N0343 N0367 vss efet w=21750 l=11600
M2203 N0362 clk2 N0368 vss efet w=8700 l=11600
M2204 vcc vcc N0368 vss efet w=6525 l=67425
M2205 XCH _OPR_0 vss vss efet w=29725 l=10875
M2206 vss _OPR_0 JCN_ISZ vss efet w=53650 l=11600
M2207 JMS _OPR_0 vss vss efet w=31175 l=10150
M2208 vss OPR_1 JUN2_JMS2 vss efet w=24650 l=11600
M2209 INC_ISZ_XCH _OPR_0 N0587 vss efet w=52200 l=13050
M2210 N0636 _OPR_0 vss vss efet w=23925 l=12325
M2211 SUB _OPR_0 vss vss efet w=31175 l=12325
M2212 vcc N0998 _OPR_0 vss efet w=39875 l=21750
M2213 vss OPA_0 FIN_FIM vss efet w=21750 l=14500
M2214 vss OPR_0 FIM_SRC vss efet w=25375 l=15225
M2215 vss OPR_0 IO vss efet w=23200 l=11600
M2216 vcc vcc N0769 vss efet w=6525 l=39875
M2217 POC vcc vcc vss efet w=7975 l=22475
M2218 _CN vcc vcc vss efet w=10150 l=28275
M2219 N0769 A12 vss vss efet w=18125 l=12325
M2220 FIN_FIM vcc vcc vss efet w=5800 l=59450
M2221 vss OPR_0 BBL vss efet w=23200 l=11600
M2222 OPR_0 N0999 vcc vss efet w=20300 l=17400
M2223 vss OPR_0 LD vss efet w=24650 l=10150
M2224 vss OPR_0 ADD vss efet w=23200 l=12325
M2225 ISZ vcc vcc vss efet w=7250 l=63800
M2226 JCN vcc vcc vss efet w=5800 l=62350
M2227 FIM_SRC vcc vcc vss efet w=5800 l=63075
M2228 IO vcc vcc vss efet w=9425 l=73225
M2229 N0493 vcc vcc vss efet w=7250 l=72500
M2230 vcc vcc OPE vss efet w=7250 l=56550
M2231 JIN_FIN vcc vcc vss efet w=7250 l=36975
M2232 vcc vcc N0510 vss efet w=7250 l=50750
M2233 JUN_JMS vcc vcc vss efet w=8700 l=39150
M2234 JCN_ISZ vcc vcc vss efet w=8700 l=34800
M2235 INC_ISZ vcc vcc vss efet w=7250 l=55100
M2236 vcc vcc DCL vss efet w=5800 l=63800
M2237 vss OPA_0 N0516 vss efet w=38425 l=10875
M2238 N0516 FIM_SRC _SRC vss efet w=23200 l=13050
M2239 vss SC N0417 vss efet w=33350 l=10150
M2240 vss reset N0327 vss efet w=35525 l=12325
M2241 vss N0397 _CN vss efet w=57275 l=13050
M2242 vss N0327 N0769 vss efet w=19575 l=12325
M2243 POC N0327 vss vss efet w=55825 l=12325
M2244 N0412 N0397 vss vss efet w=21750 l=13050
M2245 N0399 X32 vss vss efet w=13775 l=12325
M2246 N0417 X32 N0418 vss efet w=34075 l=10875
M2247 vss IO N0493 vss efet w=13775 l=11600
M2248 N0510 OPE vss vss efet w=15225 l=12325
M2249 vcc N0510 _OPE vss efet w=29000 l=11600
M2250 vss IO _I_O vss efet w=34800 l=11600
M2251 _I_O N0493 vcc vss efet w=13775 l=12325
M2252 vss ISZ N0456 vss efet w=13050 l=11600
M2253 vss JCN N0476 vss efet w=13775 l=12325
M2254 _OPE OPE vss vss efet w=29725 l=12325
M2255 vcc vcc O_IB vss efet w=7250 l=53650
M2256 vcc vcc KBP vss efet w=5800 l=65975
M2257 vcc vcc TCS vss efet w=8700 l=43500
M2258 vcc vcc DAA vss efet w=8700 l=43500
M2259 XCH vcc vcc vss efet w=5800 l=57275
M2260 BBL vcc vcc vss efet w=6525 l=57275
M2261 JMS vcc vcc vss efet w=7250 l=55100
M2262 N0636 vcc vcc vss efet w=6525 l=60900
M2263 INC_ISZ_ADD_SUB_XCH_LD vcc vcc vss efet w=10150 l=65250
M2264 vcc vcc IOW vss efet w=5800 l=56550
M2265 vcc vcc RAR vss efet w=7250 l=55100
M2266 RAL vcc vcc vss efet w=6525 l=55100
M2267 CMA vcc vcc vss efet w=6525 l=55825
M2268 vcc vcc TCC vss efet w=7250 l=56550
M2269 STC vcc vcc vss efet w=5800 l=61625
M2270 INC_ISZ_XCH vcc vcc vss efet w=5800 l=65250
M2271 LD vcc vcc vss efet w=6525 l=67425
M2272 FIN_FIM_SRC_JIN vcc vcc vss efet w=7250 l=50750
M2273 IOW _I_O vss vss efet w=38425 l=10875
M2274 vcc vcc CMC vss efet w=7250 l=53650
M2275 vcc vcc DAC vss efet w=6525 l=52925
M2276 vcc vcc IAC vss efet w=5800 l=56550
M2277 vcc vcc CLC vss efet w=7250 l=63075
M2278 SUB vcc vcc vss efet w=7250 l=60900
M2279 ADD vcc vcc vss efet w=7250 l=59450
M2280 LDM_BBL vcc vcc vss efet w=7975 l=58725
M2281 JUN2_JMS2 vcc vcc vss efet w=7250 l=63800
M2282 vcc vcc CLB vss efet w=7975 l=65250
M2283 vcc vcc SBM vss efet w=7250 l=56550
M2284 ADM vcc vcc vss efet w=5800 l=56550
M2285 OPR_0 N0998 vss vss efet w=21025 l=12325
M2286 vss N0999 _OPR_0 vss efet w=29725 l=12325
M2287 _OPR_1 N0996 vcc vss efet w=38425 l=15950
M2288 vcc N0997 OPR_1 vss efet w=24650 l=13050
M2289 N0999 N0998 vss vss efet w=27550 l=11600
M2290 vss N1010 N0996 vss efet w=58000 l=11600
M2291 N0995 N0994 vss vss efet w=29000 l=11600
M2292 N0997 N0996 vss vss efet w=29000 l=10150
M2293 D3 SC_M12_CLK2 N1008 vss efet w=10150 l=12325
M2294 N0993 N0992 vss vss efet w=26825 l=10875
M2295 N0999 vcc vcc vss efet w=13050 l=42050
M2296 _OPR_1 N0997 vss vss efet w=34075 l=13050
M2297 vss N0996 OPR_1 vss efet w=24650 l=11600
M2298 N0995 vcc vcc vss efet w=14500 l=43500
M2299 N0997 vcc vcc vss efet w=9425 l=36975
M2300 N0993 vcc vcc vss efet w=15950 l=38425
M2301 D3 OPA_IB OPA_3 vss efet w=58725 l=13775
M2302 vcc vcc IOR vss efet w=10875 l=41325
M2303 SBM _I_O vss vss efet w=31900 l=13050
M2304 ADM _I_O vss vss efet w=31900 l=12325
M2305 vcc vcc N0477 vss efet w=5800 l=49300
M2306 vss __X31__CLK2_ N0480 vss efet w=13775 l=12325
M2307 N0480 vcc vcc vss efet w=7250 l=67425
M2308 N0482 N0480 N0477 vss efet w=27550 l=11600
M2309 N0479 vcc vcc vss efet w=7250 l=77575
M2310 N0482 N0479 vss vss efet w=26825 l=10875
M2311 N0479 IOR vss vss efet w=12325 l=10150
M2312 N0412 N0399 N0413 vss efet w=20300 l=11600
M2313 N0418 N0419 N0413 vss efet w=30450 l=10150
M2314 vss N0769 N0327 vss efet w=33350 l=11600
M2315 N0297 clk2 vss vss efet w=26100 l=11600
M2317 X22 clk2 N0280 vss efet w=13775 l=12325
M2318 vcc S00678 N0297 vss efet w=7975 l=32625
M2319 vcc vcc S00678 vss efet w=5800 l=13050
M2320 N0295 N0297 N0296 vss efet w=27550 l=11600
M2321 N0296 N0280 vss vss efet w=62350 l=13050
M2322 vcc vcc N0296 vss efet w=7975 l=21025
M2323 N0739 clk1 N0296 vss efet w=11600 l=11600
M2324 N0404 clk1 N0397 vss efet w=14500 l=11600
M2325 vss N0405 N0404 vss efet w=26825 l=12325
M2326 N0413 clk2 N0405 vss efet w=8700 l=11600
M2327 vcc vcc N0399 vss efet w=7250 l=84100
M2328 vss test N0432 vss efet w=36250 l=10150
M2329 vcc vcc N0432 vss efet w=7250 l=55100
M2330 N0327 vcc vcc vss efet w=5800 l=26100
M2331 vcc vcc N0404 vss efet w=7250 l=36250
M2332 vcc vcc N0784 vss efet w=5800 l=50750
M2333 N0741 N0739 vss vss efet w=31900 l=10875
M2334 vcc vcc N0329 vss efet w=8700 l=20300
M2335 N0413 vcc vcc vss efet w=6525 l=63075
M2336 N0456 vcc vcc vss efet w=10875 l=65975
M2337 vss N0476 N0478 vss efet w=23200 l=11600
M2338 vss _OPE DCL vss efet w=23200 l=11600
M2339 O_IB _OPE vss vss efet w=23200 l=12325
M2340 vss _OPE KBP vss efet w=23925 l=12325
M2341 vss _OPE TCS vss efet w=38425 l=10875
M2342 DAA _OPE vss vss efet w=34075 l=12325
M2343 RAR _OPE vss vss efet w=23925 l=10875
M2344 vss _OPE RAL vss efet w=23925 l=10875
M2345 vss _OPE CMA vss efet w=25375 l=10875
M2346 N0478 N0487 N0481 vss efet w=44225 l=15225
M2347 N0478 _OPA_3 N0481 vss efet w=63800 l=13050
M2348 N0478 N0456 N0419 vss efet w=41325 l=13775
M2349 vss _I_O N0329 vss efet w=59450 l=11600
M2350 N0476 vcc vcc vss efet w=5800 l=58000
M2351 N0478 ADD_0 N0419 vss efet w=47125 l=13050
M2352 N0419 vcc vcc vss efet w=5800 l=50025
M2353 vcc vcc _SRC vss efet w=5800 l=68875
M2354 DCL _OPA_3 vss vss efet w=30450 l=10875
M2355 KBP _OPA_3 vss vss efet w=30450 l=11600
M2356 TCS _OPA_3 vss vss efet w=40600 l=11600
M2357 DAA _OPA_3 vss vss efet w=40600 l=13775
M2358 vss N0486 N0481 vss efet w=50750 l=14500
M2359 vss OPA_3 N0481 vss efet w=75400 l=13050
M2360 vss _OPE TCC vss efet w=23200 l=11600
M2361 STC _OPE vss vss efet w=23925 l=12325
M2362 vss _OPE CMC vss efet w=23925 l=12325
M2363 vss _OPE DAC vss efet w=23200 l=13050
M2364 vss _OPE IAC vss efet w=23925 l=12325
M2365 vss _I_O IOR vss efet w=39875 l=10875
M2366 N0477 A12 N0483 vss efet w=31900 l=11600
M2367 D2 OPA_IB OPA_2 vss efet w=61625 l=16675
M2368 vss IOR N0483 vss efet w=31175 l=15225
M2369 vss _OPE CLC vss efet w=23200 l=10150
M2370 CLB _OPE vss vss efet w=23200 l=11600
M2371 STC _OPA_3 vss vss efet w=31175 l=13050
M2372 DAC _OPA_3 vss vss efet w=30450 l=10875
M2373 SBM _OPA_3 vss vss efet w=32625 l=11600
M2374 ADM _OPA_3 vss vss efet w=30450 l=13775
M2375 IOR _OPA_3 vss vss efet w=44950 l=11600
M2376 vss N1001 _OPA_3 vss efet w=29725 l=11600
M2377 OPA_3 N1000 vss vss efet w=57275 l=12325
M2378 vss OPA_3 O_IB vss efet w=23200 l=12325
M2379 vss OPA_3 IOW vss efet w=31900 l=10150
M2380 vss OPA_3 RAR vss efet w=24650 l=10150
M2381 vss OPA_3 RAL vss efet w=23925 l=10875
M2382 vss OPA_3 CMA vss efet w=23200 l=10150
M2383 vss OPA_3 TCC vss efet w=23200 l=10150
M2384 vss OPA_3 CMC vss efet w=24650 l=11600
M2385 vss OPA_3 IAC vss efet w=23925 l=10875
M2386 vss N0486 N0487 vss efet w=13050 l=11600
M2387 DCL _OPA_2 vss vss efet w=30450 l=10875
M2388 vss OPA_2 N0501 vss efet w=44950 l=14500
M2389 N0501 ACC_0 N0486 vss efet w=29000 l=10875
M2390 N0487 vcc vcc vss efet w=5800 l=50750
M2391 vcc vcc N0398 vss efet w=6525 l=26100
M2392 KBP _OPA_2 vss vss efet w=30450 l=10875
M2393 RAR _OPA_2 vss vss efet w=31900 l=12325
M2394 RAL _OPA_2 vss vss efet w=31175 l=13050
M2395 vss OPA_3 CLC vss efet w=23200 l=11600
M2396 vss OPA_3 CLB vss efet w=24650 l=11600
M2397 CMA _OPA_2 vss vss efet w=30450 l=11600
M2398 TCC _OPA_2 vss vss efet w=31175 l=11600
M2399 N0486 vcc vcc vss efet w=5800 l=47850
M2400 vss OPA_2 TCS vss efet w=34075 l=13775
M2401 vss OPA_2 DAA vss efet w=34800 l=11600
M2402 vss N1003 _OPA_2 vss efet w=36975 l=15225
M2403 OPA_2 N1002 vss vss efet w=54375 l=15950
M2404 vcc N1000 _OPA_3 vss efet w=22475 l=10875
M2405 OPA_3 N1001 vcc vss efet w=25375 l=9425
M2406 vss OPA_2 STC vss efet w=23200 l=10150
M2407 vss OPA_2 CMC vss efet w=24650 l=10150
M2408 vss OPA_2 DAC vss efet w=23925 l=11600
M2409 vss OPA_2 IAC vss efet w=27550 l=10150
M2410 vss OPA_2 CLC vss efet w=27550 l=10150
M2411 CLB OPA_2 vss vss efet w=23200 l=13050
M2412 DAA _OPA_1 vss vss efet w=43500 l=10875
M2413 vss clk2 N0398 vss efet w=47850 l=10150
M2414 vcc vcc N0799 vss efet w=6525 l=67425
M2416 vcc S00690 N0741 vss efet w=6525 l=26825
M2417 vcc vcc S00690 vss efet w=5800 l=13050
M2418 X32 N0739 vss vss efet w=31900 l=11600
M2419 vss N0782 N0784 vss efet w=14500 l=11600
M2420 vcc N0741 X32 vss efet w=36250 l=12325
M2421 N0414 clk2 A22 vss efet w=8700 l=11600
M2422 N0799 _SRC vss vss efet w=13050 l=13050
M2423 N0407 N0414 vss vss efet w=14500 l=11600
M2424 N0407 N0398 N0408 vss efet w=8700 l=13050
M2425 vcc vcc S00685 vss efet w=6525 l=11600
M2426 vcc S00685 N0415 vss efet w=5800 l=16675
M2428 N0507 CY_1 N0486 vss efet w=27550 l=11600
M2429 RAR _OPA_1 vss vss efet w=31175 l=10150
M2430 TCC _OPA_1 vss vss efet w=30450 l=11600
M2431 vss OPA_1 N0507 vss efet w=45675 l=13050
M2432 STC _OPA_1 vss vss efet w=31900 l=11600
M2433 CMC _OPA_1 vss vss efet w=31175 l=12325
M2434 IAC _OPA_1 vss vss efet w=31900 l=11600
M2435 vss OPA_2 SBM vss efet w=28275 l=10875
M2436 vss OPA_2 ADM vss efet w=26100 l=11600
M2437 ADM _OPA_1 vss vss efet w=29725 l=12325
M2438 _COM N0782 vcc vss efet w=20300 l=11600
M2439 vss N0784 _COM vss efet w=20300 l=11600
M2440 N0800 N0801 N0782 vss efet w=30450 l=10150
M2441 vss N0329 N0800 vss efet w=27550 l=11600
M2442 N0798 N0805 vss vss efet w=27550 l=11600
M2443 N0782 N0799 N0798 vss efet w=29725 l=12325
M2444 vss N0797 N0782 vss efet w=15225 l=12325
M2445 vss clk2 N0375 vss efet w=16675 l=12325
M2446 N0797 N0408 vss vss efet w=20300 l=12325
M2447 vcc vcc N0797 vss efet w=7975 l=55100
M2448 vcc N0742 X22 vss efet w=39150 l=13050
M2449 X22 N0719 vss vss efet w=36975 l=12325
M2450 vss X22 N0288 vss efet w=25375 l=13775
M2451 N0742 N0719 vss vss efet w=30450 l=11600
M2453 vcc vcc S00710 vss efet w=6525 l=13775
M2454 vcc S00710 N0742 vss efet w=7250 l=27550
M2455 N0718 N0281 vss vss efet w=26825 l=10875
M2456 N0281 clk2 X12 vss efet w=13050 l=13775
M2457 N0719 clk1 N0718 vss efet w=14500 l=11600
M2458 vcc vcc N0718 vss efet w=8700 l=37700
M2459 N0383 X22 vss vss efet w=14500 l=11600
M2461 N0288 X12 vss vss efet w=21750 l=13775
M2462 vcc N0743 X12 vss efet w=35525 l=12325
M2463 X12 N0721 vss vss efet w=36975 l=12325
M2465 N0743 N0721 vss vss efet w=26100 l=10875
M2466 vcc vcc S00725 vss efet w=5800 l=11600
M2467 vcc S00725 N0743 vss efet w=7975 l=26825
M2468 vcc S00699 N0782 vss efet w=5800 l=39875
M2469 N0380 clk2 N0383 vss efet w=8700 l=11600
M2470 vcc vcc N0407 vss efet w=5800 l=49300
M2471 vss OPA_1 DCL vss efet w=24650 l=13050
M2472 vss OPA_1 KBP vss efet w=29000 l=11600
M2473 vss OPA_1 TCS vss efet w=33350 l=11600
M2474 vss OPA_1 RAL vss efet w=23925 l=12325
M2475 vss OPA_1 CMA vss efet w=24650 l=10875
M2476 vss OPA_1 DAC vss efet w=23200 l=10150
M2477 vss OPA_1 CLC vss efet w=23200 l=10150
M2478 vss OPA_1 CLB vss efet w=24650 l=13050
M2479 vss OPA_1 SBM vss efet w=23925 l=13050
M2480 N0512 N0432 N0486 vss efet w=27550 l=11600
M2481 vss OPA_0 N0512 vss efet w=49300 l=14500
M2482 DCL _OPA_0 vss vss efet w=30450 l=11600
M2483 TCS _OPA_0 vss vss efet w=42050 l=10875
M2484 DAA _OPA_0 vss vss efet w=41325 l=11600
M2485 RAL _OPA_0 vss vss efet w=31175 l=13775
M2486 TCC _OPA_0 vss vss efet w=30450 l=11600
M2487 CMC _OPA_0 vss vss efet w=31900 l=11600
M2488 CLC _OPA_0 vss vss efet w=31175 l=10150
M2489 ADM _OPA_0 vss vss efet w=29725 l=11600
M2490 vss OPA_0 KBP vss efet w=24650 l=10150
M2491 vss OPA_0 RAR vss efet w=24650 l=11600
M2492 vss OPA_0 DAC vss efet w=26100 l=13050
M2493 vcc N1002 _OPA_2 vss efet w=14500 l=11600
M2494 OPA_1 N1004 vss vss efet w=68875 l=12325
M2495 vss OPA_0 CMA vss efet w=23200 l=11600
M2496 vss OPA_0 STC vss efet w=23200 l=10875
M2497 vss OPA_0 IAC vss efet w=23200 l=10150
M2498 vss OPA_0 CLB vss efet w=24650 l=11600
M2499 vss OPA_0 SBM vss efet w=24650 l=10150
M2500 vss _OPE N0415 vss efet w=44225 l=10875
M2501 vss N0353 N0351 vss efet w=22475 l=10875
M2502 N0351 __X21__CLK2_ vss vss efet w=20300 l=11600
M2503 vss DCL N0353 vss efet w=14500 l=10150
M2504 WRITE_ACC_1_ KBP vss vss efet w=14500 l=10150
M2505 N0415 __X21__CLK2_ vss vss efet w=44225 l=10875
M2506 vcc vcc N0383 vss efet w=5800 l=47850
M2507 N0375 N0380 vss vss efet w=21750 l=13775
M2508 vcc vcc __X31__CLK2_ vss efet w=5800 l=15950
M2509 N0353 vcc vcc vss efet w=6525 l=64525
M2510 vss TCS WRITE_ACC_1_ vss efet w=13050 l=11600
M2511 WRITE_ACC_1_ DAA vss vss efet w=13050 l=11600
M2512 S00699 vcc vcc vss efet w=5800 l=11600
M2513 vcc vcc __X21__CLK2_ vss efet w=6525 l=18850
M2514 __X31__CLK2_ N0375 vss vss efet w=65250 l=11600
M2515 N0375 vcc vcc vss efet w=5800 l=36250
M2516 N0369 vcc vcc vss efet w=5800 l=56550
M2517 N0337 vcc vcc vss efet w=5800 l=29000
M2518 vcc vcc N0328 vss efet w=6525 l=64525
M2519 N0720 N0282 vss vss efet w=26825 l=10875
M2520 N0282 clk2 M22 vss efet w=15950 l=11600
M2521 N0721 clk1 N0720 vss efet w=14500 l=11600
M2522 vcc vcc N0720 vss efet w=7250 l=30450
M2523 N0337 N0360 vss vss efet w=34800 l=12325
M2524 vss clk2 N0337 vss efet w=28275 l=12325
M2525 __X21__CLK2_ N0337 vss vss efet w=53650 l=11600
M2526 vss N0329 N0328 vss efet w=13775 l=12325
M2527 N0328 POC vss vss efet w=11600 l=11600
M2528 N0330 X22 N0331 vss efet w=29000 l=13050
M2529 vss clk2 N0330 vss efet w=29725 l=13775
M2530 N0369 X12 vss vss efet w=15225 l=12325
M2531 N0360 clk2 N0369 vss efet w=9425 l=12325
M2532 N0335 clk1 vss vss efet w=31175 l=12325
M2533 N0336 N0337 N0335 vss efet w=31175 l=10875
M2534 N0332 N0328 N0336 vss efet w=29725 l=12325
M2535 N0331 N0329 N0332 vss efet w=30450 l=10875
M2536 vss clk2 N0423 vss efet w=21750 l=13050
M2537 N0332 POC N0331 vss efet w=29000 l=11600
M2538 N0351 vcc vcc vss efet w=7250 l=43500
M2539 vss INC_ISZ N0442 vss efet w=15950 l=10150
M2540 N0442 vcc vcc vss efet w=6525 l=58725
M2541 vss TCS WRITE_CARRY_2_ vss efet w=11600 l=11600
M2542 vss TCS ADD_GROUP_4_ vss efet w=12325 l=12325
M2543 READ_ACC_3_ DAA vss vss efet w=13050 l=11600
M2544 vss N0446 N0448 vss efet w=76125 l=10875
M2545 N0342 N0332 vcc vss efet w=21025 l=11600
M2546 vcc vcc N0423 vss efet w=6525 l=31175
M2547 vss M22 N0288 vss efet w=22475 l=13775
M2548 vcc N0744 M22 vss efet w=40600 l=11600
M2549 M22 N0723 vss vss efet w=34800 l=11600
M2551 N0744 N0723 vss vss efet w=27550 l=13050
M2552 vcc vcc S00740 vss efet w=5800 l=11600
M2553 vcc S00740 N0744 vss efet w=4350 l=31175
M2554 vcc vcc N0430 vss efet w=5800 l=49300
M2555 N0340 vcc vcc vss efet w=7250 l=72500
M2556 N0430 N0423 N0431 vss efet w=10150 l=10875
M2557 N0722 N0283 vss vss efet w=26825 l=10875
M2558 N0283 clk2 M12 vss efet w=13775 l=15225
M2559 N0723 clk1 N0722 vss efet w=14500 l=11600
M2560 M12 clk2 N0433 vss efet w=8700 l=12325
M2561 N0342 N0340 vss vss efet w=20300 l=13050
M2562 vss N0332 N0340 vss efet w=11600 l=11600
M2563 vcc S00731 N0332 vss efet w=6525 l=52925
M2564 S00731 vcc vcc vss efet w=6525 l=12325
M2566 vcc vcc N0805 vss efet w=11600 l=54375
M2567 N0853 vcc vcc vss efet w=7975 l=67425
M2568 X12 clk2 N0425 vss efet w=7975 l=13050
M2569 N0421 vcc vcc vss efet w=5800 l=56550
M2570 N0421 N0423 N0422 vss efet w=10875 l=10875
M2571 vss N0422 N0805 vss efet w=31175 l=10150
M2572 N0853 X12 vss vss efet w=13050 l=11600
M2573 vss N0433 N0430 vss efet w=15225 l=12325
M2574 vss N0425 N0421 vss efet w=15225 l=10875
M2575 N0801 vcc vcc vss efet w=6525 l=51475
M2576 vcc vcc N0722 vss efet w=7975 l=38425
M2577 vss N0431 N0801 vss efet w=23925 l=13775
M2578 N0288 M12 vss vss efet w=21750 l=13050
M2579 vcc N0745 M12 vss efet w=39150 l=21750
M2580 vss N0803 N0403 vss efet w=24650 l=10150
M2581 M12 N0725 vss vss efet w=38425 l=12325
M2583 vss POC N0717 vss efet w=70325 l=12325
M2584 N0717 S00757 vcc vss efet w=10150 l=15950
M2586 N0403 N0802 vss vss efet w=21750 l=11600
M2587 vss __X21__CLK2_ N0448 vss efet w=73950 l=11600
M2588 vss XCH WRITE_ACC_1_ vss efet w=13050 l=11600
M2589 WRITE_ACC_1_ POC vss vss efet w=13050 l=11600
M2590 INC_GROUP_5_ INC_ISZ vss vss efet w=11600 l=12325
M2591 WRITE_CARRY_2_ POC vss vss efet w=15950 l=13050
M2592 vss CMA WRITE_ACC_1_ vss efet w=13050 l=11600
M2593 WRITE_ACC_1_ TCC vss vss efet w=13775 l=10875
M2594 vss DAC WRITE_ACC_1_ vss efet w=11600 l=10150
M2595 WRITE_ACC_1_ IAC vss vss efet w=11600 l=10150
M2596 vss N1005 _OPA_1 vss efet w=34075 l=15225
M2597 WRITE_ACC_1_ CLB vss vss efet w=12325 l=10875
M2598 vcc N1004 _OPA_1 vss efet w=30450 l=26100
M2599 OPA_1 N1005 vcc vss efet w=26825 l=16675
M2600 vss LD WRITE_ACC_1_ vss efet w=14500 l=11600
M2601 WRITE_ACC_1_ SUB vss vss efet w=15225 l=10875
M2602 vss ADD WRITE_ACC_1_ vss efet w=13775 l=10875
M2603 WRITE_ACC_1_ LDM_BBL vss vss efet w=13775 l=10875
M2604 WRITE_CARRY_2_ SUB vss vss efet w=16675 l=13775
M2605 WRITE_CARRY_2_ TCC vss vss efet w=13050 l=11600
M2606 vss STC WRITE_CARRY_2_ vss efet w=13050 l=11600
M2607 WRITE_CARRY_2_ CMC vss vss efet w=13050 l=11600
M2608 vss DAC WRITE_CARRY_2_ vss efet w=13775 l=11600
M2609 WRITE_CARRY_2_ IAC vss vss efet w=15225 l=10875
M2610 vss CLC WRITE_CARRY_2_ vss efet w=13050 l=11600
M2611 WRITE_CARRY_2_ CLB vss vss efet w=13775 l=12325
M2612 vss SBM WRITE_CARRY_2_ vss efet w=13050 l=10150
M2613 WRITE_CARRY_2_ ADM vss vss efet w=13775 l=10150
M2614 vss RAR READ_ACC_3_ vss efet w=13050 l=11600
M2615 READ_ACC_3_ RAL vss vss efet w=13050 l=11600
M2616 N0448 N0445 ACB_IB vss efet w=74675 l=10875
M2617 ACB_IB __X31__CLK2_ N0448 vss efet w=76125 l=10875
M2618 vss N0442 ADD_IB vss efet w=39150 l=12325
M2619 vss XCH N0445 vss efet w=21750 l=11600
M2620 vss N0446 CY_IB vss efet w=14500 l=11600
M2621 vss IOW N0446 vss efet w=21750 l=11600
M2622 ADD_GROUP_4_ TCC vss vss efet w=13050 l=13050
M2623 READ_ACC_3_ IAC vss vss efet w=12325 l=14500
M2624 vss DAC READ_ACC_3_ vss efet w=12325 l=10875
M2625 vss SBM READ_ACC_3_ vss efet w=11600 l=10150
M2627 vss STC INC_GROUP_5_ vss efet w=11600 l=11600
M2628 N0502 RAL vss vss efet w=15225 l=10875
M2629 CY_IB __X31__CLK2_ vss vss efet w=15950 l=12325
M2630 SUB_GROUP_6_ CMC vss vss efet w=23925 l=15225
M2631 SUB_GROUP_6_ S00709 vcc vss efet w=5800 l=40600
M2632 INC_GROUP_5_ IAC vss vss efet w=14500 l=13050
M2633 INC_GROUP_5_ vcc vcc vss efet w=7250 l=66700
M2634 READ_ACC_3_ vcc vcc vss efet w=7250 l=69600
M2635 vss RAR N0490 vss efet w=15225 l=15225
M2636 vss __X31__CLK2_ ADSL vss efet w=17400 l=10875
M2637 vss __X31__CLK2_ ADD_IB vss efet w=38425 l=10875
M2639 ADD_IB S00729 vcc vss efet w=8700 l=24650
M2641 N0445 vcc vcc vss efet w=8700 l=41325
M2642 vss N0502 ADSL vss efet w=13050 l=13050
M2643 CY_IB vcc vcc vss efet w=7975 l=70325
M2644 N0446 vcc vcc vss efet w=8700 l=43500
M2645 vss __X31__CLK2_ ADSR vss efet w=14500 l=11600
M2646 ADSR N0490 vss vss efet w=15950 l=14500
M2647 vss CMA N0515 vss efet w=11600 l=11600
M2648 vcc vcc S00709 vss efet w=6525 l=13775
M2649 ACB_IB S00724 vcc vss efet w=10875 l=29725
M2650 vcc vcc ADSL vss efet w=8700 l=65250
M2651 N0502 vcc vcc vss efet w=5800 l=60900
M2652 vcc vcc N0490 vss efet w=7975 l=84825
M2653 ADSR vcc vcc vss efet w=7250 l=65250
M2654 ACC_ADAC N0515 vss vss efet w=13775 l=11600
M2655 vss N0342 ACC_ADAC vss efet w=13050 l=13050
M2656 WRITE_CARRY_2_ vcc vcc vss efet w=6525 l=63800
M2657 N0515 vcc vcc vss efet w=7250 l=84100
M2658 vss N0853 N0854 vss efet w=19575 l=13775
M2659 READ_ACC_3_ ADM vss vss efet w=13050 l=13050
M2660 ADD_GROUP_4_ ADM vss vss efet w=12325 l=16675
M2661 vss SBM SUB_GROUP_6_ vss efet w=21750 l=13050
M2662 ADD_GROUP_4_ vcc vcc vss efet w=6525 l=60175
M2663 vss ADD WRITE_CARRY_2_ vss efet w=13050 l=11600
M2664 READ_ACC_3_ SUB vss vss efet w=13050 l=13050
M2665 vss IOR WRITE_ACC_1_ vss efet w=13050 l=11600
M2666 vss ADD READ_ACC_3_ vss efet w=13775 l=12325
M2667 vss ADD ADD_GROUP_4_ vss efet w=13050 l=11600
M2668 SUB_GROUP_6_ SUB vss vss efet w=23200 l=11600
M2669 vcc vcc N1001 vss efet w=13050 l=37700
M2670 OPA_2 N1003 vcc vss efet w=32625 l=25375
M2671 N1001 N1000 vss vss efet w=27550 l=14500
M2672 vcc vcc N1005 vss efet w=13050 l=33350
M2673 D1 OPA_IB OPA_1 vss efet w=58725 l=18125
M2674 vss clk2 N0702 vss efet w=54375 l=12325
M2676 S00676 vcc vcc vss efet w=8700 l=15950
M2677 vcc vcc N0671 vss efet w=13050 l=33350
M2678 D0 OPA_IB OPA_0 vss efet w=65250 l=13050
M2679 vss N1007 _OPA_0 vss efet w=37700 l=14500
M2680 OPA_0 N1006 vss vss efet w=70325 l=12325
M2681 N0702 S00676 vcc vss efet w=13050 l=15950
M2682 N0671 N0702 N0688 vss efet w=27550 l=13775
M2683 N0671 D3 vss vss efet w=53650 l=13050
M2684 vcc N1006 _OPA_0 vss efet w=52925 l=25375
M2685 OPA_0 N1007 vcc vss efet w=29000 l=15225
M2686 vcc vcc N1003 vss efet w=12325 l=35525
M2687 N1005 N1004 vss vss efet w=26825 l=14500
M2688 vss N1012 N1000 vss efet w=56550 l=13050
M2689 vss N1014 N1004 vss efet w=55825 l=12325
M2690 vss JUN2_JMS2 N0658 vss efet w=15225 l=12325
M2691 N1003 N1002 vss vss efet w=26100 l=15225
M2692 vcc vcc N1007 vss efet w=9425 l=35525
M2693 N1007 N1006 vss vss efet w=34800 l=12325
M2694 vss N1013 N1002 vss efet w=57275 l=12325
M2695 vss N1015 N1006 vss efet w=64525 l=12325
M2696 vcc vcc S00689 vss efet w=8700 l=11600
M2697 S00687 vcc vcc vss efet w=8700 l=17400
M2699 N0687 S00687 vcc vss efet w=10150 l=14500
M2700 vcc S00689 N0689 vss efet w=10150 l=11600
M2702 vcc N0659 D0 vss efet w=47125 l=18125
M2703 N0687 N0700 vss vss efet w=253750 l=11600
M2704 vss N0700 N0689 vss efet w=228375 l=10875
M2705 N0687 N0688 vss vss efet w=98600 l=11600
M2706 vss N0687 N0689 vss efet w=74675 l=5800
M2707 D0 SC_M22_CLK2 N1015 vss efet w=10150 l=13050
M2708 vcc N0659 D2 vss efet w=47125 l=16675
M2709 N1000 vcc vcc vss efet w=19575 l=42050
M2710 N0658 LDM_BBL vss vss efet w=14500 l=10875
M2711 WRITE_ACC_1_ vcc vcc vss efet w=6525 l=71775
M2712 N1004 vcc vcc vss efet w=11600 l=30450
M2713 N1002 vcc vcc vss efet w=19575 l=42050
M2714 N1006 vcc vcc vss efet w=20300 l=40600
M2715 D2 SC_M22_CLK2 N1013 vss efet w=10875 l=13775
M2716 vss N0689 d3 vss efet w=1246275 l=6525
M2717 vss N0658 OPA_IB vss efet w=42050 l=15950
M2718 vcc vcc N0658 vss efet w=7250 l=69600
M2719 OPA_IB __X21__CLK2_ vss vss efet w=41325 l=10875
M2720 D1 SC_M22_CLK2 N1014 vss efet w=10875 l=13775
M2721 d3 N0687 vcc vss efet w=657575 l=10875
M2723 D3 SC_M22_CLK2 N1012 vss efet w=10150 l=11600
M2724 vcc S00716 OPA_IB vss efet w=8700 l=20300
M2725 D1 N0659 vcc vss efet w=46400 l=13050
M2726 D3 N0659 vcc vss efet w=39875 l=12325
M2727 vcc vcc S00716 vss efet w=7250 l=11600
M2728 N0675 vcc vcc vss efet w=7975 l=36250
M2729 N0659 vcc vcc vss efet w=11600 l=21025
M2730 N0659 N0675 vss vss efet w=53650 l=10150
M2731 vcc vcc N0678 vss efet w=11600 l=37700
M2732 vss INC_GROUP_5_ N0546 vss efet w=11600 l=12325
M2733 N0701 vcc vcc vss efet w=7250 l=20300
M2734 vss L N0686 vss efet w=57275 l=15225
M2735 vss L N0701 vss efet w=42775 l=10875
M2736 vcc vcc N0546 vss efet w=13050 l=87000
M2737 N0546 N0342 vss vss efet w=12325 l=14500
M2738 vss SUB_GROUP_6_ CY_ADAC vss efet w=14500 l=11600
M2739 vss ADD_GROUP_4_ CY_ADA vss efet w=11600 l=10875
M2740 vcc vcc N0677 vss efet w=8700 l=34075
M2741 N0685 clk1 N0701 vss efet w=21025 l=18850
M2742 CY_1 ADSR N0513 vss efet w=14500 l=11600
M2743 S00729 vcc vcc vss efet w=5800 l=11600
M2744 S00724 vcc vcc vss efet w=6525 l=15225
M2745 CY N0415 N0860 vss efet w=15950 l=10150
M2746 N0860 N0403 vcc vss efet w=13775 l=13050
M2748 CY M12 N0470 vss efet w=7975 l=12325
M2749 N0550 CY_ADA N0470 vss efet w=14500 l=11600
M2750 N0470 vcc vcc vss efet w=10150 l=34800
M2751 N0470 N0855 vss vss efet w=41325 l=11600
M2752 N0513 ADSL CY vss efet w=14500 l=11600
M2753 D0 CY_IB CY_1 vss efet w=57275 l=10150
M2754 vss N0342 CY_ADAC vss efet w=13775 l=13775
M2756 N0861 ADC_CY CY vss efet w=10150 l=13050
M2757 vss CY N0855 vss efet w=59450 l=11600
M2758 N0855 vcc vcc vss efet w=10150 l=33350
M2759 N0846 ADSR CY vss efet w=7250 l=11600
M2760 CY_ADAC S00732 vcc vss efet w=6525 l=48575
M2761 vss N0342 CY_ADA vss efet w=13050 l=11600
M2762 vss READ_ACC_3_ ACC_ADA vss efet w=14500 l=11600
M2763 vss N0342 ACC_ADA vss efet w=15225 l=14500
M2764 vss WRITE_CARRY_2_ ADC_CY vss efet w=13775 l=10875
M2765 vss WRITE_ACC_1_ ADD_ACC vss efet w=15225 l=11600
M2766 N0678 clk1 vss vss efet w=22475 l=12325
M2767 N0686 clk1 N0675 vss efet w=46400 l=11600
M2768 vss N0678 N0677 vss efet w=29000 l=15950
M2769 vss N0699 N0678 vss efet w=24650 l=14500
M2770 N0701 N0702 N0699 vss efet w=10150 l=11600
M2771 N0676 N0677 vcc vss efet w=41325 l=14500
M2772 N0678 N0685 vss vss efet w=23200 l=11600
M2773 vss N0678 N0676 vss efet w=45675 l=12325
M2774 vss N0477 ADC_CY vss efet w=13050 l=13050
M2775 vss N0477 ADD_ACC vss efet w=14500 l=13050
M2776 ADD_ACC vcc vcc vss efet w=10150 l=65250
M2777 vcc S00734 CY_ADA vss efet w=5800 l=58000
M2778 ADC_CY vcc vcc vss efet w=8700 l=79750
M2779 S00734 vcc vcc vss efet w=7250 l=11600
M2780 S00732 vcc vcc vss efet w=7975 l=10150
M2781 L clk1 N0707 vss efet w=10875 l=13050
M2782 N0675 clk2 N0684 vss efet w=44950 l=15950
M2783 N0684 N0685 vss vss efet w=56550 l=8700
M2784 N0705 N0707 vss vss efet w=59450 l=9425
M2785 N0705 L N0706 vss efet w=126150 l=13050
M2786 vss POC N0705 vss efet w=60175 l=11600
M2787 N0706 N0702 vss vss efet w=96425 l=10875
M2788 N0705 vcc vcc vss efet w=15225 l=27550
M2789 vss N0705 N0704 vss efet w=37700 l=15950
M2790 vss M12 N0550 vss efet w=10150 l=10150
M2791 N0550 N0546 vcc vss efet w=9425 l=15225
M2792 vss N0452 CY_1 vss efet w=53650 l=10150
M2793 CY_1 vcc vcc vss efet w=6525 l=29000
M2794 N0855 N0854 N0452 vss efet w=8700 l=10150
M2795 N0550 CY_ADAC N0855 vss efet w=15950 l=13050
M2796 vss SUB_GROUP_6_ N0937 vss efet w=13050 l=11600
M2797 N0937 M12 vss vss efet w=18125 l=9425
M2798 N0704 vcc vcc vss efet w=9425 l=38425
M2799 N0700 N0704 vcc vss efet w=65975 l=12325
M2800 vss M12 SUB_GROUP_6_ vss efet w=13775 l=11600
M2801 N0886 N0550 N0894 vss efet w=59450 l=11600
M2802 N0548 N0550 N0549 vss efet w=61625 l=10875
M2803 vss N0878 N0846 vss efet w=60900 l=11600
M2804 vcc vcc N0350 vss efet w=7250 l=50750
M2805 vss N0849 N0346 vss efet w=58725 l=12325
M2806 N0856 N0854 N0849 vss efet w=7975 l=12325
M2807 N0346 vcc vcc vss efet w=6525 l=32625
M2808 N0870 ACC_ADAC N0856 vss efet w=14500 l=13050
M2809 N0846 N0874 vcc vss efet w=13050 l=10150
M2810 N0894 N0870 vss vss efet w=44225 l=10875
M2811 vss CY_1 N0803 vss efet w=14500 l=17400
M2812 N0745 N0725 vss vss efet w=29000 l=13050
M2813 vcc vcc S00761 vss efet w=6525 l=11600
M2814 S00757 vcc vcc vss efet w=8700 l=13050
M2815 vss _COM N0717 vss efet w=77575 l=10875
M2816 vcc S00761 N0745 vss efet w=5800 l=27550
M2817 N0725 clk1 N0724 vss efet w=15950 l=10150
M2818 N0724 N0284 vss vss efet w=27550 l=13050
M2819 N0284 clk2 A32 vss efet w=14500 l=11600
M2820 vcc vcc N0724 vss efet w=8700 l=40600
M2821 N0288 A32 vss vss efet w=23200 l=12325
M2822 vss DAA N0802 vss efet w=13050 l=11600
M2823 N0818 N0803 vss vss efet w=28275 l=11600
M2824 N0378 DAA N0818 vss efet w=29000 l=11600
M2825 vss O_IB N0378 vss efet w=15225 l=10875
M2826 N0350 KBP vss vss efet w=17400 l=11600
M2827 N0856 vcc vcc vss efet w=10150 l=37700
M2828 N0803 N0356 N0819 vss efet w=28275 l=10150
M2829 vcc N0746 A32 vss efet w=38425 l=12325
M2830 A32 N0727 vss vss efet w=39150 l=13050
M2832 N0746 N0727 vss vss efet w=34800 l=13050
M2833 vcc vcc S00778 vss efet w=5800 l=13050
M2834 vcc S00778 N0746 vss efet w=7250 l=26100
M2835 vcc vcc N0766 vss efet w=8700 l=43500
M2836 vcc vcc N0751 vss efet w=7975 l=45675
M2837 DCL_0 vcc vcc vss efet w=7250 l=44950
M2838 vss N0348 N0819 vss efet w=34800 l=10875
M2839 N0819 N0347 vss vss efet w=37700 l=11600
M2840 N0803 vcc vcc vss efet w=5800 l=50750
M2841 N0403 vcc vcc vss efet w=6525 l=33350
M2842 N0802 vcc vcc vss efet w=6525 l=70325
M2843 N0354 vcc vcc vss efet w=7250 l=46400
M2844 N0363 vcc vcc vss efet w=9425 l=50025
M2845 N0370 vcc vcc vss efet w=7975 l=42775
M2846 vcc vcc N0345 vss efet w=7975 l=51475
M2847 N0378 vcc vcc vss efet w=7250 l=47850
M2848 N0377 N0378 N0376 vss efet w=34075 l=12325
M2849 vss N0346 ACC_0 vss efet w=21750 l=11600
M2850 CY_1 ADSL ACC_0 vss efet w=7250 l=12325
M2851 vss ACC_0 N0856 vss efet w=61625 l=11600
M2852 vss M12 N0870 vss efet w=13050 l=12325
M2853 N0471 vcc vcc vss efet w=9425 l=36975
M2854 N0346 ACB_IB D0 vss efet w=43500 l=10875
M2855 ACC_0 vcc vcc vss efet w=8700 l=44950
M2856 vss N0846 ADD_0 vss efet w=42775 l=10875
M2857 ACC_0 M12 N0471 vss efet w=7250 l=11600
M2858 N0846 ADD_ACC ACC_0 vss efet w=10150 l=11600
M2859 vss N0878 N0874 vss efet w=12325 l=13775
M2860 N0878 N0887 N0886 vss efet w=60900 l=12325
M2861 N0548 N0870 vss vss efet w=62350 l=11600
M2862 N0549 N0887 vss vss efet w=50025 l=10875
M2863 vss N0856 N0471 vss efet w=36250 l=11600
M2864 N0874 vcc vcc vss efet w=5800 l=59450
M2865 N0549 N0870 N0911 vss efet w=68875 l=17400
M2866 N0911 N0887 N0548 vss efet w=55825 l=12325
M2867 _TMP_0 N0940 vss vss efet w=22475 l=12325
M2868 vss N0705 N0700 vss efet w=95700 l=8700
M2869 _TMP_0 N0937 N0887 vss efet w=13775 l=10875
M2870 vcc N0939 _TMP_0 vss efet w=14500 l=11600
M2871 vcc vcc N0911 vss efet w=5800 l=66700
M2872 N0847 ADSR ACC_0 vss efet w=10150 l=11600
M2873 N0878 vcc vcc vss efet w=7250 l=53650
M2874 N0898 N0553 N0878 vss efet w=36250 l=13050
M2875 vss N0870 N0898 vss efet w=35525 l=13775
M2876 N0898 N0550 vss vss efet w=43500 l=13050
M2877 vss N0887 N0898 vss efet w=35525 l=12325
M2878 N0915 N0911 vss vss efet w=11600 l=11600
M2879 vcc vcc N0915 vss efet w=7250 l=63075
M2880 D0 ADD_IB N0846 vss efet w=40600 l=11600
M2881 N0870 ACC_ADA N0471 vss efet w=14500 l=13050
M2882 N0940 vcc vcc vss efet w=6525 l=45675
M2883 vss N0939 N0940 vss efet w=15225 l=12325
M2884 TMP_0 SUB_GROUP_6_ N0887 vss efet w=15225 l=12325
M2885 TMP_0 N0940 vcc vss efet w=13050 l=11600
M2886 vss N0939 TMP_0 vss efet w=23200 l=10875
M2887 vcc M12 N0604 vss efet w=7250 l=11600
M2888 N0553 N0915 vss vss efet w=20300 l=10150
M2889 D0 N0964 N0604 vss efet w=12325 l=12325
M2890 vss N0604 N0939 vss efet w=42050 l=13775
M2892 N0939 S00762 vcc vss efet w=5800 l=47850
M2893 vcc N0911 N0553 vss efet w=14500 l=11600
M2894 vss N0884 N0847 vss efet w=63075 l=13775
M2895 vcc S00764 ACC_ADAC vss efet w=5800 l=45675
M2897 ADD_0 vcc vcc vss efet w=8700 l=46400
M2898 vcc vcc N0377 vss efet w=8700 l=43500
M2899 vss DCL_0 N0751 vss efet w=35525 l=10150
M2900 N0766 N0351 vss vss efet w=22475 l=13050
M2901 vss DCL_0 N0716 vss efet w=47850 l=10150
M2902 N0751 N0766 N0767 vss efet w=12325 l=12325
M2903 DCL_0 POC vss vss efet w=23200 l=11600
M2904 vss N0350 N0376 vss efet w=37700 l=13050
M2905 vss N0767 DCL_0 vss efet w=50750 l=10150
M2906 N0345 N0350 vss vss efet w=17400 l=13050
M2907 N0354 N0350 vss vss efet w=14500 l=11600
M2908 vss N0350 N0363 vss efet w=17400 l=13050
M2909 N0370 N0350 vss vss efet w=18125 l=13775
M2910 vcc vcc N0371 vss efet w=5800 l=59450
M2911 vss N0847 ADD_0 vss efet w=39875 l=10875
M2912 N0847 ADD_IB D1 vss efet w=39875 l=11600
M2913 vcc vcc S00764 vss efet w=5800 l=11600
M2914 N0847 N0875 vcc vss efet w=15950 l=13050
M2915 vcc vcc S00767 vss efet w=9425 l=10875
M2916 D1 ACB_IB N0347 vss efet w=39875 l=11600
M2917 N0871 ACC_ADAC N0472 vss efet w=14500 l=13050
M2918 N0888 N0553 N0895 vss efet w=57275 l=10875
M2919 N0895 N0871 vss vss efet w=58000 l=11600
M2920 N0875 N0889 N0888 vss efet w=60175 l=11600
M2921 vss N0347 ACC_0 vss efet w=23200 l=10150
M2922 N0472 vcc vcc vss efet w=10875 l=35525
M2923 N0472 M12 ACC_1 vss efet w=8700 l=11600
M2924 N0472 N0857 vss vss efet w=36975 l=11600
M2925 N0846 ADSL ACC_1 vss efet w=8700 l=12325
M2926 vss N0875 N0884 vss efet w=12325 l=10875
M2927 N0551 N0553 N0552 vss efet w=60900 l=10150
M2928 N0551 N0871 vss vss efet w=65975 l=12325
M2929 N0552 N0889 vss vss efet w=48575 l=10875
M2930 N0370 N0371 vss vss efet w=17400 l=11600
M2931 N0371 N0346 vss vss efet w=14500 l=10150
M2932 vcc vcc N0364 vss efet w=6525 l=68875
M2933 N0726 N0285 vss vss efet w=27550 l=11600
M2934 N0285 clk2 A22 vss efet w=13775 l=12325
M2935 N0727 clk1 N0726 vss efet w=14500 l=11600
M2936 vcc vcc N0726 vss efet w=7975 l=37700
M2937 vss DCL_1 N0716 vss efet w=49300 l=11600
M2938 N0371 N0351 N0767 vss efet w=12325 l=10150
M2939 N0912 N0889 N0551 vss efet w=57275 l=13775
M2940 N0552 N0871 N0912 vss efet w=67425 l=15225
M2942 S00762 vcc vcc vss efet w=8700 l=11600
M2943 vss N0342 N0964 vss efet w=23925 l=13775
M2944 N0964 vcc vcc vss efet w=10875 l=35525
M2945 vss N0871 N0899 vss efet w=34800 l=14500
M2946 vss ACC_1 N0857 vss efet w=59450 l=11600
M2947 N0847 ADD_ACC ACC_1 vss efet w=8700 l=11600
M2948 N0884 vcc vcc vss efet w=10150 l=47125
M2949 N0857 vcc vcc vss efet w=10150 l=33350
M2950 N0848 ADSR ACC_1 vss efet w=7975 l=13775
M2951 N0347 vcc vcc vss efet w=7250 l=33350
M2952 vss N0850 N0347 vss efet w=58000 l=11600
M2953 N0857 N0854 N0850 vss efet w=8700 l=11600
M2954 vcc M12 N0871 vss efet w=13050 l=11600
M2955 N0875 vcc vcc vss efet w=8700 l=65250
M2956 N0899 N0556 N0875 vss efet w=35525 l=12325
M2957 N0899 N0553 vss vss efet w=43500 l=13050
M2958 vss N0889 N0899 vss efet w=36250 l=10150
M2959 N0871 ACC_ADA N0857 vss efet w=15950 l=12325
M2960 N0345 N0346 vss vss efet w=18125 l=12325
M2961 vss N0346 N0354 vss efet w=14500 l=10150
M2962 vss N0346 N0363 vss efet w=19575 l=10875
M2963 N0288 A22 vss vss efet w=23200 l=13050
M2964 vss N0765 DCL_1 vss efet w=39150 l=11600
M2965 vss N0346 N0376 vss efet w=36250 l=11600
M2966 vss N0879 N0848 vss efet w=60900 l=10150
M2967 vcc S00767 N0912 vss efet w=5800 l=51475
M2968 TMP_1 N0937 N0889 vss efet w=14500 l=11600
M2969 _TMP_1 N0942 vss vss efet w=20300 l=11600
M2970 N0672 D2 vss vss efet w=57275 l=12325
M2971 d2 POC vss vss efet w=29725 l=13775
M2972 vcc vcc N0672 vss efet w=10875 l=40600
M2973 S00765 vcc vcc vss efet w=7250 l=15950
M2974 S00766 vcc vcc vss efet w=7250 l=15225
M2976 vcc S00766 N0692 vss efet w=10150 l=12325
M2977 N0690 S00765 vcc vss efet w=12325 l=18125
M2978 vcc N0941 _TMP_1 vss efet w=13775 l=12325
M2979 N0691 N0702 N0672 vss efet w=27550 l=12325
M2980 N0942 vcc vcc vss efet w=6525 l=47125
M2981 N0916 N0912 vss vss efet w=13050 l=10150
M2982 vcc vcc N0916 vss efet w=7250 l=63075
M2983 vss N0941 N0942 vss efet w=13050 l=11600
M2985 vcc M12 N0605 vss efet w=7975 l=10150
M2986 TMP_1 N0942 vcc vss efet w=14500 l=11600
M2987 _TMP_1 SUB_GROUP_6_ N0889 vss efet w=18125 l=12325
M2988 vss N0941 TMP_1 vss efet w=20300 l=11600
M2989 N0690 N0700 vss vss efet w=262450 l=13050
M2990 D1 N0964 N0605 vss efet w=12325 l=13775
M2991 N0556 N0916 vss vss efet w=20300 l=10150
M2992 N0692 N0700 vss vss efet w=228375 l=10150
M2993 vss N0605 N0941 vss efet w=41325 l=18125
M2994 vcc N0912 N0556 vss efet w=14500 l=10150
M2996 N0941 S00781 vcc vss efet w=5800 l=43500
M2997 vss N0851 N0348 vss efet w=56550 l=11600
M2998 N0858 N0854 N0851 vss efet w=7250 l=13050
M2999 N0348 vcc vcc vss efet w=8700 l=29000
M3000 vcc N0747 A22 vss efet w=41325 l=10875
M3001 A22 N0729 vss vss efet w=37700 l=11600
M3002 vss POC DCL_1 vss efet w=23200 l=11600
M3003 DCL_1 vcc vcc vss efet w=7250 l=49300
M3004 N0364 N0351 N0765 vss efet w=12325 l=15225
M3005 vss N0364 N0363 vss efet w=17400 l=10150
M3006 vss N0347 N0345 vss efet w=24650 l=12325
M3007 N0354 N0347 vss vss efet w=13775 l=12325
M3008 N0364 N0347 vss vss efet w=14500 l=10150
M3009 N0872 ACC_ADAC N0858 vss efet w=15225 l=12325
M3010 N0848 N0876 vcc vss efet w=13775 l=15225
M3011 N0858 vcc vcc vss efet w=10150 l=41325
M3012 vss N0347 N0370 vss efet w=18850 l=10150
M3013 vss N0347 N0376 vss efet w=36250 l=10150
M3014 vss DCL_1 N0750 vss efet w=23200 l=11600
M3015 N0750 vcc vcc vss efet w=7250 l=52200
M3017 N0747 N0729 vss vss efet w=32625 l=15225
M3018 vcc vcc S00800 vss efet w=6525 l=13775
M3019 vcc S00800 N0747 vss efet w=5800 l=24650
M3020 N0750 N0766 N0765 vss efet w=10150 l=11600
M3021 vcc vcc N0355 vss efet w=6525 l=73225
M3022 N0355 N0351 N0768 vss efet w=10150 l=10150
M3023 N0354 N0355 vss vss efet w=13050 l=11600
M3024 N0355 N0348 vss vss efet w=15225 l=10875
M3025 vss N0348 ACC_0 vss efet w=23200 l=11600
M3026 N0847 ADSL ACC_2 vss efet w=7250 l=14500
M3027 vss ACC_2 N0858 vss efet w=64525 l=11600
M3028 N0473 vcc vcc vss efet w=12325 l=36975
M3029 vss N0848 ADD_0 vss efet w=42775 l=10875
M3030 N0348 ACB_IB D2 vss efet w=39150 l=13775
M3031 N0848 ADD_ACC ACC_2 vss efet w=7975 l=11600
M3032 ACC_2 M12 N0473 vss efet w=7975 l=12325
M3033 vss N0858 N0473 vss efet w=36250 l=11600
M3034 N0890 N0556 N0896 vss efet w=59450 l=11600
M3035 N0896 N0872 vss vss efet w=60900 l=10150
M3036 N0879 N0891 N0890 vss efet w=65250 l=10875
M3037 N0554 N0872 vss vss efet w=64525 l=10875
M3038 vss N0879 N0876 vss efet w=10150 l=12325
M3039 vss M12 N0872 vss efet w=15225 l=10875
M3040 N0514 ADSR ACC_2 vss efet w=9425 l=12325
M3041 N0555 N0891 vss vss efet w=52925 l=10875
M3042 N0555 N0872 N0913 vss efet w=68150 l=14500
M3043 N0913 N0891 N0554 vss efet w=56550 l=11600
M3044 N0876 vcc vcc vss efet w=8700 l=65975
M3045 D2 ADD_IB N0848 vss efet w=42775 l=11600
M3046 N0872 ACC_ADA N0473 vss efet w=14500 l=11600
M3047 N0879 vcc vcc vss efet w=9425 l=57275
M3048 vss DCL_2 N0716 vss efet w=43500 l=10150
M3049 N0728 N0286 vss vss efet w=27550 l=11600
M3050 N0729 clk1 N0728 vss efet w=13775 l=12325
M3051 N0286 clk2 A12 vss efet w=15950 l=11600
M3052 vss N0768 DCL_2 vss efet w=42050 l=10150
M3053 vss N0348 N0345 vss efet w=18850 l=11600
M3054 vss N0348 N0363 vss efet w=20300 l=11600
M3055 vss N0348 N0370 vss efet w=19575 l=10875
M3056 vss N0348 N0376 vss efet w=36250 l=10150
M3057 N0900 N0559 N0879 vss efet w=34800 l=12325
M3058 vss N0872 N0900 vss efet w=36250 l=10150
M3059 N0900 N0556 vss vss efet w=43500 l=11600
M3060 vss N0891 N0900 vss efet w=40600 l=13050
M3062 N0554 N0556 N0555 vss efet w=60900 l=11600
M3063 vss N0691 N0690 vss efet w=97875 l=9425
M3064 D2 N0964 N0606 vss efet w=19575 l=17400
M3065 vss N0690 N0692 vss efet w=73950 l=11600
M3066 S00781 vcc vcc vss efet w=9425 l=12325
M3067 vcc vcc N0913 vss efet w=5800 l=58000
M3068 _TMP_2 N0944 vss vss efet w=22475 l=11600
M3069 _TMP_2 N0937 N0891 vss efet w=15950 l=10875
M3070 vcc N0943 _TMP_2 vss efet w=14500 l=13050
M3071 vss N0692 d2 vss efet w=1202775 l=7250
M3072 N0606 M12 vcc vss efet w=8700 l=11600
M3073 N0665 N0676 vss vss efet w=26100 l=13050
M3074 N0917 N0913 vss vss efet w=13050 l=10875
M3075 vcc vcc N0917 vss efet w=5800 l=63800
M3076 N0559 N0917 vss vss efet w=20300 l=11600
M3077 vcc N0913 N0559 vss efet w=15225 l=10875
M3078 vcc vcc S00804 vss efet w=5800 l=11600
M3079 N0944 vcc vcc vss efet w=7975 l=44225
M3080 vss N0943 N0944 vss efet w=13775 l=15225
M3081 TMP_2 N0944 vcc vss efet w=15950 l=13775
M3082 vss N0943 TMP_2 vss efet w=19575 l=13775
M3083 TMP_2 SUB_GROUP_6_ N0891 vss efet w=15225 l=12325
M3084 d2 N0690 vcc vss efet w=640175 l=13775
M3085 vcc vcc N0665 vss efet w=11600 l=52200
M3086 N0665 N0666 vss vss efet w=14500 l=13050
M3087 N0943 S00801 vcc vss efet w=8700 l=53650
M3088 vcc vcc N0349 vss efet w=6525 l=61625
M3089 vcc S00803 ACC_ADA vss efet w=6525 l=45675
M3090 vcc vcc N0728 vss efet w=7250 l=38425
M3091 N0288 A12 vss vss efet w=22475 l=11600
M3092 DCL_2 vcc vcc vss efet w=8700 l=43500
M3093 N0749 vcc vcc vss efet w=7250 l=43500
M3094 vcc N0748 A12 vss efet w=39150 l=13050
M3095 vss POC DCL_2 vss efet w=26100 l=10875
M3096 vss DCL_2 N0749 vss efet w=23200 l=11600
M3097 A12 N0731 vss vss efet w=38425 l=12325
M3099 N0748 N0731 vss vss efet w=27550 l=11600
M3100 vcc vcc S00814 vss efet w=5800 l=12325
M3101 N0768 N0766 N0749 vss efet w=9425 l=13775
M3102 vss N0349 N0345 vss efet w=19575 l=13050
M3103 N0354 N0356 vss vss efet w=15225 l=10875
M3104 N0349 N0356 vss vss efet w=11600 l=10150
M3105 vss N0514 ADD_0 vss efet w=41325 l=10875
M3106 vss N0356 N0363 vss efet w=17400 l=10150
M3107 vss N0356 N0370 vss efet w=19575 l=15225
M3108 vss N0356 N0376 vss efet w=33350 l=10150
M3109 vcc S00814 N0748 vss efet w=5800 l=26100
M3110 N0514 ADD_IB D3 vss efet w=40600 l=11600
M3111 vcc vcc S00803 vss efet w=5800 l=10150
M3112 N0514 N0877 vcc vss efet w=19575 l=12325
M3113 D3 ACB_IB N0356 vss efet w=40600 l=11600
M3114 N0873 ACC_ADAC N0474 vss efet w=15950 l=13775
M3115 vss N0377 N0358 vss efet w=64525 l=13775
M3116 vss N0345 N0358 vss efet w=72500 l=11600
M3117 N0358 N0354 vss vss efet w=66700 l=11600
M3118 vss N0363 N0358 vss efet w=74675 l=12325
M3119 N0358 N0370 vss vss efet w=60175 l=10875
M3120 N0358 vcc vcc vss efet w=6525 l=65975
M3122 N0714 N0749 vss vss efet w=45675 l=12325
M3123 N0731 clk1 N0730 vss efet w=13775 l=10150
M3124 N0730 N0287 vss vss efet w=29000 l=12325
M3125 vcc vcc N0730 vss efet w=7975 l=39150
M3126 N0287 clk2 N0288 vss efet w=13050 l=11600
M3127 vss _COM N0714 vss efet w=45675 l=10875
M3128 vcc vcc S00818 vss efet w=7975 l=12325
M3129 vcc S00818 N0714 vss efet w=10150 l=24650
M3130 N0366 vcc vcc vss efet w=5800 l=66700
M3131 vcc vcc N0288 vss efet w=8700 l=34800
M3133 N0715 N0750 vss vss efet w=44950 l=11600
M3134 vcc N0714 cm_ram3 vss efet w=142100 l=11600
M3135 N0734 N0714 vss vss efet w=47850 l=18850
M3136 vss _COM N0715 vss efet w=43500 l=10150
M3137 N0366 N0354 vss vss efet w=61625 l=10875
M3138 vss N0363 N0366 vss efet w=59450 l=11600
M3139 N0366 N0370 vss vss efet w=60900 l=10875
M3140 vss N0377 N0366 vss efet w=59450 l=11600
M3141 vss N0403 N0358 vss efet w=60900 l=10150
M3142 vss N0356 ACC_0 vss efet w=23200 l=11600
M3143 N0474 vcc vcc vss efet w=10875 l=35525
M3144 N0356 N0852 vss vss efet w=53650 l=13050
M3145 N0356 vcc vcc vss efet w=8700 l=34800
M3146 N0366 TCS vss vss efet w=60175 l=10875
M3147 vcc vcc S00825 vss efet w=7975 l=12325
M3148 vcc N0715 cm_ram2 vss efet w=141375 l=12325
M3149 vcc vcc N0734 vss efet w=8700 l=20300
M3150 vcc vcc N0735 vss efet w=9425 l=19575
M3151 vss N0715 N0735 vss efet w=40600 l=13050
M3152 vcc S00825 N0715 vss efet w=10150 l=24650
M3153 N0359 vcc vcc vss efet w=6525 l=61625
M3154 vss N0345 N0359 vss efet w=61625 l=10875
M3155 N0357 vcc vcc vss efet w=6525 l=68150
M3157 cm_ram2 N0735 vss vss efet w=263900 l=14500
M3158 cm_ram3 N0734 vss vss efet w=263900 l=11600
M3159 vss _COM N0713 vss efet w=43500 l=13050
M3160 N0716 _COM vss vss efet w=59450 l=11600
M3162 S00834 vcc vcc vss efet w=7975 l=12325
M3163 N0713 N0751 vss vss efet w=47125 l=10875
M3164 N0359 N0370 vss vss efet w=65975 l=12325
M3165 vss N0377 N0359 vss efet w=60175 l=12325
M3166 D2 N0415 N0366 vss efet w=49300 l=11600
M3167 D3 N0415 N0358 vss efet w=49300 l=14500
M3168 N0359 TCS vss vss efet w=59450 l=11600
M3169 vcc vcc S00833 vss efet w=7975 l=12325
M3170 vcc S00833 N0716 vss efet w=10875 l=23925
M3171 N0713 S00834 vcc vss efet w=9425 l=22475
M3172 vss N0345 N0357 vss efet w=62350 l=13775
M3173 vss N0363 N0357 vss efet w=63800 l=15950
M3174 vss N0377 N0357 vss efet w=60175 l=12325
M3175 D1 N0415 N0359 vss efet w=50750 l=11600
M3176 D0 N0415 N0357 vss efet w=55825 l=11600
M3177 N0474 M12 ACC_3 vss efet w=8700 l=11600
M3178 N0474 N0859 vss vss efet w=36250 l=11600
M3179 N0848 ADSL ACC_3 vss efet w=8700 l=11600
M3180 vss N0885 N0514 vss efet w=65975 l=10875
M3181 vss N0606 N0943 vss efet w=41325 l=13775
M3182 N0897 N0873 vss vss efet w=60175 l=10875
M3183 vss N0877 N0885 vss efet w=13775 l=10150
M3184 N0892 N0559 N0897 vss efet w=56550 l=11600
M3185 N0877 N0893 N0892 vss efet w=65250 l=10150
M3186 N0557 N0873 vss vss efet w=76125 l=19575
M3187 vss N0893 N0558 vss efet w=61625 l=28275
M3188 vss ACC_3 N0859 vss efet w=58725 l=13775
M3189 N0514 ADD_ACC ACC_3 vss efet w=9425 l=10875
M3190 N0859 vcc vcc vss efet w=9425 l=35525
M3191 N0514 ADSL N0513 vss efet w=15225 l=12325
M3192 N0859 N0854 N0852 vss efet w=7250 l=13050
M3193 N0513 ADSR ACC_3 vss efet w=13050 l=13775
M3194 N0914 N0893 N0557 vss efet w=55825 l=12325
M3195 vss N0873 N0901 vss efet w=35525 l=12325
M3196 N0885 vcc vcc vss efet w=9425 l=54375
M3197 vcc M12 N0873 vss efet w=13775 l=12325
M3198 N0901 N0861 N0877 vss efet w=37700 l=10150
M3199 N0877 vcc vcc vss efet w=7975 l=64525
M3200 N0873 ACC_ADA N0859 vss efet w=15950 l=10875
M3201 N0558 N0873 N0914 vss efet w=65975 l=16675
M3202 N0901 N0559 vss vss efet w=43500 l=10150
M3203 vss N0893 N0901 vss efet w=37700 l=11600
M3204 N0557 N0559 N0558 vss efet w=58000 l=10150
M3207 S00801 vcc vcc vss efet w=12325 l=13050
M3208 D2 N0666 vss vss efet w=49300 l=13775
M3209 vcc N0665 D2 vss efet w=39875 l=15225
M3210 vcc S00804 N0914 vss efet w=5075 l=52200
M3211 vcc vcc N0666 vss efet w=10150 l=39150
M3212 _TMP_3 N0946 vss vss efet w=21025 l=13050
M3213 N0666 d2 vss vss efet w=71050 l=12325
M3214 _TMP_3 SUB_GROUP_6_ N0893 vss efet w=14500 l=11600
M3215 N0666 N0676 vss vss efet w=44950 l=12325
M3216 vcc N0945 _TMP_3 vss efet w=13775 l=12325
M3217 N0918 N0914 vss vss efet w=12325 l=12325
M3218 vcc vcc N0918 vss efet w=5800 l=63800
M3219 N0861 N0918 vss vss efet w=18850 l=11600
M3220 N0946 vcc vcc vss efet w=8700 l=43500
M3221 vss N0945 N0946 vss efet w=13050 l=11600
M3222 vcc M12 N0607 vss efet w=9425 l=8700
M3223 TMP_3 N0937 N0893 vss efet w=15225 l=12325
M3224 TMP_3 N0946 vcc vss efet w=13775 l=12325
M3225 vcc N0914 N0861 vss efet w=13050 l=11600
M3226 vcc vcc S00817 vss efet w=6525 l=9425
M3227 vss N0945 TMP_3 vss efet w=20300 l=11600
M3228 D3 N0964 N0607 vss efet w=14500 l=14500
M3230 vss N0607 N0945 vss efet w=38425 l=13775
M3231 d0 vss vss vss efet w=116000 l=13050
M3233 vss N0403 N0357 vss efet w=60175 l=13775
M3234 vcc vcc S00819 vss efet w=7250 l=9425
M3235 N0945 S00817 vcc vss efet w=5800 l=40600
M3237 N0670 d0 vss vss efet w=71775 l=12325
M3238 vss N0670 D0 vss efet w=49300 l=11600
M3239 vss N0670 N0669 vss efet w=13775 l=11600
M3240 d1 vss vss vss efet w=114550 l=14500
M3241 N0854 S00828 vcc vss efet w=7250 l=52200
M3242 vcc vcc S00828 vss efet w=8700 l=13050
M3243 N0670 N0676 vss vss efet w=51475 l=13775
M3244 vss N0676 N0669 vss efet w=25375 l=11600
M3245 D0 N0669 vcc vss efet w=38425 l=13050
M3246 N0670 vcc vcc vss efet w=10150 l=36975
M3247 N0669 vcc vcc vss efet w=5800 l=50750
M3248 vss D0 N0674 vss efet w=57275 l=12325
M3249 N0674 vcc vcc vss efet w=13050 l=39150
M3250 N0674 N0702 N0697 vss efet w=27550 l=11600
M3251 vss N0697 N0696 vss efet w=99325 l=10875
M3252 d0 N0696 vcc vss efet w=666275 l=10875
M3253 N0733 N0713 vss vss efet w=55100 l=14500
M3254 vcc N0713 cm_ram1 vss efet w=142100 l=11600
M3255 vcc N0716 cm_ram0 vss efet w=142100 l=11600
M3256 vcc vcc N0733 vss efet w=7250 l=23200
M3257 vcc vcc N0736 vss efet w=8700 l=21750
M3258 vss N0716 N0736 vss efet w=43500 l=11600
M3259 cm_ram1 N0733 vss vss efet w=261725 l=12325
M3260 cm_ram0 N0736 vss vss efet w=256650 l=11600
M3261 vss N0698 d0 vss efet w=1218725 l=6525
M3262 N0696 N0700 vss vss efet w=247950 l=11600
M3263 vcc vcc S00835 vss efet w=9425 l=12325
M3264 vcc S00835 N0696 vss efet w=10875 l=13775
M3266 vss N0696 N0698 vss efet w=81925 l=12325
M3267 N0698 N0700 vss vss efet w=229100 l=11600
M3268 vcc S00839 N0698 vss efet w=10150 l=11600
M3270 vcc vcc S00839 vss efet w=10150 l=13050
M3271 N0668 d1 vss vss efet w=66700 l=13050
M3272 N0937 S00819 vcc vss efet w=6525 l=33350
M3273 vss vss d2 vss efet w=99325 l=15225
M3274 vss N0668 D1 vss efet w=49300 l=11600
M3275 N0667 N0668 vss vss efet w=16675 l=10875
M3276 vss N0676 N0667 vss efet w=26825 l=12325
M3277 N0668 N0676 vss vss efet w=44225 l=13775
M3278 vcc vcc N0667 vss efet w=6525 l=55825
M3279 D1 N0667 vcc vss efet w=39150 l=11600
M3280 N0668 vcc vcc vss efet w=8700 l=35525
M3281 vss D1 N0673 vss efet w=50750 l=10875
M3282 N0673 N0702 N0694 vss efet w=27550 l=12325
M3283 N0673 vcc vcc vss efet w=10875 l=36975
M3284 D3 N0664 vss vss efet w=49300 l=12325
M3285 vcc N0663 D3 vss efet w=39875 l=12325
M3286 vss POC d3 vss efet w=29000 l=14500
M3287 vcc N0693 d1 vss efet w=681500 l=11600
M3288 d0 POC vss vss efet w=33350 l=11600
M3289 vss N0694 N0693 vss efet w=99325 l=10875
M3290 N0693 N0700 vss vss efet w=257375 l=19575
M3291 vcc vcc S00836 vss efet w=7250 l=11600
M3292 vcc S00836 N0693 vss efet w=9425 l=13775
M3293 vss N0695 d1 vss efet w=1217275 l=6525
M3295 vcc vcc N0663 vss efet w=9425 l=49300
M3296 vcc vcc N0664 vss efet w=8700 l=36250
M3297 vss N0676 N0664 vss efet w=56550 l=14500
M3298 vss N0693 N0695 vss efet w=75400 l=13050
M3299 N0695 N0700 vss vss efet w=229825 l=10875
M3300 vcc S00840 N0695 vss efet w=10150 l=14500
M3302 vcc vcc S00840 vss efet w=7250 l=13775
M3303 vss N0664 N0663 vss efet w=23200 l=15950
M3304 N0663 N0676 vss vss efet w=23925 l=11600
M3305 vss d3 N0664 vss efet w=86275 l=15225
M3306 d3 vss vss vss efet w=124700 l=13050
M3307 d1 POC vss vss efet w=30450 l=10875
