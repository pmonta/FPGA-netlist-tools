* SPICE3 converted from Lajos's format

M0 VDD VDD N0037 GND efet
M1 VDD VDD N0040 GND efet
M2 GND N0031 N0037 GND efet
M3 GND N0038 N0040 GND efet
M4 VDD VDD N0038 GND efet
M5 N0038 N0037 GND GND efet
M6 N0031 N0032 GND GND efet
M7 N0031 N0029 GND GND efet
M8 GND N0031 N0032 GND efet
M9 GND GND DATA GND efet
M10 GND N0137 Q4 GND efet
M11 GND N0119 Q3 GND efet
M12 GND N0099 Q2 GND efet
M13 GND N0079 Q1 GND efet
M14 GND N0059 Q0 GND efet
M15 N0032 N0027 GND GND efet
M16 N0127 N0128 GND GND efet
M17 N0109 N0110 GND GND efet
M18 N0089 N0090 GND GND efet
M19 N0069 N0070 GND GND efet
M20 N0049 N0050 GND GND efet
M21 VDD VDD N0031 GND efet
M22 VDD VDD N0032 GND efet
M23 GND N0027 N0029 GND efet
M24 N0127 N0021 GND GND efet
M25 N0109 N0021 GND GND efet
M26 N0089 N0021 GND GND efet
M27 N0069 N0021 GND GND efet
M28 N0049 N0021 GND GND efet
M29 VDD VDD N0029 GND efet
M30 N0027 N0024 GND GND efet
M31 GND GND CLOCK GND efet
M32 N0059 N0049 GND GND efet
M33 N0137 N0127 GND GND efet
M34 N0119 N0109 GND GND efet
M35 N0099 N0089 GND GND efet
M36 N0079 N0069 GND GND efet
M37 N0024 N0022 GND GND efet
M38 VDD VDD N0027 GND efet
M39 VDD VDD N0127 GND efet
M40 VDD VDD N0109 GND efet
M41 VDD VDD N0089 GND efet
M42 VDD VDD N0069 GND efet
M43 VDD VDD N0049 GND efet
M44 VDD VDD N0119 GND efet
M45 VDD VDD N0099 GND efet
M46 VDD VDD N0079 GND efet
M47 VDD VDD N0059 GND efet
M48 VDD VDD N0137 GND efet
M49 VDD N0049 Q0 GND efet
M50 VDD N0127 Q4 GND efet
M51 VDD N0109 Q3 GND efet
M52 VDD N0089 Q2 GND efet
M53 VDD N0069 Q1 GND efet
M54 VDD VDD N0024 GND efet
M55 VDD VDD N0019 GND efet
M56 VDD VDD N0121 GND efet
M57 VDD VDD N0101 GND efet
M58 VDD VDD N0081 GND efet
M59 VDD VDD N0061 GND efet
M60 VDD VDD N0041 GND efet
M61 N0121 N0040 N0128 GND efet
M62 N0101 N0040 N0110 GND efet
M63 N0081 N0040 N0090 GND efet
M64 N0061 N0040 N0070 GND efet
M65 N0041 N0040 N0050 GND efet
M66 N0107 N0032 N0123 GND efet
M67 N0087 N0032 N0103 GND efet
M68 N0067 N0032 N0083 GND efet
M69 N0047 N0032 N0063 GND efet
M70 GND N0019 N0022 GND efet
M71 N0131 N0040 N0121 GND efet
M72 N0113 N0040 N0101 GND efet
M73 N0093 N0040 N0081 GND efet
M74 N0073 N0040 N0061 GND efet
M75 N0053 N0040 N0041 GND efet
M76 N0042 N0031 N0041 GND efet
M77 N0122 N0031 N0121 GND efet
M78 N0102 N0031 N0101 GND efet
M79 N0082 N0031 N0081 GND efet
M80 N0062 N0031 N0061 GND efet
M81 GND CLOCK N0019 GND efet
M82 N0101 N0032 N0134 GND efet
M83 N0081 N0032 N0116 GND efet
M84 N0061 N0032 N0096 GND efet
M85 N0041 N0032 N0076 GND efet
M86 GND N0123 N0122 GND efet
M87 GND N0103 N0102 GND efet
M88 GND N0083 N0082 GND efet
M89 GND N0063 N0062 GND efet
M90 GND N0047 N0041 GND efet
M91 GND N0043 N0042 GND efet
M92 GND N0126 N0121 GND efet
M93 GND N0107 N0101 GND efet
M94 GND N0087 N0081 GND efet
M95 GND N0067 N0061 GND efet
M96 N0020 DATA GND GND efet
M97 VDD VDD N0023 GND efet
M98 N0055 N0056 GND GND efet
M99 N0133 N0134 GND GND efet
M100 N0115 N0116 GND GND efet
M101 N0095 N0096 GND GND efet
M102 N0075 N0076 GND GND efet
M103 N0047 N0053 GND GND efet
M104 N0126 N0131 GND GND efet
M105 N0107 N0113 GND GND efet
M106 N0087 N0093 GND GND efet
M107 N0067 N0073 GND GND efet
M108 GND N0020 N0023 GND efet
M109 N0087 N0031 N0095 GND efet
M110 N0067 N0031 N0075 GND efet
M111 N0047 N0031 N0055 GND efet
M112 N0126 N0031 N0133 GND efet
M113 N0107 N0031 N0115 GND efet
M114 N0023 N0032 N0043 GND efet
M115 N0126 N0039 GND GND efet
M116 GND N0039 N0107 GND efet
M117 GND N0039 N0087 GND efet
M118 GND N0039 N0067 GND efet
M119 GND N0039 N0047 GND efet
M120 VDD VDD N0126 GND efet
M121 VDD VDD N0107 GND efet
M122 VDD VDD N0087 GND efet
M123 VDD VDD N0067 GND efet
M124 VDD VDD N0047 GND efet
M125 N0020 N0032 N0056 GND efet
M126 VDD VDD N0022 GND efet
M127 VDD VDD N0020 GND efet
M128 VDD VDD N0048 GND efet
M129 VDD VDD N0068 GND efet
M130 VDD VDD N0088 GND efet
M131 VDD VDD N0108 GND efet
M132 VDD VDD N0036 GND efet
M133 VDD VDD N0039 GND efet
M134 GND N0034 N0039 GND efet
M135 VDD VDD N0030 GND efet
M136 N0058 N0032 N0121 GND efet
M137 N0046 N0032 N0126 GND efet
M138 VDD VDD N0034 GND efet
M139 N0034 N0030 GND GND efet
M140 GND N0027 N0030 GND efet
M141 N0048 N0039 GND GND efet
M142 N0068 N0039 GND GND efet
M143 N0088 N0039 GND GND efet
M144 N0108 N0039 GND GND efet
M145 N0036 N0039 GND GND efet
M146 VDD VDD N0035 GND efet
M147 N0097 N0031 N0088 GND efet
M148 N0117 N0031 N0108 GND efet
M149 N0135 N0031 N0036 GND efet
M150 N0033 N0034 N0030 GND efet
M151 N0057 N0031 N0048 GND efet
M152 N0077 N0031 N0068 GND efet
M153 GND N0132 N0036 GND efet
M154 GND N0058 N0057 GND efet
M155 GND N0035 N0033 GND efet
M156 GND N0054 N0048 GND efet
M157 GND N0078 N0077 GND efet
M158 GND N0074 N0068 GND efet
M159 GND N0098 N0097 GND efet
M160 GND N0094 N0088 GND efet
M161 GND N0118 N0117 GND efet
M162 GND N0114 N0108 GND efet
M163 GND N0136 N0135 GND efet
M164 N0028 N0017 GND GND efet
M165 N0085 N0086 GND GND efet
M166 N0105 N0106 GND GND efet
M167 N0124 N0125 GND GND efet
M168 N0045 N0046 GND GND efet
M169 N0065 N0066 GND GND efet
M170 N0044 N0048 GND GND efet
M171 N0064 N0068 GND GND efet
M172 N0084 N0088 GND GND efet
M173 N0104 N0108 GND GND efet
M174 N0026 N0036 GND GND efet
M175 N0025 N0032 GND GND efet
M176 N0017 N0028 GND GND efet
M177 N0078 N0032 N0044 GND efet
M178 N0098 N0032 N0064 GND efet
M179 N0118 N0032 N0084 GND efet
M180 N0136 N0032 N0104 GND efet
M181 N0044 N0031 N0045 GND efet
M182 N0064 N0031 N0065 GND efet
M183 N0084 N0031 N0085 GND efet
M184 N0104 N0031 N0105 GND efet
M185 N0026 N0031 N0124 GND efet
M186 N0028 N0036 N0025 GND efet
M187 N0017 N0026 N0025 GND efet
M188 N0044 N0040 N0054 GND efet
M189 N0064 N0040 N0074 GND efet
M190 N0084 N0040 N0094 GND efet
M191 N0104 N0040 N0114 GND efet
M192 N0026 N0040 N0132 GND efet
M193 N0066 N0032 N0048 GND efet
M194 N0086 N0032 N0068 GND efet
M195 N0106 N0032 N0088 GND efet
M196 N0125 N0032 N0108 GND efet
M197 VDD VDD N0028 GND efet
M198 VDD VDD N0026 GND efet
M199 VDD VDD N0044 GND efet
M200 VDD VDD N0064 GND efet
M201 VDD VDD N0084 GND efet
M202 VDD VDD N0104 GND efet
M203 VDD VDD N0017 GND efet
M204 N0130 N0040 N0026 GND efet
M205 N0052 N0040 N0044 GND efet
M206 N0072 N0040 N0064 GND efet
M207 N0092 N0040 N0084 GND efet
M208 N0112 N0040 N0104 GND efet
M209 VDD VDD N0021 GND efet
M210 VDD VDD N0100 GND efet
M211 VDD VDD N0120 GND efet
M212 VDD VDD N0138 GND efet
M213 OUT N0017 VDD GND efet
M214 VDD VDD N0060 GND efet
M215 VDD VDD N0080 GND efet
M216 VDD VDD N0091 GND efet
M217 VDD VDD N0111 GND efet
M218 VDD VDD N0129 GND efet
M219 VDD VDD N0051 GND efet
M220 VDD VDD N0071 GND efet
M221 Q5 N0051 VDD GND efet
M222 Q6 N0071 VDD GND efet
M223 Q7 N0091 VDD GND efet
M224 Q8 N0111 VDD GND efet
M225 Q9 N0129 VDD GND efet
M226 GND N0051 N0060 GND efet
M227 GND N0071 N0080 GND efet
M228 GND N0091 N0100 GND efet
M229 GND N0111 N0120 GND efet
M230 GND N0129 N0138 GND efet
M231 GND EN N0021 GND efet
M232 VDD VDD N0018 GND efet
M233 GND N0018 OUT GND efet
M234 Q5 N0060 GND GND efet
M235 GND N0021 N0051 GND efet
M236 GND N0052 N0051 GND efet
M237 Q6 N0080 GND GND efet
M238 GND N0021 N0071 GND efet
M239 GND N0072 N0071 GND efet
M240 Q7 N0100 GND GND efet
M241 GND N0021 N0091 GND efet
M242 GND N0092 N0091 GND efet
M243 Q8 N0120 GND GND efet
M244 Q9 N0138 GND GND efet
M245 GND N0021 N0129 GND efet
M246 GND N0130 N0129 GND efet
M247 GND N0021 N0111 GND efet
M248 GND N0112 N0111 GND efet
M249 GND N0017 N0018 GND efet
M250 GND GND EN GND efet
