* SPICE3 file created from 4002.ext - technology: nmos

.option scale=1u

M1000 d1 GND GND GND efet w=262 l=19
+ ad=113738 pd=7580 as=2.46415e+06 ps=180164 
M1001 diff_724_7211# diff_898_7246# GND GND efet w=191 l=16
+ ad=18994 pd=1464 as=0 ps=0 
M1002 GND diff_220_5722# diff_724_7211# GND efet w=536 l=16
+ ad=0 pd=0 as=0 ps=0 
M1003 GND d1 diff_244_7114# GND efet w=137 l=14
+ ad=0 pd=0 as=8042 ps=726 
M1004 GND diff_220_5722# diff_898_7246# GND efet w=556 l=14
+ ad=0 pd=0 as=24919 ps=1906 
M1005 diff_898_7246# diff_1144_7198# GND GND efet w=527 l=17
+ ad=0 pd=0 as=0 ps=0 
M1006 diff_724_7211# diff_724_7144# diff_724_7211# GND efet w=98 l=32
+ ad=0 pd=0 as=0 ps=0 
M1007 GND diff_244_7114# diff_413_7055# GND efet w=53 l=17
+ ad=0 pd=0 as=8711 ps=684 
M1008 diff_244_7114# diff_244_7114# diff_244_7114# GND efet w=5 l=9
+ ad=0 pd=0 as=0 ps=0 
M1009 diff_244_7114# diff_244_7114# diff_244_7114# GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M1010 diff_413_7055# diff_413_7055# diff_413_7055# GND efet w=7 l=7
+ ad=0 pd=0 as=0 ps=0 
M1011 diff_413_7055# diff_413_7055# diff_413_7055# GND efet w=2 l=9
+ ad=0 pd=0 as=0 ps=0 
M1012 diff_244_7114# Vdd Vdd GND efet w=22 l=86
+ ad=0 pd=0 as=1.05552e+06 ps=86918 
M1013 GND diff_331_7000# diff_244_7114# GND efet w=85 l=16
+ ad=0 pd=0 as=0 ps=0 
M1014 diff_413_7055# diff_331_7000# GND GND efet w=89 l=16
+ ad=0 pd=0 as=0 ps=0 
M1015 GND diff_724_7211# d1 GND efet w=2810 l=9
+ ad=0 pd=0 as=0 ps=0 
M1016 diff_898_7246# diff_967_7144# diff_898_7246# GND efet w=104 l=32
+ ad=0 pd=0 as=0 ps=0 
M1017 diff_724_7211# diff_724_7144# Vdd GND efet w=26 l=20
+ ad=0 pd=0 as=0 ps=0 
M1018 diff_724_7144# diff_724_7144# diff_724_7144# GND efet w=5 l=8
+ ad=1333 pd=184 as=0 ps=0 
M1019 diff_724_7144# diff_724_7144# diff_724_7144# GND efet w=3 l=16
+ ad=0 pd=0 as=0 ps=0 
M1020 diff_898_7246# diff_967_7144# Vdd GND efet w=26 l=20
+ ad=0 pd=0 as=0 ps=0 
M1021 diff_967_7144# diff_967_7144# diff_967_7144# GND efet w=5 l=8
+ ad=1279 pd=172 as=0 ps=0 
M1022 diff_967_7144# diff_967_7144# diff_967_7144# GND efet w=3 l=16
+ ad=0 pd=0 as=0 ps=0 
M1023 diff_724_7144# Vdd Vdd GND efet w=22 l=16
+ ad=0 pd=0 as=0 ps=0 
M1024 Vdd Vdd Vdd GND efet w=5 l=9
+ ad=0 pd=0 as=0 ps=0 
M1025 Vdd Vdd Vdd GND efet w=1 l=1
+ ad=0 pd=0 as=0 ps=0 
M1026 Vdd Vdd diff_413_7055# GND efet w=19 l=92
+ ad=0 pd=0 as=0 ps=0 
M1027 diff_629_6919# diff_413_7055# Vdd GND efet w=94 l=22
+ ad=76062 pd=6984 as=0 ps=0 
M1028 GND diff_244_7114# diff_629_6919# GND efet w=94 l=16
+ ad=0 pd=0 as=0 ps=0 
M1029 d0 GND GND GND efet w=268 l=19
+ ad=110681 pd=7622 as=0 ps=0 
M1030 GND diff_220_5722# diff_3157_7220# GND efet w=526 l=16
+ ad=0 pd=0 as=18904 ps=1446 
M1031 GND d0 diff_2359_7109# GND efet w=136 l=16
+ ad=0 pd=0 as=7791 ps=718 
M1032 diff_3157_7220# diff_3328_7249# GND GND efet w=187 l=16
+ ad=0 pd=0 as=0 ps=0 
M1033 GND diff_220_5722# diff_3328_7249# GND efet w=542 l=17
+ ad=0 pd=0 as=24580 ps=1798 
M1034 diff_3328_7249# diff_3574_7198# GND GND efet w=529 l=16
+ ad=0 pd=0 as=0 ps=0 
M1035 GND diff_2359_7109# diff_2522_7033# GND efet w=52 l=16
+ ad=0 pd=0 as=8828 ps=716 
M1036 diff_2359_7109# diff_2359_7109# diff_2359_7109# GND efet w=5 l=12
+ ad=0 pd=0 as=0 ps=0 
M1037 diff_2522_7033# diff_2522_7033# diff_2522_7033# GND efet w=12 l=11
+ ad=0 pd=0 as=0 ps=0 
M1038 d1 diff_898_7246# Vdd GND efet w=1513 l=16
+ ad=0 pd=0 as=0 ps=0 
M1039 diff_1144_7198# diff_1144_7198# diff_1144_7198# GND efet w=5 l=21
+ ad=5932 pd=554 as=0 ps=0 
M1040 diff_967_7144# Vdd Vdd GND efet w=19 l=19
+ ad=0 pd=0 as=0 ps=0 
M1041 diff_1144_7198# diff_1144_7198# diff_1144_7198# GND efet w=5 l=10
+ ad=0 pd=0 as=0 ps=0 
M1042 diff_2522_7033# diff_2522_7033# diff_2522_7033# GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M1043 diff_2359_7109# Vdd Vdd GND efet w=20 l=86
+ ad=0 pd=0 as=0 ps=0 
M1044 GND diff_331_7000# diff_2359_7109# GND efet w=85 l=16
+ ad=0 pd=0 as=0 ps=0 
M1045 diff_2522_7033# diff_331_7000# GND GND efet w=85 l=16
+ ad=0 pd=0 as=0 ps=0 
M1046 diff_3157_7220# diff_3154_7144# diff_3157_7220# GND efet w=89 l=77
+ ad=0 pd=0 as=0 ps=0 
M1047 GND diff_3157_7220# d0 GND efet w=2789 l=9
+ ad=0 pd=0 as=0 ps=0 
M1048 diff_3328_7249# diff_3397_7141# diff_3328_7249# GND efet w=83 l=82
+ ad=0 pd=0 as=0 ps=0 
M1049 diff_3157_7220# diff_3154_7144# Vdd GND efet w=23 l=17
+ ad=0 pd=0 as=0 ps=0 
M1050 o0 diff_4792_7153# GND GND efet w=493 l=16
+ ad=24276 pd=1720 as=0 ps=0 
M1051 diff_4792_7153# diff_5044_7399# GND GND efet w=274 l=16
+ ad=8484 pd=700 as=0 ps=0 
M1052 diff_4808_7162# diff_4792_7153# GND GND efet w=118 l=16
+ ad=5793 pd=424 as=0 ps=0 
M1053 diff_5039_7261# diff_4792_7153# GND GND efet w=58 l=16
+ ad=3418 pd=346 as=0 ps=0 
M1054 diff_5044_7399# diff_5128_7225# diff_5039_7261# GND efet w=31 l=16
+ ad=8675 pd=794 as=0 ps=0 
M1055 GND diff_5194_7252# diff_5044_7399# GND efet w=61 l=16
+ ad=0 pd=0 as=0 ps=0 
M1056 diff_4808_7162# diff_4808_7162# diff_4808_7162# GND efet w=7 l=10
+ ad=0 pd=0 as=0 ps=0 
M1057 diff_4808_7162# diff_4808_7162# diff_4808_7162# GND efet w=2 l=3
+ ad=0 pd=0 as=0 ps=0 
M1058 o0 diff_4808_7162# Vdd GND efet w=527 l=14
+ ad=0 pd=0 as=0 ps=0 
M1059 d0 diff_3328_7249# Vdd GND efet w=1520 l=16
+ ad=0 pd=0 as=0 ps=0 
M1060 diff_3154_7144# diff_3154_7144# diff_3154_7144# GND efet w=4 l=8
+ ad=1264 pd=166 as=0 ps=0 
M1061 diff_3154_7144# diff_3154_7144# diff_3154_7144# GND efet w=2 l=12
+ ad=0 pd=0 as=0 ps=0 
M1062 diff_3397_7141# diff_3397_7141# diff_3397_7141# GND efet w=4 l=8
+ ad=1183 pd=160 as=0 ps=0 
M1063 Vdd Vdd Vdd GND efet w=5 l=12
+ ad=0 pd=0 as=0 ps=0 
M1064 diff_1144_7198# diff_556_2707# diff_629_6919# GND efet w=71 l=16
+ ad=0 pd=0 as=0 ps=0 
M1065 Vdd Vdd diff_2522_7033# GND efet w=19 l=91
+ ad=0 pd=0 as=0 ps=0 
M1066 diff_872_2743# diff_2522_7033# Vdd GND efet w=91 l=16
+ ad=69513 pd=6156 as=0 ps=0 
M1067 GND diff_2359_7109# diff_872_2743# GND efet w=95 l=17
+ ad=0 pd=0 as=0 ps=0 
M1068 diff_3154_7144# Vdd Vdd GND efet w=23 l=20
+ ad=0 pd=0 as=0 ps=0 
M1069 diff_3397_7141# diff_3397_7141# diff_3397_7141# GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M1070 diff_3328_7249# diff_3397_7141# Vdd GND efet w=22 l=19
+ ad=0 pd=0 as=0 ps=0 
M1071 Vdd Vdd diff_3397_7141# GND efet w=17 l=19
+ ad=0 pd=0 as=0 ps=0 
M1072 Vdd Vdd Vdd GND efet w=1 l=1
+ ad=0 pd=0 as=0 ps=0 
M1073 diff_4808_7162# Vdd Vdd GND efet w=22 l=46
+ ad=0 pd=0 as=0 ps=0 
M1074 diff_5039_7261# Vdd Vdd GND efet w=16 l=73
+ ad=0 pd=0 as=0 ps=0 
M1075 GND diff_5188_6931# diff_5128_7225# GND efet w=31 l=16
+ ad=0 pd=0 as=1766 ps=186 
M1076 diff_5128_7225# Vdd Vdd GND efet w=17 l=140
+ ad=0 pd=0 as=0 ps=0 
M1077 Vdd Vdd Vdd GND efet w=10 l=19
+ ad=0 pd=0 as=0 ps=0 
M1078 Vdd Vdd Vdd GND efet w=10 l=9
+ ad=0 pd=0 as=0 ps=0 
M1079 diff_4792_7153# Vdd Vdd GND efet w=26 l=44
+ ad=0 pd=0 as=0 ps=0 
M1080 GND diff_6040_7132# diff_5935_6883# GND efet w=121 l=16
+ ad=0 pd=0 as=7081 ps=464 
M1081 GND diff_6040_7132# o1 GND efet w=505 l=13
+ ad=0 pd=0 as=26088 ps=1762 
M1082 diff_5044_7399# diff_5188_6931# diff_5263_6937# GND efet w=46 l=14
+ ad=0 pd=0 as=1784 ps=198 
M1083 Vdd diff_172_5905# d2 GND efet w=1556 l=14
+ ad=0 pd=0 as=120149 ps=7670 
M1084 GND diff_175_6337# d2 GND efet w=2861 l=9
+ ad=0 pd=0 as=0 ps=0 
M1085 diff_3574_7198# diff_556_2707# diff_872_2743# GND efet w=64 l=16
+ ad=4836 pd=422 as=0 ps=0 
M1086 diff_5263_6937# clk2 diff_872_2743# GND efet w=43 l=16
+ ad=0 pd=0 as=0 ps=0 
M1087 diff_5935_6883# Vdd Vdd GND efet w=25 l=46
+ ad=0 pd=0 as=0 ps=0 
M1088 diff_5935_6883# diff_5935_6883# diff_5935_6883# GND efet w=8 l=8
+ ad=0 pd=0 as=0 ps=0 
M1089 o1 diff_5935_6883# Vdd GND efet w=521 l=14
+ ad=0 pd=0 as=0 ps=0 
M1090 GND diff_6040_7132# diff_6134_6844# GND efet w=64 l=19
+ ad=0 pd=0 as=4012 ps=370 
M1091 diff_6134_6844# Vdd Vdd GND efet w=25 l=70
+ ad=0 pd=0 as=0 ps=0 
M1092 Vdd Vdd Vdd GND efet w=7 l=19
+ ad=0 pd=0 as=0 ps=0 
M1093 Vdd Vdd Vdd GND efet w=7 l=19
+ ad=0 pd=0 as=0 ps=0 
M1094 diff_6134_6844# diff_6059_6787# diff_5864_6631# GND efet w=34 l=19
+ ad=0 pd=0 as=9695 ps=812 
M1095 diff_6059_6787# Vdd Vdd GND efet w=19 l=142
+ ad=2072 pd=198 as=0 ps=0 
M1096 GND diff_5864_6631# diff_6040_7132# GND efet w=277 l=11
+ ad=0 pd=0 as=8748 ps=682 
M1097 diff_6059_6787# diff_5188_6931# GND GND efet w=35 l=14
+ ad=0 pd=0 as=0 ps=0 
M1098 diff_5864_6631# diff_5194_7252# GND GND efet w=61 l=14
+ ad=0 pd=0 as=0 ps=0 
M1099 Vdd Vdd Vdd GND efet w=5 l=8
+ ad=0 pd=0 as=0 ps=0 
M1100 diff_1217_6508# diff_817_6145# diff_872_2743# GND efet w=94 l=16
+ ad=6227 pd=566 as=0 ps=0 
M1101 diff_1217_6508# diff_1309_3670# diff_1267_6511# GND efet w=94 l=16
+ ad=0 pd=0 as=10577 ps=848 
M1102 diff_1370_6508# diff_1066_3979# diff_1217_6508# GND efet w=113 l=17
+ ad=19066 pd=2152 as=0 ps=0 
M1103 Vdd Vdd Vdd GND efet w=5 l=15
+ ad=0 pd=0 as=0 ps=0 
M1104 diff_5813_6613# clk2 diff_629_6919# GND efet w=49 l=16
+ ad=2003 pd=204 as=0 ps=0 
M1105 diff_5864_6631# diff_5188_6931# diff_5813_6613# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M1106 diff_1418_6481# Vdd Vdd GND efet w=19 l=73
+ ad=5480 pd=564 as=0 ps=0 
M1107 Vdd diff_1660_6529# diff_1267_6511# GND efet w=37 l=16
+ ad=0 pd=0 as=0 ps=0 
M1108 diff_1418_6481# diff_1060_6050# diff_1370_6508# GND efet w=79 l=16
+ ad=0 pd=0 as=0 ps=0 
M1109 diff_1217_6388# diff_817_6145# diff_629_6919# GND efet w=94 l=16
+ ad=6221 pd=566 as=0 ps=0 
M1110 diff_1418_6383# diff_1060_6050# diff_1370_6335# GND efet w=77 l=17
+ ad=5498 pd=546 as=19147 ps=2206 
M1111 diff_1267_6511# diff_1418_6481# GND GND efet w=136 l=19
+ ad=0 pd=0 as=0 ps=0 
M1112 diff_1418_6481# diff_1660_6529# GND GND efet w=65 l=17
+ ad=0 pd=0 as=0 ps=0 
M1113 GND diff_1418_6383# diff_1267_6334# GND efet w=133 l=19
+ ad=0 pd=0 as=10535 ps=830 
M1114 diff_2033_6463# diff_2011_6529# GND GND efet w=55 l=16
+ ad=1541 pd=180 as=0 ps=0 
M1115 diff_1370_6508# diff_2110_3745# diff_2011_6529# GND efet w=22 l=16
+ ad=0 pd=0 as=1545 ps=182 
M1116 diff_1660_6529# diff_2020_3610# diff_2033_6463# GND efet w=52 l=19
+ ad=38820 pd=3768 as=0 ps=0 
M1117 diff_1663_6337# diff_2020_3610# diff_2033_6358# GND efet w=53 l=22
+ ad=36930 pd=3786 as=1544 ps=186 
M1118 diff_172_5905# diff_220_6232# GND GND efet w=536 l=14
+ ad=25279 pd=1968 as=0 ps=0 
M1119 diff_220_6232# diff_220_6232# diff_220_6232# GND efet w=3 l=13
+ ad=6925 pd=538 as=0 ps=0 
M1120 diff_220_6232# diff_220_6232# diff_220_6232# GND efet w=6 l=7
+ ad=0 pd=0 as=0 ps=0 
M1121 diff_577_5317# diff_556_2707# diff_220_6232# GND efet w=67 l=16
+ ad=69359 pd=6174 as=0 ps=0 
M1122 diff_1217_6229# diff_817_6145# diff_577_5317# GND efet w=94 l=16
+ ad=6035 pd=566 as=0 ps=0 
M1123 diff_1217_6388# diff_1309_3670# diff_1267_6334# GND efet w=94 l=16
+ ad=0 pd=0 as=0 ps=0 
M1124 diff_1370_6335# diff_1066_3979# diff_1217_6388# GND efet w=110 l=17
+ ad=0 pd=0 as=0 ps=0 
M1125 GND diff_1663_6337# diff_1418_6383# GND efet w=64 l=16
+ ad=0 pd=0 as=0 ps=0 
M1126 GND diff_817_6145# diff_1102_6116# GND efet w=128 l=17
+ ad=0 pd=0 as=3785 ps=318 
M1127 diff_1217_6229# diff_1309_3670# diff_1267_6169# GND efet w=91 l=16
+ ad=0 pd=0 as=10418 ps=806 
M1128 diff_1370_6154# diff_1066_3979# diff_1217_6229# GND efet w=110 l=17
+ ad=18610 pd=2140 as=0 ps=0 
M1129 Vdd diff_1663_6337# diff_1267_6334# GND efet w=35 l=16
+ ad=0 pd=0 as=0 ps=0 
M1130 diff_2033_6358# diff_2011_6322# GND GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1131 diff_1418_6383# Vdd Vdd GND efet w=16 l=67
+ ad=0 pd=0 as=0 ps=0 
M1132 Vdd Vdd Vdd GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M1133 Vdd Vdd Vdd GND efet w=8 l=26
+ ad=0 pd=0 as=0 ps=0 
M1134 diff_1418_6127# Vdd Vdd GND efet w=16 l=67
+ ad=5765 pd=582 as=0 ps=0 
M1135 diff_1418_6127# diff_1060_6050# diff_1370_6154# GND efet w=79 l=16
+ ad=0 pd=0 as=0 ps=0 
M1136 diff_1102_6116# diff_1066_3979# diff_1060_6050# GND efet w=119 l=17
+ ad=0 pd=0 as=5945 ps=510 
M1137 diff_172_5905# diff_220_5722# GND GND efet w=536 l=17
+ ad=0 pd=0 as=0 ps=0 
M1138 Vdd diff_406_5971# diff_172_5905# GND efet w=25 l=19
+ ad=0 pd=0 as=0 ps=0 
M1139 Vdd Vdd diff_1060_6050# GND efet w=28 l=95
+ ad=0 pd=0 as=0 ps=0 
M1140 diff_172_5905# diff_406_5971# diff_172_5905# GND efet w=118 l=44
+ ad=0 pd=0 as=0 ps=0 
M1141 diff_406_5971# diff_406_5971# diff_406_5971# GND efet w=6 l=16
+ ad=1429 pd=188 as=0 ps=0 
M1142 Vdd Vdd diff_406_5971# GND efet w=22 l=19
+ ad=0 pd=0 as=0 ps=0 
M1143 diff_406_5971# diff_406_5971# diff_406_5971# GND efet w=3 l=7
+ ad=0 pd=0 as=0 ps=0 
M1144 Vdd Vdd Vdd GND efet w=5 l=15
+ ad=0 pd=0 as=0 ps=0 
M1145 Vdd Vdd Vdd GND efet w=3 l=7
+ ad=0 pd=0 as=0 ps=0 
M1146 Vdd diff_1660_6178# diff_1267_6169# GND efet w=31 l=14
+ ad=0 pd=0 as=0 ps=0 
M1147 diff_1267_6169# diff_1418_6127# GND GND efet w=128 l=17
+ ad=0 pd=0 as=0 ps=0 
M1148 diff_2201_6535# diff_2182_3644# diff_1370_6508# GND efet w=22 l=16
+ ad=1500 pd=182 as=0 ps=0 
M1149 diff_2378_6463# diff_2353_6529# GND GND efet w=55 l=22
+ ad=1517 pd=186 as=0 ps=0 
M1150 diff_2261_6454# diff_2236_3644# diff_1660_6529# GND efet w=52 l=16
+ ad=1682 pd=192 as=0 ps=0 
M1151 GND diff_2201_6535# diff_2261_6454# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1152 diff_1370_6508# diff_2455_3644# diff_2353_6529# GND efet w=23 l=16
+ ad=0 pd=0 as=1536 ps=182 
M1153 diff_1660_6529# diff_2365_3607# diff_2378_6463# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1154 diff_2261_6370# diff_2236_3644# diff_1663_6337# GND efet w=52 l=16
+ ad=1706 pd=192 as=0 ps=0 
M1155 diff_1663_6337# diff_2365_3607# diff_2377_6413# GND efet w=52 l=20
+ ad=0 pd=0 as=1547 ps=194 
M1156 GND diff_2201_6322# diff_2261_6370# GND efet w=56 l=17
+ ad=0 pd=0 as=0 ps=0 
M1157 diff_1370_6335# diff_2110_3745# diff_2011_6322# GND efet w=19 l=16
+ ad=0 pd=0 as=1533 ps=188 
M1158 diff_2201_6322# diff_2182_3644# diff_1370_6335# GND efet w=19 l=16
+ ad=1386 pd=182 as=0 ps=0 
M1159 diff_1418_6127# diff_1660_6178# GND GND efet w=64 l=16
+ ad=0 pd=0 as=0 ps=0 
M1160 diff_1418_6026# diff_1060_6050# diff_1370_5981# GND efet w=79 l=17
+ ad=5756 pd=582 as=18841 ps=2158 
M1161 diff_2033_6109# diff_2011_6175# GND GND efet w=55 l=16
+ ad=1487 pd=180 as=0 ps=0 
M1162 diff_1370_6154# diff_2110_3745# diff_2011_6175# GND efet w=19 l=16
+ ad=0 pd=0 as=1440 ps=182 
M1163 diff_1660_6178# diff_2020_3610# diff_2033_6109# GND efet w=52 l=19
+ ad=38946 pd=3774 as=0 ps=0 
M1164 diff_1663_5983# diff_2020_3610# diff_2033_6004# GND efet w=53 l=17
+ ad=37776 pd=3798 as=1559 ps=192 
M1165 GND diff_1418_6026# diff_1267_5983# GND efet w=124 l=16
+ ad=0 pd=0 as=10229 ps=812 
M1166 GND diff_1663_5983# diff_1418_6026# GND efet w=64 l=19
+ ad=0 pd=0 as=0 ps=0 
M1167 diff_175_6337# diff_172_5905# GND GND efet w=196 l=13
+ ad=20149 pd=1524 as=0 ps=0 
M1168 diff_1217_5923# diff_817_6145# diff_580_3394# GND efet w=94 l=16
+ ad=6086 pd=566 as=74853 ps=6748 
M1169 diff_1217_5923# diff_1309_3670# diff_1267_5983# GND efet w=92 l=17
+ ad=0 pd=0 as=0 ps=0 
M1170 diff_1370_5981# diff_1066_3979# diff_1217_5923# GND efet w=112 l=19
+ ad=0 pd=0 as=0 ps=0 
M1171 Vdd diff_1663_5983# diff_1267_5983# GND efet w=32 l=17
+ ad=0 pd=0 as=0 ps=0 
M1172 diff_2033_6004# diff_2011_5968# GND GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M1173 diff_175_6337# diff_220_5722# GND GND efet w=537 l=20
+ ad=0 pd=0 as=0 ps=0 
M1174 Vdd diff_406_5716# diff_175_6337# GND efet w=26 l=17
+ ad=0 pd=0 as=0 ps=0 
M1175 diff_175_6337# diff_406_5716# diff_175_6337# GND efet w=98 l=41
+ ad=0 pd=0 as=0 ps=0 
M1176 diff_406_5716# diff_406_5716# diff_406_5716# GND efet w=5 l=15
+ ad=1348 pd=184 as=0 ps=0 
M1177 Vdd Vdd diff_406_5716# GND efet w=19 l=19
+ ad=0 pd=0 as=0 ps=0 
M1178 diff_1217_5782# diff_820_3511# diff_872_2743# GND efet w=94 l=16
+ ad=6887 pd=626 as=0 ps=0 
M1179 diff_1217_5782# diff_1309_3670# diff_1267_5803# GND efet w=97 l=16
+ ad=0 pd=0 as=10160 ps=836 
M1180 diff_1418_6026# Vdd Vdd GND efet w=16 l=67
+ ad=0 pd=0 as=0 ps=0 
M1181 Vdd Vdd Vdd GND efet w=7 l=25
+ ad=0 pd=0 as=0 ps=0 
M1182 Vdd Vdd Vdd GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M1183 diff_1370_5800# diff_1066_3979# diff_1217_5782# GND efet w=110 l=17
+ ad=18574 pd=2158 as=0 ps=0 
M1184 diff_1418_5773# Vdd Vdd GND efet w=16 l=70
+ ad=5330 pd=546 as=0 ps=0 
M1185 Vdd diff_1663_5821# diff_1267_5803# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M1186 diff_1418_5773# diff_1060_5345# diff_1370_5800# GND efet w=79 l=16
+ ad=0 pd=0 as=0 ps=0 
M1187 diff_406_5716# diff_406_5716# diff_406_5716# GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M1188 diff_1217_5647# diff_820_3511# diff_629_6919# GND efet w=91 l=16
+ ad=6020 pd=572 as=0 ps=0 
M1189 diff_1418_5684# diff_1060_5345# diff_1370_5630# GND efet w=77 l=17
+ ad=5309 pd=540 as=18571 ps=2140 
M1190 diff_1267_5803# diff_1418_5773# GND GND efet w=134 l=17
+ ad=0 pd=0 as=0 ps=0 
M1191 diff_2201_6181# diff_2182_3644# diff_1370_6154# GND efet w=19 l=16
+ ad=1422 pd=182 as=0 ps=0 
M1192 diff_2377_6413# diff_2353_6322# GND GND efet w=55 l=17
+ ad=0 pd=0 as=0 ps=0 
M1193 diff_2261_6100# diff_2236_3644# diff_1660_6178# GND efet w=52 l=16
+ ad=1679 pd=186 as=0 ps=0 
M1194 GND diff_2201_6181# diff_2261_6100# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1195 diff_2375_6109# diff_2353_6178# GND GND efet w=56 l=17
+ ad=1658 pd=186 as=0 ps=0 
M1196 diff_2543_6535# diff_2524_3644# diff_1370_6508# GND efet w=22 l=16
+ ad=1476 pd=188 as=0 ps=0 
M1197 diff_2606_6454# diff_2581_3644# diff_1660_6529# GND efet w=52 l=16
+ ad=1526 pd=186 as=0 ps=0 
M1198 GND diff_2543_6535# diff_2606_6454# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1199 diff_2720_6463# diff_2698_6529# GND GND efet w=55 l=16
+ ad=1523 pd=180 as=0 ps=0 
M1200 diff_1370_6508# diff_2797_3745# diff_2698_6529# GND efet w=22 l=16
+ ad=0 pd=0 as=1545 ps=182 
M1201 diff_2888_6535# diff_2869_3644# diff_1370_6508# GND efet w=26 l=14
+ ad=1479 pd=176 as=0 ps=0 
M1202 diff_1660_6529# diff_2707_3610# diff_2720_6463# GND efet w=52 l=19
+ ad=0 pd=0 as=0 ps=0 
M1203 diff_2606_6370# diff_2581_3644# diff_1663_6337# GND efet w=52 l=19
+ ad=1526 pd=186 as=0 ps=0 
M1204 diff_1663_6337# diff_2707_3610# diff_2720_6358# GND efet w=52 l=20
+ ad=0 pd=0 as=1523 ps=180 
M1205 diff_1370_6335# diff_2455_3644# diff_2353_6322# GND efet w=19 l=19
+ ad=0 pd=0 as=1551 ps=188 
M1206 diff_2543_6322# diff_2524_3644# diff_1370_6335# GND efet w=19 l=16
+ ad=1470 pd=188 as=0 ps=0 
M1207 diff_1370_6154# diff_2455_3644# diff_2353_6178# GND efet w=19 l=19
+ ad=0 pd=0 as=1416 ps=188 
M1208 diff_1660_6178# diff_2365_3607# diff_2375_6109# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1209 diff_2261_6019# diff_2236_3644# diff_1663_5983# GND efet w=52 l=16
+ ad=1718 pd=192 as=0 ps=0 
M1210 GND diff_2201_5968# diff_2261_6019# GND efet w=56 l=17
+ ad=0 pd=0 as=0 ps=0 
M1211 diff_1370_5981# diff_2110_3745# diff_2011_5968# GND efet w=19 l=16
+ ad=0 pd=0 as=1542 ps=188 
M1212 diff_2201_5968# diff_2182_3644# diff_1370_5981# GND efet w=19 l=16
+ ad=1464 pd=176 as=0 ps=0 
M1213 diff_1370_5800# diff_2110_3745# diff_2011_5821# GND efet w=19 l=16
+ ad=0 pd=0 as=1548 ps=182 
M1214 diff_1418_5773# diff_1663_5821# GND GND efet w=65 l=17
+ ad=0 pd=0 as=0 ps=0 
M1215 diff_2033_5755# diff_2011_5821# GND GND efet w=55 l=16
+ ad=1496 pd=180 as=0 ps=0 
M1216 GND diff_1418_5684# diff_1267_5629# GND efet w=124 l=19
+ ad=0 pd=0 as=10007 ps=800 
M1217 diff_1663_5821# diff_2020_3610# diff_2033_5755# GND efet w=52 l=19
+ ad=38886 pd=3774 as=0 ps=0 
M1218 diff_1217_5524# diff_820_3511# diff_577_5317# GND efet w=91 l=16
+ ad=6113 pd=566 as=0 ps=0 
M1219 diff_1217_5647# diff_1309_3670# diff_1267_5629# GND efet w=91 l=16
+ ad=0 pd=0 as=0 ps=0 
M1220 diff_1370_5630# diff_1066_3979# diff_1217_5647# GND efet w=115 l=16
+ ad=0 pd=0 as=0 ps=0 
M1221 GND diff_820_3511# diff_1102_5408# GND efet w=139 l=16
+ ad=0 pd=0 as=3494 ps=306 
M1222 diff_1217_5524# diff_1309_3670# diff_1267_5467# GND efet w=94 l=16
+ ad=0 pd=0 as=10199 ps=818 
M1223 diff_1370_5446# diff_1066_3979# diff_1217_5524# GND efet w=112 l=16
+ ad=18790 pd=2158 as=0 ps=0 
M1224 GND diff_1663_5629# diff_1418_5684# GND efet w=64 l=16
+ ad=0 pd=0 as=0 ps=0 
M1225 diff_1267_5629# diff_1663_5629# Vdd GND efet w=32 l=16
+ ad=0 pd=0 as=0 ps=0 
M1226 diff_2033_5650# diff_2011_5614# GND GND efet w=58 l=16
+ ad=1550 pd=186 as=0 ps=0 
M1227 diff_1663_5629# diff_2020_3610# diff_2033_5650# GND efet w=52 l=19
+ ad=36654 pd=3738 as=0 ps=0 
M1228 diff_1418_5684# Vdd Vdd GND efet w=13 l=64
+ ad=0 pd=0 as=0 ps=0 
M1229 Vdd Vdd Vdd GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M1230 Vdd Vdd Vdd GND efet w=7 l=19
+ ad=0 pd=0 as=0 ps=0 
M1231 diff_1421_5419# Vdd Vdd GND efet w=13 l=64
+ ad=5759 pd=582 as=0 ps=0 
M1232 diff_1421_5419# diff_1060_5345# diff_1370_5446# GND efet w=82 l=19
+ ad=0 pd=0 as=0 ps=0 
M1233 diff_1102_5408# diff_1066_3979# diff_1060_5345# GND efet w=115 l=19
+ ad=0 pd=0 as=5786 ps=510 
M1234 GND diff_407_5030# diff_577_5317# GND efet w=94 l=16
+ ad=0 pd=0 as=0 ps=0 
M1235 d2 GND GND GND efet w=262 l=16
+ ad=0 pd=0 as=0 ps=0 
M1236 diff_577_5317# diff_425_5110# Vdd GND efet w=94 l=16
+ ad=0 pd=0 as=0 ps=0 
M1237 Vdd Vdd diff_1060_5345# GND efet w=28 l=94
+ ad=0 pd=0 as=0 ps=0 
M1238 Vdd Vdd Vdd GND efet w=5 l=15
+ ad=0 pd=0 as=0 ps=0 
M1239 Vdd Vdd Vdd GND efet w=3 l=7
+ ad=0 pd=0 as=0 ps=0 
M1240 Vdd diff_1663_5467# diff_1267_5467# GND efet w=32 l=17
+ ad=0 pd=0 as=0 ps=0 
M1241 diff_1267_5467# diff_1421_5419# GND GND efet w=130 l=19
+ ad=0 pd=0 as=0 ps=0 
M1242 diff_2201_5827# diff_2182_3644# diff_1370_5800# GND efet w=19 l=16
+ ad=1482 pd=176 as=0 ps=0 
M1243 diff_2375_6020# diff_2353_5968# GND GND efet w=62 l=20
+ ad=1655 pd=198 as=0 ps=0 
M1244 diff_1663_5983# diff_2365_3607# diff_2375_6020# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1245 diff_2261_5746# diff_2236_3644# diff_1663_5821# GND efet w=52 l=16
+ ad=1682 pd=192 as=0 ps=0 
M1246 GND diff_2201_5827# diff_2261_5746# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1247 diff_2378_5755# diff_2353_5824# GND GND efet w=55 l=19
+ ad=1514 pd=180 as=0 ps=0 
M1248 diff_2543_6181# diff_2524_3644# diff_1370_6154# GND efet w=19 l=16
+ ad=1455 pd=194 as=0 ps=0 
M1249 GND diff_2543_6322# diff_2606_6370# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1250 diff_2720_6358# diff_2695_6331# GND GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1251 diff_2606_6100# diff_2581_3644# diff_1660_6178# GND efet w=52 l=16
+ ad=1523 pd=180 as=0 ps=0 
M1252 GND diff_2543_6181# diff_2606_6100# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1253 diff_2720_6109# diff_2698_6175# GND GND efet w=55 l=16
+ ad=1505 pd=180 as=0 ps=0 
M1254 diff_2948_6454# diff_2923_3644# diff_1660_6529# GND efet w=52 l=16
+ ad=1688 pd=186 as=0 ps=0 
M1255 GND diff_2888_6535# diff_2948_6454# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1256 diff_3065_6463# diff_3040_6529# GND GND efet w=55 l=19
+ ad=1517 pd=186 as=0 ps=0 
M1257 diff_1370_6508# diff_3142_3644# diff_3040_6529# GND efet w=22 l=17
+ ad=0 pd=0 as=1467 ps=188 
M1258 diff_1660_6529# diff_3052_3607# diff_3065_6463# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1259 diff_2948_6370# diff_2923_3644# diff_1663_6337# GND efet w=52 l=16
+ ad=1688 pd=186 as=0 ps=0 
M1260 diff_1370_6335# diff_2797_3745# diff_2695_6331# GND efet w=19 l=16
+ ad=0 pd=0 as=1521 ps=182 
M1261 diff_2888_6322# diff_2869_3644# diff_1370_6335# GND efet w=22 l=16
+ ad=1446 pd=176 as=0 ps=0 
M1262 diff_1370_6154# diff_2797_3745# diff_2698_6175# GND efet w=19 l=16
+ ad=0 pd=0 as=1530 ps=182 
M1263 diff_2888_6181# diff_2869_3644# diff_1370_6154# GND efet w=20 l=16
+ ad=1422 pd=182 as=0 ps=0 
M1264 diff_1660_6178# diff_2707_3610# diff_2720_6109# GND efet w=52 l=19
+ ad=0 pd=0 as=0 ps=0 
M1265 diff_2606_6019# diff_2581_3644# diff_1663_5983# GND efet w=52 l=16
+ ad=1571 pd=186 as=0 ps=0 
M1266 diff_2720_6004# diff_2698_5968# GND GND efet w=56 l=17
+ ad=1565 pd=186 as=0 ps=0 
M1267 diff_2543_5968# diff_2524_3644# diff_1370_5981# GND efet w=19 l=17
+ ad=1470 pd=188 as=0 ps=0 
M1268 diff_1370_5981# diff_2455_3644# diff_2353_5968# GND efet w=19 l=19
+ ad=0 pd=0 as=1515 ps=188 
M1269 diff_1370_5800# diff_2455_3644# diff_2353_5824# GND efet w=19 l=19
+ ad=0 pd=0 as=1488 ps=188 
M1270 diff_1663_5821# diff_2365_3607# diff_2378_5755# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1271 diff_2261_5665# diff_2236_3644# diff_1663_5629# GND efet w=49 l=16
+ ad=1682 pd=186 as=0 ps=0 
M1272 diff_1663_5629# diff_2365_3607# diff_2378_5650# GND efet w=50 l=20
+ ad=0 pd=0 as=1541 ps=186 
M1273 GND diff_2201_5614# diff_2261_5665# GND efet w=56 l=17
+ ad=0 pd=0 as=0 ps=0 
M1274 diff_1370_5630# diff_2110_3745# diff_2011_5614# GND efet w=19 l=16
+ ad=0 pd=0 as=1503 ps=182 
M1275 diff_2201_5614# diff_2182_3644# diff_1370_5630# GND efet w=19 l=16
+ ad=1467 pd=182 as=0 ps=0 
M1276 diff_1370_5446# diff_2110_3745# diff_2011_5470# GND efet w=22 l=16
+ ad=0 pd=0 as=1491 ps=182 
M1277 diff_1421_5419# diff_1663_5467# GND GND efet w=65 l=17
+ ad=0 pd=0 as=0 ps=0 
M1278 diff_1421_5318# diff_1060_5345# diff_1370_5273# GND efet w=82 l=19
+ ad=5570 pd=582 as=18733 ps=2182 
M1279 GND diff_1421_5318# diff_1267_5275# GND efet w=128 l=16
+ ad=0 pd=0 as=10235 ps=806 
M1280 diff_2033_5401# diff_2011_5470# GND GND efet w=58 l=19
+ ad=1661 pd=186 as=0 ps=0 
M1281 diff_1663_5467# diff_2020_3610# diff_2033_5401# GND efet w=50 l=17
+ ad=38223 pd=3768 as=0 ps=0 
M1282 diff_1217_5215# diff_820_3511# diff_580_3394# GND efet w=95 l=17
+ ad=6257 pd=566 as=0 ps=0 
M1283 diff_425_5110# diff_407_5030# GND GND efet w=52 l=16
+ ad=9140 pd=690 as=0 ps=0 
M1284 diff_425_5110# diff_425_5110# diff_425_5110# GND efet w=4 l=7
+ ad=0 pd=0 as=0 ps=0 
M1285 diff_425_5110# diff_425_5110# diff_425_5110# GND efet w=5 l=18
+ ad=0 pd=0 as=0 ps=0 
M1286 Vdd Vdd diff_425_5110# GND efet w=19 l=91
+ ad=0 pd=0 as=0 ps=0 
M1287 diff_1217_5215# diff_1309_3670# diff_1267_5275# GND efet w=94 l=16
+ ad=0 pd=0 as=0 ps=0 
M1288 diff_1370_5273# diff_1066_3979# diff_1217_5215# GND efet w=110 l=17
+ ad=0 pd=0 as=0 ps=0 
M1289 GND diff_1663_5275# diff_1421_5318# GND efet w=67 l=19
+ ad=0 pd=0 as=0 ps=0 
M1290 diff_2033_5299# diff_2011_5260# GND GND efet w=55 l=16
+ ad=1661 pd=186 as=0 ps=0 
M1291 diff_1663_5275# diff_2020_3610# diff_2033_5299# GND efet w=52 l=16
+ ad=38679 pd=3792 as=0 ps=0 
M1292 diff_2201_5473# diff_2182_3644# diff_1370_5446# GND efet w=22 l=16
+ ad=1470 pd=176 as=0 ps=0 
M1293 diff_1267_5275# diff_1663_5275# Vdd GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M1294 diff_1421_5318# Vdd Vdd GND efet w=13 l=64
+ ad=0 pd=0 as=0 ps=0 
M1295 diff_407_5030# diff_407_5030# diff_407_5030# GND efet w=5 l=15
+ ad=7358 pd=706 as=0 ps=0 
M1296 diff_407_5030# diff_407_5030# diff_407_5030# GND efet w=3 l=16
+ ad=0 pd=0 as=0 ps=0 
M1297 diff_407_5030# d2 GND GND efet w=139 l=19
+ ad=0 pd=0 as=0 ps=0 
M1298 diff_425_5110# diff_331_7000# GND GND efet w=85 l=14
+ ad=0 pd=0 as=0 ps=0 
M1299 diff_1217_5074# diff_829_3778# diff_872_2743# GND efet w=94 l=16
+ ad=6842 pd=614 as=0 ps=0 
M1300 diff_1217_5074# diff_1309_3670# diff_1267_5095# GND efet w=94 l=16
+ ad=0 pd=0 as=10202 ps=812 
M1301 Vdd Vdd Vdd GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M1302 diff_1370_5092# diff_1066_3979# diff_1217_5074# GND efet w=110 l=17
+ ad=19078 pd=2152 as=0 ps=0 
M1303 Vdd Vdd Vdd GND efet w=7 l=19
+ ad=0 pd=0 as=0 ps=0 
M1304 diff_1421_5065# Vdd Vdd GND efet w=14 l=65
+ ad=5216 pd=546 as=0 ps=0 
M1305 Vdd diff_1663_5113# diff_1267_5095# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M1306 diff_1421_5065# diff_1060_4634# diff_1370_5092# GND efet w=77 l=17
+ ad=0 pd=0 as=0 ps=0 
M1307 GND diff_331_7000# diff_407_5030# GND efet w=85 l=14
+ ad=0 pd=0 as=0 ps=0 
M1308 GND GND GND GND efet w=0 l=1
+ ad=0 pd=0 as=0 ps=0 
M1309 Vdd Vdd Vdd GND efet w=5 l=18
+ ad=0 pd=0 as=0 ps=0 
M1310 Vdd Vdd Vdd GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M1311 Vdd Vdd diff_407_5030# GND efet w=19 l=88
+ ad=0 pd=0 as=0 ps=0 
M1312 diff_1217_4939# diff_829_3778# diff_629_6919# GND efet w=91 l=16
+ ad=6116 pd=554 as=0 ps=0 
M1313 diff_1267_5095# diff_1421_5065# GND GND efet w=130 l=19
+ ad=0 pd=0 as=0 ps=0 
M1314 diff_1421_5065# diff_1663_5113# GND GND efet w=68 l=17
+ ad=0 pd=0 as=0 ps=0 
M1315 diff_2033_5047# diff_2011_5113# GND GND efet w=59 l=17
+ ad=1694 pd=192 as=0 ps=0 
M1316 diff_2378_5650# diff_2353_5617# GND GND efet w=58 l=21
+ ad=0 pd=0 as=0 ps=0 
M1317 diff_2261_5392# diff_2236_3644# diff_1663_5467# GND efet w=55 l=18
+ ad=1559 pd=192 as=0 ps=0 
M1318 GND diff_2201_5473# diff_2261_5392# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1319 diff_2378_5401# diff_2353_5470# GND GND efet w=55 l=19
+ ad=1499 pd=186 as=0 ps=0 
M1320 diff_2543_5827# diff_2524_3644# diff_1370_5800# GND efet w=19 l=16
+ ad=1488 pd=188 as=0 ps=0 
M1321 GND diff_2543_5968# diff_2606_6019# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1322 diff_1663_5983# diff_2707_3610# diff_2720_6004# GND efet w=56 l=20
+ ad=0 pd=0 as=0 ps=0 
M1323 GND diff_2888_6322# diff_2948_6370# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1324 diff_3065_6358# diff_3040_6322# GND GND efet w=55 l=19
+ ad=1517 pd=186 as=0 ps=0 
M1325 diff_1663_6337# diff_3052_3607# diff_3065_6358# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1326 diff_2948_6100# diff_2923_3644# diff_1660_6178# GND efet w=52 l=16
+ ad=1670 pd=186 as=0 ps=0 
M1327 GND diff_2888_6181# diff_2948_6100# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1328 diff_3065_6109# diff_3040_6178# GND GND efet w=55 l=19
+ ad=1505 pd=180 as=0 ps=0 
M1329 diff_3230_6535# diff_3211_3644# diff_1370_6508# GND efet w=22 l=16
+ ad=1446 pd=182 as=0 ps=0 
M1330 diff_3293_6454# diff_3268_3644# diff_1660_6529# GND efet w=52 l=16
+ ad=1526 pd=186 as=0 ps=0 
M1331 GND diff_3230_6535# diff_3293_6454# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1332 diff_3407_6463# diff_3385_6529# GND GND efet w=55 l=16
+ ad=1505 pd=180 as=0 ps=0 
M1333 diff_1370_6508# diff_3484_3742# diff_3385_6529# GND efet w=22 l=16
+ ad=0 pd=0 as=1545 ps=182 
M1334 diff_1660_6529# diff_3394_3613# diff_3407_6463# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1335 diff_3293_6370# diff_3268_3644# diff_1663_6337# GND efet w=50 l=17
+ ad=1517 pd=186 as=0 ps=0 
M1336 diff_1370_6335# diff_3142_3644# diff_3040_6322# GND efet w=19 l=22
+ ad=0 pd=0 as=1422 ps=182 
M1337 diff_3230_6322# diff_3211_3644# diff_1370_6335# GND efet w=19 l=19
+ ad=1443 pd=188 as=0 ps=0 
M1338 diff_1370_6154# diff_3142_3644# diff_3040_6178# GND efet w=19 l=19
+ ad=0 pd=0 as=1431 ps=182 
M1339 diff_1660_6178# diff_3052_3607# diff_3065_6109# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1340 diff_2948_6019# diff_2923_3644# diff_1663_5983# GND efet w=50 l=16
+ ad=1691 pd=186 as=0 ps=0 
M1341 diff_1663_5983# diff_3052_3607# diff_3065_6004# GND efet w=52 l=22
+ ad=0 pd=0 as=1526 ps=186 
M1342 diff_1370_5981# diff_2797_3745# diff_2698_5968# GND efet w=19 l=16
+ ad=0 pd=0 as=1521 ps=182 
M1343 diff_2888_5968# diff_2869_3644# diff_1370_5981# GND efet w=22 l=19
+ ad=1464 pd=176 as=0 ps=0 
M1344 diff_2606_5746# diff_2581_3644# diff_1663_5821# GND efet w=52 l=16
+ ad=1526 pd=186 as=0 ps=0 
M1345 GND diff_2543_5827# diff_2606_5746# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1346 diff_2720_5755# diff_2698_5821# GND GND efet w=55 l=16
+ ad=1526 pd=186 as=0 ps=0 
M1347 diff_1370_5800# diff_2797_3745# diff_2698_5821# GND efet w=19 l=16
+ ad=0 pd=0 as=1539 ps=182 
M1348 diff_1663_5821# diff_2707_3610# diff_2720_5755# GND efet w=52 l=19
+ ad=0 pd=0 as=0 ps=0 
M1349 diff_2606_5662# diff_2581_3644# diff_1663_5629# GND efet w=52 l=22
+ ad=1544 pd=186 as=0 ps=0 
M1350 diff_1663_5629# diff_2707_3610# diff_2720_5650# GND efet w=50 l=23
+ ad=0 pd=0 as=1559 ps=186 
M1351 GND diff_2543_5614# diff_2606_5662# GND efet w=59 l=20
+ ad=0 pd=0 as=0 ps=0 
M1352 diff_2720_5650# diff_2698_5614# GND GND efet w=58 l=22
+ ad=0 pd=0 as=0 ps=0 
M1353 diff_1370_5630# diff_2455_3644# diff_2353_5617# GND efet w=22 l=19
+ ad=0 pd=0 as=1533 ps=200 
M1354 diff_2543_5614# diff_2524_3644# diff_1370_5630# GND efet w=19 l=16
+ ad=1554 pd=194 as=0 ps=0 
M1355 diff_1370_5446# diff_2455_3644# diff_2353_5470# GND efet w=25 l=17
+ ad=0 pd=0 as=1521 ps=200 
M1356 diff_2543_5473# diff_2524_3644# diff_1370_5446# GND efet w=22 l=16
+ ad=1476 pd=188 as=0 ps=0 
M1357 diff_1663_5467# diff_2365_3607# diff_2378_5401# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1358 diff_2261_5345# diff_2236_3644# diff_1663_5275# GND efet w=58 l=19
+ ad=1580 pd=192 as=0 ps=0 
M1359 GND diff_2201_5263# diff_2261_5345# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1360 diff_2378_5299# diff_2353_5260# GND GND efet w=55 l=19
+ ad=1514 pd=180 as=0 ps=0 
M1361 diff_1663_5275# diff_2365_3607# diff_2378_5299# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1362 diff_1370_5273# diff_2110_3745# diff_2011_5260# GND efet w=22 l=17
+ ad=0 pd=0 as=1548 ps=182 
M1363 diff_2201_5263# diff_2182_3644# diff_1370_5273# GND efet w=19 l=16
+ ad=1455 pd=176 as=0 ps=0 
M1364 diff_1370_5092# diff_2110_3745# diff_2011_5113# GND efet w=20 l=20
+ ad=0 pd=0 as=1542 ps=188 
M1365 diff_2201_5119# diff_2182_3644# diff_1370_5092# GND efet w=20 l=17
+ ad=1479 pd=176 as=0 ps=0 
M1366 diff_1421_4961# diff_1060_4634# diff_1370_4919# GND efet w=79 l=22
+ ad=5312 pd=540 as=19012 ps=2260 
M1367 GND diff_1421_4961# diff_1267_4921# GND efet w=127 l=16
+ ad=0 pd=0 as=9920 ps=812 
M1368 diff_1663_5113# diff_2020_3610# diff_2033_5047# GND efet w=52 l=16
+ ad=38595 pd=3768 as=0 ps=0 
M1369 Vdd diff_172_3988# d3 GND efet w=1529 l=14
+ ad=0 pd=0 as=118679 ps=7568 
M1370 GND diff_175_4780# d3 GND efet w=2867 l=9
+ ad=0 pd=0 as=0 ps=0 
M1371 diff_1217_4813# diff_829_3778# diff_577_5317# GND efet w=94 l=16
+ ad=6323 pd=578 as=0 ps=0 
M1372 diff_1217_4939# diff_1309_3670# diff_1267_4921# GND efet w=91 l=16
+ ad=0 pd=0 as=0 ps=0 
M1373 diff_1370_4919# diff_1066_3979# diff_1217_4939# GND efet w=110 l=17
+ ad=0 pd=0 as=0 ps=0 
M1374 diff_1217_4813# diff_1309_3670# diff_1267_4756# GND efet w=100 l=16
+ ad=0 pd=0 as=10130 ps=818 
M1375 GND diff_829_3778# diff_1102_4697# GND efet w=130 l=14
+ ad=0 pd=0 as=3593 ps=312 
M1376 GND diff_1663_4918# diff_1421_4961# GND efet w=64 l=16
+ ad=0 pd=0 as=0 ps=0 
M1377 diff_1267_4921# diff_1663_4918# Vdd GND efet w=34 l=14
+ ad=0 pd=0 as=0 ps=0 
M1378 diff_2033_4942# diff_2011_4906# GND GND efet w=58 l=16
+ ad=1724 pd=192 as=0 ps=0 
M1379 diff_1663_4918# diff_2020_3610# diff_2033_4942# GND efet w=52 l=16
+ ad=36900 pd=3756 as=0 ps=0 
M1380 Vdd Vdd Vdd GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M1381 diff_1370_4735# diff_1066_3979# diff_1217_4813# GND efet w=113 l=17
+ ad=18979 pd=2182 as=0 ps=0 
M1382 diff_1421_4961# Vdd Vdd GND efet w=16 l=64
+ ad=0 pd=0 as=0 ps=0 
M1383 Vdd Vdd Vdd GND efet w=7 l=19
+ ad=0 pd=0 as=0 ps=0 
M1384 diff_1421_4708# Vdd Vdd GND efet w=17 l=65
+ ad=5855 pd=582 as=0 ps=0 
M1385 diff_1102_4697# diff_1066_3979# diff_1060_4634# GND efet w=125 l=17
+ ad=0 pd=0 as=5954 ps=528 
M1386 Vdd Vdd diff_1060_4634# GND efet w=26 l=95
+ ad=0 pd=0 as=0 ps=0 
M1387 Vdd Vdd Vdd GND efet w=5 l=15
+ ad=0 pd=0 as=0 ps=0 
M1388 Vdd Vdd Vdd GND efet w=4 l=7
+ ad=0 pd=0 as=0 ps=0 
M1389 diff_1421_4708# diff_1060_4634# diff_1370_4735# GND efet w=80 l=17
+ ad=0 pd=0 as=0 ps=0 
M1390 Vdd diff_1663_4756# diff_1267_4756# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M1391 diff_1267_4756# diff_1421_4708# GND GND efet w=127 l=19
+ ad=0 pd=0 as=0 ps=0 
M1392 diff_1421_4708# diff_1663_4756# GND GND efet w=65 l=17
+ ad=0 pd=0 as=0 ps=0 
M1393 diff_2033_4693# diff_2011_4759# GND GND efet w=55 l=16
+ ad=1673 pd=186 as=0 ps=0 
M1394 diff_1370_4919# diff_2110_3745# diff_2011_4906# GND efet w=29 l=37
+ ad=0 pd=0 as=1503 ps=182 
M1395 diff_2264_5038# diff_2236_3644# diff_1663_5113# GND efet w=52 l=19
+ ad=1526 pd=186 as=0 ps=0 
M1396 GND diff_2201_5119# diff_2264_5038# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1397 diff_2378_5047# diff_2353_5113# GND GND efet w=59 l=17
+ ad=1517 pd=186 as=0 ps=0 
M1398 diff_2606_5392# diff_2581_3644# diff_1663_5467# GND efet w=52 l=16
+ ad=1514 pd=180 as=0 ps=0 
M1399 GND diff_2543_5473# diff_2606_5392# GND efet w=56 l=17
+ ad=0 pd=0 as=0 ps=0 
M1400 diff_2720_5401# diff_2698_5470# GND GND efet w=55 l=16
+ ad=1496 pd=180 as=0 ps=0 
M1401 diff_2888_5827# diff_2869_3644# diff_1370_5800# GND efet w=19 l=19
+ ad=1482 pd=176 as=0 ps=0 
M1402 GND diff_2888_5968# diff_2948_6019# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1403 diff_3065_6004# diff_3040_5968# GND GND efet w=55 l=19
+ ad=0 pd=0 as=0 ps=0 
M1404 diff_2948_5746# diff_2923_3644# diff_1663_5821# GND efet w=64 l=16
+ ad=1676 pd=210 as=0 ps=0 
M1405 GND diff_2888_5827# diff_2948_5746# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1406 diff_3065_5755# diff_3040_5824# GND GND efet w=55 l=19
+ ad=1505 pd=180 as=0 ps=0 
M1407 diff_3230_6181# diff_3211_3644# diff_1370_6154# GND efet w=19 l=16
+ ad=1461 pd=188 as=0 ps=0 
M1408 GND diff_3230_6322# diff_3293_6370# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1409 diff_3407_6358# diff_3385_6322# GND GND efet w=55 l=16
+ ad=1505 pd=180 as=0 ps=0 
M1410 diff_1663_6337# diff_3394_3613# diff_3407_6358# GND efet w=50 l=17
+ ad=0 pd=0 as=0 ps=0 
M1411 diff_3293_6100# diff_3268_3644# diff_1660_6178# GND efet w=52 l=16
+ ad=1514 pd=180 as=0 ps=0 
M1412 GND diff_3230_6181# diff_3293_6100# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1413 diff_3407_6109# diff_3385_6175# GND GND efet w=55 l=16
+ ad=1505 pd=180 as=0 ps=0 
M1414 diff_3575_6535# diff_3556_3644# diff_1370_6508# GND efet w=22 l=17
+ ad=1479 pd=176 as=0 ps=0 
M1415 diff_1370_6335# diff_3484_3742# diff_3385_6322# GND efet w=19 l=16
+ ad=0 pd=0 as=1494 ps=182 
M1416 diff_3635_6454# diff_3610_3644# diff_1660_6529# GND efet w=52 l=16
+ ad=1679 pd=186 as=0 ps=0 
M1417 GND diff_3575_6535# diff_3635_6454# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1418 diff_3752_6463# diff_3727_6532# GND GND efet w=55 l=19
+ ad=1505 pd=180 as=0 ps=0 
M1419 diff_1370_6508# diff_3829_3644# diff_3727_6532# GND efet w=23 l=19
+ ad=0 pd=0 as=1467 ps=188 
M1420 diff_3917_6535# diff_3898_3644# diff_1370_6508# GND efet w=20 l=17
+ ad=1536 pd=182 as=0 ps=0 
M1421 diff_1660_6529# diff_3739_3610# diff_3752_6463# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1422 diff_3635_6370# diff_3610_3644# diff_1663_6337# GND efet w=50 l=17
+ ad=1670 pd=186 as=0 ps=0 
M1423 diff_3575_6322# diff_3556_3644# diff_1370_6335# GND efet w=19 l=19
+ ad=1449 pd=182 as=0 ps=0 
M1424 diff_1370_6154# diff_3484_3742# diff_3385_6175# GND efet w=19 l=16
+ ad=0 pd=0 as=1503 ps=182 
M1425 diff_1660_6178# diff_3394_3613# diff_3407_6109# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1426 diff_3293_6019# diff_3268_3644# diff_1663_5983# GND efet w=52 l=16
+ ad=1553 pd=186 as=0 ps=0 
M1427 diff_1663_5983# diff_3394_3613# diff_3407_6004# GND efet w=52 l=22
+ ad=0 pd=0 as=1526 ps=186 
M1428 diff_1370_5981# diff_3142_3644# diff_3040_5968# GND efet w=19 l=19
+ ad=0 pd=0 as=1452 ps=188 
M1429 diff_3230_5968# diff_3211_3644# diff_1370_5981# GND efet w=19 l=16
+ ad=1470 pd=188 as=0 ps=0 
M1430 diff_1370_5800# diff_3142_3644# diff_3040_5824# GND efet w=19 l=19
+ ad=0 pd=0 as=1479 ps=188 
M1431 diff_1663_5821# diff_3052_3607# diff_3065_5755# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1432 diff_2948_5669# diff_2923_3644# diff_1663_5629# GND efet w=55 l=19
+ ad=1664 pd=192 as=0 ps=0 
M1433 GND diff_2888_5614# diff_2948_5669# GND efet w=56 l=17
+ ad=0 pd=0 as=0 ps=0 
M1434 diff_3065_5650# diff_3040_5617# GND GND efet w=58 l=19
+ ad=1493 pd=186 as=0 ps=0 
M1435 diff_1663_5629# diff_3052_3607# diff_3065_5650# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M1436 diff_1370_5630# diff_2797_3745# diff_2698_5614# GND efet w=19 l=16
+ ad=0 pd=0 as=1542 ps=188 
M1437 diff_2888_5614# diff_2869_3644# diff_1370_5630# GND efet w=22 l=17
+ ad=1455 pd=176 as=0 ps=0 
M1438 diff_1370_5446# diff_2797_3745# diff_2698_5470# GND efet w=22 l=16
+ ad=0 pd=0 as=1575 ps=188 
M1439 diff_1663_5467# diff_2707_3610# diff_2720_5401# GND efet w=52 l=19
+ ad=0 pd=0 as=0 ps=0 
M1440 diff_2606_5311# diff_2581_3644# diff_1663_5275# GND efet w=52 l=16
+ ad=1505 pd=180 as=0 ps=0 
M1441 diff_1370_5273# diff_2455_3644# diff_2353_5260# GND efet w=23 l=16
+ ad=0 pd=0 as=1539 ps=200 
M1442 diff_2543_5263# diff_2524_3644# diff_1370_5273# GND efet w=19 l=16
+ ad=1452 pd=188 as=0 ps=0 
M1443 diff_1370_5092# diff_2455_3644# diff_2353_5113# GND efet w=19 l=16
+ ad=0 pd=0 as=1530 ps=182 
M1444 diff_1663_5113# diff_2365_3607# diff_2378_5047# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1445 diff_2264_4954# diff_2236_3644# diff_1663_4918# GND efet w=53 l=20
+ ad=1568 pd=186 as=0 ps=0 
M1446 GND diff_2201_4906# diff_2264_4954# GND efet w=56 l=17
+ ad=0 pd=0 as=0 ps=0 
M1447 diff_2201_4906# diff_2182_3644# diff_1370_4919# GND efet w=19 l=16
+ ad=1512 pd=182 as=0 ps=0 
M1448 diff_1370_4735# diff_2110_3745# diff_2011_4759# GND efet w=19 l=19
+ ad=0 pd=0 as=1512 ps=182 
M1449 diff_1421_4607# diff_1060_4634# diff_1370_4565# GND efet w=77 l=16
+ ad=5759 pd=582 as=18682 ps=2164 
M1450 diff_1663_4756# diff_2020_3610# diff_2033_4693# GND efet w=49 l=16
+ ad=38025 pd=3738 as=0 ps=0 
M1451 GND diff_1421_4607# diff_1267_4564# GND efet w=127 l=19
+ ad=0 pd=0 as=10238 ps=806 
M1452 GND diff_1663_4564# diff_1421_4607# GND efet w=67 l=16
+ ad=0 pd=0 as=0 ps=0 
M1453 diff_1217_4504# diff_829_3778# diff_580_3394# GND efet w=95 l=17
+ ad=6350 pd=572 as=0 ps=0 
M1454 diff_1217_4504# diff_1309_3670# diff_1267_4564# GND efet w=94 l=16
+ ad=0 pd=0 as=0 ps=0 
M1455 diff_1370_4565# diff_1066_3979# diff_1217_4504# GND efet w=110 l=17
+ ad=0 pd=0 as=0 ps=0 
M1456 diff_1267_4564# diff_1663_4564# Vdd GND efet w=32 l=17
+ ad=0 pd=0 as=0 ps=0 
M1457 diff_2033_4588# diff_2011_4549# GND GND efet w=55 l=16
+ ad=1661 pd=186 as=0 ps=0 
M1458 diff_1663_4564# diff_2020_3610# diff_2033_4588# GND efet w=52 l=16
+ ad=38637 pd=3762 as=0 ps=0 
M1459 diff_172_3988# diff_223_4213# GND GND efet w=544 l=16
+ ad=25771 pd=1992 as=0 ps=0 
M1460 diff_1217_4351# diff_1093_4033# diff_872_2743# GND efet w=91 l=16
+ ad=7169 pd=644 as=0 ps=0 
M1461 diff_1217_4351# diff_1309_3670# diff_1267_4369# GND efet w=97 l=16
+ ad=0 pd=0 as=10331 ps=836 
M1462 diff_1421_4607# Vdd Vdd GND efet w=14 l=67
+ ad=0 pd=0 as=0 ps=0 
M1463 Vdd Vdd Vdd GND efet w=13 l=9
+ ad=0 pd=0 as=0 ps=0 
M1464 diff_1370_4381# diff_1066_3979# diff_1217_4351# GND efet w=110 l=17
+ ad=18874 pd=2140 as=0 ps=0 
M1465 Vdd Vdd Vdd GND efet w=7 l=19
+ ad=0 pd=0 as=0 ps=0 
M1466 diff_1421_4354# Vdd Vdd GND efet w=13 l=64
+ ad=5255 pd=540 as=0 ps=0 
M1467 Vdd diff_1663_4402# diff_1267_4369# GND efet w=32 l=16
+ ad=0 pd=0 as=0 ps=0 
M1468 diff_223_4213# diff_223_4213# diff_223_4213# GND efet w=5 l=9
+ ad=7060 pd=532 as=0 ps=0 
M1469 diff_223_4213# diff_223_4213# diff_223_4213# GND efet w=7 l=10
+ ad=0 pd=0 as=0 ps=0 
M1470 diff_580_3394# diff_556_2707# diff_223_4213# GND efet w=67 l=16
+ ad=0 pd=0 as=0 ps=0 
M1471 diff_1217_4228# diff_1093_4033# diff_629_6919# GND efet w=91 l=16
+ ad=6110 pd=566 as=0 ps=0 
M1472 diff_1421_4354# diff_1060_3926# diff_1370_4381# GND efet w=76 l=16
+ ad=0 pd=0 as=0 ps=0 
M1473 diff_1421_4253# diff_1060_3926# diff_1370_4211# GND efet w=77 l=17
+ ad=5219 pd=540 as=18889 ps=2158 
M1474 diff_1267_4369# diff_1421_4354# GND GND efet w=124 l=16
+ ad=0 pd=0 as=0 ps=0 
M1475 diff_1421_4354# diff_1663_4402# GND GND efet w=64 l=16
+ ad=0 pd=0 as=0 ps=0 
M1476 GND diff_1421_4253# diff_1267_4210# GND efet w=127 l=16
+ ad=0 pd=0 as=9950 ps=806 
M1477 diff_2033_4336# diff_2011_4402# GND GND efet w=62 l=17
+ ad=1718 pd=198 as=0 ps=0 
M1478 diff_2201_4765# diff_2182_3644# diff_1370_4735# GND efet w=19 l=16
+ ad=1464 pd=176 as=0 ps=0 
M1479 diff_2378_4942# diff_2353_4906# GND GND efet w=64 l=16
+ ad=1559 pd=186 as=0 ps=0 
M1480 diff_1663_4918# diff_2365_3607# diff_2378_4942# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1481 diff_2264_4681# diff_2236_3644# diff_1663_4756# GND efet w=53 l=20
+ ad=1592 pd=186 as=0 ps=0 
M1482 GND diff_2201_4765# diff_2264_4681# GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M1483 diff_2378_4690# diff_2353_4759# GND GND efet w=62 l=17
+ ad=1541 pd=186 as=0 ps=0 
M1484 diff_2543_5122# diff_2524_3644# diff_1370_5092# GND efet w=19 l=16
+ ad=1431 pd=182 as=0 ps=0 
M1485 diff_1370_4919# diff_2455_3644# diff_2353_4906# GND efet w=19 l=16
+ ad=0 pd=0 as=1599 ps=194 
M1486 GND diff_2543_5263# diff_2606_5311# GND efet w=55 l=17
+ ad=0 pd=0 as=0 ps=0 
M1487 diff_2720_5299# diff_2698_5260# GND GND efet w=55 l=16
+ ad=1505 pd=180 as=0 ps=0 
M1488 diff_1663_5275# diff_2707_3610# diff_2720_5299# GND efet w=52 l=19
+ ad=0 pd=0 as=0 ps=0 
M1489 diff_2888_5473# diff_2869_3644# diff_1370_5446# GND efet w=22 l=16
+ ad=1395 pd=170 as=0 ps=0 
M1490 diff_2951_5392# diff_2923_3644# diff_1663_5467# GND efet w=52 l=19
+ ad=1523 pd=180 as=0 ps=0 
M1491 GND diff_2888_5473# diff_2951_5392# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1492 diff_3065_5401# diff_3040_5470# GND GND efet w=55 l=19
+ ad=1499 pd=186 as=0 ps=0 
M1493 diff_3230_5827# diff_3211_3644# diff_1370_5800# GND efet w=19 l=16
+ ad=1461 pd=188 as=0 ps=0 
M1494 GND diff_3230_5968# diff_3293_6019# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1495 diff_3407_6004# diff_3385_5968# GND GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1496 diff_3293_5746# diff_3268_3644# diff_1663_5821# GND efet w=52 l=16
+ ad=1517 pd=186 as=0 ps=0 
M1497 GND diff_3230_5827# diff_3293_5746# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1498 diff_3407_5755# diff_3385_5821# GND GND efet w=55 l=16
+ ad=1496 pd=180 as=0 ps=0 
M1499 diff_3575_6181# diff_3556_3644# diff_1370_6154# GND efet w=19 l=19
+ ad=1455 pd=176 as=0 ps=0 
M1500 GND diff_3575_6322# diff_3635_6370# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1501 diff_3752_6358# diff_3727_6322# GND GND efet w=55 l=19
+ ad=1505 pd=180 as=0 ps=0 
M1502 diff_1663_6337# diff_3739_3610# diff_3752_6358# GND efet w=50 l=17
+ ad=0 pd=0 as=0 ps=0 
M1503 diff_3635_6100# diff_3610_3644# diff_1660_6178# GND efet w=52 l=16
+ ad=1661 pd=186 as=0 ps=0 
M1504 GND diff_3575_6181# diff_3635_6100# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1505 diff_3752_6109# diff_3727_6178# GND GND efet w=55 l=19
+ ad=1505 pd=180 as=0 ps=0 
M1506 diff_3980_6454# diff_3955_3644# diff_1660_6529# GND efet w=52 l=16
+ ad=1505 pd=180 as=0 ps=0 
M1507 GND diff_3917_6535# diff_3980_6454# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1508 diff_4094_6463# diff_4072_6529# GND GND efet w=55 l=16
+ ad=1514 pd=180 as=0 ps=0 
M1509 diff_1370_6508# diff_4171_3745# diff_4072_6529# GND efet w=20 l=17
+ ad=0 pd=0 as=1452 ps=188 
M1510 diff_4262_6535# diff_4243_3644# diff_1370_6508# GND efet w=20 l=17
+ ad=1455 pd=182 as=0 ps=0 
M1511 diff_1660_6529# diff_4084_3607# diff_4094_6463# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1512 diff_3980_6370# diff_3955_3644# diff_1663_6337# GND efet w=50 l=17
+ ad=1505 pd=180 as=0 ps=0 
M1513 diff_1370_6335# diff_3829_3644# diff_3727_6322# GND efet w=19 l=19
+ ad=0 pd=0 as=1437 ps=176 
M1514 diff_3917_6322# diff_3898_3644# diff_1370_6335# GND efet w=19 l=16
+ ad=1512 pd=182 as=0 ps=0 
M1515 diff_1370_6154# diff_3829_3644# diff_3727_6178# GND efet w=19 l=19
+ ad=0 pd=0 as=1398 ps=188 
M1516 diff_3917_6181# diff_3898_3644# diff_1370_6154# GND efet w=19 l=16
+ ad=1440 pd=182 as=0 ps=0 
M1517 diff_1660_6178# diff_3739_3610# diff_3752_6109# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1518 diff_3635_6019# diff_3610_3644# diff_1663_5983# GND efet w=49 l=16
+ ad=1655 pd=186 as=0 ps=0 
M1519 diff_1370_5981# diff_3484_3742# diff_3385_5968# GND efet w=19 l=16
+ ad=0 pd=0 as=1503 ps=182 
M1520 diff_3575_5968# diff_3556_3644# diff_1370_5981# GND efet w=19 l=19
+ ad=1446 pd=176 as=0 ps=0 
M1521 diff_1370_5800# diff_3484_3742# diff_3385_5821# GND efet w=19 l=16
+ ad=0 pd=0 as=1521 ps=182 
M1522 diff_1663_5821# diff_3394_3613# diff_3407_5755# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1523 diff_3293_5665# diff_3268_3644# diff_1663_5629# GND efet w=49 l=16
+ ad=1511 pd=186 as=0 ps=0 
M1524 diff_1370_5630# diff_3142_3644# diff_3040_5617# GND efet w=19 l=19
+ ad=0 pd=0 as=1443 ps=188 
M1525 diff_3230_5614# diff_3211_3644# diff_1370_5630# GND efet w=19 l=16
+ ad=1443 pd=188 as=0 ps=0 
M1526 diff_1370_5446# diff_3142_3644# diff_3040_5470# GND efet w=19 l=19
+ ad=0 pd=0 as=1461 ps=188 
M1527 diff_1663_5467# diff_3052_3607# diff_3065_5401# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1528 diff_2951_5311# diff_2923_3644# diff_1663_5275# GND efet w=52 l=19
+ ad=1514 pd=180 as=0 ps=0 
M1529 diff_1370_5273# diff_2797_3745# diff_2698_5260# GND efet w=19 l=16
+ ad=0 pd=0 as=1512 ps=182 
M1530 diff_2606_5038# diff_2581_3644# diff_1663_5113# GND efet w=52 l=16
+ ad=1526 pd=186 as=0 ps=0 
M1531 GND diff_2543_5122# diff_2606_5038# GND efet w=55 l=19
+ ad=0 pd=0 as=0 ps=0 
M1532 diff_2720_5047# diff_2698_5113# GND GND efet w=55 l=16
+ ad=1505 pd=180 as=0 ps=0 
M1533 diff_2888_5263# diff_2869_3644# diff_1370_5273# GND efet w=19 l=16
+ ad=1464 pd=176 as=0 ps=0 
M1534 diff_1370_5092# diff_2797_3745# diff_2698_5113# GND efet w=19 l=16
+ ad=0 pd=0 as=1530 ps=182 
M1535 diff_1663_5113# diff_2707_3610# diff_2720_5047# GND efet w=52 l=19
+ ad=0 pd=0 as=0 ps=0 
M1536 diff_2606_4954# diff_2581_3644# diff_1663_4918# GND efet w=53 l=17
+ ad=1565 pd=186 as=0 ps=0 
M1537 diff_1663_4918# diff_2707_3610# diff_2720_4942# GND efet w=53 l=20
+ ad=0 pd=0 as=1568 ps=192 
M1538 GND diff_2543_4906# diff_2606_4954# GND efet w=56 l=23
+ ad=0 pd=0 as=0 ps=0 
M1539 diff_2720_4942# diff_2698_4903# GND GND efet w=55 l=19
+ ad=0 pd=0 as=0 ps=0 
M1540 diff_2543_4906# diff_2524_3644# diff_1370_4919# GND efet w=19 l=16
+ ad=1482 pd=194 as=0 ps=0 
M1541 diff_1370_4735# diff_2455_3644# diff_2353_4759# GND efet w=20 l=17
+ ad=0 pd=0 as=1530 ps=200 
M1542 diff_2543_4765# diff_2524_3644# diff_1370_4735# GND efet w=19 l=16
+ ad=1443 pd=188 as=0 ps=0 
M1543 diff_1663_4756# diff_2365_3607# diff_2378_4690# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1544 diff_2264_4600# diff_2236_3644# diff_1663_4564# GND efet w=52 l=19
+ ad=1514 pd=180 as=0 ps=0 
M1545 diff_1370_4565# diff_2110_3745# diff_2011_4549# GND efet w=19 l=19
+ ad=0 pd=0 as=1533 ps=188 
M1546 diff_2201_4552# diff_2182_3644# diff_1370_4565# GND efet w=19 l=16
+ ad=1485 pd=182 as=0 ps=0 
M1547 GND diff_2201_4552# diff_2264_4600# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1548 diff_2378_4588# diff_2353_4549# GND GND efet w=55 l=16
+ ad=1514 pd=180 as=0 ps=0 
M1549 diff_1663_4564# diff_2365_3607# diff_2378_4588# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1550 diff_1370_4381# diff_2110_3745# diff_2011_4402# GND efet w=19 l=19
+ ad=0 pd=0 as=1521 ps=182 
M1551 diff_1663_4402# diff_2020_3610# diff_2033_4336# GND efet w=52 l=16
+ ad=38430 pd=3762 as=0 ps=0 
M1552 diff_1217_4228# diff_1309_3670# diff_1267_4210# GND efet w=95 l=17
+ ad=0 pd=0 as=0 ps=0 
M1553 diff_172_3988# diff_220_5722# GND GND efet w=544 l=16
+ ad=0 pd=0 as=0 ps=0 
M1554 Vdd diff_406_4054# diff_172_3988# GND efet w=25 l=17
+ ad=0 pd=0 as=0 ps=0 
M1555 diff_172_3988# diff_406_4054# diff_172_3988# GND efet w=121 l=41
+ ad=0 pd=0 as=0 ps=0 
M1556 diff_406_4054# diff_406_4054# diff_406_4054# GND efet w=5 l=18
+ ad=1381 pd=196 as=0 ps=0 
M1557 Vdd Vdd diff_406_4054# GND efet w=19 l=16
+ ad=0 pd=0 as=0 ps=0 
M1558 diff_406_4054# diff_406_4054# diff_406_4054# GND efet w=7 l=8
+ ad=0 pd=0 as=0 ps=0 
M1559 diff_175_4780# diff_172_3988# GND GND efet w=196 l=13
+ ad=19903 pd=1518 as=0 ps=0 
M1560 diff_175_4780# diff_220_5722# GND GND efet w=535 l=17
+ ad=0 pd=0 as=0 ps=0 
M1561 diff_175_4780# diff_406_3802# diff_175_4780# GND efet w=95 l=45
+ ad=0 pd=0 as=0 ps=0 
M1562 Vdd diff_406_3802# diff_175_4780# GND efet w=25 l=19
+ ad=0 pd=0 as=0 ps=0 
M1563 diff_406_3802# diff_406_3802# diff_406_3802# GND efet w=5 l=21
+ ad=1273 pd=170 as=0 ps=0 
M1564 Vdd Vdd diff_406_3802# GND efet w=19 l=19
+ ad=0 pd=0 as=0 ps=0 
M1565 diff_406_3802# diff_406_3802# diff_406_3802# GND efet w=0 l=5
+ ad=0 pd=0 as=0 ps=0 
M1566 diff_1217_4105# diff_1093_4033# diff_577_5317# GND efet w=91 l=16
+ ad=5918 pd=560 as=0 ps=0 
M1567 diff_1370_4211# diff_1066_3979# diff_1217_4228# GND efet w=112 l=19
+ ad=0 pd=0 as=0 ps=0 
M1568 GND diff_1093_4033# diff_1102_3989# GND efet w=130 l=14
+ ad=0 pd=0 as=3656 ps=312 
M1569 diff_1217_4105# diff_1309_3670# diff_1267_4048# GND efet w=94 l=19
+ ad=0 pd=0 as=10160 ps=812 
M1570 diff_1370_4027# diff_1066_3979# diff_1217_4105# GND efet w=110 l=17
+ ad=18385 pd=2146 as=0 ps=0 
M1571 GND diff_1663_4210# diff_1421_4253# GND efet w=68 l=17
+ ad=0 pd=0 as=0 ps=0 
M1572 diff_1267_4210# diff_1663_4210# Vdd GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M1573 diff_2033_4231# diff_2011_4195# GND GND efet w=61 l=16
+ ad=1703 pd=198 as=0 ps=0 
M1574 diff_1663_4210# diff_2020_3610# diff_2033_4231# GND efet w=52 l=16
+ ad=36825 pd=3804 as=0 ps=0 
M1575 diff_1421_4253# Vdd Vdd GND efet w=13 l=64
+ ad=0 pd=0 as=0 ps=0 
M1576 Vdd Vdd Vdd GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M1577 Vdd Vdd Vdd GND efet w=7 l=19
+ ad=0 pd=0 as=0 ps=0 
M1578 diff_1421_4000# Vdd Vdd GND efet w=16 l=67
+ ad=5516 pd=570 as=0 ps=0 
M1579 diff_1421_4000# diff_1060_3926# diff_1370_4027# GND efet w=83 l=20
+ ad=0 pd=0 as=0 ps=0 
M1580 diff_1102_3989# diff_1066_3979# diff_1060_3926# GND efet w=115 l=16
+ ad=0 pd=0 as=6035 ps=510 
M1581 Vdd Vdd diff_1060_3926# GND efet w=28 l=97
+ ad=0 pd=0 as=0 ps=0 
M1582 Vdd Vdd Vdd GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M1583 Vdd Vdd Vdd GND efet w=1 l=1
+ ad=0 pd=0 as=0 ps=0 
M1584 Vdd Vdd Vdd GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M1585 Vdd diff_1663_4051# diff_1267_4048# GND efet w=32 l=17
+ ad=0 pd=0 as=0 ps=0 
M1586 diff_1267_4048# diff_1421_4000# GND GND efet w=127 l=16
+ ad=0 pd=0 as=0 ps=0 
M1587 diff_1421_4000# diff_1663_4051# GND GND efet w=64 l=19
+ ad=0 pd=0 as=0 ps=0 
M1588 diff_1421_3899# diff_1060_3926# diff_1370_3857# GND efet w=79 l=16
+ ad=5744 pd=576 as=18844 ps=2146 
M1589 diff_2033_3992# diff_2011_4051# GND GND efet w=61 l=17
+ ad=1520 pd=192 as=0 ps=0 
M1590 diff_2201_4411# diff_2182_3644# diff_1370_4381# GND efet w=19 l=16
+ ad=1473 pd=176 as=0 ps=0 
M1591 diff_1370_4211# diff_2110_3745# diff_2011_4195# GND efet w=19 l=19
+ ad=0 pd=0 as=1512 ps=182 
M1592 GND diff_2201_4411# diff_2264_4327# GND efet w=56 l=17
+ ad=0 pd=0 as=1523 ps=186 
M1593 diff_2378_4336# diff_2353_4405# GND GND efet w=62 l=17
+ ad=1559 pd=186 as=0 ps=0 
M1594 diff_2264_4327# diff_2236_3644# diff_1663_4402# GND efet w=56 l=20
+ ad=0 pd=0 as=0 ps=0 
M1595 diff_2888_5122# diff_2869_3644# diff_1370_5092# GND efet w=19 l=16
+ ad=1464 pd=176 as=0 ps=0 
M1596 diff_1370_4919# diff_2797_3745# diff_2698_4903# GND efet w=19 l=16
+ ad=0 pd=0 as=1578 ps=188 
M1597 GND diff_2888_5263# diff_2951_5311# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1598 diff_3065_5299# diff_3040_5260# GND GND efet w=55 l=17
+ ad=1496 pd=180 as=0 ps=0 
M1599 diff_1663_5275# diff_3052_3607# diff_3065_5299# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1600 diff_2951_5038# diff_2923_3644# diff_1663_5113# GND efet w=52 l=19
+ ad=1505 pd=180 as=0 ps=0 
M1601 GND diff_2888_5122# diff_2951_5038# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1602 diff_3065_5047# diff_3040_5113# GND GND efet w=62 l=17
+ ad=1508 pd=186 as=0 ps=0 
M1603 diff_3230_5473# diff_3211_3644# diff_1370_5446# GND efet w=19 l=16
+ ad=1479 pd=188 as=0 ps=0 
M1604 GND diff_3230_5614# diff_3293_5665# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1605 diff_3407_5650# diff_3385_5614# GND GND efet w=55 l=16
+ ad=1517 pd=180 as=0 ps=0 
M1606 diff_1663_5629# diff_3394_3613# diff_3407_5650# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M1607 diff_3575_5827# diff_3556_3644# diff_1370_5800# GND efet w=19 l=19
+ ad=1449 pd=182 as=0 ps=0 
M1608 GND diff_3575_5968# diff_3635_6019# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1609 diff_3749_6050# diff_3727_5968# GND GND efet w=58 l=17
+ ad=1490 pd=192 as=0 ps=0 
M1610 diff_1663_5983# diff_3739_3610# diff_3749_6050# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M1611 diff_3635_5746# diff_3610_3644# diff_1663_5821# GND efet w=52 l=16
+ ad=1652 pd=186 as=0 ps=0 
M1612 GND diff_3575_5827# diff_3635_5746# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1613 diff_3752_5755# diff_3727_5824# GND GND efet w=55 l=19
+ ad=1514 pd=180 as=0 ps=0 
M1614 GND diff_3917_6322# diff_3980_6370# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1615 diff_4094_6358# diff_4072_6322# GND GND efet w=55 l=16
+ ad=1517 pd=186 as=0 ps=0 
M1616 diff_1663_6337# diff_4084_3607# diff_4094_6358# GND efet w=50 l=17
+ ad=0 pd=0 as=0 ps=0 
M1617 diff_3980_6100# diff_3955_3644# diff_1660_6178# GND efet w=52 l=16
+ ad=1514 pd=180 as=0 ps=0 
M1618 GND diff_3917_6181# diff_3980_6100# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1619 diff_4094_6109# diff_4072_6178# GND GND efet w=55 l=16
+ ad=1514 pd=180 as=0 ps=0 
M1620 diff_1370_6335# diff_4171_3745# diff_4072_6322# GND efet w=19 l=16
+ ad=0 pd=0 as=1422 ps=182 
M1621 diff_4322_6470# diff_4300_3644# diff_1660_6529# GND efet w=62 l=17
+ ad=1598 pd=210 as=0 ps=0 
M1622 GND diff_4262_6535# diff_4322_6470# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1623 diff_4439_6463# diff_4414_6532# GND GND efet w=55 l=16
+ ad=1517 pd=186 as=0 ps=0 
M1624 diff_1370_6508# diff_4516_3742# diff_4414_6532# GND efet w=22 l=16
+ ad=0 pd=0 as=1521 ps=188 
M1625 diff_4604_6554# diff_4588_3644# diff_1370_6508# GND efet w=23 l=17
+ ad=1476 pd=194 as=0 ps=0 
M1626 diff_1660_6529# diff_4426_3610# diff_4439_6463# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1627 diff_4322_6370# diff_4300_3644# diff_1663_6337# GND efet w=61 l=17
+ ad=1661 pd=210 as=0 ps=0 
M1628 diff_4262_6322# diff_4243_3644# diff_1370_6335# GND efet w=19 l=16
+ ad=1443 pd=188 as=0 ps=0 
M1629 diff_1370_6154# diff_4171_3745# diff_4072_6178# GND efet w=19 l=16
+ ad=0 pd=0 as=1425 ps=188 
M1630 diff_1660_6178# diff_4084_3607# diff_4094_6109# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1631 diff_3980_6019# diff_3955_3644# diff_1663_5983# GND efet w=49 l=17
+ ad=1529 pd=186 as=0 ps=0 
M1632 GND diff_3917_5968# diff_3980_6019# GND efet w=55 l=19
+ ad=0 pd=0 as=0 ps=0 
M1633 diff_1370_5981# diff_3829_3644# diff_3727_5968# GND efet w=19 l=17
+ ad=0 pd=0 as=1455 ps=176 
M1634 diff_3917_5968# diff_3898_3644# diff_1370_5981# GND efet w=19 l=16
+ ad=1512 pd=182 as=0 ps=0 
M1635 diff_1370_5800# diff_3829_3644# diff_3727_5824# GND efet w=19 l=19
+ ad=0 pd=0 as=1476 ps=182 
M1636 diff_1663_5821# diff_3739_3610# diff_3752_5755# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1637 diff_3635_5665# diff_3610_3644# diff_1663_5629# GND efet w=49 l=16
+ ad=1664 pd=186 as=0 ps=0 
M1638 diff_1370_5630# diff_3484_3742# diff_3385_5614# GND efet w=19 l=16
+ ad=0 pd=0 as=1506 ps=188 
M1639 diff_3575_5614# diff_3556_3644# diff_1370_5630# GND efet w=19 l=19
+ ad=1437 pd=176 as=0 ps=0 
M1640 diff_3293_5392# diff_3268_3644# diff_1663_5467# GND efet w=52 l=16
+ ad=1508 pd=186 as=0 ps=0 
M1641 GND diff_3230_5473# diff_3293_5392# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1642 diff_3407_5401# diff_3385_5470# GND GND efet w=55 l=16
+ ad=1496 pd=180 as=0 ps=0 
M1643 diff_1370_5446# diff_3484_3742# diff_3385_5470# GND efet w=19 l=16
+ ad=0 pd=0 as=1464 ps=194 
M1644 diff_1663_5467# diff_3394_3613# diff_3407_5401# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1645 diff_3293_5311# diff_3268_3644# diff_1663_5275# GND efet w=52 l=16
+ ad=1514 pd=180 as=0 ps=0 
M1646 diff_3230_5263# diff_3211_3644# diff_1370_5273# GND efet w=25 l=30
+ ad=1470 pd=206 as=0 ps=0 
M1647 diff_1370_5273# diff_3142_3644# diff_3040_5260# GND efet w=19 l=19
+ ad=0 pd=0 as=1470 ps=188 
M1648 diff_1370_5092# diff_3142_3644# diff_3040_5113# GND efet w=19 l=16
+ ad=0 pd=0 as=1536 ps=194 
M1649 diff_1663_5113# diff_3052_3607# diff_3065_5047# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1650 diff_2951_4954# diff_2923_3644# diff_1663_4918# GND efet w=52 l=22
+ ad=1514 pd=180 as=0 ps=0 
M1651 diff_1663_4918# diff_3052_3607# diff_3065_4942# GND efet w=50 l=20
+ ad=0 pd=0 as=1508 ps=186 
M1652 diff_2888_4906# diff_2869_3644# diff_1370_4919# GND efet w=19 l=16
+ ad=1512 pd=182 as=0 ps=0 
M1653 diff_2606_4681# diff_2581_3644# diff_1663_4756# GND efet w=52 l=16
+ ad=1577 pd=186 as=0 ps=0 
M1654 GND diff_2543_4765# diff_2606_4681# GND efet w=58 l=19
+ ad=0 pd=0 as=0 ps=0 
M1655 diff_2720_4690# diff_2698_4759# GND GND efet w=58 l=16
+ ad=1583 pd=192 as=0 ps=0 
M1656 diff_1370_4735# diff_2797_3745# diff_2698_4759# GND efet w=20 l=16
+ ad=0 pd=0 as=1533 ps=188 
M1657 diff_1663_4756# diff_2707_3610# diff_2720_4690# GND efet w=55 l=19
+ ad=0 pd=0 as=0 ps=0 
M1658 diff_2606_4600# diff_2581_3644# diff_1663_4564# GND efet w=52 l=16
+ ad=1523 pd=180 as=0 ps=0 
M1659 diff_1370_4565# diff_2455_3644# diff_2353_4549# GND efet w=19 l=16
+ ad=0 pd=0 as=1521 ps=200 
M1660 diff_2543_4552# diff_2524_3644# diff_1370_4565# GND efet w=19 l=16
+ ad=1446 pd=194 as=0 ps=0 
M1661 diff_1370_4381# diff_2455_3644# diff_2353_4405# GND efet w=19 l=16
+ ad=0 pd=0 as=1536 ps=194 
M1662 diff_1663_4402# diff_2365_3607# diff_2378_4336# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1663 diff_2264_4243# diff_2236_3644# diff_1663_4210# GND efet w=55 l=23
+ ad=1556 pd=180 as=0 ps=0 
M1664 diff_2201_4195# diff_2182_3644# diff_1370_4211# GND efet w=19 l=16
+ ad=1455 pd=176 as=0 ps=0 
M1665 GND diff_2201_4195# diff_2264_4243# GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M1666 diff_2378_4231# diff_2353_4195# GND GND efet w=62 l=17
+ ad=1565 pd=186 as=0 ps=0 
M1667 diff_1663_4210# diff_2365_3607# diff_2378_4231# GND efet w=53 l=17
+ ad=0 pd=0 as=0 ps=0 
M1668 diff_1370_4027# diff_2110_3745# diff_2011_4051# GND efet w=19 l=19
+ ad=0 pd=0 as=1512 ps=182 
M1669 diff_1663_4051# diff_2020_3610# diff_2033_3992# GND efet w=52 l=16
+ ad=37203 pd=3738 as=0 ps=0 
M1670 GND diff_1421_3899# diff_1267_3856# GND efet w=127 l=16
+ ad=0 pd=0 as=10433 ps=812 
M1671 diff_1217_3803# diff_1093_4033# diff_580_3394# GND efet w=98 l=20
+ ad=5855 pd=566 as=0 ps=0 
M1672 diff_1217_3803# diff_1309_3670# diff_1267_3856# GND efet w=91 l=19
+ ad=0 pd=0 as=0 ps=0 
M1673 diff_1370_3857# diff_1066_3979# diff_1217_3803# GND efet w=110 l=17
+ ad=0 pd=0 as=0 ps=0 
M1674 GND diff_1663_3859# diff_1421_3899# GND efet w=64 l=19
+ ad=0 pd=0 as=0 ps=0 
M1675 diff_1267_3856# diff_1663_3859# Vdd GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M1676 diff_2036_3880# diff_2011_3844# GND GND efet w=55 l=19
+ ad=1505 pd=180 as=0 ps=0 
M1677 diff_1663_3859# diff_2020_3610# diff_2036_3880# GND efet w=52 l=16
+ ad=37644 pd=3774 as=0 ps=0 
M1678 diff_1421_3899# Vdd Vdd GND efet w=14 l=65
+ ad=0 pd=0 as=0 ps=0 
M1679 Vdd Vdd Vdd GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M1680 Vdd Vdd Vdd GND efet w=3 l=13
+ ad=0 pd=0 as=0 ps=0 
M1681 diff_2201_4054# diff_2182_3644# diff_1370_4027# GND efet w=19 l=16
+ ad=1473 pd=176 as=0 ps=0 
M1682 diff_2264_3973# diff_2236_3644# diff_1663_4051# GND efet w=52 l=19
+ ad=1523 pd=180 as=0 ps=0 
M1683 GND diff_2201_4054# diff_2264_3973# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1684 diff_2378_3982# diff_2353_4051# GND GND efet w=62 l=17
+ ad=1505 pd=180 as=0 ps=0 
M1685 diff_2543_4411# diff_2524_3644# diff_1370_4381# GND efet w=19 l=16
+ ad=1512 pd=182 as=0 ps=0 
M1686 GND diff_2543_4552# diff_2606_4600# GND efet w=55 l=19
+ ad=0 pd=0 as=0 ps=0 
M1687 diff_2720_4588# diff_2698_4549# GND GND efet w=55 l=16
+ ad=1514 pd=180 as=0 ps=0 
M1688 diff_1663_4564# diff_2707_3610# diff_2720_4588# GND efet w=52 l=19
+ ad=0 pd=0 as=0 ps=0 
M1689 diff_2888_4765# diff_2869_3644# diff_1370_4735# GND efet w=19 l=16
+ ad=1464 pd=176 as=0 ps=0 
M1690 GND diff_2888_4906# diff_2951_4954# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1691 diff_3065_4942# diff_3040_4906# GND GND efet w=61 l=17
+ ad=0 pd=0 as=0 ps=0 
M1692 diff_3230_5122# diff_3211_3644# diff_1370_5092# GND efet w=19 l=16
+ ad=1467 pd=182 as=0 ps=0 
M1693 GND diff_3230_5263# diff_3293_5311# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1694 diff_3407_5299# diff_3385_5260# GND GND efet w=55 l=16
+ ad=1505 pd=180 as=0 ps=0 
M1695 diff_1663_5275# diff_3394_3613# diff_3407_5299# GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M1696 diff_3575_5473# diff_3556_3644# diff_1370_5446# GND efet w=19 l=19
+ ad=1464 pd=176 as=0 ps=0 
M1697 GND diff_3575_5614# diff_3635_5665# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1698 diff_3752_5650# diff_3727_5617# GND GND efet w=55 l=19
+ ad=1484 pd=186 as=0 ps=0 
M1699 diff_1663_5629# diff_3739_3610# diff_3752_5650# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M1700 diff_3917_5827# diff_3898_3644# diff_1370_5800# GND efet w=19 l=16
+ ad=1479 pd=188 as=0 ps=0 
M1701 diff_3635_5392# diff_3610_3644# diff_1663_5467# GND efet w=52 l=16
+ ad=1661 pd=186 as=0 ps=0 
M1702 GND diff_3575_5473# diff_3635_5392# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1703 diff_3752_5401# diff_3727_5470# GND GND efet w=55 l=19
+ ad=1499 pd=186 as=0 ps=0 
M1704 diff_4094_6004# diff_4072_5968# GND GND efet w=55 l=16
+ ad=1502 pd=186 as=0 ps=0 
M1705 diff_1663_5983# diff_4084_3607# diff_4094_6004# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M1706 diff_3980_5746# diff_3955_3644# diff_1663_5821# GND efet w=52 l=16
+ ad=1505 pd=180 as=0 ps=0 
M1707 GND diff_3917_5827# diff_3980_5746# GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M1708 diff_4094_5755# diff_4072_5821# GND GND efet w=55 l=16
+ ad=1514 pd=180 as=0 ps=0 
M1709 diff_4262_6181# diff_4243_3644# diff_1370_6154# GND efet w=19 l=16
+ ad=1422 pd=182 as=0 ps=0 
M1710 GND diff_4262_6322# diff_4322_6370# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1711 diff_4439_6358# diff_4414_6325# GND GND efet w=55 l=16
+ ad=1517 pd=186 as=0 ps=0 
M1712 diff_1663_6337# diff_4426_3610# diff_4439_6358# GND efet w=50 l=17
+ ad=0 pd=0 as=0 ps=0 
M1713 diff_4322_6100# diff_4300_3644# diff_1660_6178# GND efet w=52 l=16
+ ad=1670 pd=186 as=0 ps=0 
M1714 GND diff_4262_6181# diff_4322_6100# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1715 diff_4439_6109# diff_4414_6178# GND GND efet w=55 l=16
+ ad=1514 pd=180 as=0 ps=0 
M1716 diff_4667_6454# diff_4642_3644# diff_1660_6529# GND efet w=52 l=16
+ ad=1664 pd=192 as=0 ps=0 
M1717 GND diff_4604_6554# diff_4667_6454# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1718 diff_4784_6463# diff_4759_6532# GND GND efet w=55 l=16
+ ad=1517 pd=186 as=0 ps=0 
M1719 diff_1370_6508# diff_4861_3742# diff_4759_6532# GND efet w=17 l=17
+ ad=0 pd=0 as=1506 ps=182 
M1720 diff_1660_6529# diff_4771_3607# diff_4784_6463# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1721 diff_4667_6373# diff_4642_3644# diff_1663_6337# GND efet w=49 l=16
+ ad=1685 pd=192 as=0 ps=0 
M1722 diff_1370_6335# diff_4516_3742# diff_4414_6325# GND efet w=19 l=16
+ ad=0 pd=0 as=1512 ps=182 
M1723 diff_4607_6322# diff_4588_3644# diff_1370_6335# GND efet w=19 l=19
+ ad=1443 pd=188 as=0 ps=0 
M1724 diff_1370_6154# diff_4516_3742# diff_4414_6178# GND efet w=19 l=16
+ ad=0 pd=0 as=1512 ps=182 
M1725 diff_1660_6178# diff_4426_3610# diff_4439_6109# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1726 diff_4322_6019# diff_4300_3644# diff_1663_5983# GND efet w=49 l=16
+ ad=1649 pd=192 as=0 ps=0 
M1727 diff_1663_5983# diff_4426_3610# diff_4439_6004# GND efet w=52 l=19
+ ad=0 pd=0 as=1526 ps=186 
M1728 diff_1370_5981# diff_4171_3745# diff_4072_5968# GND efet w=19 l=16
+ ad=0 pd=0 as=1434 ps=188 
M1729 diff_4262_5968# diff_4243_3644# diff_1370_5981# GND efet w=19 l=16
+ ad=1470 pd=188 as=0 ps=0 
M1730 diff_1370_5800# diff_4171_3745# diff_4072_5821# GND efet w=19 l=16
+ ad=0 pd=0 as=1359 ps=182 
M1731 diff_1663_5821# diff_4084_3607# diff_4094_5755# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1732 diff_3980_5665# diff_3955_3644# diff_1663_5629# GND efet w=49 l=16
+ ad=1502 pd=186 as=0 ps=0 
M1733 GND diff_3917_5614# diff_3980_5665# GND efet w=62 l=17
+ ad=0 pd=0 as=0 ps=0 
M1734 diff_1370_5630# diff_3829_3644# diff_3727_5617# GND efet w=19 l=19
+ ad=0 pd=0 as=1422 ps=182 
M1735 diff_3917_5614# diff_3898_3644# diff_1370_5630# GND efet w=19 l=16
+ ad=1485 pd=182 as=0 ps=0 
M1736 diff_1370_5446# diff_3829_3644# diff_3727_5470# GND efet w=22 l=16
+ ad=0 pd=0 as=1425 ps=182 
M1737 diff_1663_5467# diff_3739_3610# diff_3752_5401# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1738 diff_3635_5311# diff_3610_3644# diff_1663_5275# GND efet w=52 l=16
+ ad=1652 pd=186 as=0 ps=0 
M1739 diff_1370_5273# diff_3484_3742# diff_3385_5260# GND efet w=19 l=16
+ ad=0 pd=0 as=1503 ps=182 
M1740 diff_3575_5263# diff_3556_3644# diff_1370_5273# GND efet w=22 l=16
+ ad=1494 pd=182 as=0 ps=0 
M1741 GND diff_3230_5122# diff_3293_5038# GND efet w=65 l=17
+ ad=0 pd=0 as=1526 ps=186 
M1742 diff_3293_5038# diff_3268_3644# diff_1663_5113# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1743 diff_3407_5047# diff_3385_5113# GND GND efet w=55 l=16
+ ad=1505 pd=180 as=0 ps=0 
M1744 diff_1370_5092# diff_3484_3742# diff_3385_5113# GND efet w=19 l=16
+ ad=0 pd=0 as=1521 ps=182 
M1745 diff_1663_5113# diff_3394_3613# diff_3407_5047# GND efet w=52 l=19
+ ad=0 pd=0 as=0 ps=0 
M1746 diff_3293_4954# diff_3268_3644# diff_1663_4918# GND efet w=52 l=17
+ ad=1526 pd=186 as=0 ps=0 
M1747 GND diff_3230_4906# diff_3293_4954# GND efet w=65 l=17
+ ad=0 pd=0 as=0 ps=0 
M1748 diff_1370_4919# diff_3142_3644# diff_3040_4906# GND efet w=19 l=16
+ ad=0 pd=0 as=1497 ps=188 
M1749 diff_3230_4906# diff_3211_3644# diff_1370_4919# GND efet w=19 l=16
+ ad=1533 pd=188 as=0 ps=0 
M1750 diff_2951_4681# diff_2923_3644# diff_1663_4756# GND efet w=52 l=19
+ ad=1568 pd=186 as=0 ps=0 
M1751 GND diff_2888_4765# diff_2951_4681# GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M1752 diff_3065_4690# diff_3040_4759# GND GND efet w=59 l=17
+ ad=1541 pd=186 as=0 ps=0 
M1753 diff_1370_4735# diff_3142_3644# diff_3040_4759# GND efet w=22 l=16
+ ad=0 pd=0 as=1560 ps=194 
M1754 diff_1663_4756# diff_3052_3607# diff_3065_4690# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1755 diff_2951_4597# diff_2923_3644# diff_1663_4564# GND efet w=53 l=20
+ ad=1520 pd=180 as=0 ps=0 
M1756 diff_1370_4565# diff_2797_3745# diff_2698_4549# GND efet w=19 l=16
+ ad=0 pd=0 as=1521 ps=182 
M1757 diff_2888_4552# diff_2869_3644# diff_1370_4565# GND efet w=19 l=16
+ ad=1485 pd=182 as=0 ps=0 
M1758 diff_2606_4327# diff_2581_3644# diff_1663_4402# GND efet w=52 l=16
+ ad=1526 pd=186 as=0 ps=0 
M1759 GND diff_2543_4411# diff_2606_4327# GND efet w=55 l=19
+ ad=0 pd=0 as=0 ps=0 
M1760 diff_2720_4336# diff_2698_4405# GND GND efet w=55 l=16
+ ad=1547 pd=186 as=0 ps=0 
M1761 diff_1370_4381# diff_2797_3745# diff_2698_4405# GND efet w=19 l=16
+ ad=0 pd=0 as=1530 ps=182 
M1762 diff_1663_4402# diff_2707_3610# diff_2720_4336# GND efet w=55 l=19
+ ad=0 pd=0 as=0 ps=0 
M1763 diff_2606_4243# diff_2581_3644# diff_1663_4210# GND efet w=52 l=17
+ ad=1574 pd=186 as=0 ps=0 
M1764 diff_1370_4211# diff_2455_3644# diff_2353_4195# GND efet w=19 l=16
+ ad=0 pd=0 as=1488 ps=188 
M1765 diff_2543_4195# diff_2524_3644# diff_1370_4211# GND efet w=20 l=16
+ ad=1509 pd=182 as=0 ps=0 
M1766 diff_1370_4027# diff_2455_3644# diff_2353_4051# GND efet w=19 l=16
+ ad=0 pd=0 as=1527 ps=194 
M1767 diff_1663_4051# diff_2365_3607# diff_2378_3982# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1768 diff_2264_3889# diff_2236_3644# diff_1663_3859# GND efet w=58 l=19
+ ad=1574 pd=186 as=0 ps=0 
M1769 diff_1370_3857# diff_2110_3745# diff_2011_3844# GND efet w=19 l=19
+ ad=0 pd=0 as=1512 ps=182 
M1770 diff_2201_3841# diff_2182_3644# diff_1370_3857# GND efet w=20 l=17
+ ad=1470 pd=176 as=0 ps=0 
M1771 GND diff_2201_3841# diff_2264_3889# GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M1772 diff_2378_3877# diff_2353_3844# GND GND efet w=59 l=17
+ ad=1550 pd=186 as=0 ps=0 
M1773 diff_1663_3859# diff_2365_3607# diff_2378_3877# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1774 diff_2546_4054# diff_2524_3644# diff_1370_4027# GND efet w=19 l=19
+ ad=1461 pd=188 as=0 ps=0 
M1775 GND diff_2543_4195# diff_2606_4243# GND efet w=58 l=19
+ ad=0 pd=0 as=0 ps=0 
M1776 diff_2720_4231# diff_2698_4195# GND GND efet w=58 l=16
+ ad=1574 pd=186 as=0 ps=0 
M1777 diff_1663_4210# diff_2707_3610# diff_2720_4231# GND efet w=53 l=20
+ ad=0 pd=0 as=0 ps=0 
M1778 diff_2888_4411# diff_2869_3644# diff_1370_4381# GND efet w=19 l=16
+ ad=1449 pd=182 as=0 ps=0 
M1779 diff_1370_4211# diff_2797_3745# diff_2698_4195# GND efet w=19 l=16
+ ad=0 pd=0 as=1512 ps=182 
M1780 GND diff_2888_4552# diff_2951_4597# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1781 diff_3065_4588# diff_3040_4549# GND GND efet w=59 l=17
+ ad=1496 pd=180 as=0 ps=0 
M1782 diff_1663_4564# diff_3052_3607# diff_3065_4588# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1783 diff_2951_4327# diff_2923_3644# diff_1663_4402# GND efet w=52 l=19
+ ad=1514 pd=180 as=0 ps=0 
M1784 GND diff_2888_4411# diff_2951_4327# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1785 diff_3065_4336# diff_3040_4405# GND GND efet w=65 l=17
+ ad=1517 pd=186 as=0 ps=0 
M1786 diff_3230_4762# diff_3211_3644# diff_1370_4735# GND efet w=22 l=16
+ ad=1569 pd=194 as=0 ps=0 
M1787 diff_3407_4942# diff_3385_4906# GND GND efet w=55 l=16
+ ad=1541 pd=180 as=0 ps=0 
M1788 diff_1663_4918# diff_3394_3613# diff_3407_4942# GND efet w=52 l=19
+ ad=0 pd=0 as=0 ps=0 
M1789 diff_3575_5122# diff_3556_3644# diff_1370_5092# GND efet w=19 l=16
+ ad=1476 pd=182 as=0 ps=0 
M1790 diff_1370_4919# diff_3484_3742# diff_3385_4906# GND efet w=22 l=16
+ ad=0 pd=0 as=1560 ps=194 
M1791 GND diff_3575_5263# diff_3635_5311# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1792 diff_3752_5299# diff_3727_5260# GND GND efet w=55 l=17
+ ad=1496 pd=180 as=0 ps=0 
M1793 diff_1663_5275# diff_3739_3610# diff_3752_5299# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1794 diff_3635_5038# diff_3610_3644# diff_1663_5113# GND efet w=52 l=16
+ ad=1661 pd=186 as=0 ps=0 
M1795 GND diff_3575_5122# diff_3635_5038# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1796 diff_3752_5047# diff_3727_5113# GND GND efet w=58 l=17
+ ad=1496 pd=180 as=0 ps=0 
M1797 diff_3917_5473# diff_3898_3644# diff_1370_5446# GND efet w=19 l=16
+ ad=1512 pd=182 as=0 ps=0 
M1798 diff_1370_5273# diff_3829_3644# diff_3727_5260# GND efet w=16 l=16
+ ad=0 pd=0 as=1527 ps=188 
M1799 diff_4094_5650# diff_4072_5614# GND GND efet w=55 l=16
+ ad=1517 pd=186 as=0 ps=0 
M1800 diff_1663_5629# diff_4084_3607# diff_4094_5650# GND efet w=50 l=17
+ ad=0 pd=0 as=0 ps=0 
M1801 diff_4262_5827# diff_4243_3644# diff_1370_5800# GND efet w=19 l=16
+ ad=1356 pd=176 as=0 ps=0 
M1802 GND diff_4262_5968# diff_4322_6019# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1803 diff_4439_6004# diff_4414_5971# GND GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1804 diff_4322_5746# diff_4300_3644# diff_1663_5821# GND efet w=55 l=16
+ ad=1649 pd=192 as=0 ps=0 
M1805 GND diff_4262_5827# diff_4322_5746# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1806 diff_4439_5755# diff_4414_5824# GND GND efet w=55 l=16
+ ad=1523 pd=180 as=0 ps=0 
M1807 diff_4604_6181# diff_4588_3644# diff_1370_6154# GND efet w=20 l=17
+ ad=1422 pd=206 as=0 ps=0 
M1808 GND diff_4607_6322# diff_4667_6373# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1809 diff_4784_6358# diff_4759_6325# GND GND efet w=55 l=16
+ ad=1529 pd=186 as=0 ps=0 
M1810 diff_1663_6337# diff_4771_3607# diff_4784_6358# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M1811 diff_4667_6100# diff_4642_3644# diff_1660_6178# GND efet w=52 l=16
+ ad=1673 pd=192 as=0 ps=0 
M1812 GND diff_4604_6181# diff_4667_6100# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1813 diff_4784_6109# diff_4759_6178# GND GND efet w=56 l=17
+ ad=1505 pd=180 as=0 ps=0 
M1814 diff_4949_6538# diff_4933_3644# diff_1370_6508# GND efet w=19 l=16
+ ad=1482 pd=194 as=0 ps=0 
M1815 diff_5012_6454# diff_4987_3652# diff_1660_6529# GND efet w=52 l=16
+ ad=1655 pd=192 as=0 ps=0 
M1816 GND diff_4949_6538# diff_5012_6454# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1817 diff_5129_6463# diff_5104_6532# GND GND efet w=61 l=16
+ ad=1487 pd=180 as=0 ps=0 
M1818 diff_1370_6508# diff_5206_3742# diff_5104_6532# GND efet w=16 l=16
+ ad=0 pd=0 as=1461 ps=182 
M1819 diff_1660_6529# diff_5116_3613# diff_5129_6463# GND efet w=50 l=17
+ ad=0 pd=0 as=0 ps=0 
M1820 diff_5012_6373# diff_4987_3652# diff_1663_6337# GND efet w=49 l=16
+ ad=1649 pd=192 as=0 ps=0 
M1821 diff_5294_6538# diff_5278_3644# diff_1370_6508# GND efet w=16 l=16
+ ad=1437 pd=188 as=0 ps=0 
M1822 diff_1370_6335# diff_4861_3742# diff_4759_6325# GND efet w=19 l=16
+ ad=0 pd=0 as=1485 ps=182 
M1823 diff_4949_6322# diff_4933_3644# diff_1370_6335# GND efet w=19 l=16
+ ad=1461 pd=188 as=0 ps=0 
M1824 diff_1370_6154# diff_4861_3742# diff_4759_6178# GND efet w=19 l=16
+ ad=0 pd=0 as=1455 ps=194 
M1825 diff_1660_6178# diff_4771_3607# diff_4784_6109# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1826 diff_1663_5983# diff_4771_3607# diff_4784_6004# GND efet w=52 l=19
+ ad=0 pd=0 as=1505 ps=186 
M1827 diff_4667_6019# diff_4642_3644# diff_1663_5983# GND efet w=49 l=16
+ ad=1631 pd=192 as=0 ps=0 
M1828 GND diff_4604_5972# diff_4667_6019# GND efet w=56 l=20
+ ad=0 pd=0 as=0 ps=0 
M1829 diff_4784_6004# diff_4759_5968# GND GND efet w=58 l=19
+ ad=0 pd=0 as=0 ps=0 
M1830 diff_1370_5981# diff_4516_3742# diff_4414_5971# GND efet w=19 l=16
+ ad=0 pd=0 as=1569 ps=188 
M1831 diff_4604_5972# diff_4588_3644# diff_1370_5981# GND efet w=25 l=17
+ ad=1473 pd=200 as=0 ps=0 
M1832 diff_1370_5800# diff_4516_3742# diff_4414_5824# GND efet w=19 l=16
+ ad=0 pd=0 as=1443 ps=188 
M1833 diff_4604_5834# diff_4588_3644# diff_1370_5800# GND efet w=22 l=16
+ ad=1446 pd=188 as=0 ps=0 
M1834 diff_1663_5821# diff_4426_3610# diff_4439_5755# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1835 diff_4322_5665# diff_4300_3644# diff_1663_5629# GND efet w=52 l=16
+ ad=1601 pd=198 as=0 ps=0 
M1836 diff_1370_5630# diff_4171_3745# diff_4072_5614# GND efet w=19 l=16
+ ad=0 pd=0 as=1434 ps=188 
M1837 diff_4262_5614# diff_4243_3644# diff_1370_5630# GND efet w=19 l=16
+ ad=1506 pd=188 as=0 ps=0 
M1838 diff_1370_5446# diff_4171_3745# diff_4072_5470# GND efet w=19 l=16
+ ad=0 pd=0 as=1422 ps=182 
M1839 diff_3980_5392# diff_3955_3644# diff_1663_5467# GND efet w=52 l=16
+ ad=1505 pd=180 as=0 ps=0 
M1840 GND diff_3917_5473# diff_3980_5392# GND efet w=59 l=17
+ ad=0 pd=0 as=0 ps=0 
M1841 diff_4094_5401# diff_4072_5470# GND GND efet w=55 l=16
+ ad=1508 pd=186 as=0 ps=0 
M1842 diff_1663_5467# diff_4084_3607# diff_4094_5401# GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M1843 diff_3980_5311# diff_3955_3644# diff_1663_5275# GND efet w=52 l=16
+ ad=1523 pd=180 as=0 ps=0 
M1844 diff_1663_5275# diff_4084_3607# diff_4094_5299# GND efet w=58 l=16
+ ad=0 pd=0 as=1592 ps=192 
M1845 diff_3917_5263# diff_3898_3644# diff_1370_5273# GND efet w=16 l=16
+ ad=1515 pd=182 as=0 ps=0 
M1846 diff_1370_5092# diff_3829_3644# diff_3727_5113# GND efet w=22 l=16
+ ad=0 pd=0 as=1536 ps=182 
M1847 diff_1663_5113# diff_3739_3610# diff_3752_5047# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1848 diff_3635_4954# diff_3610_3644# diff_1663_4918# GND efet w=50 l=17
+ ad=1670 pd=186 as=0 ps=0 
M1849 diff_3575_4906# diff_3556_3644# diff_1370_4919# GND efet w=19 l=16
+ ad=1560 pd=188 as=0 ps=0 
M1850 diff_3293_4681# diff_3268_3644# diff_1663_4756# GND efet w=52 l=16
+ ad=1433 pd=186 as=0 ps=0 
M1851 GND diff_3230_4762# diff_3293_4681# GND efet w=59 l=17
+ ad=0 pd=0 as=0 ps=0 
M1852 diff_3407_4690# diff_3385_4759# GND GND efet w=58 l=16
+ ad=1577 pd=186 as=0 ps=0 
M1853 diff_1370_4735# diff_3484_3742# diff_3385_4759# GND efet w=22 l=16
+ ad=0 pd=0 as=1536 ps=182 
M1854 diff_1663_4756# diff_3394_3613# diff_3407_4690# GND efet w=52 l=19
+ ad=0 pd=0 as=0 ps=0 
M1855 diff_3293_4600# diff_3268_3644# diff_1663_4564# GND efet w=52 l=16
+ ad=1523 pd=180 as=0 ps=0 
M1856 GND diff_3230_4552# diff_3293_4600# GND efet w=56 l=17
+ ad=0 pd=0 as=0 ps=0 
M1857 diff_1370_4565# diff_3142_3644# diff_3040_4549# GND efet w=19 l=16
+ ad=0 pd=0 as=1509 ps=194 
M1858 diff_3230_4552# diff_3211_3644# diff_1370_4565# GND efet w=19 l=16
+ ad=1458 pd=182 as=0 ps=0 
M1859 diff_1370_4381# diff_3142_3644# diff_3040_4405# GND efet w=20 l=16
+ ad=0 pd=0 as=1479 ps=194 
M1860 diff_3230_4411# diff_3211_3644# diff_1370_4381# GND efet w=19 l=16
+ ad=1359 pd=182 as=0 ps=0 
M1861 diff_1663_4402# diff_3052_3607# diff_3065_4336# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1862 diff_2951_4243# diff_2923_3644# diff_1663_4210# GND efet w=52 l=22
+ ad=1532 pd=180 as=0 ps=0 
M1863 GND diff_2888_4195# diff_2951_4243# GND efet w=56 l=20
+ ad=0 pd=0 as=0 ps=0 
M1864 diff_2888_4195# diff_2869_3644# diff_1370_4211# GND efet w=19 l=16
+ ad=1485 pd=182 as=0 ps=0 
M1865 diff_2606_3973# diff_2581_3644# diff_1663_4051# GND efet w=52 l=16
+ ad=1514 pd=180 as=0 ps=0 
M1866 GND diff_2546_4054# diff_2606_3973# GND efet w=55 l=19
+ ad=0 pd=0 as=0 ps=0 
M1867 diff_2720_3982# diff_2698_4051# GND GND efet w=55 l=16
+ ad=1505 pd=180 as=0 ps=0 
M1868 diff_1370_4027# diff_2797_3745# diff_2698_4051# GND efet w=19 l=16
+ ad=0 pd=0 as=1521 ps=182 
M1869 diff_1663_4051# diff_2707_3610# diff_2720_3982# GND efet w=52 l=19
+ ad=0 pd=0 as=0 ps=0 
M1870 diff_2888_4054# diff_2869_3644# diff_1370_4027# GND efet w=19 l=16
+ ad=1455 pd=176 as=0 ps=0 
M1871 diff_2606_3892# diff_2581_3644# diff_1663_3859# GND efet w=52 l=16
+ ad=1559 pd=186 as=0 ps=0 
M1872 diff_1370_3857# diff_2455_3644# diff_2353_3844# GND efet w=22 l=19
+ ad=0 pd=0 as=1542 ps=194 
M1873 diff_2546_3841# diff_2524_3644# diff_1370_3857# GND efet w=20 l=20
+ ad=1473 pd=182 as=0 ps=0 
M1874 GND diff_2546_3841# diff_2606_3892# GND efet w=58 l=19
+ ad=0 pd=0 as=0 ps=0 
M1875 diff_2720_3877# diff_2698_3844# GND GND efet w=58 l=16
+ ad=1607 pd=198 as=0 ps=0 
M1876 diff_1663_3859# diff_2707_3610# diff_2720_3877# GND efet w=58 l=19
+ ad=0 pd=0 as=0 ps=0 
M1877 diff_3065_4231# diff_3040_4195# GND GND efet w=58 l=22
+ ad=1535 pd=186 as=0 ps=0 
M1878 diff_1663_4210# diff_3052_3607# diff_3065_4231# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M1879 diff_2951_3973# diff_2923_3644# diff_1663_4051# GND efet w=52 l=19
+ ad=1505 pd=180 as=0 ps=0 
M1880 GND diff_2888_4054# diff_2951_3973# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1881 diff_3065_3982# diff_3040_4051# GND GND efet w=55 l=17
+ ad=1505 pd=180 as=0 ps=0 
M1882 diff_1370_4211# diff_3142_3644# diff_3040_4195# GND efet w=22 l=19
+ ad=0 pd=0 as=1476 ps=194 
M1883 diff_3407_4588# diff_3385_4549# GND GND efet w=55 l=16
+ ad=1514 pd=180 as=0 ps=0 
M1884 diff_1663_4564# diff_3394_3613# diff_3407_4588# GND efet w=52 l=19
+ ad=0 pd=0 as=0 ps=0 
M1885 diff_3575_4762# diff_3556_3644# diff_1370_4735# GND efet w=22 l=16
+ ad=1485 pd=188 as=0 ps=0 
M1886 GND diff_3575_4906# diff_3635_4954# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1887 diff_3752_4942# diff_3727_4906# GND GND efet w=55 l=17
+ ad=1499 pd=180 as=0 ps=0 
M1888 diff_1663_4918# diff_3739_3610# diff_3752_4942# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M1889 diff_3635_4681# diff_3610_3644# diff_1663_4756# GND efet w=52 l=16
+ ad=1733 pd=192 as=0 ps=0 
M1890 GND diff_3575_4762# diff_3635_4681# GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M1891 diff_3752_4690# diff_3727_4759# GND GND efet w=59 l=17
+ ad=1550 pd=186 as=0 ps=0 
M1892 diff_3917_5119# diff_3898_3644# diff_1370_5092# GND efet w=19 l=16
+ ad=1521 pd=182 as=0 ps=0 
M1893 GND diff_3917_5263# diff_3980_5311# GND efet w=55 l=17
+ ad=0 pd=0 as=0 ps=0 
M1894 diff_4094_5299# diff_4072_5260# GND GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1895 GND diff_3917_5119# diff_3980_5038# GND efet w=58 l=17
+ ad=0 pd=0 as=1517 ps=186 
M1896 diff_3980_5038# diff_3955_3644# diff_1663_5113# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1897 diff_4094_5047# diff_4072_5113# GND GND efet w=55 l=16
+ ad=1673 pd=192 as=0 ps=0 
M1898 diff_4262_5473# diff_4243_3644# diff_1370_5446# GND efet w=19 l=16
+ ad=1440 pd=182 as=0 ps=0 
M1899 diff_1370_5273# diff_4171_3745# diff_4072_5260# GND efet w=17 l=17
+ ad=0 pd=0 as=1440 ps=182 
M1900 GND diff_4262_5614# diff_4322_5665# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1901 diff_4439_5650# diff_4414_5617# GND GND efet w=55 l=16
+ ad=1508 pd=180 as=0 ps=0 
M1902 diff_1663_5629# diff_4426_3610# diff_4439_5650# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M1903 diff_4322_5396# diff_4300_3644# diff_1663_5467# GND efet w=55 l=17
+ ad=1541 pd=192 as=0 ps=0 
M1904 GND diff_4262_5473# diff_4322_5396# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1905 diff_4439_5401# diff_4414_5473# GND GND efet w=55 l=16
+ ad=1514 pd=180 as=0 ps=0 
M1906 diff_4667_5746# diff_4642_3644# diff_1663_5821# GND efet w=52 l=16
+ ad=1673 pd=192 as=0 ps=0 
M1907 GND diff_4604_5834# diff_4667_5746# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1908 diff_4784_5755# diff_4759_5824# GND GND efet w=58 l=16
+ ad=1505 pd=180 as=0 ps=0 
M1909 diff_4949_6181# diff_4933_3644# diff_1370_6154# GND efet w=19 l=16
+ ad=1470 pd=188 as=0 ps=0 
M1910 GND diff_4949_6322# diff_5012_6373# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1911 diff_5129_6358# diff_5104_6322# GND GND efet w=59 l=17
+ ad=1520 pd=186 as=0 ps=0 
M1912 diff_1663_6337# diff_5116_3613# diff_5129_6358# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M1913 diff_5012_6100# diff_4987_3652# diff_1660_6178# GND efet w=52 l=16
+ ad=1655 pd=192 as=0 ps=0 
M1914 GND diff_4949_6181# diff_5012_6100# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1915 diff_5126_6140# diff_5104_6178# GND GND efet w=61 l=17
+ ad=1517 pd=192 as=0 ps=0 
M1916 Vdd diff_4732_1658# diff_1370_6508# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M1917 diff_5357_6454# diff_5335_3644# diff_1660_6529# GND efet w=52 l=16
+ ad=1715 pd=192 as=0 ps=0 
M1918 GND diff_5294_6538# diff_5357_6454# GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M1919 Vdd diff_5563_3961# diff_1660_6529# GND efet w=34 l=14
+ ad=0 pd=0 as=0 ps=0 
M1920 diff_6040_7132# Vdd Vdd GND efet w=25 l=46
+ ad=0 pd=0 as=0 ps=0 
M1921 Vdd Vdd Vdd GND efet w=10 l=6
+ ad=0 pd=0 as=0 ps=0 
M1922 Vdd Vdd Vdd GND efet w=8 l=17
+ ad=0 pd=0 as=0 ps=0 
M1923 diff_6035_6505# Vdd Vdd GND efet w=31 l=44
+ ad=7827 pd=646 as=0 ps=0 
M1924 diff_5813_6445# clk2 diff_577_5317# GND efet w=46 l=16
+ ad=1706 pd=192 as=0 ps=0 
M1925 diff_5861_6427# diff_5188_6931# diff_5813_6445# GND efet w=46 l=16
+ ad=9929 pd=812 as=0 ps=0 
M1926 diff_5357_6373# diff_5335_3644# diff_1663_6337# GND efet w=49 l=16
+ ad=1334 pd=162 as=0 ps=0 
M1927 GND diff_5294_6322# diff_5357_6373# GND efet w=40 l=16
+ ad=0 pd=0 as=0 ps=0 
M1928 diff_1370_6335# diff_5206_3742# diff_5104_6322# GND efet w=19 l=19
+ ad=0 pd=0 as=1467 ps=182 
M1929 diff_5294_6322# diff_5278_3644# diff_1370_6335# GND efet w=19 l=16
+ ad=1461 pd=188 as=0 ps=0 
M1930 diff_1370_6154# diff_5206_3742# diff_5104_6178# GND efet w=17 l=20
+ ad=0 pd=0 as=1334 ps=220 
M1931 diff_5294_6181# diff_5278_3644# diff_1370_6154# GND efet w=19 l=19
+ ad=1440 pd=182 as=0 ps=0 
M1932 diff_1660_6178# diff_5116_3613# diff_5126_6140# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1933 diff_5012_6019# diff_4987_3652# diff_1663_5983# GND efet w=50 l=17
+ ad=1589 pd=192 as=0 ps=0 
M1934 diff_1370_5981# diff_4861_3742# diff_4759_5968# GND efet w=19 l=16
+ ad=0 pd=0 as=1503 ps=182 
M1935 diff_4949_5968# diff_4933_3644# diff_1370_5981# GND efet w=19 l=16
+ ad=1488 pd=188 as=0 ps=0 
M1936 diff_1370_5800# diff_4861_3742# diff_4759_5824# GND efet w=20 l=17
+ ad=0 pd=0 as=1536 ps=182 
M1937 diff_1663_5821# diff_4771_3607# diff_4784_5755# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1938 diff_4667_5665# diff_4642_3644# diff_1663_5629# GND efet w=49 l=16
+ ad=1646 pd=186 as=0 ps=0 
M1939 diff_1370_5630# diff_4516_3742# diff_4414_5617# GND efet w=19 l=16
+ ad=0 pd=0 as=1488 ps=188 
M1940 diff_4604_5627# diff_4588_3644# diff_1370_5630# GND efet w=23 l=16
+ ad=1461 pd=194 as=0 ps=0 
M1941 diff_1370_5446# diff_4516_3742# diff_4414_5473# GND efet w=19 l=16
+ ad=0 pd=0 as=1512 ps=182 
M1942 diff_1663_5467# diff_4426_3610# diff_4439_5401# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1943 diff_4325_5311# diff_4300_3644# diff_1663_5275# GND efet w=52 l=19
+ ad=1559 pd=186 as=0 ps=0 
M1944 diff_4262_5260# diff_4243_3644# diff_1370_5273# GND efet w=19 l=19
+ ad=1449 pd=182 as=0 ps=0 
M1945 GND diff_4262_5260# diff_4325_5311# GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M1946 diff_4439_5296# diff_4414_5275# GND GND efet w=58 l=16
+ ad=1541 pd=186 as=0 ps=0 
M1947 diff_1663_5275# diff_4426_3610# diff_4439_5296# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1948 diff_4262_5119# diff_4243_3644# diff_1370_5092# GND efet w=22 l=19
+ ad=1437 pd=182 as=0 ps=0 
M1949 diff_1370_5092# diff_4171_3745# diff_4072_5113# GND efet w=19 l=16
+ ad=0 pd=0 as=1440 ps=182 
M1950 diff_1663_5113# diff_4084_3607# diff_4094_5047# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1951 diff_3980_4957# diff_3955_3644# diff_1663_4918# GND efet w=49 l=16
+ ad=1499 pd=180 as=0 ps=0 
M1952 diff_1370_4919# diff_3829_3644# diff_3727_4906# GND efet w=19 l=16
+ ad=0 pd=0 as=1476 ps=182 
M1953 diff_3917_4906# diff_3898_3644# diff_1370_4919# GND efet w=19 l=16
+ ad=1473 pd=194 as=0 ps=0 
M1954 diff_1370_4735# diff_3829_3644# diff_3727_4759# GND efet w=20 l=17
+ ad=0 pd=0 as=1530 ps=182 
M1955 diff_3917_4762# diff_3898_3644# diff_1370_4735# GND efet w=22 l=16
+ ad=1542 pd=194 as=0 ps=0 
M1956 diff_1663_4756# diff_3739_3610# diff_3752_4690# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1957 diff_3635_4600# diff_3610_3644# diff_1663_4564# GND efet w=52 l=16
+ ad=1670 pd=186 as=0 ps=0 
M1958 diff_1370_4565# diff_3484_3742# diff_3385_4549# GND efet w=19 l=16
+ ad=0 pd=0 as=1512 ps=182 
M1959 diff_3575_4552# diff_3556_3644# diff_1370_4565# GND efet w=19 l=16
+ ad=1494 pd=182 as=0 ps=0 
M1960 GND diff_3230_4411# diff_3293_4327# GND efet w=62 l=17
+ ad=0 pd=0 as=1526 ps=186 
M1961 diff_3293_4327# diff_3268_3644# diff_1663_4402# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1962 diff_3407_4336# diff_3385_4402# GND GND efet w=55 l=16
+ ad=1505 pd=180 as=0 ps=0 
M1963 diff_1370_4381# diff_3484_3742# diff_3385_4402# GND efet w=19 l=16
+ ad=0 pd=0 as=1503 ps=182 
M1964 diff_1663_4402# diff_3394_3613# diff_3407_4336# GND efet w=52 l=19
+ ad=0 pd=0 as=0 ps=0 
M1965 diff_3293_4246# diff_3268_3644# diff_1663_4210# GND efet w=49 l=16
+ ad=1520 pd=186 as=0 ps=0 
M1966 diff_3230_4195# diff_3211_3644# diff_1370_4211# GND efet w=19 l=16
+ ad=1479 pd=188 as=0 ps=0 
M1967 diff_1370_4027# diff_3142_3644# diff_3040_4051# GND efet w=23 l=17
+ ad=0 pd=0 as=1470 ps=206 
M1968 diff_1663_4051# diff_3052_3607# diff_3065_3982# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1969 diff_3230_4054# diff_3211_3644# diff_1370_4027# GND efet w=19 l=16
+ ad=1419 pd=194 as=0 ps=0 
M1970 diff_2951_3892# diff_2923_3644# diff_1663_3859# GND efet w=52 l=19
+ ad=1550 pd=186 as=0 ps=0 
M1971 diff_1370_3857# diff_2797_3745# diff_2698_3844# GND efet w=20 l=17
+ ad=0 pd=0 as=1545 ps=182 
M1972 diff_2888_3841# diff_2869_3644# diff_1370_3857# GND efet w=22 l=16
+ ad=1470 pd=176 as=0 ps=0 
M1973 GND diff_2888_3841# diff_2951_3892# GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M1974 diff_3065_3877# diff_3040_3844# GND GND efet w=62 l=17
+ ad=1517 pd=192 as=0 ps=0 
M1975 diff_1663_3859# diff_3052_3607# diff_3065_3877# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1976 GND diff_3230_4195# diff_3293_4246# GND efet w=56 l=17
+ ad=0 pd=0 as=0 ps=0 
M1977 diff_3407_4231# diff_3385_4195# GND GND efet w=55 l=16
+ ad=1517 pd=180 as=0 ps=0 
M1978 diff_1663_4210# diff_3394_3613# diff_3407_4231# GND efet w=49 l=19
+ ad=0 pd=0 as=0 ps=0 
M1979 diff_3293_3973# diff_3268_3644# diff_1663_4051# GND efet w=52 l=16
+ ad=1514 pd=180 as=0 ps=0 
M1980 GND diff_3230_4054# diff_3293_3973# GND efet w=58 l=17
+ ad=0 pd=0 as=0 ps=0 
M1981 diff_3407_3982# diff_3385_4051# GND GND efet w=55 l=16
+ ad=1496 pd=180 as=0 ps=0 
M1982 diff_3575_4411# diff_3556_3644# diff_1370_4381# GND efet w=19 l=16
+ ad=1422 pd=182 as=0 ps=0 
M1983 GND diff_3575_4552# diff_3635_4600# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1984 diff_3752_4588# diff_3727_4549# GND GND efet w=61 l=17
+ ad=1490 pd=186 as=0 ps=0 
M1985 diff_1663_4564# diff_3739_3610# diff_3752_4588# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1986 diff_3635_4327# diff_3610_3644# diff_1663_4402# GND efet w=55 l=16
+ ad=1658 pd=192 as=0 ps=0 
M1987 GND diff_3575_4411# diff_3635_4327# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1988 diff_3752_4336# diff_3727_4405# GND GND efet w=55 l=19
+ ad=1496 pd=180 as=0 ps=0 
M1989 GND diff_3917_4906# diff_3980_4957# GND efet w=55 l=19
+ ad=0 pd=0 as=0 ps=0 
M1990 diff_4094_4942# diff_4072_4906# GND GND efet w=55 l=16
+ ad=1634 pd=192 as=0 ps=0 
M1991 diff_1663_4918# diff_4084_3607# diff_4094_4942# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M1992 diff_3980_4681# diff_3955_3644# diff_1663_4756# GND efet w=52 l=16
+ ad=1577 pd=186 as=0 ps=0 
M1993 GND diff_3917_4762# diff_3980_4681# GND efet w=58 l=19
+ ad=0 pd=0 as=0 ps=0 
M1994 diff_4094_4690# diff_4072_4759# GND GND efet w=58 l=16
+ ad=1721 pd=198 as=0 ps=0 
M1995 diff_1370_4919# diff_4171_3745# diff_4072_4906# GND efet w=19 l=16
+ ad=0 pd=0 as=1359 ps=182 
M1996 diff_4325_5038# diff_4300_3644# diff_1663_5113# GND efet w=52 l=19
+ ad=1406 pd=180 as=0 ps=0 
M1997 GND diff_4262_5119# diff_4325_5038# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M1998 diff_4439_5047# diff_4417_5113# GND GND efet w=55 l=16
+ ad=1517 pd=186 as=0 ps=0 
M1999 diff_4607_5473# diff_4588_3644# diff_1370_5446# GND efet w=19 l=19
+ ad=1452 pd=188 as=0 ps=0 
M2000 GND diff_4604_5627# diff_4667_5665# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2001 diff_4784_5650# diff_4759_5617# GND GND efet w=65 l=17
+ ad=1526 pd=180 as=0 ps=0 
M2002 diff_1663_5629# diff_4771_3607# diff_4784_5650# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M2003 diff_4667_5392# diff_4642_3644# diff_1663_5467# GND efet w=52 l=16
+ ad=1637 pd=192 as=0 ps=0 
M2004 GND diff_4607_5473# diff_4667_5392# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2005 diff_4784_5401# diff_4759_5470# GND GND efet w=61 l=16
+ ad=1487 pd=180 as=0 ps=0 
M2006 diff_4949_5827# diff_4933_3644# diff_1370_5800# GND efet w=19 l=16
+ ad=1488 pd=188 as=0 ps=0 
M2007 GND diff_4949_5968# diff_5012_6019# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2008 diff_5129_6007# diff_5104_5968# GND GND efet w=53 l=17
+ ad=1427 pd=174 as=0 ps=0 
M2009 diff_1663_5983# diff_5116_3613# diff_5129_6007# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M2010 diff_5012_5746# diff_4987_3652# diff_1663_5821# GND efet w=52 l=16
+ ad=1664 pd=192 as=0 ps=0 
M2011 GND diff_4949_5827# diff_5012_5746# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2012 diff_5129_5755# diff_5104_5824# GND GND efet w=65 l=17
+ ad=1487 pd=180 as=0 ps=0 
M2013 Vdd diff_5563_3961# diff_1663_6337# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M2014 Vdd diff_4732_1658# diff_1370_6335# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M2015 GND diff_5188_6931# diff_6059_6298# GND efet w=37 l=13
+ ad=0 pd=0 as=2327 ps=210 
M2016 GND diff_5194_7252# diff_5861_6427# GND efet w=68 l=14
+ ad=0 pd=0 as=0 ps=0 
M2017 diff_6059_6298# Vdd Vdd GND efet w=19 l=142
+ ad=0 pd=0 as=0 ps=0 
M2018 Vdd Vdd Vdd GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M2019 diff_5861_6427# diff_6059_6298# diff_6137_6238# GND efet w=34 l=16
+ ad=0 pd=0 as=3877 ps=352 
M2020 diff_6035_6505# diff_5861_6427# GND GND efet w=278 l=14
+ ad=0 pd=0 as=0 ps=0 
M2021 Vdd Vdd Vdd GND efet w=8 l=20
+ ad=0 pd=0 as=0 ps=0 
M2022 diff_6137_6238# Vdd Vdd GND efet w=25 l=68
+ ad=0 pd=0 as=0 ps=0 
M2023 Vdd diff_4732_1658# diff_1370_6154# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M2024 diff_5357_6100# diff_5335_3644# diff_1660_6178# GND efet w=52 l=16
+ ad=1661 pd=186 as=0 ps=0 
M2025 GND diff_5294_6181# diff_5357_6100# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2026 Vdd diff_5563_3961# diff_1660_6178# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M2027 o2 diff_5938_6088# Vdd GND efet w=515 l=14
+ ad=24765 pd=1738 as=0 ps=0 
M2028 diff_5357_6019# diff_5335_3644# diff_1663_5983# GND efet w=52 l=16
+ ad=1646 pd=192 as=0 ps=0 
M2029 diff_1370_5981# diff_5206_3742# diff_5104_5968# GND efet w=19 l=16
+ ad=0 pd=0 as=1494 ps=182 
M2030 diff_5294_5968# diff_5278_3644# diff_1370_5981# GND efet w=19 l=16
+ ad=1470 pd=188 as=0 ps=0 
M2031 diff_1370_5800# diff_5206_3742# diff_5104_5824# GND efet w=19 l=16
+ ad=0 pd=0 as=1503 ps=182 
M2032 diff_1663_5821# diff_5116_3613# diff_5129_5755# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2033 diff_5294_5827# diff_5278_3644# diff_1370_5800# GND efet w=19 l=16
+ ad=1470 pd=188 as=0 ps=0 
M2034 diff_5012_5665# diff_4987_3652# diff_1663_5629# GND efet w=49 l=16
+ ad=1649 pd=192 as=0 ps=0 
M2035 diff_1370_5630# diff_4861_3742# diff_4759_5617# GND efet w=19 l=16
+ ad=0 pd=0 as=1515 ps=188 
M2036 diff_4949_5614# diff_4933_3644# diff_1370_5630# GND efet w=19 l=16
+ ad=1461 pd=188 as=0 ps=0 
M2037 diff_1370_5446# diff_4861_3742# diff_4759_5470# GND efet w=19 l=16
+ ad=0 pd=0 as=1503 ps=182 
M2038 diff_4949_5476# diff_4933_3644# diff_1370_5446# GND efet w=16 l=16
+ ad=1473 pd=188 as=0 ps=0 
M2039 diff_1663_5467# diff_4771_3607# diff_4784_5401# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2040 diff_4667_5311# diff_4642_3644# diff_1663_5275# GND efet w=52 l=16
+ ad=1661 pd=186 as=0 ps=0 
M2041 diff_1370_5273# diff_4516_3742# diff_4414_5275# GND efet w=19 l=16
+ ad=0 pd=0 as=1500 ps=194 
M2042 diff_4607_5263# diff_4588_3644# diff_1370_5273# GND efet w=20 l=19
+ ad=1479 pd=188 as=0 ps=0 
M2043 diff_1370_5092# diff_4516_3742# diff_4417_5113# GND efet w=22 l=16
+ ad=0 pd=0 as=1548 ps=188 
M2044 diff_1663_5113# diff_4426_3610# diff_4439_5047# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2045 diff_4325_4954# diff_4300_3644# diff_1663_4918# GND efet w=50 l=20
+ ad=1517 pd=186 as=0 ps=0 
M2046 diff_4262_4906# diff_4243_3644# diff_1370_4919# GND efet w=19 l=16
+ ad=1350 pd=182 as=0 ps=0 
M2047 diff_1370_4735# diff_4171_3745# diff_4072_4759# GND efet w=19 l=16
+ ad=0 pd=0 as=1431 ps=182 
M2048 diff_1663_4756# diff_4084_3607# diff_4094_4690# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2049 diff_3980_4600# diff_3955_3644# diff_1663_4564# GND efet w=52 l=16
+ ad=1541 pd=186 as=0 ps=0 
M2050 diff_1663_4564# diff_4084_3607# diff_4094_4585# GND efet w=65 l=16
+ ad=0 pd=0 as=1664 ps=216 
M2051 diff_1370_4565# diff_3829_3644# diff_3727_4549# GND efet w=20 l=17
+ ad=0 pd=0 as=1521 ps=182 
M2052 diff_3917_4549# diff_3898_3644# diff_1370_4565# GND efet w=22 l=19
+ ad=1527 pd=182 as=0 ps=0 
M2053 diff_1370_4381# diff_3829_3644# diff_3727_4405# GND efet w=19 l=16
+ ad=0 pd=0 as=1494 ps=182 
M2054 diff_1663_4402# diff_3739_3610# diff_3752_4336# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2055 diff_3635_4246# diff_3610_3644# diff_1663_4210# GND efet w=49 l=16
+ ad=1664 pd=186 as=0 ps=0 
M2056 diff_1370_4211# diff_3484_3742# diff_3385_4195# GND efet w=19 l=16
+ ad=0 pd=0 as=1533 ps=188 
M2057 diff_3575_4195# diff_3556_3644# diff_1370_4211# GND efet w=20 l=17
+ ad=1446 pd=176 as=0 ps=0 
M2058 diff_1370_4027# diff_3484_3742# diff_3385_4051# GND efet w=19 l=16
+ ad=0 pd=0 as=1512 ps=182 
M2059 diff_1663_4051# diff_3394_3613# diff_3407_3982# GND efet w=52 l=19
+ ad=0 pd=0 as=0 ps=0 
M2060 diff_3293_3892# diff_3268_3644# diff_1663_3859# GND efet w=52 l=16
+ ad=1508 pd=186 as=0 ps=0 
M2061 diff_1370_3857# diff_3142_3644# diff_3040_3844# GND efet w=19 l=16
+ ad=0 pd=0 as=1527 ps=194 
M2062 diff_3230_3844# diff_3211_3644# diff_1370_3857# GND efet w=19 l=16
+ ad=1461 pd=188 as=0 ps=0 
M2063 GND diff_3230_3844# diff_3293_3892# GND efet w=55 l=19
+ ad=0 pd=0 as=0 ps=0 
M2064 diff_3407_3880# diff_3385_3844# GND GND efet w=55 l=16
+ ad=1487 pd=180 as=0 ps=0 
M2065 diff_1663_3859# diff_3394_3613# diff_3407_3880# GND efet w=52 l=19
+ ad=0 pd=0 as=0 ps=0 
M2066 diff_3575_4054# diff_3556_3644# diff_1370_4027# GND efet w=19 l=16
+ ad=1446 pd=176 as=0 ps=0 
M2067 GND diff_3575_4195# diff_3635_4246# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2068 diff_3752_4231# diff_3727_4195# GND GND efet w=55 l=19
+ ad=1484 pd=186 as=0 ps=0 
M2069 diff_1663_4210# diff_3739_3610# diff_3752_4231# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M2070 diff_3635_3973# diff_3610_3644# diff_1663_4051# GND efet w=52 l=16
+ ad=1670 pd=186 as=0 ps=0 
M2071 GND diff_3575_4054# diff_3635_3973# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2072 diff_3752_3982# diff_3727_4051# GND GND efet w=55 l=19
+ ad=1496 pd=180 as=0 ps=0 
M2073 diff_3917_4411# diff_3898_3644# diff_1370_4381# GND efet w=19 l=16
+ ad=1512 pd=182 as=0 ps=0 
M2074 diff_1370_4211# diff_3829_3644# diff_3727_4195# GND efet w=19 l=16
+ ad=0 pd=0 as=1503 ps=182 
M2075 GND diff_3917_4549# diff_3980_4600# GND efet w=56 l=20
+ ad=0 pd=0 as=0 ps=0 
M2076 diff_4094_4585# diff_4072_4549# GND GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M2077 diff_4262_4765# diff_4243_3644# diff_1370_4735# GND efet w=19 l=16
+ ad=1509 pd=194 as=0 ps=0 
M2078 GND diff_4262_4906# diff_4325_4954# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2079 diff_4439_4942# diff_4417_4903# GND GND efet w=55 l=16
+ ad=1508 pd=186 as=0 ps=0 
M2080 diff_1663_4918# diff_4426_3610# diff_4439_4942# GND efet w=50 l=17
+ ad=0 pd=0 as=0 ps=0 
M2081 diff_4325_4681# diff_4300_3644# diff_1663_4756# GND efet w=52 l=19
+ ad=1568 pd=186 as=0 ps=0 
M2082 GND diff_4262_4765# diff_4325_4681# GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M2083 diff_4439_4690# diff_4414_4762# GND GND efet w=58 l=16
+ ad=1577 pd=186 as=0 ps=0 
M2084 diff_4607_5119# diff_4588_3644# diff_1370_5092# GND efet w=22 l=16
+ ad=1494 pd=188 as=0 ps=0 
M2085 GND diff_4607_5263# diff_4667_5311# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2086 diff_4784_5299# diff_4759_5260# GND GND efet w=55 l=16
+ ad=1505 pd=180 as=0 ps=0 
M2087 diff_1663_5275# diff_4771_3607# diff_4784_5299# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2088 diff_4667_5038# diff_4642_3644# diff_1663_5113# GND efet w=52 l=16
+ ad=1664 pd=192 as=0 ps=0 
M2089 GND diff_4607_5119# diff_4667_5038# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2090 diff_4784_5047# diff_4759_5113# GND GND efet w=55 l=16
+ ad=1505 pd=180 as=0 ps=0 
M2091 GND diff_4949_5614# diff_5012_5665# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2092 diff_5129_5650# diff_5104_5617# GND GND efet w=59 l=17
+ ad=1481 pd=180 as=0 ps=0 
M2093 diff_1663_5629# diff_5116_3613# diff_5129_5650# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M2094 diff_5012_5395# diff_4987_3652# diff_1663_5467# GND efet w=49 l=16
+ ad=1619 pd=186 as=0 ps=0 
M2095 GND diff_4949_5476# diff_5012_5395# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2096 diff_5129_5401# diff_5104_5470# GND GND efet w=55 l=17
+ ad=1442 pd=174 as=0 ps=0 
M2097 GND diff_5294_5968# diff_5357_6019# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2098 diff_6137_6238# diff_6035_6505# GND GND efet w=61 l=16
+ ad=0 pd=0 as=0 ps=0 
M2099 o2 diff_6035_6505# GND GND efet w=490 l=13
+ ad=0 pd=0 as=0 ps=0 
M2100 Vdd diff_5563_3961# diff_1663_5983# GND efet w=34 l=19
+ ad=0 pd=0 as=0 ps=0 
M2101 Vdd diff_4732_1658# diff_1370_5981# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M2102 diff_5938_6088# diff_5938_6088# diff_5938_6088# GND efet w=2 l=7
+ ad=6075 pd=412 as=0 ps=0 
M2103 diff_5938_6088# diff_5938_6088# diff_5938_6088# GND efet w=4 l=4
+ ad=0 pd=0 as=0 ps=0 
M2104 diff_5938_6088# Vdd Vdd GND efet w=25 l=46
+ ad=0 pd=0 as=0 ps=0 
M2105 diff_5938_6088# diff_6035_6505# GND GND efet w=122 l=14
+ ad=0 pd=0 as=0 ps=0 
M2106 Vdd diff_4732_1658# diff_1370_5800# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M2107 diff_5357_5746# diff_5335_3644# diff_1663_5821# GND efet w=52 l=16
+ ad=1664 pd=192 as=0 ps=0 
M2108 GND diff_5294_5827# diff_5357_5746# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2109 Vdd diff_5563_3961# diff_1663_5821# GND efet w=34 l=14
+ ad=0 pd=0 as=0 ps=0 
M2110 diff_5357_5665# diff_5335_3644# diff_1663_5629# GND efet w=49 l=16
+ ad=1589 pd=192 as=0 ps=0 
M2111 diff_1370_5630# diff_5206_3742# diff_5104_5617# GND efet w=19 l=16
+ ad=0 pd=0 as=1485 ps=182 
M2112 diff_5294_5614# diff_5278_3644# diff_1370_5630# GND efet w=19 l=16
+ ad=1467 pd=182 as=0 ps=0 
M2113 diff_1370_5446# diff_5206_3742# diff_5104_5470# GND efet w=16 l=16
+ ad=0 pd=0 as=1488 ps=182 
M2114 diff_1663_5467# diff_5116_3613# diff_5129_5401# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M2115 diff_5012_5311# diff_4987_3652# diff_1663_5275# GND efet w=52 l=16
+ ad=1652 pd=186 as=0 ps=0 
M2116 diff_1370_5273# diff_4861_3742# diff_4759_5260# GND efet w=16 l=16
+ ad=0 pd=0 as=1527 ps=188 
M2117 diff_4949_5263# diff_4933_3644# diff_1370_5273# GND efet w=16 l=16
+ ad=1494 pd=194 as=0 ps=0 
M2118 diff_1370_5092# diff_4861_3742# diff_4759_5113# GND efet w=22 l=16
+ ad=0 pd=0 as=1557 ps=188 
M2119 diff_4949_5122# diff_4933_3644# diff_1370_5092# GND efet w=19 l=16
+ ad=1467 pd=182 as=0 ps=0 
M2120 diff_1663_5113# diff_4771_3607# diff_4784_5047# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2121 diff_4667_4957# diff_4642_3644# diff_1663_4918# GND efet w=49 l=16
+ ad=1658 pd=192 as=0 ps=0 
M2122 diff_1370_4919# diff_4516_3742# diff_4417_4903# GND efet w=19 l=16
+ ad=0 pd=0 as=1458 ps=200 
M2123 diff_4607_4906# diff_4588_3644# diff_1370_4919# GND efet w=19 l=16
+ ad=1392 pd=194 as=0 ps=0 
M2124 diff_1370_4735# diff_4516_3742# diff_4414_4762# GND efet w=19 l=16
+ ad=0 pd=0 as=1437 ps=194 
M2125 diff_4607_4765# diff_4588_3644# diff_1370_4735# GND efet w=23 l=17
+ ad=1437 pd=194 as=0 ps=0 
M2126 diff_1663_4756# diff_4426_3610# diff_4439_4690# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2127 diff_4325_4600# diff_4300_3644# diff_1663_4564# GND efet w=52 l=19
+ ad=1550 pd=186 as=0 ps=0 
M2128 diff_1370_4565# diff_4171_3745# diff_4072_4549# GND efet w=22 l=16
+ ad=0 pd=0 as=1464 ps=182 
M2129 diff_4262_4549# diff_4243_3644# diff_1370_4565# GND efet w=22 l=16
+ ad=1476 pd=188 as=0 ps=0 
M2130 GND diff_4262_4549# diff_4325_4600# GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M2131 diff_4439_4585# diff_4414_4558# GND GND efet w=58 l=16
+ ad=1550 pd=186 as=0 ps=0 
M2132 diff_1663_4564# diff_4426_3610# diff_4439_4585# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2133 diff_1370_4381# diff_4171_3745# diff_4072_4402# GND efet w=16 l=17
+ ad=0 pd=0 as=1428 ps=188 
M2134 diff_4262_4411# diff_4243_3644# diff_1370_4381# GND efet w=17 l=17
+ ad=1452 pd=188 as=0 ps=0 
M2135 diff_3980_4327# diff_3955_3644# diff_1663_4402# GND efet w=52 l=16
+ ad=1517 pd=186 as=0 ps=0 
M2136 GND diff_3917_4411# diff_3980_4327# GND efet w=55 l=19
+ ad=0 pd=0 as=0 ps=0 
M2137 diff_4094_4336# diff_4072_4402# GND GND efet w=55 l=16
+ ad=1574 pd=204 as=0 ps=0 
M2138 diff_1663_4402# diff_4084_3607# diff_4094_4336# GND efet w=59 l=17
+ ad=0 pd=0 as=0 ps=0 
M2139 diff_3980_4246# diff_3955_3644# diff_1663_4210# GND efet w=49 l=16
+ ad=1499 pd=180 as=0 ps=0 
M2140 diff_3917_4195# diff_3898_3644# diff_1370_4211# GND efet w=19 l=16
+ ad=1521 pd=182 as=0 ps=0 
M2141 diff_1370_4027# diff_3829_3644# diff_3727_4051# GND efet w=19 l=19
+ ad=0 pd=0 as=1500 ps=194 
M2142 diff_1663_4051# diff_3739_3610# diff_3752_3982# GND efet w=50 l=19
+ ad=0 pd=0 as=0 ps=0 
M2143 diff_3635_3892# diff_3610_3644# diff_1663_3859# GND efet w=58 l=19
+ ad=1625 pd=198 as=0 ps=0 
M2144 diff_1370_3857# diff_3484_3742# diff_3385_3844# GND efet w=19 l=16
+ ad=0 pd=0 as=1521 ps=182 
M2145 diff_3575_3844# diff_3556_3644# diff_1370_3857# GND efet w=19 l=16
+ ad=1446 pd=176 as=0 ps=0 
M2146 GND diff_3575_3844# diff_3635_3892# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2147 diff_3752_3880# diff_3727_3844# GND GND efet w=52 l=19
+ ad=1469 pd=192 as=0 ps=0 
M2148 diff_1663_3859# diff_3739_3610# diff_3752_3880# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2149 diff_3917_4054# diff_3898_3644# diff_1370_4027# GND efet w=19 l=16
+ ad=1431 pd=182 as=0 ps=0 
M2150 GND diff_3917_4195# diff_3980_4246# GND efet w=55 l=19
+ ad=0 pd=0 as=0 ps=0 
M2151 diff_4094_4231# diff_4072_4195# GND GND efet w=55 l=16
+ ad=1502 pd=186 as=0 ps=0 
M2152 diff_1663_4210# diff_4084_3607# diff_4094_4231# GND efet w=49 l=19
+ ad=0 pd=0 as=0 ps=0 
M2153 diff_1370_4211# diff_4171_3745# diff_4072_4195# GND efet w=19 l=16
+ ad=0 pd=0 as=1434 ps=188 
M2154 diff_4325_4327# diff_4300_3644# diff_1663_4402# GND efet w=52 l=19
+ ad=1409 pd=186 as=0 ps=0 
M2155 GND diff_4262_4411# diff_4325_4327# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2156 diff_4439_4336# diff_4414_4408# GND GND efet w=55 l=16
+ ad=1517 pd=186 as=0 ps=0 
M2157 GND diff_4607_4906# diff_4667_4957# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2158 diff_4784_4942# diff_4759_4906# GND GND efet w=55 l=16
+ ad=1499 pd=180 as=0 ps=0 
M2159 diff_1663_4918# diff_4771_3607# diff_4784_4942# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M2160 diff_4667_4681# diff_4642_3644# diff_1663_4756# GND efet w=52 l=16
+ ad=1715 pd=192 as=0 ps=0 
M2161 GND diff_4607_4765# diff_4667_4681# GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M2162 diff_4784_4690# diff_4759_4759# GND GND efet w=58 l=16
+ ad=1568 pd=186 as=0 ps=0 
M2163 GND diff_4949_5263# diff_5012_5311# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2164 diff_5129_5299# diff_5104_5260# GND GND efet w=62 l=17
+ ad=1487 pd=180 as=0 ps=0 
M2165 diff_1663_5275# diff_5116_3613# diff_5129_5299# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2166 diff_5012_5038# diff_4987_3652# diff_1663_5113# GND efet w=52 l=16
+ ad=1664 pd=192 as=0 ps=0 
M2167 GND diff_4949_5122# diff_5012_5038# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2168 diff_5129_5047# diff_5104_5113# GND GND efet w=56 l=17
+ ad=1487 pd=180 as=0 ps=0 
M2169 diff_5294_5476# diff_5278_3644# diff_1370_5446# GND efet w=16 l=16
+ ad=1446 pd=188 as=0 ps=0 
M2170 GND diff_5294_5614# diff_5357_5665# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2171 Vdd diff_5563_3961# diff_1663_5629# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M2172 Vdd diff_4732_1658# diff_1370_5630# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M2173 Vdd diff_4732_1658# diff_1370_5446# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M2174 GND diff_5294_5476# diff_5357_5395# GND efet w=53 l=17
+ ad=0 pd=0 as=1595 ps=186 
M2175 diff_5357_5395# diff_5335_3644# diff_1663_5467# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M2176 Vdd diff_5563_3961# diff_1663_5467# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M2177 diff_6043_4888# Vdd Vdd GND efet w=25 l=46
+ ad=8184 pd=646 as=0 ps=0 
M2178 diff_5813_5371# clk2 diff_580_3394# GND efet w=46 l=16
+ ad=1679 pd=192 as=0 ps=0 
M2179 diff_5357_5311# diff_5335_3644# diff_1663_5275# GND efet w=52 l=16
+ ad=1661 pd=186 as=0 ps=0 
M2180 diff_1370_5273# diff_5206_3742# diff_5104_5260# GND efet w=16 l=16
+ ad=0 pd=0 as=1470 ps=182 
M2181 diff_5294_5263# diff_5278_3644# diff_1370_5273# GND efet w=16 l=16
+ ad=1464 pd=188 as=0 ps=0 
M2182 diff_1370_5092# diff_5206_3742# diff_5104_5113# GND efet w=19 l=19
+ ad=0 pd=0 as=1476 ps=182 
M2183 diff_1663_5113# diff_5116_3613# diff_5129_5047# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2184 diff_5294_5122# diff_5278_3644# diff_1370_5092# GND efet w=16 l=16
+ ad=1473 pd=188 as=0 ps=0 
M2185 diff_5012_4957# diff_4987_3652# diff_1663_4918# GND efet w=49 l=16
+ ad=1646 pd=186 as=0 ps=0 
M2186 diff_1370_4919# diff_4861_3742# diff_4759_4906# GND efet w=19 l=16
+ ad=0 pd=0 as=1452 ps=188 
M2187 diff_4949_4906# diff_4933_3644# diff_1370_4919# GND efet w=19 l=16
+ ad=1470 pd=188 as=0 ps=0 
M2188 diff_1370_4735# diff_4861_3742# diff_4759_4759# GND efet w=19 l=16
+ ad=0 pd=0 as=1515 ps=188 
M2189 diff_1663_4756# diff_4771_3607# diff_4784_4690# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2190 diff_4667_4600# diff_4642_3644# diff_1663_4564# GND efet w=52 l=16
+ ad=1679 pd=186 as=0 ps=0 
M2191 diff_1370_4565# diff_4516_3742# diff_4414_4558# GND efet w=22 l=16
+ ad=0 pd=0 as=1506 ps=194 
M2192 diff_4607_4549# diff_4588_3644# diff_1370_4565# GND efet w=26 l=17
+ ad=1467 pd=188 as=0 ps=0 
M2193 diff_1370_4381# diff_4516_3742# diff_4414_4408# GND efet w=19 l=16
+ ad=0 pd=0 as=1542 ps=188 
M2194 diff_1663_4402# diff_4426_3610# diff_4439_4336# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2195 diff_4325_4246# diff_4300_3644# diff_1663_4210# GND efet w=49 l=19
+ ad=1502 pd=186 as=0 ps=0 
M2196 diff_1663_4210# diff_4426_3610# diff_4439_4231# GND efet w=52 l=19
+ ad=0 pd=0 as=1517 ps=180 
M2197 diff_4262_4195# diff_4243_3644# diff_1370_4211# GND efet w=19 l=16
+ ad=1449 pd=182 as=0 ps=0 
M2198 diff_3980_3973# diff_3955_3644# diff_1663_4051# GND efet w=50 l=17
+ ad=1514 pd=180 as=0 ps=0 
M2199 GND diff_3917_4054# diff_3980_3973# GND efet w=55 l=19
+ ad=0 pd=0 as=0 ps=0 
M2200 diff_4094_3982# diff_4072_4051# GND GND efet w=55 l=16
+ ad=1538 pd=186 as=0 ps=0 
M2201 GND diff_4262_4195# diff_4325_4246# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2202 diff_4439_4231# diff_4414_4198# GND GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2203 diff_1370_4027# diff_4171_3745# diff_4072_4051# GND efet w=19 l=16
+ ad=0 pd=0 as=1422 ps=182 
M2204 diff_1663_4051# diff_4084_3607# diff_4094_3982# GND efet w=53 l=20
+ ad=0 pd=0 as=0 ps=0 
M2205 diff_3980_3892# diff_3955_3644# diff_1663_3859# GND efet w=49 l=16
+ ad=1493 pd=186 as=0 ps=0 
M2206 diff_1663_3859# diff_4084_3607# diff_4094_3877# GND efet w=50 l=17
+ ad=0 pd=0 as=1520 ps=192 
M2207 diff_1370_3857# diff_3829_3644# diff_3727_3844# GND efet w=22 l=16
+ ad=0 pd=0 as=1551 ps=194 
M2208 diff_3917_3841# diff_3898_3644# diff_1370_3857# GND efet w=22 l=16
+ ad=1536 pd=182 as=0 ps=0 
M2209 GND diff_3917_3841# diff_3980_3892# GND efet w=55 l=19
+ ad=0 pd=0 as=0 ps=0 
M2210 diff_4094_3877# diff_4072_3844# GND GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2211 diff_4262_4054# diff_4243_3644# diff_1370_4027# GND efet w=19 l=16
+ ad=1371 pd=188 as=0 ps=0 
M2212 diff_4325_3973# diff_4300_3644# diff_1663_4051# GND efet w=50 l=20
+ ad=1514 pd=180 as=0 ps=0 
M2213 GND diff_4262_4054# diff_4325_3973# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2214 diff_4439_3982# diff_4414_4054# GND GND efet w=55 l=16
+ ad=1514 pd=180 as=0 ps=0 
M2215 diff_4607_4411# diff_4588_3644# diff_1370_4381# GND efet w=19 l=19
+ ad=1488 pd=188 as=0 ps=0 
M2216 GND diff_4607_4549# diff_4667_4600# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2217 diff_4784_4588# diff_4759_4552# GND GND efet w=55 l=16
+ ad=1514 pd=180 as=0 ps=0 
M2218 diff_1663_4564# diff_4771_3607# diff_4784_4588# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2219 diff_1370_4211# diff_4516_3742# diff_4414_4198# GND efet w=19 l=16
+ ad=0 pd=0 as=1521 ps=182 
M2220 diff_4667_4327# diff_4642_3644# diff_1663_4402# GND efet w=52 l=16
+ ad=1673 pd=192 as=0 ps=0 
M2221 GND diff_4607_4411# diff_4667_4327# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2222 diff_4784_4336# diff_4759_4405# GND GND efet w=55 l=16
+ ad=1505 pd=180 as=0 ps=0 
M2223 diff_4949_4765# diff_4933_3644# diff_1370_4735# GND efet w=19 l=16
+ ad=1482 pd=194 as=0 ps=0 
M2224 GND diff_4949_4906# diff_5012_4957# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2225 diff_5129_4942# diff_5104_4906# GND GND efet w=55 l=16
+ ad=1484 pd=186 as=0 ps=0 
M2226 diff_1663_4918# diff_5116_3613# diff_5129_4942# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M2227 diff_5012_4684# diff_4987_3652# diff_1663_4756# GND efet w=49 l=16
+ ad=1670 pd=186 as=0 ps=0 
M2228 GND diff_4949_4765# diff_5012_4684# GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M2229 diff_5129_4690# diff_5104_4759# GND GND efet w=55 l=16
+ ad=1442 pd=174 as=0 ps=0 
M2230 diff_1370_4919# diff_5206_3742# diff_5104_4906# GND efet w=19 l=16
+ ad=0 pd=0 as=1431 ps=182 
M2231 GND diff_5294_5263# diff_5357_5311# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2232 diff_5861_5353# diff_5188_6931# diff_5813_5371# GND efet w=46 l=16
+ ad=10067 pd=836 as=0 ps=0 
M2233 Vdd diff_5563_3961# diff_1663_5275# GND efet w=37 l=16
+ ad=0 pd=0 as=0 ps=0 
M2234 GND diff_5188_6931# diff_6062_5224# GND efet w=34 l=14
+ ad=0 pd=0 as=2087 ps=198 
M2235 GND diff_5194_7252# diff_5861_5353# GND efet w=67 l=13
+ ad=0 pd=0 as=0 ps=0 
M2236 Vdd diff_4732_1658# diff_1370_5273# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M2237 diff_6062_5224# Vdd Vdd GND efet w=20 l=143
+ ad=0 pd=0 as=0 ps=0 
M2238 Vdd Vdd Vdd GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M2239 Vdd diff_4732_1658# diff_1370_5092# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M2240 diff_5861_5353# diff_6062_5224# diff_6137_5167# GND efet w=34 l=13
+ ad=0 pd=0 as=4012 ps=370 
M2241 diff_6043_4888# diff_5861_5353# GND GND efet w=277 l=16
+ ad=0 pd=0 as=0 ps=0 
M2242 Vdd Vdd Vdd GND efet w=10 l=19
+ ad=0 pd=0 as=0 ps=0 
M2243 diff_6137_5167# Vdd Vdd GND efet w=22 l=74
+ ad=0 pd=0 as=0 ps=0 
M2244 diff_5357_5038# diff_5335_3644# diff_1663_5113# GND efet w=52 l=16
+ ad=1664 pd=192 as=0 ps=0 
M2245 GND diff_5294_5122# diff_5357_5038# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2246 Vdd diff_5563_3961# diff_1663_5113# GND efet w=37 l=13
+ ad=0 pd=0 as=0 ps=0 
M2247 diff_5357_4957# diff_5335_3644# diff_1663_4918# GND efet w=49 l=16
+ ad=1640 pd=192 as=0 ps=0 
M2248 diff_5294_4906# diff_5278_3644# diff_1370_4919# GND efet w=19 l=16
+ ad=1419 pd=194 as=0 ps=0 
M2249 diff_1370_4735# diff_5206_3742# diff_5104_4759# GND efet w=19 l=16
+ ad=0 pd=0 as=1458 ps=182 
M2250 diff_1663_4756# diff_5116_3613# diff_5129_4690# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M2251 diff_5012_4600# diff_4987_3652# diff_1663_4564# GND efet w=52 l=16
+ ad=1661 pd=186 as=0 ps=0 
M2252 diff_1370_4565# diff_4861_3742# diff_4759_4552# GND efet w=19 l=16
+ ad=0 pd=0 as=1521 ps=182 
M2253 diff_4949_4552# diff_4933_3644# diff_1370_4565# GND efet w=22 l=16
+ ad=1410 pd=188 as=0 ps=0 
M2254 diff_1370_4381# diff_4861_3742# diff_4759_4405# GND efet w=19 l=16
+ ad=0 pd=0 as=1494 ps=182 
M2255 diff_1663_4402# diff_4771_3607# diff_4784_4336# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2256 diff_4667_4246# diff_4642_3644# diff_1663_4210# GND efet w=49 l=16
+ ad=1658 pd=192 as=0 ps=0 
M2257 diff_4607_4195# diff_4588_3644# diff_1370_4211# GND efet w=19 l=19
+ ad=1452 pd=188 as=0 ps=0 
M2258 diff_1370_4027# diff_4516_3742# diff_4414_4054# GND efet w=19 l=16
+ ad=0 pd=0 as=1512 ps=182 
M2259 diff_1663_4051# diff_4426_3610# diff_4439_3982# GND efet w=50 l=17
+ ad=0 pd=0 as=0 ps=0 
M2260 diff_4325_3892# diff_4300_3644# diff_1663_3859# GND efet w=49 l=19
+ ad=1502 pd=186 as=0 ps=0 
M2261 diff_1663_3859# diff_4426_3610# diff_4439_3877# GND efet w=49 l=19
+ ad=0 pd=0 as=1517 ps=180 
M2262 diff_1370_3857# diff_4171_3745# diff_4072_3844# GND efet w=22 l=16
+ ad=0 pd=0 as=1455 ps=182 
M2263 diff_4262_3841# diff_4243_3644# diff_1370_3857# GND efet w=22 l=16
+ ad=1455 pd=182 as=0 ps=0 
M2264 GND diff_4262_3841# diff_4325_3892# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2265 diff_4439_3877# diff_4414_3847# GND GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2266 diff_4607_4054# diff_4588_3644# diff_1370_4027# GND efet w=19 l=19
+ ad=1401 pd=194 as=0 ps=0 
M2267 GND diff_4607_4195# diff_4667_4246# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2268 diff_4784_4231# diff_4759_4198# GND GND efet w=61 l=19
+ ad=1517 pd=180 as=0 ps=0 
M2269 diff_1663_4210# diff_4771_3607# diff_4784_4231# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M2270 diff_4667_3973# diff_4642_3644# diff_1663_4051# GND efet w=50 l=17
+ ad=1661 pd=186 as=0 ps=0 
M2271 GND diff_4607_4054# diff_4667_3973# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2272 diff_4784_3982# diff_4759_4051# GND GND efet w=56 l=17
+ ad=1505 pd=180 as=0 ps=0 
M2273 diff_4949_4411# diff_4933_3644# diff_1370_4381# GND efet w=19 l=16
+ ad=1452 pd=188 as=0 ps=0 
M2274 diff_1370_4211# diff_4861_3742# diff_4759_4198# GND efet w=19 l=16
+ ad=0 pd=0 as=1512 ps=182 
M2275 GND diff_4949_4552# diff_5012_4600# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2276 diff_5129_4588# diff_5104_4552# GND GND efet w=55 l=16
+ ad=1487 pd=180 as=0 ps=0 
M2277 diff_1663_4564# diff_5116_3613# diff_5129_4588# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2278 diff_5012_4327# diff_4987_3652# diff_1663_4402# GND efet w=52 l=16
+ ad=1664 pd=192 as=0 ps=0 
M2279 GND diff_4949_4411# diff_5012_4327# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2280 diff_5129_4336# diff_5104_4405# GND GND efet w=61 l=17
+ ad=1487 pd=180 as=0 ps=0 
M2281 diff_5294_4765# diff_5278_3644# diff_1370_4735# GND efet w=19 l=16
+ ad=1434 pd=188 as=0 ps=0 
M2282 GND diff_5294_4906# diff_5357_4957# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2283 o3 diff_5938_5011# Vdd GND efet w=514 l=16
+ ad=25515 pd=1702 as=0 ps=0 
M2284 diff_6137_5167# diff_6043_4888# GND GND efet w=67 l=16
+ ad=0 pd=0 as=0 ps=0 
M2285 o3 diff_6043_4888# GND GND efet w=482 l=14
+ ad=0 pd=0 as=0 ps=0 
M2286 Vdd diff_5563_3961# diff_1663_4918# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M2287 Vdd diff_4732_1658# diff_1370_4919# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M2288 diff_5938_5011# diff_5938_5011# diff_5938_5011# GND efet w=2 l=5
+ ad=6102 pd=424 as=0 ps=0 
M2289 diff_5938_5011# Vdd Vdd GND efet w=28 l=44
+ ad=0 pd=0 as=0 ps=0 
M2290 diff_5938_5011# diff_5938_5011# diff_5938_5011# GND efet w=4 l=4
+ ad=0 pd=0 as=0 ps=0 
M2291 diff_5938_5011# diff_6043_4888# GND GND efet w=125 l=14
+ ad=0 pd=0 as=0 ps=0 
M2292 Vdd diff_4732_1658# diff_1370_4735# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M2293 diff_5357_4684# diff_5335_3644# diff_1663_4756# GND efet w=49 l=16
+ ad=1646 pd=186 as=0 ps=0 
M2294 GND diff_5294_4765# diff_5357_4684# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2295 Vdd diff_5563_3961# diff_1663_4756# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M2296 diff_5357_4600# diff_5335_3644# diff_1663_4564# GND efet w=50 l=17
+ ad=1661 pd=186 as=0 ps=0 
M2297 diff_1370_4565# diff_5206_3742# diff_5104_4552# GND efet w=19 l=16
+ ad=0 pd=0 as=1494 ps=182 
M2298 diff_5294_4552# diff_5278_3644# diff_1370_4565# GND efet w=19 l=16
+ ad=1518 pd=194 as=0 ps=0 
M2299 diff_1370_4381# diff_5206_3742# diff_5104_4405# GND efet w=19 l=16
+ ad=0 pd=0 as=1524 ps=188 
M2300 diff_1663_4402# diff_5116_3613# diff_5129_4336# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2301 diff_5294_4411# diff_5278_3644# diff_1370_4381# GND efet w=19 l=16
+ ad=1452 pd=188 as=0 ps=0 
M2302 diff_5012_4246# diff_4987_3652# diff_1663_4210# GND efet w=49 l=16
+ ad=1640 pd=192 as=0 ps=0 
M2303 diff_4949_4195# diff_4933_3644# diff_1370_4211# GND efet w=19 l=16
+ ad=1500 pd=194 as=0 ps=0 
M2304 diff_1370_4027# diff_4861_3742# diff_4759_4051# GND efet w=19 l=16
+ ad=0 pd=0 as=1494 ps=182 
M2305 diff_1663_4051# diff_4771_3607# diff_4784_3982# GND efet w=50 l=17
+ ad=0 pd=0 as=0 ps=0 
M2306 diff_4667_3892# diff_4642_3644# diff_1663_3859# GND efet w=49 l=16
+ ad=1649 pd=192 as=0 ps=0 
M2307 diff_1370_3857# diff_4516_3742# diff_4414_3847# GND efet w=22 l=16
+ ad=0 pd=0 as=1536 ps=182 
M2308 diff_4607_3841# diff_4588_3644# diff_1370_3857# GND efet w=25 l=19
+ ad=1461 pd=176 as=0 ps=0 
M2309 GND diff_4607_3841# diff_4667_3892# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2310 diff_4784_3877# diff_4759_3844# GND GND efet w=55 l=19
+ ad=1490 pd=180 as=0 ps=0 
M2311 diff_1663_3859# diff_4771_3607# diff_4784_3877# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M2312 diff_4949_4054# diff_4933_3644# diff_1370_4027# GND efet w=19 l=16
+ ad=1461 pd=188 as=0 ps=0 
M2313 GND diff_4949_4195# diff_5012_4246# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2314 diff_5129_4231# diff_5104_4198# GND GND efet w=56 l=17
+ ad=1472 pd=180 as=0 ps=0 
M2315 diff_1663_4210# diff_5116_3613# diff_5129_4231# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M2316 diff_5012_3973# diff_4987_3652# diff_1663_4051# GND efet w=50 l=17
+ ad=1652 pd=186 as=0 ps=0 
M2317 GND diff_4949_4054# diff_5012_3973# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2318 diff_5129_3982# diff_5104_4051# GND GND efet w=55 l=19
+ ad=1487 pd=180 as=0 ps=0 
M2319 diff_1370_4211# diff_5206_3742# diff_5104_4198# GND efet w=22 l=16
+ ad=0 pd=0 as=1491 ps=188 
M2320 GND diff_5294_4552# diff_5357_4600# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2321 Vdd diff_5563_3961# diff_1663_4564# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M2322 Vdd diff_4732_1658# diff_1370_4565# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M2323 Vdd diff_4732_1658# diff_1370_4381# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M2324 diff_5357_4327# diff_5335_3644# diff_1663_4402# GND efet w=52 l=16
+ ad=1697 pd=192 as=0 ps=0 
M2325 GND diff_5294_4411# diff_5357_4327# GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M2326 Vdd diff_5563_3961# diff_1663_4402# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M2327 GND diff_4481_442# diff_5194_7252# GND efet w=130 l=13
+ ad=0 pd=0 as=4619 ps=372 
M2328 diff_5357_4246# diff_5335_3644# diff_1663_4210# GND efet w=52 l=16
+ ad=1652 pd=186 as=0 ps=0 
M2329 diff_5294_4195# diff_5278_3644# diff_1370_4211# GND efet w=19 l=16
+ ad=1500 pd=194 as=0 ps=0 
M2330 diff_1370_4027# diff_5206_3742# diff_5104_4051# GND efet w=19 l=16
+ ad=0 pd=0 as=1488 ps=188 
M2331 diff_1663_4051# diff_5116_3613# diff_5129_3982# GND efet w=50 l=17
+ ad=0 pd=0 as=0 ps=0 
M2332 diff_5012_3892# diff_4987_3652# diff_1663_3859# GND efet w=49 l=16
+ ad=1583 pd=180 as=0 ps=0 
M2333 diff_5294_4054# diff_5278_3644# diff_1370_4027# GND efet w=19 l=16
+ ad=1512 pd=182 as=0 ps=0 
M2334 diff_1370_3857# diff_4861_3742# diff_4759_3844# GND efet w=19 l=16
+ ad=0 pd=0 as=1530 ps=182 
M2335 diff_4949_3844# diff_4933_3644# diff_1370_3857# GND efet w=19 l=16
+ ad=1503 pd=182 as=0 ps=0 
M2336 GND diff_4949_3844# diff_5012_3892# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2337 diff_5129_3880# diff_5104_3844# GND GND efet w=52 l=19
+ ad=1427 pd=174 as=0 ps=0 
M2338 diff_1663_3859# diff_5116_3613# diff_5129_3880# GND efet w=49 l=16
+ ad=0 pd=0 as=0 ps=0 
M2339 GND diff_5294_4195# diff_5357_4246# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2340 Vdd diff_5563_3961# diff_1663_4210# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M2341 Vdd diff_4732_1658# diff_1370_4211# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M2342 diff_5194_7252# Vdd Vdd GND efet w=25 l=44
+ ad=0 pd=0 as=0 ps=0 
M2343 Vdd diff_4732_1658# diff_1370_4027# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M2344 diff_5563_3961# diff_5705_4015# diff_5563_3961# GND efet w=74 l=77
+ ad=9419 pd=652 as=0 ps=0 
M2345 diff_5357_3973# diff_5335_3644# diff_1663_4051# GND efet w=52 l=16
+ ad=1634 pd=186 as=0 ps=0 
M2346 GND diff_5294_4054# diff_5357_3973# GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2347 Vdd diff_5563_3961# diff_1663_4051# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M2348 diff_5705_4015# Vdd Vdd GND efet w=19 l=16
+ ad=1561 pd=196 as=0 ps=0 
M2349 diff_5705_4015# diff_5705_4015# diff_5705_4015# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M2350 diff_5705_4015# diff_5705_4015# diff_5705_4015# GND efet w=5 l=15
+ ad=0 pd=0 as=0 ps=0 
M2351 GND diff_5855_3847# diff_5563_3961# GND efet w=184 l=16
+ ad=0 pd=0 as=0 ps=0 
M2352 diff_5563_3961# diff_5705_4015# Vdd GND efet w=25 l=28
+ ad=0 pd=0 as=0 ps=0 
M2353 diff_5563_3961# diff_5563_3961# diff_5563_3961# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M2354 diff_5563_3961# diff_5563_3961# diff_5563_3961# GND efet w=8 l=8
+ ad=0 pd=0 as=0 ps=0 
M2355 diff_5357_3892# diff_5335_3644# diff_1663_3859# GND efet w=52 l=16
+ ad=1628 pd=186 as=0 ps=0 
M2356 diff_1370_3857# diff_5206_3742# diff_5104_3844# GND efet w=19 l=16
+ ad=0 pd=0 as=1404 ps=182 
M2357 diff_5294_3844# diff_5278_3644# diff_1370_3857# GND efet w=16 l=19
+ ad=1479 pd=182 as=0 ps=0 
M2358 GND diff_5294_3844# diff_5357_3892# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2359 Vdd diff_5563_3961# diff_1663_3859# GND efet w=32 l=16
+ ad=0 pd=0 as=0 ps=0 
M2360 diff_5855_3847# Vdd Vdd GND efet w=25 l=46
+ ad=5897 pd=436 as=0 ps=0 
M2361 Vdd diff_4732_1658# diff_1370_3857# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M2362 diff_5855_3847# clk1 diff_5866_3757# GND efet w=181 l=16
+ ad=0 pd=0 as=8360 ps=662 
M2363 GND diff_5849_3703# diff_5866_3757# GND efet w=283 l=16
+ ad=0 pd=0 as=0 ps=0 
M2364 GND diff_1996_3562# diff_2020_3610# GND efet w=43 l=19
+ ad=0 pd=0 as=3344 ps=296 
M2365 GND diff_1996_3562# diff_2110_3745# GND efet w=28 l=19
+ ad=0 pd=0 as=1232 ps=144 
M2366 GND diff_2170_3691# diff_2182_3644# GND efet w=28 l=19
+ ad=0 pd=0 as=1232 ps=144 
M2367 GND diff_2170_3691# diff_2236_3644# GND efet w=43 l=19
+ ad=0 pd=0 as=3068 ps=290 
M2368 Vdd Vdd diff_1093_4033# GND efet w=25 l=94
+ ad=0 pd=0 as=6459 ps=660 
M2369 Vdd Vdd diff_829_3778# GND efet w=25 l=103
+ ad=0 pd=0 as=9084 ps=858 
M2370 diff_820_3511# diff_820_3511# diff_820_3511# GND efet w=7 l=7
+ ad=7995 pd=694 as=0 ps=0 
M2371 Vdd Vdd diff_820_3511# GND efet w=25 l=91
+ ad=0 pd=0 as=0 ps=0 
M2372 diff_820_3511# diff_820_3511# diff_820_3511# GND efet w=3 l=7
+ ad=0 pd=0 as=0 ps=0 
M2373 diff_1066_3979# diff_1786_2191# Vdd GND efet w=94 l=16
+ ad=15472 pd=1082 as=0 ps=0 
M2374 GND diff_1829_3439# diff_1066_3979# GND efet w=94 l=16
+ ad=0 pd=0 as=0 ps=0 
M2375 diff_2053_3553# diff_2026_2897# diff_2020_3610# GND efet w=76 l=24
+ ad=54830 pd=5644 as=0 ps=0 
M2376 diff_2110_3745# diff_2026_2897# diff_2113_3589# GND efet w=29 l=17
+ ad=0 pd=0 as=51738 ps=5000 
M2377 diff_2182_3644# diff_2170_3631# diff_2113_3589# GND efet w=29 l=17
+ ad=0 pd=0 as=0 ps=0 
M2378 diff_817_6145# diff_817_6145# diff_817_6145# GND efet w=8 l=8
+ ad=6655 pd=700 as=0 ps=0 
M2379 Vdd Vdd diff_817_6145# GND efet w=25 l=94
+ ad=0 pd=0 as=0 ps=0 
M2380 diff_817_6145# diff_817_6145# diff_817_6145# GND efet w=7 l=7
+ ad=0 pd=0 as=0 ps=0 
M2381 GND diff_407_3110# diff_580_3394# GND efet w=95 l=14
+ ad=0 pd=0 as=0 ps=0 
M2382 diff_1829_3439# Vdd Vdd GND efet w=19 l=94
+ ad=2915 pd=270 as=0 ps=0 
M2383 diff_2236_3644# diff_2170_3631# diff_2053_3553# GND efet w=76 l=24
+ ad=0 pd=0 as=0 ps=0 
M2384 GND diff_2344_3556# diff_2365_3607# GND efet w=43 l=19
+ ad=0 pd=0 as=3170 ps=290 
M2385 GND diff_2344_3556# diff_2455_3644# GND efet w=31 l=19
+ ad=0 pd=0 as=1364 ps=150 
M2386 GND diff_2515_3691# diff_2524_3644# GND efet w=31 l=19
+ ad=0 pd=0 as=1232 ps=144 
M2387 GND diff_2515_3691# diff_2581_3644# GND efet w=40 l=19
+ ad=0 pd=0 as=3035 ps=290 
M2388 diff_2053_3553# diff_2368_2803# diff_2365_3607# GND efet w=76 l=24
+ ad=0 pd=0 as=0 ps=0 
M2389 diff_2455_3644# diff_2368_2803# diff_2113_3589# GND efet w=34 l=19
+ ad=0 pd=0 as=0 ps=0 
M2390 diff_2524_3644# diff_2515_3628# diff_2113_3589# GND efet w=29 l=17
+ ad=0 pd=0 as=0 ps=0 
M2391 diff_2581_3644# diff_2515_3628# diff_2053_3553# GND efet w=75 l=26
+ ad=0 pd=0 as=0 ps=0 
M2392 GND diff_2689_3475# diff_2707_3610# GND efet w=43 l=19
+ ad=0 pd=0 as=3320 ps=302 
M2393 GND diff_2689_3475# diff_2797_3745# GND efet w=28 l=19
+ ad=0 pd=0 as=1232 ps=144 
M2394 GND diff_2857_3691# diff_2869_3644# GND efet w=28 l=19
+ ad=0 pd=0 as=1232 ps=144 
M2395 GND diff_2857_3691# diff_2923_3644# GND efet w=43 l=19
+ ad=0 pd=0 as=3215 ps=296 
M2396 diff_2053_3553# diff_2713_2900# diff_2707_3610# GND efet w=82 l=24
+ ad=0 pd=0 as=0 ps=0 
M2397 diff_2797_3745# diff_2713_2900# diff_2113_3589# GND efet w=29 l=17
+ ad=0 pd=0 as=0 ps=0 
M2398 diff_2869_3644# diff_2857_3628# diff_2113_3589# GND efet w=29 l=17
+ ad=0 pd=0 as=0 ps=0 
M2399 diff_2923_3644# diff_2857_3628# diff_2053_3553# GND efet w=76 l=24
+ ad=0 pd=0 as=0 ps=0 
M2400 GND diff_3031_3556# diff_3052_3607# GND efet w=40 l=19
+ ad=0 pd=0 as=3119 ps=290 
M2401 GND diff_3031_3556# diff_3142_3644# GND efet w=31 l=19
+ ad=0 pd=0 as=1364 ps=150 
M2402 GND diff_3202_3691# diff_3211_3644# GND efet w=31 l=19
+ ad=0 pd=0 as=1364 ps=150 
M2403 GND diff_3202_3691# diff_3268_3644# GND efet w=40 l=19
+ ad=0 pd=0 as=3098 ps=290 
M2404 diff_2053_3553# diff_3055_2897# diff_3052_3607# GND efet w=73 l=24
+ ad=0 pd=0 as=0 ps=0 
M2405 diff_3142_3644# diff_3055_2897# diff_2113_3589# GND efet w=32 l=17
+ ad=0 pd=0 as=0 ps=0 
M2406 diff_3211_3644# diff_3202_3628# diff_2113_3589# GND efet w=35 l=17
+ ad=0 pd=0 as=0 ps=0 
M2407 diff_3268_3644# diff_3202_3628# diff_2053_3553# GND efet w=75 l=26
+ ad=0 pd=0 as=0 ps=0 
M2408 GND diff_3376_3475# diff_3394_3613# GND efet w=43 l=19
+ ad=0 pd=0 as=3215 ps=296 
M2409 GND diff_3376_3475# diff_3484_3742# GND efet w=28 l=19
+ ad=0 pd=0 as=1232 ps=144 
M2410 GND diff_3544_3691# diff_3556_3644# GND efet w=28 l=19
+ ad=0 pd=0 as=1232 ps=144 
M2411 GND diff_3544_3691# diff_3610_3644# GND efet w=43 l=19
+ ad=0 pd=0 as=3233 ps=296 
M2412 diff_2053_3553# diff_3400_2897# diff_3394_3613# GND efet w=79 l=24
+ ad=0 pd=0 as=0 ps=0 
M2413 diff_3484_3742# diff_3400_2897# diff_2113_3589# GND efet w=29 l=17
+ ad=0 pd=0 as=0 ps=0 
M2414 diff_3556_3644# diff_3544_3628# diff_2113_3589# GND efet w=29 l=17
+ ad=0 pd=0 as=0 ps=0 
M2415 diff_3610_3644# diff_3544_3628# diff_2053_3553# GND efet w=76 l=24
+ ad=0 pd=0 as=0 ps=0 
M2416 GND diff_3718_3556# diff_3739_3610# GND efet w=43 l=19
+ ad=0 pd=0 as=3110 ps=296 
M2417 GND diff_3718_3556# diff_3829_3644# GND efet w=31 l=17
+ ad=0 pd=0 as=1364 ps=150 
M2418 GND diff_3889_3691# diff_3898_3644# GND efet w=29 l=19
+ ad=0 pd=0 as=1364 ps=150 
M2419 GND diff_3889_3691# diff_3955_3644# GND efet w=43 l=19
+ ad=0 pd=0 as=3095 ps=290 
M2420 diff_2053_3553# diff_3745_2897# diff_3739_3610# GND efet w=76 l=24
+ ad=0 pd=0 as=0 ps=0 
M2421 diff_3829_3644# diff_3745_2897# diff_2113_3589# GND efet w=32 l=17
+ ad=0 pd=0 as=0 ps=0 
M2422 diff_3898_3644# diff_3889_3628# diff_2113_3589# GND efet w=32 l=17
+ ad=0 pd=0 as=0 ps=0 
M2423 diff_3955_3644# diff_3889_3628# diff_2053_3553# GND efet w=78 l=26
+ ad=0 pd=0 as=0 ps=0 
M2424 GND diff_4063_3493# diff_4084_3607# GND efet w=43 l=19
+ ad=0 pd=0 as=3104 ps=290 
M2425 GND diff_4063_3493# diff_4171_3745# GND efet w=29 l=17
+ ad=0 pd=0 as=1232 ps=144 
M2426 GND diff_4231_3691# diff_4243_3644# GND efet w=28 l=19
+ ad=0 pd=0 as=1232 ps=144 
M2427 GND diff_4231_3691# diff_4300_3644# GND efet w=40 l=19
+ ad=0 pd=0 as=3101 ps=290 
M2428 diff_2053_3553# diff_4087_2900# diff_4084_3607# GND efet w=79 l=24
+ ad=0 pd=0 as=0 ps=0 
M2429 diff_4171_3745# diff_4087_2900# diff_2113_3589# GND efet w=29 l=17
+ ad=0 pd=0 as=0 ps=0 
M2430 diff_4243_3644# diff_4231_3628# diff_2113_3589# GND efet w=29 l=17
+ ad=0 pd=0 as=0 ps=0 
M2431 diff_4300_3644# diff_4231_3628# diff_2053_3553# GND efet w=76 l=24
+ ad=0 pd=0 as=0 ps=0 
M2432 GND diff_4405_3556# diff_4426_3610# GND efet w=43 l=19
+ ad=0 pd=0 as=3224 ps=296 
M2433 GND diff_4405_3556# diff_4516_3742# GND efet w=28 l=17
+ ad=0 pd=0 as=1232 ps=144 
M2434 GND diff_4576_3691# diff_4588_3644# GND efet w=28 l=19
+ ad=0 pd=0 as=1232 ps=144 
M2435 GND diff_4576_3691# diff_4642_3644# GND efet w=46 l=19
+ ad=0 pd=0 as=3257 ps=302 
M2436 diff_2053_3553# diff_4399_2803# diff_4426_3610# GND efet w=79 l=24
+ ad=0 pd=0 as=0 ps=0 
M2437 diff_4516_3742# diff_4399_2803# diff_2113_3589# GND efet w=29 l=17
+ ad=0 pd=0 as=0 ps=0 
M2438 diff_4588_3644# diff_4552_2860# diff_2113_3589# GND efet w=29 l=17
+ ad=0 pd=0 as=0 ps=0 
M2439 diff_4642_3644# diff_4552_2860# diff_2053_3553# GND efet w=79 l=24
+ ad=0 pd=0 as=0 ps=0 
M2440 GND diff_4750_3556# diff_4771_3607# GND efet w=47 l=17
+ ad=0 pd=0 as=3164 ps=314 
M2441 GND diff_4750_3556# diff_4861_3742# GND efet w=28 l=16
+ ad=0 pd=0 as=1316 ps=150 
M2442 GND diff_4921_3691# diff_4933_3644# GND efet w=31 l=16
+ ad=0 pd=0 as=1304 ps=156 
M2443 diff_4987_3652# diff_4921_3691# GND GND efet w=41 l=17
+ ad=3260 pd=302 as=0 ps=0 
M2444 diff_2053_3553# diff_4732_2900# diff_4771_3607# GND efet w=75 l=26
+ ad=0 pd=0 as=0 ps=0 
M2445 diff_4861_3742# diff_4732_2900# diff_2113_3589# GND efet w=28 l=16
+ ad=0 pd=0 as=0 ps=0 
M2446 diff_4933_3644# diff_4915_3191# diff_2113_3589# GND efet w=29 l=17
+ ad=0 pd=0 as=0 ps=0 
M2447 diff_4987_3652# diff_4915_3191# diff_2053_3553# GND efet w=75 l=24
+ ad=0 pd=0 as=0 ps=0 
M2448 GND diff_5095_3556# diff_5116_3613# GND efet w=47 l=16
+ ad=0 pd=0 as=3248 ps=308 
M2449 GND diff_5095_3556# diff_5206_3742# GND efet w=28 l=16
+ ad=0 pd=0 as=1316 ps=150 
M2450 GND diff_5266_3691# diff_5278_3644# GND efet w=28 l=16
+ ad=0 pd=0 as=1316 ps=150 
M2451 GND diff_5266_3691# diff_5335_3644# GND efet w=40 l=16
+ ad=0 pd=0 as=3212 ps=296 
M2452 diff_5849_3703# Vdd Vdd GND efet w=25 l=67
+ ad=5736 pd=524 as=0 ps=0 
M2453 diff_5849_3703# diff_5849_3703# diff_5849_3703# GND efet w=4 l=10
+ ad=0 pd=0 as=0 ps=0 
M2454 diff_5849_3703# diff_5849_3703# diff_5849_3703# GND efet w=5 l=18
+ ad=0 pd=0 as=0 ps=0 
M2455 diff_2053_3553# diff_5029_3068# diff_5116_3613# GND efet w=79 l=24
+ ad=0 pd=0 as=0 ps=0 
M2456 diff_5206_3742# diff_5029_3068# diff_2113_3589# GND efet w=28 l=16
+ ad=0 pd=0 as=0 ps=0 
M2457 diff_5278_3644# diff_5134_2953# diff_2113_3589# GND efet w=28 l=16
+ ad=0 pd=0 as=0 ps=0 
M2458 diff_5335_3644# diff_5134_2953# diff_2053_3553# GND efet w=75 l=23
+ ad=0 pd=0 as=0 ps=0 
M2459 diff_1996_3562# diff_1996_3562# diff_1996_3562# GND efet w=10 l=16
+ ad=3267 pd=354 as=0 ps=0 
M2460 diff_1996_3562# diff_1996_3562# diff_1996_3562# GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M2461 GND diff_2026_2897# diff_1996_3562# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M2462 diff_2170_3691# diff_2170_3631# GND GND efet w=34 l=16
+ ad=3072 pd=342 as=0 ps=0 
M2463 diff_2170_3691# diff_2170_3691# diff_2170_3691# GND efet w=10 l=16
+ ad=0 pd=0 as=0 ps=0 
M2464 diff_2170_3691# diff_2170_3691# diff_2170_3691# GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M2465 Vdd Vdd diff_1996_3562# GND efet w=16 l=94
+ ad=0 pd=0 as=0 ps=0 
M2466 GND diff_1786_2191# diff_1829_3439# GND efet w=46 l=16
+ ad=0 pd=0 as=0 ps=0 
M2467 d3 GND GND GND efet w=256 l=19
+ ad=0 pd=0 as=0 ps=0 
M2468 diff_580_3394# diff_425_3187# Vdd GND efet w=94 l=16
+ ad=0 pd=0 as=0 ps=0 
M2469 diff_2026_2897# diff_2026_2897# diff_2026_2897# GND efet w=5 l=5
+ ad=11418 pd=1152 as=0 ps=0 
M2470 diff_829_3778# diff_1291_3346# GND GND efet w=61 l=16
+ ad=0 pd=0 as=0 ps=0 
M2471 diff_817_6145# diff_1291_3346# GND GND efet w=61 l=16
+ ad=0 pd=0 as=0 ps=0 
M2472 diff_425_3187# diff_407_3110# GND GND efet w=55 l=16
+ ad=8522 pd=690 as=0 ps=0 
M2473 diff_425_3187# diff_425_3187# diff_425_3187# GND efet w=4 l=4
+ ad=0 pd=0 as=0 ps=0 
M2474 diff_425_3187# diff_425_3187# diff_425_3187# GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M2475 Vdd Vdd diff_425_3187# GND efet w=19 l=89
+ ad=0 pd=0 as=0 ps=0 
M2476 diff_2026_2897# diff_2026_2897# diff_2026_2897# GND efet w=5 l=10
+ ad=0 pd=0 as=0 ps=0 
M2477 diff_2344_3556# diff_2344_3556# diff_2344_3556# GND efet w=10 l=13
+ ad=3216 pd=342 as=0 ps=0 
M2478 diff_2344_3556# diff_2344_3556# diff_2344_3556# GND efet w=10 l=6
+ ad=0 pd=0 as=0 ps=0 
M2479 GND diff_2368_2803# diff_2344_3556# GND efet w=34 l=19
+ ad=0 pd=0 as=0 ps=0 
M2480 diff_2515_3691# diff_2515_3628# GND GND efet w=40 l=16
+ ad=3138 pd=354 as=0 ps=0 
M2481 diff_2515_3691# diff_2515_3691# diff_2515_3691# GND efet w=10 l=13
+ ad=0 pd=0 as=0 ps=0 
M2482 diff_2515_3691# diff_2515_3691# diff_2515_3691# GND efet w=10 l=6
+ ad=0 pd=0 as=0 ps=0 
M2483 Vdd Vdd diff_2170_3691# GND efet w=20 l=124
+ ad=0 pd=0 as=0 ps=0 
M2484 diff_2344_3556# Vdd Vdd GND efet w=20 l=111
+ ad=0 pd=0 as=0 ps=0 
M2485 diff_2170_3631# diff_2170_3631# diff_2170_3631# GND efet w=4 l=7
+ ad=11873 pd=1120 as=0 ps=0 
M2486 diff_2170_3631# diff_2170_3631# diff_2170_3631# GND efet w=7 l=8
+ ad=0 pd=0 as=0 ps=0 
M2487 diff_2368_2803# diff_2368_2803# diff_2368_2803# GND efet w=5 l=5
+ ad=10775 pd=1216 as=0 ps=0 
M2488 diff_2368_2803# diff_2368_2803# diff_2368_2803# GND efet w=5 l=13
+ ad=0 pd=0 as=0 ps=0 
M2489 diff_2689_3475# diff_2689_3475# diff_2689_3475# GND efet w=10 l=16
+ ad=3279 pd=354 as=0 ps=0 
M2490 diff_2689_3475# diff_2689_3475# diff_2689_3475# GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M2491 GND diff_2713_2900# diff_2689_3475# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M2492 diff_2857_3691# diff_2857_3628# GND GND efet w=34 l=16
+ ad=3159 pd=348 as=0 ps=0 
M2493 diff_2857_3691# diff_2857_3691# diff_2857_3691# GND efet w=10 l=16
+ ad=0 pd=0 as=0 ps=0 
M2494 diff_3031_3556# diff_3031_3556# diff_3031_3556# GND efet w=10 l=16
+ ad=3177 pd=342 as=0 ps=0 
M2495 diff_2857_3691# diff_2857_3691# diff_2857_3691# GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M2496 Vdd Vdd diff_2515_3691# GND efet w=20 l=117
+ ad=0 pd=0 as=0 ps=0 
M2497 diff_2689_3475# Vdd Vdd GND efet w=20 l=117
+ ad=0 pd=0 as=0 ps=0 
M2498 diff_2515_3628# diff_2515_3628# diff_2515_3628# GND efet w=4 l=5
+ ad=11462 pd=1114 as=0 ps=0 
M2499 diff_2515_3628# diff_2515_3628# diff_2515_3628# GND efet w=8 l=8
+ ad=0 pd=0 as=0 ps=0 
M2500 diff_2713_2900# diff_2713_2900# diff_2713_2900# GND efet w=7 l=7
+ ad=11316 pd=1152 as=0 ps=0 
M2501 diff_2713_2900# diff_2713_2900# diff_2713_2900# GND efet w=5 l=10
+ ad=0 pd=0 as=0 ps=0 
M2502 GND diff_3055_2897# diff_3031_3556# GND efet w=37 l=16
+ ad=0 pd=0 as=0 ps=0 
M2503 diff_3031_3556# diff_3031_3556# diff_3031_3556# GND efet w=10 l=6
+ ad=0 pd=0 as=0 ps=0 
M2504 diff_3202_3691# diff_3202_3628# GND GND efet w=34 l=16
+ ad=3174 pd=348 as=0 ps=0 
M2505 diff_3202_3691# diff_3202_3691# diff_3202_3691# GND efet w=10 l=16
+ ad=0 pd=0 as=0 ps=0 
M2506 diff_3202_3691# diff_3202_3691# diff_3202_3691# GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M2507 diff_2857_3691# Vdd Vdd GND efet w=22 l=115
+ ad=0 pd=0 as=0 ps=0 
M2508 diff_3031_3556# Vdd Vdd GND efet w=23 l=115
+ ad=0 pd=0 as=0 ps=0 
M2509 diff_2857_3628# diff_2857_3628# diff_2857_3628# GND efet w=4 l=7
+ ad=11645 pd=1090 as=0 ps=0 
M2510 diff_2857_3628# diff_2857_3628# diff_2857_3628# GND efet w=8 l=8
+ ad=0 pd=0 as=0 ps=0 
M2511 diff_3055_2897# diff_3055_2897# diff_3055_2897# GND efet w=5 l=5
+ ad=11229 pd=1158 as=0 ps=0 
M2512 diff_3055_2897# diff_3055_2897# diff_3055_2897# GND efet w=6 l=13
+ ad=0 pd=0 as=0 ps=0 
M2513 diff_3376_3475# diff_3376_3475# diff_3376_3475# GND efet w=11 l=14
+ ad=3246 pd=366 as=0 ps=0 
M2514 GND diff_3400_2897# diff_3376_3475# GND efet w=41 l=17
+ ad=0 pd=0 as=0 ps=0 
M2515 diff_3544_3691# diff_3544_3628# GND GND efet w=40 l=17
+ ad=3183 pd=342 as=0 ps=0 
M2516 diff_3544_3691# diff_3544_3691# diff_3544_3691# GND efet w=10 l=13
+ ad=0 pd=0 as=0 ps=0 
M2517 diff_3376_3475# diff_3376_3475# diff_3376_3475# GND efet w=10 l=6
+ ad=0 pd=0 as=0 ps=0 
M2518 diff_3544_3691# diff_3544_3691# diff_3544_3691# GND efet w=10 l=6
+ ad=0 pd=0 as=0 ps=0 
M2519 Vdd Vdd diff_3202_3691# GND efet w=20 l=114
+ ad=0 pd=0 as=0 ps=0 
M2520 diff_3376_3475# Vdd Vdd GND efet w=20 l=112
+ ad=0 pd=0 as=0 ps=0 
M2521 diff_3202_3628# diff_3202_3628# diff_3202_3628# GND efet w=4 l=5
+ ad=11369 pd=1102 as=0 ps=0 
M2522 diff_3202_3628# diff_3202_3628# diff_3202_3628# GND efet w=8 l=8
+ ad=0 pd=0 as=0 ps=0 
M2523 diff_3400_2897# diff_3400_2897# diff_3400_2897# GND efet w=4 l=7
+ ad=11319 pd=1140 as=0 ps=0 
M2524 diff_3400_2897# diff_3400_2897# diff_3400_2897# GND efet w=5 l=10
+ ad=0 pd=0 as=0 ps=0 
M2525 diff_3718_3556# diff_3718_3556# diff_3718_3556# GND efet w=10 l=16
+ ad=3156 pd=348 as=0 ps=0 
M2526 GND diff_3745_2897# diff_3718_3556# GND efet w=37 l=16
+ ad=0 pd=0 as=0 ps=0 
M2527 diff_3889_3691# diff_3889_3628# GND GND efet w=37 l=16
+ ad=3165 pd=348 as=0 ps=0 
M2528 diff_3718_3556# diff_3718_3556# diff_3718_3556# GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M2529 diff_3889_3691# diff_3889_3691# diff_3889_3691# GND efet w=10 l=16
+ ad=0 pd=0 as=0 ps=0 
M2530 diff_4063_3493# diff_4063_3493# diff_4063_3493# GND efet w=10 l=16
+ ad=3195 pd=354 as=0 ps=0 
M2531 diff_3889_3691# diff_3889_3691# diff_3889_3691# GND efet w=10 l=6
+ ad=0 pd=0 as=0 ps=0 
M2532 diff_4063_3493# diff_4063_3493# diff_4063_3493# GND efet w=10 l=6
+ ad=0 pd=0 as=0 ps=0 
M2533 GND diff_4087_2900# diff_4063_3493# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M2534 diff_4231_3691# diff_4231_3628# GND GND efet w=34 l=16
+ ad=3174 pd=348 as=0 ps=0 
M2535 diff_4231_3691# diff_4231_3691# diff_4231_3691# GND efet w=10 l=16
+ ad=0 pd=0 as=0 ps=0 
M2536 diff_4231_3691# diff_4231_3691# diff_4231_3691# GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M2537 Vdd Vdd diff_3544_3691# GND efet w=19 l=115
+ ad=0 pd=0 as=0 ps=0 
M2538 diff_3544_3628# diff_3544_3628# diff_3544_3628# GND efet w=5 l=5
+ ad=11726 pd=1094 as=0 ps=0 
M2539 diff_3544_3628# diff_3544_3628# diff_3544_3628# GND efet w=7 l=7
+ ad=0 pd=0 as=0 ps=0 
M2540 diff_3718_3556# Vdd Vdd GND efet w=21 l=119
+ ad=0 pd=0 as=0 ps=0 
M2541 diff_3745_2897# diff_3745_2897# diff_3745_2897# GND efet w=5 l=5
+ ad=10433 pd=1042 as=0 ps=0 
M2542 diff_3745_2897# diff_3745_2897# diff_3745_2897# GND efet w=4 l=7
+ ad=0 pd=0 as=0 ps=0 
M2543 Vdd Vdd diff_3889_3691# GND efet w=21 l=116
+ ad=0 pd=0 as=0 ps=0 
M2544 diff_3889_3628# diff_3889_3628# diff_3889_3628# GND efet w=4 l=5
+ ad=11762 pd=1284 as=0 ps=0 
M2545 diff_3889_3628# diff_3889_3628# diff_3889_3628# GND efet w=8 l=9
+ ad=0 pd=0 as=0 ps=0 
M2546 diff_4063_3493# Vdd Vdd GND efet w=17 l=115
+ ad=0 pd=0 as=0 ps=0 
M2547 diff_4087_2900# diff_4087_2900# diff_4087_2900# GND efet w=5 l=5
+ ad=11460 pd=1170 as=0 ps=0 
M2548 diff_4087_2900# diff_4087_2900# diff_4087_2900# GND efet w=5 l=10
+ ad=0 pd=0 as=0 ps=0 
M2549 diff_4405_3556# diff_4405_3556# diff_4405_3556# GND efet w=10 l=13
+ ad=3201 pd=342 as=0 ps=0 
M2550 diff_4405_3556# diff_4405_3556# diff_4405_3556# GND efet w=10 l=6
+ ad=0 pd=0 as=0 ps=0 
M2551 GND diff_4399_2803# diff_4405_3556# GND efet w=34 l=19
+ ad=0 pd=0 as=0 ps=0 
M2552 diff_4576_3691# diff_4552_2860# GND GND efet w=38 l=17
+ ad=3210 pd=342 as=0 ps=0 
M2553 diff_4576_3691# diff_4576_3691# diff_4576_3691# GND efet w=10 l=13
+ ad=0 pd=0 as=0 ps=0 
M2554 diff_4576_3691# diff_4576_3691# diff_4576_3691# GND efet w=10 l=6
+ ad=0 pd=0 as=0 ps=0 
M2555 Vdd Vdd diff_4231_3691# GND efet w=20 l=114
+ ad=0 pd=0 as=0 ps=0 
M2556 diff_4231_3628# diff_4231_3628# diff_4231_3628# GND efet w=2 l=8
+ ad=12905 pd=1302 as=0 ps=0 
M2557 diff_4231_3628# diff_4231_3628# diff_4231_3628# GND efet w=7 l=7
+ ad=0 pd=0 as=0 ps=0 
M2558 diff_4405_3556# Vdd Vdd GND efet w=19 l=112
+ ad=0 pd=0 as=0 ps=0 
M2559 diff_4399_2803# diff_4399_2803# diff_4399_2803# GND efet w=7 l=10
+ ad=13371 pd=1370 as=0 ps=0 
M2560 diff_4399_2803# diff_4399_2803# diff_4399_2803# GND efet w=3 l=8
+ ad=0 pd=0 as=0 ps=0 
M2561 diff_4750_3556# diff_4750_3556# diff_4750_3556# GND efet w=10 l=16
+ ad=3285 pd=354 as=0 ps=0 
M2562 diff_4750_3556# diff_4750_3556# diff_4750_3556# GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M2563 GND diff_4732_2900# diff_4750_3556# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M2564 diff_4921_3691# diff_4915_3191# GND GND efet w=34 l=16
+ ad=3159 pd=348 as=0 ps=0 
M2565 diff_4921_3691# diff_4921_3691# diff_4921_3691# GND efet w=10 l=13
+ ad=0 pd=0 as=0 ps=0 
M2566 diff_5095_3556# diff_5095_3556# diff_5095_3556# GND efet w=10 l=16
+ ad=3183 pd=348 as=0 ps=0 
M2567 diff_4921_3691# diff_4921_3691# diff_4921_3691# GND efet w=10 l=6
+ ad=0 pd=0 as=0 ps=0 
M2568 Vdd Vdd diff_4576_3691# GND efet w=20 l=115
+ ad=0 pd=0 as=0 ps=0 
M2569 diff_4750_3556# Vdd Vdd GND efet w=20 l=114
+ ad=0 pd=0 as=0 ps=0 
M2570 diff_4552_2860# diff_4552_2860# diff_4552_2860# GND efet w=2 l=4
+ ad=14136 pd=1492 as=0 ps=0 
M2571 diff_4552_2860# diff_4552_2860# diff_4552_2860# GND efet w=7 l=7
+ ad=0 pd=0 as=0 ps=0 
M2572 diff_2026_2897# diff_2062_3349# GND GND efet w=37 l=17
+ ad=0 pd=0 as=0 ps=0 
M2573 diff_2170_3631# diff_2062_3349# GND GND efet w=40 l=19
+ ad=0 pd=0 as=0 ps=0 
M2574 diff_2368_2803# diff_2062_3349# GND GND efet w=38 l=20
+ ad=0 pd=0 as=0 ps=0 
M2575 diff_2515_3628# diff_2062_3349# GND GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2576 diff_2713_2900# diff_2062_3349# GND GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2577 diff_2857_3628# diff_2062_3349# GND GND efet w=38 l=20
+ ad=0 pd=0 as=0 ps=0 
M2578 diff_3055_2897# diff_2062_3349# GND GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2579 diff_3202_3628# diff_2062_3349# GND GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2580 diff_3400_2897# diff_3254_2623# GND GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2581 diff_3544_3628# diff_3254_2623# GND GND efet w=38 l=20
+ ad=0 pd=0 as=0 ps=0 
M2582 diff_3745_2897# diff_3254_2623# GND GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2583 diff_3889_3628# diff_3254_2623# GND GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2584 GND diff_3254_2623# diff_4087_2900# GND efet w=40 l=19
+ ad=0 pd=0 as=0 ps=0 
M2585 diff_4231_3628# diff_3254_2623# GND GND efet w=37 l=16
+ ad=0 pd=0 as=0 ps=0 
M2586 diff_4399_2803# diff_3254_2623# GND GND efet w=40 l=16
+ ad=0 pd=0 as=0 ps=0 
M2587 diff_4552_2860# diff_3254_2623# GND GND efet w=37 l=16
+ ad=0 pd=0 as=0 ps=0 
M2588 diff_5095_3556# diff_5095_3556# diff_5095_3556# GND efet w=12 l=8
+ ad=0 pd=0 as=0 ps=0 
M2589 GND diff_5029_3068# diff_5095_3556# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M2590 diff_5849_3703# diff_673_1115# diff_5875_3626# GND efet w=170 l=14
+ ad=0 pd=0 as=6299 ps=500 
M2591 diff_5875_3626# diff_1960_562# GND GND efet w=178 l=14
+ ad=0 pd=0 as=0 ps=0 
M2592 diff_5266_3691# diff_5266_3691# diff_5266_3691# GND efet w=2 l=4
+ ad=3444 pd=482 as=0 ps=0 
M2593 Vdd Vdd diff_4921_3691# GND efet w=17 l=113
+ ad=0 pd=0 as=0 ps=0 
M2594 diff_5095_3556# Vdd Vdd GND efet w=21 l=115
+ ad=0 pd=0 as=0 ps=0 
M2595 diff_5266_3691# diff_5266_3691# diff_5266_3691# GND efet w=4 l=4
+ ad=0 pd=0 as=0 ps=0 
M2596 diff_2053_3553# diff_5776_3412# Vdd GND efet w=94 l=19
+ ad=0 pd=0 as=0 ps=0 
M2597 GND diff_1291_3280# diff_820_3511# GND efet w=61 l=16
+ ad=0 pd=0 as=0 ps=0 
M2598 GND diff_1291_3280# diff_1093_4033# GND efet w=61 l=16
+ ad=0 pd=0 as=0 ps=0 
M2599 diff_1309_3670# diff_550_2356# Vdd GND efet w=71 l=16
+ ad=8967 pd=634 as=0 ps=0 
M2600 GND diff_1829_3133# diff_1309_3670# GND efet w=67 l=16
+ ad=0 pd=0 as=0 ps=0 
M2601 GND diff_2056_3301# diff_2026_2897# GND efet w=40 l=19
+ ad=0 pd=0 as=0 ps=0 
M2602 GND diff_2056_3301# diff_2170_3631# GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2603 GND diff_2056_3301# diff_2368_2803# GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2604 GND diff_2056_3301# diff_2515_3628# GND efet w=41 l=17
+ ad=0 pd=0 as=0 ps=0 
M2605 GND diff_2056_3301# diff_3400_2897# GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2606 GND diff_2056_3301# diff_3544_3628# GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2607 GND diff_2056_3301# diff_3745_2897# GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2608 GND diff_2056_3301# diff_3889_3628# GND efet w=38 l=17
+ ad=0 pd=0 as=0 ps=0 
M2609 diff_5266_3691# diff_5134_2953# GND GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M2610 Vdd Vdd diff_5266_3691# GND efet w=14 l=110
+ ad=0 pd=0 as=0 ps=0 
M2611 GND diff_5837_3124# diff_2053_3553# GND efet w=107 l=13
+ ad=0 pd=0 as=0 ps=0 
M2612 GND diff_5837_3124# diff_5776_3412# GND efet w=100 l=16
+ ad=0 pd=0 as=9542 ps=948 
M2613 diff_5134_2953# diff_5191_3280# diff_5134_2953# GND efet w=207 l=8
+ ad=12340 pd=1428 as=0 ps=0 
M2614 diff_2713_2900# diff_2743_3241# GND GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2615 diff_2857_3628# diff_2743_3241# GND GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2616 diff_3055_2897# diff_2743_3241# GND GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2617 diff_3202_3628# diff_2743_3241# GND GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2618 diff_4087_2900# diff_2743_3241# GND GND efet w=38 l=17
+ ad=0 pd=0 as=0 ps=0 
M2619 diff_4231_3628# diff_2743_3241# GND GND efet w=41 l=17
+ ad=0 pd=0 as=0 ps=0 
M2620 diff_820_3511# diff_1291_3169# GND GND efet w=61 l=16
+ ad=0 pd=0 as=0 ps=0 
M2621 diff_817_6145# diff_1291_3169# GND GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M2622 diff_425_3187# diff_331_7000# GND GND efet w=88 l=16
+ ad=0 pd=0 as=0 ps=0 
M2623 diff_407_3110# diff_407_3110# diff_407_3110# GND efet w=5 l=15
+ ad=7394 pd=724 as=0 ps=0 
M2624 diff_407_3110# diff_407_3110# diff_407_3110# GND efet w=5 l=13
+ ad=0 pd=0 as=0 ps=0 
M2625 diff_407_3110# d3 GND GND efet w=136 l=16
+ ad=0 pd=0 as=0 ps=0 
M2626 diff_1829_3133# Vdd Vdd GND efet w=19 l=95
+ ad=2261 pd=228 as=0 ps=0 
M2627 diff_2026_2897# diff_2056_3184# GND GND efet w=41 l=17
+ ad=0 pd=0 as=0 ps=0 
M2628 diff_4399_2803# diff_2743_3241# GND GND efet w=37 l=16
+ ad=0 pd=0 as=0 ps=0 
M2629 diff_4552_2860# diff_2743_3241# GND GND efet w=37 l=17
+ ad=0 pd=0 as=0 ps=0 
M2630 Vdd diff_5191_3280# diff_5134_2953# GND efet w=19 l=88
+ ad=0 pd=0 as=0 ps=0 
M2631 diff_5191_3280# diff_5191_3280# diff_5191_3280# GND efet w=2 l=7
+ ad=1471 pd=190 as=0 ps=0 
M2632 diff_5191_3280# diff_5191_3280# diff_5191_3280# GND efet w=4 l=8
+ ad=0 pd=0 as=0 ps=0 
M2633 Vdd Vdd diff_5191_3280# GND efet w=19 l=16
+ ad=0 pd=0 as=0 ps=0 
M2634 diff_5776_3412# diff_5762_3178# Vdd GND efet w=22 l=46
+ ad=0 pd=0 as=0 ps=0 
M2635 diff_4732_2900# diff_4756_3238# GND GND efet w=49 l=17
+ ad=11221 pd=964 as=0 ps=0 
M2636 diff_2170_3631# diff_2056_3184# GND GND efet w=37 l=16
+ ad=0 pd=0 as=0 ps=0 
M2637 GND diff_2056_3184# diff_2713_2900# GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2638 GND diff_550_2356# diff_1829_3133# GND efet w=47 l=20
+ ad=0 pd=0 as=0 ps=0 
M2639 GND diff_1291_3103# diff_829_3778# GND efet w=61 l=16
+ ad=0 pd=0 as=0 ps=0 
M2640 GND diff_1291_3103# diff_1093_4033# GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M2641 GND diff_2056_3184# diff_2857_3628# GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2642 diff_5134_2953# diff_4756_3238# GND GND efet w=46 l=19
+ ad=0 pd=0 as=0 ps=0 
M2643 diff_3400_2897# diff_2056_3184# GND GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2644 diff_3544_3628# diff_2056_3184# GND GND efet w=41 l=17
+ ad=0 pd=0 as=0 ps=0 
M2645 GND diff_2056_3184# diff_4087_2900# GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2646 GND diff_2056_3184# diff_4231_3628# GND efet w=41 l=17
+ ad=0 pd=0 as=0 ps=0 
M2647 diff_5776_3412# diff_5762_3178# diff_5776_3412# GND efet w=132 l=26
+ ad=0 pd=0 as=0 ps=0 
M2648 diff_5762_3178# diff_5762_3178# diff_5762_3178# GND efet w=5 l=5
+ ad=1477 pd=190 as=0 ps=0 
M2649 diff_5762_3178# diff_5762_3178# diff_5762_3178# GND efet w=3 l=16
+ ad=0 pd=0 as=0 ps=0 
M2650 diff_4915_3191# diff_4903_3178# GND GND efet w=76 l=16
+ ad=11017 pd=1200 as=0 ps=0 
M2651 GND diff_4903_3178# diff_5029_3068# GND efet w=79 l=16
+ ad=0 pd=0 as=12829 ps=1242 
M2652 diff_5762_3178# Vdd Vdd GND efet w=20 l=19
+ ad=0 pd=0 as=0 ps=0 
M2653 GND diff_2101_2551# diff_2368_2803# GND efet w=37 l=17
+ ad=0 pd=0 as=0 ps=0 
M2654 GND diff_2101_2551# diff_2515_3628# GND efet w=40 l=19
+ ad=0 pd=0 as=0 ps=0 
M2655 diff_3055_2897# diff_2101_2551# GND GND efet w=38 l=20
+ ad=0 pd=0 as=0 ps=0 
M2656 diff_3202_3628# diff_2101_2551# GND GND efet w=38 l=20
+ ad=0 pd=0 as=0 ps=0 
M2657 GND diff_2101_2551# diff_3745_2897# GND efet w=40 l=22
+ ad=0 pd=0 as=0 ps=0 
M2658 GND diff_2101_2551# diff_3889_3628# GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2659 diff_4399_2803# diff_2101_2551# GND GND efet w=38 l=16
+ ad=0 pd=0 as=0 ps=0 
M2660 diff_4552_2860# diff_2101_2551# GND GND efet w=37 l=16
+ ad=0 pd=0 as=0 ps=0 
M2661 GND diff_331_7000# diff_407_3110# GND efet w=88 l=16
+ ad=0 pd=0 as=0 ps=0 
M2662 diff_2026_2897# diff_2056_3070# GND GND efet w=37 l=16
+ ad=0 pd=0 as=0 ps=0 
M2663 diff_2368_2803# diff_2056_3070# GND GND efet w=37 l=16
+ ad=0 pd=0 as=0 ps=0 
M2664 diff_2713_2900# diff_2056_3070# GND GND efet w=41 l=17
+ ad=0 pd=0 as=0 ps=0 
M2665 GND diff_2056_3070# diff_3055_2897# GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2666 diff_3400_2897# diff_2056_3070# GND GND efet w=37 l=19
+ ad=0 pd=0 as=0 ps=0 
M2667 GND diff_4936_3115# diff_4915_3191# GND efet w=46 l=19
+ ad=0 pd=0 as=0 ps=0 
M2668 GND diff_4936_3115# diff_5134_2953# GND efet w=46 l=19
+ ad=0 pd=0 as=0 ps=0 
M2669 diff_5837_3124# Vdd Vdd GND efet w=25 l=46
+ ad=5453 pd=460 as=0 ps=0 
M2670 diff_3745_2897# diff_2056_3070# GND GND efet w=44 l=22
+ ad=0 pd=0 as=0 ps=0 
M2671 Vdd Vdd Vdd GND efet w=2 l=13
+ ad=0 pd=0 as=0 ps=0 
M2672 Vdd Vdd Vdd GND efet w=9 l=16
+ ad=0 pd=0 as=0 ps=0 
M2673 Vdd Vdd diff_407_3110# GND efet w=20 l=89
+ ad=0 pd=0 as=0 ps=0 
M2674 diff_2515_3628# diff_2209_3019# GND GND efet w=41 l=17
+ ad=0 pd=0 as=0 ps=0 
M2675 GND diff_2209_3019# diff_2857_3628# GND efet w=43 l=16
+ ad=0 pd=0 as=0 ps=0 
M2676 diff_4087_2900# diff_2056_3070# GND GND efet w=46 l=19
+ ad=0 pd=0 as=0 ps=0 
M2677 GND diff_2056_3070# diff_4399_2803# GND efet w=38 l=17
+ ad=0 pd=0 as=0 ps=0 
M2678 diff_5837_3124# clk2 diff_5848_3025# GND efet w=178 l=16
+ ad=0 pd=0 as=9059 ps=650 
M2679 GND diff_5771_2965# diff_5848_3025# GND efet w=280 l=16
+ ad=0 pd=0 as=0 ps=0 
M2680 diff_4732_2900# diff_4723_3052# GND GND efet w=79 l=16
+ ad=0 pd=0 as=0 ps=0 
M2681 diff_5029_3068# diff_4723_3052# GND GND efet w=79 l=16
+ ad=0 pd=0 as=0 ps=0 
M2682 GND diff_2209_3019# diff_3889_3628# GND efet w=40 l=16
+ ad=0 pd=0 as=0 ps=0 
M2683 GND diff_2209_3019# diff_2170_3631# GND efet w=37 l=16
+ ad=0 pd=0 as=0 ps=0 
M2684 GND diff_2209_3019# diff_3202_3628# GND efet w=37 l=16
+ ad=0 pd=0 as=0 ps=0 
M2685 GND diff_2209_3019# diff_3544_3628# GND efet w=38 l=17
+ ad=0 pd=0 as=0 ps=0 
M2686 diff_4231_3628# diff_2209_3019# GND GND efet w=38 l=17
+ ad=0 pd=0 as=0 ps=0 
M2687 diff_4552_2860# diff_2209_3019# GND GND efet w=37 l=16
+ ad=0 pd=0 as=0 ps=0 
M2688 diff_220_5722# diff_550_2755# GND GND efet w=163 l=16
+ ad=9128 pd=438 as=0 ps=0 
M2689 Vdd diff_622_2720# diff_220_5722# GND efet w=172 l=16
+ ad=0 pd=0 as=0 ps=0 
M2690 diff_1291_3280# diff_1291_3346# GND GND efet w=46 l=16
+ ad=4990 pd=364 as=0 ps=0 
M2691 Vdd Vdd diff_1291_3280# GND efet w=26 l=116
+ ad=0 pd=0 as=0 ps=0 
M2692 diff_1291_3280# diff_1417_2311# diff_1436_2722# GND efet w=19 l=16
+ ad=0 pd=0 as=3940 ps=396 
M2693 diff_2026_2897# diff_2023_2797# diff_2026_2897# GND efet w=79 l=118
+ ad=0 pd=0 as=0 ps=0 
M2694 diff_550_2755# diff_550_2755# diff_550_2755# GND efet w=5 l=15
+ ad=1240 pd=152 as=0 ps=0 
M2695 diff_550_2755# diff_550_2755# diff_550_2755# GND efet w=2 l=15
+ ad=0 pd=0 as=0 ps=0 
M2696 diff_622_2720# diff_622_2720# diff_622_2720# GND efet w=5 l=11
+ ad=1309 pd=164 as=0 ps=0 
M2697 diff_622_2720# diff_622_2720# diff_622_2720# GND efet w=5 l=14
+ ad=0 pd=0 as=0 ps=0 
M2698 diff_872_2743# diff_508_1279# Vdd GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2699 diff_1291_3346# diff_1436_2722# GND GND efet w=79 l=16
+ ad=6782 pd=576 as=0 ps=0 
M2700 Vdd Vdd diff_1291_3346# GND efet w=25 l=115
+ ad=0 pd=0 as=0 ps=0 
M2701 diff_2170_3631# diff_2176_2758# diff_2170_3631# GND efet w=76 l=121
+ ad=0 pd=0 as=0 ps=0 
M2702 diff_550_2755# diff_556_2707# diff_562_2665# GND efet w=35 l=14
+ ad=0 pd=0 as=6620 ps=524 
M2703 diff_622_2720# diff_556_2707# diff_550_2479# GND efet w=34 l=19
+ ad=0 pd=0 as=4985 ps=456 
M2704 diff_1436_2722# diff_1405_2629# diff_872_2743# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M2705 diff_1436_2722# diff_1436_2722# diff_1436_2722# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M2706 diff_1436_2722# diff_1436_2722# diff_1436_2722# GND efet w=3 l=7
+ ad=0 pd=0 as=0 ps=0 
M2707 diff_2023_2797# diff_2023_2797# diff_2023_2797# GND efet w=5 l=5
+ ad=1144 pd=166 as=0 ps=0 
M2708 diff_2023_2797# diff_2023_2797# diff_2023_2797# GND efet w=3 l=7
+ ad=0 pd=0 as=0 ps=0 
M2709 diff_2026_2897# diff_2023_2797# Vdd GND efet w=19 l=91
+ ad=0 pd=0 as=0 ps=0 
M2710 diff_2170_3631# diff_2176_2758# Vdd GND efet w=19 l=91
+ ad=0 pd=0 as=0 ps=0 
M2711 diff_2176_2758# diff_2176_2758# diff_2176_2758# GND efet w=5 l=5
+ ad=1168 pd=166 as=0 ps=0 
M2712 diff_2023_2797# Vdd Vdd GND efet w=16 l=16
+ ad=0 pd=0 as=0 ps=0 
M2713 diff_562_2665# diff_550_2479# GND GND efet w=124 l=16
+ ad=0 pd=0 as=0 ps=0 
M2714 diff_629_6919# diff_508_1279# Vdd GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2715 diff_1436_2665# diff_1405_2629# diff_629_6919# GND efet w=31 l=16
+ ad=3706 pd=396 as=0 ps=0 
M2716 diff_1436_2665# diff_1436_2665# diff_1436_2665# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M2717 diff_1436_2665# diff_1436_2665# diff_1436_2665# GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M2718 diff_2176_2758# diff_2176_2758# diff_2176_2758# GND efet w=3 l=7
+ ad=0 pd=0 as=0 ps=0 
M2719 diff_2176_2758# Vdd Vdd GND efet w=19 l=16
+ ad=0 pd=0 as=0 ps=0 
M2720 Vdd Vdd diff_2101_2551# GND efet w=23 l=70
+ ad=0 pd=0 as=12845 ps=1580 
M2721 Vdd Vdd diff_562_2665# GND efet w=25 l=46
+ ad=0 pd=0 as=0 ps=0 
M2722 diff_577_5317# diff_508_1279# Vdd GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M2723 diff_1291_3169# diff_1436_2665# GND GND efet w=79 l=16
+ ad=6794 pd=564 as=0 ps=0 
M2724 Vdd Vdd diff_1291_3169# GND efet w=25 l=115
+ ad=0 pd=0 as=0 ps=0 
M2725 GND diff_2062_2569# diff_2101_2551# GND efet w=122 l=17
+ ad=0 pd=0 as=0 ps=0 
M2726 diff_2368_2803# diff_2371_2794# diff_2368_2803# GND efet w=124 l=68
+ ad=0 pd=0 as=0 ps=0 
M2727 diff_2515_3628# diff_2521_2758# diff_2515_3628# GND efet w=74 l=116
+ ad=0 pd=0 as=0 ps=0 
M2728 diff_2371_2794# diff_2371_2794# diff_2371_2794# GND efet w=5 l=5
+ ad=1213 pd=180 as=0 ps=0 
M2729 diff_2371_2794# diff_2371_2794# diff_2371_2794# GND efet w=4 l=8
+ ad=0 pd=0 as=0 ps=0 
M2730 diff_2368_2803# diff_2371_2794# Vdd GND efet w=19 l=91
+ ad=0 pd=0 as=0 ps=0 
M2731 diff_2515_3628# diff_2521_2758# Vdd GND efet w=19 l=91
+ ad=0 pd=0 as=0 ps=0 
M2732 diff_2521_2758# diff_2521_2758# diff_2521_2758# GND efet w=5 l=5
+ ad=1231 pd=180 as=0 ps=0 
M2733 diff_2521_2758# diff_2521_2758# diff_2521_2758# GND efet w=4 l=8
+ ad=0 pd=0 as=0 ps=0 
M2734 diff_2371_2794# Vdd Vdd GND efet w=20 l=17
+ ad=0 pd=0 as=0 ps=0 
M2735 diff_2521_2758# Vdd Vdd GND efet w=19 l=19
+ ad=0 pd=0 as=0 ps=0 
M2736 diff_2056_3184# Vdd Vdd GND efet w=19 l=76
+ ad=8474 pd=1038 as=0 ps=0 
M2737 diff_2713_2900# diff_2710_2797# diff_2713_2900# GND efet w=74 l=118
+ ad=0 pd=0 as=0 ps=0 
M2738 diff_2857_3628# diff_2863_2758# diff_2857_3628# GND efet w=76 l=115
+ ad=0 pd=0 as=0 ps=0 
M2739 diff_2710_2797# diff_2710_2797# diff_2710_2797# GND efet w=5 l=5
+ ad=1126 pd=172 as=0 ps=0 
M2740 diff_2710_2797# diff_2710_2797# diff_2710_2797# GND efet w=3 l=7
+ ad=0 pd=0 as=0 ps=0 
M2741 diff_2713_2900# diff_2710_2797# Vdd GND efet w=19 l=91
+ ad=0 pd=0 as=0 ps=0 
M2742 diff_2857_3628# diff_2863_2758# Vdd GND efet w=19 l=91
+ ad=0 pd=0 as=0 ps=0 
M2743 diff_2863_2758# diff_2863_2758# diff_2863_2758# GND efet w=5 l=5
+ ad=1120 pd=166 as=0 ps=0 
M2744 diff_2710_2797# Vdd Vdd GND efet w=19 l=20
+ ad=0 pd=0 as=0 ps=0 
M2745 diff_2863_2758# diff_2863_2758# diff_2863_2758# GND efet w=3 l=7
+ ad=0 pd=0 as=0 ps=0 
M2746 diff_2863_2758# Vdd Vdd GND efet w=20 l=17
+ ad=0 pd=0 as=0 ps=0 
M2747 diff_3055_2897# diff_3055_2803# diff_3055_2897# GND efet w=79 l=84
+ ad=0 pd=0 as=0 ps=0 
M2748 diff_3202_3628# diff_3205_2761# diff_3202_3628# GND efet w=77 l=68
+ ad=0 pd=0 as=0 ps=0 
M2749 diff_3400_2897# diff_3397_2791# diff_3400_2897# GND efet w=77 l=115
+ ad=0 pd=0 as=0 ps=0 
M2750 diff_3055_2803# diff_3055_2803# diff_3055_2803# GND efet w=5 l=5
+ ad=1171 pd=172 as=0 ps=0 
M2751 diff_3055_2803# diff_3055_2803# diff_3055_2803# GND efet w=3 l=7
+ ad=0 pd=0 as=0 ps=0 
M2752 diff_3055_2897# diff_3055_2803# Vdd GND efet w=19 l=91
+ ad=0 pd=0 as=0 ps=0 
M2753 diff_3202_3628# diff_3205_2761# Vdd GND efet w=19 l=91
+ ad=0 pd=0 as=0 ps=0 
M2754 diff_3205_2761# diff_3205_2761# diff_3205_2761# GND efet w=5 l=5
+ ad=1213 pd=168 as=0 ps=0 
M2755 diff_3205_2761# diff_3205_2761# diff_3205_2761# GND efet w=2 l=8
+ ad=0 pd=0 as=0 ps=0 
M2756 diff_3055_2803# Vdd Vdd GND efet w=19 l=16
+ ad=0 pd=0 as=0 ps=0 
M2757 diff_3205_2761# Vdd Vdd GND efet w=19 l=17
+ ad=0 pd=0 as=0 ps=0 
M2758 diff_3544_3628# diff_3550_2758# diff_3544_3628# GND efet w=77 l=116
+ ad=0 pd=0 as=0 ps=0 
M2759 diff_3397_2791# diff_3397_2791# diff_3397_2791# GND efet w=4 l=7
+ ad=1111 pd=160 as=0 ps=0 
M2760 diff_3397_2791# diff_3397_2791# diff_3397_2791# GND efet w=3 l=7
+ ad=0 pd=0 as=0 ps=0 
M2761 diff_3400_2897# diff_3397_2791# Vdd GND efet w=19 l=91
+ ad=0 pd=0 as=0 ps=0 
M2762 diff_3544_3628# diff_3550_2758# Vdd GND efet w=19 l=91
+ ad=0 pd=0 as=0 ps=0 
M2763 GND diff_4243_2545# diff_4732_2900# GND efet w=46 l=16
+ ad=0 pd=0 as=0 ps=0 
M2764 GND diff_4243_2545# diff_4915_3191# GND efet w=46 l=17
+ ad=0 pd=0 as=0 ps=0 
M2765 GND diff_4243_2545# diff_5029_3068# GND efet w=52 l=16
+ ad=0 pd=0 as=0 ps=0 
M2766 GND diff_4243_2545# diff_5134_2953# GND efet w=46 l=16
+ ad=0 pd=0 as=0 ps=0 
M2767 diff_3745_2897# diff_3742_2791# diff_3745_2897# GND efet w=77 l=115
+ ad=0 pd=0 as=0 ps=0 
M2768 diff_3889_3628# diff_3892_2761# diff_3889_3628# GND efet w=120 l=68
+ ad=0 pd=0 as=0 ps=0 
M2769 diff_3550_2758# diff_3550_2758# diff_3550_2758# GND efet w=5 l=5
+ ad=1120 pd=160 as=0 ps=0 
M2770 diff_3397_2791# Vdd Vdd GND efet w=17 l=20
+ ad=0 pd=0 as=0 ps=0 
M2771 Vdd Vdd diff_550_2479# GND efet w=23 l=47
+ ad=0 pd=0 as=0 ps=0 
M2772 diff_550_2479# diff_550_2356# GND GND efet w=127 l=16
+ ad=0 pd=0 as=0 ps=0 
M2773 diff_580_3394# diff_508_1279# Vdd GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M2774 Vdd Vdd diff_1291_3103# GND efet w=22 l=115
+ ad=0 pd=0 as=5959 ps=640 
M2775 diff_2056_3184# diff_2101_2551# GND GND efet w=64 l=19
+ ad=0 pd=0 as=0 ps=0 
M2776 diff_2062_3349# diff_2818_2438# GND GND efet w=94 l=19
+ ad=9068 pd=1008 as=0 ps=0 
M2777 Vdd Vdd diff_2062_3349# GND efet w=19 l=73
+ ad=0 pd=0 as=0 ps=0 
M2778 diff_3254_2623# Vdd Vdd GND efet w=19 l=76
+ ad=8423 pd=1074 as=0 ps=0 
M2779 diff_3550_2758# diff_3550_2758# diff_3550_2758# GND efet w=3 l=7
+ ad=0 pd=0 as=0 ps=0 
M2780 diff_3550_2758# Vdd Vdd GND efet w=19 l=19
+ ad=0 pd=0 as=0 ps=0 
M2781 diff_3742_2791# diff_3742_2791# diff_3742_2791# GND efet w=5 l=5
+ ad=1246 pd=174 as=0 ps=0 
M2782 diff_3742_2791# diff_3742_2791# diff_3742_2791# GND efet w=4 l=8
+ ad=0 pd=0 as=0 ps=0 
M2783 diff_3745_2897# diff_3742_2791# Vdd GND efet w=19 l=91
+ ad=0 pd=0 as=0 ps=0 
M2784 diff_3889_3628# diff_3892_2761# Vdd GND efet w=19 l=91
+ ad=0 pd=0 as=0 ps=0 
M2785 diff_3892_2761# diff_3892_2761# diff_3892_2761# GND efet w=2 l=8
+ ad=1237 pd=174 as=0 ps=0 
M2786 diff_3742_2791# Vdd Vdd GND efet w=22 l=17
+ ad=0 pd=0 as=0 ps=0 
M2787 diff_3892_2761# diff_3892_2761# diff_3892_2761# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M2788 diff_3892_2761# Vdd Vdd GND efet w=22 l=16
+ ad=0 pd=0 as=0 ps=0 
M2789 diff_3254_2623# diff_2062_3349# GND GND efet w=61 l=16
+ ad=0 pd=0 as=0 ps=0 
M2790 diff_2743_3241# diff_3505_2438# GND GND efet w=94 l=19
+ ad=9125 pd=1062 as=0 ps=0 
M2791 Vdd Vdd diff_2743_3241# GND efet w=19 l=76
+ ad=0 pd=0 as=0 ps=0 
M2792 diff_2056_3301# Vdd Vdd GND efet w=17 l=74
+ ad=7841 pd=1002 as=0 ps=0 
M2793 diff_4087_2900# diff_4084_2797# diff_4087_2900# GND efet w=74 l=118
+ ad=0 pd=0 as=0 ps=0 
M2794 diff_4231_3628# diff_4237_2758# diff_4231_3628# GND efet w=118 l=60
+ ad=0 pd=0 as=0 ps=0 
M2795 diff_4084_2797# diff_4084_2797# diff_4084_2797# GND efet w=4 l=7
+ ad=1129 pd=160 as=0 ps=0 
M2796 diff_4084_2797# diff_4084_2797# diff_4084_2797# GND efet w=3 l=7
+ ad=0 pd=0 as=0 ps=0 
M2797 diff_4087_2900# diff_4084_2797# Vdd GND efet w=19 l=91
+ ad=0 pd=0 as=0 ps=0 
M2798 diff_4231_3628# diff_4237_2758# Vdd GND efet w=19 l=91
+ ad=0 pd=0 as=0 ps=0 
M2799 diff_4237_2758# diff_4237_2758# diff_4237_2758# GND efet w=4 l=5
+ ad=1204 pd=174 as=0 ps=0 
M2800 diff_4084_2797# Vdd Vdd GND efet w=19 l=17
+ ad=0 pd=0 as=0 ps=0 
M2801 diff_4237_2758# diff_4237_2758# diff_4237_2758# GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M2802 diff_4399_2803# diff_4417_2732# diff_4399_2803# GND efet w=117 l=59
+ ad=0 pd=0 as=0 ps=0 
M2803 diff_4552_2860# diff_4549_2758# diff_4552_2860# GND efet w=118 l=60
+ ad=0 pd=0 as=0 ps=0 
M2804 diff_4417_2732# diff_4417_2732# diff_4417_2732# GND efet w=4 l=7
+ ad=1324 pd=178 as=0 ps=0 
M2805 diff_4417_2732# diff_4417_2732# diff_4417_2732# GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M2806 diff_4399_2803# diff_4417_2732# Vdd GND efet w=19 l=91
+ ad=0 pd=0 as=0 ps=0 
M2807 diff_4552_2860# diff_4549_2758# Vdd GND efet w=19 l=91
+ ad=0 pd=0 as=0 ps=0 
M2808 diff_4549_2758# diff_4549_2758# diff_4549_2758# GND efet w=4 l=5
+ ad=1213 pd=174 as=0 ps=0 
M2809 diff_4237_2758# Vdd Vdd GND efet w=20 l=17
+ ad=0 pd=0 as=0 ps=0 
M2810 Vdd Vdd Vdd GND efet w=7 l=22
+ ad=0 pd=0 as=0 ps=0 
M2811 Vdd Vdd Vdd GND efet w=7 l=22
+ ad=0 pd=0 as=0 ps=0 
M2812 Vdd Vdd Vdd GND efet w=13 l=9
+ ad=0 pd=0 as=0 ps=0 
M2813 Vdd Vdd Vdd GND efet w=7 l=19
+ ad=0 pd=0 as=0 ps=0 
M2814 Vdd Vdd diff_2056_3070# GND efet w=22 l=76
+ ad=0 pd=0 as=3201 ps=364 
M2815 diff_2056_3301# diff_2743_3241# GND GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M2816 diff_4417_2732# Vdd Vdd GND efet w=19 l=19
+ ad=0 pd=0 as=0 ps=0 
M2817 diff_4549_2758# diff_4549_2758# diff_4549_2758# GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M2818 diff_4549_2758# Vdd Vdd GND efet w=20 l=16
+ ad=0 pd=0 as=0 ps=0 
M2819 Vdd Vdd Vdd GND efet w=3 l=13
+ ad=0 pd=0 as=0 ps=0 
M2820 Vdd Vdd Vdd GND efet w=5 l=20
+ ad=0 pd=0 as=0 ps=0 
M2821 Vdd Vdd Vdd GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M2822 Vdd Vdd Vdd GND efet w=13 l=9
+ ad=0 pd=0 as=0 ps=0 
M2823 diff_2056_3070# diff_2056_3070# diff_2056_3070# GND efet w=4 l=5
+ ad=0 pd=0 as=0 ps=0 
M2824 diff_2056_3070# diff_2056_3070# diff_2056_3070# GND efet w=5 l=8
+ ad=0 pd=0 as=0 ps=0 
M2825 Vdd Vdd diff_2209_3019# GND efet w=19 l=73
+ ad=0 pd=0 as=2988 ps=350 
M2826 diff_4732_2900# diff_4726_2803# diff_4732_2900# GND efet w=76 l=121
+ ad=0 pd=0 as=0 ps=0 
M2827 diff_4726_2803# diff_4726_2803# diff_4726_2803# GND efet w=5 l=5
+ ad=1186 pd=174 as=0 ps=0 
M2828 diff_4726_2803# diff_4726_2803# diff_4726_2803# GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M2829 diff_4732_2900# diff_4726_2803# Vdd GND efet w=19 l=91
+ ad=0 pd=0 as=0 ps=0 
M2830 diff_4726_2803# Vdd Vdd GND efet w=19 l=19
+ ad=0 pd=0 as=0 ps=0 
M2831 diff_5771_2965# Vdd Vdd GND efet w=25 l=67
+ ad=3176 pd=282 as=0 ps=0 
M2832 GND diff_5821_2920# diff_5771_2965# GND efet w=95 l=14
+ ad=0 pd=0 as=0 ps=0 
M2833 diff_4915_3191# diff_4927_2758# diff_4915_3191# GND efet w=130 l=63
+ ad=0 pd=0 as=0 ps=0 
M2834 diff_4915_3191# diff_4927_2758# Vdd GND efet w=19 l=94
+ ad=0 pd=0 as=0 ps=0 
M2835 diff_5029_3068# diff_5053_2732# diff_5029_3068# GND efet w=123 l=69
+ ad=0 pd=0 as=0 ps=0 
M2836 diff_5821_2920# diff_5821_2920# diff_5821_2920# GND efet w=2 l=9
+ ad=3540 pd=272 as=0 ps=0 
M2837 diff_4927_2758# diff_4927_2758# diff_4927_2758# GND efet w=4 l=7
+ ad=1087 pd=166 as=0 ps=0 
M2838 diff_4927_2758# diff_4927_2758# diff_4927_2758# GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M2839 diff_4243_2545# Vdd Vdd GND efet w=20 l=77
+ ad=5235 pd=518 as=0 ps=0 
M2840 diff_2209_3019# diff_2209_3019# diff_2209_3019# GND efet w=2 l=7
+ ad=0 pd=0 as=0 ps=0 
M2841 diff_2209_3019# diff_2209_3019# diff_2209_3019# GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M2842 diff_5053_2732# diff_5053_2732# diff_5053_2732# GND efet w=4 l=7
+ ad=1114 pd=160 as=0 ps=0 
M2843 diff_5053_2732# diff_5053_2732# diff_5053_2732# GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M2844 diff_5029_3068# diff_5053_2732# Vdd GND efet w=19 l=91
+ ad=0 pd=0 as=0 ps=0 
M2845 diff_4927_2758# Vdd Vdd GND efet w=16 l=17
+ ad=0 pd=0 as=0 ps=0 
M2846 diff_5053_2732# Vdd Vdd GND efet w=16 l=16
+ ad=0 pd=0 as=0 ps=0 
M2847 Vdd Vdd Vdd GND efet w=13 l=9
+ ad=0 pd=0 as=0 ps=0 
M2848 Vdd Vdd Vdd GND efet w=5 l=19
+ ad=0 pd=0 as=0 ps=0 
M2849 Vdd Vdd Vdd GND efet w=13 l=9
+ ad=0 pd=0 as=0 ps=0 
M2850 diff_4936_3115# diff_4936_3115# diff_4936_3115# GND efet w=8 l=12
+ ad=6141 pd=484 as=0 ps=0 
M2851 Vdd Vdd Vdd GND efet w=7 l=19
+ ad=0 pd=0 as=0 ps=0 
M2852 Vdd Vdd diff_4936_3115# GND efet w=19 l=88
+ ad=0 pd=0 as=0 ps=0 
M2853 diff_4936_3115# diff_4723_3052# GND GND efet w=103 l=16
+ ad=0 pd=0 as=0 ps=0 
M2854 diff_4936_3115# diff_4936_3115# diff_4936_3115# GND efet w=4 l=4
+ ad=0 pd=0 as=0 ps=0 
M2855 diff_4243_2545# diff_4243_2545# diff_4243_2545# GND efet w=3 l=15
+ ad=0 pd=0 as=0 ps=0 
M2856 diff_4243_2545# diff_4243_2545# diff_4243_2545# GND efet w=5 l=10
+ ad=0 pd=0 as=0 ps=0 
M2857 diff_4756_3238# Vdd Vdd GND efet w=20 l=89
+ ad=4023 pd=350 as=0 ps=0 
M2858 diff_4756_3238# diff_4756_3238# diff_4756_3238# GND efet w=8 l=18
+ ad=0 pd=0 as=0 ps=0 
M2859 diff_4756_3238# diff_4756_3238# diff_4756_3238# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M2860 diff_4243_2545# diff_4699_2554# GND GND efet w=115 l=17
+ ad=0 pd=0 as=0 ps=0 
M2861 diff_1436_2665# diff_1417_2311# diff_1291_3103# GND efet w=19 l=16
+ ad=0 pd=0 as=0 ps=0 
M2862 diff_1291_3103# diff_1291_3169# GND GND efet w=46 l=16
+ ad=0 pd=0 as=0 ps=0 
M2863 diff_2056_3070# diff_4243_2545# diff_4252_2516# GND efet w=121 l=16
+ ad=0 pd=0 as=3146 ps=294 
M2864 diff_2209_3019# diff_4243_2545# diff_4447_2516# GND efet w=121 l=16
+ ad=0 pd=0 as=4127 ps=402 
M2865 GND diff_4903_3178# diff_4756_3238# GND efet w=91 l=16
+ ad=0 pd=0 as=0 ps=0 
M2866 diff_5821_2920# diff_5821_2920# diff_5821_2920# GND efet w=7 l=7
+ ad=0 pd=0 as=0 ps=0 
M2867 diff_5821_2920# Vdd Vdd GND efet w=20 l=143
+ ad=0 pd=0 as=0 ps=0 
M2868 diff_5987_2827# diff_4481_442# diff_5821_2920# GND efet w=64 l=16
+ ad=5546 pd=458 as=0 ps=0 
M2869 diff_5987_2827# diff_2203_2482# GND GND efet w=67 l=16
+ ad=0 pd=0 as=0 ps=0 
M2870 GND diff_2122_2422# diff_5987_2827# GND efet w=73 l=14
+ ad=0 pd=0 as=0 ps=0 
M2871 diff_673_1115# clk1 diff_6091_2533# GND efet w=35 l=14
+ ad=6566 pd=590 as=1503 ps=158 
M2872 diff_4435_2500# diff_4435_2500# diff_4435_2500# GND efet w=3 l=7
+ ad=5079 pd=500 as=0 ps=0 
M2873 diff_4699_2554# diff_4699_2554# diff_4699_2554# GND efet w=3 l=7
+ ad=5280 pd=500 as=0 ps=0 
M2874 diff_4723_3052# diff_4723_3052# diff_4723_3052# GND efet w=3 l=7
+ ad=5004 pd=482 as=0 ps=0 
M2875 diff_4435_2500# diff_4435_2500# diff_4435_2500# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M2876 diff_4699_2554# diff_4699_2554# diff_4699_2554# GND efet w=4 l=4
+ ad=0 pd=0 as=0 ps=0 
M2877 diff_4723_3052# diff_4723_3052# diff_4723_3052# GND efet w=4 l=4
+ ad=0 pd=0 as=0 ps=0 
M2878 diff_2062_2569# diff_2203_2482# diff_2203_2368# GND efet w=31 l=16
+ ad=4865 pd=420 as=9395 ps=770 
M2879 diff_2818_2438# diff_2203_2482# diff_2890_2341# GND efet w=34 l=16
+ ad=6002 pd=522 as=8805 ps=772 
M2880 diff_4252_2516# diff_2209_3019# GND GND efet w=125 l=17
+ ad=0 pd=0 as=0 ps=0 
M2881 diff_3505_2438# diff_2203_2482# diff_3577_2338# GND efet w=31 l=16
+ ad=5678 pd=516 as=8688 ps=760 
M2882 diff_4447_2516# diff_4435_2500# GND GND efet w=187 l=16
+ ad=0 pd=0 as=0 ps=0 
M2883 diff_2062_2569# diff_2122_2422# diff_1921_2057# GND efet w=31 l=16
+ ad=0 pd=0 as=7827 ps=818 
M2884 diff_1405_2629# diff_1417_2311# GND GND efet w=34 l=16
+ ad=2540 pd=270 as=0 ps=0 
M2885 Vdd Vdd diff_1405_2629# GND efet w=19 l=145
+ ad=0 pd=0 as=0 ps=0 
M2886 diff_2818_2438# diff_2122_2422# diff_2608_2057# GND efet w=31 l=16
+ ad=0 pd=0 as=7942 ps=848 
M2887 diff_4435_2500# diff_2203_2482# diff_4462_2026# GND efet w=34 l=16
+ ad=0 pd=0 as=9372 ps=794 
M2888 GND diff_6091_2533# diff_2122_2422# GND efet w=130 l=13
+ ad=0 pd=0 as=10491 ps=898 
M2889 diff_4903_3178# diff_4903_3178# diff_4903_3178# GND efet w=7 l=19
+ ad=6273 pd=540 as=0 ps=0 
M2890 diff_4699_2554# diff_2203_2482# diff_4231_1556# GND efet w=31 l=16
+ ad=0 pd=0 as=7711 ps=720 
M2891 diff_3505_2438# diff_2122_2422# diff_3310_2065# GND efet w=32 l=16
+ ad=0 pd=0 as=5377 ps=622 
M2892 diff_2608_2057# diff_2608_2057# diff_2608_2057# GND efet w=5 l=8
+ ad=0 pd=0 as=0 ps=0 
M2893 diff_2608_2057# diff_2608_2057# diff_2608_2057# GND efet w=2 l=9
+ ad=0 pd=0 as=0 ps=0 
M2894 Vdd Vdd diff_595_2158# GND efet w=19 l=22
+ ad=0 pd=0 as=1054 ps=154 
M2895 diff_595_2158# diff_595_2158# diff_595_2158# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M2896 diff_595_2158# diff_595_2158# diff_595_2158# GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M2897 Vdd diff_595_2158# diff_556_2707# GND efet w=22 l=22
+ ad=0 pd=0 as=9055 ps=630 
M2898 diff_556_2707# diff_595_2158# diff_556_2707# GND efet w=89 l=66
+ ad=0 pd=0 as=0 ps=0 
M2899 diff_2890_2341# diff_2890_2341# diff_2890_2341# GND efet w=4 l=10
+ ad=0 pd=0 as=0 ps=0 
M2900 diff_2890_2341# diff_2890_2341# diff_2890_2341# GND efet w=2 l=9
+ ad=0 pd=0 as=0 ps=0 
M2901 diff_4435_2500# diff_2122_2422# diff_3997_2065# GND efet w=31 l=16
+ ad=0 pd=0 as=5563 ps=638 
M2902 diff_4723_3052# diff_2203_2482# diff_3722_1087# GND efet w=34 l=16
+ ad=0 pd=0 as=7243 ps=696 
M2903 Vdd Vdd Vdd GND efet w=3 l=7
+ ad=0 pd=0 as=0 ps=0 
M2904 diff_4903_3178# diff_4903_3178# diff_4903_3178# GND efet w=10 l=9
+ ad=0 pd=0 as=0 ps=0 
M2905 diff_4699_2554# diff_2122_2422# diff_4684_2065# GND efet w=34 l=16
+ ad=0 pd=0 as=5995 ps=668 
M2906 diff_4723_3052# diff_2122_2422# diff_2608_2057# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M2907 diff_3310_2065# diff_3310_2065# diff_3310_2065# GND efet w=5 l=14
+ ad=0 pd=0 as=0 ps=0 
M2908 diff_3310_2065# diff_3310_2065# diff_3310_2065# GND efet w=2 l=6
+ ad=0 pd=0 as=0 ps=0 
M2909 diff_556_2707# clk2 GND GND efet w=125 l=14
+ ad=0 pd=0 as=0 ps=0 
M2910 Vdd Vdd diff_1921_2057# GND efet w=25 l=58
+ ad=0 pd=0 as=0 ps=0 
M2911 diff_1912_2041# Vdd Vdd GND efet w=16 l=112
+ ad=4410 pd=470 as=0 ps=0 
M2912 diff_1921_2057# diff_1912_2041# GND GND efet w=82 l=19
+ ad=0 pd=0 as=0 ps=0 
M2913 diff_1912_2041# diff_1912_2041# diff_1912_2041# GND efet w=5 l=15
+ ad=0 pd=0 as=0 ps=0 
M2914 diff_1912_2041# diff_1912_2041# diff_1912_2041# GND efet w=3 l=8
+ ad=0 pd=0 as=0 ps=0 
M2915 Vdd Vdd diff_2098_1949# GND efet w=19 l=142
+ ad=0 pd=0 as=3737 ps=374 
M2916 diff_1939_1963# Vdd Vdd GND efet w=16 l=112
+ ad=4617 pd=446 as=0 ps=0 
M2917 diff_1939_1963# diff_1939_1963# diff_1939_1963# GND efet w=5 l=15
+ ad=0 pd=0 as=0 ps=0 
M2918 diff_1939_1963# diff_1939_1963# diff_1939_1963# GND efet w=5 l=10
+ ad=0 pd=0 as=0 ps=0 
M2919 GND diff_1939_1963# diff_2098_1949# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M2920 GND diff_965_1612# diff_1358_1843# GND efet w=34 l=16
+ ad=0 pd=0 as=4913 ps=520 
M2921 GND diff_1939_1963# diff_1912_2041# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M2922 diff_1358_1843# diff_1358_1843# diff_1358_1843# GND efet w=13 l=9
+ ad=0 pd=0 as=0 ps=0 
M2923 diff_1358_1843# diff_1358_1843# diff_1358_1843# GND efet w=7 l=19
+ ad=0 pd=0 as=0 ps=0 
M2924 diff_1921_2057# diff_1921_2057# diff_1921_2057# GND efet w=5 l=8
+ ad=0 pd=0 as=0 ps=0 
M2925 diff_1921_2057# diff_1921_2057# diff_1921_2057# GND efet w=5 l=14
+ ad=0 pd=0 as=0 ps=0 
M2926 diff_2098_1949# diff_965_1612# diff_1912_1771# GND efet w=35 l=17
+ ad=0 pd=0 as=2634 ps=224 
M2927 Vdd Vdd diff_2203_2368# GND efet w=25 l=91
+ ad=0 pd=0 as=0 ps=0 
M2928 Vdd Vdd diff_2479_1856# GND efet w=19 l=142
+ ad=0 pd=0 as=2956 ps=358 
M2929 Vdd Vdd diff_2608_2057# GND efet w=26 l=59
+ ad=0 pd=0 as=0 ps=0 
M2930 diff_2203_2368# diff_2203_2368# diff_2203_2368# GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M2931 GND diff_1912_2041# diff_1939_1963# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M2932 diff_2203_2368# diff_2203_2368# diff_2203_2368# GND efet w=7 l=7
+ ad=0 pd=0 as=0 ps=0 
M2933 diff_2479_1856# diff_2479_1856# diff_2479_1856# GND efet w=3 l=13
+ ad=0 pd=0 as=0 ps=0 
M2934 diff_2479_1856# diff_2479_1856# diff_2479_1856# GND efet w=6 l=10
+ ad=0 pd=0 as=0 ps=0 
M2935 diff_1921_2057# diff_965_1612# diff_2158_1852# GND efet w=34 l=16
+ ad=0 pd=0 as=2643 ps=224 
M2936 diff_1912_2041# diff_1358_1843# diff_1888_1780# GND efet w=74 l=17
+ ad=0 pd=0 as=4346 ps=416 
M2937 diff_944_1837# clk2 sync GND efet w=19 l=16
+ ad=1666 pd=190 as=25237 ps=2506 
M2938 diff_944_1837# diff_944_1837# diff_944_1837# GND efet w=4 l=4
+ ad=0 pd=0 as=0 ps=0 
M2939 diff_944_1837# diff_944_1837# diff_944_1837# GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M2940 diff_989_1735# diff_944_1837# GND GND efet w=76 l=16
+ ad=3814 pd=334 as=0 ps=0 
M2941 Vdd Vdd diff_989_1735# GND efet w=19 l=142
+ ad=0 pd=0 as=0 ps=0 
M2942 diff_1358_1843# Vdd Vdd GND efet w=22 l=145
+ ad=0 pd=0 as=0 ps=0 
M2943 GND diff_1361_1756# diff_1358_1843# GND efet w=32 l=17
+ ad=0 pd=0 as=0 ps=0 
M2944 GND diff_1912_1771# diff_1888_1780# GND efet w=125 l=17
+ ad=0 pd=0 as=0 ps=0 
M2945 diff_1361_1756# diff_1361_1756# diff_1361_1756# GND efet w=5 l=5
+ ad=2919 pd=316 as=0 ps=0 
M2946 diff_1361_1756# diff_1361_1756# diff_1361_1756# GND efet w=5 l=13
+ ad=0 pd=0 as=0 ps=0 
M2947 diff_949_1603# clk1 diff_989_1735# GND efet w=20 l=17
+ ad=1992 pd=224 as=0 ps=0 
M2948 diff_1361_1756# Vdd Vdd GND efet w=14 l=134
+ ad=0 pd=0 as=0 ps=0 
M2949 diff_965_1612# diff_949_1603# GND GND efet w=49 l=16
+ ad=2632 pd=274 as=0 ps=0 
M2950 diff_1361_1756# diff_989_1735# GND GND efet w=28 l=19
+ ad=0 pd=0 as=0 ps=0 
M2951 Vdd Vdd diff_965_1612# GND efet w=19 l=101
+ ad=0 pd=0 as=0 ps=0 
M2952 diff_965_1612# clk2 diff_886_1528# GND efet w=20 l=14
+ ad=0 pd=0 as=1323 ps=164 
M2953 GND diff_886_1528# diff_892_1507# GND efet w=35 l=14
+ ad=0 pd=0 as=3655 ps=382 
M2954 diff_2203_2368# diff_2377_1729# diff_2416_1697# GND efet w=31 l=19
+ ad=0 pd=0 as=6270 ps=610 
M2955 diff_1939_1963# diff_1358_1843# diff_2263_1867# GND efet w=67 l=16
+ ad=0 pd=0 as=4916 ps=446 
M2956 diff_2263_1867# diff_2158_1852# GND GND efet w=127 l=16
+ ad=0 pd=0 as=0 ps=0 
M2957 GND diff_2479_1856# diff_2203_2368# GND efet w=61 l=16
+ ad=0 pd=0 as=0 ps=0 
M2958 diff_2599_2041# Vdd Vdd GND efet w=16 l=112
+ ad=4578 pd=482 as=0 ps=0 
M2959 diff_2608_2057# diff_2599_2041# GND GND efet w=82 l=19
+ ad=0 pd=0 as=0 ps=0 
M2960 diff_2599_2041# diff_2599_2041# diff_2599_2041# GND efet w=5 l=15
+ ad=0 pd=0 as=0 ps=0 
M2961 diff_2599_2041# diff_2599_2041# diff_2599_2041# GND efet w=5 l=8
+ ad=0 pd=0 as=0 ps=0 
M2962 Vdd Vdd diff_2785_1949# GND efet w=19 l=142
+ ad=0 pd=0 as=3584 ps=374 
M2963 diff_2626_1963# Vdd Vdd GND efet w=17 l=110
+ ad=4509 pd=440 as=0 ps=0 
M2964 diff_2626_1963# diff_2626_1963# diff_2626_1963# GND efet w=3 l=13
+ ad=0 pd=0 as=0 ps=0 
M2965 diff_2626_1963# diff_2626_1963# diff_2626_1963# GND efet w=5 l=10
+ ad=0 pd=0 as=0 ps=0 
M2966 GND diff_2626_1963# diff_2785_1949# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M2967 GND diff_2626_1963# diff_2599_2041# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M2968 diff_2608_2057# diff_2608_2057# diff_2608_2057# GND efet w=5 l=8
+ ad=0 pd=0 as=0 ps=0 
M2969 diff_2608_2057# diff_2608_2057# diff_2608_2057# GND efet w=5 l=11
+ ad=0 pd=0 as=0 ps=0 
M2970 diff_2785_1949# diff_1912_2041# diff_2599_1771# GND efet w=35 l=20
+ ad=0 pd=0 as=2598 ps=224 
M2971 diff_3577_2338# diff_3577_2338# diff_3577_2338# GND efet w=4 l=7
+ ad=0 pd=0 as=0 ps=0 
M2972 diff_3997_2065# diff_3997_2065# diff_3997_2065# GND efet w=8 l=8
+ ad=0 pd=0 as=0 ps=0 
M2973 diff_4462_2026# diff_4462_2026# diff_4462_2026# GND efet w=5 l=10
+ ad=0 pd=0 as=0 ps=0 
M2974 diff_3577_2338# diff_3577_2338# diff_3577_2338# GND efet w=2 l=9
+ ad=0 pd=0 as=0 ps=0 
M2975 diff_3997_2065# diff_3997_2065# diff_3997_2065# GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M2976 diff_4462_2026# diff_4462_2026# diff_4462_2026# GND efet w=2 l=9
+ ad=0 pd=0 as=0 ps=0 
M2977 diff_4684_2065# diff_4684_2065# diff_4684_2065# GND efet w=8 l=8
+ ad=0 pd=0 as=0 ps=0 
M2978 diff_4231_1556# diff_4231_1556# diff_4231_1556# GND efet w=6 l=10
+ ad=0 pd=0 as=0 ps=0 
M2979 diff_4684_2065# diff_4684_2065# diff_4684_2065# GND efet w=2 l=9
+ ad=0 pd=0 as=0 ps=0 
M2980 diff_4231_1556# diff_4231_1556# diff_4231_1556# GND efet w=2 l=9
+ ad=0 pd=0 as=0 ps=0 
M2981 Vdd Vdd Vdd GND efet w=8 l=10
+ ad=0 pd=0 as=0 ps=0 
M2982 diff_2122_2422# Vdd Vdd GND efet w=25 l=46
+ ad=0 pd=0 as=0 ps=0 
M2983 diff_4903_3178# diff_2203_2482# diff_3962_1084# GND efet w=31 l=16
+ ad=0 pd=0 as=7303 ps=718 
M2984 diff_3722_1087# diff_3722_1087# diff_3722_1087# GND efet w=4 l=8
+ ad=0 pd=0 as=0 ps=0 
M2985 diff_4903_3178# diff_2122_2422# diff_1921_2057# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M2986 diff_2890_2341# Vdd Vdd GND efet w=23 l=92
+ ad=0 pd=0 as=0 ps=0 
M2987 Vdd Vdd diff_3166_1856# GND efet w=19 l=142
+ ad=0 pd=0 as=2956 ps=354 
M2988 Vdd Vdd diff_3310_2065# GND efet w=25 l=91
+ ad=0 pd=0 as=0 ps=0 
M2989 diff_3289_1904# Vdd Vdd GND efet w=16 l=124
+ ad=4488 pd=494 as=0 ps=0 
M2990 diff_2890_2341# diff_2890_2341# diff_2890_2341# GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M2991 GND diff_2599_2041# diff_2626_1963# GND efet w=35 l=17
+ ad=0 pd=0 as=0 ps=0 
M2992 diff_2890_2341# diff_2890_2341# diff_2890_2341# GND efet w=7 l=7
+ ad=0 pd=0 as=0 ps=0 
M2993 diff_3166_1856# diff_3166_1856# diff_3166_1856# GND efet w=3 l=13
+ ad=0 pd=0 as=0 ps=0 
M2994 diff_3166_1856# diff_3166_1856# diff_3166_1856# GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M2995 diff_2608_2057# diff_1912_2041# diff_2845_1858# GND efet w=37 l=16
+ ad=0 pd=0 as=2625 ps=224 
M2996 diff_2599_2041# diff_1939_1963# diff_2569_1822# GND efet w=71 l=16
+ ad=0 pd=0 as=5078 ps=458 
M2997 diff_2416_1697# diff_2416_1697# diff_2416_1697# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M2998 diff_2416_1697# diff_2416_1697# diff_2416_1697# GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M2999 diff_2479_1856# diff_2416_1697# GND GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M3000 GND diff_2599_1771# diff_2569_1822# GND efet w=143 l=17
+ ad=0 pd=0 as=0 ps=0 
M3001 diff_2890_2341# diff_2377_1729# diff_3103_1685# GND efet w=31 l=17
+ ad=0 pd=0 as=6489 ps=634 
M3002 diff_2626_1963# diff_1939_1963# diff_2950_1870# GND efet w=67 l=16
+ ad=0 pd=0 as=4934 ps=440 
M3003 GND diff_2845_1858# diff_2950_1870# GND efet w=125 l=17
+ ad=0 pd=0 as=0 ps=0 
M3004 GND diff_3166_1856# diff_2890_2341# GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M3005 diff_3310_2065# diff_3289_1904# GND GND efet w=61 l=17
+ ad=0 pd=0 as=0 ps=0 
M3006 diff_3289_1904# diff_3289_1904# diff_3289_1904# GND efet w=2 l=12
+ ad=0 pd=0 as=0 ps=0 
M3007 diff_3289_1904# diff_3289_1904# diff_3289_1904# GND efet w=6 l=10
+ ad=0 pd=0 as=0 ps=0 
M3008 Vdd Vdd diff_3475_1949# GND efet w=19 l=142
+ ad=0 pd=0 as=3299 ps=350 
M3009 diff_3313_1963# Vdd Vdd GND efet w=16 l=112
+ ad=4488 pd=446 as=0 ps=0 
M3010 diff_3313_1963# diff_3313_1963# diff_3313_1963# GND efet w=2 l=12
+ ad=0 pd=0 as=0 ps=0 
M3011 diff_3313_1963# diff_3313_1963# diff_3313_1963# GND efet w=5 l=10
+ ad=0 pd=0 as=0 ps=0 
M3012 GND diff_3313_1963# diff_3475_1949# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M3013 GND diff_3313_1963# diff_3289_1904# GND efet w=34 l=19
+ ad=0 pd=0 as=0 ps=0 
M3014 diff_3310_2065# diff_3310_2065# diff_3310_2065# GND efet w=4 l=8
+ ad=0 pd=0 as=0 ps=0 
M3015 diff_3310_2065# diff_3310_2065# diff_3310_2065# GND efet w=4 l=5
+ ad=0 pd=0 as=0 ps=0 
M3016 diff_3722_1087# diff_3722_1087# diff_3722_1087# GND efet w=2 l=12
+ ad=0 pd=0 as=0 ps=0 
M3017 diff_2122_2422# diff_2122_2422# diff_2122_2422# GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M3018 diff_2122_2422# diff_2122_2422# diff_2122_2422# GND efet w=7 l=7
+ ad=0 pd=0 as=0 ps=0 
M3019 diff_3962_1084# diff_3962_1084# diff_3962_1084# GND efet w=5 l=10
+ ad=0 pd=0 as=0 ps=0 
M3020 diff_2122_2422# clk2 diff_6091_2320# GND efet w=34 l=16
+ ad=0 pd=0 as=1512 ps=158 
M3021 diff_3962_1084# diff_3962_1084# diff_3962_1084# GND efet w=2 l=9
+ ad=0 pd=0 as=0 ps=0 
M3022 Vdd Vdd diff_3577_2338# GND efet w=22 l=91
+ ad=0 pd=0 as=0 ps=0 
M3023 Vdd Vdd diff_3853_1856# GND efet w=19 l=142
+ ad=0 pd=0 as=3556 ps=366 
M3024 Vdd Vdd diff_3997_2065# GND efet w=22 l=91
+ ad=0 pd=0 as=0 ps=0 
M3025 diff_3577_2338# diff_3577_2338# diff_3577_2338# GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M3026 GND diff_3289_1904# diff_3313_1963# GND efet w=35 l=16
+ ad=0 pd=0 as=0 ps=0 
M3027 diff_3577_2338# diff_3577_2338# diff_3577_2338# GND efet w=7 l=7
+ ad=0 pd=0 as=0 ps=0 
M3028 diff_3853_1856# diff_3853_1856# diff_3853_1856# GND efet w=3 l=13
+ ad=0 pd=0 as=0 ps=0 
M3029 diff_3853_1856# diff_3853_1856# diff_3853_1856# GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M3030 diff_3475_1949# diff_2599_2041# diff_3286_1771# GND efet w=31 l=19
+ ad=0 pd=0 as=2517 ps=236 
M3031 diff_3310_2065# diff_2599_2041# diff_3532_1855# GND efet w=34 l=19
+ ad=0 pd=0 as=2634 ps=224 
M3032 diff_3103_1685# diff_3103_1685# diff_3103_1685# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M3033 diff_3289_1904# diff_2626_1963# diff_3259_1780# GND efet w=77 l=17
+ ad=0 pd=0 as=4961 ps=458 
M3034 diff_3103_1685# diff_3103_1685# diff_3103_1685# GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M3035 diff_3166_1856# diff_3103_1685# GND GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M3036 GND diff_3286_1771# diff_3259_1780# GND efet w=145 l=16
+ ad=0 pd=0 as=0 ps=0 
M3037 diff_3577_2338# diff_2377_1729# diff_3781_1697# GND efet w=31 l=17
+ ad=0 pd=0 as=6144 ps=610 
M3038 diff_3637_1879# diff_2626_1963# diff_3313_1963# GND efet w=67 l=19
+ ad=4769 pd=446 as=0 ps=0 
M3039 diff_3637_1879# diff_3532_1855# GND GND efet w=124 l=16
+ ad=0 pd=0 as=0 ps=0 
M3040 GND diff_3853_1856# diff_3577_2338# GND efet w=58 l=16
+ ad=0 pd=0 as=0 ps=0 
M3041 diff_3976_1904# Vdd Vdd GND efet w=16 l=112
+ ad=4434 pd=488 as=0 ps=0 
M3042 diff_3997_2065# diff_3976_1904# GND GND efet w=58 l=17
+ ad=0 pd=0 as=0 ps=0 
M3043 diff_3976_1904# diff_3976_1904# diff_3976_1904# GND efet w=2 l=12
+ ad=0 pd=0 as=0 ps=0 
M3044 diff_3976_1904# diff_3976_1904# diff_3976_1904# GND efet w=5 l=8
+ ad=0 pd=0 as=0 ps=0 
M3045 Vdd Vdd diff_4162_1949# GND efet w=19 l=142
+ ad=0 pd=0 as=3371 ps=356 
M3046 diff_4000_1963# Vdd Vdd GND efet w=16 l=112
+ ad=4386 pd=434 as=0 ps=0 
M3047 diff_4000_1963# diff_4000_1963# diff_4000_1963# GND efet w=3 l=13
+ ad=0 pd=0 as=0 ps=0 
M3048 diff_4000_1963# diff_4000_1963# diff_4000_1963# GND efet w=5 l=8
+ ad=0 pd=0 as=0 ps=0 
M3049 GND diff_4000_1963# diff_4162_1949# GND efet w=32 l=20
+ ad=0 pd=0 as=0 ps=0 
M3050 GND diff_4000_1963# diff_3976_1904# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M3051 diff_3997_2065# diff_3997_2065# diff_3997_2065# GND efet w=5 l=8
+ ad=0 pd=0 as=0 ps=0 
M3052 diff_3997_2065# diff_3997_2065# diff_3997_2065# GND efet w=5 l=11
+ ad=0 pd=0 as=0 ps=0 
M3053 diff_4162_1949# diff_3289_1904# diff_3973_1771# GND efet w=32 l=17
+ ad=0 pd=0 as=2418 ps=218 
M3054 Vdd Vdd diff_4462_2026# GND efet w=22 l=94
+ ad=0 pd=0 as=0 ps=0 
M3055 Vdd Vdd diff_4543_1856# GND efet w=19 l=142
+ ad=0 pd=0 as=3472 ps=352 
M3056 Vdd Vdd diff_4684_2065# GND efet w=25 l=91
+ ad=0 pd=0 as=0 ps=0 
M3057 diff_4666_1904# Vdd Vdd GND efet w=14 l=113
+ ad=4386 pd=496 as=0 ps=0 
M3058 diff_4462_2026# diff_4462_2026# diff_4462_2026# GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M3059 diff_4462_2026# diff_4462_2026# diff_4462_2026# GND efet w=6 l=7
+ ad=0 pd=0 as=0 ps=0 
M3060 GND diff_3976_1904# diff_4000_1963# GND efet w=32 l=16
+ ad=0 pd=0 as=0 ps=0 
M3061 diff_4543_1856# diff_4543_1856# diff_4543_1856# GND efet w=2 l=12
+ ad=0 pd=0 as=0 ps=0 
M3062 diff_4543_1856# diff_4543_1856# diff_4543_1856# GND efet w=5 l=10
+ ad=0 pd=0 as=0 ps=0 
M3063 GND diff_4543_1856# diff_4462_2026# GND efet w=68 l=17
+ ad=0 pd=0 as=0 ps=0 
M3064 diff_3997_2065# diff_3289_1904# diff_4222_1852# GND efet w=31 l=16
+ ad=0 pd=0 as=2418 ps=218 
M3065 diff_3976_1904# diff_3313_1963# diff_3946_1780# GND efet w=71 l=17
+ ad=0 pd=0 as=4937 ps=440 
M3066 diff_3781_1697# diff_3781_1697# diff_3781_1697# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M3067 diff_3781_1697# diff_3781_1697# diff_3781_1697# GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M3068 diff_2416_1697# diff_2407_1684# diff_872_2743# GND efet w=31 l=13
+ ad=0 pd=0 as=0 ps=0 
M3069 diff_3103_1685# diff_2407_1684# diff_629_6919# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M3070 Vdd Vdd diff_892_1507# GND efet w=19 l=145
+ ad=0 pd=0 as=0 ps=0 
M3071 GND GND diff_1387_1337# GND efet w=94 l=17
+ ad=0 pd=0 as=10638 ps=1002 
M3072 diff_892_1507# clk1 diff_886_1384# GND efet w=20 l=14
+ ad=0 pd=0 as=1471 ps=216 
M3073 GND diff_580_3394# diff_1387_1337# GND efet w=211 l=16
+ ad=0 pd=0 as=0 ps=0 
M3074 diff_886_1384# diff_886_1384# diff_886_1384# GND efet w=8 l=8
+ ad=0 pd=0 as=0 ps=0 
M3075 GND diff_886_1384# diff_892_1357# GND efet w=34 l=14
+ ad=0 pd=0 as=3919 ps=400 
M3076 diff_886_1384# diff_886_1384# diff_886_1384# GND efet w=5 l=10
+ ad=0 pd=0 as=0 ps=0 
M3077 diff_1387_1249# Vdd diff_1387_1337# GND efet w=101 l=17
+ ad=13750 pd=1250 as=0 ps=0 
M3078 Vdd Vdd diff_892_1357# GND efet w=19 l=142
+ ad=0 pd=0 as=0 ps=0 
M3079 GND diff_577_5317# diff_1582_1201# GND efet w=220 l=19
+ ad=0 pd=0 as=15343 ps=1238 
M3080 diff_1513_1009# diff_577_5317# GND GND efet w=115 l=19
+ ad=5508 pd=574 as=0 ps=0 
M3081 diff_1387_1337# diff_1378_1321# diff_1387_1249# GND efet w=133 l=16
+ ad=0 pd=0 as=0 ps=0 
M3082 clk1 GND GND GND efet w=262 l=13
+ ad=22314 pd=1600 as=0 ps=0 
M3083 GND diff_715_1141# diff_673_1115# GND efet w=124 l=16
+ ad=0 pd=0 as=0 ps=0 
M3084 diff_892_1357# clk2 diff_883_1234# GND efet w=19 l=13
+ ad=0 pd=0 as=1510 ps=216 
M3085 diff_883_1234# diff_883_1234# diff_883_1234# GND efet w=7 l=7
+ ad=0 pd=0 as=0 ps=0 
M3086 GND diff_883_1234# diff_892_1207# GND efet w=34 l=14
+ ad=0 pd=0 as=3583 ps=370 
M3087 GND diff_580_3394# diff_1378_1321# GND efet w=100 l=19
+ ad=0 pd=0 as=3059 ps=300 
M3088 diff_1417_2311# diff_1417_2311# diff_1417_2311# GND efet w=8 l=8
+ ad=16044 pd=2080 as=0 ps=0 
M3089 diff_1417_2311# diff_1417_2311# diff_1417_2311# GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M3090 diff_1859_1291# diff_1834_1103# GND GND efet w=34 l=16
+ ad=3602 pd=356 as=0 ps=0 
M3091 diff_883_1234# diff_883_1234# diff_883_1234# GND efet w=5 l=10
+ ad=0 pd=0 as=0 ps=0 
M3092 GND diff_769_1192# diff_778_1165# GND efet w=85 l=13
+ ad=0 pd=0 as=4690 ps=430 
M3093 Vdd Vdd diff_892_1207# GND efet w=19 l=142
+ ad=0 pd=0 as=0 ps=0 
M3094 diff_1378_1321# Vdd Vdd GND efet w=25 l=94
+ ad=0 pd=0 as=0 ps=0 
M3095 GND p0 diff_1582_1201# GND efet w=101 l=17
+ ad=0 pd=0 as=0 ps=0 
M3096 GND p0 diff_1642_1000# GND efet w=34 l=16
+ ad=0 pd=0 as=3255 ps=364 
M3097 diff_1859_1291# diff_1417_2311# diff_1825_1156# GND efet w=32 l=17
+ ad=0 pd=0 as=3339 ps=364 
M3098 GND diff_1417_2311# diff_1942_1112# GND efet w=31 l=20
+ ad=0 pd=0 as=3117 ps=318 
M3099 diff_892_1207# clk1 diff_769_1192# GND efet w=35 l=14
+ ad=0 pd=0 as=1323 ps=146 
M3100 diff_715_1141# diff_715_1141# diff_715_1141# GND efet w=5 l=15
+ ad=1492 pd=184 as=0 ps=0 
M3101 diff_673_1115# Vdd Vdd GND efet w=22 l=43
+ ad=0 pd=0 as=0 ps=0 
M3102 diff_715_1141# diff_715_1141# diff_715_1141# GND efet w=7 l=7
+ ad=0 pd=0 as=0 ps=0 
M3103 diff_778_1165# clk2 diff_715_1141# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M3104 diff_1582_1201# diff_1513_1009# diff_1387_1249# GND efet w=136 l=19
+ ad=0 pd=0 as=0 ps=0 
M3105 diff_778_1165# Vdd Vdd GND efet w=23 l=65
+ ad=0 pd=0 as=0 ps=0 
M3106 diff_1642_1000# diff_1642_1000# diff_1642_1000# GND efet w=7 l=10
+ ad=0 pd=0 as=0 ps=0 
M3107 GND diff_1825_1156# diff_1834_1103# GND efet w=59 l=17
+ ad=0 pd=0 as=2111 ps=210 
M3108 diff_1642_1000# diff_1642_1000# diff_1642_1000# GND efet w=5 l=13
+ ad=0 pd=0 as=0 ps=0 
M3109 diff_1942_1112# diff_1942_1112# diff_1942_1112# GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M3110 diff_2026_1181# diff_1942_1112# diff_1387_1249# GND efet w=31 l=19
+ ad=2619 pd=292 as=0 ps=0 
M3111 diff_1387_1249# diff_1642_1000# diff_1582_1201# GND efet w=133 l=19
+ ad=0 pd=0 as=0 ps=0 
M3112 Vdd Vdd diff_847_706# GND efet w=20 l=14
+ ad=0 pd=0 as=1516 ps=202 
M3113 diff_508_1279# diff_847_706# diff_508_1279# GND efet w=126 l=27
+ ad=9343 pd=914 as=0 ps=0 
M3114 diff_847_706# diff_847_706# diff_847_706# GND efet w=5 l=11
+ ad=0 pd=0 as=0 ps=0 
M3115 diff_847_706# diff_847_706# diff_847_706# GND efet w=2 l=9
+ ad=0 pd=0 as=0 ps=0 
M3116 diff_508_1279# diff_847_706# Vdd GND efet w=28 l=49
+ ad=0 pd=0 as=0 ps=0 
M3117 Vdd Vdd diff_916_577# GND efet w=19 l=142
+ ad=0 pd=0 as=2408 ps=234 
M3118 Vdd diff_1195_823# diff_331_7000# GND efet w=49 l=14
+ ad=0 pd=0 as=21139 ps=2348 
M3119 diff_331_7000# diff_1153_682# GND GND efet w=46 l=16
+ ad=0 pd=0 as=0 ps=0 
M3120 diff_916_577# clk1 diff_1036_647# GND efet w=67 l=19
+ ad=0 pd=0 as=2726 ps=240 
M3121 diff_508_1279# diff_916_577# GND GND efet w=109 l=14
+ ad=0 pd=0 as=0 ps=0 
M3122 diff_1036_647# diff_1027_631# GND GND efet w=64 l=16
+ ad=0 pd=0 as=0 ps=0 
M3123 Vdd Vdd diff_1153_682# GND efet w=19 l=142
+ ad=0 pd=0 as=2348 ps=228 
M3124 diff_1513_1009# Vdd Vdd GND efet w=22 l=76
+ ad=0 pd=0 as=0 ps=0 
M3125 Vdd Vdd diff_1387_1249# GND efet w=25 l=97
+ ad=0 pd=0 as=0 ps=0 
M3126 diff_1642_1000# Vdd Vdd GND efet w=19 l=143
+ ad=0 pd=0 as=0 ps=0 
M3127 diff_1942_1112# diff_1942_1112# diff_1942_1112# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M3128 diff_3853_1856# diff_3781_1697# GND GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M3129 GND diff_3973_1771# diff_3946_1780# GND efet w=140 l=17
+ ad=0 pd=0 as=0 ps=0 
M3130 diff_4462_2026# diff_2377_1729# diff_4477_1730# GND efet w=34 l=17
+ ad=0 pd=0 as=6126 ps=574 
M3131 diff_4000_1963# diff_3313_1963# diff_4327_1867# GND efet w=64 l=16
+ ad=0 pd=0 as=4487 ps=434 
M3132 diff_4327_1867# diff_4222_1852# GND GND efet w=124 l=16
+ ad=0 pd=0 as=0 ps=0 
M3133 diff_4684_2065# diff_4666_1904# GND GND efet w=61 l=16
+ ad=0 pd=0 as=0 ps=0 
M3134 diff_4666_1904# diff_4666_1904# diff_4666_1904# GND efet w=3 l=13
+ ad=0 pd=0 as=0 ps=0 
M3135 diff_4666_1904# diff_4666_1904# diff_4666_1904# GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M3136 Vdd Vdd diff_4852_1946# GND efet w=19 l=142
+ ad=0 pd=0 as=3290 ps=350 
M3137 diff_4687_1963# Vdd Vdd GND efet w=16 l=125
+ ad=4641 pd=466 as=0 ps=0 
M3138 diff_4687_1963# diff_4687_1963# diff_4687_1963# GND efet w=2 l=12
+ ad=0 pd=0 as=0 ps=0 
M3139 diff_4687_1963# diff_4687_1963# diff_4687_1963# GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M3140 GND diff_4687_1963# diff_4852_1946# GND efet w=31 l=19
+ ad=0 pd=0 as=0 ps=0 
M3141 GND diff_4687_1963# diff_4666_1904# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M3142 diff_4684_2065# diff_4684_2065# diff_4684_2065# GND efet w=3 l=5
+ ad=0 pd=0 as=0 ps=0 
M3143 diff_4684_2065# diff_4684_2065# diff_4684_2065# GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M3144 GND diff_4666_1904# diff_4687_1963# GND efet w=34 l=16
+ ad=0 pd=0 as=0 ps=0 
M3145 diff_4852_1946# diff_3976_1904# diff_4663_1771# GND efet w=32 l=17
+ ad=0 pd=0 as=2445 ps=224 
M3146 diff_4684_2065# diff_3976_1904# diff_4909_1861# GND efet w=34 l=16
+ ad=0 pd=0 as=2616 ps=224 
M3147 diff_4666_1904# diff_4000_1963# diff_4633_1837# GND efet w=64 l=16
+ ad=0 pd=0 as=5033 ps=446 
M3148 diff_4477_1730# diff_4477_1730# diff_4477_1730# GND efet w=7 l=7
+ ad=0 pd=0 as=0 ps=0 
M3149 diff_4477_1730# diff_4477_1730# diff_4477_1730# GND efet w=4 l=4
+ ad=0 pd=0 as=0 ps=0 
M3150 diff_4543_1856# diff_4477_1730# GND GND efet w=55 l=16
+ ad=0 pd=0 as=0 ps=0 
M3151 GND diff_4663_1771# diff_4633_1837# GND efet w=142 l=16
+ ad=0 pd=0 as=0 ps=0 
M3152 diff_4687_1963# diff_4000_1963# diff_5017_1867# GND efet w=64 l=16
+ ad=0 pd=0 as=4520 ps=446 
M3153 diff_5017_1867# diff_4909_1861# GND GND efet w=130 l=16
+ ad=0 pd=0 as=0 ps=0 
M3154 diff_4477_1730# diff_2407_1684# diff_580_3394# GND efet w=41 l=16
+ ad=0 pd=0 as=0 ps=0 
M3155 GND diff_4720_1750# diff_4732_1658# GND efet w=160 l=16
+ ad=0 pd=0 as=14528 ps=1440 
M3156 diff_3781_1697# diff_2407_1684# diff_577_5317# GND efet w=31 l=16
+ ad=0 pd=0 as=0 ps=0 
M3157 diff_4732_1658# diff_4720_1633# diff_4732_1658# GND efet w=105 l=53
+ ad=0 pd=0 as=0 ps=0 
M3158 GND diff_6091_2320# diff_5470_1585# GND efet w=62 l=16
+ ad=0 pd=0 as=16764 ps=2040 
M3159 diff_4102_1499# Vdd Vdd GND efet w=26 l=85
+ ad=4296 pd=368 as=0 ps=0 
M3160 diff_4732_1658# diff_4720_1633# Vdd GND efet w=23 l=26
+ ad=0 pd=0 as=0 ps=0 
M3161 GND diff_1834_1103# diff_2128_1144# GND efet w=85 l=16
+ ad=0 pd=0 as=5813 ps=518 
M3162 diff_2714_1150# diff_2026_1181# GND GND efet w=58 l=16
+ ad=5066 pd=532 as=0 ps=0 
M3163 GND diff_965_1612# diff_2026_1181# GND efet w=35 l=17
+ ad=0 pd=0 as=0 ps=0 
M3164 diff_2714_1150# diff_2714_1150# diff_2714_1150# GND efet w=13 l=9
+ ad=0 pd=0 as=0 ps=0 
M3165 diff_2714_1150# diff_2452_1015# GND GND efet w=34 l=19
+ ad=0 pd=0 as=0 ps=0 
M3166 GND clk2 diff_2929_1223# GND efet w=55 l=19
+ ad=0 pd=0 as=1973 ps=204 
M3167 Vdd Vdd diff_4231_1556# GND efet w=25 l=46
+ ad=0 pd=0 as=0 ps=0 
M3168 diff_4720_1633# diff_4720_1633# diff_4720_1633# GND efet w=2 l=9
+ ad=1309 pd=178 as=0 ps=0 
M3169 diff_4720_1633# diff_4720_1633# diff_4720_1633# GND efet w=5 l=8
+ ad=0 pd=0 as=0 ps=0 
M3170 diff_4345_1120# Vdd Vdd GND efet w=25 l=94
+ ad=6782 pd=724 as=0 ps=0 
M3171 Vdd Vdd diff_4477_1126# GND efet w=23 l=92
+ ad=0 pd=0 as=8986 ps=898 
M3172 diff_3971_1525# diff_2128_1144# diff_577_5317# GND efet w=31 l=16
+ ad=1212 pd=146 as=0 ps=0 
M3173 diff_4102_1499# diff_4102_1499# diff_4102_1499# GND efet w=3 l=5
+ ad=0 pd=0 as=0 ps=0 
M3174 diff_4231_1556# diff_4102_1499# GND GND efet w=143 l=17
+ ad=0 pd=0 as=0 ps=0 
M3175 diff_4231_1556# diff_4231_1556# diff_4231_1556# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M3176 diff_4102_1499# diff_4102_1499# diff_4102_1499# GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M3177 diff_629_6919# diff_2128_1144# diff_3562_1297# GND efet w=31 l=16
+ ad=0 pd=0 as=1488 ps=158 
M3178 diff_872_2743# diff_2128_1144# diff_3709_1297# GND efet w=31 l=16
+ ad=0 pd=0 as=1488 ps=158 
M3179 diff_2377_1729# diff_2377_1729# diff_2377_1729# GND efet w=3 l=10
+ ad=5499 pd=604 as=0 ps=0 
M3180 diff_2714_1150# diff_2714_1150# diff_2714_1150# GND efet w=8 l=20
+ ad=0 pd=0 as=0 ps=0 
M3181 GND diff_2714_1150# diff_2797_1142# GND efet w=32 l=17
+ ad=0 pd=0 as=1556 ps=174 
M3182 diff_2929_1223# diff_1654_625# diff_2929_1181# GND efet w=74 l=17
+ ad=0 pd=0 as=1688 ps=198 
M3183 diff_2929_1181# diff_2797_1142# diff_2929_1138# GND efet w=73 l=19
+ ad=0 pd=0 as=4262 ps=390 
M3184 diff_1834_1103# Vdd Vdd GND efet w=19 l=142
+ ad=0 pd=0 as=0 ps=0 
M3185 diff_1859_1291# Vdd Vdd GND efet w=19 l=140
+ ad=0 pd=0 as=0 ps=0 
M3186 diff_1942_1112# Vdd Vdd GND efet w=19 l=142
+ ad=0 pd=0 as=0 ps=0 
M3187 diff_1387_1249# diff_1942_1112# diff_1825_1156# GND efet w=34 l=19
+ ad=0 pd=0 as=0 ps=0 
M3188 GND diff_2185_1084# diff_2128_1144# GND efet w=82 l=16
+ ad=0 pd=0 as=0 ps=0 
M3189 diff_2378_1045# clk2 diff_1417_2311# GND efet w=76 l=19
+ ad=2717 pd=252 as=0 ps=0 
M3190 diff_2128_1144# Vdd Vdd GND efet w=22 l=70
+ ad=0 pd=0 as=0 ps=0 
M3191 diff_1417_2311# Vdd Vdd GND efet w=19 l=142
+ ad=0 pd=0 as=0 ps=0 
M3192 diff_1153_682# diff_1195_823# GND GND efet w=34 l=19
+ ad=0 pd=0 as=0 ps=0 
M3193 Vdd Vdd diff_1195_823# GND efet w=19 l=142
+ ad=0 pd=0 as=5758 ps=484 
M3194 diff_1375_760# Vdd Vdd GND efet w=16 l=136
+ ad=1733 pd=204 as=0 ps=0 
M3195 Vdd Vdd diff_1471_625# GND efet w=16 l=112
+ ad=0 pd=0 as=5517 ps=430 
M3196 diff_1568_757# diff_1027_631# Vdd GND efet w=32 l=17
+ ad=1655 pd=186 as=0 ps=0 
M3197 diff_1568_757# clk1 diff_1531_577# GND efet w=19 l=16
+ ad=0 pd=0 as=3810 ps=352 
M3198 GND diff_1744_715# diff_1375_760# GND efet w=29 l=20
+ ad=0 pd=0 as=0 ps=0 
M3199 diff_1531_577# diff_1531_577# diff_1531_577# GND efet w=8 l=8
+ ad=0 pd=0 as=0 ps=0 
M3200 diff_1531_577# diff_1531_577# diff_1531_577# GND efet w=4 l=12
+ ad=0 pd=0 as=0 ps=0 
M3201 diff_1471_625# diff_1471_625# diff_1471_625# GND efet w=8 l=8
+ ad=0 pd=0 as=0 ps=0 
M3202 GND diff_1531_577# diff_1471_625# GND efet w=104 l=17
+ ad=0 pd=0 as=0 ps=0 
M3203 diff_1471_625# diff_1471_625# diff_1471_625# GND efet w=3 l=21
+ ad=0 pd=0 as=0 ps=0 
M3204 GND diff_1654_625# diff_1531_577# GND efet w=38 l=17
+ ad=0 pd=0 as=0 ps=0 
M3205 diff_2426_1021# diff_2407_757# diff_2378_1045# GND efet w=98 l=20
+ ad=2600 pd=252 as=0 ps=0 
M3206 GND diff_2452_1015# diff_2426_1021# GND efet w=100 l=19
+ ad=0 pd=0 as=0 ps=0 
M3207 diff_2714_1150# Vdd Vdd GND efet w=19 l=148
+ ad=0 pd=0 as=0 ps=0 
M3208 Vdd Vdd diff_1027_631# GND efet w=22 l=92
+ ad=0 pd=0 as=3629 ps=324 
M3209 diff_2600_1012# diff_2452_1015# diff_2185_1084# GND efet w=76 l=19
+ ad=1976 pd=204 as=3098 ps=282 
M3210 diff_2642_1015# diff_2626_631# diff_2600_1012# GND efet w=74 l=17
+ ad=1790 pd=204 as=0 ps=0 
M3211 GND clk2 diff_2642_1015# GND efet w=56 l=20
+ ad=0 pd=0 as=0 ps=0 
M3212 diff_2185_1084# Vdd Vdd GND efet w=19 l=184
+ ad=0 pd=0 as=0 ps=0 
M3213 GND diff_1960_562# diff_1027_631# GND efet w=53 l=23
+ ad=0 pd=0 as=0 ps=0 
M3214 diff_1195_823# diff_1375_760# GND GND efet w=37 l=16
+ ad=0 pd=0 as=0 ps=0 
M3215 GND diff_1471_625# diff_1195_823# GND efet w=37 l=16
+ ad=0 pd=0 as=0 ps=0 
M3216 clk2 GND GND GND efet w=262 l=19
+ ad=31430 pd=2274 as=0 ps=0 
M3217 diff_2797_1142# Vdd Vdd GND efet w=19 l=145
+ ad=0 pd=0 as=0 ps=0 
M3218 Vdd Vdd diff_2929_1138# GND efet w=19 l=181
+ ad=0 pd=0 as=0 ps=0 
M3219 diff_2407_1684# diff_2929_1138# GND GND efet w=85 l=19
+ ad=3672 pd=386 as=0 ps=0 
M3220 diff_2377_1729# diff_2377_1729# diff_2377_1729# GND efet w=7 l=7
+ ad=0 pd=0 as=0 ps=0 
M3221 diff_2377_1729# diff_2407_1684# GND GND efet w=106 l=19
+ ad=0 pd=0 as=0 ps=0 
M3222 diff_4102_1499# diff_3971_1525# GND GND efet w=100 l=16
+ ad=0 pd=0 as=0 ps=0 
M3223 diff_4231_1556# diff_4231_1556# diff_4231_1556# GND efet w=4 l=7
+ ad=0 pd=0 as=0 ps=0 
M3224 diff_4345_1120# diff_4231_1556# GND GND efet w=79 l=16
+ ad=0 pd=0 as=0 ps=0 
M3225 Vdd Vdd Vdd GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M3226 Vdd Vdd Vdd GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M3227 Vdd diff_5311_1888# diff_2113_3589# GND efet w=53 l=14
+ ad=0 pd=0 as=0 ps=0 
M3228 Vdd Vdd Vdd GND efet w=2 l=5
+ ad=0 pd=0 as=0 ps=0 
M3229 diff_5470_1585# Vdd Vdd GND efet w=25 l=91
+ ad=0 pd=0 as=0 ps=0 
M3230 Vdd Vdd Vdd GND efet w=6 l=9
+ ad=0 pd=0 as=0 ps=0 
M3231 Vdd Vdd diff_5428_2056# GND efet w=25 l=67
+ ad=0 pd=0 as=4788 ps=446 
M3232 diff_5470_1585# clk1 diff_6046_2134# GND efet w=34 l=16
+ ad=0 pd=0 as=1452 ps=164 
M3233 GND diff_6046_2134# diff_2626_631# GND efet w=125 l=14
+ ad=0 pd=0 as=12714 ps=1480 
M3234 Vdd Vdd diff_5308_1972# GND efet w=19 l=16
+ ad=0 pd=0 as=1294 ps=184 
M3235 diff_2113_3589# diff_5428_2056# GND GND efet w=49 l=13
+ ad=0 pd=0 as=0 ps=0 
M3236 diff_5428_2056# diff_5428_2056# diff_5428_2056# GND efet w=5 l=12
+ ad=0 pd=0 as=0 ps=0 
M3237 diff_5308_1972# diff_5308_1972# diff_5308_1972# GND efet w=5 l=12
+ ad=0 pd=0 as=0 ps=0 
M3238 diff_5308_1972# diff_5308_1972# diff_5308_1972# GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M3239 diff_5491_1889# clk2 diff_5428_2056# GND efet w=128 l=14
+ ad=8309 pd=636 as=0 ps=0 
M3240 diff_5428_2056# diff_5428_2056# diff_5428_2056# GND efet w=3 l=7
+ ad=0 pd=0 as=0 ps=0 
M3241 GND diff_5428_2056# diff_5311_1888# GND efet w=55 l=16
+ ad=0 pd=0 as=7421 ps=828 
M3242 Vdd diff_5308_1972# diff_5311_1888# GND efet w=22 l=64
+ ad=0 pd=0 as=0 ps=0 
M3243 Vdd Vdd Vdd GND efet w=5 l=8
+ ad=0 pd=0 as=0 ps=0 
M3244 Vdd Vdd Vdd GND efet w=8 l=16
+ ad=0 pd=0 as=0 ps=0 
M3245 diff_2626_631# Vdd Vdd GND efet w=25 l=46
+ ad=0 pd=0 as=0 ps=0 
M3246 GND diff_2626_631# diff_5491_1889# GND efet w=178 l=16
+ ad=0 pd=0 as=0 ps=0 
M3247 diff_2626_631# diff_2626_631# diff_2626_631# GND efet w=3 l=12
+ ad=0 pd=0 as=0 ps=0 
M3248 diff_2626_631# diff_2626_631# diff_2626_631# GND efet w=7 l=10
+ ad=0 pd=0 as=0 ps=0 
M3249 diff_2626_631# clk2 diff_6037_1948# GND efet w=34 l=14
+ ad=0 pd=0 as=1503 ps=158 
M3250 diff_5311_1888# diff_5308_1972# diff_5311_1888# GND efet w=130 l=45
+ ad=0 pd=0 as=0 ps=0 
M3251 GND diff_6037_1948# diff_1960_562# GND efet w=128 l=14
+ ad=0 pd=0 as=6497 ps=572 
M3252 Vdd Vdd Vdd GND efet w=3 l=7
+ ad=0 pd=0 as=0 ps=0 
M3253 diff_5491_1889# diff_1786_2191# GND GND efet w=115 l=16
+ ad=0 pd=0 as=0 ps=0 
M3254 GND diff_5266_1684# diff_5305_1636# GND efet w=253 l=16
+ ad=0 pd=0 as=9458 ps=806 
M3255 Vdd Vdd Vdd GND efet w=6 l=18
+ ad=0 pd=0 as=0 ps=0 
M3256 diff_1960_562# Vdd Vdd GND efet w=25 l=46
+ ad=0 pd=0 as=0 ps=0 
M3257 diff_1960_562# clk1 diff_5992_1762# GND efet w=34 l=16
+ ad=0 pd=0 as=1461 ps=164 
M3258 diff_5482_1601# diff_5089_1069# GND GND efet w=199 l=16
+ ad=12215 pd=928 as=0 ps=0 
M3259 Vdd Vdd Vdd GND efet w=3 l=5
+ ad=0 pd=0 as=0 ps=0 
M3260 GND diff_5992_1762# diff_2203_2482# GND efet w=124 l=16
+ ad=0 pd=0 as=6239 ps=548 
M3261 Vdd Vdd Vdd GND efet w=5 l=10
+ ad=0 pd=0 as=0 ps=0 
M3262 diff_2203_2482# Vdd Vdd GND efet w=25 l=46
+ ad=0 pd=0 as=0 ps=0 
M3263 diff_5482_1601# diff_4759_1004# GND GND efet w=196 l=16
+ ad=0 pd=0 as=0 ps=0 
M3264 diff_4720_1750# clk1 diff_5305_1636# GND efet w=190 l=16
+ ad=5525 pd=456 as=0 ps=0 
M3265 diff_4720_1633# Vdd Vdd GND efet w=19 l=16
+ ad=0 pd=0 as=0 ps=0 
M3266 Vdd Vdd Vdd GND efet w=8 l=23
+ ad=0 pd=0 as=0 ps=0 
M3267 diff_4477_1126# diff_4231_1556# GND GND efet w=74 l=17
+ ad=0 pd=0 as=0 ps=0 
M3268 Vdd Vdd Vdd GND efet w=13 l=9
+ ad=0 pd=0 as=0 ps=0 
M3269 GND diff_3722_1087# diff_4477_1126# GND efet w=74 l=16
+ ad=0 pd=0 as=0 ps=0 
M3270 diff_4345_1120# diff_3587_1105# GND GND efet w=77 l=17
+ ad=0 pd=0 as=0 ps=0 
M3271 diff_5018_1444# Vdd Vdd GND efet w=17 l=17
+ ad=1432 pd=182 as=0 ps=0 
M3272 diff_5018_1444# diff_5018_1444# diff_5018_1444# GND efet w=2 l=9
+ ad=0 pd=0 as=0 ps=0 
M3273 diff_5018_1444# diff_5018_1444# diff_5018_1444# GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M3274 diff_550_2356# diff_5018_1444# diff_550_2356# GND efet w=167 l=56
+ ad=24980 pd=2684 as=0 ps=0 
M3275 diff_4720_1750# Vdd Vdd GND efet w=22 l=46
+ ad=0 pd=0 as=0 ps=0 
M3276 diff_5482_1601# diff_5470_1585# diff_5266_1684# GND efet w=164 l=17
+ ad=0 pd=0 as=4523 ps=388 
M3277 diff_1786_2191# diff_5206_1351# diff_1786_2191# GND efet w=162 l=82
+ ad=21167 pd=2300 as=0 ps=0 
M3278 diff_550_2356# diff_5018_1444# Vdd GND efet w=22 l=25
+ ad=0 pd=0 as=0 ps=0 
M3279 GND diff_3962_1084# diff_4345_1120# GND efet w=58 l=26
+ ad=0 pd=0 as=0 ps=0 
M3280 GND diff_965_1612# diff_3346_1166# GND efet w=32 l=17
+ ad=0 pd=0 as=1643 ps=168 
M3281 diff_2407_1684# diff_2407_1684# diff_2407_1684# GND efet w=4 l=7
+ ad=0 pd=0 as=0 ps=0 
M3282 diff_2407_1684# diff_2407_1684# diff_2407_1684# GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M3283 GND diff_3175_1156# diff_2377_1729# GND efet w=88 l=16
+ ad=0 pd=0 as=0 ps=0 
M3284 diff_4019_1288# diff_2128_1144# diff_580_3394# GND efet w=31 l=16
+ ad=1246 pd=178 as=0 ps=0 
M3285 diff_4019_1288# diff_4019_1288# diff_4019_1288# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M3286 diff_4019_1288# diff_4019_1288# diff_4019_1288# GND efet w=6 l=7
+ ad=0 pd=0 as=0 ps=0 
M3287 GND diff_3790_1090# diff_4477_1126# GND efet w=74 l=17
+ ad=0 pd=0 as=0 ps=0 
M3288 diff_4477_1126# diff_4019_1288# GND GND efet w=125 l=17
+ ad=0 pd=0 as=0 ps=0 
M3289 GND diff_3461_1093# diff_4477_1126# GND efet w=59 l=17
+ ad=0 pd=0 as=0 ps=0 
M3290 Vdd Vdd diff_5206_1351# GND efet w=17 l=17
+ ad=0 pd=0 as=1414 ps=194 
M3291 diff_5266_1684# Vdd Vdd GND efet w=23 l=68
+ ad=0 pd=0 as=0 ps=0 
M3292 diff_2203_2482# clk2 diff_6004_1579# GND efet w=34 l=13
+ ad=0 pd=0 as=1494 ps=158 
M3293 GND diff_6004_1579# diff_5089_1069# GND efet w=101 l=14
+ ad=0 pd=0 as=23254 ps=2866 
M3294 Vdd Vdd Vdd GND efet w=2 l=4
+ ad=0 pd=0 as=0 ps=0 
M3295 Vdd Vdd Vdd GND efet w=4 l=5
+ ad=0 pd=0 as=0 ps=0 
M3296 diff_5089_1069# Vdd Vdd GND efet w=26 l=68
+ ad=0 pd=0 as=0 ps=0 
M3297 diff_5206_1351# diff_5206_1351# diff_5206_1351# GND efet w=2 l=12
+ ad=0 pd=0 as=0 ps=0 
M3298 diff_5206_1351# diff_5206_1351# diff_5206_1351# GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M3299 Vdd Vdd Vdd GND efet w=11 l=23
+ ad=0 pd=0 as=0 ps=0 
M3300 Vdd Vdd Vdd GND efet w=5 l=23
+ ad=0 pd=0 as=0 ps=0 
M3301 diff_5089_1069# clk1 diff_5947_1387# GND efet w=32 l=13
+ ad=0 pd=0 as=1329 ps=152 
M3302 Vdd Vdd diff_5188_6931# GND efet w=23 l=46
+ ad=0 pd=0 as=20436 ps=2072 
M3303 Vdd diff_5206_1351# diff_1786_2191# GND efet w=22 l=46
+ ad=0 pd=0 as=0 ps=0 
M3304 diff_550_2356# diff_4936_1297# GND GND efet w=187 l=16
+ ad=0 pd=0 as=0 ps=0 
M3305 diff_1786_2191# diff_4936_1297# GND GND efet w=113 l=14
+ ad=0 pd=0 as=0 ps=0 
M3306 Vdd Vdd diff_5179_1243# GND efet w=22 l=67
+ ad=0 pd=0 as=3686 ps=362 
M3307 GND diff_5947_1387# diff_2407_757# GND efet w=131 l=14
+ ad=0 pd=0 as=15771 ps=1626 
M3308 Vdd Vdd Vdd GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M3309 Vdd Vdd Vdd GND efet w=8 l=17
+ ad=0 pd=0 as=0 ps=0 
M3310 diff_2407_757# Vdd Vdd GND efet w=25 l=46
+ ad=0 pd=0 as=0 ps=0 
M3311 diff_5188_6931# diff_4936_1297# GND GND efet w=142 l=16
+ ad=0 pd=0 as=0 ps=0 
M3312 diff_3346_1166# diff_2128_1144# Vdd GND efet w=34 l=17
+ ad=0 pd=0 as=0 ps=0 
M3313 diff_2407_1684# Vdd Vdd GND efet w=23 l=71
+ ad=0 pd=0 as=0 ps=0 
M3314 diff_2377_1729# Vdd Vdd GND efet w=25 l=76
+ ad=0 pd=0 as=0 ps=0 
M3315 diff_3175_1156# diff_1960_562# GND GND efet w=92 l=23
+ ad=2147 pd=220 as=0 ps=0 
M3316 diff_3461_1093# diff_3346_1166# GND GND efet w=155 l=17
+ ad=4247 pd=402 as=0 ps=0 
M3317 diff_3587_1105# diff_3562_1297# GND GND efet w=121 l=16
+ ad=4737 pd=418 as=0 ps=0 
M3318 diff_3587_1105# diff_3587_1105# diff_3587_1105# GND efet w=7 l=7
+ ad=0 pd=0 as=0 ps=0 
M3319 diff_3722_1087# diff_3587_1105# GND GND efet w=79 l=19
+ ad=0 pd=0 as=0 ps=0 
M3320 diff_4483_1244# diff_4019_1288# GND GND efet w=121 l=16
+ ad=9820 pd=968 as=0 ps=0 
M3321 GND diff_4676_991# diff_550_2356# GND efet w=178 l=16
+ ad=0 pd=0 as=0 ps=0 
M3322 GND diff_5179_1243# diff_1786_2191# GND efet w=106 l=16
+ ad=0 pd=0 as=0 ps=0 
M3323 diff_3722_1087# diff_3722_1087# diff_3722_1087# GND efet w=5 l=12
+ ad=0 pd=0 as=0 ps=0 
M3324 GND diff_3709_1297# diff_3790_1090# GND efet w=110 l=17
+ ad=0 pd=0 as=5319 ps=492 
M3325 diff_3587_1105# diff_3587_1105# diff_3587_1105# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M3326 Vdd Vdd diff_3175_1156# GND efet w=23 l=74
+ ad=0 pd=0 as=0 ps=0 
M3327 diff_3461_1093# Vdd Vdd GND efet w=22 l=70
+ ad=0 pd=0 as=0 ps=0 
M3328 diff_3722_1087# diff_3722_1087# diff_3722_1087# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M3329 diff_3790_1090# diff_3790_1090# diff_3790_1090# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M3330 diff_3962_1084# diff_3790_1090# GND GND efet w=82 l=19
+ ad=0 pd=0 as=0 ps=0 
M3331 GND diff_4019_1288# diff_4066_1042# GND efet w=112 l=16
+ ad=0 pd=0 as=4434 ps=424 
M3332 diff_3962_1084# diff_3962_1084# diff_3962_1084# GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M3333 diff_3587_1105# Vdd Vdd GND efet w=22 l=94
+ ad=0 pd=0 as=0 ps=0 
M3334 diff_3790_1090# diff_3790_1090# diff_3790_1090# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M3335 diff_3962_1084# diff_3962_1084# diff_3962_1084# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M3336 diff_1744_715# diff_4066_1042# GND GND efet w=61 l=16
+ ad=6936 pd=680 as=0 ps=0 
M3337 GND diff_3461_1093# diff_1744_715# GND efet w=80 l=16
+ ad=0 pd=0 as=0 ps=0 
M3338 diff_1744_715# diff_4345_1120# GND GND efet w=61 l=19
+ ad=0 pd=0 as=0 ps=0 
M3339 GND diff_3461_1093# diff_4483_1244# GND efet w=76 l=16
+ ad=0 pd=0 as=0 ps=0 
M3340 diff_4483_1244# diff_4477_1126# GND GND efet w=77 l=23
+ ad=0 pd=0 as=0 ps=0 
M3341 diff_1744_715# diff_1744_715# diff_1744_715# GND efet w=4 l=5
+ ad=0 pd=0 as=0 ps=0 
M3342 diff_4066_1042# diff_4066_1042# diff_4066_1042# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M3343 diff_1744_715# diff_1744_715# diff_1744_715# GND efet w=4 l=5
+ ad=0 pd=0 as=0 ps=0 
M3344 diff_3722_1087# Vdd Vdd GND efet w=25 l=70
+ ad=0 pd=0 as=0 ps=0 
M3345 diff_4066_1042# diff_4066_1042# diff_4066_1042# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M3346 diff_3962_1084# Vdd Vdd GND efet w=23 l=76
+ ad=0 pd=0 as=0 ps=0 
M3347 Vdd Vdd diff_4066_1042# GND efet w=25 l=97
+ ad=0 pd=0 as=0 ps=0 
M3348 Vdd Vdd diff_3790_1090# GND efet w=22 l=97
+ ad=0 pd=0 as=0 ps=0 
M3349 diff_1744_715# Vdd Vdd GND efet w=22 l=94
+ ad=0 pd=0 as=0 ps=0 
M3350 GND diff_5179_1243# diff_5188_6931# GND efet w=133 l=16
+ ad=0 pd=0 as=0 ps=0 
M3351 diff_4936_1297# diff_4481_442# GND GND efet w=76 l=16
+ ad=3740 pd=396 as=0 ps=0 
M3352 GND diff_5089_1069# diff_550_2356# GND efet w=146 l=30
+ ad=0 pd=0 as=0 ps=0 
M3353 diff_1786_2191# diff_4759_1004# GND GND efet w=109 l=16
+ ad=0 pd=0 as=0 ps=0 
M3354 GND diff_4345_1120# diff_4483_1244# GND efet w=62 l=17
+ ad=0 pd=0 as=0 ps=0 
M3355 GND diff_4483_1244# diff_4759_1004# GND efet w=52 l=16
+ ad=0 pd=0 as=2858 ps=252 
M3356 GND diff_2407_757# diff_5179_1243# GND efet w=94 l=16
+ ad=0 pd=0 as=0 ps=0 
M3357 diff_5188_6931# diff_4879_1024# GND GND efet w=140 l=17
+ ad=0 pd=0 as=0 ps=0 
M3358 GND diff_4477_1126# diff_4879_1024# GND efet w=52 l=16
+ ad=0 pd=0 as=2450 ps=246 
M3359 diff_4483_1244# Vdd Vdd GND efet w=22 l=91
+ ad=0 pd=0 as=0 ps=0 
M3360 diff_4676_991# diff_1744_715# GND GND efet w=49 l=19
+ ad=3071 pd=240 as=0 ps=0 
M3361 Vdd Vdd diff_4676_991# GND efet w=25 l=124
+ ad=0 pd=0 as=0 ps=0 
M3362 Vdd Vdd diff_4759_1004# GND efet w=25 l=115
+ ad=0 pd=0 as=0 ps=0 
M3363 diff_4879_1024# Vdd Vdd GND efet w=25 l=115
+ ad=0 pd=0 as=0 ps=0 
M3364 diff_4936_1297# Vdd Vdd GND efet w=16 l=56
+ ad=0 pd=0 as=0 ps=0 
M3365 diff_2407_757# clk2 diff_5959_1177# GND efet w=34 l=13
+ ad=0 pd=0 as=1419 ps=152 
M3366 Vdd Vdd Vdd GND efet w=2 l=4
+ ad=0 pd=0 as=0 ps=0 
M3367 diff_5897_1123# Vdd Vdd GND efet w=26 l=137
+ ad=4222 pd=412 as=0 ps=0 
M3368 GND diff_5959_1177# diff_5897_1123# GND efet w=43 l=16
+ ad=0 pd=0 as=0 ps=0 
M3369 Vdd Vdd Vdd GND efet w=5 l=7
+ ad=0 pd=0 as=0 ps=0 
M3370 diff_5897_1123# clk1 diff_5947_1054# GND efet w=31 l=16
+ ad=0 pd=0 as=1302 ps=146 
M3371 GND diff_5947_1054# diff_1654_625# GND efet w=125 l=14
+ ad=0 pd=0 as=5099 ps=438 
M3372 Vdd Vdd Vdd GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M3373 Vdd Vdd Vdd GND efet w=6 l=7
+ ad=0 pd=0 as=0 ps=0 
M3374 Vdd Vdd Vdd GND efet w=5 l=12
+ ad=0 pd=0 as=0 ps=0 
M3375 Vdd Vdd Vdd GND efet w=2 l=2
+ ad=0 pd=0 as=0 ps=0 
M3376 diff_4481_442# Vdd Vdd GND efet w=25 l=47
+ ad=15713 pd=1386 as=0 ps=0 
M3377 Vdd Vdd diff_2452_1015# GND efet w=25 l=67
+ ad=0 pd=0 as=4547 ps=438 
M3378 diff_1654_625# Vdd Vdd GND efet w=25 l=47
+ ad=0 pd=0 as=0 ps=0 
M3379 Vdd Vdd diff_5359_406# GND efet w=31 l=110
+ ad=0 pd=0 as=5340 ps=482 
M3380 diff_4481_442# reset GND GND efet w=313 l=16
+ ad=0 pd=0 as=0 ps=0 
M3381 sync GND GND GND efet w=262 l=19
+ ad=0 pd=0 as=0 ps=0 
M3382 reset GND GND GND efet w=268 l=19
+ ad=20616 pd=1936 as=0 ps=0 
M3383 GND GND p0 GND efet w=262 l=19
+ ad=0 pd=0 as=18030 ps=1876 
M3384 diff_5359_406# diff_5359_406# diff_5359_406# GND efet w=5 l=5
+ ad=0 pd=0 as=0 ps=0 
M3385 diff_5359_406# diff_5359_406# diff_5359_406# GND efet w=3 l=10
+ ad=0 pd=0 as=0 ps=0 
M3386 diff_2452_1015# diff_5359_406# GND GND efet w=94 l=13
+ ad=0 pd=0 as=0 ps=0 
M3387 GND cm diff_5359_406# GND efet w=124 l=16
+ ad=0 pd=0 as=0 ps=0 
M3388 cm GND GND GND efet w=263 l=17
+ ad=19623 pd=1948 as=0 ps=0 
C0 metal_6031_103# gnd! 245.1fF ;**FLOATING
C1 metal_5893_124# gnd! 263.4fF ;**FLOATING
C2 metal_5755_130# gnd! 276.8fF ;**FLOATING
C3 metal_5617_157# gnd! 243.7fF ;**FLOATING
C4 metal_1741_139# gnd! 35.8fF ;**FLOATING
C5 metal_1690_160# gnd! 19.8fF ;**FLOATING
C6 metal_1651_193# gnd! 59.3fF ;**FLOATING
C7 metal_1687_193# gnd! 147.4fF ;**FLOATING
C8 metal_1795_280# gnd! 426.1fF ;**FLOATING
C9 metal_1651_319# gnd! 8.0fF ;**FLOATING
C10 metal_391_406# gnd! 48.9fF ;**FLOATING
C11 metal_5887_7378# gnd! 313.1fF ;**FLOATING
C12 diff_5359_406# gnd! 730.2fF
C13 cm gnd! 7259.6fF
C14 reset gnd! 5467.7fF
C15 diff_5947_1054# gnd! 398.1fF
C16 diff_5897_1123# gnd! 463.4fF
C17 diff_5959_1177# gnd! 341.9fF
C18 diff_4879_1024# gnd! 1038.1fF
C19 diff_4066_1042# gnd! 768.2fF
C20 diff_4676_991# gnd! 937.2fF
C21 diff_4483_1244# gnd! 1695.7fF
C22 diff_5179_1243# gnd! 766.7fF
C23 diff_4936_1297# gnd! 1042.2fF
C24 diff_5947_1387# gnd! 379.9fF
C25 diff_6004_1579# gnd! 365.5fF
C26 diff_3346_1166# gnd! 577.2fF
C27 diff_3175_1156# gnd! 542.6fF
C28 diff_3461_1093# gnd! 1921.2fF
C29 diff_4019_1288# gnd! 1166.7fF
C30 diff_3790_1090# gnd! 1557.0fF
C31 diff_5206_1351# gnd! 722.5fF
C32 diff_3587_1105# gnd! 1562.5fF
C33 diff_5018_1444# gnd! 676.5fF
C34 diff_4759_1004# gnd! 1833.2fF
C35 diff_5992_1762# gnd! 401.0fF
C36 diff_5089_1069# gnd! 4413.2fF
C37 diff_5482_1601# gnd! 1457.3fF
C38 diff_5305_1636# gnd! 1026.4fF
C39 diff_5266_1684# gnd! 998.5fF
C40 diff_6037_1948# gnd! 393.6fF
C41 diff_5491_1889# gnd! 1067.3fF
C42 diff_5308_1972# gnd! 689.7fF
C43 diff_5428_2056# gnd! 747.9fF
C44 diff_6046_2134# gnd! 387.9fF
C45 diff_5311_1888# gnd! 1323.0fF
C46 diff_4477_1126# gnd! 2066.4fF
C47 diff_3709_1297# gnd! 511.8fF
C48 diff_2642_1015# gnd! 199.4fF
C49 diff_2600_1012# gnd! 218.0fF
C50 diff_2626_631# gnd! 6052.8fF
C51 diff_2426_1021# gnd! 285.2fF
C52 diff_1471_625# gnd! 747.8fF
C53 diff_1531_577# gnd! 613.4fF
C54 diff_1744_715# gnd! 3882.6fF
C55 diff_1568_757# gnd! 184.1fF
C56 diff_409_424# gnd! 68.9fF ;**FLOATING
C57 diff_397_451# gnd! 103.2fF ;**FLOATING
C58 diff_388_469# gnd! 583.6fF ;**FLOATING
C59 diff_1375_760# gnd! 783.2fF
C60 diff_2378_1045# gnd! 296.9fF
C61 diff_2407_757# gnd! 6100.6fF
C62 diff_2185_1084# gnd! 777.0fF
C63 diff_2929_1181# gnd! 188.6fF
C64 diff_1654_625# gnd! 4803.9fF
C65 diff_2929_1223# gnd! 217.7fF
C66 diff_2797_1142# gnd! 459.6fF
C67 diff_2929_1138# gnd! 722.0fF
C68 diff_3562_1297# gnd! 436.1fF
C69 diff_4345_1120# gnd! 1489.6fF
C70 diff_3971_1525# gnd! 404.2fF
C71 diff_4102_1499# gnd! 678.3fF
C72 diff_2452_1015# gnd! 4705.4fF
C73 diff_2714_1150# gnd! 736.7fF
C74 diff_2128_1144# gnd! 3205.1fF
C75 diff_5470_1585# gnd! 3169.8fF
C76 diff_4720_1633# gnd! 622.1fF
C77 diff_4720_1750# gnd! 1288.4fF
C78 diff_5017_1867# gnd! 496.6fF
C79 diff_4909_1861# gnd! 559.9fF
C80 diff_4633_1837# gnd! 547.9fF
C81 diff_4663_1771# gnd! 567.3fF
C82 diff_4852_1946# gnd! 529.8fF
C83 diff_4687_1963# gnd! 1158.3fF
C84 diff_4666_1904# gnd! 1380.3fF
C85 diff_4327_1867# gnd! 492.1fF
C86 diff_4477_1730# gnd! 821.8fF
C87 diff_4222_1852# gnd! 542.2fF
C88 diff_1027_631# gnd! 1411.0fF
C89 diff_1036_647# gnd! 296.6fF
C90 diff_916_577# gnd! 584.9fF
C91 diff_1153_682# gnd! 569.2fF
C92 diff_1195_823# gnd! 1090.1fF
C93 diff_847_706# gnd! 666.8fF
C94 diff_2026_1181# gnd! 1045.2fF
C95 diff_1942_1112# gnd! 576.7fF
C96 diff_1642_1000# gnd! 607.6fF
C97 diff_1825_1156# gnd! 707.4fF
C98 p0 gnd! 8683.7fF
C99 diff_778_1165# gnd! 512.0fF
C100 diff_769_1192# gnd! 392.8fF
C101 diff_892_1207# gnd! 395.3fF
C102 diff_1859_1291# gnd! 760.9fF
C103 diff_883_1234# gnd! 284.4fF
C104 diff_715_1141# gnd! 372.1fF
C105 diff_1378_1321# gnd! 679.2fF
C106 diff_1513_1009# gnd! 1214.4fF
C107 diff_1834_1103# gnd! 1122.3fF
C108 diff_1582_1201# gnd! 1829.2fF
C109 diff_892_1357# gnd! 431.9fF
C110 diff_1387_1249# gnd! 2639.4fF
C111 diff_886_1384# gnd! 281.9fF
C112 diff_1387_1337# gnd! 1164.0fF
C113 diff_892_1507# gnd! 403.7fF
C114 diff_2407_1684# gnd! 3030.7fF
C115 diff_3973_1771# gnd! 579.7fF
C116 diff_3946_1780# gnd! 537.7fF
C117 diff_4543_1856# gnd! 694.1fF
C118 diff_4162_1949# gnd! 525.5fF
C119 diff_4000_1963# gnd! 2138.2fF
C120 diff_3976_1904# gnd! 2119.7fF
C121 diff_3781_1697# gnd! 831.9fF
C122 diff_3637_1879# gnd! 521.5fF
C123 diff_3532_1855# gnd! 587.1fF
C124 diff_3259_1780# gnd! 541.9fF
C125 diff_3286_1771# gnd! 596.4fF
C126 diff_3853_1856# gnd! 699.5fF
C127 diff_6091_2320# gnd! 347.7fF
C128 diff_3475_1949# gnd! 517.9fF
C129 diff_3313_1963# gnd! 2172.1fF
C130 diff_3289_1904# gnd! 2117.5fF
C131 diff_3103_1685# gnd! 872.1fF
C132 diff_2950_1870# gnd! 537.4fF
C133 diff_2845_1858# gnd! 585.8fF
C134 diff_2599_1771# gnd! 625.7fF
C135 diff_2569_1822# gnd! 553.6fF
C136 diff_3166_1856# gnd! 639.3fF
C137 diff_3962_1084# gnd! 3264.8fF
C138 diff_2785_1949# gnd! 550.5fF
C139 diff_2626_1963# gnd! 2181.1fF
C140 diff_2599_2041# gnd! 2156.4fF
C141 diff_2416_1697# gnd! 845.8fF
C142 diff_2263_1867# gnd! 536.2fF
C143 diff_2158_1852# gnd! 588.2fF
C144 diff_886_1528# gnd! 310.8fF
C145 diff_949_1603# gnd! 420.6fF
C146 diff_1912_1771# gnd! 593.2fF
C147 diff_1361_1756# gnd! 521.3fF
C148 diff_944_1837# gnd! 332.8fF
C149 sync gnd! 9291.7fF
C150 diff_1888_1780# gnd! 476.2fF
C151 diff_2377_1729# gnd! 3986.7fF
C152 diff_2479_1856# gnd! 640.2fF
C153 diff_989_1735# gnd! 1199.6fF
C154 diff_1358_1843# gnd! 1619.7fF
C155 diff_2098_1949# gnd! 567.5fF
C156 diff_1939_1963# gnd! 2165.2fF
C157 diff_1912_2041# gnd! 2128.2fF
C158 diff_965_1612# gnd! 4723.8fF
C159 diff_3722_1087# gnd! 3270.4fF
C160 diff_4684_2065# gnd! 1627.7fF
C161 diff_4231_1556# gnd! 2503.3fF
C162 diff_3997_2065# gnd! 2131.8fF
C163 diff_3310_2065# gnd! 1407.1fF
C164 diff_10_2008# gnd! 10514.5fF ;**FLOATING
C165 diff_595_2158# gnd! 616.4fF
C166 diff_4462_2026# gnd! 1978.6fF
C167 diff_3577_2338# gnd! 1589.1fF
C168 diff_2608_2057# gnd! 3989.4fF
C169 diff_1921_2057# gnd! 4225.4fF
C170 diff_2890_2341# gnd! 1545.5fF
C171 diff_2203_2368# gnd! 1610.0fF
C172 diff_6091_2533# gnd! 380.3fF
C173 diff_4447_2516# gnd! 452.9fF
C174 diff_4252_2516# gnd! 344.0fF
C175 diff_4435_2500# gnd! 1172.8fF
C176 diff_5987_2827# gnd! 735.2fF
C177 diff_4699_2554# gnd! 1139.3fF
C178 diff_2122_2422# gnd! 5998.2fF
C179 diff_5053_2732# gnd! 846.2fF
C180 diff_2203_2482# gnd! 5880.4fF
C181 diff_4927_2758# gnd! 798.6fF
C182 diff_4726_2803# gnd! 863.8fF
C183 diff_4549_2758# gnd! 759.2fF
C184 diff_4417_2732# gnd! 765.8fF
C185 diff_4237_2758# gnd! 761.4fF
C186 diff_4084_2797# gnd! 859.2fF
C187 diff_3505_2438# gnd! 902.5fF
C188 diff_3892_2761# gnd! 835.8fF
C189 diff_3742_2791# gnd! 861.9fF
C190 diff_5821_2920# gnd! 593.2fF
C191 diff_4243_2545# gnd! 1879.4fF
C192 diff_3550_2758# gnd! 851.7fF
C193 diff_3397_2791# gnd! 861.9fF
C194 diff_3205_2761# gnd! 830.8fF
C195 diff_3055_2803# gnd! 848.8fF
C196 diff_2818_2438# gnd! 966.2fF
C197 diff_2863_2758# gnd! 850.2fF
C198 diff_2710_2797# gnd! 866.3fF
C199 diff_2521_2758# gnd! 840.4fF
C200 diff_2371_2794# gnd! 843.4fF
C201 diff_2062_2569# gnd! 829.6fF
C202 diff_1436_2665# gnd! 770.1fF
C203 diff_550_2479# gnd! 1030.0fF
C204 diff_562_2665# gnd! 811.4fF
C205 diff_1405_2629# gnd! 686.5fF
C206 diff_2176_2758# gnd! 870.4fF
C207 diff_508_1279# gnd! 3676.4fF
C208 diff_2023_2797# gnd! 862.1fF
C209 diff_1436_2722# gnd! 758.0fF
C210 diff_1417_2311# gnd! 4280.1fF
C211 diff_622_2720# gnd! 370.0fF
C212 diff_550_2755# gnd! 385.8fF
C213 diff_4723_3052# gnd! 2160.5fF
C214 diff_5848_3025# gnd! 970.9fF
C215 diff_2209_3019# gnd! 3284.1fF
C216 diff_2056_3070# gnd! 3435.0fF
C217 diff_4936_3115# gnd! 1557.3fF
C218 diff_5771_2965# gnd! 834.2fF
C219 diff_2101_2551# gnd! 4306.0fF
C220 diff_4903_3178# gnd! 1895.4fF
C221 diff_1291_3103# gnd! 1597.4fF
C222 diff_4756_3238# gnd! 1610.7fF
C223 diff_5762_3178# gnd! 681.2fF
C224 diff_2056_3184# gnd! 3537.1fF
C225 diff_1291_3169# gnd! 1809.2fF
C226 diff_2743_3241# gnd! 3446.8fF
C227 diff_5191_3280# gnd! 815.0fF
C228 diff_2056_3301# gnd! 3343.8fF
C229 diff_1291_3280# gnd! 1160.6fF
C230 diff_1829_3133# gnd! 522.6fF
C231 diff_550_2356# gnd! 9035.2fF
C232 diff_5837_3124# gnd! 1085.5fF
C233 diff_5776_3412# gnd! 1393.4fF
C234 diff_1960_562# gnd! 7529.9fF
C235 diff_5875_3626# gnd! 679.9fF
C236 diff_673_1115# gnd! 8732.3fF
C237 diff_2062_3349# gnd! 2942.2fF
C238 diff_3254_2623# gnd! 2511.0fF
C239 diff_1291_3346# gnd! 1713.1fF
C240 diff_425_3187# gnd! 1320.8fF
C241 diff_5134_2953# gnd! 2244.2fF
C242 diff_5029_3068# gnd! 2271.8fF
C243 diff_5266_3691# gnd! 659.3fF
C244 diff_4915_3191# gnd! 1954.5fF
C245 diff_4732_2900# gnd! 2011.3fF
C246 diff_5095_3556# gnd! 690.7fF
C247 diff_4921_3691# gnd! 674.8fF
C248 diff_4552_2860# gnd! 2288.6fF
C249 diff_4399_2803# gnd! 2194.6fF
C250 diff_4750_3556# gnd! 723.1fF
C251 diff_4576_3691# gnd! 694.5fF
C252 diff_4231_3628# gnd! 2087.7fF
C253 diff_4087_2900# gnd! 1985.2fF
C254 diff_4405_3556# gnd! 719.3fF
C255 diff_4231_3691# gnd! 719.6fF
C256 diff_3889_3628# gnd! 1993.1fF
C257 diff_3745_2897# gnd! 1854.3fF
C258 diff_4063_3493# gnd! 700.7fF
C259 diff_3889_3691# gnd! 700.8fF
C260 diff_3544_3628# gnd! 1987.7fF
C261 diff_3400_2897# gnd! 1979.4fF
C262 diff_3718_3556# gnd! 722.9fF
C263 diff_3544_3691# gnd! 719.1fF
C264 diff_3376_3475# gnd! 707.6fF
C265 diff_3202_3628# gnd! 1934.5fF
C266 diff_3055_2897# gnd! 1961.1fF
C267 diff_3202_3691# gnd! 718.4fF
C268 diff_2857_3628# gnd! 1972.6fF
C269 diff_2713_2900# gnd! 1970.5fF
C270 diff_3031_3556# gnd! 724.7fF
C271 diff_2857_3691# gnd! 720.6fF
C272 diff_2515_3628# gnd! 1954.2fF
C273 diff_2368_2803# gnd! 1937.0fF
C274 diff_2689_3475# gnd! 720.8fF
C275 diff_2515_3691# gnd! 694.3fF
C276 diff_407_3110# gnd! 1355.3fF
C277 diff_2053_3553# gnd! 9247.3fF
C278 diff_2113_3589# gnd! 9166.3fF
C279 diff_2170_3631# gnd! 1972.5fF
C280 diff_2026_2897# gnd! 1970.1fF
C281 diff_1829_3439# gnd! 593.0fF
C282 diff_1786_2191# gnd! 8302.4fF
C283 diff_2344_3556# gnd! 723.2fF
C284 diff_2170_3691# gnd! 712.2fF
C285 diff_1996_3562# gnd! 749.6fF
C286 diff_5866_3757# gnd! 902.2fF
C287 diff_5849_3703# gnd! 1056.4fF
C288 clk1 gnd! 15700.0fF
C289 diff_5357_3892# gnd! 181.4fF
C290 diff_5855_3847# gnd! 1006.2fF
C291 diff_5294_3844# gnd! 368.5fF
C292 diff_5357_3973# gnd! 182.0fF
C293 diff_5705_4015# gnd! 653.3fF
C294 diff_5129_3880# gnd! 160.1fF
C295 diff_5104_3844# gnd! 371.9fF
C296 diff_4949_3844# gnd! 365.4fF
C297 diff_5012_3892# gnd! 176.3fF
C298 diff_5294_4054# gnd! 363.9fF
C299 diff_5294_4195# gnd! 365.9fF
C300 diff_5357_4246# gnd! 183.8fF
C301 diff_4481_442# gnd! 6414.5fF
C302 diff_5357_4327# gnd! 188.9fF
C303 diff_5129_3982# gnd! 166.7fF
C304 diff_5012_3973# gnd! 183.8fF
C305 diff_5104_4051# gnd! 373.2fF
C306 diff_4784_3877# gnd! 167.0fF
C307 diff_4759_3844# gnd! 387.3fF
C308 diff_4607_3841# gnd! 371.4fF
C309 diff_4667_3892# gnd! 184.1fF
C310 diff_4949_4054# gnd! 361.3fF
C311 diff_5129_4231# gnd! 165.2fF
C312 diff_5104_4198# gnd! 372.2fF
C313 diff_4949_4195# gnd! 366.9fF
C314 diff_5012_4246# gnd! 183.2fF
C315 diff_5294_4411# gnd! 365.2fF
C316 diff_5294_4552# gnd! 370.7fF
C317 diff_5357_4600# gnd! 184.7fF
C318 diff_5357_4684# gnd! 183.2fF
C319 o3 gnd! 6027.5fF
C320 diff_5129_4336# gnd! 166.7fF
C321 diff_5012_4327# gnd! 185.6fF
C322 diff_5104_4405# gnd! 382.0fF
C323 diff_4784_3982# gnd! 168.5fF
C324 diff_4667_3973# gnd! 184.7fF
C325 diff_4759_4051# gnd! 372.5fF
C326 diff_4439_3877# gnd! 169.7fF
C327 diff_4414_3847# gnd! 380.9fF
C328 diff_4325_3892# gnd! 168.8fF
C329 diff_4262_3841# gnd! 370.2fF
C330 diff_4607_4054# gnd! 356.3fF
C331 diff_4784_4231# gnd! 169.7fF
C332 diff_4759_4198# gnd! 373.4fF
C333 diff_4607_4195# gnd! 361.1fF
C334 diff_4667_4246# gnd! 185.0fF
C335 diff_4949_4411# gnd! 368.5fF
C336 diff_5129_4588# gnd! 166.7fF
C337 diff_5012_4600# gnd! 184.7fF
C338 diff_5104_4552# gnd! 370.6fF
C339 diff_4949_4552# gnd! 362.9fF
C340 diff_5294_4765# gnd! 355.0fF
C341 diff_5294_4906# gnd! 357.2fF
C342 diff_5357_4957# gnd! 183.2fF
C343 diff_5938_5011# gnd! 1252.0fF
C344 diff_6137_5167# gnd! 438.2fF
C345 diff_6062_5224# gnd! 385.2fF
C346 diff_5357_5038# gnd! 185.6fF
C347 diff_5129_4690# gnd! 161.6fF
C348 diff_5012_4684# gnd! 185.6fF
C349 diff_5104_4759# gnd! 362.5fF
C350 diff_4784_4336# gnd! 168.5fF
C351 diff_4667_4327# gnd! 186.5fF
C352 diff_4759_4405# gnd! 373.7fF
C353 diff_4439_3982# gnd! 169.4fF
C354 diff_4325_3973# gnd! 169.4fF
C355 diff_4414_4054# gnd! 367.1fF
C356 diff_4094_3877# gnd! 171.2fF
C357 diff_3980_3892# gnd! 167.9fF
C358 diff_4072_3844# gnd! 370.6fF
C359 diff_3917_3841# gnd! 389.2fF
C360 diff_4262_4054# gnd! 349.9fF
C361 diff_4094_3982# gnd! 172.4fF
C362 diff_3980_3973# gnd! 169.4fF
C363 diff_4072_4051# gnd! 359.1fF
C364 diff_4439_4231# gnd! 169.7fF
C365 diff_4414_4198# gnd! 366.4fF
C366 diff_4262_4195# gnd! 358.4fF
C367 diff_4325_4246# gnd! 168.8fF
C368 diff_4607_4411# gnd! 373.3fF
C369 diff_4784_4588# gnd! 169.4fF
C370 diff_4607_4549# gnd! 368.9fF
C371 diff_4667_4600# gnd! 186.5fF
C372 diff_4759_4552# gnd! 371.9fF
C373 diff_4949_4765# gnd! 364.5fF
C374 diff_5129_4942# gnd! 167.0fF
C375 diff_5104_4906# gnd! 360.9fF
C376 diff_5012_4957# gnd! 183.2fF
C377 diff_4949_4906# gnd! 363.6fF
C378 diff_5294_5122# gnd! 359.6fF
C379 diff_5357_5311# gnd! 184.7fF
C380 diff_5861_5353# gnd! 1699.6fF
C381 diff_5813_5371# gnd! 187.1fF
C382 diff_5294_5263# gnd! 363.9fF
C383 diff_6043_4888# gnd! 2212.8fF
C384 diff_5357_5395# gnd! 178.1fF
C385 diff_5129_5047# gnd! 166.7fF
C386 diff_5012_5038# gnd! 185.6fF
C387 diff_5104_5113# gnd! 364.8fF
C388 diff_4784_4690# gnd! 175.4fF
C389 diff_4667_4681# gnd! 190.7fF
C390 diff_4759_4759# gnd! 370.3fF
C391 diff_4439_4336# gnd! 170.3fF
C392 diff_4325_4327# gnd! 159.5fF
C393 diff_4414_4408# gnd! 376.9fF
C394 diff_3752_3880# gnd! 166.1fF
C395 diff_3727_3844# gnd! 391.3fF
C396 diff_3635_3892# gnd! 182.3fF
C397 diff_3575_3844# gnd! 371.0fF
C398 diff_3917_4054# gnd! 371.0fF
C399 diff_4094_4231# gnd! 168.8fF
C400 diff_4072_4195# gnd! 359.5fF
C401 diff_3980_4246# gnd! 167.9fF
C402 diff_3917_4195# gnd! 379.4fF
C403 diff_4094_4336# gnd! 177.8fF
C404 diff_4262_4411# gnd! 365.6fF
C405 diff_3980_4327# gnd! 170.3fF
C406 diff_4072_4402# gnd! 367.0fF
C407 diff_4439_4585# gnd! 173.6fF
C408 diff_4414_4558# gnd! 372.5fF
C409 diff_4262_4549# gnd! 366.1fF
C410 diff_4325_4600# gnd! 173.6fF
C411 diff_4607_4765# gnd! 361.0fF
C412 diff_4784_4942# gnd! 167.9fF
C413 diff_4759_4906# gnd! 362.6fF
C414 diff_4607_4906# gnd! 357.7fF
C415 diff_4667_4957# gnd! 185.0fF
C416 diff_4949_5122# gnd! 361.4fF
C417 diff_5129_5299# gnd! 166.7fF
C418 diff_5012_5311# gnd! 183.8fF
C419 diff_5104_5260# gnd! 369.8fF
C420 diff_4949_5263# gnd! 368.8fF
C421 diff_5294_5476# gnd! 357.1fF
C422 diff_5294_5614# gnd! 362.5fF
C423 diff_5357_5665# gnd! 178.1fF
C424 diff_5357_5746# gnd! 185.6fF
C425 diff_5129_5401# gnd! 161.6fF
C426 diff_5012_5395# gnd! 180.5fF
C427 diff_5104_5470# gnd! 371.8fF
C428 diff_4784_5047# gnd! 168.5fF
C429 diff_4667_5038# gnd! 185.6fF
C430 diff_4759_5113# gnd! 373.3fF
C431 diff_4439_4690# gnd! 176.3fF
C432 diff_4325_4681# gnd! 175.4fF
C433 diff_4414_4762# gnd! 358.3fF
C434 diff_3752_3982# gnd! 167.6fF
C435 diff_3635_3973# gnd! 185.6fF
C436 diff_3727_4051# gnd! 380.4fF
C437 diff_3407_3880# gnd! 166.7fF
C438 diff_3385_3844# gnd! 379.0fF
C439 diff_3230_3844# gnd! 381.5fF
C440 diff_3293_3892# gnd! 169.4fF
C441 diff_3575_4054# gnd! 367.8fF
C442 diff_3752_4231# gnd! 167.0fF
C443 diff_3727_4195# gnd! 376.4fF
C444 diff_3575_4195# gnd! 360.2fF
C445 diff_3635_4246# gnd! 185.0fF
C446 diff_3917_4411# gnd! 387.2fF
C447 diff_4094_4585# gnd! 188.0fF
C448 diff_4072_4549# gnd! 366.2fF
C449 diff_3917_4549# gnd! 382.1fF
C450 diff_3980_4600# gnd! 172.7fF
C451 diff_4262_4765# gnd! 365.8fF
C452 diff_4439_4942# gnd! 169.4fF
C453 diff_4417_4903# gnd! 363.6fF
C454 diff_4262_4906# gnd! 349.8fF
C455 diff_4325_4954# gnd! 170.3fF
C456 diff_4607_5119# gnd! 364.2fF
C457 diff_4784_5299# gnd! 168.5fF
C458 diff_4759_5260# gnd! 369.7fF
C459 diff_4607_5263# gnd! 364.2fF
C460 diff_4667_5311# gnd! 184.7fF
C461 diff_4949_5476# gnd! 361.7fF
C462 diff_5129_5650# gnd! 166.1fF
C463 diff_5104_5617# gnd! 373.1fF
C464 diff_5012_5665# gnd! 184.1fF
C465 diff_4949_5614# gnd! 367.3fF
C466 diff_5294_5827# gnd! 358.2fF
C467 diff_5294_5968# gnd! 358.4fF
C468 diff_5357_6019# gnd! 183.8fF
C469 o2 gnd! 5968.9fF
C470 diff_5938_6088# gnd! 1230.8fF
C471 diff_5357_6100# gnd! 184.7fF
C472 diff_6137_6238# gnd! 422.9fF
C473 diff_6059_6298# gnd! 414.1fF
C474 diff_5129_5755# gnd! 166.7fF
C475 diff_5012_5746# gnd! 185.6fF
C476 diff_5104_5824# gnd! 368.2fF
C477 diff_4784_5401# gnd! 166.7fF
C478 diff_4667_5392# gnd! 182.9fF
C479 diff_4759_5470# gnd! 366.4fF
C480 diff_4325_5038# gnd! 158.6fF
C481 diff_4439_5047# gnd! 170.3fF
C482 diff_4417_5113# gnd! 369.2fF
C483 diff_4094_4690# gnd! 191.9fF
C484 diff_3980_4681# gnd! 176.3fF
C485 diff_4072_4759# gnd! 357.8fF
C486 diff_3752_4336# gnd! 167.6fF
C487 diff_3635_4327# gnd! 185.0fF
C488 diff_3727_4405# gnd! 382.5fF
C489 diff_3407_3982# gnd! 167.6fF
C490 diff_3293_3973# gnd! 169.4fF
C491 diff_3385_4051# gnd! 375.7fF
C492 diff_3065_3877# gnd! 170.9fF
C493 diff_3040_3844# gnd! 386.6fF
C494 diff_2951_3892# gnd! 173.6fF
C495 diff_2888_3841# gnd! 373.7fF
C496 diff_3230_4054# gnd! 375.3fF
C497 diff_3407_4231# gnd! 169.7fF
C498 diff_3385_4195# gnd! 369.8fF
C499 diff_3230_4195# gnd! 364.6fF
C500 diff_3293_4246# gnd! 170.6fF
C501 diff_3575_4411# gnd! 365.5fF
C502 diff_3407_4336# gnd! 168.5fF
C503 diff_3293_4327# gnd! 171.2fF
C504 diff_3385_4402# gnd! 373.7fF
C505 diff_3752_4588# gnd! 167.6fF
C506 diff_3727_4549# gnd! 377.4fF
C507 diff_3575_4552# gnd! 371.7fF
C508 diff_3635_4600# gnd! 185.6fF
C509 diff_3917_4762# gnd! 380.1fF
C510 diff_4094_4942# gnd! 182.6fF
C511 diff_4072_4906# gnd! 351.1fF
C512 diff_3980_4957# gnd! 167.9fF
C513 diff_3917_4906# gnd! 375.7fF
C514 diff_4262_5119# gnd! 358.8fF
C515 diff_4439_5296# gnd! 172.7fF
C516 diff_4414_5275# gnd! 364.6fF
C517 diff_4262_5260# gnd! 357.7fF
C518 diff_4325_5311# gnd! 174.5fF
C519 diff_4607_5473# gnd! 360.0fF
C520 diff_4784_5650# gnd! 170.6fF
C521 diff_4759_5617# gnd! 374.9fF
C522 diff_4604_5627# gnd! 368.9fF
C523 diff_4667_5665# gnd! 183.2fF
C524 diff_4949_5827# gnd! 362.0fF
C525 diff_5129_6007# gnd! 160.1fF
C526 diff_5104_5968# gnd! 370.5fF
C527 diff_4949_5968# gnd! 363.3fF
C528 diff_5012_6019# gnd! 178.1fF
C529 diff_5294_6181# gnd! 354.9fF
C530 diff_5294_6322# gnd! 359.8fF
C531 diff_5357_6373# gnd! 149.6fF
C532 diff_5861_6427# gnd! 1682.4fF
C533 diff_5813_6445# gnd! 189.8fF
C534 diff_6035_6505# gnd! 2174.2fF
C535 diff_5563_3961# gnd! 4525.4fF
C536 diff_5357_6454# gnd! 190.7fF
C537 diff_5126_6140# gnd! 170.9fF
C538 diff_5012_6100# gnd! 184.7fF
C539 diff_5104_6178# gnd! 356.4fF
C540 diff_4784_5755# gnd! 168.5fF
C541 diff_4667_5746# gnd! 186.5fF
C542 diff_4759_5824# gnd! 368.8fF
C543 diff_4439_5401# gnd! 169.4fF
C544 diff_4322_5396# gnd! 173.3fF
C545 diff_4414_5473# gnd! 364.3fF
C546 diff_4094_5047# gnd! 186.5fF
C547 diff_3980_5038# gnd! 170.3fF
C548 diff_4072_5113# gnd! 360.9fF
C549 diff_3752_4690# gnd! 173.6fF
C550 diff_3635_4681# gnd! 192.5fF
C551 diff_3727_4759# gnd! 375.9fF
C552 diff_3065_3982# gnd! 168.5fF
C553 diff_2951_3973# gnd! 168.5fF
C554 diff_3040_4051# gnd! 382.1fF
C555 diff_2720_3877# gnd! 180.5fF
C556 diff_2606_3892# gnd! 174.5fF
C557 diff_2698_3844# gnd! 382.1fF
C558 diff_2546_3841# gnd! 385.5fF
C559 diff_2888_4054# gnd! 370.8fF
C560 diff_2720_3982# gnd! 168.5fF
C561 diff_2606_3973# gnd! 169.4fF
C562 diff_2698_4051# gnd! 376.9fF
C563 diff_3065_4231# gnd! 172.1fF
C564 diff_3040_4195# gnd! 375.1fF
C565 diff_2888_4195# gnd! 364.2fF
C566 diff_2951_4243# gnd! 171.2fF
C567 diff_3230_4411# gnd! 364.4fF
C568 diff_3407_4588# gnd! 169.4fF
C569 diff_3385_4549# gnd! 373.9fF
C570 diff_3230_4552# gnd! 375.3fF
C571 diff_3293_4600# gnd! 170.3fF
C572 diff_3575_4762# gnd! 364.9fF
C573 diff_3407_4690# gnd! 176.3fF
C574 diff_3293_4681# gnd! 161.9fF
C575 diff_3385_4759# gnd! 369.8fF
C576 diff_3752_4942# gnd! 167.9fF
C577 diff_3727_4906# gnd! 372.5fF
C578 diff_3635_4954# gnd! 185.6fF
C579 diff_3575_4906# gnd! 373.3fF
C580 diff_3917_5119# gnd! 375.4fF
C581 diff_4094_5299# gnd! 178.4fF
C582 diff_4072_5260# gnd! 362.1fF
C583 diff_3917_5263# gnd! 378.1fF
C584 diff_3980_5311# gnd! 170.3fF
C585 diff_3980_5392# gnd! 168.5fF
C586 diff_4094_5401# gnd! 169.4fF
C587 diff_4262_5473# gnd! 355.0fF
C588 diff_4072_5470# gnd! 357.8fF
C589 diff_4439_5650# gnd! 168.8fF
C590 diff_4414_5617# gnd! 367.2fF
C591 diff_4262_5614# gnd! 369.8fF
C592 diff_4322_5665# gnd! 179.9fF
C593 diff_4604_5834# gnd! 358.2fF
C594 diff_4784_6004# gnd! 169.1fF
C595 diff_4759_5968# gnd! 365.4fF
C596 diff_4604_5972# gnd! 361.9fF
C597 diff_4667_6019# gnd! 182.3fF
C598 diff_4949_6181# gnd! 359.8fF
C599 diff_5129_6358# gnd! 170.6fF
C600 diff_5104_6322# gnd! 369.8fF
C601 diff_4949_6322# gnd! 361.4fF
C602 diff_5012_6373# gnd! 184.1fF
C603 diff_5335_3644# gnd! 2745.0fF
C604 diff_5278_3644# gnd! 2538.4fF
C605 diff_5206_3742# gnd! 2556.7fF
C606 diff_5129_6463# gnd! 166.7fF
C607 diff_5012_6454# gnd! 184.7fF
C608 diff_5116_3613# gnd! 2745.0fF
C609 diff_5294_6538# gnd! 349.5fF
C610 diff_5104_6532# gnd! 355.1fF
C611 diff_4732_1658# gnd! 7521.2fF
C612 diff_4987_3652# gnd! 2752.2fF
C613 diff_4784_6109# gnd! 168.5fF
C614 diff_4667_6100# gnd! 186.5fF
C615 diff_4759_6178# gnd! 361.1fF
C616 diff_4439_5755# gnd! 170.3fF
C617 diff_4322_5746# gnd! 184.1fF
C618 diff_4414_5824# gnd! 362.1fF
C619 diff_3752_5047# gnd! 167.6fF
C620 diff_3635_5038# gnd! 184.7fF
C621 diff_3727_5113# gnd! 379.1fF
C622 diff_2951_4327# gnd! 169.4fF
C623 diff_3065_4336# gnd! 170.3fF
C624 diff_3040_4405# gnd! 378.7fF
C625 diff_2378_3877# gnd! 173.6fF
C626 diff_2264_3889# gnd! 176.0fF
C627 diff_2353_3844# gnd! 381.8fF
C628 diff_2201_3841# gnd! 369.3fF
C629 diff_2546_4054# gnd! 380.1fF
C630 diff_2720_4231# gnd! 176.0fF
C631 diff_2698_4195# gnd! 367.3fF
C632 diff_2543_4195# gnd! 376.2fF
C633 diff_2606_4243# gnd! 176.0fF
C634 diff_2888_4411# gnd! 368.3fF
C635 diff_2720_4336# gnd! 173.3fF
C636 diff_2606_4327# gnd! 171.2fF
C637 diff_2698_4405# gnd! 376.7fF
C638 diff_3065_4588# gnd! 167.6fF
C639 diff_2888_4552# gnd! 369.7fF
C640 diff_2951_4597# gnd! 170.0fF
C641 diff_3040_4549# gnd! 378.8fF
C642 diff_3230_4762# gnd! 383.1fF
C643 diff_3065_4690# gnd! 172.7fF
C644 diff_2951_4681# gnd! 175.4fF
C645 diff_3040_4759# gnd! 381.6fF
C646 diff_3407_4942# gnd! 172.1fF
C647 diff_3385_4906# gnd! 374.3fF
C648 diff_3230_4906# gnd! 375.1fF
C649 diff_3293_4954# gnd! 171.2fF
C650 diff_3575_5122# gnd! 365.6fF
C651 diff_3407_5047# gnd! 168.5fF
C652 diff_3293_5038# gnd! 171.2fF
C653 diff_3385_5113# gnd! 370.6fF
C654 diff_3752_5299# gnd! 167.6fF
C655 diff_3727_5260# gnd! 378.6fF
C656 diff_3635_5311# gnd! 183.8fF
C657 diff_3575_5263# gnd! 369.1fF
C658 diff_3917_5473# gnd! 375.2fF
C659 diff_4094_5650# gnd! 170.3fF
C660 diff_4072_5614# gnd! 362.8fF
C661 diff_3917_5614# gnd! 373.3fF
C662 diff_3980_5665# gnd! 168.8fF
C663 diff_4262_5827# gnd! 349.5fF
C664 diff_4439_6004# gnd! 171.2fF
C665 diff_4414_5971# gnd! 371.1fF
C666 diff_4262_5968# gnd! 361.7fF
C667 diff_4322_6019# gnd! 184.1fF
C668 diff_4604_6181# gnd! 354.6fF
C669 diff_4784_6358# gnd! 171.5fF
C670 diff_4759_6325# gnd! 363.3fF
C671 diff_4607_6322# gnd! 359.4fF
C672 diff_4667_6373# gnd! 187.7fF
C673 diff_4933_3644# gnd! 2560.4fF
C674 diff_4861_3742# gnd! 2542.4fF
C675 diff_4784_6463# gnd! 170.3fF
C676 diff_4667_6454# gnd! 185.6fF
C677 diff_4949_6538# gnd! 356.9fF
C678 diff_4759_6532# gnd! 358.5fF
C679 diff_4771_3607# gnd! 2734.7fF
C680 diff_4439_6109# gnd! 169.4fF
C681 diff_4322_6100# gnd! 185.6fF
C682 diff_4414_6178# gnd! 364.0fF
C683 diff_4094_5755# gnd! 169.4fF
C684 diff_3980_5746# gnd! 168.5fF
C685 diff_4072_5821# gnd! 353.3fF
C686 diff_3635_5392# gnd! 184.7fF
C687 diff_3752_5401# gnd! 168.5fF
C688 diff_3727_5470# gnd! 367.8fF
C689 diff_2378_3982# gnd! 168.5fF
C690 diff_2264_3973# gnd! 170.3fF
C691 diff_2353_4051# gnd! 379.7fF
C692 diff_1217_3803# gnd! 766.0fF
C693 diff_1267_3856# gnd! 1360.6fF
C694 diff_1663_3859# gnd! 7709.1fF
C695 diff_2036_3880# gnd! 168.5fF
C696 diff_2011_3844# gnd! 387.3fF
C697 diff_2201_4054# gnd! 368.2fF
C698 diff_2378_4231# gnd! 175.1fF
C699 diff_2353_4195# gnd! 368.4fF
C700 diff_2201_4195# gnd! 359.3fF
C701 diff_2264_4243# gnd! 173.6fF
C702 diff_2543_4411# gnd! 386.7fF
C703 diff_2720_4588# gnd! 169.4fF
C704 diff_2698_4549# gnd! 371.4fF
C705 diff_2543_4552# gnd! 373.2fF
C706 diff_2606_4600# gnd! 170.3fF
C707 diff_2888_4765# gnd! 360.0fF
C708 diff_2720_4690# gnd! 177.5fF
C709 diff_2606_4681# gnd! 176.3fF
C710 diff_2698_4759# gnd! 367.2fF
C711 diff_3065_4942# gnd! 169.4fF
C712 diff_3040_4906# gnd! 375.2fF
C713 diff_2951_4954# gnd! 169.4fF
C714 diff_2888_4906# gnd! 367.4fF
C715 diff_3230_5122# gnd! 369.9fF
C716 diff_3407_5299# gnd! 168.5fF
C717 diff_3385_5260# gnd! 369.5fF
C718 diff_3230_5263# gnd! 366.9fF
C719 diff_3293_5311# gnd! 169.4fF
C720 diff_3575_5473# gnd! 360.4fF
C721 diff_3407_5401# gnd! 167.6fF
C722 diff_3293_5392# gnd! 169.4fF
C723 diff_3385_5470# gnd! 362.2fF
C724 diff_3752_5650# gnd! 167.0fF
C725 diff_3727_5617# gnd! 370.6fF
C726 diff_3635_5665# gnd! 185.0fF
C727 diff_3575_5614# gnd! 362.9fF
C728 diff_3917_5827# gnd! 364.1fF
C729 diff_4094_6004# gnd! 168.8fF
C730 diff_4072_5968# gnd! 357.7fF
C731 diff_3917_5968# gnd! 363.9fF
C732 diff_3980_6019# gnd! 171.5fF
C733 diff_4262_6181# gnd! 353.1fF
C734 diff_4439_6358# gnd! 170.3fF
C735 diff_4414_6325# gnd! 365.6fF
C736 diff_4262_6322# gnd! 358.0fF
C737 diff_4322_6370# gnd! 187.1fF
C738 diff_4642_3644# gnd! 2746.6fF
C739 diff_4588_3644# gnd! 2782.6fF
C740 diff_4516_3742# gnd! 2531.3fF
C741 diff_4426_3610# gnd! 2737.9fF
C742 diff_4439_6463# gnd! 170.3fF
C743 diff_4604_6554# gnd! 352.1fF
C744 diff_4414_6532# gnd! 358.8fF
C745 diff_4322_6470# gnd! 180.8fF
C746 diff_4094_6109# gnd! 169.4fF
C747 diff_3980_6100# gnd! 169.4fF
C748 diff_4072_6178# gnd! 353.9fF
C749 diff_3752_5755# gnd! 169.4fF
C750 diff_3635_5746# gnd! 183.8fF
C751 diff_3727_5824# gnd! 372.5fF
C752 diff_2951_5038# gnd! 168.5fF
C753 diff_3065_5047# gnd! 169.4fF
C754 diff_3040_5113# gnd! 378.4fF
C755 diff_2378_4336# gnd! 174.5fF
C756 diff_2264_4327# gnd! 170.9fF
C757 diff_2353_4405# gnd! 378.9fF
C758 diff_2033_3992# gnd! 171.2fF
C759 diff_1370_3857# gnd! 6166.2fF
C760 diff_1421_3899# gnd! 1072.5fF
C761 diff_2011_4051# gnd! 383.1fF
C762 diff_1663_4051# gnd! 7739.0fF
C763 diff_1421_4000# gnd! 1042.7fF
C764 diff_1370_4027# gnd! 6185.8fF
C765 diff_1102_3989# gnd! 396.8fF
C766 diff_1267_4048# gnd! 1331.7fF
C767 diff_1217_4105# gnd! 780.5fF
C768 diff_406_3802# gnd! 659.4fF
C769 diff_406_4054# gnd! 647.4fF
C770 diff_1267_4210# gnd! 1315.9fF
C771 diff_1663_4210# gnd! 7631.8fF
C772 diff_2033_4231# gnd! 190.1fF
C773 diff_2011_4195# gnd! 367.2fF
C774 diff_2201_4411# gnd! 369.0fF
C775 diff_2378_4588# gnd! 169.4fF
C776 diff_2353_4549# gnd! 375.2fF
C777 diff_2201_4552# gnd! 367.5fF
C778 diff_2264_4600# gnd! 169.4fF
C779 diff_2543_4765# gnd! 368.6fF
C780 diff_2720_4942# gnd! 176.0fF
C781 diff_2698_4903# gnd! 377.9fF
C782 diff_2543_4906# gnd! 379.0fF
C783 diff_2606_4954# gnd! 175.1fF
C784 diff_2888_5122# gnd! 360.7fF
C785 diff_2720_5047# gnd! 168.5fF
C786 diff_2606_5038# gnd! 171.2fF
C787 diff_2698_5113# gnd! 370.5fF
C788 diff_3065_5299# gnd! 167.6fF
C789 diff_3040_5260# gnd! 374.9fF
C790 diff_2888_5263# gnd! 363.6fF
C791 diff_2951_5311# gnd! 169.4fF
C792 diff_3230_5473# gnd! 364.0fF
C793 diff_3407_5650# gnd! 169.7fF
C794 diff_3385_5614# gnd! 372.8fF
C795 diff_3293_5665# gnd! 169.7fF
C796 diff_3230_5614# gnd! 367.4fF
C797 diff_3575_5827# gnd! 360.2fF
C798 diff_3749_6050# gnd! 168.2fF
C799 diff_3727_5968# gnd! 367.4fF
C800 diff_3635_6019# gnd! 184.1fF
C801 diff_3575_5968# gnd! 358.7fF
C802 diff_3917_6181# gnd! 355.1fF
C803 diff_4094_6358# gnd! 170.3fF
C804 diff_4072_6322# gnd! 355.5fF
C805 diff_3917_6322# gnd! 365.6fF
C806 diff_3980_6370# gnd! 168.5fF
C807 diff_4300_3644# gnd! 2974.0fF
C808 diff_4243_3644# gnd! 2532.9fF
C809 diff_4171_3745# gnd! 2533.8fF
C810 diff_4094_6463# gnd! 169.4fF
C811 diff_3980_6454# gnd! 168.5fF
C812 diff_4084_3607# gnd! 2799.8fF
C813 diff_4262_6535# gnd! 350.6fF
C814 diff_4072_6529# gnd! 353.7fF
C815 diff_3955_3644# gnd! 2727.4fF
C816 diff_3752_6109# gnd! 168.5fF
C817 diff_3635_6100# gnd! 184.7fF
C818 diff_3727_6178# gnd! 359.8fF
C819 diff_3407_5755# gnd! 167.6fF
C820 diff_3293_5746# gnd! 170.3fF
C821 diff_3385_5821# gnd! 366.3fF
C822 diff_2951_5392# gnd! 170.3fF
C823 diff_3065_5401# gnd! 168.5fF
C824 diff_3040_5470# gnd! 372.4fF
C825 diff_2378_4690# gnd! 172.7fF
C826 diff_2264_4681# gnd! 177.8fF
C827 diff_2353_4759# gnd! 372.2fF
C828 diff_2033_4336# gnd! 191.6fF
C829 diff_2011_4402# gnd! 377.0fF
C830 diff_1370_4211# gnd! 6089.9fF
C831 diff_1421_4253# gnd! 1028.7fF
C832 diff_1060_3926# gnd! 1596.2fF
C833 diff_1217_4228# gnd! 876.1fF
C834 diff_1663_4402# gnd! 7889.8fF
C835 diff_1421_4354# gnd! 1037.5fF
C836 diff_1370_4381# gnd! 6090.7fF
C837 diff_1093_4033# gnd! 2384.5fF
C838 diff_223_4213# gnd! 1377.5fF
C839 diff_1267_4369# gnd! 1365.8fF
C840 diff_1217_4351# gnd! 898.7fF
C841 diff_1217_4504# gnd! 814.9fF
C842 diff_1267_4564# gnd! 1338.3fF
C843 diff_2033_4588# gnd! 184.7fF
C844 diff_2011_4549# gnd! 374.7fF
C845 diff_1663_4564# gnd! 7788.6fF
C846 diff_1370_4565# gnd! 6072.2fF
C847 diff_1421_4607# gnd! 1095.3fF
C848 diff_2201_4765# gnd! 361.5fF
C849 diff_2353_4906# gnd! 377.6fF
C850 diff_2378_4942# gnd! 174.5fF
C851 diff_2201_4906# gnd! 365.8fF
C852 diff_2264_4954# gnd! 175.4fF
C853 diff_2543_5122# gnd! 370.2fF
C854 diff_2720_5299# gnd! 168.5fF
C855 diff_2698_5260# gnd! 369.4fF
C856 diff_2543_5263# gnd! 374.0fF
C857 diff_2606_5311# gnd! 168.5fF
C858 diff_2888_5473# gnd! 352.8fF
C859 diff_3065_5650# gnd! 167.9fF
C860 diff_3040_5617# gnd! 375.2fF
C861 diff_2888_5614# gnd! 367.7fF
C862 diff_2948_5669# gnd! 185.6fF
C863 diff_3230_5827# gnd! 361.2fF
C864 diff_3407_6004# gnd! 171.2fF
C865 diff_3385_5968# gnd! 364.9fF
C866 diff_3230_5968# gnd! 362.3fF
C867 diff_3293_6019# gnd! 173.9fF
C868 diff_3575_6181# gnd! 357.7fF
C869 diff_3752_6358# gnd! 168.5fF
C870 diff_3635_6370# gnd! 185.6fF
C871 diff_3575_6322# gnd! 360.0fF
C872 diff_3727_6322# gnd! 364.2fF
C873 diff_3898_3644# gnd! 2542.8fF
C874 diff_3829_3644# gnd! 2685.2fF
C875 diff_3739_3610# gnd! 2729.0fF
C876 diff_3752_6463# gnd! 168.5fF
C877 diff_3635_6454# gnd! 186.5fF
C878 diff_3917_6535# gnd! 363.0fF
C879 diff_3727_6532# gnd! 364.8fF
C880 diff_3407_6109# gnd! 168.5fF
C881 diff_3293_6100# gnd! 169.4fF
C882 diff_3385_6175# gnd! 365.2fF
C883 diff_3065_5755# gnd! 168.5fF
C884 diff_2948_5746# gnd! 188.6fF
C885 diff_3040_5824# gnd! 372.7fF
C886 diff_2720_5401# gnd! 167.6fF
C887 diff_2606_5392# gnd! 169.4fF
C888 diff_2698_5470# gnd! 377.6fF
C889 diff_2378_5047# gnd! 170.3fF
C890 diff_2264_5038# gnd! 171.2fF
C891 diff_2353_5113# gnd! 368.9fF
C892 diff_2033_4693# gnd! 185.9fF
C893 diff_2011_4759# gnd! 366.1fF
C894 diff_1663_4756# gnd! 7716.3fF
C895 diff_1421_4708# gnd! 1106.1fF
C896 diff_1370_4735# gnd! 6372.6fF
C897 diff_1102_4697# gnd! 390.5fF
C898 diff_1267_4756# gnd! 1327.8fF
C899 diff_1217_4813# gnd! 822.8fF
C900 diff_175_4780# gnd! 5106.0fF
C901 d3 gnd! 18244.3fF
C902 diff_172_3988# gnd! 4758.6fF
C903 diff_1267_4921# gnd! 1308.2fF
C904 diff_1663_4918# gnd! 7602.5fF
C905 diff_2033_4942# gnd! 191.6fF
C906 diff_2011_4906# gnd! 369.1fF
C907 diff_1370_4919# gnd! 6147.9fF
C908 diff_1421_4961# gnd! 1039.1fF
C909 diff_2201_5119# gnd! 361.8fF
C910 diff_2378_5299# gnd! 169.4fF
C911 diff_2353_5260# gnd! 382.0fF
C912 diff_2201_5263# gnd! 363.3fF
C913 diff_2261_5345# gnd! 177.2fF
C914 diff_2543_5473# gnd! 375.2fF
C915 diff_2720_5650# gnd! 174.5fF
C916 diff_2698_5614# gnd! 378.3fF
C917 diff_2543_5614# gnd! 380.8fF
C918 diff_2606_5662# gnd! 173.0fF
C919 diff_2888_5827# gnd! 362.1fF
C920 diff_2720_5755# gnd! 171.2fF
C921 diff_2606_5746# gnd! 171.2fF
C922 diff_2698_5821# gnd! 368.5fF
C923 diff_3065_6004# gnd! 171.2fF
C924 diff_3040_5968# gnd! 370.1fF
C925 diff_2948_6019# gnd! 187.7fF
C926 diff_2888_5968# gnd! 359.7fF
C927 diff_3230_6181# gnd! 361.2fF
C928 diff_3407_6358# gnd! 168.5fF
C929 diff_3385_6322# gnd! 363.9fF
C930 diff_3230_6322# gnd! 359.7fF
C931 diff_3293_6370# gnd! 170.3fF
C932 diff_3610_3644# gnd! 2752.6fF
C933 diff_3575_6535# gnd! 360.3fF
C934 diff_3556_3644# gnd! 2697.3fF
C935 diff_3484_3742# gnd! 2533.9fF
C936 diff_3407_6463# gnd! 168.5fF
C937 diff_3293_6454# gnd! 171.2fF
C938 diff_3385_6529# gnd! 363.0fF
C939 diff_3394_3613# gnd! 2958.7fF
C940 diff_3065_6109# gnd! 168.5fF
C941 diff_2948_6100# gnd! 185.6fF
C942 diff_3040_6178# gnd! 363.4fF
C943 diff_2378_5401# gnd! 168.5fF
C944 diff_2261_5392# gnd! 175.1fF
C945 diff_2353_5470# gnd! 379.5fF
C946 diff_2033_5047# gnd! 188.6fF
C947 diff_2011_5113# gnd! 371.9fF
C948 diff_1217_4939# gnd! 870.4fF
C949 diff_1060_4634# gnd! 1586.6fF
C950 diff_1663_5113# gnd! 7780.5fF
C951 diff_1421_5065# gnd! 1049.6fF
C952 diff_1370_5092# gnd! 6076.5fF
C953 diff_1267_5095# gnd! 1337.0fF
C954 diff_829_3778# gnd! 3618.1fF
C955 diff_1217_5074# gnd! 867.1fF
C956 diff_1217_5215# gnd! 805.0fF
C957 diff_1267_5275# gnd! 1336.6fF
C958 diff_1663_5275# gnd! 7991.1fF
C959 diff_2033_5299# gnd! 184.7fF
C960 diff_2011_5260# gnd! 373.4fF
C961 diff_2033_5401# gnd! 184.7fF
C962 diff_1370_5273# gnd! 6057.8fF
C963 diff_1421_5318# gnd! 1055.5fF
C964 diff_2201_5473# gnd! 361.3fF
C965 diff_2378_5650# gnd! 172.7fF
C966 diff_2353_5617# gnd! 382.1fF
C967 diff_2201_5614# gnd! 366.0fF
C968 diff_2261_5665# gnd! 186.8fF
C969 diff_2543_5827# gnd! 362.8fF
C970 diff_2543_5968# gnd! 359.9fF
C971 diff_2720_6004# gnd! 175.1fF
C972 diff_2698_5968# gnd! 366.8fF
C973 diff_2606_6019# gnd! 175.7fF
C974 diff_2888_6181# gnd! 353.2fF
C975 diff_2888_6322# gnd! 356.0fF
C976 diff_2948_6370# gnd! 187.4fF
C977 diff_3065_6358# gnd! 170.3fF
C978 diff_3040_6322# gnd! 365.4fF
C979 diff_3268_3644# gnd! 2729.0fF
C980 diff_3211_3644# gnd! 2542.7fF
C981 diff_3142_3644# gnd! 2769.9fF
C982 diff_3052_3607# gnd! 2726.1fF
C983 diff_2948_6454# gnd! 187.4fF
C984 diff_3065_6463# gnd! 170.3fF
C985 diff_3230_6535# gnd! 353.1fF
C986 diff_3040_6529# gnd! 367.9fF
C987 diff_2923_3644# gnd! 3013.1fF
C988 diff_2720_6109# gnd! 168.5fF
C989 diff_2606_6100# gnd! 170.3fF
C990 diff_2698_6175# gnd! 366.3fF
C991 diff_2378_5755# gnd! 169.4fF
C992 diff_2261_5746# gnd! 187.4fF
C993 diff_2353_5824# gnd! 373.8fF
C994 diff_2011_5470# gnd! 364.5fF
C995 diff_1663_5467# gnd! 7866.9fF
C996 diff_425_5110# gnd! 1378.1fF
C997 diff_407_5030# gnd! 1351.8fF
C998 diff_1421_5419# gnd! 1095.8fF
C999 diff_1370_5446# gnd! 6070.3fF
C1000 diff_1102_5408# gnd! 380.0fF
C1001 diff_1267_5467# gnd! 1336.5fF
C1002 diff_1217_5524# gnd! 800.2fF
C1003 diff_1267_5629# gnd! 1313.2fF
C1004 diff_1663_5629# gnd! 7725.0fF
C1005 diff_2033_5650# gnd! 173.6fF
C1006 diff_2011_5614# gnd! 368.6fF
C1007 diff_2033_5755# gnd! 167.6fF
C1008 diff_2201_5827# gnd! 362.7fF
C1009 diff_2011_5821# gnd! 368.1fF
C1010 diff_2375_6020# gnd! 185.3fF
C1011 diff_2353_5968# gnd! 371.6fF
C1012 diff_2201_5968# gnd! 363.6fF
C1013 diff_2261_6019# gnd! 191.0fF
C1014 diff_2543_6181# gnd! 360.2fF
C1015 diff_2720_6358# gnd! 170.3fF
C1016 diff_2695_6331# gnd! 366.9fF
C1017 diff_2543_6322# gnd! 362.9fF
C1018 diff_2606_6370# gnd! 171.2fF
C1019 diff_2720_6463# gnd! 170.3fF
C1020 diff_2869_3644# gnd! 2626.2fF
C1021 diff_2797_3745# gnd! 2547.7fF
C1022 diff_2707_3610# gnd! 3123.2fF
C1023 diff_2888_6535# gnd! 356.8fF
C1024 diff_2698_6529# gnd! 364.2fF
C1025 diff_2606_6454# gnd! 171.2fF
C1026 diff_2375_6109# gnd! 184.4fF
C1027 diff_2261_6100# gnd! 186.5fF
C1028 diff_2353_6178# gnd! 355.0fF
C1029 diff_1370_5630# gnd! 6043.9fF
C1030 diff_1418_5684# gnd! 1051.6fF
C1031 diff_1217_5647# gnd! 870.5fF
C1032 diff_1060_5345# gnd! 1551.8fF
C1033 diff_1663_5821# gnd! 7935.3fF
C1034 diff_1418_5773# gnd! 1041.7fF
C1035 diff_1370_5800# gnd! 6024.6fF
C1036 diff_1267_5803# gnd! 1331.8fF
C1037 diff_406_5716# gnd! 655.5fF
C1038 diff_820_3511# gnd! 4146.3fF
C1039 diff_1217_5782# gnd! 880.6fF
C1040 diff_1217_5923# gnd! 790.1fF
C1041 diff_580_3394# gnd! 20543.1fF
C1042 diff_1267_5983# gnd! 1343.6fF
C1043 diff_1663_5983# gnd! 7725.8fF
C1044 diff_2033_6004# gnd! 175.1fF
C1045 diff_2011_5968# gnd! 370.8fF
C1046 diff_2201_6181# gnd! 357.5fF
C1047 diff_2033_6109# gnd! 166.7fF
C1048 diff_1370_5981# gnd! 6035.6fF
C1049 diff_1418_6026# gnd! 1076.8fF
C1050 diff_2011_6175# gnd! 356.9fF
C1051 diff_2377_6413# gnd! 174.1fF
C1052 diff_2353_6322# gnd! 378.4fF
C1053 diff_2261_6370# gnd! 189.8fF
C1054 diff_2201_6322# gnd! 353.8fF
C1055 diff_2581_3644# gnd! 2724.6fF
C1056 diff_2524_3644# gnd! 2584.1fF
C1057 diff_2455_3644# gnd! 2717.3fF
C1058 diff_2365_3607# gnd! 2733.4fF
C1059 diff_2378_6463# gnd! 170.3fF
C1060 diff_2261_6454# gnd! 187.4fF
C1061 diff_2543_6535# gnd! 357.6fF
C1062 diff_2353_6529# gnd! 374.0fF
C1063 diff_2236_3644# gnd! 2940.1fF
C1064 diff_406_5971# gnd! 643.1fF
C1065 diff_1660_6178# gnd! 8034.6fF
C1066 diff_1418_6127# gnd! 1076.6fF
C1067 diff_1370_6154# gnd! 6018.0fF
C1068 diff_1102_6116# gnd! 410.3fF
C1069 diff_1267_6169# gnd! 1359.4fF
C1070 diff_1217_6229# gnd! 795.9fF
C1071 diff_220_6232# gnd! 1352.2fF
C1072 diff_1267_6334# gnd! 1374.0fF
C1073 diff_1663_6337# gnd! 7611.2fF
C1074 diff_2033_6358# gnd! 173.0fF
C1075 diff_2011_6322# gnd! 366.6fF
C1076 diff_2033_6463# gnd! 172.1fF
C1077 diff_2182_3644# gnd! 2548.9fF
C1078 diff_2110_3745# gnd! 2759.0fF
C1079 diff_2020_3610# gnd! 2870.5fF
C1080 diff_2201_6535# gnd! 360.3fF
C1081 diff_2011_6529# gnd! 362.9fF
C1082 diff_1370_6335# gnd! 6282.2fF
C1083 diff_1418_6383# gnd! 1076.4fF
C1084 diff_1217_6388# gnd! 890.2fF
C1085 diff_577_5317# gnd! 18468.9fF
C1086 diff_1060_6050# gnd! 1549.4fF
C1087 diff_1660_6529# gnd! 7792.3fF
C1088 diff_1418_6481# gnd! 1060.5fF
C1089 diff_1066_3979# gnd! 7710.6fF
C1090 diff_1370_6508# gnd! 5867.5fF
C1091 diff_1267_6511# gnd! 1390.1fF
C1092 diff_1217_6508# gnd! 805.9fF
C1093 diff_1309_3670# gnd! 4119.1fF
C1094 diff_817_6145# gnd! 4741.6fF
C1095 diff_5813_6613# gnd! 220.7fF
C1096 diff_6059_6787# gnd! 389.1fF
C1097 diff_5864_6631# gnd! 1637.1fF
C1098 diff_6134_6844# gnd! 438.2fF
C1099 clk2 gnd! 21241.5fF
C1100 diff_5263_6937# gnd! 198.2fF
C1101 diff_175_6337# gnd! 5120.9fF
C1102 d2 gnd! 18375.1fF
C1103 diff_172_5905# gnd! 4746.8fF
C1104 o1 gnd! 6367.2fF
C1105 diff_5935_6883# gnd! 1325.5fF
C1106 diff_6040_7132# gnd! 2267.8fF
C1107 diff_5188_6931# gnd! 8706.0fF
C1108 diff_556_2707# gnd! 7483.1fF
C1109 diff_872_2743# gnd! 16628.2fF
C1110 diff_5128_7225# gnd! 360.1fF
C1111 diff_5039_7261# gnd! 376.4fF
C1112 diff_4808_7162# gnd! 1223.8fF
C1113 diff_5194_7252# gnd! 4437.2fF
C1114 o0 gnd! 6043.2fF
C1115 diff_3397_7141# gnd! 650.9fF
C1116 diff_3154_7144# gnd! 667.7fF
C1117 diff_2522_7033# gnd! 1351.2fF
C1118 diff_3574_7198# gnd! 1234.9fF
C1119 diff_2359_7109# gnd! 1423.7fF
C1120 diff_3157_7220# gnd! 5172.1fF
C1121 diff_3328_7249# gnd! 4674.4fF
C1122 diff_629_6919# gnd! 17868.3fF
C1123 diff_967_7144# gnd! 665.6fF
C1124 Vdd gnd! 227187.0fF
C1125 diff_331_7000# gnd! 10517.2fF
C1126 diff_413_7055# gnd! 1356.5fF
C1127 diff_724_7144# gnd! 681.3fF
C1128 diff_244_7114# gnd! 1445.6fF
C1129 diff_1144_7198# gnd! 1335.9fF
C1130 diff_220_5722# gnd! 11948.0fF
C1131 diff_724_7211# gnd! 5160.9fF
C1132 diff_898_7246# gnd! 4749.7fF
C1133 diff_4792_7153# gnd! 2307.5fF
C1134 d0 gnd! 17129.8fF
C1135 d1 gnd! 17052.3fF
C1136 diff_5044_7399# gnd! 1568.4fF
