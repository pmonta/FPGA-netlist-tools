* SPICE3 file created from 4003.ext - technology: nmos

.option scale=0.001u

M1000 vcc vcc diff_258130_451520# vss efet w=10790 l=9960
M1003 vcc vcc diff_1540480_996000# vss efet w=6640 l=143590
M1004 diff_1540480_996000# diff_232400_451520# vss vss efet w=14940 l=7470
M1005 vss diff_1466610_1008450# diff_258130_451520# vss efet w=247340 l=14110
M1006 vcc vcc diff_1466610_1008450# vss efet w=6640 l=146080
M1007 diff_1466610_1008450# diff_1540480_996000# vss vss efet w=174300 l=22410
M1008 vss diff_273900_560250# diff_232400_451520# vss efet w=150230 l=7470
M1009 diff_273900_560250# diff_232400_451520# vss vss efet w=61420 l=7470
M1010 q4 diff_404210_938730# vss vss efet w=351505 l=7885
M1011 vss diff_312080_771900# diff_296310_846600# vss efet w=66815 l=7885
M1012 diff_296310_846600# diff_207500_451520# vss vss efet w=37765 l=7885
M1017 diff_296310_846600# vcc vcc vss efet w=8300 l=24900
M1020 q3 diff_644910_939560# vss vss efet w=350260 l=7470
M1021 vss diff_551950_771900# diff_536180_846600# vss efet w=67645 l=7885
M1022 diff_536180_846600# diff_207500_451520# vss vss efet w=39010 l=7470
M1025 diff_404210_938730# diff_296310_846600# vss vss efet w=54780 l=7470
M1030 q4 diff_296310_846600# vcc vss efet w=24900 l=7470
M1031 diff_404210_938730# vcc vcc vss efet w=9960 l=19920
M1032 diff_536180_846600# vcc vcc vss efet w=8300 l=24070
M1039 diff_312080_771900# diff_258130_451520# diff_278050_567720# vss efet w=14110 l=8300
M1040 diff_292990_681430# diff_258130_451520# diff_278050_567720# vss efet w=14110 l=7470
M1043 diff_278050_567720# diff_273900_607560# vss vss efet w=21995 l=7885
M1044 vcc vcc diff_278050_567720# vss efet w=8300 l=40670
M1045 q2 diff_884780_939560# vss vss efet w=350260 l=7470
M1046 vss diff_792650_771900# diff_776880_846600# vss efet w=68060 l=7470
M1047 diff_776880_846600# diff_207500_451520# vss vss efet w=39010 l=7470
M1050 diff_644910_939560# diff_536180_846600# vss vss efet w=54780 l=7470
M1055 q3 diff_536180_846600# vcc vss efet w=24070 l=7470
M1056 diff_644910_939560# vcc vcc vss efet w=9960 l=20750
M1057 diff_776880_846600# vcc vcc vss efet w=8300 l=24070
M1064 diff_551950_771900# diff_258130_451520# diff_510450_712970# vss efet w=14110 l=7470
M1067 diff_278050_567720# diff_232400_451520# diff_395080_711310# vss efet w=48970 l=7470
M1068 diff_510450_738700# diff_273900_560250# diff_390930_703840# vss efet w=14110 l=7470
M1071 vss diff_292990_681430# diff_273900_607560# vss efet w=37350 l=7470
M1072 diff_395080_711310# diff_390930_703840# vss vss efet w=78020 l=7470
M1073 vss diff_390930_685580# diff_395080_673960# vss efet w=78020 l=7470
M1076 diff_510450_712970# diff_273900_560250# diff_390930_685580# vss efet w=14110 l=7470
M1077 diff_532860_681430# diff_258130_451520# diff_510450_712970# vss efet w=14110 l=7470
M1080 diff_510450_712970# diff_510450_738700# vss vss efet w=22410 l=7470
M1081 vcc vcc diff_510450_712970# vss efet w=8300 l=39840
M1082 q1 diff_1125480_939560# vss vss efet w=351090 l=7470
M1083 vss diff_1032520_771900# diff_1016750_846600# vss efet w=68060 l=7470
M1084 diff_1016750_846600# diff_207500_451520# vss vss efet w=39010 l=7470
M1087 diff_884780_939560# diff_776880_846600# vss vss efet w=54780 l=7470
M1092 q2 diff_776880_846600# vcc vss efet w=24900 l=7470
M1093 diff_884780_939560# vcc vcc vss efet w=9960 l=19920
M1094 diff_1016750_846600# vcc vcc vss efet w=8300 l=24070
M1101 diff_792650_771900# diff_258130_451520# diff_751150_712970# vss efet w=14110 l=7470
M1104 diff_510450_712970# diff_232400_451520# diff_634950_712140# vss efet w=49800 l=7470
M1105 diff_751150_738700# diff_273900_560250# diff_630800_705500# vss efet w=14110 l=7470
M1108 diff_395080_673960# diff_232400_451520# diff_273900_607560# vss efet w=48970 l=7470
M1109 vss diff_341130_652380# diff_273900_607560# vss efet w=27390 l=7470
M1112 diff_273900_607560# vcc vcc vss efet w=8300 l=43160
M1113 vss diff_532860_681430# diff_510450_738700# vss efet w=37350 l=7470
M1114 diff_634950_712140# diff_630800_705500# vss vss efet w=78020 l=7470
M1115 vss diff_630800_686410# diff_634950_673960# vss efet w=78850 l=7470
M1118 diff_751150_712970# diff_273900_560250# diff_630800_686410# vss efet w=14110 l=7470
M1119 diff_773560_682260# diff_258130_451520# diff_751150_712970# vss efet w=14110 l=6640
M1122 diff_751150_712970# diff_751150_738700# vss vss efet w=22410 l=7470
M1123 diff_634950_673960# diff_232400_451520# diff_510450_738700# vss efet w=49800 l=7470
M1124 vss diff_341130_652380# diff_510450_738700# vss efet w=22410 l=7470
M1125 diff_510450_738700# vcc vcc vss efet w=8300 l=42330
M1126 vcc vcc diff_751150_712970# vss efet w=8300 l=39840
M1127 q0 diff_1365350_939560# vss vss efet w=350260 l=7470
M1128 vss diff_1273220_771900# diff_1257450_846600# vss efet w=67645 l=7055
M1129 diff_1257450_846600# diff_207500_451520# vss vss efet w=39010 l=7470
M1132 diff_1125480_939560# diff_1016750_846600# vss vss efet w=55195 l=7055
M1137 q1 diff_1016750_846600# vcc vss efet w=24900 l=7470
M1138 diff_1125480_939560# vcc vcc vss efet w=10790 l=19920
M1139 diff_1257450_846600# vcc vcc vss efet w=8300 l=24070
M1146 diff_1032520_771900# diff_258130_451520# diff_991020_712970# vss efet w=14110 l=7470
M1149 diff_751150_712970# diff_232400_451520# diff_875650_712140# vss efet w=48970 l=7470
M1150 diff_991020_738700# diff_273900_560250# diff_871500_704670# vss efet w=14110 l=7470
M1153 vss diff_773560_682260# diff_751150_738700# vss efet w=38180 l=7470
M1154 diff_875650_712140# diff_871500_704670# vss vss efet w=77190 l=7470
M1155 vss diff_871500_685580# diff_875650_674790# vss efet w=77605 l=7055
M1158 diff_991020_712970# diff_273900_560250# diff_871500_685580# vss efet w=14110 l=7470
M1159 diff_1013430_682260# diff_258130_451520# diff_991020_712970# vss efet w=14110 l=7470
M1162 diff_991020_712970# diff_991020_738700# vss vss efet w=22410 l=6640
M1163 vcc vcc diff_991020_712970# vss efet w=8300 l=39840
M1164 diff_1365350_939560# diff_1257450_846600# vss vss efet w=55610 l=7470
M1167 q0 diff_1257450_846600# vcc vss efet w=24900 l=7470
M1168 diff_1365350_939560# vcc vcc vss efet w=10375 l=20335
M1173 vss diff_1621820_879800# diff_232400_451520# vss efet w=149400 l=7470
M1174 vss diff_1505620_931260# diff_273900_560250# vss efet w=64740 l=7470
M1175 diff_273900_560250# vcc vcc vss efet w=10790 l=20750
M1176 diff_232400_451520# vcc vcc vss efet w=10790 l=9960
M1179 diff_1621820_879800# vcc vcc vss efet w=8300 l=24070
M1180 vss diff_1505620_931260# diff_1621820_879800# vss efet w=34030 l=7470
M1183 vss diff_1588620_812570# diff_1505620_931260# vss efet w=34030 l=8300
M1184 diff_1588620_812570# diff_1566210_789330# vss vss efet w=170150 l=22410
M1185 diff_1273220_771900# diff_258130_451520# diff_1231720_712970# vss efet w=14110 l=7470
M1188 diff_991020_712970# diff_232400_451520# diff_1115520_712140# vss efet w=49385 l=7055
M1189 diff_1231720_738700# diff_273900_560250# diff_1111370_704670# vss efet w=14110 l=7470
M1192 diff_875650_674790# diff_232400_451520# diff_751150_738700# vss efet w=49385 l=7055
M1193 vss diff_341130_652380# diff_751150_738700# vss efet w=22410 l=7470
M1194 diff_751150_738700# vcc vcc vss efet w=8300 l=41500
M1195 vss diff_1013430_682260# diff_991020_738700# vss efet w=38180 l=7470
M1196 diff_1115520_712140# diff_1111370_704670# vss vss efet w=78020 l=7470
M1197 vss diff_1111370_685580# diff_1115520_674790# vss efet w=78435 l=7885
M1200 diff_1231720_712970# diff_273900_560250# diff_1111370_685580# vss efet w=14110 l=7470
M1201 diff_1254960_682260# diff_258130_451520# diff_1231720_712970# vss efet w=14110 l=7470
M1204 diff_1231720_712970# diff_1231720_738700# vss vss efet w=22410 l=7470
M1205 vcc vcc diff_1231720_712970# vss efet w=8300 l=39840
M1206 diff_1477400_740360# vcc vcc vss efet w=6640 l=180940
M1207 diff_1505620_931260# vcc vcc vss efet w=8300 l=24900
M1208 vcc vcc diff_1588620_812570# vss efet w=8300 l=24070
M1211 data_in vss vss vss efet w=112880 l=8300
M1212 cp vss vss vss efet w=112880 l=8300
M1213 diff_1231720_712970# diff_232400_451520# diff_1355390_712140# vss efet w=50215 l=7885
M1214 diff_1115520_674790# diff_232400_451520# diff_991020_738700# vss efet w=49385 l=7055
M1215 vss diff_341130_652380# diff_991020_738700# vss efet w=22410 l=7470
M1216 diff_991020_738700# vcc vcc vss efet w=8300 l=41500
M1217 vss diff_1254960_682260# diff_1231720_738700# vss efet w=38180 l=7470
M1218 diff_1355390_712140# diff_1352070_704670# vss vss efet w=79680 l=7470
M1219 diff_1566210_789330# diff_1477400_740360# vss vss efet w=164340 l=23240
M1220 vss cp diff_1477400_740360# vss efet w=14110 l=7470
M1221 vss diff_1352070_685580# diff_1355390_674790# vss efet w=80925 l=7885
M1222 diff_1355390_674790# diff_232400_451520# diff_1231720_738700# vss efet w=49800 l=7470
M1223 vss diff_341130_652380# diff_1231720_738700# vss efet w=21580 l=7470
M1224 diff_1466610_655700# vcc vcc vss efet w=8300 l=22410
M1225 vss data_in diff_1466610_629970# vss efet w=163095 l=7885
M1226 vss diff_1466610_629970# diff_1466610_655700# vss efet w=50630 l=8300
M1229 diff_1466610_655700# diff_273900_560250# diff_1352070_704670# vss efet w=14110 l=7470
M1230 diff_1231720_738700# vcc vcc vss efet w=8300 l=41500
M1233 diff_1466610_629970# diff_273900_560250# diff_1352070_685580# vss efet w=14110 l=7470
M1236 diff_1466610_629970# vcc vcc vss efet w=10790 l=19920
M1238 vcc vcc diff_336150_519580# vss efet w=7885 l=42745
M1256 diff_278050_567720# diff_273900_560250# diff_278050_543650# vss efet w=14110 l=7470
M1257 diff_273900_607560# diff_273900_560250# diff_289670_464800# vss efet w=14110 l=7470
M1260 diff_336150_519580# diff_232400_451520# diff_322040_502150# vss efet w=48970 l=7470
M1261 diff_336150_519580# diff_341130_652380# vss vss efet w=21580 l=8300
M1262 diff_322040_502150# diff_278050_543650# vss vss efet w=77605 l=7885
M1263 vss diff_289670_464800# diff_305440_456500# vss efet w=78020 l=7470
M1264 diff_336150_519580# diff_415830_432430# vss vss efet w=37350 l=8300
M1265 diff_336150_427450# diff_232400_451520# diff_305440_456500# vss efet w=49385 l=7885
M1266 diff_336150_427450# vcc vcc vss efet w=8300 l=39840
M1267 vcc vcc diff_576020_519580# vss efet w=8300 l=42330
M1268 diff_576020_519580# diff_232400_451520# diff_544480_499660# vss efet w=49800 l=7470
M1269 diff_576020_519580# diff_341130_652380# vss vss efet w=22410 l=7470
M1270 diff_544480_499660# diff_512940_454840# vss vss efet w=79680 l=7470
M1271 vss diff_336150_519580# diff_336150_427450# vss efet w=21580 l=8300
M1274 diff_336150_427450# diff_258130_451520# diff_415830_432430# vss efet w=14110 l=7470
M1275 diff_512940_454840# diff_273900_560250# diff_336150_427450# vss efet w=12450 l=7470
M1277 diff_563570_456500# diff_512940_429940# vss vss efet w=76775 l=7885
M1278 diff_576020_519580# diff_656530_432430# vss vss efet w=38595 l=7885
M1279 diff_576020_427450# diff_232400_451520# diff_563570_456500# vss efet w=49800 l=7470
M1283 diff_512940_429940# diff_273900_560250# diff_336150_519580# vss efet w=12450 l=7470
M1286 diff_336150_427450# diff_258130_451520# diff_444050_322040# vss efet w=14110 l=7470
M1291 vcc vcc diff_275560_234060# vss efet w=10375 l=19920
M1292 vcc diff_314570_311250# q5 vss efet w=24900 l=8300
M1295 diff_275560_234060# diff_314570_311250# vss vss efet w=56025 l=7885
M1296 vss diff_275560_234060# q5 vss efet w=347355 l=7885
M1297 diff_576020_427450# vcc vcc vss efet w=8300 l=39840
M1298 vcc vcc diff_816720_520410# vss efet w=9130 l=42330
M1299 diff_816720_520410# diff_232400_451520# diff_786010_499660# vss efet w=49800 l=7470
M1300 diff_816720_520410# diff_341130_652380# vss vss efet w=22410 l=6640
M1301 diff_786010_499660# diff_754470_454010# vss vss efet w=78850 l=7470
M1302 vss diff_576020_519580# diff_576020_427450# vss efet w=21580 l=7470
M1305 diff_576020_427450# diff_258130_451520# diff_656530_432430# vss efet w=14110 l=7470
M1306 diff_754470_454010# diff_273900_560250# diff_576020_427450# vss efet w=13280 l=7470
M1308 diff_804270_456500# diff_754470_429110# vss vss efet w=77190 l=7470
M1309 diff_816720_520410# diff_896400_434090# vss vss efet w=38180 l=7470
M1310 diff_816720_427450# diff_232400_451520# diff_804270_456500# vss efet w=49800 l=7470
M1314 diff_754470_429110# diff_273900_560250# diff_576020_519580# vss efet w=13280 l=7470
M1317 diff_576020_427450# diff_258130_451520# diff_684750_321210# vss efet w=14110 l=7470
M1324 vcc vcc diff_314570_311250# vss efet w=7885 l=24485
M1325 vcc vcc diff_517090_234060# vss efet w=10790 l=19920
M1326 vcc diff_556100_312080# q6 vss efet w=24900 l=7470
M1331 diff_517090_234060# diff_556100_312080# vss vss efet w=56440 l=7470
M1334 vss diff_207500_451520# diff_314570_311250# vss efet w=39010 l=8300
M1335 diff_314570_311250# diff_444050_322040# vss vss efet w=67230 l=7470
M1336 vss diff_517090_234060# q6 vss efet w=347355 l=7885
M1337 diff_816720_427450# vcc vcc vss efet w=8300 l=39840
M1338 vcc vcc diff_1056590_520410# vss efet w=9130 l=42330
M1339 diff_1056590_520410# diff_232400_451520# diff_1025050_499660# vss efet w=49800 l=7470
M1340 diff_1056590_520410# diff_341130_652380# vss vss efet w=22410 l=7470
M1341 diff_1025050_499660# diff_993510_454010# vss vss efet w=79680 l=7470
M1342 vss diff_816720_520410# diff_816720_427450# vss efet w=21580 l=7470
M1345 diff_816720_427450# diff_258130_451520# diff_896400_434090# vss efet w=14110 l=7470
M1346 diff_993510_454010# diff_273900_560250# diff_816720_427450# vss efet w=13280 l=6640
M1348 diff_1043310_456500# diff_993510_429110# vss vss efet w=77605 l=7055
M1349 diff_1056590_520410# diff_1137100_433260# vss vss efet w=38180 l=7470
M1350 diff_1056590_427450# diff_232400_451520# diff_1043310_456500# vss efet w=49800 l=7470
M1354 diff_993510_429110# diff_273900_560250# diff_816720_520410# vss efet w=13280 l=6640
M1357 diff_816720_427450# diff_258130_451520# diff_924620_321210# vss efet w=14110 l=7470
M1364 vcc vcc diff_556100_312080# vss efet w=7885 l=25315
M1365 vcc vcc diff_756130_234890# vss efet w=10790 l=20750
M1366 vcc diff_795140_312080# q7 vss efet w=24900 l=7470
M1371 diff_756130_234890# diff_795140_312080# vss vss efet w=56025 l=7885
M1374 vss diff_207500_451520# diff_556100_312080# vss efet w=39010 l=7470
M1375 diff_556100_312080# diff_684750_321210# vss vss efet w=66815 l=7885
M1376 vss diff_756130_234890# q7 vss efet w=347355 l=7885
M1377 diff_1056590_427450# vcc vcc vss efet w=8300 l=39840
M1378 vcc vcc diff_1297290_520410# vss efet w=8300 l=42330
M1379 diff_341130_652380# vcc vcc vss efet w=8300 l=16600
M1380 vss diff_1483210_498830# diff_341130_652380# vss efet w=61835 l=7885
M1381 vcc vcc diff_1509770_516260# vss efet w=8300 l=62250
M1382 vcc vcc diff_1483210_498830# vss efet w=8715 l=23655
M1383 diff_1297290_520410# diff_232400_451520# diff_1266580_499660# vss efet w=48970 l=7470
M1384 diff_1297290_520410# diff_341130_652380# vss vss efet w=22410 l=8300
M1385 diff_1266580_499660# diff_1235040_454010# vss vss efet w=78020 l=7470
M1386 vss diff_1056590_520410# diff_1056590_427450# vss efet w=22410 l=7470
M1389 diff_1056590_427450# diff_258130_451520# diff_1137100_433260# vss efet w=14110 l=7470
M1390 diff_1235040_454010# diff_273900_560250# diff_1056590_427450# vss efet w=13280 l=7470
M1392 diff_1284840_456500# diff_1235040_429110# vss vss efet w=76360 l=7470
M1393 diff_1297290_520410# diff_1376970_433260# vss vss efet w=39840 l=7470
M1394 diff_1297290_428280# diff_232400_451520# diff_1284840_456500# vss efet w=48970 l=7470
M1398 diff_1235040_429110# diff_273900_560250# diff_1056590_520410# vss efet w=13280 l=7470
M1401 diff_1056590_427450# diff_258130_451520# diff_1165320_321210# vss efet w=14110 l=7470
M1408 vcc vcc diff_795140_312080# vss efet w=8300 l=24900
M1409 vcc vcc diff_994340_234060# vss efet w=9960 l=20750
M1410 vcc diff_1033350_312080# q8 vss efet w=24900 l=7470
M1415 diff_994340_234060# diff_1033350_312080# vss vss efet w=55610 l=7470
M1418 vss diff_207500_451520# diff_795140_312080# vss efet w=38595 l=7885
M1419 diff_795140_312080# diff_924620_321210# vss vss efet w=67230 l=7470
M1420 vss diff_994340_234060# q8 vss efet w=347770 l=7470
M1421 diff_1297290_428280# vcc vcc vss efet w=8300 l=40670
M1422 vss diff_1297290_520410# diff_1297290_428280# vss efet w=22410 l=7470
M1423 diff_1483210_498830# diff_1509770_516260# vss vss efet w=38180 l=7470
M1424 vcc vcc diff_1566210_789330# vss efet w=7885 l=180525
M1425 vss diff_1505620_931260# diff_1509770_516260# vss efet w=20335 l=7885
M1426 diff_1509770_516260# diff_1483210_498830# diff_1552100_502150# vss efet w=28220 l=7470
M1427 diff_1552100_502150# diff_1548780_494680# vss vss efet w=28220 l=8300
M1428 vss diff_1505620_352750# diff_1472420_424130# vss efet w=27805 l=7885
M1429 vss diff_273900_560250# diff_1472420_449860# vss efet w=68890 l=7470
M1430 vss diff_1472420_424130# diff_1505620_352750# vss efet w=34030 l=7470
M1434 diff_1297290_428280# diff_258130_451520# diff_1376970_433260# vss efet w=14110 l=7470
M1435 diff_1472420_449860# diff_1297290_520410# diff_1472420_424130# vss efet w=43990 l=7470
M1436 diff_1472420_449860# diff_1297290_428280# diff_1505620_352750# vss efet w=76360 l=7470
M1438 diff_1297290_428280# diff_258130_451520# diff_1405190_321210# vss efet w=14110 l=7470
M1439 vcc vcc diff_1505620_352750# vss efet w=8715 l=21995
M1440 diff_1472420_424130# vcc vcc vss efet w=8715 l=40255
M1447 vcc vcc diff_1033350_312080# vss efet w=8300 l=24900
M1448 vcc vcc diff_1236700_234890# vss efet w=10790 l=20750
M1449 vcc diff_1276540_312080# q9 vss efet w=24900 l=7470
M1454 diff_1236700_234890# diff_1276540_312080# vss vss efet w=55610 l=7470
M1457 vss diff_207500_451520# diff_1033350_312080# vss efet w=39010 l=7470
M1458 diff_1033350_312080# diff_1165320_321210# vss vss efet w=66400 l=7470
M1459 vss diff_1236700_234890# q9 vss efet w=349015 l=7885
M1464 diff_1548780_494680# vcc vcc vss efet w=6640 l=120350
M1469 vcc vcc diff_1276540_312080# vss efet w=8300 l=24900
M1470 vcc vcc diff_207500_451520# vss efet w=9960 l=18260
M1473 vcc diff_1505620_352750# serial_out vss efet w=49800 l=7470
M1476 diff_207500_451520# e vss vss efet w=166830 l=7470
M1479 vss diff_207500_451520# diff_1276540_312080# vss efet w=39425 l=7885
M1480 diff_1276540_312080# diff_1405190_321210# vss vss efet w=67230 l=7470
M1483 diff_1534670_282200# vcc vcc vss efet w=8300 l=16600
M1485 serial_out diff_1534670_282200# vss vss efet w=228665 l=7885
M1487 diff_1534670_282200# diff_1505620_352750# vss vss efet w=53120 l=7470
M1488 e vss vss vss efet w=111220 l=9130
