* SPICE3 file created from 4004.ext - technology: nmos

.option scale=0.01u

M1000 GND diff_51480_235440# diff_51960_227760# GND efet w=7440 l=960
+ ad=1.39029e+08 pd=2.33335e+07 as=5.17968e+07 ps=172080 
M1001 GND GND test GND efet w=9900 l=1260
+ ad=0 pd=0 as=5.60592e+07 ps=151200 
M1002 reset GND GND GND efet w=9780 l=1260
+ ad=5.69952e+07 pd=160080 as=0 ps=0 
M1003 GND diff_36720_291840# diff_42000_294000# GND efet w=2160 l=1080
+ ad=0 pd=0 as=2.48112e+07 ps=73200 
M1004 GND diff_75840_295200# diff_75240_295200# GND efet w=2520 l=1020
+ ad=0 pd=0 as=1.0944e+06 ps=5520 
M1005 diff_75240_295200# diff_73440_237000# diff_51480_235440# GND efet w=2160 l=1080
+ ad=0 pd=0 as=1.37506e+08 ps=438480 
M1006 GND diff_28560_293760# diff_36720_291840# GND efet w=1800 l=960
+ ad=0 pd=0 as=4.5648e+06 ps=11520 
M1007 diff_42000_294000# diff_28560_293760# diff_40800_290280# GND efet w=6480 l=960
+ ad=0 pd=0 as=6.9264e+06 ps=22080 
M1008 diff_36720_291840# GND GND GND efet w=600 l=5760
+ ad=0 pd=0 as=0 ps=0 
M1009 diff_36720_291840# GND GND GND efet w=1980 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1010 GND GND diff_42000_294000# GND efet w=720 l=2520
+ ad=0 pd=0 as=0 ps=0 
M1011 diff_40800_290280# GND GND GND efet w=10440 l=2520
+ ad=0 pd=0 as=0 ps=0 
M1012 GND diff_52080_238440# diff_50160_238320# GND efet w=3660 l=1140
+ ad=0 pd=0 as=7.4808e+07 ps=232080 
M1013 diff_51960_227760# diff_51960_227760# GND GND efet w=3660 l=1440
+ ad=0 pd=0 as=0 ps=0 
M1014 diff_51480_235440# diff_64920_237000# diff_42000_294000# GND efet w=1200 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1015 GND GND diff_27600_280080# GND efet w=1260 l=1020
+ ad=0 pd=0 as=6.1056e+06 ps=21120 
M1016 GND GND diff_28560_293760# GND efet w=420 l=1500
+ ad=0 pd=0 as=3.0528e+06 ps=12720 
M1017 GND diff_26520_220920# GND GND efet w=1740 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1018 diff_50160_238320# diff_50160_238320# GND GND efet w=2820 l=1800
+ ad=0 pd=0 as=0 ps=0 
M1019 diff_27240_279000# diff_26520_220920# GND GND efet w=1680 l=960
+ ad=2.2176e+06 pd=7200 as=0 ps=0 
M1020 diff_27600_280080# diff_27240_279000# diff_24720_257280# GND efet w=1200 l=1020
+ ad=0 pd=0 as=6.8832e+06 ps=20400 
M1021 diff_28560_293760# diff_27240_279000# diff_26760_257280# GND efet w=2160 l=960
+ ad=0 pd=0 as=4.4784e+06 ps=13680 
M1022 GND diff_27240_279000# diff_40800_274440# GND efet w=10200 l=960
+ ad=0 pd=0 as=6.6528e+06 ps=20160 
M1023 GND diff_4200_259560# GND GND efet w=101340 l=900
+ ad=0 pd=0 as=0 ps=0 
M1024 diff_4200_259560# diff_4200_259560# diff_4200_259560# GND efet w=5220 l=1680
+ ad=1.14336e+07 pd=44640 as=0 ps=0 
M1025 GND GND diff_4200_259560# GND efet w=480 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1026 GND diff_4200_259560# diff_4200_259560# GND efet w=840 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1027 GND GND GND GND efet w=5520 l=1320
+ ad=0 pd=0 as=0 ps=0 
M1028 GND GND GND GND efet w=960 l=960
+ ad=0 pd=0 as=0 ps=0 
M1029 GND GND GND GND efet w=540 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1030 GND GND GND GND efet w=51360 l=5940
+ ad=0 pd=0 as=0 ps=0 
M1031 diff_50160_238320# diff_50160_238320# GND GND efet w=2580 l=1860
+ ad=0 pd=0 as=0 ps=0 
M1032 GND GND diff_29880_257280# GND efet w=660 l=1620
+ ad=0 pd=0 as=3.0096e+06 ps=11040 
M1033 diff_42000_270960# diff_29880_257280# diff_40800_274440# GND efet w=5640 l=960
+ ad=2.39904e+07 pd=74160 as=0 ps=0 
M1034 GND diff_27240_279000# GND GND efet w=1920 l=840
+ ad=0 pd=0 as=0 ps=0 
M1035 GND GND GND GND efet w=600 l=5640
+ ad=0 pd=0 as=0 ps=0 
M1036 GND GND diff_42000_270960# GND efet w=600 l=2280
+ ad=0 pd=0 as=0 ps=0 
M1037 GND diff_29880_257280# GND GND efet w=1980 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1038 diff_42000_270960# GND GND GND efet w=1920 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1039 GND diff_36600_265200# diff_42000_267240# GND efet w=2160 l=960
+ ad=0 pd=0 as=2.33568e+07 ps=72960 
M1040 GND diff_31320_260160# diff_36600_265200# GND efet w=1980 l=960
+ ad=0 pd=0 as=5.1408e+06 ps=12000 
M1041 diff_42000_267240# diff_31320_260160# diff_40680_263760# GND efet w=5820 l=1020
+ ad=0 pd=0 as=6.3504e+06 ps=20640 
M1042 diff_36600_265200# GND GND GND efet w=660 l=5580
+ ad=0 pd=0 as=0 ps=0 
M1043 diff_36600_265200# GND GND GND efet w=1740 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1044 GND GND diff_42000_267240# GND efet w=660 l=2460
+ ad=0 pd=0 as=0 ps=0 
M1045 diff_40680_263760# GND GND GND efet w=9600 l=1800
+ ad=0 pd=0 as=0 ps=0 
M1046 diff_29880_257280# GND diff_29760_255720# GND efet w=1920 l=1560
+ ad=0 pd=0 as=864000 ps=4080 
M1047 diff_24720_257280# GND diff_24720_255720# GND efet w=1080 l=960
+ ad=0 pd=0 as=648000 ps=3360 
M1048 diff_26760_257280# GND diff_26760_255720# GND efet w=1920 l=960
+ ad=0 pd=0 as=1.152e+06 ps=5040 
M1049 GND GND diff_31320_260160# GND efet w=780 l=1140
+ ad=0 pd=0 as=5.7456e+06 ps=18960 
M1050 GND diff_26520_220920# GND GND efet w=1680 l=960
+ ad=0 pd=0 as=0 ps=0 
M1051 diff_42000_294000# diff_60240_235200# diff_51480_235440# GND efet w=1200 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1052 diff_51480_235440# diff_51480_235440# diff_42000_294000# GND efet w=780 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1053 diff_51480_235440# diff_51480_235440# diff_42000_270960# GND efet w=1320 l=960
+ ad=0 pd=0 as=0 ps=0 
M1054 diff_42000_270960# diff_60240_235200# diff_51480_235440# GND efet w=1320 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1055 GND diff_52080_238440# diff_54240_272160# GND efet w=3660 l=1020
+ ad=0 pd=0 as=1.27728e+07 ps=38400 
M1056 diff_51960_227760# diff_51960_227760# GND GND efet w=3480 l=1320
+ ad=0 pd=0 as=0 ps=0 
M1057 GND diff_52080_238440# diff_54240_263880# GND efet w=3660 l=1200
+ ad=0 pd=0 as=1.31472e+07 ps=38400 
M1058 diff_51960_227760# diff_51960_227760# GND GND efet w=4260 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1059 diff_50160_238320# diff_50160_238320# GND GND efet w=2640 l=1920
+ ad=0 pd=0 as=0 ps=0 
M1060 diff_24720_255720# diff_24240_254880# diff_24720_254040# GND efet w=1080 l=960
+ ad=0 pd=0 as=7.5312e+06 ps=25200 
M1061 diff_26760_255720# diff_24240_254880# diff_26760_254160# GND efet w=1920 l=960
+ ad=0 pd=0 as=9.3312e+06 ps=24720 
M1062 diff_29760_255720# diff_24240_254880# diff_26760_254160# GND efet w=1440 l=960
+ ad=0 pd=0 as=0 ps=0 
M1063 diff_31320_260160# diff_24240_254880# diff_26760_254160# GND efet w=720 l=960
+ ad=0 pd=0 as=0 ps=0 
M1064 diff_24240_254880# diff_26520_220920# GND GND efet w=1920 l=1020
+ ad=1.296e+06 pd=5280 as=0 ps=0 
M1065 GND diff_24240_254880# diff_40680_247920# GND efet w=10380 l=1020
+ ad=0 pd=0 as=6.552e+06 ps=20640 
M1066 diff_24720_254040# GND GND GND efet w=660 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1067 diff_50160_238320# diff_50160_238320# GND GND efet w=2760 l=1980
+ ad=0 pd=0 as=0 ps=0 
M1068 GND GND diff_36120_243120# GND efet w=900 l=1200
+ ad=0 pd=0 as=2.088e+06 ps=9360 
M1069 diff_42000_244200# diff_36120_243120# diff_40680_247920# GND efet w=5760 l=960
+ ad=2.39472e+07 pd=72960 as=0 ps=0 
M1070 GND diff_24240_254880# GND GND efet w=2400 l=960
+ ad=0 pd=0 as=0 ps=0 
M1071 GND GND GND GND efet w=660 l=5580
+ ad=0 pd=0 as=0 ps=0 
M1072 GND GND diff_42000_244200# GND efet w=600 l=2280
+ ad=0 pd=0 as=0 ps=0 
M1073 GND GND diff_26760_254160# GND efet w=2160 l=1560
+ ad=0 pd=0 as=0 ps=0 
M1074 GND diff_36120_243120# GND GND efet w=1800 l=840
+ ad=0 pd=0 as=0 ps=0 
M1075 diff_36120_243120# GND GND GND efet w=1200 l=960
+ ad=0 pd=0 as=0 ps=0 
M1076 diff_42000_244200# GND GND GND efet w=2160 l=960
+ ad=0 pd=0 as=0 ps=0 
M1077 GND GND diff_4200_259560# GND efet w=7500 l=1980
+ ad=0 pd=0 as=0 ps=0 
M1078 diff_24720_254040# GND diff_28320_238920# GND efet w=1200 l=960
+ ad=0 pd=0 as=3.1248e+06 ps=11040 
M1079 GND GND GND GND efet w=8160 l=2280
+ ad=0 pd=0 as=0 ps=0 
M1080 GND diff_87000_295200# diff_86400_294960# GND efet w=2160 l=1200
+ ad=0 pd=0 as=950400 ps=5520 
M1081 diff_82800_293280# diff_81000_291840# GND GND efet w=1620 l=900
+ ad=1.2096e+06 pd=5520 as=0 ps=0 
M1082 diff_51480_235440# diff_51480_235440# diff_82800_293280# GND efet w=2220 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1083 diff_86400_294960# diff_85440_237000# diff_51480_235440# GND efet w=2160 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1084 diff_51480_235440# diff_51480_235440# diff_93960_293280# GND efet w=2280 l=1080
+ ad=0 pd=0 as=1.2096e+06 ps=6000 
M1085 diff_93960_293280# diff_92280_291840# GND GND efet w=1920 l=960
+ ad=0 pd=0 as=0 ps=0 
M1086 diff_50160_238320# diff_51480_235440# GND GND efet w=6000 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1087 diff_51960_227760# diff_75720_237120# diff_75840_295200# GND efet w=540 l=1020
+ ad=0 pd=0 as=360000 ps=2640 
M1088 diff_81000_291840# diff_78120_238200# diff_51960_227760# GND efet w=660 l=900
+ ad=316800 pd=2640 as=0 ps=0 
M1089 diff_50160_238320# diff_75720_237120# diff_75840_287400# GND efet w=540 l=1020
+ ad=0 pd=0 as=345600 ps=2400 
M1090 diff_81000_290400# diff_78120_238200# diff_50160_238320# GND efet w=480 l=840
+ ad=345600 pd=2400 as=0 ps=0 
M1091 diff_75120_287520# diff_73440_237000# diff_51480_235440# GND efet w=2280 l=960
+ ad=1.1664e+06 pd=5760 as=0 ps=0 
M1092 GND diff_75840_287400# diff_75120_287520# GND efet w=2100 l=1260
+ ad=0 pd=0 as=0 ps=0 
M1093 diff_51960_227760# diff_50160_238320# diff_87000_295200# GND efet w=540 l=1020
+ ad=0 pd=0 as=360000 ps=2640 
M1094 diff_92280_291840# diff_51480_235440# diff_51960_227760# GND efet w=480 l=960
+ ad=302400 pd=2400 as=0 ps=0 
M1095 diff_50160_238320# diff_50160_238320# diff_87000_287520# GND efet w=420 l=1140
+ ad=0 pd=0 as=345600 ps=2400 
M1096 GND diff_51480_235440# diff_50160_238320# GND efet w=6000 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1097 diff_75240_286080# diff_73440_237000# diff_51480_235440# GND efet w=2040 l=900
+ ad=1.0512e+06 pd=5520 as=0 ps=0 
M1098 GND diff_75840_286320# diff_75240_286080# GND efet w=2040 l=1260
+ ad=0 pd=0 as=0 ps=0 
M1099 diff_82800_287520# diff_81000_290400# GND GND efet w=1860 l=1140
+ ad=1.2816e+06 pd=6000 as=0 ps=0 
M1100 diff_51480_235440# diff_51480_235440# diff_82800_287520# GND efet w=1860 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1101 diff_86400_287400# diff_85440_237000# diff_51480_235440# GND efet w=2220 l=900
+ ad=1.3824e+06 pd=5760 as=0 ps=0 
M1102 GND diff_87000_287520# diff_86400_287400# GND efet w=1980 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1103 diff_50160_238320# diff_51480_235440# GND GND efet w=5880 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1104 diff_50160_238320# diff_75720_237120# diff_75840_286320# GND efet w=660 l=1020
+ ad=0 pd=0 as=388800 ps=3120 
M1105 diff_82800_284400# diff_81000_282960# GND GND efet w=1980 l=1260
+ ad=1.2816e+06 pd=5760 as=0 ps=0 
M1106 diff_92280_290400# diff_51480_235440# diff_50160_238320# GND efet w=480 l=1080
+ ad=360000 pd=2880 as=0 ps=0 
M1107 GND diff_86760_205920# diff_51480_235440# GND efet w=720 l=960
+ ad=0 pd=0 as=0 ps=0 
M1108 GND diff_26520_220920# GND GND efet w=1200 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1109 GND diff_123240_258000# diff_117960_263280# GND efet w=1440 l=1080
+ ad=0 pd=0 as=2.72376e+08 ps=860160 
M1110 GND diff_117960_263280# diff_117840_290880# GND efet w=5280 l=960
+ ad=0 pd=0 as=1.48032e+07 ps=48000 
M1111 GND GND diff_51960_227760# GND efet w=540 l=2580
+ ad=0 pd=0 as=0 ps=0 
M1112 GND GND GND GND efet w=8400 l=1680
+ ad=0 pd=0 as=0 ps=0 
M1113 GND GND diff_50160_238320# GND efet w=540 l=2580
+ ad=0 pd=0 as=0 ps=0 
M1114 GND diff_87120_286080# diff_86400_286080# GND efet w=2100 l=1020
+ ad=0 pd=0 as=1.3104e+06 ps=5760 
M1115 diff_51480_235440# diff_51480_235440# diff_82800_284400# GND efet w=1620 l=1440
+ ad=0 pd=0 as=0 ps=0 
M1116 diff_86400_286080# diff_85440_237000# diff_51480_235440# GND efet w=2220 l=900
+ ad=0 pd=0 as=0 ps=0 
M1117 diff_93960_288000# diff_92280_290400# GND GND efet w=1980 l=1140
+ ad=1.2528e+06 pd=5520 as=0 ps=0 
M1118 diff_51480_235440# diff_51480_235440# diff_93960_288000# GND efet w=2220 l=900
+ ad=0 pd=0 as=0 ps=0 
M1119 GND diff_86760_205920# diff_51480_235440# GND efet w=780 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1120 GND GND diff_117840_290880# GND efet w=3600 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1121 diff_117960_263280# diff_117960_263280# GND GND efet w=3420 l=1440
+ ad=0 pd=0 as=0 ps=0 
M1122 GND GND GND GND efet w=660 l=1860
+ ad=0 pd=0 as=0 ps=0 
M1123 diff_93960_284400# diff_92280_282960# GND GND efet w=1980 l=1140
+ ad=1.296e+06 pd=5760 as=0 ps=0 
M1124 diff_51480_235440# diff_51480_235440# diff_93960_284400# GND efet w=2340 l=900
+ ad=0 pd=0 as=0 ps=0 
M1125 diff_81000_282960# diff_78120_238200# diff_50160_238320# GND efet w=540 l=840
+ ad=374400 pd=2640 as=0 ps=0 
M1126 diff_50160_238320# diff_75720_237120# diff_75840_278520# GND efet w=480 l=840
+ ad=0 pd=0 as=345600 ps=2400 
M1127 diff_81000_281520# diff_78120_238200# diff_50160_238320# GND efet w=480 l=840
+ ad=345600 pd=2400 as=0 ps=0 
M1128 diff_75120_278520# diff_73440_237000# diff_51480_235440# GND efet w=2340 l=900
+ ad=1.1808e+06 pd=6000 as=0 ps=0 
M1129 GND diff_75840_278520# diff_75120_278520# GND efet w=2040 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1130 diff_50160_238320# diff_50160_238320# diff_87120_286080# GND efet w=360 l=1200
+ ad=0 pd=0 as=374400 ps=2880 
M1131 GND diff_86760_205920# diff_51480_235440# GND efet w=780 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1132 GND GND GND GND efet w=660 l=1740
+ ad=0 pd=0 as=0 ps=0 
M1133 diff_92280_282960# diff_51480_235440# diff_50160_238320# GND efet w=480 l=960
+ ad=345600 pd=2400 as=0 ps=0 
M1134 diff_50160_238320# diff_50160_238320# diff_87000_278520# GND efet w=420 l=960
+ ad=0 pd=0 as=345600 ps=2400 
M1135 diff_92280_281520# diff_51480_235440# diff_50160_238320# GND efet w=480 l=960
+ ad=374400 pd=2640 as=0 ps=0 
M1136 GND diff_51480_235440# diff_54240_272160# GND efet w=5280 l=960
+ ad=0 pd=0 as=0 ps=0 
M1137 GND diff_51480_235440# diff_51960_227760# GND efet w=5700 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1138 diff_51480_235440# diff_64920_237000# diff_42000_270960# GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M1139 diff_75240_277200# diff_73440_237000# diff_51480_235440# GND efet w=2040 l=900
+ ad=1.0512e+06 pd=5280 as=0 ps=0 
M1140 GND diff_75840_277320# diff_75240_277200# GND efet w=2040 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1141 diff_82680_279240# diff_81000_281520# GND GND efet w=1980 l=1140
+ ad=1.2096e+06 pd=5760 as=0 ps=0 
M1142 diff_51480_235440# diff_51480_235440# diff_82680_279240# GND efet w=1740 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1143 diff_86400_278520# diff_85440_237000# diff_51480_235440# GND efet w=2220 l=900
+ ad=1.3536e+06 pd=5760 as=0 ps=0 
M1144 GND diff_87000_278520# diff_86400_278520# GND efet w=2040 l=960
+ ad=0 pd=0 as=0 ps=0 
M1145 GND GND GND GND efet w=9180 l=1260
+ ad=0 pd=0 as=0 ps=0 
M1146 GND GND diff_50160_238320# GND efet w=600 l=2640
+ ad=0 pd=0 as=0 ps=0 
M1147 GND GND diff_50160_238320# GND efet w=540 l=2580
+ ad=0 pd=0 as=0 ps=0 
M1148 diff_93960_279120# diff_92280_281520# GND GND efet w=1980 l=1500
+ ad=1.2816e+06 pd=5760 as=0 ps=0 
M1149 diff_82800_275640# diff_81000_274080# GND GND efet w=1860 l=1260
+ ad=1.1232e+06 pd=5520 as=0 ps=0 
M1150 GND diff_87000_277320# diff_86400_276960# GND efet w=1980 l=1020
+ ad=0 pd=0 as=1.2816e+06 ps=5520 
M1151 diff_51480_235440# diff_51480_235440# diff_82800_275640# GND efet w=1800 l=1320
+ ad=0 pd=0 as=0 ps=0 
M1152 diff_86400_276960# diff_85440_237000# diff_51480_235440# GND efet w=2100 l=900
+ ad=0 pd=0 as=0 ps=0 
M1153 diff_51480_235440# diff_51480_235440# diff_93960_279120# GND efet w=1800 l=1320
+ ad=0 pd=0 as=0 ps=0 
M1154 GND diff_86760_205920# diff_51480_235440# GND efet w=720 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1155 GND GND diff_117960_280920# GND efet w=3600 l=1080
+ ad=0 pd=0 as=1.42416e+07 ps=46320 
M1156 diff_117960_263280# diff_117960_263280# GND GND efet w=3420 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1157 diff_117960_263280# diff_117960_263280# GND GND efet w=720 l=1500
+ ad=0 pd=0 as=0 ps=0 
M1158 diff_117960_263280# diff_117960_263280# GND GND efet w=4920 l=960
+ ad=0 pd=0 as=0 ps=0 
M1159 diff_138480_294720# diff_117960_263280# diff_117960_263280# GND efet w=1560 l=1560
+ ad=964800 pd=5280 as=0 ps=0 
M1160 GND GND diff_138480_294720# GND efet w=2100 l=1260
+ ad=0 pd=0 as=0 ps=0 
M1161 diff_146040_293280# diff_144240_291720# GND GND efet w=2040 l=1200
+ ad=921600 pd=5040 as=0 ps=0 
M1162 diff_117960_263280# diff_117960_263280# diff_146040_293280# GND efet w=1620 l=1500
+ ad=0 pd=0 as=0 ps=0 
M1163 diff_149640_294720# diff_117960_263280# diff_117960_263280# GND efet w=1800 l=1440
+ ad=1.152e+06 pd=5280 as=0 ps=0 
M1164 GND diff_150240_291840# diff_149640_294720# GND efet w=1980 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1165 diff_157200_293280# diff_155400_291720# GND GND efet w=2100 l=1380
+ ad=892800 pd=5040 as=0 ps=0 
M1166 diff_117960_263280# diff_117960_263280# diff_157200_293280# GND efet w=1680 l=1500
+ ad=0 pd=0 as=0 ps=0 
M1167 diff_160800_294960# diff_117960_263280# diff_117960_263280# GND efet w=1740 l=1620
+ ad=936000 pd=5520 as=0 ps=0 
M1168 GND diff_161280_294840# diff_160800_294960# GND efet w=2220 l=1620
+ ad=0 pd=0 as=0 ps=0 
M1169 diff_168360_293160# diff_166560_291720# GND GND efet w=2100 l=1140
+ ad=864000 pd=5760 as=0 ps=0 
M1170 diff_117840_290880# diff_139680_254520# GND GND efet w=480 l=960
+ ad=0 pd=0 as=0 ps=0 
M1171 diff_144240_291720# diff_142200_254520# diff_117840_290880# GND efet w=480 l=960
+ ad=302400 pd=2400 as=0 ps=0 
M1172 diff_117840_290880# diff_151440_254520# diff_150240_291840# GND efet w=540 l=1020
+ ad=0 pd=0 as=316800 ps=2640 
M1173 diff_117960_263280# diff_139680_254520# diff_138960_287280# GND efet w=480 l=960
+ ad=0 pd=0 as=288000 ps=2160 
M1174 diff_144240_290280# diff_142200_254520# diff_117960_263280# GND efet w=480 l=960
+ ad=316800 pd=2640 as=0 ps=0 
M1175 diff_138360_287280# diff_117960_263280# diff_117960_263280# GND efet w=2280 l=1080
+ ad=1.2096e+06 pd=5760 as=0 ps=0 
M1176 GND diff_138960_287280# diff_138360_287280# GND efet w=2040 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1177 diff_155400_291720# diff_153840_254520# diff_117840_290880# GND efet w=480 l=960
+ ad=345600 pd=2400 as=0 ps=0 
M1178 GND diff_138960_286080# diff_138360_286080# GND efet w=1980 l=1140
+ ad=0 pd=0 as=1.1232e+06 ps=5520 
M1179 GND diff_26520_220920# GND GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M1180 diff_93960_275640# diff_92160_274080# GND GND efet w=2040 l=1380
+ ad=1.2096e+06 pd=5520 as=0 ps=0 
M1181 diff_51480_235440# diff_51480_235440# diff_93960_275640# GND efet w=1620 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1182 diff_54240_272160# diff_75720_237120# diff_75840_277320# GND efet w=660 l=1020
+ ad=0 pd=0 as=460800 ps=2880 
M1183 diff_81000_274080# diff_78120_238200# diff_54240_272160# GND efet w=480 l=1020
+ ad=403200 pd=3120 as=0 ps=0 
M1184 diff_51960_227760# diff_75720_237120# diff_75840_269640# GND efet w=480 l=840
+ ad=0 pd=0 as=403200 ps=2640 
M1185 diff_81000_272640# diff_78120_238200# diff_51960_227760# GND efet w=480 l=840
+ ad=345600 pd=2400 as=0 ps=0 
M1186 diff_75120_269640# diff_73440_237000# diff_51480_235440# GND efet w=2280 l=900
+ ad=1.1952e+06 pd=5760 as=0 ps=0 
M1187 GND diff_75840_269640# diff_75120_269640# GND efet w=1980 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1188 diff_54240_272160# diff_50160_238320# diff_87000_277320# GND efet w=540 l=900
+ ad=0 pd=0 as=374400 ps=2880 
M1189 diff_92160_274080# diff_51480_235440# diff_54240_272160# GND efet w=480 l=840
+ ad=403200 pd=2640 as=0 ps=0 
M1190 diff_51960_227760# diff_50160_238320# diff_87000_269640# GND efet w=480 l=840
+ ad=0 pd=0 as=345600 ps=2400 
M1191 diff_92160_272640# diff_51480_235440# diff_51960_227760# GND efet w=480 l=840
+ ad=403200 pd=2640 as=0 ps=0 
M1192 GND diff_51480_235440# diff_51960_227760# GND efet w=6060 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1193 diff_51480_235440# diff_64920_237000# diff_42000_267240# GND efet w=1200 l=900
+ ad=0 pd=0 as=0 ps=0 
M1194 diff_42000_267240# diff_60240_235200# diff_51480_235440# GND efet w=1200 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1195 diff_75120_268440# diff_73440_237000# diff_51480_235440# GND efet w=2220 l=900
+ ad=1.0944e+06 pd=5520 as=0 ps=0 
M1196 GND diff_75840_268440# diff_75120_268440# GND efet w=2040 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1197 diff_82800_269880# diff_81000_272640# GND GND efet w=1920 l=1200
+ ad=1.2528e+06 pd=5520 as=0 ps=0 
M1198 diff_51480_235440# diff_51480_235440# diff_82800_269880# GND efet w=2160 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1199 diff_86400_269640# diff_85440_237000# diff_51480_235440# GND efet w=2280 l=960
+ ad=1.368e+06 pd=5760 as=0 ps=0 
M1200 GND diff_87000_269640# diff_86400_269640# GND efet w=2040 l=960
+ ad=0 pd=0 as=0 ps=0 
M1201 GND diff_86760_205920# diff_51480_235440# GND efet w=720 l=960
+ ad=0 pd=0 as=0 ps=0 
M1202 GND diff_26520_220920# GND GND efet w=1200 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1203 diff_51480_235440# diff_51480_235440# diff_42000_267240# GND efet w=1200 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1204 diff_51480_235440# diff_51480_235440# diff_42000_244200# GND efet w=1260 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1205 diff_54240_263880# diff_51480_235440# GND GND efet w=5460 l=900
+ ad=0 pd=0 as=0 ps=0 
M1206 diff_51960_227760# diff_75720_237120# diff_75840_268440# GND efet w=540 l=1080
+ ad=0 pd=0 as=388800 ps=2880 
M1207 diff_82680_266760# diff_81000_265200# GND GND efet w=1920 l=1200
+ ad=1.3392e+06 pd=5520 as=0 ps=0 
M1208 GND diff_87000_268440# diff_86280_268320# GND efet w=2160 l=1080
+ ad=0 pd=0 as=1.2528e+06 ps=5760 
M1209 diff_51480_235440# diff_51480_235440# diff_82680_266760# GND efet w=2040 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1210 diff_86280_268320# diff_85440_237000# diff_51480_235440# GND efet w=2160 l=960
+ ad=0 pd=0 as=0 ps=0 
M1211 diff_93960_270120# diff_92160_272640# GND GND efet w=2040 l=1080
+ ad=1.2384e+06 pd=5520 as=0 ps=0 
M1212 diff_51480_235440# diff_51480_235440# diff_93960_270120# GND efet w=1800 l=1320
+ ad=0 pd=0 as=0 ps=0 
M1213 GND GND diff_54240_272160# GND efet w=540 l=2460
+ ad=0 pd=0 as=0 ps=0 
M1214 GND GND diff_117960_263280# GND efet w=3600 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1215 GND GND GND GND efet w=8340 l=1620
+ ad=0 pd=0 as=0 ps=0 
M1216 GND GND diff_51960_227760# GND efet w=540 l=2460
+ ad=0 pd=0 as=0 ps=0 
M1217 GND diff_86760_205920# diff_51480_235440# GND efet w=840 l=960
+ ad=0 pd=0 as=0 ps=0 
M1218 diff_117960_263280# diff_117960_263280# GND GND efet w=660 l=1500
+ ad=0 pd=0 as=0 ps=0 
M1219 GND diff_123240_258000# diff_117960_263280# GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M1220 GND diff_123240_258000# diff_117960_263280# GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M1221 diff_93960_266640# diff_92160_265200# GND GND efet w=2100 l=1140
+ ad=1.224e+06 pd=5520 as=0 ps=0 
M1222 diff_81000_265200# diff_78120_238200# diff_51960_227760# GND efet w=480 l=960
+ ad=360000 pd=2640 as=0 ps=0 
M1223 diff_81000_263760# diff_78120_238200# diff_54240_263880# GND efet w=480 l=1080
+ ad=345600 pd=2400 as=0 ps=0 
M1224 diff_54240_263880# diff_75720_237120# diff_75840_260760# GND efet w=480 l=960
+ ad=0 pd=0 as=345600 ps=2400 
M1225 diff_75120_260760# diff_73440_237000# diff_51480_235440# GND efet w=2340 l=900
+ ad=1.2384e+06 pd=5760 as=0 ps=0 
M1226 GND diff_75840_260760# diff_75120_260760# GND efet w=1980 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1227 diff_51960_227760# diff_50160_238320# diff_87000_268440# GND efet w=480 l=840
+ ad=0 pd=0 as=360000 ps=2640 
M1228 diff_51480_235440# diff_51480_235440# diff_93960_266640# GND efet w=1740 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1229 diff_92160_265200# diff_51480_235440# diff_51960_227760# GND efet w=480 l=840
+ ad=360000 pd=2640 as=0 ps=0 
M1230 diff_54240_263880# diff_50160_238320# diff_87000_260760# GND efet w=480 l=840
+ ad=0 pd=0 as=345600 ps=2400 
M1231 diff_82680_261240# diff_81000_263760# GND GND efet w=1980 l=1020
+ ad=1.3968e+06 pd=6000 as=0 ps=0 
M1232 GND diff_75840_259440# diff_75120_259560# GND efet w=2100 l=1140
+ ad=0 pd=0 as=1.1088e+06 ps=5520 
M1233 GND diff_51480_235440# diff_50160_238320# GND efet w=5760 l=960
+ ad=0 pd=0 as=0 ps=0 
M1234 diff_75120_259560# diff_73440_237000# diff_51480_235440# GND efet w=2100 l=900
+ ad=0 pd=0 as=0 ps=0 
M1235 diff_51480_235440# diff_51480_235440# diff_82680_261240# GND efet w=2220 l=900
+ ad=0 pd=0 as=0 ps=0 
M1236 diff_86400_260760# diff_85440_237000# diff_51480_235440# GND efet w=2160 l=960
+ ad=1.2816e+06 pd=6000 as=0 ps=0 
M1237 GND diff_87000_260760# diff_86400_260760# GND efet w=2160 l=960
+ ad=0 pd=0 as=0 ps=0 
M1238 diff_92160_263760# diff_51480_235440# diff_54240_263880# GND efet w=480 l=960
+ ad=345600 pd=2400 as=0 ps=0 
M1239 diff_93960_261240# diff_92160_263760# GND GND efet w=1980 l=1140
+ ad=1.152e+06 pd=5280 as=0 ps=0 
M1240 diff_51480_235440# diff_51480_235440# diff_93960_261240# GND efet w=1620 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1241 diff_50160_238320# diff_51480_235440# GND GND efet w=5640 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1242 diff_50160_238320# diff_75720_237120# diff_75840_259440# GND efet w=480 l=960
+ ad=0 pd=0 as=345600 ps=2400 
M1243 diff_82680_258240# diff_81000_256320# GND GND efet w=2040 l=1080
+ ad=1.3104e+06 pd=6000 as=0 ps=0 
M1244 GND diff_87000_259560# diff_86400_259200# GND efet w=1980 l=1020
+ ad=0 pd=0 as=1.296e+06 ps=5520 
M1245 diff_51480_235440# diff_51480_235440# diff_82680_258240# GND efet w=2100 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1246 diff_86400_259200# diff_85440_237000# diff_51480_235440# GND efet w=2160 l=960
+ ad=0 pd=0 as=0 ps=0 
M1247 GND GND GND GND efet w=600 l=1680
+ ad=0 pd=0 as=0 ps=0 
M1248 GND diff_86760_205920# diff_51480_235440# GND efet w=780 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1249 GND GND diff_51960_227760# GND efet w=480 l=2520
+ ad=0 pd=0 as=0 ps=0 
M1250 diff_109920_264000# GND GND GND efet w=660 l=1680
+ ad=1.35936e+07 pd=41520 as=0 ps=0 
M1251 GND diff_109920_264000# diff_109920_264000# GND efet w=9180 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1252 diff_117960_263280# diff_117960_263280# GND GND efet w=3300 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1253 GND diff_117960_263280# diff_117960_263280# GND efet w=4920 l=960
+ ad=0 pd=0 as=0 ps=0 
M1254 diff_117960_280920# diff_117960_263280# GND GND efet w=4980 l=900
+ ad=0 pd=0 as=0 ps=0 
M1255 diff_138360_286080# diff_117960_263280# diff_117960_263280# GND efet w=2160 l=960
+ ad=0 pd=0 as=0 ps=0 
M1256 diff_145920_287880# diff_144240_290280# GND GND efet w=2400 l=1200
+ ad=1.1232e+06 pd=6000 as=0 ps=0 
M1257 diff_117960_263280# diff_117960_263280# diff_145920_287880# GND efet w=2280 l=960
+ ad=0 pd=0 as=0 ps=0 
M1258 diff_149520_287400# diff_117960_263280# diff_117960_263280# GND efet w=2160 l=1080
+ ad=1.152e+06 pd=5520 as=0 ps=0 
M1259 diff_117960_263280# diff_151440_254520# diff_150240_287160# GND efet w=480 l=960
+ ad=0 pd=0 as=288000 ps=2160 
M1260 GND diff_150240_287160# diff_149520_287400# GND efet w=1800 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1261 diff_145920_284400# diff_144240_282840# GND GND efet w=2220 l=1260
+ ad=1.152e+06 pd=6240 as=0 ps=0 
M1262 diff_117960_263280# diff_139680_254520# diff_138960_286080# GND efet w=480 l=960
+ ad=0 pd=0 as=331200 ps=2640 
M1263 diff_155400_290280# diff_153840_254520# diff_117960_263280# GND efet w=480 l=960
+ ad=345600 pd=2400 as=0 ps=0 
M1264 diff_157200_287760# diff_155400_290280# GND GND efet w=2040 l=1320
+ ad=921600 pd=5280 as=0 ps=0 
M1265 diff_117960_263280# diff_167640_254400# diff_168360_293160# GND efet w=2520 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1266 diff_171960_294720# diff_117960_263280# diff_117960_263280# GND efet w=2280 l=1080
+ ad=892800 pd=5520 as=0 ps=0 
M1267 GND diff_172440_294840# diff_171960_294720# GND efet w=2220 l=1560
+ ad=0 pd=0 as=0 ps=0 
M1268 diff_179520_293160# diff_177840_291720# GND GND efet w=2280 l=1080
+ ad=820800 pd=5520 as=0 ps=0 
M1269 diff_117960_263280# diff_179280_254400# diff_179520_293160# GND efet w=2400 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1270 diff_117960_263280# diff_117960_263280# diff_157200_287760# GND efet w=1980 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1271 diff_117840_290880# diff_117960_263280# diff_161280_294840# GND efet w=480 l=1080
+ ad=0 pd=0 as=302400 ps=2400 
M1272 diff_166560_291720# diff_117960_263280# diff_117840_290880# GND efet w=660 l=1020
+ ad=273600 pd=2400 as=0 ps=0 
M1273 diff_117960_263280# diff_117960_263280# diff_161400_287160# GND efet w=600 l=1080
+ ad=0 pd=0 as=288000 ps=2160 
M1274 GND diff_161400_287160# diff_160800_287280# GND efet w=1800 l=1200
+ ad=0 pd=0 as=1.152e+06 ps=5280 
M1275 diff_166560_290280# diff_117960_263280# diff_117960_263280# GND efet w=540 l=1020
+ ad=316800 pd=2400 as=0 ps=0 
M1276 diff_160800_287280# diff_117960_263280# diff_117960_263280# GND efet w=1680 l=1320
+ ad=0 pd=0 as=0 ps=0 
M1277 GND diff_150240_286080# diff_149520_286080# GND efet w=1920 l=1260
+ ad=0 pd=0 as=1.1664e+06 ps=5760 
M1278 diff_117960_263280# diff_117960_263280# diff_145920_284400# GND efet w=2280 l=960
+ ad=0 pd=0 as=0 ps=0 
M1279 diff_149520_286080# diff_117960_263280# diff_117960_263280# GND efet w=2100 l=900
+ ad=0 pd=0 as=0 ps=0 
M1280 diff_117840_290880# diff_174360_263520# diff_172440_294840# GND efet w=480 l=1080
+ ad=0 pd=0 as=288000 ps=2160 
M1281 diff_177840_291720# diff_117960_263280# diff_117840_290880# GND efet w=480 l=1200
+ ad=230400 pd=1920 as=0 ps=0 
M1282 diff_117960_263280# diff_174360_263520# diff_172680_287040# GND efet w=600 l=1140
+ ad=0 pd=0 as=316800 ps=2400 
M1283 diff_157080_284280# diff_155400_282840# GND GND efet w=2100 l=1380
+ ad=1.1376e+06 pd=6240 as=0 ps=0 
M1284 diff_117960_263280# diff_117960_263280# diff_157080_284280# GND efet w=2280 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1285 diff_144240_282840# diff_142200_254520# diff_117960_263280# GND efet w=480 l=960
+ ad=345600 pd=2400 as=0 ps=0 
M1286 diff_117960_280920# diff_139680_254520# diff_139080_278280# GND efet w=480 l=960
+ ad=0 pd=0 as=288000 ps=2160 
M1287 diff_144240_281400# diff_142200_254520# diff_117960_280920# GND efet w=480 l=960
+ ad=345600 pd=2400 as=0 ps=0 
M1288 diff_138360_278640# diff_117960_263280# diff_117960_263280# GND efet w=2280 l=960
+ ad=1.1376e+06 pd=5520 as=0 ps=0 
M1289 GND diff_139080_278280# diff_138360_278640# GND efet w=1920 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1290 diff_117960_263280# diff_151440_254520# diff_150240_286080# GND efet w=540 l=900
+ ad=0 pd=0 as=331200 ps=2640 
M1291 diff_160800_285840# diff_117960_263280# diff_117960_263280# GND efet w=1740 l=1440
+ ad=1.1952e+06 pd=5520 as=0 ps=0 
M1292 GND diff_161400_286080# diff_160800_285840# GND efet w=1860 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1293 diff_168360_287640# diff_166560_290280# GND GND efet w=2220 l=1140
+ ad=878400 pd=5280 as=0 ps=0 
M1294 diff_117960_263280# diff_167640_254400# diff_168360_287640# GND efet w=2100 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1295 diff_171960_287280# diff_117960_263280# diff_117960_263280# GND efet w=1740 l=1380
+ ad=1.2096e+06 pd=5280 as=0 ps=0 
M1296 GND diff_172680_287040# diff_171960_287280# GND efet w=1680 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1297 GND diff_117960_263280# diff_117960_263280# GND efet w=660 l=1260
+ ad=0 pd=0 as=0 ps=0 
M1298 diff_168360_284280# diff_166560_282840# GND GND efet w=2160 l=1080
+ ad=936000 pd=5520 as=0 ps=0 
M1299 diff_117960_263280# diff_167640_254400# diff_168360_284280# GND efet w=2160 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1300 diff_179520_287640# GND GND GND efet w=2100 l=1140
+ ad=849600 pd=5280 as=0 ps=0 
M1301 diff_117960_263280# diff_179280_254400# diff_179520_287640# GND efet w=2160 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1302 diff_155400_282840# diff_153840_254520# diff_117960_263280# GND efet w=480 l=960
+ ad=345600 pd=2400 as=0 ps=0 
M1303 diff_117960_280920# diff_151440_254520# diff_150240_278280# GND efet w=480 l=900
+ ad=0 pd=0 as=288000 ps=2160 
M1304 diff_155400_281400# diff_153840_254520# diff_117960_280920# GND efet w=480 l=960
+ ad=345600 pd=2400 as=0 ps=0 
M1305 diff_145920_280320# diff_144240_281400# GND GND efet w=2040 l=1080
+ ad=1.1088e+06 pd=6000 as=0 ps=0 
M1306 GND diff_139080_277080# diff_138480_276960# GND efet w=1980 l=1140
+ ad=0 pd=0 as=1.1232e+06 ps=5280 
M1307 GND diff_117960_263280# diff_117960_263280# GND efet w=4440 l=1440
+ ad=0 pd=0 as=0 ps=0 
M1308 diff_138480_276960# diff_117960_263280# diff_117960_263280# GND efet w=2100 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1309 diff_117960_263280# diff_117960_263280# diff_145920_280320# GND efet w=2340 l=960
+ ad=0 pd=0 as=0 ps=0 
M1310 diff_149640_278400# diff_117960_263280# diff_117960_263280# GND efet w=2160 l=960
+ ad=1.2096e+06 pd=5520 as=0 ps=0 
M1311 GND diff_150240_278280# diff_149640_278400# GND efet w=1920 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1312 diff_117960_263280# diff_117960_263280# diff_161400_286080# GND efet w=480 l=1080
+ ad=0 pd=0 as=302400 ps=2400 
M1313 diff_171960_285840# diff_117960_263280# diff_117960_263280# GND efet w=1680 l=1320
+ ad=1.1952e+06 pd=5520 as=0 ps=0 
M1314 GND diff_172680_282840# diff_171960_285840# GND efet w=1740 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1315 GND diff_171480_208680# diff_117960_263280# GND efet w=960 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1316 GND GND diff_117840_290880# GND efet w=720 l=2760
+ ad=0 pd=0 as=0 ps=0 
M1317 GND GND diff_117960_263280# GND efet w=720 l=2760
+ ad=0 pd=0 as=0 ps=0 
M1318 GND diff_171480_208680# diff_117960_263280# GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M1319 diff_179520_284280# diff_177840_282840# GND GND efet w=2160 l=1080
+ ad=907200 pd=5280 as=0 ps=0 
M1320 diff_166560_282840# diff_117960_263280# diff_117960_263280# GND efet w=480 l=960
+ ad=345600 pd=2400 as=0 ps=0 
M1321 diff_117960_280920# diff_117960_263280# diff_161400_278280# GND efet w=480 l=1200
+ ad=0 pd=0 as=288000 ps=2160 
M1322 diff_117960_263280# diff_117960_263280# GND GND efet w=5160 l=960
+ ad=0 pd=0 as=0 ps=0 
M1323 diff_117960_263280# diff_117960_263280# GND GND efet w=660 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1324 diff_146040_275520# diff_144240_273960# GND GND efet w=1920 l=1080
+ ad=1.1376e+06 pd=5280 as=0 ps=0 
M1325 diff_117960_263280# diff_117960_263280# diff_146040_275520# GND efet w=2100 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1326 diff_149640_276960# diff_117960_263280# diff_117960_263280# GND efet w=2040 l=960
+ ad=1.1376e+06 pd=5280 as=0 ps=0 
M1327 GND diff_150240_277080# diff_149640_276960# GND efet w=1920 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1328 diff_157200_278880# diff_155400_281400# GND GND efet w=1980 l=1140
+ ad=1.0368e+06 pd=5760 as=0 ps=0 
M1329 diff_117960_263280# diff_117960_263280# diff_157200_278880# GND efet w=2220 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1330 diff_160800_278400# diff_117960_263280# diff_117960_263280# GND efet w=1800 l=1320
+ ad=1.2528e+06 pd=5520 as=0 ps=0 
M1331 GND diff_161400_278280# diff_160800_278400# GND efet w=1920 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1332 diff_166560_281400# diff_117960_263280# diff_117960_280920# GND efet w=600 l=1080
+ ad=345600 pd=2640 as=0 ps=0 
M1333 diff_117960_263280# diff_174360_263520# diff_172680_282840# GND efet w=480 l=1080
+ ad=0 pd=0 as=288000 ps=2160 
M1334 diff_117960_263280# diff_179280_254400# diff_179520_284280# GND efet w=2160 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1335 diff_177840_282840# diff_117960_263280# diff_117960_263280# GND efet w=540 l=1140
+ ad=288000 pd=2160 as=0 ps=0 
M1336 diff_117960_280920# diff_174360_263520# diff_172680_278280# GND efet w=600 l=1080
+ ad=0 pd=0 as=360000 ps=2400 
M1337 diff_168360_278880# diff_166560_281400# GND GND efet w=1920 l=1140
+ ad=936000 pd=5520 as=0 ps=0 
M1338 diff_117960_263280# diff_167640_254400# diff_168360_278880# GND efet w=2100 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1339 diff_171960_278400# diff_117960_263280# diff_117960_263280# GND efet w=1680 l=1380
+ ad=1.224e+06 pd=5520 as=0 ps=0 
M1340 GND diff_172680_278280# diff_171960_278400# GND efet w=1680 l=960
+ ad=0 pd=0 as=0 ps=0 
M1341 diff_157200_275520# diff_155400_274320# GND GND efet w=1920 l=1200
+ ad=1.1088e+06 pd=5280 as=0 ps=0 
M1342 diff_117960_263280# diff_139680_254520# diff_139080_277080# GND efet w=480 l=1020
+ ad=0 pd=0 as=259200 ps=2400 
M1343 diff_144240_273960# diff_142200_254520# diff_117960_263280# GND efet w=540 l=1020
+ ad=374400 pd=2880 as=0 ps=0 
M1344 diff_117960_263280# diff_139680_254520# diff_139080_269520# GND efet w=660 l=900
+ ad=0 pd=0 as=316800 ps=2640 
M1345 diff_144240_272520# diff_142200_254520# diff_117960_263280# GND efet w=480 l=960
+ ad=345600 pd=2400 as=0 ps=0 
M1346 diff_138480_269640# diff_117960_263280# diff_117960_263280# GND efet w=2040 l=960
+ ad=1.1232e+06 pd=5280 as=0 ps=0 
M1347 GND diff_139080_269520# diff_138480_269640# GND efet w=1920 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1348 diff_117960_263280# diff_117960_263280# diff_157200_275520# GND efet w=2040 l=960
+ ad=0 pd=0 as=0 ps=0 
M1349 diff_160800_276960# diff_117960_263280# diff_117960_263280# GND efet w=1680 l=1320
+ ad=1.152e+06 pd=5280 as=0 ps=0 
M1350 GND diff_161400_277200# diff_160800_276960# GND efet w=1980 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1351 diff_177840_281280# diff_117960_263280# diff_117960_280920# GND efet w=660 l=1260
+ ad=374400 pd=2640 as=0 ps=0 
M1352 diff_179520_278760# diff_177840_281280# GND GND efet w=2280 l=1200
+ ad=864000 pd=5280 as=0 ps=0 
M1353 diff_168360_275520# diff_166680_273960# GND GND efet w=1920 l=1200
+ ad=1.0512e+06 pd=5280 as=0 ps=0 
M1354 diff_117960_263280# diff_151440_254520# diff_150240_277080# GND efet w=480 l=1080
+ ad=0 pd=0 as=302400 ps=2400 
M1355 diff_155400_274320# diff_153840_254520# diff_117960_263280# GND efet w=600 l=900
+ ad=302400 pd=2400 as=0 ps=0 
M1356 diff_117960_263280# diff_151440_254520# diff_150360_269400# GND efet w=480 l=960
+ ad=0 pd=0 as=345600 ps=2400 
M1357 GND diff_139080_268320# diff_138480_268200# GND efet w=1980 l=1140
+ ad=0 pd=0 as=1.1088e+06 ps=5280 
M1358 GND GND diff_54240_263880# GND efet w=480 l=2520
+ ad=0 pd=0 as=0 ps=0 
M1359 GND diff_86760_205920# diff_51480_235440# GND efet w=900 l=960
+ ad=0 pd=0 as=0 ps=0 
M1360 diff_109920_264000# diff_26520_220920# GND GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M1361 GND GND diff_117960_263280# GND efet w=3840 l=960
+ ad=0 pd=0 as=0 ps=0 
M1362 diff_117960_263280# diff_117960_263280# GND GND efet w=3300 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1363 diff_93960_257880# diff_92160_256320# GND GND efet w=1980 l=1260
+ ad=1.1808e+06 pd=5520 as=0 ps=0 
M1364 diff_81000_256320# diff_78120_238200# diff_50160_238320# GND efet w=480 l=960
+ ad=360000 pd=2640 as=0 ps=0 
M1365 diff_51480_235440# diff_51480_235440# diff_93960_257880# GND efet w=1680 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1366 diff_50160_238320# diff_50160_238320# diff_87000_259560# GND efet w=480 l=840
+ ad=0 pd=0 as=374400 ps=2640 
M1367 diff_92160_256320# diff_51480_235440# diff_50160_238320# GND efet w=480 l=840
+ ad=360000 pd=2640 as=0 ps=0 
M1368 diff_50160_238320# diff_75720_237120# diff_75840_251880# GND efet w=480 l=960
+ ad=0 pd=0 as=345600 ps=2400 
M1369 diff_75120_251880# diff_73440_237000# diff_51480_235440# GND efet w=2280 l=900
+ ad=1.2384e+06 pd=5760 as=0 ps=0 
M1370 GND diff_75840_251880# diff_75120_251880# GND efet w=1980 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1371 diff_81000_254880# diff_78120_238200# diff_50160_238320# GND efet w=480 l=960
+ ad=345600 pd=2400 as=0 ps=0 
M1372 diff_82680_252360# diff_81000_254880# GND GND efet w=1980 l=1140
+ ad=1.224e+06 pd=5760 as=0 ps=0 
M1373 diff_50160_238320# diff_50160_238320# diff_87000_251880# GND efet w=480 l=840
+ ad=0 pd=0 as=345600 ps=2400 
M1374 GND diff_51480_235440# diff_54240_245520# GND efet w=5640 l=960
+ ad=0 pd=0 as=1.35072e+07 ps=39360 
M1375 GND diff_75840_250680# diff_75120_250560# GND efet w=2040 l=1200
+ ad=0 pd=0 as=1.152e+06 ps=5520 
M1376 diff_42000_244200# diff_60240_235200# diff_51480_235440# GND efet w=1200 l=960
+ ad=0 pd=0 as=0 ps=0 
M1377 GND diff_52080_238440# diff_54240_245520# GND efet w=3600 l=960
+ ad=0 pd=0 as=0 ps=0 
M1378 diff_51960_227760# diff_51960_227760# GND GND efet w=3600 l=1320
+ ad=0 pd=0 as=0 ps=0 
M1379 GND GND diff_28320_238920# GND efet w=600 l=960
+ ad=0 pd=0 as=0 ps=0 
M1380 diff_40440_238080# diff_28320_238920# GND GND efet w=2400 l=960
+ ad=3.9168e+06 pd=13440 as=0 ps=0 
M1381 diff_75120_250560# diff_73440_237000# diff_51480_235440# GND efet w=2160 l=960
+ ad=0 pd=0 as=0 ps=0 
M1382 diff_51480_235440# diff_51480_235440# diff_82680_252360# GND efet w=2100 l=900
+ ad=0 pd=0 as=0 ps=0 
M1383 diff_86400_251880# diff_85440_237000# diff_51480_235440# GND efet w=2160 l=960
+ ad=1.1952e+06 pd=6000 as=0 ps=0 
M1384 GND diff_87000_251880# diff_86400_251880# GND efet w=1980 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1385 diff_92160_254880# diff_51480_235440# diff_50160_238320# GND efet w=480 l=900
+ ad=345600 pd=2400 as=0 ps=0 
M1386 diff_93960_252240# diff_92160_254880# GND GND efet w=1860 l=1260
+ ad=1.1664e+06 pd=5280 as=0 ps=0 
M1387 diff_82800_249000# diff_81000_247440# GND GND efet w=1800 l=1200
+ ad=1.1232e+06 pd=5280 as=0 ps=0 
M1388 diff_51480_235440# diff_51480_235440# diff_82800_249000# GND efet w=1980 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1389 GND diff_51480_235440# diff_51960_227760# GND efet w=5700 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1390 diff_51480_235440# diff_64920_237000# diff_42000_244200# GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M1391 diff_54240_245520# diff_75720_237120# diff_75840_250680# GND efet w=540 l=1140
+ ad=0 pd=0 as=360000 ps=2640 
M1392 diff_86400_250320# diff_85440_237000# diff_51480_235440# GND efet w=2040 l=960
+ ad=1.1088e+06 pd=5520 as=0 ps=0 
M1393 GND diff_87000_250680# diff_86400_250320# GND efet w=1920 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1394 diff_51480_235440# diff_51480_235440# diff_93960_252240# GND efet w=1680 l=1320
+ ad=0 pd=0 as=0 ps=0 
M1395 GND diff_86760_205920# diff_51480_235440# GND efet w=720 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1396 diff_117960_263280# diff_117960_263280# diff_109920_264000# GND efet w=720 l=1320
+ ad=0 pd=0 as=0 ps=0 
M1397 diff_109920_264000# diff_123240_258000# diff_117960_263280# GND efet w=1260 l=840
+ ad=0 pd=0 as=0 ps=0 
M1398 GND diff_117960_263280# diff_117960_263280# GND efet w=4920 l=960
+ ad=0 pd=0 as=0 ps=0 
M1399 diff_138480_268200# diff_117960_263280# diff_117960_263280# GND efet w=2040 l=960
+ ad=0 pd=0 as=0 ps=0 
M1400 diff_146040_270000# diff_144240_272520# GND GND efet w=1980 l=1140
+ ad=1.1376e+06 pd=5280 as=0 ps=0 
M1401 diff_117960_263280# diff_117960_263280# diff_146040_270000# GND efet w=1740 l=1260
+ ad=0 pd=0 as=0 ps=0 
M1402 diff_149640_269640# diff_117960_263280# diff_117960_263280# GND efet w=2040 l=1080
+ ad=1.224e+06 pd=5760 as=0 ps=0 
M1403 GND diff_150360_269400# diff_149640_269640# GND efet w=2100 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1404 diff_146040_266640# diff_144240_265200# GND GND efet w=1920 l=1080
+ ad=1.1664e+06 pd=5280 as=0 ps=0 
M1405 diff_155520_272520# diff_153840_254520# diff_117960_263280# GND efet w=480 l=960
+ ad=302400 pd=2400 as=0 ps=0 
M1406 diff_117960_263280# diff_167640_254400# diff_168360_275520# GND efet w=2100 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1407 diff_171960_276960# diff_117960_263280# diff_117960_263280# GND efet w=1860 l=1380
+ ad=1.224e+06 pd=5760 as=0 ps=0 
M1408 GND diff_172680_273960# diff_171960_276960# GND efet w=1680 l=960
+ ad=0 pd=0 as=0 ps=0 
M1409 diff_117960_263280# diff_117960_263280# diff_161400_277200# GND efet w=480 l=960
+ ad=0 pd=0 as=345600 ps=2400 
M1410 diff_166680_273960# diff_117960_263280# diff_117960_263280# GND efet w=540 l=1080
+ ad=288000 pd=2160 as=0 ps=0 
M1411 diff_117960_263280# diff_179280_254400# diff_179520_278760# GND efet w=2100 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1412 GND diff_171480_208680# diff_117960_263280# GND efet w=960 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1413 GND GND diff_117960_263280# GND efet w=600 l=3120
+ ad=0 pd=0 as=0 ps=0 
M1414 GND GND diff_117960_280920# GND efet w=660 l=2940
+ ad=0 pd=0 as=0 ps=0 
M1415 GND diff_171480_208680# diff_117960_263280# GND efet w=1020 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1416 diff_179520_275400# diff_177840_273960# GND GND efet w=2280 l=1200
+ ad=936000 pd=5520 as=0 ps=0 
M1417 diff_117960_263280# diff_179280_254400# diff_179520_275400# GND efet w=2160 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1418 diff_117960_263280# diff_117960_263280# diff_161400_269520# GND efet w=480 l=960
+ ad=0 pd=0 as=345600 ps=2400 
M1419 diff_117960_263280# diff_117960_263280# GND GND efet w=4920 l=960
+ ad=0 pd=0 as=0 ps=0 
M1420 diff_117960_263280# diff_117960_263280# diff_146040_266640# GND efet w=1740 l=1260
+ ad=0 pd=0 as=0 ps=0 
M1421 diff_149640_268200# diff_117960_263280# diff_117960_263280# GND efet w=2040 l=960
+ ad=1.152e+06 pd=5520 as=0 ps=0 
M1422 GND diff_150240_268320# diff_149640_268200# GND efet w=2220 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1423 diff_157200_270000# diff_155520_272520# GND GND efet w=1980 l=1260
+ ad=1.1808e+06 pd=5760 as=0 ps=0 
M1424 diff_117960_263280# diff_117960_263280# diff_157200_270000# GND efet w=2340 l=900
+ ad=0 pd=0 as=0 ps=0 
M1425 diff_160800_269520# diff_117960_263280# diff_117960_263280# GND efet w=2400 l=960
+ ad=1.224e+06 pd=6240 as=0 ps=0 
M1426 GND diff_161400_269520# diff_160800_269520# GND efet w=2100 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1427 diff_166680_272520# diff_117960_263280# diff_117960_263280# GND efet w=480 l=960
+ ad=302400 pd=2400 as=0 ps=0 
M1428 diff_117960_263280# diff_174360_263520# diff_172680_273960# GND efet w=480 l=1020
+ ad=0 pd=0 as=288000 ps=2160 
M1429 diff_177840_273960# diff_117960_263280# diff_117960_263280# GND efet w=300 l=1380
+ ad=288000 pd=2160 as=0 ps=0 
M1430 diff_117960_263280# diff_174360_263520# diff_172680_269400# GND efet w=540 l=1140
+ ad=0 pd=0 as=316800 ps=2400 
M1431 diff_177840_272520# diff_117960_263280# diff_117960_263280# GND efet w=300 l=1500
+ ad=302400 pd=2400 as=0 ps=0 
M1432 diff_168360_270000# diff_166680_272520# GND GND efet w=2040 l=1080
+ ad=1.0944e+06 pd=5520 as=0 ps=0 
M1433 diff_117960_263280# diff_167640_254400# diff_168360_270000# GND efet w=2220 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1434 diff_171960_269520# diff_117960_263280# diff_117960_263280# GND efet w=2160 l=1200
+ ad=1.0944e+06 pd=5760 as=0 ps=0 
M1435 diff_157200_266640# diff_155520_265080# GND GND efet w=1920 l=1140
+ ad=1.152e+06 pd=5520 as=0 ps=0 
M1436 diff_117960_263280# diff_139680_254520# diff_139080_268320# GND efet w=540 l=1140
+ ad=0 pd=0 as=388800 ps=3120 
M1437 diff_144240_265200# diff_142200_254520# diff_117960_263280# GND efet w=360 l=1020
+ ad=259200 pd=2160 as=0 ps=0 
M1438 diff_117960_263280# diff_139680_254520# diff_139080_260640# GND efet w=600 l=960
+ ad=0 pd=0 as=316800 ps=2640 
M1439 diff_144240_263640# diff_142200_254520# diff_117960_263280# GND efet w=480 l=960
+ ad=345600 pd=2400 as=0 ps=0 
M1440 diff_138480_260760# diff_117960_263280# diff_117960_263280# GND efet w=2040 l=1140
+ ad=1.1088e+06 pd=5280 as=0 ps=0 
M1441 GND diff_139080_260640# diff_138480_260760# GND efet w=1920 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1442 diff_117960_263280# diff_151440_254520# diff_150240_268320# GND efet w=600 l=960
+ ad=0 pd=0 as=417600 ps=2640 
M1443 diff_117960_263280# diff_117960_263280# diff_157200_266640# GND efet w=2220 l=960
+ ad=0 pd=0 as=0 ps=0 
M1444 diff_160800_268080# diff_117960_263280# diff_117960_263280# GND efet w=2040 l=1200
+ ad=1.0512e+06 pd=5760 as=0 ps=0 
M1445 GND diff_161520_265080# diff_160800_268080# GND efet w=2160 l=1320
+ ad=0 pd=0 as=0 ps=0 
M1446 GND diff_172680_269400# diff_171960_269520# GND efet w=1740 l=1260
+ ad=0 pd=0 as=0 ps=0 
M1447 diff_168360_266520# diff_166680_265080# GND GND efet w=2040 l=1200
+ ad=1.1232e+06 pd=5520 as=0 ps=0 
M1448 diff_155520_265080# diff_153840_254520# diff_117960_263280# GND efet w=540 l=1140
+ ad=302400 pd=2400 as=0 ps=0 
M1449 diff_117960_263280# diff_151440_254520# diff_150360_260520# GND efet w=480 l=960
+ ad=0 pd=0 as=345600 ps=2400 
M1450 GND GND diff_50160_238320# GND efet w=480 l=2520
+ ad=0 pd=0 as=0 ps=0 
M1451 GND diff_110040_234240# diff_109800_255840# GND efet w=1080 l=1080
+ ad=0 pd=0 as=3.8016e+06 ps=14880 
M1452 diff_109800_255840# GND GND GND efet w=720 l=5400
+ ad=0 pd=0 as=0 ps=0 
M1453 diff_110040_234240# diff_109800_255840# GND GND efet w=960 l=960
+ ad=9.2592e+06 pd=29280 as=0 ps=0 
M1454 diff_146040_261120# diff_144240_263640# GND GND efet w=1980 l=1140
+ ad=1.2096e+06 pd=5760 as=0 ps=0 
M1455 diff_117960_263280# diff_117960_263280# diff_146040_261120# GND efet w=2040 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1456 diff_149640_260640# diff_117960_263280# diff_117960_263280# GND efet w=2160 l=1200
+ ad=1.2672e+06 pd=5760 as=0 ps=0 
M1457 GND diff_150360_260520# diff_149640_260640# GND efet w=2280 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1458 diff_155520_263640# diff_153840_254520# diff_117960_263280# GND efet w=480 l=960
+ ad=302400 pd=2400 as=0 ps=0 
M1459 diff_117960_263280# diff_167640_254400# diff_168360_266520# GND efet w=2160 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1460 diff_171960_268200# diff_117960_263280# diff_117960_263280# GND efet w=2280 l=1440
+ ad=1.0656e+06 pd=5520 as=0 ps=0 
M1461 GND diff_172560_268320# diff_171960_268200# GND efet w=1860 l=1440
+ ad=0 pd=0 as=0 ps=0 
M1462 diff_179520_270000# diff_177840_272520# GND GND efet w=2460 l=1260
+ ad=864000 pd=5760 as=0 ps=0 
M1463 diff_117960_263280# diff_179280_254400# diff_179520_270000# GND efet w=2280 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1464 GND diff_171480_208680# diff_117960_263280# GND efet w=1200 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1465 GND GND diff_117960_263280# GND efet w=720 l=2820
+ ad=0 pd=0 as=0 ps=0 
M1466 GND GND diff_117960_263280# GND efet w=660 l=2700
+ ad=0 pd=0 as=0 ps=0 
M1467 GND diff_171480_208680# diff_117960_263280# GND efet w=960 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1468 diff_179520_266520# diff_177840_265080# GND GND efet w=2400 l=1080
+ ad=1.08e+06 pd=6240 as=0 ps=0 
M1469 diff_117960_263280# diff_179280_254400# diff_179520_266520# GND efet w=2400 l=960
+ ad=0 pd=0 as=0 ps=0 
M1470 diff_117960_263280# diff_117960_263280# diff_161520_265080# GND efet w=480 l=960
+ ad=0 pd=0 as=331200 ps=2400 
M1471 diff_166680_265080# diff_117960_263280# diff_117960_263280# GND efet w=420 l=1200
+ ad=288000 pd=2160 as=0 ps=0 
M1472 diff_117960_263280# diff_117960_263280# diff_161520_260520# GND efet w=480 l=960
+ ad=0 pd=0 as=331200 ps=2400 
M1473 diff_157200_261120# diff_155520_263640# GND GND efet w=1980 l=1140
+ ad=1.224e+06 pd=5760 as=0 ps=0 
M1474 diff_117960_263280# diff_117960_263280# diff_157200_261120# GND efet w=2280 l=960
+ ad=0 pd=0 as=0 ps=0 
M1475 diff_160800_260640# diff_117960_263280# diff_117960_263280# GND efet w=2280 l=960
+ ad=1.2096e+06 pd=6000 as=0 ps=0 
M1476 GND diff_161520_260520# diff_160800_260640# GND efet w=2100 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1477 diff_166680_263640# diff_117960_263280# diff_117960_263280# GND efet w=480 l=960
+ ad=302400 pd=2400 as=0 ps=0 
M1478 diff_168360_261840# diff_166680_263640# GND GND efet w=2220 l=1200
+ ad=1.008e+06 pd=5760 as=0 ps=0 
M1479 diff_117960_263280# diff_174360_263520# diff_172560_268320# GND efet w=480 l=960
+ ad=0 pd=0 as=302400 ps=2400 
M1480 GND diff_171480_208680# diff_117960_263280# GND efet w=960 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1481 diff_177840_265080# diff_117960_263280# diff_117960_263280# GND efet w=300 l=1260
+ ad=288000 pd=2160 as=0 ps=0 
M1482 diff_117960_263280# diff_174360_263520# diff_172680_260520# GND efet w=480 l=1080
+ ad=0 pd=0 as=331200 ps=2640 
M1483 diff_177840_263520# diff_117960_263280# diff_117960_263280# GND efet w=360 l=1440
+ ad=360000 pd=2640 as=0 ps=0 
M1484 diff_117960_263280# diff_167640_254400# diff_168360_261840# GND efet w=2160 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1485 diff_172080_260640# diff_117960_263280# diff_117960_263280# GND efet w=2160 l=1080
+ ad=1.0944e+06 pd=5760 as=0 ps=0 
M1486 GND diff_172680_260520# diff_172080_260640# GND efet w=2280 l=1320
+ ad=0 pd=0 as=0 ps=0 
M1487 GND GND diff_117960_263280# GND efet w=720 l=2820
+ ad=0 pd=0 as=0 ps=0 
M1488 GND GND GND GND efet w=9780 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1489 GND GND GND GND efet w=8940 l=1500
+ ad=0 pd=0 as=0 ps=0 
M1490 GND GND diff_117960_263280# GND efet w=720 l=2820
+ ad=0 pd=0 as=0 ps=0 
M1491 diff_179520_261120# diff_177840_263520# GND GND efet w=2160 l=1320
+ ad=950400 pd=5280 as=0 ps=0 
M1492 diff_117960_263280# diff_179280_254400# diff_179520_261120# GND efet w=2220 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1493 GND diff_171480_208680# diff_117960_263280# GND efet w=960 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1494 GND GND diff_50160_238320# GND efet w=480 l=2400
+ ad=0 pd=0 as=0 ps=0 
M1495 GND GND diff_110040_234240# GND efet w=480 l=5400
+ ad=0 pd=0 as=0 ps=0 
M1496 diff_94080_217680# GND GND GND efet w=720 l=5520
+ ad=1.17216e+07 pd=40560 as=0 ps=0 
M1497 GND diff_110040_234240# diff_94080_217680# GND efet w=1260 l=900
+ ad=0 pd=0 as=0 ps=0 
M1498 diff_117120_254520# diff_109800_255840# GND GND efet w=1200 l=960
+ ad=3.6432e+06 pd=13440 as=0 ps=0 
M1499 GND diff_134880_253320# diff_117960_263280# GND efet w=1200 l=960
+ ad=0 pd=0 as=0 ps=0 
M1500 GND diff_134880_253320# diff_139680_254520# GND efet w=960 l=960
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M1501 GND diff_141600_255960# diff_142200_254520# GND efet w=960 l=960
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M1502 GND diff_141600_255960# diff_117960_263280# GND efet w=1200 l=960
+ ad=0 pd=0 as=0 ps=0 
M1503 GND GND diff_117120_254520# GND efet w=780 l=5460
+ ad=0 pd=0 as=0 ps=0 
M1504 GND diff_86760_205920# diff_51480_235440# GND efet w=780 l=900
+ ad=0 pd=0 as=0 ps=0 
M1505 diff_134880_253320# GND GND GND efet w=540 l=5100
+ ad=4.6944e+06 pd=18480 as=0 ps=0 
M1506 diff_117960_263280# diff_133560_235080# diff_133560_235080# GND efet w=1320 l=960
+ ad=0 pd=0 as=9.7776e+07 ps=313680 
M1507 diff_139680_254520# diff_133560_235080# diff_139680_251040# GND efet w=1140 l=1080
+ ad=0 pd=0 as=4.49424e+07 ps=111360 
M1508 diff_142200_254520# diff_133560_235080# diff_139680_251040# GND efet w=1020 l=900
+ ad=0 pd=0 as=0 ps=0 
M1509 diff_117960_263280# diff_133560_235080# diff_133560_235080# GND efet w=1320 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1510 diff_93960_249000# diff_92160_247440# GND GND efet w=1860 l=1500
+ ad=1.1232e+06 pd=5280 as=0 ps=0 
M1511 diff_94080_217680# diff_105120_208440# diff_110640_249960# GND efet w=720 l=840
+ ad=0 pd=0 as=475200 ps=2880 
M1512 diff_117120_254520# diff_105120_208440# diff_115080_246600# GND efet w=720 l=1080
+ ad=0 pd=0 as=518400 ps=2880 
M1513 diff_81000_247440# diff_78120_238200# diff_54240_245520# GND efet w=540 l=1020
+ ad=345600 pd=2400 as=0 ps=0 
M1514 diff_51960_227760# diff_75720_237120# diff_75840_243000# GND efet w=480 l=960
+ ad=0 pd=0 as=345600 ps=2400 
M1515 diff_75120_243120# diff_73440_237000# diff_51480_235440# GND efet w=2280 l=1080
+ ad=1.152e+06 pd=5520 as=0 ps=0 
M1516 GND GND diff_40440_238080# GND efet w=600 l=5400
+ ad=0 pd=0 as=0 ps=0 
M1517 GND diff_11280_215400# diff_35040_230160# GND efet w=2040 l=960
+ ad=0 pd=0 as=4.7808e+06 ps=13680 
M1518 diff_40440_238080# GND diff_39480_236280# GND efet w=1080 l=1200
+ ad=0 pd=0 as=576000 ps=4080 
M1519 GND GND GND GND efet w=33240 l=2280
+ ad=0 pd=0 as=0 ps=0 
M1520 GND GND GND GND efet w=46620 l=4560
+ ad=0 pd=0 as=0 ps=0 
M1521 diff_35040_230160# diff_21360_57480# GND GND efet w=2220 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1522 GND GND GND GND efet w=2460 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1523 GND GND diff_60240_235200# GND efet w=480 l=2280
+ ad=0 pd=0 as=4.0464e+06 ps=15840 
M1524 GND diff_21360_45480# diff_32040_231840# GND efet w=1080 l=1020
+ ad=0 pd=0 as=4.896e+06 ps=16560 
M1525 diff_40560_232800# diff_39480_236280# GND GND efet w=1680 l=960
+ ad=3.7872e+06 pd=10080 as=0 ps=0 
M1526 diff_51480_235440# GND GND GND efet w=600 l=2280
+ ad=0 pd=0 as=0 ps=0 
M1527 GND diff_44400_224400# diff_51480_235440# GND efet w=2400 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1528 GND GND diff_40560_232800# GND efet w=540 l=4260
+ ad=0 pd=0 as=0 ps=0 
M1529 diff_32040_231840# GND GND GND efet w=540 l=5580
+ ad=0 pd=0 as=0 ps=0 
M1530 diff_39480_231000# GND diff_40560_232800# GND efet w=720 l=960
+ ad=1.4688e+06 pd=6480 as=0 ps=0 
M1531 GND GND diff_51480_235440# GND efet w=2760 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1532 GND diff_75840_243000# diff_75120_243120# GND efet w=1980 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1533 diff_81000_246000# diff_78120_238200# diff_51960_227760# GND efet w=480 l=960
+ ad=345600 pd=2400 as=0 ps=0 
M1534 diff_51480_235440# diff_51480_235440# diff_93960_249000# GND efet w=1620 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1535 diff_54240_245520# diff_50160_238320# diff_87000_250680# GND efet w=540 l=900
+ ad=0 pd=0 as=388800 ps=2880 
M1536 diff_92160_247440# diff_51480_235440# diff_54240_245520# GND efet w=480 l=840
+ ad=345600 pd=2400 as=0 ps=0 
M1537 diff_51960_227760# diff_50160_238320# diff_87000_243000# GND efet w=480 l=840
+ ad=0 pd=0 as=345600 ps=2400 
M1538 diff_92160_246000# diff_51480_235440# diff_51960_227760# GND efet w=480 l=840
+ ad=345600 pd=2400 as=0 ps=0 
M1539 diff_82680_243840# diff_81000_246000# GND GND efet w=2160 l=1080
+ ad=1.2672e+06 pd=6240 as=0 ps=0 
M1540 diff_51480_235440# diff_51480_235440# diff_82680_243840# GND efet w=1920 l=1440
+ ad=0 pd=0 as=0 ps=0 
M1541 diff_86400_243000# diff_85440_237000# diff_51480_235440# GND efet w=2100 l=1020
+ ad=1.1808e+06 pd=6000 as=0 ps=0 
M1542 diff_64920_237000# GND GND GND efet w=660 l=2580
+ ad=5.976e+06 pd=15120 as=0 ps=0 
M1543 GND diff_87000_243000# diff_86400_243000# GND efet w=2100 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1544 diff_93960_243360# diff_92160_246000# GND GND efet w=1980 l=1260
+ ad=1.1952e+06 pd=5520 as=0 ps=0 
M1545 diff_51480_235440# diff_51480_235440# diff_93960_243360# GND efet w=1740 l=1620
+ ad=0 pd=0 as=0 ps=0 
M1546 GND diff_86760_205920# diff_51480_235440# GND efet w=720 l=960
+ ad=0 pd=0 as=0 ps=0 
M1547 diff_112200_247080# diff_110040_234240# diff_109800_255840# GND efet w=1800 l=1020
+ ad=1.5408e+06 pd=6720 as=0 ps=0 
M1548 GND GND diff_54240_245520# GND efet w=540 l=2700
+ ad=0 pd=0 as=0 ps=0 
M1549 GND diff_110640_249960# diff_112200_247080# GND efet w=2820 l=960
+ ad=0 pd=0 as=0 ps=0 
M1550 diff_116040_246960# diff_115080_246600# GND GND efet w=2880 l=960
+ ad=1.5696e+06 pd=6960 as=0 ps=0 
M1551 diff_110040_234240# diff_110040_234240# diff_116040_246960# GND efet w=1080 l=1560
+ ad=0 pd=0 as=0 ps=0 
M1552 GND GND diff_51960_227760# GND efet w=540 l=2580
+ ad=0 pd=0 as=0 ps=0 
M1553 GND diff_147480_249360# diff_117960_263280# GND efet w=1200 l=840
+ ad=0 pd=0 as=0 ps=0 
M1554 GND diff_147480_249360# diff_151440_254520# GND efet w=960 l=840
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M1555 GND diff_117960_263280# diff_153840_254520# GND efet w=1080 l=840
+ ad=0 pd=0 as=1.4256e+06 ps=4800 
M1556 GND diff_117960_263280# diff_117960_263280# GND efet w=1260 l=900
+ ad=0 pd=0 as=0 ps=0 
M1557 GND diff_117960_263280# diff_117960_263280# GND efet w=840 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1558 diff_117960_263280# diff_133560_235080# diff_133560_235080# GND efet w=1140 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1559 diff_151440_254520# diff_133560_235080# diff_139680_251040# GND efet w=1020 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1560 diff_153840_254520# diff_133560_235080# diff_139680_251040# GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M1561 diff_117960_263280# diff_133560_235080# diff_133560_235080# GND efet w=1200 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1562 GND diff_133560_235080# diff_134880_253320# GND efet w=960 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1563 diff_141600_255960# diff_133560_235080# GND GND efet w=840 l=960
+ ad=2.9232e+06 pd=10080 as=0 ps=0 
M1564 GND diff_133560_235080# diff_147480_249360# GND efet w=900 l=1020
+ ad=0 pd=0 as=3.024e+06 ps=10080 
M1565 diff_117960_263280# diff_133560_235080# GND GND efet w=840 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1566 GND diff_117960_263280# diff_117960_263280# GND efet w=660 l=1320
+ ad=0 pd=0 as=0 ps=0 
M1567 GND diff_117960_263280# diff_117960_263280# GND efet w=900 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1568 GND diff_117960_263280# diff_167640_254400# GND efet w=1080 l=1020
+ ad=0 pd=0 as=1.4256e+06 ps=4800 
M1569 diff_117960_263280# diff_156720_230520# diff_133560_235080# GND efet w=1200 l=900
+ ad=0 pd=0 as=0 ps=0 
M1570 diff_139680_251040# diff_156720_230520# diff_117960_263280# GND efet w=1020 l=900
+ ad=0 pd=0 as=0 ps=0 
M1571 diff_117960_263280# diff_161160_232920# diff_139680_251040# GND efet w=1020 l=900
+ ad=0 pd=0 as=0 ps=0 
M1572 diff_167640_254400# diff_161160_232920# diff_133560_235080# GND efet w=1080 l=840
+ ad=0 pd=0 as=0 ps=0 
M1573 GND diff_156720_230520# diff_117960_263280# GND efet w=1020 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1574 GND diff_128520_245400# GND GND efet w=6420 l=540
+ ad=0 pd=0 as=0 ps=0 
M1575 GND diff_128520_245400# GND GND efet w=840 l=1920
+ ad=0 pd=0 as=0 ps=0 
M1576 diff_128520_245400# GND GND GND efet w=540 l=1140
+ ad=230400 pd=1920 as=0 ps=0 
M1577 GND diff_86760_205920# diff_51480_235440# GND efet w=840 l=960
+ ad=0 pd=0 as=0 ps=0 
M1578 diff_110040_234240# GND GND GND efet w=540 l=5940
+ ad=0 pd=0 as=0 ps=0 
M1579 GND diff_105120_208440# diff_110040_234240# GND efet w=960 l=960
+ ad=0 pd=0 as=0 ps=0 
M1580 diff_105120_208440# diff_110040_234240# GND GND efet w=1080 l=960
+ ad=9.4896e+06 pd=29520 as=0 ps=0 
M1581 diff_141600_255960# GND GND GND efet w=540 l=3780
+ ad=0 pd=0 as=0 ps=0 
M1582 GND GND diff_147480_249360# GND efet w=540 l=4380
+ ad=0 pd=0 as=0 ps=0 
M1583 diff_117960_263280# diff_161160_232920# GND GND efet w=960 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1584 GND diff_117960_263280# diff_117960_263280# GND efet w=840 l=1320
+ ad=0 pd=0 as=0 ps=0 
M1585 GND diff_117960_263280# diff_174360_263520# GND efet w=960 l=960
+ ad=0 pd=0 as=1.2672e+06 ps=4560 
M1586 GND diff_176640_255840# diff_117960_263280# GND efet w=960 l=960
+ ad=0 pd=0 as=0 ps=0 
M1587 GND diff_176640_255840# diff_179280_254400# GND efet w=1200 l=960
+ ad=0 pd=0 as=1.5408e+06 ps=5280 
M1588 diff_117960_263280# diff_165720_226080# diff_133560_235080# GND efet w=1260 l=900
+ ad=0 pd=0 as=0 ps=0 
M1589 diff_174360_263520# diff_165720_226080# diff_139680_251040# GND efet w=1020 l=900
+ ad=0 pd=0 as=0 ps=0 
M1590 diff_117960_263280# diff_133560_235080# diff_139680_251040# GND efet w=1020 l=900
+ ad=0 pd=0 as=0 ps=0 
M1591 diff_179280_254400# diff_133560_235080# diff_133560_235080# GND efet w=840 l=1320
+ ad=0 pd=0 as=0 ps=0 
M1592 diff_117960_263280# GND GND GND efet w=480 l=3960
+ ad=0 pd=0 as=0 ps=0 
M1593 GND GND diff_117960_263280# GND efet w=540 l=4380
+ ad=0 pd=0 as=0 ps=0 
M1594 GND diff_165720_226080# diff_117960_263280# GND efet w=840 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1595 diff_176640_255840# diff_133560_235080# GND GND efet w=840 l=1080
+ ad=2.6928e+06 pd=9600 as=0 ps=0 
M1596 GND GND GND GND efet w=1080 l=3780
+ ad=0 pd=0 as=0 ps=0 
M1597 diff_117960_263280# GND GND GND efet w=540 l=4020
+ ad=0 pd=0 as=0 ps=0 
M1598 GND GND diff_117960_263280# GND efet w=480 l=3960
+ ad=0 pd=0 as=0 ps=0 
M1599 diff_176640_255840# GND GND GND efet w=480 l=3960
+ ad=0 pd=0 as=0 ps=0 
M1600 diff_133560_235080# diff_133560_235080# GND GND efet w=1860 l=1500
+ ad=0 pd=0 as=0 ps=0 
M1601 GND GND diff_133560_235080# GND efet w=600 l=2400
+ ad=0 pd=0 as=0 ps=0 
M1602 GND GND diff_105120_208440# GND efet w=540 l=5700
+ ad=0 pd=0 as=0 ps=0 
M1603 diff_94080_215520# GND GND GND efet w=780 l=6120
+ ad=1.14048e+07 pd=40080 as=0 ps=0 
M1604 GND diff_105120_208440# diff_94080_215520# GND efet w=1140 l=900
+ ad=0 pd=0 as=0 ps=0 
M1605 diff_117120_241680# diff_110040_234240# GND GND efet w=1080 l=960
+ ad=3.5856e+06 pd=13200 as=0 ps=0 
M1606 GND GND diff_117120_241680# GND efet w=720 l=5520
+ ad=0 pd=0 as=0 ps=0 
M1607 diff_128520_243360# GND GND GND efet w=540 l=1140
+ ad=273600 pd=2640 as=0 ps=0 
M1608 diff_117960_263280# diff_128520_243360# diff_117960_263280# GND efet w=4740 l=1260
+ ad=0 pd=0 as=0 ps=0 
M1609 diff_117960_263280# diff_128520_243360# GND GND efet w=600 l=1800
+ ad=0 pd=0 as=0 ps=0 
M1610 diff_60240_235200# GND GND GND efet w=2280 l=960
+ ad=0 pd=0 as=0 ps=0 
M1611 GND diff_41520_198840# diff_64920_237000# GND efet w=2400 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1612 GND diff_44400_224400# diff_60240_235200# GND efet w=2280 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1613 diff_64920_237000# diff_44400_224400# GND GND efet w=2460 l=900
+ ad=0 pd=0 as=0 ps=0 
M1614 GND diff_71760_233040# diff_73440_237000# GND efet w=1320 l=840
+ ad=0 pd=0 as=1.7424e+06 ps=5280 
M1615 GND diff_71760_233040# diff_75720_237120# GND efet w=960 l=840
+ ad=0 pd=0 as=1.2528e+06 ps=4560 
M1616 GND diff_77640_238440# diff_78120_238200# GND efet w=960 l=960
+ ad=0 pd=0 as=1.2816e+06 ps=4800 
M1617 GND diff_77640_238440# diff_51480_235440# GND efet w=1320 l=840
+ ad=0 pd=0 as=0 ps=0 
M1618 diff_73440_237000# diff_72840_236280# diff_63960_210840# GND efet w=1320 l=960
+ ad=0 pd=0 as=2.20896e+07 ps=74160 
M1619 diff_75720_237120# diff_72840_236280# diff_69480_207240# GND efet w=840 l=960
+ ad=0 pd=0 as=2.0808e+07 ps=51840 
M1620 diff_78120_238200# diff_77640_236160# diff_69480_207240# GND efet w=1020 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1621 diff_51480_235440# diff_77640_236160# diff_63960_210840# GND efet w=1320 l=960
+ ad=0 pd=0 as=0 ps=0 
M1622 GND GND GND GND efet w=780 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1623 diff_32040_231840# diff_34560_231000# diff_35040_230160# GND efet w=1920 l=840
+ ad=0 pd=0 as=0 ps=0 
M1624 GND diff_50160_238320# diff_85440_237000# GND efet w=1320 l=840
+ ad=0 pd=0 as=1.7424e+06 ps=5280 
M1625 diff_50160_238320# diff_50160_238320# GND GND efet w=780 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1626 GND diff_51480_235440# diff_51480_235440# GND efet w=660 l=1260
+ ad=0 pd=0 as=0 ps=0 
M1627 diff_51480_235440# diff_51480_235440# GND GND efet w=1260 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1628 diff_94080_215520# GND diff_110640_237120# GND efet w=600 l=960
+ ad=0 pd=0 as=374400 ps=2640 
M1629 diff_133560_235080# diff_133560_235080# GND GND efet w=1200 l=840
+ ad=0 pd=0 as=0 ps=0 
M1630 diff_133560_235080# diff_133560_235080# GND GND efet w=1200 l=960
+ ad=0 pd=0 as=0 ps=0 
M1631 diff_133560_235080# diff_133560_235080# GND GND efet w=1140 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1632 diff_156720_230520# GND GND GND efet w=1140 l=1140
+ ad=9.2304e+06 pd=30720 as=0 ps=0 
M1633 GND GND diff_133560_235080# GND efet w=2400 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1634 diff_161160_232920# GND GND GND efet w=1260 l=1020
+ ad=8.7696e+06 pd=30240 as=0 ps=0 
M1635 diff_165720_226080# GND GND GND efet w=1140 l=1140
+ ad=1.04832e+07 pd=36240 as=0 ps=0 
M1636 diff_133560_235080# GND GND GND efet w=1380 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1637 GND diff_183360_241080# GND GND efet w=4380 l=1260
+ ad=0 pd=0 as=0 ps=0 
M1638 diff_133560_235080# diff_138120_242040# GND GND efet w=2280 l=840
+ ad=0 pd=0 as=0 ps=0 
M1639 diff_133560_235080# diff_138120_242040# GND GND efet w=1200 l=900
+ ad=0 pd=0 as=0 ps=0 
M1640 GND diff_138120_242040# diff_156720_230520# GND efet w=1140 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1641 GND diff_138120_242040# diff_161160_232920# GND efet w=1140 l=900
+ ad=0 pd=0 as=0 ps=0 
M1642 diff_133560_235080# diff_148080_240000# GND GND efet w=1140 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1643 GND diff_133560_235080# diff_133560_235080# GND efet w=2040 l=1320
+ ad=0 pd=0 as=0 ps=0 
M1644 diff_133560_235080# diff_148080_240000# GND GND efet w=1140 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1645 diff_117120_241680# GND diff_115080_234840# GND efet w=600 l=1080
+ ad=0 pd=0 as=374400 ps=2640 
M1646 diff_165720_226080# diff_148080_240000# GND GND efet w=1080 l=840
+ ad=0 pd=0 as=0 ps=0 
M1647 diff_133560_235080# diff_148080_240000# GND GND efet w=1320 l=1320
+ ad=0 pd=0 as=0 ps=0 
M1648 GND GND diff_138120_242040# GND efet w=420 l=3540
+ ad=0 pd=0 as=3.9312e+06 ps=13680 
M1649 diff_133560_235080# diff_133560_235080# GND GND efet w=1080 l=1440
+ ad=0 pd=0 as=0 ps=0 
M1650 diff_85440_237000# diff_83160_218280# diff_63960_210840# GND efet w=1320 l=960
+ ad=0 pd=0 as=0 ps=0 
M1651 diff_50160_238320# diff_83160_218280# diff_69480_207240# GND efet w=900 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1652 diff_51480_235440# diff_63960_210840# diff_69480_207240# GND efet w=960 l=960
+ ad=0 pd=0 as=0 ps=0 
M1653 diff_51480_235440# diff_63960_210840# diff_63960_210840# GND efet w=1320 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1654 GND diff_110640_237120# diff_112200_234120# GND efet w=3360 l=960
+ ad=0 pd=0 as=1.5696e+06 ps=7440 
M1655 GND diff_72840_236280# diff_71760_233040# GND efet w=1020 l=1020
+ ad=0 pd=0 as=3.4416e+06 ps=12000 
M1656 diff_77640_238440# diff_77640_236160# GND GND efet w=960 l=960
+ ad=1.9296e+06 pd=6240 as=0 ps=0 
M1657 diff_112200_234120# diff_105120_208440# diff_110040_234240# GND efet w=1800 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1658 diff_116040_234240# diff_115080_234840# GND GND efet w=3180 l=1020
+ ad=1.5552e+06 pd=7200 as=0 ps=0 
M1659 GND diff_133560_235080# diff_156720_230520# GND efet w=1200 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1660 GND diff_133560_235080# diff_165720_226080# GND efet w=1080 l=840
+ ad=0 pd=0 as=0 ps=0 
M1661 diff_138120_242040# diff_148080_240000# GND GND efet w=2160 l=960
+ ad=0 pd=0 as=0 ps=0 
M1662 diff_148080_240000# diff_164160_221520# GND GND efet w=4320 l=1080
+ ad=4.536e+06 pd=15120 as=0 ps=0 
M1663 diff_105120_208440# diff_105120_208440# diff_116040_234240# GND efet w=960 l=1740
+ ad=0 pd=0 as=0 ps=0 
M1664 diff_133560_235080# GND diff_133560_235080# GND efet w=3420 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1665 diff_133560_235080# GND GND GND efet w=720 l=3360
+ ad=0 pd=0 as=0 ps=0 
M1666 GND GND diff_133560_235080# GND efet w=1620 l=1740
+ ad=0 pd=0 as=0 ps=0 
M1667 GND GND diff_51480_235440# GND efet w=480 l=5040
+ ad=0 pd=0 as=0 ps=0 
M1668 GND diff_83160_218280# diff_50160_238320# GND efet w=960 l=900
+ ad=0 pd=0 as=0 ps=0 
M1669 diff_51480_235440# diff_63960_210840# GND GND efet w=960 l=960
+ ad=0 pd=0 as=0 ps=0 
M1670 diff_34560_231000# diff_39480_231000# GND GND efet w=1620 l=1020
+ ad=2.2176e+06 pd=7680 as=0 ps=0 
M1671 GND GND diff_34560_231000# GND efet w=720 l=5400
+ ad=0 pd=0 as=0 ps=0 
M1672 GND diff_32040_231840# GND GND efet w=1140 l=960
+ ad=0 pd=0 as=0 ps=0 
M1673 GND diff_58200_222720# diff_50160_238320# GND efet w=3600 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1674 diff_51960_227760# GND GND GND efet w=660 l=1920
+ ad=0 pd=0 as=0 ps=0 
M1675 diff_44400_224400# GND GND GND efet w=2160 l=1080
+ ad=1.29888e+07 pd=40560 as=0 ps=0 
M1676 GND GND GND GND efet w=840 l=4200
+ ad=0 pd=0 as=0 ps=0 
M1677 GND GND GND GND efet w=1260 l=900
+ ad=0 pd=0 as=0 ps=0 
M1678 GND GND diff_44400_224400# GND efet w=540 l=2460
+ ad=0 pd=0 as=0 ps=0 
M1679 GND GND GND GND efet w=6600 l=2280
+ ad=0 pd=0 as=0 ps=0 
M1680 diff_26520_220920# diff_22800_212640# GND GND efet w=1980 l=1260
+ ad=1.21536e+07 pd=32400 as=0 ps=0 
M1681 GND diff_23400_208080# diff_26520_220920# GND efet w=1680 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1682 diff_22800_212640# diff_20760_213720# diff_22800_212640# GND efet w=4740 l=1200
+ ad=5.04e+06 pd=25680 as=0 ps=0 
M1683 diff_20760_213720# GND GND GND efet w=600 l=960
+ ad=360000 pd=2400 as=0 ps=0 
M1684 GND diff_23400_208080# diff_22800_212640# GND efet w=1200 l=960
+ ad=0 pd=0 as=0 ps=0 
M1685 diff_38760_219600# GND GND GND efet w=660 l=5040
+ ad=4.9536e+06 pd=16320 as=0 ps=0 
M1686 GND GND diff_38760_219600# GND efet w=1320 l=840
+ ad=0 pd=0 as=0 ps=0 
M1687 diff_52080_238440# GND GND GND efet w=660 l=2220
+ ad=4.176e+06 pd=13920 as=0 ps=0 
M1688 diff_50160_238320# GND GND GND efet w=720 l=1800
+ ad=0 pd=0 as=0 ps=0 
M1689 diff_52080_238440# GND GND GND efet w=4200 l=960
+ ad=0 pd=0 as=0 ps=0 
M1690 GND diff_62040_223560# diff_52080_238440# GND efet w=3540 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1691 diff_51960_227760# GND GND GND efet w=4440 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1692 GND diff_65760_223560# diff_51960_227760# GND efet w=4140 l=960
+ ad=0 pd=0 as=0 ps=0 
M1693 GND GND diff_71760_233040# GND efet w=480 l=5160
+ ad=0 pd=0 as=0 ps=0 
M1694 GND GND diff_77640_238440# GND efet w=540 l=4140
+ ad=0 pd=0 as=0 ps=0 
M1695 diff_50160_238320# GND GND GND efet w=480 l=4320
+ ad=0 pd=0 as=0 ps=0 
M1696 GND GND GND GND efet w=1980 l=900
+ ad=0 pd=0 as=0 ps=0 
M1697 GND diff_143160_236160# diff_133560_235080# GND efet w=1260 l=900
+ ad=0 pd=0 as=0 ps=0 
M1698 diff_133560_235080# diff_143160_236160# GND GND efet w=1200 l=960
+ ad=0 pd=0 as=0 ps=0 
M1699 diff_161160_232920# diff_143160_236160# GND GND efet w=1200 l=840
+ ad=0 pd=0 as=0 ps=0 
M1700 diff_133560_235080# diff_143160_236160# GND GND efet w=1200 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1701 diff_133560_235080# diff_133560_235080# GND GND efet w=840 l=1500
+ ad=0 pd=0 as=0 ps=0 
M1702 diff_133560_235080# diff_133560_235080# GND GND efet w=960 l=1440
+ ad=0 pd=0 as=0 ps=0 
M1703 diff_133560_235080# diff_133560_235080# GND GND efet w=1140 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1704 diff_156720_230520# diff_133560_235080# GND GND efet w=1380 l=960
+ ad=0 pd=0 as=0 ps=0 
M1705 diff_161160_232920# diff_133560_235080# GND GND efet w=1260 l=900
+ ad=0 pd=0 as=0 ps=0 
M1706 diff_165720_226080# diff_133560_235080# GND GND efet w=1200 l=960
+ ad=0 pd=0 as=0 ps=0 
M1707 diff_133560_235080# diff_133560_235080# GND GND efet w=1200 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1708 diff_133560_235080# diff_142320_226920# diff_133560_235080# GND efet w=4860 l=2460
+ ad=0 pd=0 as=0 ps=0 
M1709 GND GND GND GND efet w=720 l=5400
+ ad=0 pd=0 as=0 ps=0 
M1710 diff_133560_235080# diff_137400_226080# diff_133560_235080# GND efet w=1320 l=4200
+ ad=0 pd=0 as=0 ps=0 
M1711 diff_83160_218280# GND GND GND efet w=720 l=1320
+ ad=7.4592e+06 pd=22080 as=0 ps=0 
M1712 diff_110040_229200# GND GND GND efet w=600 l=5400
+ ad=3.7584e+06 pd=13680 as=0 ps=0 
M1713 GND diff_110040_208680# diff_110040_229200# GND efet w=1200 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1714 diff_99360_217440# GND GND GND efet w=720 l=5640
+ ad=1.18944e+07 pd=37200 as=0 ps=0 
M1715 GND diff_110040_208680# diff_99360_217440# GND efet w=1260 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1716 diff_110040_208680# diff_110040_229200# GND GND efet w=1080 l=960
+ ad=8.352e+06 pd=28560 as=0 ps=0 
M1717 GND GND diff_110040_208680# GND efet w=540 l=5580
+ ad=0 pd=0 as=0 ps=0 
M1718 diff_117120_227880# diff_110040_229200# GND GND efet w=1200 l=1080
+ ad=3.5712e+06 pd=13440 as=0 ps=0 
M1719 GND GND diff_117120_227880# GND efet w=720 l=5520
+ ad=0 pd=0 as=0 ps=0 
M1720 diff_63960_210840# GND GND GND efet w=1380 l=1260
+ ad=0 pd=0 as=0 ps=0 
M1721 diff_99360_217440# diff_110160_224880# diff_110640_223320# GND efet w=720 l=960
+ ad=0 pd=0 as=446400 ps=2880 
M1722 diff_117120_227880# diff_110160_224880# diff_115080_221040# GND efet w=780 l=1020
+ ad=0 pd=0 as=417600 ps=3360 
M1723 diff_38760_219600# GND diff_58200_222720# GND efet w=600 l=1080
+ ad=0 pd=0 as=388800 ps=2880 
M1724 diff_62040_223560# GND diff_35040_214560# GND efet w=600 l=960
+ ad=374400 pd=2640 as=3.6432e+06 ps=12480 
M1725 diff_65760_223560# GND diff_30480_212760# GND efet w=660 l=1140
+ ad=374400 pd=2640 as=6.2496e+06 ps=19680 
M1726 diff_22800_212640# diff_20760_213720# GND GND efet w=660 l=3120
+ ad=0 pd=0 as=0 ps=0 
M1727 diff_35040_214560# diff_21360_45480# GND GND efet w=1200 l=960
+ ad=0 pd=0 as=0 ps=0 
M1728 GND diff_21360_57480# diff_30480_212760# GND efet w=1320 l=840
+ ad=0 pd=0 as=0 ps=0 
M1729 GND GND diff_30480_212760# GND efet w=780 l=4620
+ ad=0 pd=0 as=0 ps=0 
M1730 GND GND diff_23400_208080# GND efet w=540 l=3060
+ ad=0 pd=0 as=7.3728e+06 ps=36000 
M1731 diff_23400_208080# GND diff_21960_203880# GND efet w=4020 l=1260
+ ad=0 pd=0 as=2.232e+06 ps=8640 
M1732 diff_21960_203880# diff_19080_201840# GND GND efet w=3660 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1733 GND GND diff_16920_200160# GND efet w=540 l=3420
+ ad=0 pd=0 as=5.5008e+06 ps=22320 
M1734 GND GND diff_23400_208080# GND efet w=1440 l=1500
+ ad=0 pd=0 as=0 ps=0 
M1735 diff_23400_208080# diff_20640_113640# GND GND efet w=1920 l=720
+ ad=0 pd=0 as=0 ps=0 
M1736 GND GND diff_35040_214560# GND efet w=540 l=4380
+ ad=0 pd=0 as=0 ps=0 
M1737 diff_19080_201840# GND diff_16920_200160# GND efet w=1200 l=960
+ ad=1.6704e+06 pd=6240 as=0 ps=0 
M1738 GND GND diff_16920_200160# GND efet w=1740 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1739 diff_50160_238320# GND GND GND efet w=3600 l=960
+ ad=0 pd=0 as=0 ps=0 
M1740 diff_72840_236280# GND GND GND efet w=1080 l=840
+ ad=9.3168e+06 pd=27360 as=0 ps=0 
M1741 diff_77640_236160# GND GND GND efet w=1680 l=840
+ ad=7.1136e+06 pd=30480 as=0 ps=0 
M1742 diff_72840_236280# diff_74880_222120# GND GND efet w=1020 l=840
+ ad=0 pd=0 as=0 ps=0 
M1743 diff_77640_236160# diff_74880_222120# GND GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M1744 GND diff_83400_222240# diff_83160_218280# GND efet w=1680 l=840
+ ad=0 pd=0 as=0 ps=0 
M1745 diff_63960_210840# diff_83400_222240# GND GND efet w=1680 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1746 diff_72840_236280# diff_73200_214320# diff_72840_236280# GND efet w=2520 l=2940
+ ad=0 pd=0 as=0 ps=0 
M1747 GND diff_11280_215400# diff_16920_200160# GND efet w=1920 l=960
+ ad=0 pd=0 as=0 ps=0 
M1748 GND GND diff_41520_198840# GND efet w=600 l=5760
+ ad=0 pd=0 as=1.36512e+07 ps=45360 
M1749 diff_72840_236280# diff_73200_214320# GND GND efet w=600 l=4680
+ ad=0 pd=0 as=0 ps=0 
M1750 diff_77640_236160# diff_78120_219240# diff_77640_236160# GND efet w=5040 l=2520
+ ad=0 pd=0 as=0 ps=0 
M1751 diff_83160_218280# diff_82680_213840# diff_83160_218280# GND efet w=2460 l=4980
+ ad=0 pd=0 as=0 ps=0 
M1752 GND diff_110640_223320# diff_112200_220320# GND efet w=3240 l=960
+ ad=0 pd=0 as=1.584e+06 ps=7200 
M1753 diff_63960_210840# diff_87600_213720# diff_63960_210840# GND efet w=5160 l=2640
+ ad=0 pd=0 as=0 ps=0 
M1754 diff_77640_236160# diff_78120_219240# GND GND efet w=600 l=4560
+ ad=0 pd=0 as=0 ps=0 
M1755 diff_83160_218280# diff_82680_213840# GND GND efet w=600 l=4680
+ ad=0 pd=0 as=0 ps=0 
M1756 diff_74880_222120# diff_83400_222240# GND GND efet w=2040 l=960
+ ad=2.7936e+06 pd=9360 as=0 ps=0 
M1757 GND GND diff_74880_222120# GND efet w=720 l=5520
+ ad=0 pd=0 as=0 ps=0 
M1758 diff_112200_220320# diff_110040_208680# diff_110040_229200# GND efet w=1800 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1759 diff_116040_220560# diff_115080_221040# GND GND efet w=3240 l=1080
+ ad=1.5408e+06 pd=6720 as=0 ps=0 
M1760 diff_110040_208680# diff_110040_208680# diff_116040_220560# GND efet w=1080 l=1680
+ ad=0 pd=0 as=0 ps=0 
M1761 diff_133560_235080# diff_137400_226080# GND GND efet w=840 l=4620
+ ad=0 pd=0 as=0 ps=0 
M1762 diff_133560_235080# diff_146760_226200# diff_133560_235080# GND efet w=2340 l=2580
+ ad=0 pd=0 as=0 ps=0 
M1763 diff_133560_235080# diff_142320_226920# GND GND efet w=660 l=4980
+ ad=0 pd=0 as=0 ps=0 
M1764 diff_133560_235080# diff_146760_226200# GND GND efet w=600 l=4680
+ ad=0 pd=0 as=0 ps=0 
M1765 diff_133560_235080# diff_151680_228720# diff_133560_235080# GND efet w=2460 l=4560
+ ad=0 pd=0 as=0 ps=0 
M1766 diff_156720_230520# diff_156120_226800# diff_156720_230520# GND efet w=2460 l=4380
+ ad=0 pd=0 as=0 ps=0 
M1767 diff_161160_232920# diff_161040_229440# diff_161160_232920# GND efet w=2460 l=4380
+ ad=0 pd=0 as=0 ps=0 
M1768 diff_165720_226080# diff_165720_226080# diff_165720_226080# GND efet w=2400 l=2700
+ ad=0 pd=0 as=0 ps=0 
M1769 diff_133560_235080# diff_151680_228720# GND GND efet w=600 l=4680
+ ad=0 pd=0 as=0 ps=0 
M1770 diff_156720_230520# diff_156120_226800# GND GND efet w=720 l=4920
+ ad=0 pd=0 as=0 ps=0 
M1771 diff_161160_232920# diff_161040_229440# GND GND efet w=780 l=4500
+ ad=0 pd=0 as=0 ps=0 
M1772 diff_165720_226080# diff_165720_226080# GND GND efet w=780 l=4620
+ ad=0 pd=0 as=0 ps=0 
M1773 GND GND diff_148080_240000# GND efet w=420 l=3420
+ ad=0 pd=0 as=0 ps=0 
M1774 GND GND diff_133560_235080# GND efet w=960 l=3540
+ ad=0 pd=0 as=0 ps=0 
M1775 diff_133560_235080# diff_170640_228120# diff_133560_235080# GND efet w=2520 l=2580
+ ad=0 pd=0 as=0 ps=0 
M1776 diff_133560_235080# diff_143160_236160# GND GND efet w=2160 l=840
+ ad=0 pd=0 as=0 ps=0 
M1777 diff_143160_236160# diff_133560_222480# GND GND efet w=4020 l=900
+ ad=4.104e+06 pd=14880 as=0 ps=0 
M1778 GND GND diff_143160_236160# GND efet w=840 l=3660
+ ad=0 pd=0 as=0 ps=0 
M1779 diff_133560_235080# diff_170640_228120# GND GND efet w=600 l=4440
+ ad=0 pd=0 as=0 ps=0 
M1780 GND diff_188880_226560# diff_133560_222480# GND efet w=720 l=1080
+ ad=0 pd=0 as=1.00656e+07 ps=36960 
M1781 GND diff_188880_226560# diff_164160_221520# GND efet w=600 l=1080
+ ad=0 pd=0 as=1.06848e+07 ps=27840 
M1782 diff_137400_226080# GND GND GND efet w=720 l=960
+ ad=619200 pd=3600 as=0 ps=0 
M1783 diff_142320_226920# GND GND GND efet w=720 l=1020
+ ad=532800 pd=3120 as=0 ps=0 
M1784 diff_146760_226200# GND GND GND efet w=840 l=840
+ ad=633600 pd=3360 as=0 ps=0 
M1785 diff_151680_228720# GND GND GND efet w=840 l=840
+ ad=619200 pd=3360 as=0 ps=0 
M1786 diff_156120_226800# GND GND GND efet w=720 l=840
+ ad=532800 pd=3120 as=0 ps=0 
M1787 diff_161040_229440# GND GND GND efet w=780 l=900
+ ad=518400 pd=2880 as=0 ps=0 
M1788 diff_165720_226080# GND GND GND efet w=900 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1789 diff_170640_228120# GND GND GND efet w=840 l=960
+ ad=604800 pd=3120 as=0 ps=0 
M1790 GND GND diff_134880_217080# GND efet w=480 l=5700
+ ad=0 pd=0 as=7.8192e+06 ps=19440 
M1791 GND GND diff_140640_215520# GND efet w=540 l=5460
+ ad=0 pd=0 as=8.5968e+06 ps=23760 
M1792 GND GND diff_148200_217200# GND efet w=480 l=5520
+ ad=0 pd=0 as=2.6352e+06 ps=10800 
M1793 GND GND diff_158880_215640# GND efet w=480 l=5280
+ ad=0 pd=0 as=7.3728e+06 ps=17280 
M1794 diff_133560_222480# diff_138120_220200# diff_140160_216480# GND efet w=720 l=960
+ ad=0 pd=0 as=7.0272e+06 ps=19440 
M1795 GND GND diff_140160_216480# GND efet w=480 l=2760
+ ad=0 pd=0 as=0 ps=0 
M1796 GND GND diff_164520_215520# GND efet w=480 l=6000
+ ad=0 pd=0 as=8.9568e+06 ps=24240 
M1797 GND GND diff_172080_217080# GND efet w=480 l=5280
+ ad=0 pd=0 as=2.736e+06 ps=10320 
M1798 GND GND diff_164040_216360# GND efet w=540 l=3420
+ ad=0 pd=0 as=7.4016e+06 ps=19200 
M1799 diff_164160_221520# diff_138120_220200# diff_164040_216360# GND efet w=900 l=900
+ ad=0 pd=0 as=0 ps=0 
M1800 diff_63960_210840# diff_87600_213720# GND GND efet w=600 l=4440
+ ad=0 pd=0 as=0 ps=0 
M1801 GND diff_20640_113640# diff_94080_217680# GND efet w=720 l=960
+ ad=0 pd=0 as=0 ps=0 
M1802 diff_99360_217440# GND GND GND efet w=720 l=960
+ ad=0 pd=0 as=0 ps=0 
M1803 diff_83400_222240# diff_20640_113640# diff_94080_215520# GND efet w=720 l=960
+ ad=892800 pd=6480 as=0 ps=0 
M1804 diff_99360_215760# GND diff_83400_222240# GND efet w=660 l=1080
+ ad=1.39248e+07 pd=41520 as=0 ps=0 
M1805 diff_57000_209520# diff_56520_205560# diff_57000_209520# GND efet w=6120 l=2400
+ ad=1.31904e+07 pd=51600 as=0 ps=0 
M1806 GND GND diff_64080_204360# GND efet w=540 l=4980
+ ad=0 pd=0 as=1.1664e+06 ps=6720 
M1807 diff_73200_214320# GND GND GND efet w=840 l=960
+ ad=604800 pd=3120 as=0 ps=0 
M1808 diff_78120_219240# GND GND GND efet w=960 l=840
+ ad=590400 pd=3120 as=0 ps=0 
M1809 diff_82680_213840# GND GND GND efet w=900 l=840
+ ad=604800 pd=3360 as=0 ps=0 
M1810 diff_87600_213720# GND GND GND efet w=960 l=960
+ ad=561600 pd=3360 as=0 ps=0 
M1811 diff_63960_210840# diff_57000_209520# GND GND efet w=3420 l=1740
+ ad=0 pd=0 as=0 ps=0 
M1812 GND GND diff_56520_205560# GND efet w=660 l=1020
+ ad=0 pd=0 as=331200 ps=2640 
M1813 GND GND diff_49320_199200# GND efet w=2820 l=1140
+ ad=0 pd=0 as=1.512e+06 ps=6240 
M1814 GND diff_56520_205560# diff_57000_209520# GND efet w=480 l=3600
+ ad=0 pd=0 as=0 ps=0 
M1815 GND diff_64080_204360# diff_63960_210840# GND efet w=2460 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1816 GND GND GND GND efet w=540 l=5700
+ ad=0 pd=0 as=0 ps=0 
M1817 diff_47040_199200# GND diff_41520_198840# GND efet w=2520 l=960
+ ad=3.3264e+06 pd=7680 as=0 ps=0 
M1818 diff_49320_199200# diff_45720_176880# diff_47040_199200# GND efet w=2520 l=960
+ ad=0 pd=0 as=0 ps=0 
M1819 diff_50880_194400# GND GND GND efet w=2700 l=1020
+ ad=4.608e+06 pd=19680 as=0 ps=0 
M1820 diff_41520_198840# diff_11280_215400# GND GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M1821 diff_50880_194400# GND diff_49320_194400# GND efet w=3060 l=1680
+ ad=0 pd=0 as=1.44e+06 ps=6000 
M1822 diff_43800_194280# GND GND GND efet w=2520 l=1080
+ ad=1.7712e+06 pd=6480 as=0 ps=0 
M1823 diff_45480_194400# diff_44520_186120# diff_43800_194280# GND efet w=2400 l=1080
+ ad=1.4976e+06 pd=6240 as=0 ps=0 
M1824 GND GND diff_45480_194400# GND efet w=2100 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1825 diff_49320_194400# diff_45720_176880# GND GND efet w=2400 l=960
+ ad=0 pd=0 as=0 ps=0 
M1826 diff_52440_194280# diff_51480_191880# diff_50880_194400# GND efet w=2520 l=960
+ ad=1.512e+06 pd=6240 as=0 ps=0 
M1827 GND diff_53040_193920# diff_52440_194280# GND efet w=2580 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1828 diff_64080_204360# diff_57000_209520# GND GND efet w=1080 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1829 GND GND diff_70800_207960# GND efet w=720 l=4260
+ ad=0 pd=0 as=1.512e+06 ps=8880 
M1830 GND diff_70800_207960# diff_69480_207240# GND efet w=1680 l=840
+ ad=0 pd=0 as=0 ps=0 
M1831 GND diff_80640_207120# diff_70800_206280# GND efet w=600 l=3360
+ ad=0 pd=0 as=9.4752e+06 ps=48000 
M1832 GND GND diff_80640_207120# GND efet w=480 l=840
+ ad=0 pd=0 as=345600 ps=2400 
M1833 diff_86640_208320# GND GND GND efet w=480 l=960
+ ad=388800 pd=2880 as=0 ps=0 
M1834 GND diff_86640_208320# diff_86760_205920# GND efet w=660 l=1500
+ ad=0 pd=0 as=1.9944e+07 ps=62400 
M1835 diff_70800_206280# diff_80640_207120# diff_70800_206280# GND efet w=4020 l=1920
+ ad=0 pd=0 as=0 ps=0 
M1836 GND diff_70800_206280# diff_69480_207240# GND efet w=1740 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1837 GND diff_70800_206280# diff_70800_207960# GND efet w=1140 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1838 diff_86760_205920# diff_86640_208320# diff_86760_205920# GND efet w=6780 l=1860
+ ad=0 pd=0 as=0 ps=0 
M1839 diff_86760_205920# diff_92760_202560# GND GND efet w=2940 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1840 GND GND diff_86760_205920# GND efet w=1860 l=2100
+ ad=0 pd=0 as=0 ps=0 
M1841 GND diff_95880_204840# diff_86760_205920# GND efet w=2880 l=960
+ ad=0 pd=0 as=0 ps=0 
M1842 GND GND diff_66840_200160# GND efet w=480 l=4200
+ ad=0 pd=0 as=1.224e+06 ps=7680 
M1843 diff_57000_209520# GND GND GND efet w=1140 l=900
+ ad=0 pd=0 as=0 ps=0 
M1844 diff_70800_206280# diff_77400_204960# GND GND efet w=1140 l=900
+ ad=0 pd=0 as=0 ps=0 
M1845 diff_70800_206280# diff_75120_202800# diff_74040_202080# GND efet w=2460 l=900
+ ad=0 pd=0 as=2.4192e+06 ps=9360 
M1846 diff_57000_209520# GND GND GND efet w=1260 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1847 GND diff_64920_198240# diff_57000_209520# GND efet w=1200 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1848 diff_57000_209520# diff_66840_200160# GND GND efet w=1200 l=960
+ ad=0 pd=0 as=0 ps=0 
M1849 diff_74040_202080# diff_44520_186120# GND GND efet w=2460 l=900
+ ad=0 pd=0 as=0 ps=0 
M1850 GND diff_73200_192960# diff_70800_206280# GND efet w=1260 l=900
+ ad=0 pd=0 as=0 ps=0 
M1851 GND diff_21360_57480# GND GND efet w=1500 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1852 diff_66840_200160# GND GND GND efet w=1200 l=840
+ ad=0 pd=0 as=0 ps=0 
M1853 GND diff_44520_147840# diff_53040_193920# GND efet w=2820 l=1140
+ ad=0 pd=0 as=8.5392e+06 ps=33600 
M1854 diff_53040_193920# GND GND GND efet w=2220 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1855 diff_45600_181560# GND GND GND efet w=2700 l=840
+ ad=1.8144e+06 pd=6480 as=0 ps=0 
M1856 GND diff_21360_45480# GND GND efet w=1020 l=900
+ ad=0 pd=0 as=0 ps=0 
M1857 diff_47160_181560# diff_44520_186120# diff_45600_181560# GND efet w=2640 l=840
+ ad=1.7424e+06 pd=6720 as=0 ps=0 
M1858 GND GND diff_47160_181560# GND efet w=1980 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1859 GND GND GND GND efet w=660 l=5340
+ ad=0 pd=0 as=0 ps=0 
M1860 diff_52440_182520# diff_45720_176880# diff_50880_179400# GND efet w=3000 l=960
+ ad=1.9728e+06 pd=7680 as=1.11888e+07 ps=31680 
M1861 GND GND diff_52440_182520# GND efet w=3180 l=900
+ ad=0 pd=0 as=0 ps=0 
M1862 diff_56280_181320# diff_51480_191880# GND GND efet w=2760 l=960
+ ad=1.656e+06 pd=6720 as=0 ps=0 
M1863 diff_50880_179400# diff_53040_193920# diff_56280_181320# GND efet w=2760 l=960
+ ad=0 pd=0 as=0 ps=0 
M1864 GND diff_20640_113640# diff_50880_179400# GND efet w=2880 l=840
+ ad=0 pd=0 as=0 ps=0 
M1865 GND GND diff_45720_176880# GND efet w=2280 l=900
+ ad=0 pd=0 as=2.0448e+06 ps=8640 
M1866 diff_45720_176880# GND GND GND efet w=480 l=2280
+ ad=0 pd=0 as=0 ps=0 
M1867 diff_53040_193920# GND GND GND efet w=540 l=2340
+ ad=0 pd=0 as=0 ps=0 
M1868 diff_44040_172320# diff_49320_172200# GND GND efet w=540 l=2340
+ ad=5.8752e+06 pd=30000 as=0 ps=0 
M1869 GND diff_44040_172320# GND GND efet w=3120 l=960
+ ad=0 pd=0 as=0 ps=0 
M1870 GND GND diff_49320_172200# GND efet w=480 l=1140
+ ad=0 pd=0 as=316800 ps=2400 
M1871 GND diff_20640_113640# diff_64920_198240# GND efet w=1260 l=1020
+ ad=0 pd=0 as=6.336e+06 ps=24720 
M1872 GND GND diff_64920_198240# GND efet w=1020 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1873 GND GND diff_77400_204960# GND efet w=540 l=4260
+ ad=0 pd=0 as=2.376e+06 ps=8160 
M1874 diff_64920_198240# GND GND GND efet w=480 l=5520
+ ad=0 pd=0 as=0 ps=0 
M1875 diff_77400_204960# GND GND GND efet w=1200 l=840
+ ad=0 pd=0 as=0 ps=0 
M1876 GND GND diff_72240_189360# GND efet w=480 l=2280
+ ad=0 pd=0 as=4.896e+06 ps=18480 
M1877 GND GND GND GND efet w=480 l=2400
+ ad=0 pd=0 as=0 ps=0 
M1878 diff_90840_198360# GND GND GND efet w=660 l=4500
+ ad=9.5328e+06 pd=28080 as=0 ps=0 
M1879 diff_92760_202560# GND diff_90840_198360# GND efet w=780 l=1260
+ ad=1.0224e+06 pd=5520 as=0 ps=0 
M1880 diff_110040_208680# GND GND GND efet w=540 l=6060
+ ad=0 pd=0 as=0 ps=0 
M1881 GND diff_110160_224880# diff_110040_208680# GND efet w=960 l=960
+ ad=0 pd=0 as=0 ps=0 
M1882 GND diff_110160_224880# diff_99360_215760# GND efet w=1560 l=840
+ ad=0 pd=0 as=0 ps=0 
M1883 diff_99360_215760# GND GND GND efet w=660 l=5700
+ ad=0 pd=0 as=0 ps=0 
M1884 diff_110160_224880# diff_110040_208680# GND GND efet w=1080 l=960
+ ad=1.78704e+07 pd=66720 as=0 ps=0 
M1885 GND GND diff_110160_224880# GND efet w=540 l=5400
+ ad=0 pd=0 as=0 ps=0 
M1886 diff_117120_215640# diff_110040_208680# GND GND efet w=1200 l=960
+ ad=3.5424e+06 pd=13680 as=0 ps=0 
M1887 GND GND diff_117120_215640# GND efet w=780 l=6300
+ ad=0 pd=0 as=0 ps=0 
M1888 diff_110640_210960# GND diff_99360_215760# GND efet w=720 l=900
+ ad=417600 pd=2880 as=0 ps=0 
M1889 diff_117120_215640# GND diff_115080_208680# GND efet w=600 l=840
+ ad=0 pd=0 as=432000 ps=2640 
M1890 diff_140160_216480# GND diff_134040_213360# GND efet w=660 l=1260
+ ad=0 pd=0 as=345600 ps=2400 
M1891 diff_134880_217080# diff_133320_215640# diff_134640_214200# GND efet w=2040 l=1020
+ ad=0 pd=0 as=1.6416e+06 ps=7200 
M1892 diff_134640_214200# diff_134040_213360# GND GND efet w=2820 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1893 GND diff_140640_215520# diff_140160_216480# GND efet w=1800 l=960
+ ad=0 pd=0 as=0 ps=0 
M1894 GND diff_140640_215520# diff_134880_217080# GND efet w=1020 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1895 GND GND diff_148200_217200# GND efet w=660 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1896 diff_148200_217200# diff_134880_217080# GND GND efet w=1020 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1897 diff_140640_215520# diff_134880_217080# GND GND efet w=1020 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1898 diff_164040_216360# diff_134880_217080# diff_157920_213240# GND efet w=840 l=1020
+ ad=0 pd=0 as=273600 ps=2400 
M1899 GND diff_110640_210960# diff_112200_208080# GND efet w=3240 l=1080
+ ad=0 pd=0 as=1.5408e+06 ps=6960 
M1900 GND GND diff_102600_202200# GND efet w=600 l=5400
+ ad=0 pd=0 as=2.88e+06 ps=14160 
M1901 diff_105120_208440# GND GND GND efet w=540 l=2340
+ ad=0 pd=0 as=0 ps=0 
M1902 diff_112200_208080# diff_110160_224880# diff_110040_208680# GND efet w=1620 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1903 diff_116040_208080# diff_115080_208680# GND GND efet w=3240 l=960
+ ad=1.5408e+06 pd=6720 as=0 ps=0 
M1904 diff_110160_224880# diff_110160_224880# diff_116040_208080# GND efet w=1380 l=1380
+ ad=0 pd=0 as=0 ps=0 
M1905 GND diff_124200_197520# GND GND efet w=3360 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1906 GND diff_102600_202200# diff_105120_208440# GND efet w=2160 l=960
+ ad=0 pd=0 as=0 ps=0 
M1907 GND GND diff_95880_204840# GND efet w=480 l=3000
+ ad=0 pd=0 as=3.888e+06 ps=15120 
M1908 diff_110160_224880# diff_109680_203520# GND GND efet w=2220 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1909 GND diff_89040_188280# GND GND efet w=2580 l=1260
+ ad=0 pd=0 as=0 ps=0 
M1910 diff_140640_215520# diff_133320_215640# diff_152280_214200# GND efet w=1740 l=1020
+ ad=0 pd=0 as=1.6704e+06 ps=6960 
M1911 diff_175200_217320# diff_134880_217080# diff_172080_217080# GND efet w=720 l=1080
+ ad=403200 pd=2880 as=0 ps=0 
M1912 GND diff_158880_215640# diff_172080_217080# GND efet w=1080 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1913 diff_158880_215640# diff_140640_215520# diff_158520_214320# GND efet w=1800 l=1080
+ ad=0 pd=0 as=1.6848e+06 ps=6960 
M1914 GND diff_164520_215520# diff_164040_216360# GND efet w=1800 l=840
+ ad=0 pd=0 as=0 ps=0 
M1915 diff_158880_215640# diff_164520_215520# GND GND efet w=960 l=840
+ ad=0 pd=0 as=0 ps=0 
M1916 diff_152280_214200# GND GND GND efet w=2100 l=1920
+ ad=0 pd=0 as=0 ps=0 
M1917 diff_158520_214320# diff_157920_213240# GND GND efet w=2760 l=960
+ ad=0 pd=0 as=0 ps=0 
M1918 GND GND GND GND efet w=2400 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1919 GND GND diff_110160_224880# GND efet w=780 l=2520
+ ad=0 pd=0 as=0 ps=0 
M1920 GND GND diff_106680_199920# GND efet w=2460 l=1260
+ ad=0 pd=0 as=2.0304e+06 ps=7440 
M1921 diff_106680_199920# GND diff_105120_200040# GND efet w=2580 l=1020
+ ad=0 pd=0 as=1.4688e+06 ps=6240 
M1922 GND GND diff_72240_189360# GND efet w=2160 l=1140
+ ad=0 pd=0 as=0 ps=0 
M1923 GND diff_84720_180000# GND GND efet w=2160 l=960
+ ad=0 pd=0 as=0 ps=0 
M1924 GND diff_20640_113640# diff_90840_198360# GND efet w=1560 l=960
+ ad=0 pd=0 as=0 ps=0 
M1925 diff_95880_204840# GND GND GND efet w=1920 l=960
+ ad=0 pd=0 as=0 ps=0 
M1926 diff_105120_200040# diff_72240_189360# diff_102600_202200# GND efet w=2400 l=960
+ ad=0 pd=0 as=0 ps=0 
M1927 diff_71760_186600# diff_20640_113640# GND GND efet w=1800 l=1080
+ ad=1.08e+06 pd=4800 as=0 ps=0 
M1928 diff_73200_192960# GND diff_71640_183960# GND efet w=660 l=1020
+ ad=518400 pd=4080 as=5.76e+06 ps=22560 
M1929 diff_71640_183960# diff_72240_189360# diff_71760_186600# GND efet w=1800 l=960
+ ad=0 pd=0 as=0 ps=0 
M1930 diff_75120_202800# GND GND GND efet w=1200 l=900
+ ad=3.2976e+06 pd=13680 as=0 ps=0 
M1931 GND GND diff_83040_186840# GND efet w=480 l=4320
+ ad=0 pd=0 as=2.088e+06 ps=9360 
M1932 diff_71640_183960# GND GND GND efet w=480 l=5400
+ ad=0 pd=0 as=0 ps=0 
M1933 diff_71640_183960# diff_11280_215400# GND GND efet w=1200 l=900
+ ad=0 pd=0 as=0 ps=0 
M1934 diff_75120_202800# GND GND GND efet w=600 l=3960
+ ad=0 pd=0 as=0 ps=0 
M1935 GND GND diff_90840_198360# GND efet w=1260 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1936 GND diff_89040_188280# diff_84720_183480# GND efet w=2460 l=1020
+ ad=0 pd=0 as=1.07136e+07 ps=35040 
M1937 GND diff_44520_147840# diff_83040_186840# GND efet w=1380 l=960
+ ad=0 pd=0 as=0 ps=0 
M1938 GND GND diff_90600_186120# GND efet w=1800 l=960
+ ad=0 pd=0 as=1.08e+06 ps=4800 
M1939 diff_90600_186120# diff_44520_186120# diff_84720_180000# GND efet w=2100 l=900
+ ad=0 pd=0 as=1.13328e+07 ps=34320 
M1940 diff_84720_183480# diff_83040_186840# diff_84720_181920# GND efet w=2460 l=1020
+ ad=0 pd=0 as=1.44e+06 ps=6000 
M1941 diff_109680_203520# GND diff_109680_203520# GND efet w=240 l=5520
+ ad=1.17072e+07 pd=48960 as=0 ps=0 
M1942 diff_109080_192240# GND GND GND efet w=2520 l=960
+ ad=1.512e+06 pd=6240 as=0 ps=0 
M1943 diff_110640_192240# diff_20640_113640# diff_109080_192240# GND efet w=2640 l=960
+ ad=1.4976e+06 pd=6480 as=0 ps=0 
M1944 diff_109680_203520# diff_89040_188280# diff_110640_192240# GND efet w=2520 l=960
+ ad=0 pd=0 as=0 ps=0 
M1945 GND GND diff_115200_193800# GND efet w=480 l=2760
+ ad=0 pd=0 as=2.4192e+06 ps=10800 
M1946 GND GND diff_119880_192240# GND efet w=480 l=5820
+ ad=0 pd=0 as=6.7824e+06 ps=22800 
M1947 diff_124200_197520# GND diff_119880_192240# GND efet w=1080 l=1080
+ ad=619200 pd=3600 as=0 ps=0 
M1948 GND GND diff_115200_193800# GND efet w=1800 l=960
+ ad=0 pd=0 as=0 ps=0 
M1949 diff_164520_215520# diff_158880_215640# GND GND efet w=1020 l=900
+ ad=0 pd=0 as=0 ps=0 
M1950 diff_164520_215520# diff_140640_215520# diff_176640_214080# GND efet w=1800 l=1080
+ ad=0 pd=0 as=1.656e+06 ps=7200 
M1951 diff_176640_214080# diff_175200_217320# GND GND efet w=3000 l=960
+ ad=0 pd=0 as=0 ps=0 
M1952 GND diff_188880_226560# diff_183360_241080# GND efet w=840 l=1080
+ ad=0 pd=0 as=9.2016e+06 ps=27120 
M1953 GND GND diff_183120_215520# GND efet w=480 l=5400
+ ad=0 pd=0 as=7.56e+06 ps=17760 
M1954 GND GND diff_188760_215400# GND efet w=540 l=5580
+ ad=0 pd=0 as=9.2736e+06 ps=24000 
M1955 GND GND diff_196440_216960# GND efet w=600 l=5760
+ ad=0 pd=0 as=2.7072e+06 ps=10320 
M1956 diff_183360_241080# diff_138120_220200# diff_188280_216360# GND efet w=600 l=960
+ ad=0 pd=0 as=7.0272e+06 ps=18480 
M1957 GND GND diff_188280_216360# GND efet w=420 l=2820
+ ad=0 pd=0 as=0 ps=0 
M1958 diff_188280_216360# diff_158880_215640# diff_182160_213240# GND efet w=660 l=1020
+ ad=0 pd=0 as=273600 ps=2880 
M1959 diff_183120_215520# diff_164520_215520# diff_182880_214080# GND efet w=1740 l=1020
+ ad=0 pd=0 as=1.8864e+06 ps=7200 
M1960 GND diff_188760_215400# diff_188280_216360# GND efet w=1800 l=960
+ ad=0 pd=0 as=0 ps=0 
M1961 diff_183120_215520# diff_188760_215400# GND GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M1962 diff_182880_214080# diff_182160_213240# GND GND efet w=3000 l=960
+ ad=0 pd=0 as=0 ps=0 
M1963 GND diff_158880_215640# diff_196440_216960# GND efet w=900 l=1260
+ ad=0 pd=0 as=0 ps=0 
M1964 diff_196440_216960# diff_183120_215520# GND GND efet w=960 l=840
+ ad=0 pd=0 as=0 ps=0 
M1965 diff_188760_215400# diff_183120_215520# GND GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M1966 GND GND GND GND efet w=480 l=4260
+ ad=0 pd=0 as=0 ps=0 
M1967 GND diff_162960_208080# diff_123240_258000# GND efet w=2040 l=960
+ ad=0 pd=0 as=8.3952e+06 ps=22560 
M1968 GND diff_167280_200280# diff_133320_215640# GND efet w=1740 l=1020
+ ad=0 pd=0 as=4.7088e+06 ps=17280 
M1969 diff_171480_208680# diff_170760_206520# diff_171480_208680# GND efet w=4620 l=2280
+ ad=1.81296e+07 pd=72480 as=0 ps=0 
M1970 diff_117960_263280# diff_89040_188280# GND GND efet w=3240 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1971 GND GND diff_137400_197640# GND efet w=480 l=5880
+ ad=0 pd=0 as=6.5952e+06 ps=21600 
M1972 GND diff_141240_199080# diff_117960_263280# GND efet w=3060 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1973 GND diff_115200_193800# diff_110160_224880# GND efet w=2460 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1974 diff_137400_197640# GND diff_141240_199080# GND efet w=1380 l=900
+ ad=0 pd=0 as=792000 ps=4560 
M1975 diff_118320_192240# GND GND GND efet w=1860 l=1020
+ ad=1.0656e+06 pd=4800 as=0 ps=0 
M1976 diff_121680_193680# diff_120240_185760# diff_119880_192240# GND efet w=2700 l=1140
+ ad=1.4976e+06 pd=6480 as=0 ps=0 
M1977 diff_119880_192240# GND diff_118320_192240# GND efet w=1800 l=1020
+ ad=0 pd=0 as=0 ps=0 
M1978 diff_123480_192240# diff_20640_113640# diff_121680_193680# GND efet w=2460 l=1140
+ ad=1.2096e+06 pd=6000 as=0 ps=0 
M1979 diff_20640_113640# GND GND GND efet w=1980 l=1020
+ ad=1.14638e+08 pd=326160 as=0 ps=0 
M1980 diff_84720_181920# diff_51480_191880# diff_84720_180000# GND efet w=2400 l=960
+ ad=0 pd=0 as=0 ps=0 
M1981 diff_84720_180000# GND diff_84720_183480# GND efet w=1800 l=960
+ ad=0 pd=0 as=0 ps=0 
M1982 diff_20640_113640# diff_20640_113640# diff_109680_203520# GND efet w=1980 l=1260
+ ad=0 pd=0 as=0 ps=0 
M1983 diff_109680_203520# GND diff_20640_113640# GND efet w=1920 l=960
+ ad=0 pd=0 as=0 ps=0 
M1984 diff_109680_203520# diff_20640_113640# diff_20640_113640# GND efet w=1800 l=1080
+ ad=0 pd=0 as=0 ps=0 
M1985 GND GND diff_123480_192240# GND efet w=1440 l=2160
+ ad=0 pd=0 as=0 ps=0 
M1986 GND GND diff_117960_263280# GND efet w=2880 l=1320
+ ad=0 pd=0 as=0 ps=0 
M1987 diff_137400_197640# diff_20640_113640# diff_135600_195960# GND efet w=2580 l=1260
+ ad=0 pd=0 as=9.0288e+06 ps=31680 
M1988 GND diff_20640_113640# diff_128520_190200# GND efet w=3540 l=1140
+ ad=0 pd=0 as=4.9392e+06 ps=22320 
M1989 GND GND diff_89040_188280# GND efet w=720 l=2040
+ ad=0 pd=0 as=7.0128e+06 ps=28560 
M1990 diff_123240_258000# GND GND GND efet w=480 l=2760
+ ad=0 pd=0 as=0 ps=0 
M1991 diff_156600_191160# GND GND GND efet w=480 l=5760
+ ad=4.9824e+06 pd=23040 as=0 ps=0 
M1992 GND GND diff_117960_263280# GND efet w=600 l=2400
+ ad=0 pd=0 as=0 ps=0 
M1993 diff_133320_215640# GND GND GND efet w=480 l=3000
+ ad=0 pd=0 as=0 ps=0 
M1994 diff_171480_208680# diff_170760_206520# GND GND efet w=840 l=2280
+ ad=0 pd=0 as=0 ps=0 
M1995 diff_171480_208680# diff_174480_199320# GND GND efet w=3120 l=1200
+ ad=0 pd=0 as=0 ps=0 
M1996 diff_188760_215400# diff_164520_215520# diff_200880_213960# GND efet w=2040 l=1320
+ ad=0 pd=0 as=1.6704e+06 ps=6960 
M1997 diff_200880_213960# GND GND GND efet w=1800 l=1920
+ ad=0 pd=0 as=0 ps=0 
M1998 GND diff_180360_195360# diff_182160_210000# GND efet w=1020 l=1020
+ ad=0 pd=0 as=5.6448e+06 ps=24720 
M1999 diff_182160_210000# diff_181440_206520# diff_182160_210000# GND efet w=4380 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2000 GND diff_181440_206520# diff_182160_210000# GND efet w=540 l=4500
+ ad=0 pd=0 as=0 ps=0 
M2001 GND diff_180360_195360# diff_139680_251040# GND efet w=1680 l=960
+ ad=0 pd=0 as=0 ps=0 
M2002 GND diff_192240_207600# diff_198960_207240# GND efet w=960 l=960
+ ad=0 pd=0 as=2.3472e+06 ps=11760 
M2003 diff_192240_207600# diff_191520_202680# diff_192240_207600# GND efet w=4380 l=1500
+ ad=1.60704e+07 pd=57120 as=0 ps=0 
M2004 diff_139680_251040# diff_182160_210000# GND GND efet w=1560 l=960
+ ad=0 pd=0 as=0 ps=0 
M2005 diff_133560_235080# diff_198960_207240# GND GND efet w=2040 l=960
+ ad=0 pd=0 as=0 ps=0 
M2006 diff_170760_206520# GND GND GND efet w=540 l=900
+ ad=388800 pd=2880 as=0 ps=0 
M2007 diff_117960_263280# diff_156600_191160# GND GND efet w=2760 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2008 diff_135600_195960# diff_89400_129240# diff_135600_194640# GND efet w=4380 l=1020
+ ad=0 pd=0 as=2.5488e+06 ps=9840 
M2009 diff_130080_189840# diff_89400_129240# diff_128520_190200# GND efet w=6660 l=1080
+ ad=2.4336e+06 pd=11040 as=0 ps=0 
M2010 GND GND diff_130080_189840# GND efet w=3180 l=1500
+ ad=0 pd=0 as=0 ps=0 
M2011 GND GND diff_135600_194640# GND efet w=2100 l=1380
+ ad=0 pd=0 as=0 ps=0 
M2012 GND GND diff_143400_188160# GND efet w=2460 l=1140
+ ad=0 pd=0 as=4.2768e+06 ps=15600 
M2013 diff_89040_188280# GND GND GND efet w=4980 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2014 GND GND diff_135600_195960# GND efet w=1800 l=840
+ ad=0 pd=0 as=0 ps=0 
M2015 diff_120240_185760# diff_89400_129240# GND GND efet w=4560 l=960
+ ad=6.6528e+06 pd=21120 as=0 ps=0 
M2016 GND diff_89040_188280# diff_153120_192360# GND efet w=2520 l=960
+ ad=0 pd=0 as=1.512e+06 ps=6240 
M2017 diff_153120_192360# GND diff_153120_191040# GND efet w=2580 l=900
+ ad=0 pd=0 as=4.9392e+06 ps=17040 
M2018 diff_167280_200280# GND GND GND efet w=480 l=5880
+ ad=2.9376e+06 pd=10800 as=0 ps=0 
M2019 GND GND diff_174480_199320# GND efet w=480 l=5880
+ ad=0 pd=0 as=8.208e+06 ps=28560 
M2020 diff_181440_206520# GND GND GND efet w=600 l=960
+ ad=432000 pd=2640 as=0 ps=0 
M2021 diff_174480_199320# GND diff_174480_194280# GND efet w=2520 l=840
+ ad=0 pd=0 as=3.528e+06 ps=13680 
M2022 diff_167280_200280# GND diff_169320_193320# GND efet w=2520 l=960
+ ad=0 pd=0 as=2.9808e+06 ps=13440 
M2023 diff_192240_207600# diff_191520_202680# GND GND efet w=480 l=4320
+ ad=0 pd=0 as=0 ps=0 
M2024 diff_143400_188160# GND diff_143400_186720# GND efet w=3060 l=1020
+ ad=0 pd=0 as=4.896e+06 ps=21360 
M2025 diff_149880_184080# diff_148680_185160# GND GND efet w=2460 l=1200
+ ad=4.9248e+06 pd=14640 as=0 ps=0 
M2026 diff_84720_180000# GND GND GND efet w=480 l=5040
+ ad=0 pd=0 as=0 ps=0 
M2027 GND GND GND GND efet w=2640 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2028 diff_82080_164400# GND GND GND efet w=2700 l=900
+ ad=1.32336e+07 pd=50880 as=0 ps=0 
M2029 GND diff_89040_188280# diff_89160_121200# GND efet w=2040 l=960
+ ad=0 pd=0 as=1.60272e+07 ps=58320 
M2030 diff_120240_185760# GND GND GND efet w=480 l=2280
+ ad=0 pd=0 as=0 ps=0 
M2031 GND diff_145200_181200# diff_141720_184920# GND efet w=2340 l=1200
+ ad=0 pd=0 as=3.1248e+06 ps=13200 
M2032 diff_153120_191040# diff_89400_129240# diff_148680_185160# GND efet w=4500 l=1020
+ ad=0 pd=0 as=3.8016e+06 ps=14640 
M2033 diff_141720_184920# GND GND GND efet w=480 l=2280
+ ad=0 pd=0 as=0 ps=0 
M2034 diff_159960_191040# diff_149880_184080# diff_158400_186360# GND efet w=2820 l=1320
+ ad=1.2384e+06 pd=6480 as=4.1472e+06 ps=21600 
M2035 GND GND diff_159960_191040# GND efet w=2820 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2036 diff_163800_191040# diff_20640_113640# GND GND efet w=2580 l=1140
+ ad=1.2096e+06 pd=6000 as=0 ps=0 
M2037 diff_165360_185160# diff_149880_184080# diff_163800_191040# GND efet w=2520 l=1080
+ ad=4.608e+06 pd=18960 as=0 ps=0 
M2038 diff_158400_186360# GND diff_156600_191160# GND efet w=2820 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2039 diff_159960_184200# diff_89400_129240# diff_158400_186360# GND efet w=4440 l=1140
+ ad=1.728e+06 pd=9360 as=0 ps=0 
M2040 diff_145200_181200# GND diff_143400_186720# GND efet w=2580 l=1020
+ ad=2.0016e+06 pd=8400 as=0 ps=0 
M2041 GND GND diff_145200_181200# GND efet w=540 l=5340
+ ad=0 pd=0 as=0 ps=0 
M2042 diff_149880_184080# GND GND GND efet w=480 l=2280
+ ad=0 pd=0 as=0 ps=0 
M2043 diff_163800_185160# diff_141720_184920# GND GND efet w=2580 l=1140
+ ad=1.2096e+06 pd=6000 as=0 ps=0 
M2044 GND diff_141720_184920# diff_159960_184200# GND efet w=2520 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2045 diff_165360_185160# diff_120240_185760# diff_163800_185160# GND efet w=2520 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2046 diff_176040_194040# GND diff_174480_194280# GND efet w=2700 l=1260
+ ad=4.2912e+06 pd=15360 as=0 ps=0 
M2047 diff_170880_192840# diff_21360_45480# diff_169320_193320# GND efet w=2700 l=1140
+ ad=1.2096e+06 pd=6000 as=0 ps=0 
M2048 GND GND diff_170880_192840# GND efet w=2520 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2049 GND diff_20640_113640# diff_176040_194040# GND efet w=2580 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2050 GND GND diff_180360_195360# GND efet w=600 l=5640
+ ad=0 pd=0 as=1.1232e+07 ps=41520 
M2051 diff_191520_202680# GND GND GND efet w=540 l=900
+ ad=345600 pd=2400 as=0 ps=0 
M2052 GND GND diff_198960_207240# GND efet w=480 l=4320
+ ad=0 pd=0 as=0 ps=0 
M2053 diff_180360_195360# GND diff_180360_194040# GND efet w=3060 l=900
+ ad=0 pd=0 as=2.664e+06 ps=14400 
M2054 GND GND diff_180120_190560# GND efet w=2520 l=960
+ ad=0 pd=0 as=1.1088e+07 ps=28800 
M2055 diff_183600_181920# diff_20640_113640# diff_179760_181440# GND efet w=7020 l=1380
+ ad=1.65312e+07 pd=55680 as=1.58544e+07 ps=55200 
M2056 diff_180120_190560# diff_21360_45480# GND GND efet w=3000 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2057 GND diff_21360_57480# diff_176040_194040# GND efet w=2460 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2058 diff_162960_208080# GND diff_165360_185160# GND efet w=2640 l=1080
+ ad=3.0672e+06 pd=9840 as=0 ps=0 
M2059 GND GND diff_162960_208080# GND efet w=660 l=5580
+ ad=0 pd=0 as=0 ps=0 
M2060 diff_148680_185160# GND GND GND efet w=480 l=5400
+ ad=0 pd=0 as=0 ps=0 
M2061 diff_180120_190560# GND diff_180360_194040# GND efet w=2820 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2062 GND GND diff_179760_181440# GND efet w=7140 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2063 GND GND diff_138120_220200# GND efet w=480 l=2880
+ ad=0 pd=0 as=1.6704e+07 ps=49680 
M2064 diff_133560_235080# diff_192240_207600# GND GND efet w=1800 l=840
+ ad=0 pd=0 as=0 ps=0 
M2065 GND GND diff_205680_198000# GND efet w=780 l=5460
+ ad=0 pd=0 as=2.232e+06 ps=8400 
M2066 GND GND diff_188880_226560# GND efet w=660 l=2100
+ ad=0 pd=0 as=5.6448e+06 ps=19200 
M2067 diff_188880_226560# diff_205680_198000# GND GND efet w=3120 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2068 diff_192240_207600# diff_193320_187440# GND GND efet w=1140 l=900
+ ad=0 pd=0 as=0 ps=0 
M2069 GND GND diff_192240_207600# GND efet w=1380 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2070 diff_205680_198000# diff_20640_113640# diff_205680_196560# GND efet w=2700 l=1020
+ ad=0 pd=0 as=1.9152e+06 ps=7920 
M2071 GND diff_201120_185760# diff_138120_220200# GND efet w=2100 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2072 diff_178920_94920# GND diff_183600_181920# GND efet w=1200 l=1080
+ ad=2.45664e+07 pd=64800 as=0 ps=0 
M2073 diff_206520_194880# GND diff_205680_196560# GND efet w=2520 l=960
+ ad=1.512e+06 pd=6240 as=0 ps=0 
M2074 diff_206520_194880# GND GND GND efet w=2340 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2075 diff_196920_186240# diff_20640_113640# GND GND efet w=2580 l=1020
+ ad=5.1696e+06 pd=18240 as=0 ps=0 
M2076 diff_97800_109440# GND GND GND efet w=2520 l=1260
+ ad=1.66176e+07 pd=60480 as=0 ps=0 
M2077 GND GND GND GND efet w=2520 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2078 GND GND GND GND efet w=4380 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2079 GND GND diff_69720_171360# GND efet w=3960 l=960
+ ad=0 pd=0 as=2.5992e+07 ps=82800 
M2080 GND GND GND GND efet w=2580 l=960
+ ad=0 pd=0 as=0 ps=0 
M2081 GND GND GND GND efet w=2520 l=900
+ ad=0 pd=0 as=0 ps=0 
M2082 GND GND GND GND efet w=2580 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2083 diff_51480_191880# GND GND GND efet w=4140 l=960
+ ad=2.05056e+07 pd=62880 as=0 ps=0 
M2084 GND GND GND GND efet w=2100 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2085 GND GND GND GND efet w=1980 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2086 diff_52080_163800# GND GND GND efet w=540 l=2940
+ ad=4.3056e+06 pd=18720 as=0 ps=0 
M2087 diff_44040_172320# diff_49320_172200# diff_44040_172320# GND efet w=5760 l=420
+ ad=0 pd=0 as=0 ps=0 
M2088 GND diff_47160_165840# GND GND efet w=2520 l=960
+ ad=0 pd=0 as=0 ps=0 
M2089 diff_44040_172320# diff_47160_165840# GND GND efet w=2400 l=960
+ ad=0 pd=0 as=0 ps=0 
M2090 GND GND diff_65520_142080# GND efet w=2040 l=960
+ ad=0 pd=0 as=1.2888e+07 ps=47520 
M2091 GND GND GND GND efet w=1980 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2092 GND GND diff_44520_186120# GND efet w=3720 l=960
+ ad=0 pd=0 as=2.24496e+07 ps=62640 
M2093 GND GND GND GND efet w=3660 l=960
+ ad=0 pd=0 as=0 ps=0 
M2094 GND GND diff_89160_121200# GND efet w=1920 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2095 diff_65520_142080# diff_69720_171360# GND GND efet w=2580 l=960
+ ad=0 pd=0 as=0 ps=0 
M2096 GND diff_69720_171360# GND GND efet w=2460 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2097 diff_82080_164400# diff_69720_171360# GND GND efet w=2580 l=960
+ ad=0 pd=0 as=0 ps=0 
M2098 GND diff_69720_171360# GND GND efet w=4620 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2099 GND GND GND GND efet w=1980 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2100 GND GND GND GND efet w=1920 l=960
+ ad=0 pd=0 as=0 ps=0 
M2101 GND GND GND GND efet w=2640 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2102 GND diff_11280_215400# diff_196920_186240# GND efet w=2460 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2103 diff_196920_186240# GND diff_195360_185760# GND efet w=2820 l=1140
+ ad=0 pd=0 as=1.584e+06 ps=7200 
M2104 GND GND diff_179760_181440# GND efet w=6780 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2105 GND diff_11280_215400# diff_183600_181920# GND efet w=4260 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2106 diff_183600_181920# GND GND GND efet w=3060 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2107 GND diff_178920_94920# diff_178920_94920# GND efet w=3960 l=1560
+ ad=0 pd=0 as=0 ps=0 
M2108 diff_178920_94920# diff_178920_94920# GND GND efet w=5040 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2109 diff_195360_185760# GND diff_193320_187440# GND efet w=2520 l=720
+ ad=0 pd=0 as=3.9024e+06 ps=15360 
M2110 GND GND diff_207360_188640# GND efet w=2460 l=900
+ ad=0 pd=0 as=2.0736e+06 ps=6720 
M2111 diff_207360_188640# GND diff_207360_187080# GND efet w=2460 l=900
+ ad=0 pd=0 as=1.7712e+06 ps=6480 
M2112 diff_203520_184560# diff_21360_57480# diff_201120_185760# GND efet w=1980 l=780
+ ad=1.152e+06 pd=5040 as=2.5344e+06 ps=10560 
M2113 GND GND diff_203520_184560# GND efet w=1920 l=960
+ ad=0 pd=0 as=0 ps=0 
M2114 diff_207360_187080# GND diff_207360_185520# GND efet w=2520 l=840
+ ad=0 pd=0 as=2.3616e+06 ps=9600 
M2115 diff_183600_181920# GND GND GND efet w=600 l=3120
+ ad=0 pd=0 as=0 ps=0 
M2116 GND GND diff_193320_187440# GND efet w=540 l=5340
+ ad=0 pd=0 as=0 ps=0 
M2117 GND GND GND GND efet w=3540 l=1500
+ ad=0 pd=0 as=0 ps=0 
M2118 diff_69720_171360# GND GND GND efet w=2940 l=1500
+ ad=0 pd=0 as=0 ps=0 
M2119 GND diff_69720_171360# diff_95160_164880# GND efet w=7620 l=900
+ ad=0 pd=0 as=1.46016e+07 ps=35280 
M2120 diff_89160_121200# diff_69720_171360# GND GND efet w=2520 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2121 GND diff_69720_171360# GND GND efet w=2520 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2122 diff_58200_162360# diff_51480_191880# diff_56040_162240# GND efet w=3000 l=1320
+ ad=1.04976e+07 pd=36960 as=9.4464e+06 ps=30000 
M2123 diff_56040_162240# GND diff_58200_162360# GND efet w=2760 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2124 GND diff_69720_171360# GND GND efet w=2640 l=960
+ ad=0 pd=0 as=0 ps=0 
M2125 GND GND GND GND efet w=2040 l=960
+ ad=0 pd=0 as=0 ps=0 
M2126 GND GND GND GND efet w=1980 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2127 GND diff_69720_171360# GND GND efet w=4680 l=960
+ ad=0 pd=0 as=0 ps=0 
M2128 diff_69720_171360# diff_69720_171360# GND GND efet w=3780 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2129 GND diff_69720_171360# GND GND efet w=2700 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2130 diff_95160_164880# GND diff_51480_191880# GND efet w=8160 l=960
+ ad=0 pd=0 as=0 ps=0 
M2131 GND GND GND GND efet w=1560 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2132 GND GND GND GND efet w=1740 l=1380
+ ad=0 pd=0 as=0 ps=0 
M2133 GND GND GND GND efet w=1680 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2134 GND diff_69720_171360# GND GND efet w=2700 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2135 GND GND diff_44520_186120# GND efet w=3720 l=840
+ ad=0 pd=0 as=0 ps=0 
M2136 GND GND GND GND efet w=2580 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2137 diff_65520_142080# GND GND GND efet w=2640 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2138 GND GND diff_97800_109440# GND efet w=1920 l=960
+ ad=0 pd=0 as=0 ps=0 
M2139 GND GND GND GND efet w=1740 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2140 GND GND GND GND efet w=3840 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2141 GND diff_173280_163200# GND GND efet w=3960 l=1680
+ ad=0 pd=0 as=0 ps=0 
M2142 GND GND diff_69720_171360# GND efet w=2760 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2143 diff_69720_171360# GND GND GND efet w=3000 l=1440
+ ad=0 pd=0 as=0 ps=0 
M2144 GND GND GND GND efet w=1860 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2145 GND GND GND GND efet w=2460 l=960
+ ad=0 pd=0 as=0 ps=0 
M2146 GND GND GND GND efet w=2460 l=960
+ ad=0 pd=0 as=0 ps=0 
M2147 diff_82080_164400# GND GND GND efet w=2520 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2148 diff_44520_186120# GND GND GND efet w=4440 l=960
+ ad=0 pd=0 as=0 ps=0 
M2149 diff_89160_121200# GND GND GND efet w=2460 l=900
+ ad=0 pd=0 as=0 ps=0 
M2150 diff_95160_164880# GND GND GND efet w=7380 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2151 diff_97800_109440# GND GND GND efet w=2520 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2152 GND GND GND GND efet w=1680 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2153 GND GND GND GND efet w=1620 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2154 GND GND GND GND efet w=1740 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2155 GND GND GND GND efet w=4740 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2156 GND GND diff_69720_171360# GND efet w=3780 l=960
+ ad=0 pd=0 as=0 ps=0 
M2157 diff_52080_163800# GND diff_47160_165840# GND efet w=1200 l=1080
+ ad=0 pd=0 as=2.1024e+06 ps=7200 
M2158 diff_56040_162240# GND GND GND efet w=3120 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2159 diff_43800_159360# GND GND GND efet w=660 l=5340
+ ad=979200 pd=6240 as=0 ps=0 
M2160 GND diff_52680_161880# diff_52080_163800# GND efet w=1860 l=900
+ ad=0 pd=0 as=0 ps=0 
M2161 diff_58200_162360# GND diff_56040_162240# GND efet w=2640 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2162 diff_51360_158880# GND diff_58200_162360# GND efet w=2880 l=960
+ ad=9.7488e+06 pd=31440 as=0 ps=0 
M2163 GND GND GND GND efet w=1980 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2164 GND GND GND GND efet w=3420 l=1500
+ ad=0 pd=0 as=0 ps=0 
M2165 GND GND GND GND efet w=1920 l=840
+ ad=0 pd=0 as=0 ps=0 
M2166 diff_95160_164880# GND diff_51480_191880# GND efet w=7980 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2167 GND GND GND GND efet w=1920 l=960
+ ad=0 pd=0 as=0 ps=0 
M2168 GND GND GND GND efet w=1800 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2169 GND GND diff_69720_171360# GND efet w=3540 l=1380
+ ad=0 pd=0 as=0 ps=0 
M2170 GND GND GND GND efet w=2520 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2171 GND GND GND GND efet w=2640 l=960
+ ad=0 pd=0 as=0 ps=0 
M2172 GND diff_173280_163200# diff_69720_171360# GND efet w=2700 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2173 GND GND GND GND efet w=2460 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2174 diff_178920_94920# GND GND GND efet w=840 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2175 GND diff_182760_168000# GND GND efet w=3240 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2176 GND diff_182160_172680# GND GND efet w=1680 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2177 GND GND diff_201120_185760# GND efet w=600 l=5040
+ ad=0 pd=0 as=0 ps=0 
M2178 diff_207360_185520# GND GND GND efet w=540 l=5220
+ ad=0 pd=0 as=0 ps=0 
M2179 GND diff_207360_185520# diff_209760_180360# GND efet w=3060 l=780
+ ad=0 pd=0 as=2.4768e+06 ps=10320 
M2180 diff_209760_180360# GND GND GND efet w=540 l=2160
+ ad=0 pd=0 as=0 ps=0 
M2181 GND diff_209760_180360# diff_191760_165240# GND efet w=960 l=1020
+ ad=0 pd=0 as=1.9152e+06 ps=6720 
M2182 GND diff_209760_180360# diff_197160_165000# GND efet w=900 l=960
+ ad=0 pd=0 as=1.8e+06 ps=6960 
M2183 GND diff_182160_172680# GND GND efet w=2460 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2184 GND diff_182760_168000# GND GND efet w=1680 l=960
+ ad=0 pd=0 as=0 ps=0 
M2185 GND GND GND GND efet w=720 l=2520
+ ad=0 pd=0 as=0 ps=0 
M2186 GND GND GND GND efet w=840 l=2700
+ ad=0 pd=0 as=0 ps=0 
M2187 GND diff_191760_165240# GND GND efet w=4860 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2188 GND diff_208440_168000# diff_182160_172680# GND efet w=5160 l=960
+ ad=0 pd=0 as=4.4784e+06 ps=20880 
M2189 GND diff_209760_180360# diff_202560_165000# GND efet w=900 l=1020
+ ad=0 pd=0 as=1.9008e+06 ps=6720 
M2190 diff_178200_154800# GND GND GND efet w=1020 l=2400
+ ad=3.96e+06 pd=16800 as=0 ps=0 
M2191 GND diff_197160_165000# GND GND efet w=5100 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2192 diff_182160_172680# GND GND GND efet w=720 l=2760
+ ad=0 pd=0 as=0 ps=0 
M2193 GND GND GND GND efet w=1980 l=900
+ ad=0 pd=0 as=0 ps=0 
M2194 GND GND GND GND efet w=1860 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2195 GND GND GND GND efet w=1800 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2196 diff_65520_142080# GND GND GND efet w=2640 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2197 GND GND GND GND efet w=2520 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2198 diff_82080_164400# GND GND GND efet w=2520 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2199 diff_44520_186120# GND GND GND efet w=4320 l=900
+ ad=0 pd=0 as=0 ps=0 
M2200 GND GND diff_43800_159360# GND efet w=1020 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2201 diff_49800_158880# diff_43800_159360# GND GND efet w=1800 l=960
+ ad=1.08e+06 pd=4800 as=0 ps=0 
M2202 diff_51360_158880# diff_47160_165840# diff_49800_158880# GND efet w=1800 l=960
+ ad=0 pd=0 as=0 ps=0 
M2203 diff_52680_161880# GND diff_51360_158880# GND efet w=720 l=960
+ ad=777600 pd=3600 as=0 ps=0 
M2204 diff_51360_158880# GND diff_51360_158880# GND efet w=300 l=5820
+ ad=0 pd=0 as=0 ps=0 
M2205 diff_97800_109440# GND GND GND efet w=2460 l=900
+ ad=0 pd=0 as=0 ps=0 
M2206 GND GND diff_51480_191880# GND efet w=4380 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2207 GND GND GND GND efet w=2580 l=840
+ ad=0 pd=0 as=0 ps=0 
M2208 GND GND GND GND efet w=1740 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2209 GND GND diff_69720_171360# GND efet w=4320 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2210 GND GND GND GND efet w=1980 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2211 GND GND GND GND efet w=2580 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2212 GND GND GND GND efet w=3300 l=1800
+ ad=0 pd=0 as=0 ps=0 
M2213 GND diff_66000_145440# GND GND efet w=1800 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2214 GND GND GND GND efet w=1800 l=1560
+ ad=0 pd=0 as=0 ps=0 
M2215 GND GND GND GND efet w=1680 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2216 GND GND diff_43560_137160# GND efet w=540 l=3300
+ ad=0 pd=0 as=2.2176e+06 ps=9600 
M2217 GND GND GND GND efet w=660 l=1860
+ ad=0 pd=0 as=0 ps=0 
M2218 diff_44520_147840# GND GND GND efet w=840 l=2340
+ ad=4.5072e+06 pd=15120 as=0 ps=0 
M2219 diff_43560_137160# diff_21360_45480# GND GND efet w=1500 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2220 GND GND GND GND efet w=480 l=4920
+ ad=0 pd=0 as=0 ps=0 
M2221 GND GND GND GND efet w=1560 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2222 GND diff_168480_155400# GND GND efet w=1680 l=1440
+ ad=0 pd=0 as=0 ps=0 
M2223 GND GND GND GND efet w=2040 l=840
+ ad=0 pd=0 as=0 ps=0 
M2224 GND GND GND GND efet w=1560 l=1380
+ ad=0 pd=0 as=0 ps=0 
M2225 diff_65520_142080# GND GND GND efet w=600 l=5280
+ ad=0 pd=0 as=0 ps=0 
M2226 GND GND GND GND efet w=480 l=5160
+ ad=0 pd=0 as=0 ps=0 
M2227 GND GND GND GND efet w=480 l=5220
+ ad=0 pd=0 as=0 ps=0 
M2228 GND GND GND GND efet w=780 l=6060
+ ad=0 pd=0 as=0 ps=0 
M2229 diff_55080_128160# GND GND GND efet w=600 l=6000
+ ad=3.312e+06 pd=12720 as=0 ps=0 
M2230 GND GND diff_82080_164400# GND efet w=600 l=4680
+ ad=0 pd=0 as=0 ps=0 
M2231 diff_44520_186120# GND GND GND efet w=600 l=3060
+ ad=0 pd=0 as=0 ps=0 
M2232 GND GND diff_84840_148440# GND efet w=600 l=4200
+ ad=0 pd=0 as=1.4976e+06 ps=7440 
M2233 GND GND GND GND efet w=720 l=3240
+ ad=0 pd=0 as=0 ps=0 
M2234 diff_51480_191880# GND GND GND efet w=720 l=2880
+ ad=0 pd=0 as=0 ps=0 
M2235 diff_89160_121200# GND GND GND efet w=600 l=4560
+ ad=0 pd=0 as=0 ps=0 
M2236 GND GND GND GND efet w=480 l=5280
+ ad=0 pd=0 as=0 ps=0 
M2237 GND diff_66000_145440# diff_74760_145920# GND efet w=3180 l=900
+ ad=0 pd=0 as=1.8144e+06 ps=7920 
M2238 diff_74760_145920# GND diff_57000_124920# GND efet w=1920 l=1080
+ ad=0 pd=0 as=5.112e+06 ps=19440 
M2239 GND GND diff_61320_143040# GND efet w=2760 l=840
+ ad=0 pd=0 as=1.8576e+06 ps=7200 
M2240 GND reset diff_41160_139680# GND efet w=2940 l=1020
+ ad=0 pd=0 as=6.696e+06 ps=20880 
M2241 GND GND diff_44520_147840# GND efet w=4260 l=1560
+ ad=0 pd=0 as=0 ps=0 
M2242 GND diff_41160_139680# diff_43560_137160# GND efet w=1620 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2243 GND diff_41160_139680# GND GND efet w=4620 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2244 diff_55320_141960# GND GND GND efet w=1800 l=1080
+ ad=1.728e+06 pd=7440 as=0 ps=0 
M2245 diff_55800_140760# GND GND GND efet w=1140 l=1020
+ ad=1.2096e+06 pd=7200 as=0 ps=0 
M2246 diff_61320_143040# GND diff_61320_141480# GND efet w=2820 l=900
+ ad=0 pd=0 as=1.8144e+06 ps=6480 
M2247 GND GND diff_55080_128160# GND efet w=1140 l=960
+ ad=0 pd=0 as=0 ps=0 
M2248 diff_84840_148440# diff_82080_164400# GND GND efet w=1260 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2249 GND diff_84840_148440# GND GND efet w=2400 l=960
+ ad=0 pd=0 as=0 ps=0 
M2250 GND GND diff_55080_128160# GND efet w=2880 l=960
+ ad=0 pd=0 as=0 ps=0 
M2251 diff_55080_128160# diff_55080_128160# GND GND efet w=660 l=1500
+ ad=0 pd=0 as=0 ps=0 
M2252 GND diff_65520_142080# diff_66000_140160# GND efet w=1080 l=960
+ ad=0 pd=0 as=2.736e+06 ps=7920 
M2253 GND GND diff_68400_139200# GND efet w=720 l=1440
+ ad=0 pd=0 as=2.8944e+06 ps=12240 
M2254 GND diff_82080_164400# GND GND efet w=2460 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2255 GND GND GND GND efet w=600 l=4440
+ ad=0 pd=0 as=0 ps=0 
M2256 GND GND GND GND efet w=480 l=5460
+ ad=0 pd=0 as=0 ps=0 
M2257 GND GND GND GND efet w=720 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2258 GND GND GND GND efet w=720 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2259 diff_97800_109440# GND GND GND efet w=480 l=4740
+ ad=0 pd=0 as=0 ps=0 
M2260 GND GND GND GND efet w=540 l=4740
+ ad=0 pd=0 as=0 ps=0 
M2261 GND GND GND GND efet w=600 l=4560
+ ad=0 pd=0 as=0 ps=0 
M2262 GND GND GND GND efet w=540 l=5040
+ ad=0 pd=0 as=0 ps=0 
M2263 GND GND GND GND efet w=840 l=5400
+ ad=0 pd=0 as=0 ps=0 
M2264 GND GND diff_106440_110160# GND efet w=480 l=4680
+ ad=0 pd=0 as=4.8096e+06 ps=15600 
M2265 GND GND diff_115920_125040# GND efet w=600 l=4560
+ ad=0 pd=0 as=8.9424e+06 ps=33120 
M2266 GND GND GND GND efet w=540 l=4560
+ ad=0 pd=0 as=0 ps=0 
M2267 GND GND GND GND efet w=540 l=4620
+ ad=0 pd=0 as=0 ps=0 
M2268 GND GND GND GND efet w=600 l=4680
+ ad=0 pd=0 as=0 ps=0 
M2269 GND GND GND GND efet w=480 l=5100
+ ad=0 pd=0 as=0 ps=0 
M2270 GND GND GND GND efet w=480 l=5400
+ ad=0 pd=0 as=0 ps=0 
M2271 GND GND GND GND efet w=540 l=5580
+ ad=0 pd=0 as=0 ps=0 
M2272 GND GND GND GND efet w=600 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2273 diff_106440_110160# diff_55080_128160# GND GND efet w=3180 l=900
+ ad=0 pd=0 as=0 ps=0 
M2274 GND GND GND GND efet w=600 l=4440
+ ad=0 pd=0 as=0 ps=0 
M2275 GND GND GND GND efet w=540 l=4380
+ ad=0 pd=0 as=0 ps=0 
M2276 GND GND GND GND efet w=480 l=4680
+ ad=0 pd=0 as=0 ps=0 
M2277 GND GND GND GND efet w=600 l=5220
+ ad=0 pd=0 as=0 ps=0 
M2278 GND GND GND GND efet w=600 l=5040
+ ad=0 pd=0 as=0 ps=0 
M2279 GND GND GND GND efet w=600 l=4920
+ ad=0 pd=0 as=0 ps=0 
M2280 GND GND GND GND efet w=660 l=4860
+ ad=0 pd=0 as=0 ps=0 
M2281 GND GND GND GND efet w=600 l=5280
+ ad=0 pd=0 as=0 ps=0 
M2282 GND GND GND GND efet w=660 l=5400
+ ad=0 pd=0 as=0 ps=0 
M2283 GND GND GND GND efet w=600 l=4680
+ ad=0 pd=0 as=0 ps=0 
M2284 GND GND GND GND efet w=480 l=4680
+ ad=0 pd=0 as=0 ps=0 
M2285 GND GND GND GND efet w=1740 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2286 GND diff_168480_155400# GND GND efet w=2460 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2287 GND diff_178200_154800# GND GND efet w=3180 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2288 GND diff_178200_162000# GND GND efet w=2040 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2289 diff_168480_155400# GND GND GND efet w=1800 l=1440
+ ad=3.9456e+06 pd=15600 as=0 ps=0 
M2290 GND diff_202560_165000# diff_178200_154800# GND efet w=4800 l=960
+ ad=0 pd=0 as=0 ps=0 
M2291 diff_173280_163200# GND GND GND efet w=1920 l=1440
+ ad=6.7392e+06 pd=21840 as=0 ps=0 
M2292 diff_178200_162000# diff_178200_154800# GND GND efet w=2400 l=840
+ ad=4.5072e+06 pd=14400 as=0 ps=0 
M2293 GND diff_209760_180360# diff_208440_168000# GND efet w=840 l=1020
+ ad=0 pd=0 as=1.8432e+06 ps=6480 
M2294 diff_182760_168000# diff_182160_172680# GND GND efet w=2220 l=900
+ ad=4.248e+06 pd=14880 as=0 ps=0 
M2295 diff_168480_155400# diff_189960_159840# diff_168480_155400# GND efet w=300 l=4260
+ ad=0 pd=0 as=0 ps=0 
M2296 GND diff_178200_162000# GND GND efet w=2820 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2297 GND diff_178200_154800# GND GND efet w=2040 l=960
+ ad=0 pd=0 as=0 ps=0 
M2298 diff_173280_163200# GND diff_173280_163200# GND efet w=360 l=4440
+ ad=0 pd=0 as=0 ps=0 
M2299 diff_178200_162000# GND diff_178200_162000# GND efet w=300 l=3540
+ ad=0 pd=0 as=0 ps=0 
M2300 diff_182760_168000# GND diff_182760_168000# GND efet w=240 l=4260
+ ad=0 pd=0 as=0 ps=0 
M2301 GND diff_165480_110160# GND GND efet w=4860 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2302 GND GND GND GND efet w=900 l=3420
+ ad=0 pd=0 as=0 ps=0 
M2303 GND diff_55080_128160# GND GND efet w=2640 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2304 GND diff_55080_128160# GND GND efet w=2640 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2305 GND GND diff_159360_93840# GND efet w=480 l=4080
+ ad=0 pd=0 as=4.536e+06 ps=15600 
M2306 GND diff_70080_105840# diff_178560_149760# GND efet w=1140 l=1020
+ ad=0 pd=0 as=2.1888e+06 ps=10080 
M2307 diff_178560_149760# GND GND GND efet w=600 l=5580
+ ad=0 pd=0 as=0 ps=0 
M2308 diff_183600_148680# diff_178560_149760# diff_159360_93840# GND efet w=2280 l=960
+ ad=1.2672e+06 pd=5760 as=0 ps=0 
M2309 diff_180360_148200# GND GND GND efet w=600 l=6420
+ ad=1.44e+06 pd=7440 as=0 ps=0 
M2310 diff_183600_148680# diff_180360_148200# GND GND efet w=2220 l=900
+ ad=0 pd=0 as=0 ps=0 
M2311 diff_180360_148200# GND GND GND efet w=780 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2312 diff_55320_141960# diff_55800_140760# diff_56400_140040# GND efet w=1680 l=960
+ ad=0 pd=0 as=4.9104e+06 ps=15600 
M2313 diff_61320_141480# diff_60720_140760# diff_56400_140040# GND efet w=2520 l=840
+ ad=0 pd=0 as=0 ps=0 
M2314 GND diff_43560_137160# diff_41160_139680# GND efet w=2760 l=960
+ ad=0 pd=0 as=0 ps=0 
M2315 diff_30000_135120# GND GND GND efet w=2160 l=960
+ ad=9.0576e+06 pd=34080 as=0 ps=0 
M2316 diff_30000_135120# diff_30720_135000# diff_30000_135120# GND efet w=6180 l=420
+ ad=0 pd=0 as=0 ps=0 
M2317 GND GND diff_26040_133800# GND efet w=900 l=1260
+ ad=0 pd=0 as=950400 ps=4800 
M2318 GND diff_30720_135000# diff_30000_135120# GND efet w=660 l=2700
+ ad=0 pd=0 as=0 ps=0 
M2319 GND GND diff_30720_135000# GND efet w=480 l=1080
+ ad=0 pd=0 as=316800 ps=2400 
M2320 GND diff_30000_135120# diff_27480_130800# GND efet w=2280 l=960
+ ad=0 pd=0 as=7.1712e+06 ps=23520 
M2321 diff_27480_130800# diff_26040_133800# GND GND efet w=5160 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2322 GND GND diff_27480_130800# GND efet w=660 l=1740
+ ad=0 pd=0 as=0 ps=0 
M2323 GND GND diff_27480_130800# GND efet w=960 l=960
+ ad=0 pd=0 as=0 ps=0 
M2324 diff_52440_136080# GND GND GND efet w=1200 l=960
+ ad=2.6496e+06 pd=9600 as=0 ps=0 
M2325 GND diff_53040_136920# diff_52440_136080# GND efet w=2220 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2326 diff_56400_140040# GND diff_53040_136920# GND efet w=720 l=960
+ ad=0 pd=0 as=979200 ps=5280 
M2327 GND GND diff_55800_140760# GND efet w=600 l=6960
+ ad=0 pd=0 as=0 ps=0 
M2328 GND test diff_42960_134880# GND efet w=3000 l=840
+ ad=0 pd=0 as=1.05984e+07 ps=34800 
M2329 GND GND diff_42960_134880# GND efet w=360 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2330 diff_41160_139680# GND GND GND efet w=480 l=2160
+ ad=0 pd=0 as=0 ps=0 
M2331 GND GND diff_52440_136080# GND efet w=600 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2332 GND GND diff_46320_121200# GND efet w=480 l=4200
+ ad=0 pd=0 as=2.3904e+06 ps=10320 
M2333 diff_27840_125040# GND GND GND efet w=2640 l=900
+ ad=7.8192e+06 pd=30000 as=0 ps=0 
M2334 GND GND GND GND efet w=720 l=1680
+ ad=0 pd=0 as=0 ps=0 
M2335 diff_56400_140040# GND GND GND efet w=540 l=5220
+ ad=0 pd=0 as=0 ps=0 
M2336 diff_66000_140160# GND GND GND efet w=900 l=5460
+ ad=0 pd=0 as=0 ps=0 
M2337 GND diff_68400_139200# diff_70560_140880# GND efet w=1920 l=960
+ ad=0 pd=0 as=1.48464e+07 ps=53760 
M2338 GND GND GND GND efet w=1620 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2339 GND GND GND GND efet w=1680 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2340 GND GND GND GND efet w=1980 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2341 GND GND GND GND efet w=3180 l=900
+ ad=0 pd=0 as=0 ps=0 
M2342 GND GND GND GND efet w=2820 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2343 diff_115920_125040# GND GND GND efet w=1980 l=900
+ ad=0 pd=0 as=0 ps=0 
M2344 GND GND GND GND efet w=1980 l=900
+ ad=0 pd=0 as=0 ps=0 
M2345 GND GND GND GND efet w=2040 l=960
+ ad=0 pd=0 as=0 ps=0 
M2346 diff_70560_140880# diff_75840_138120# diff_77400_140520# GND efet w=3660 l=1260
+ ad=0 pd=0 as=7.272e+06 ps=27360 
M2347 diff_70560_140880# GND diff_77400_140520# GND efet w=5280 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2348 diff_70560_140880# diff_66000_140160# diff_60720_140760# GND efet w=3420 l=1140
+ ad=0 pd=0 as=5.6448e+06 ps=15360 
M2349 GND diff_55080_128160# GND GND efet w=4920 l=960
+ ad=0 pd=0 as=0 ps=0 
M2350 diff_68400_139200# GND GND GND efet w=480 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2351 diff_70560_140880# diff_72120_132600# diff_60720_140760# GND efet w=3900 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2352 diff_60720_140760# GND GND GND efet w=480 l=4140
+ ad=0 pd=0 as=0 ps=0 
M2353 GND GND diff_57000_124920# GND efet w=480 l=5700
+ ad=0 pd=0 as=0 ps=0 
M2354 GND GND GND GND efet w=2520 l=900
+ ad=0 pd=0 as=0 ps=0 
M2355 GND GND GND GND efet w=2520 l=960
+ ad=0 pd=0 as=0 ps=0 
M2356 GND GND GND GND efet w=3360 l=960
+ ad=0 pd=0 as=0 ps=0 
M2357 GND GND GND GND efet w=3360 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2358 GND GND diff_77400_140520# GND efet w=3840 l=1560
+ ad=0 pd=0 as=0 ps=0 
M2359 GND GND diff_77400_140520# GND efet w=6240 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2360 GND GND GND GND efet w=1560 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2361 GND GND GND GND efet w=1620 l=1380
+ ad=0 pd=0 as=0 ps=0 
M2362 GND GND GND GND efet w=1620 l=1380
+ ad=0 pd=0 as=0 ps=0 
M2363 GND GND GND GND efet w=1560 l=1440
+ ad=0 pd=0 as=0 ps=0 
M2364 GND GND GND GND efet w=1620 l=1380
+ ad=0 pd=0 as=0 ps=0 
M2365 GND diff_55080_128160# GND GND efet w=3300 l=900
+ ad=0 pd=0 as=0 ps=0 
M2366 diff_159360_93840# diff_21360_45480# diff_168960_143880# GND efet w=2640 l=960
+ ad=0 pd=0 as=2.2752e+06 ps=8400 
M2367 GND diff_165480_110160# GND GND efet w=5100 l=1380
+ ad=0 pd=0 as=0 ps=0 
M2368 GND GND diff_168960_143880# GND efet w=2400 l=1440
+ ad=0 pd=0 as=0 ps=0 
M2369 GND GND GND GND efet w=1620 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2370 GND GND GND GND efet w=1620 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2371 GND GND GND GND efet w=2580 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2372 GND GND GND GND efet w=2460 l=960
+ ad=0 pd=0 as=0 ps=0 
M2373 GND GND GND GND efet w=2700 l=960
+ ad=0 pd=0 as=0 ps=0 
M2374 GND GND GND GND efet w=2520 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2375 GND GND GND GND efet w=3420 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2376 GND diff_172560_117720# GND GND efet w=2460 l=960
+ ad=0 pd=0 as=0 ps=0 
M2377 GND GND GND GND efet w=4680 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2378 GND GND GND GND efet w=1620 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2379 GND GND diff_106440_110160# GND efet w=2640 l=840
+ ad=0 pd=0 as=0 ps=0 
M2380 GND GND diff_115920_125040# GND efet w=2040 l=840
+ ad=0 pd=0 as=0 ps=0 
M2381 GND GND GND GND efet w=1980 l=900
+ ad=0 pd=0 as=0 ps=0 
M2382 GND GND GND GND efet w=1920 l=840
+ ad=0 pd=0 as=0 ps=0 
M2383 GND GND GND GND efet w=1920 l=840
+ ad=0 pd=0 as=0 ps=0 
M2384 GND GND GND GND efet w=2040 l=960
+ ad=0 pd=0 as=0 ps=0 
M2385 GND GND GND GND efet w=1620 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2386 GND GND diff_75840_138120# GND efet w=1080 l=960
+ ad=0 pd=0 as=2.2176e+06 ps=10560 
M2387 GND diff_89400_137160# GND GND efet w=2520 l=900
+ ad=0 pd=0 as=0 ps=0 
M2388 GND GND diff_84120_135360# GND efet w=3720 l=1200
+ ad=0 pd=0 as=3.8736e+06 ps=12240 
M2389 diff_84120_135360# diff_76560_120480# GND GND efet w=2400 l=900
+ ad=0 pd=0 as=0 ps=0 
M2390 diff_75840_138120# GND GND GND efet w=480 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2391 GND GND diff_64680_127080# GND efet w=540 l=2160
+ ad=0 pd=0 as=5.04e+06 ps=20640 
M2392 GND diff_89400_137160# GND GND efet w=2520 l=900
+ ad=0 pd=0 as=0 ps=0 
M2393 diff_115920_125040# diff_89400_137160# GND GND efet w=2640 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2394 GND diff_89400_137160# GND GND efet w=2580 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2395 GND GND GND GND efet w=1560 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2396 GND GND GND GND efet w=1680 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2397 GND diff_89400_137160# GND GND efet w=2520 l=960
+ ad=0 pd=0 as=0 ps=0 
M2398 GND diff_89400_137160# GND GND efet w=2580 l=960
+ ad=0 pd=0 as=0 ps=0 
M2399 GND GND GND GND efet w=480 l=3960
+ ad=0 pd=0 as=0 ps=0 
M2400 GND GND GND GND efet w=2580 l=1380
+ ad=0 pd=0 as=0 ps=0 
M2401 GND GND GND GND efet w=2520 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2402 GND diff_183360_117720# diff_89400_137160# GND efet w=3060 l=1260
+ ad=0 pd=0 as=5.6448e+06 ps=18720 
M2403 GND GND GND GND efet w=4020 l=1800
+ ad=0 pd=0 as=0 ps=0 
M2404 GND GND GND GND efet w=1860 l=900
+ ad=0 pd=0 as=0 ps=0 
M2405 GND diff_172560_117720# GND GND efet w=2100 l=780
+ ad=0 pd=0 as=0 ps=0 
M2406 GND GND GND GND efet w=1620 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2407 GND GND GND GND efet w=1800 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2408 GND GND GND GND efet w=1860 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2409 GND GND GND GND efet w=2100 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2410 GND GND GND GND efet w=2100 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2411 GND GND GND GND efet w=1500 l=1500
+ ad=0 pd=0 as=0 ps=0 
M2412 GND diff_102000_133320# GND GND efet w=3600 l=900
+ ad=0 pd=0 as=0 ps=0 
M2413 GND GND diff_64680_127080# GND efet w=3960 l=840
+ ad=0 pd=0 as=0 ps=0 
M2414 GND GND diff_41160_121200# GND efet w=540 l=5580
+ ad=0 pd=0 as=1.10016e+07 ps=39840 
M2415 diff_27840_125040# diff_28560_123960# diff_27840_125040# GND efet w=6000 l=480
+ ad=0 pd=0 as=0 ps=0 
M2416 GND diff_28560_123960# diff_27840_125040# GND efet w=540 l=2220
+ ad=0 pd=0 as=0 ps=0 
M2417 GND GND diff_28560_123960# GND efet w=480 l=1080
+ ad=0 pd=0 as=360000 ps=2880 
M2418 GND GND GND GND efet w=2580 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2419 GND diff_41160_121200# diff_46320_121200# GND efet w=1200 l=960
+ ad=0 pd=0 as=0 ps=0 
M2420 GND diff_27840_125040# GND GND efet w=3000 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2421 diff_71040_129240# GND diff_21360_57480# GND efet w=720 l=960
+ ad=475200 pd=2880 as=9.58032e+07 ps=246960 
M2422 diff_41160_121200# diff_57000_124920# GND GND efet w=1080 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2423 diff_70080_125040# diff_71040_129240# GND GND efet w=1200 l=960
+ ad=3.2688e+06 pd=12960 as=0 ps=0 
M2424 diff_70080_125040# diff_64680_127080# diff_67080_124440# GND efet w=720 l=1080
+ ad=0 pd=0 as=1.1808e+06 ps=5760 
M2425 GND GND diff_74160_129960# GND efet w=540 l=960
+ ad=0 pd=0 as=2.2032e+06 ps=8880 
M2426 GND diff_74160_129960# GND GND efet w=480 l=1380
+ ad=0 pd=0 as=0 ps=0 
M2427 GND diff_74160_129960# GND GND efet w=5760 l=2220
+ ad=0 pd=0 as=0 ps=0 
M2428 diff_84000_131040# diff_55200_81120# GND GND efet w=2280 l=960
+ ad=3.168e+06 pd=12960 as=0 ps=0 
M2429 diff_115920_125040# diff_102000_133320# GND GND efet w=2580 l=840
+ ad=0 pd=0 as=0 ps=0 
M2430 GND diff_102000_133320# GND GND efet w=2520 l=960
+ ad=0 pd=0 as=0 ps=0 
M2431 GND GND diff_84000_131040# GND efet w=3780 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2432 GND diff_102000_133320# GND GND efet w=2640 l=960
+ ad=0 pd=0 as=0 ps=0 
M2433 GND diff_102000_133320# GND GND efet w=2580 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2434 GND diff_102000_133320# GND GND efet w=2640 l=960
+ ad=0 pd=0 as=0 ps=0 
M2435 GND GND GND GND efet w=2340 l=900
+ ad=0 pd=0 as=0 ps=0 
M2436 GND GND GND GND efet w=1800 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2437 GND diff_102000_133320# GND GND efet w=2460 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2438 GND diff_41160_121200# GND GND efet w=1680 l=960
+ ad=0 pd=0 as=0 ps=0 
M2439 GND diff_46320_121200# GND GND efet w=1680 l=960
+ ad=0 pd=0 as=0 ps=0 
M2440 diff_52200_120960# diff_43560_89160# diff_41160_121200# GND efet w=2520 l=840
+ ad=1.368e+06 pd=5760 as=0 ps=0 
M2441 GND GND diff_52200_120960# GND efet w=2280 l=960
+ ad=0 pd=0 as=0 ps=0 
M2442 diff_56040_120960# diff_45720_111480# GND GND efet w=2280 l=960
+ ad=3.6864e+06 pd=12960 as=0 ps=0 
M2443 diff_41160_121200# diff_41160_121200# diff_56040_120960# GND efet w=1980 l=1500
+ ad=0 pd=0 as=0 ps=0 
M2444 GND diff_60720_122640# diff_41160_121200# GND efet w=1260 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2445 GND GND diff_65040_121200# GND efet w=1380 l=1020
+ ad=0 pd=0 as=6.1344e+06 ps=25440 
M2446 diff_60720_122640# diff_67080_124440# GND GND efet w=1680 l=1020
+ ad=2.0016e+06 pd=7680 as=0 ps=0 
M2447 GND GND diff_60720_122640# GND efet w=660 l=4560
+ ad=0 pd=0 as=0 ps=0 
M2448 GND diff_27840_112800# GND GND efet w=3240 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2449 GND diff_24000_117480# GND GND efet w=3060 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2450 GND GND diff_20640_113640# GND efet w=2100 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2451 diff_27840_112800# diff_24000_117480# GND GND efet w=2520 l=960
+ ad=8.0064e+06 pd=28320 as=0 ps=0 
M2452 diff_27840_112800# diff_28560_113400# diff_27840_112800# GND efet w=5820 l=480
+ ad=0 pd=0 as=0 ps=0 
M2453 GND GND diff_28560_113400# GND efet w=540 l=1140
+ ad=0 pd=0 as=244800 ps=2160 
M2454 GND diff_28560_113400# diff_27840_112800# GND efet w=600 l=2280
+ ad=0 pd=0 as=0 ps=0 
M2455 diff_30240_108840# diff_27960_108600# GND GND efet w=2220 l=900
+ ad=4.7952e+06 pd=17520 as=0 ps=0 
M2456 diff_27960_108600# GND diff_20640_113640# GND efet w=1080 l=1140
+ ad=1.1232e+06 pd=5040 as=0 ps=0 
M2457 diff_24000_117480# GND diff_30240_108840# GND efet w=1200 l=960
+ ad=993600 pd=5040 as=0 ps=0 
M2458 GND GND diff_30240_108840# GND efet w=720 l=3120
+ ad=0 pd=0 as=0 ps=0 
M2459 diff_63480_120120# GND GND GND efet w=1200 l=960
+ ad=1.7856e+06 pd=7920 as=0 ps=0 
M2460 diff_41160_121200# diff_54720_116400# diff_41160_121200# GND efet w=1320 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2461 diff_20640_113640# diff_20640_113640# GND GND efet w=1500 l=1440
+ ad=0 pd=0 as=0 ps=0 
M2462 GND GND diff_20640_113640# GND efet w=2340 l=1620
+ ad=0 pd=0 as=0 ps=0 
M2463 diff_20640_113640# diff_24120_105360# GND GND efet w=3060 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2464 GND diff_28560_101520# GND GND efet w=6240 l=480
+ ad=0 pd=0 as=0 ps=0 
M2465 GND diff_24120_105360# GND GND efet w=2160 l=900
+ ad=0 pd=0 as=0 ps=0 
M2466 GND GND diff_28560_101520# GND efet w=480 l=960
+ ad=0 pd=0 as=316800 ps=2400 
M2467 GND diff_28560_101520# GND GND efet w=660 l=2220
+ ad=0 pd=0 as=0 ps=0 
M2468 GND diff_54720_116400# diff_41160_121200# GND efet w=480 l=3300
+ ad=0 pd=0 as=0 ps=0 
M2469 diff_65160_119400# GND diff_63480_120120# GND efet w=720 l=960
+ ad=403200 pd=2640 as=0 ps=0 
M2470 GND GND diff_70080_125040# GND efet w=480 l=4080
+ ad=0 pd=0 as=0 ps=0 
M2471 GND GND GND GND efet w=1620 l=1500
+ ad=0 pd=0 as=0 ps=0 
M2472 GND GND GND GND efet w=2100 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2473 GND GND GND GND efet w=2580 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2474 GND GND GND GND efet w=1680 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2475 GND GND GND GND efet w=1680 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2476 GND GND GND GND efet w=1560 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2477 GND GND GND GND efet w=1680 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2478 GND GND GND GND efet w=2040 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2479 GND GND GND GND efet w=1620 l=1440
+ ad=0 pd=0 as=0 ps=0 
M2480 diff_86760_128040# diff_42960_134880# GND GND efet w=2280 l=960
+ ad=3.6e+06 pd=13920 as=0 ps=0 
M2481 GND diff_66000_145440# diff_86760_128040# GND efet w=4080 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2482 GND diff_89400_129240# GND GND efet w=2520 l=960
+ ad=0 pd=0 as=0 ps=0 
M2483 GND diff_89400_129240# GND GND efet w=3480 l=900
+ ad=0 pd=0 as=0 ps=0 
M2484 GND diff_89400_129240# GND GND efet w=3420 l=960
+ ad=0 pd=0 as=0 ps=0 
M2485 GND diff_89400_129240# GND GND efet w=2580 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2486 GND diff_89400_129240# GND GND efet w=2520 l=960
+ ad=0 pd=0 as=0 ps=0 
M2487 GND diff_89400_129240# GND GND efet w=2640 l=960
+ ad=0 pd=0 as=0 ps=0 
M2488 GND diff_89400_129240# GND GND efet w=2580 l=840
+ ad=0 pd=0 as=0 ps=0 
M2489 GND diff_89400_129240# GND GND efet w=2460 l=960
+ ad=0 pd=0 as=0 ps=0 
M2490 GND diff_66000_145440# GND GND efet w=2040 l=840
+ ad=0 pd=0 as=0 ps=0 
M2491 GND diff_66000_145440# diff_115920_125040# GND efet w=2040 l=960
+ ad=0 pd=0 as=0 ps=0 
M2492 GND diff_66000_145440# GND GND efet w=2160 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2493 GND GND diff_89400_137160# GND efet w=1200 l=960
+ ad=0 pd=0 as=0 ps=0 
M2494 GND GND GND GND efet w=5700 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2495 GND diff_66000_145440# GND GND efet w=1920 l=960
+ ad=0 pd=0 as=0 ps=0 
M2496 GND diff_66000_145440# GND GND efet w=1920 l=900
+ ad=0 pd=0 as=0 ps=0 
M2497 GND diff_66000_145440# GND GND efet w=1920 l=840
+ ad=0 pd=0 as=0 ps=0 
M2498 GND diff_66000_145440# GND GND efet w=2040 l=960
+ ad=0 pd=0 as=0 ps=0 
M2499 GND diff_66000_145440# GND GND efet w=2040 l=840
+ ad=0 pd=0 as=0 ps=0 
M2500 GND GND GND GND efet w=3660 l=900
+ ad=0 pd=0 as=0 ps=0 
M2501 GND diff_84120_123480# diff_44280_73320# GND efet w=1860 l=900
+ ad=0 pd=0 as=3.08016e+07 ps=84960 
M2502 diff_44280_73320# GND GND GND efet w=1680 l=960
+ ad=0 pd=0 as=0 ps=0 
M2503 GND GND diff_84120_123480# GND efet w=1200 l=840
+ ad=0 pd=0 as=2.1168e+06 ps=10560 
M2504 diff_98880_123960# GND GND GND efet w=1200 l=840
+ ad=2.69136e+07 pd=102480 as=0 ps=0 
M2505 GND GND GND GND efet w=3660 l=900
+ ad=0 pd=0 as=0 ps=0 
M2506 GND GND diff_63480_120120# GND efet w=480 l=3960
+ ad=0 pd=0 as=0 ps=0 
M2507 diff_65040_121200# diff_65160_119400# GND GND efet w=1800 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2508 GND GND diff_70080_105840# GND efet w=480 l=1320
+ ad=0 pd=0 as=1.25712e+07 ps=41280 
M2509 diff_84120_123480# GND GND GND efet w=540 l=5340
+ ad=0 pd=0 as=0 ps=0 
M2510 GND GND diff_98880_123960# GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M2511 diff_98880_123960# GND GND GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M2512 diff_54720_116400# GND GND GND efet w=480 l=960
+ ad=820800 pd=4560 as=0 ps=0 
M2513 GND GND GND GND efet w=540 l=1560
+ ad=0 pd=0 as=0 ps=0 
M2514 diff_70080_105840# diff_65040_121200# GND GND efet w=5400 l=960
+ ad=0 pd=0 as=0 ps=0 
M2515 diff_65040_121200# GND GND GND efet w=480 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2516 diff_49560_105120# GND GND GND efet w=480 l=4680
+ ad=3.3264e+06 pd=15600 as=0 ps=0 
M2517 diff_54240_108720# GND GND GND efet w=480 l=2400
+ ad=6.2928e+06 pd=22560 as=0 ps=0 
M2518 GND GND diff_60720_104520# GND efet w=540 l=5340
+ ad=0 pd=0 as=6.4224e+06 ps=26880 
M2519 diff_30240_96720# diff_27960_96720# GND GND efet w=2220 l=900
+ ad=4.7664e+06 pd=16800 as=0 ps=0 
M2520 diff_27960_96720# GND diff_20640_113640# GND efet w=1320 l=960
+ ad=1.2096e+06 pd=5040 as=0 ps=0 
M2521 diff_24120_105360# GND diff_30240_96720# GND efet w=1200 l=960
+ ad=1.1232e+06 pd=5040 as=0 ps=0 
M2522 GND GND diff_30240_96720# GND efet w=600 l=2520
+ ad=0 pd=0 as=0 ps=0 
M2523 diff_54240_108720# diff_51120_105120# GND GND efet w=2880 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2524 GND GND diff_54240_108720# GND efet w=1800 l=1560
+ ad=0 pd=0 as=0 ps=0 
M2525 GND diff_54240_108720# GND GND efet w=4440 l=960
+ ad=0 pd=0 as=0 ps=0 
M2526 GND GND diff_60720_104520# GND efet w=840 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2527 diff_60720_104520# GND GND GND efet w=960 l=960
+ ad=0 pd=0 as=0 ps=0 
M2528 diff_55200_105000# GND GND GND efet w=2400 l=1080
+ ad=1.44e+06 pd=6000 as=0 ps=0 
M2529 GND GND diff_55200_105000# GND efet w=2460 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2530 diff_49560_105120# diff_20640_113640# GND GND efet w=1260 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2531 diff_51120_105120# GND diff_49560_105120# GND efet w=780 l=1020
+ ad=792000 pd=4320 as=0 ps=0 
M2532 diff_58440_105000# GND GND GND efet w=2580 l=1020
+ ad=1.5984e+06 pd=6720 as=0 ps=0 
M2533 diff_60000_105000# diff_54240_108720# diff_58440_105000# GND efet w=2580 l=900
+ ad=1.6848e+06 pd=6240 as=0 ps=0 
M2534 diff_58800_94080# diff_60720_104520# diff_60000_105000# GND efet w=2460 l=1020
+ ad=1.35792e+07 pd=64080 as=0 ps=0 
M2535 GND GND diff_58800_94080# GND efet w=2280 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2536 GND GND diff_46680_91560# GND efet w=1800 l=1080
+ ad=0 pd=0 as=4.1904e+06 ps=13680 
M2537 diff_58800_94080# GND GND GND efet w=2400 l=960
+ ad=0 pd=0 as=0 ps=0 
M2538 diff_44280_73320# GND GND GND efet w=600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2539 GND diff_89160_121200# diff_87480_109680# GND efet w=1320 l=840
+ ad=0 pd=0 as=1.728e+06 ps=6240 
M2540 diff_87480_109680# GND GND GND efet w=540 l=4860
+ ad=0 pd=0 as=0 ps=0 
M2541 GND GND GND GND efet w=960 l=960
+ ad=0 pd=0 as=0 ps=0 
M2542 GND GND diff_99120_118920# GND efet w=1020 l=1020
+ ad=0 pd=0 as=7.128e+06 ps=30240 
M2543 diff_104880_119520# GND GND GND efet w=1080 l=960
+ ad=1.20672e+07 pd=49680 as=0 ps=0 
M2544 GND diff_94440_117120# diff_91800_105960# GND efet w=6300 l=900
+ ad=0 pd=0 as=1.476e+07 ps=46800 
M2545 GND diff_58800_94080# GND GND efet w=1740 l=960
+ ad=0 pd=0 as=0 ps=0 
M2546 GND GND diff_46680_91560# GND efet w=540 l=2580
+ ad=0 pd=0 as=0 ps=0 
M2547 GND diff_20640_113640# diff_20640_113640# GND efet w=1440 l=1560
+ ad=0 pd=0 as=0 ps=0 
M2548 GND diff_27840_93120# diff_20640_113640# GND efet w=3360 l=960
+ ad=0 pd=0 as=0 ps=0 
M2549 diff_20640_113640# diff_24120_93360# GND GND efet w=2880 l=960
+ ad=0 pd=0 as=0 ps=0 
M2550 diff_27840_93120# diff_28560_89520# diff_27840_93120# GND efet w=5820 l=480
+ ad=7.7184e+06 pd=28080 as=0 ps=0 
M2551 diff_27840_93120# diff_24120_93360# GND GND efet w=2280 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2552 GND GND diff_28560_89520# GND efet w=480 l=960
+ ad=0 pd=0 as=460800 ps=2880 
M2553 GND diff_28560_89520# diff_27840_93120# GND efet w=360 l=2580
+ ad=0 pd=0 as=0 ps=0 
M2554 GND GND diff_47760_87000# GND efet w=480 l=4080
+ ad=0 pd=0 as=4.32e+06 ps=17280 
M2555 diff_58680_100920# GND diff_58680_100920# GND efet w=360 l=6240
+ ad=2.8368e+06 pd=10560 as=0 ps=0 
M2556 diff_47760_87000# diff_46680_91560# diff_45240_90120# GND efet w=840 l=900
+ ad=0 pd=0 as=403200 ps=3360 
M2557 diff_30240_84720# diff_28080_84600# GND GND efet w=2220 l=900
+ ad=4.6512e+06 pd=17520 as=0 ps=0 
M2558 diff_28080_84600# GND GND GND efet w=1140 l=1260
+ ad=1.1088e+06 pd=4800 as=0 ps=0 
M2559 diff_24120_93360# GND diff_30240_84720# GND efet w=1200 l=960
+ ad=1.0944e+06 pd=5520 as=0 ps=0 
M2560 GND GND diff_48240_86520# GND efet w=720 l=1020
+ ad=0 pd=0 as=432000 ps=3120 
M2561 GND diff_58680_100920# GND GND efet w=1680 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2562 GND diff_58800_94080# diff_58680_100920# GND efet w=960 l=960
+ ad=0 pd=0 as=0 ps=0 
M2563 GND diff_59040_94320# diff_58800_94080# GND efet w=540 l=4380
+ ad=0 pd=0 as=0 ps=0 
M2564 diff_59040_94320# GND GND GND efet w=540 l=1020
+ ad=950400 pd=5280 as=0 ps=0 
M2565 diff_58800_94080# diff_59040_94320# diff_58800_94080# GND efet w=5820 l=420
+ ad=0 pd=0 as=0 ps=0 
M2566 GND GND diff_45720_111480# GND efet w=960 l=4500
+ ad=0 pd=0 as=2.66688e+07 ps=81840 
M2567 GND GND GND GND efet w=300 l=5940
+ ad=0 pd=0 as=0 ps=0 
M2568 diff_20640_113640# GND diff_66480_87720# GND efet w=660 l=1080
+ ad=0 pd=0 as=950400 ps=4560 
M2569 diff_62160_91320# GND GND GND efet w=480 l=4680
+ ad=5.328e+06 pd=17280 as=0 ps=0 
M2570 diff_62160_91320# diff_46680_91560# GND GND efet w=900 l=900
+ ad=0 pd=0 as=0 ps=0 
M2571 GND GND diff_45720_111480# GND efet w=2220 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2572 GND diff_20640_113640# GND GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M2573 GND diff_48240_86520# diff_47760_87000# GND efet w=1260 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2574 GND diff_66480_87720# diff_62160_91320# GND efet w=1260 l=900
+ ad=0 pd=0 as=0 ps=0 
M2575 diff_43560_89160# GND GND GND efet w=540 l=4260
+ ad=9.2448e+06 pd=33600 as=0 ps=0 
M2576 GND GND diff_30240_84720# GND efet w=660 l=3180
+ ad=0 pd=0 as=0 ps=0 
M2577 GND diff_45240_90120# diff_43560_89160# GND efet w=1980 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2578 diff_20640_113640# GND GND GND efet w=1800 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2579 GND GND GND GND efet w=2880 l=2160
+ ad=0 pd=0 as=0 ps=0 
M2580 GND diff_56400_79440# GND GND efet w=2040 l=840
+ ad=0 pd=0 as=0 ps=0 
M2581 GND diff_24120_80040# GND GND efet w=3180 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2582 GND diff_41040_77520# GND GND efet w=5460 l=600
+ ad=0 pd=0 as=0 ps=0 
M2583 GND GND GND GND efet w=5820 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2584 GND diff_41040_77520# GND GND efet w=840 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2585 GND diff_28560_76560# GND GND efet w=6480 l=720
+ ad=0 pd=0 as=0 ps=0 
M2586 GND diff_62400_80640# GND GND efet w=1800 l=960
+ ad=0 pd=0 as=0 ps=0 
M2587 GND GND diff_91800_105960# GND efet w=6120 l=960
+ ad=0 pd=0 as=0 ps=0 
M2588 GND diff_97800_109440# diff_98880_123960# GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M2589 diff_98880_123960# GND GND GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M2590 diff_108000_115920# diff_89160_121200# GND GND efet w=960 l=1020
+ ad=4.1904e+06 pd=16080 as=0 ps=0 
M2591 GND GND GND GND efet w=1200 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2592 GND GND diff_98880_123960# GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M2593 diff_98880_123960# GND GND GND efet w=1140 l=900
+ ad=0 pd=0 as=0 ps=0 
M2594 GND GND diff_98880_123960# GND efet w=960 l=840
+ ad=0 pd=0 as=0 ps=0 
M2595 diff_98880_123960# GND GND GND efet w=960 l=840
+ ad=0 pd=0 as=0 ps=0 
M2596 GND diff_177960_117720# diff_102000_133320# GND efet w=2820 l=1260
+ ad=0 pd=0 as=4.4928e+06 ps=17040 
M2597 diff_98880_123960# GND GND GND efet w=1020 l=900
+ ad=0 pd=0 as=0 ps=0 
M2598 GND GND diff_102000_133320# GND efet w=2520 l=2160
+ ad=0 pd=0 as=0 ps=0 
M2599 GND diff_177960_117720# GND GND efet w=2220 l=1380
+ ad=0 pd=0 as=0 ps=0 
M2600 GND GND diff_98880_123960# GND efet w=1200 l=960
+ ad=0 pd=0 as=0 ps=0 
M2601 diff_98880_123960# GND GND GND efet w=1260 l=900
+ ad=0 pd=0 as=0 ps=0 
M2602 GND GND diff_98880_123960# GND efet w=1140 l=900
+ ad=0 pd=0 as=0 ps=0 
M2603 diff_98880_123960# GND GND GND efet w=1140 l=900
+ ad=0 pd=0 as=0 ps=0 
M2604 GND GND GND GND efet w=1380 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2605 GND GND GND GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M2606 GND GND GND GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M2607 GND GND GND GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M2608 GND GND GND GND efet w=1140 l=960
+ ad=0 pd=0 as=0 ps=0 
M2609 GND GND GND GND efet w=1260 l=900
+ ad=0 pd=0 as=0 ps=0 
M2610 GND GND GND GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M2611 GND GND GND GND efet w=1140 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2612 GND GND GND GND efet w=1080 l=840
+ ad=0 pd=0 as=0 ps=0 
M2613 GND GND GND GND efet w=1140 l=840
+ ad=0 pd=0 as=0 ps=0 
M2614 GND diff_115920_125040# diff_104880_119520# GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M2615 diff_104880_119520# GND GND GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M2616 diff_91800_105960# diff_94440_111840# diff_90000_47280# GND efet w=6180 l=900
+ ad=0 pd=0 as=2.81232e+07 ps=78720 
M2617 diff_90000_47280# diff_70080_105840# diff_91800_105960# GND efet w=6300 l=900
+ ad=0 pd=0 as=0 ps=0 
M2618 GND diff_87480_109680# diff_87360_101640# GND efet w=3240 l=1020
+ ad=0 pd=0 as=1.96704e+07 ps=65520 
M2619 GND diff_97800_109440# diff_94440_111840# GND efet w=1800 l=960
+ ad=0 pd=0 as=1.9152e+06 ps=9600 
M2620 GND diff_94440_117120# diff_97440_92520# GND efet w=1200 l=960
+ ad=0 pd=0 as=4.3056e+06 ps=14160 
M2621 GND diff_106440_110160# diff_94440_117120# GND efet w=1800 l=960
+ ad=0 pd=0 as=3.24e+06 ps=13440 
M2622 diff_99120_118920# GND GND GND efet w=1080 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2623 diff_104880_119520# GND GND GND efet w=1020 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2624 GND GND diff_104880_119520# GND efet w=1020 l=900
+ ad=0 pd=0 as=0 ps=0 
M2625 GND GND diff_104880_119520# GND efet w=960 l=840
+ ad=0 pd=0 as=0 ps=0 
M2626 GND diff_131760_114840# GND GND efet w=5400 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2627 GND GND diff_108000_115920# GND efet w=960 l=960
+ ad=0 pd=0 as=0 ps=0 
M2628 diff_111720_106680# GND GND GND efet w=1260 l=900
+ ad=3.0528e+06 pd=12480 as=0 ps=0 
M2629 diff_97440_92520# diff_70080_105840# GND GND efet w=1320 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2630 GND GND GND GND efet w=1980 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2631 GND diff_131760_114840# GND GND efet w=480 l=3360
+ ad=0 pd=0 as=0 ps=0 
M2632 diff_108000_115920# GND GND GND efet w=1200 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2633 diff_108000_115920# GND GND GND efet w=600 l=5520
+ ad=0 pd=0 as=0 ps=0 
M2634 diff_104880_119520# GND GND GND efet w=600 l=5760
+ ad=0 pd=0 as=0 ps=0 
M2635 GND diff_115920_125040# diff_117480_108840# GND efet w=1260 l=1260
+ ad=0 pd=0 as=3.7152e+06 ps=15600 
M2636 GND diff_70080_105840# diff_110280_107400# GND efet w=1440 l=900
+ ad=0 pd=0 as=4.5216e+06 ps=15600 
M2637 GND diff_70080_105840# diff_87360_101640# GND efet w=3180 l=900
+ ad=0 pd=0 as=0 ps=0 
M2638 diff_87360_101640# diff_86760_94560# diff_87360_101640# GND efet w=6960 l=2340
+ ad=0 pd=0 as=0 ps=0 
M2639 diff_87360_101640# diff_86760_94560# GND GND efet w=720 l=2040
+ ad=0 pd=0 as=0 ps=0 
M2640 diff_90000_47280# diff_92160_93720# diff_90000_47280# GND efet w=6180 l=4140
+ ad=0 pd=0 as=0 ps=0 
M2641 diff_94440_111840# GND diff_94440_111840# GND efet w=300 l=3840
+ ad=0 pd=0 as=0 ps=0 
M2642 GND diff_111720_106680# diff_110280_107400# GND efet w=1080 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2643 diff_97440_92520# GND GND GND efet w=480 l=6000
+ ad=0 pd=0 as=0 ps=0 
M2644 diff_94440_117120# GND GND GND efet w=720 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2645 GND diff_70080_105840# diff_118080_91560# GND efet w=1200 l=960
+ ad=0 pd=0 as=1.6056e+07 ps=52800 
M2646 diff_118080_91560# diff_117480_108840# GND GND efet w=1320 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2647 GND GND diff_126240_106680# GND efet w=960 l=960
+ ad=0 pd=0 as=1.08e+06 ps=6480 
M2648 GND GND diff_131760_114840# GND efet w=540 l=1140
+ ad=0 pd=0 as=1.0944e+06 ps=5520 
M2649 diff_90000_47280# diff_92160_93720# GND GND efet w=900 l=2460
+ ad=0 pd=0 as=0 ps=0 
M2650 GND GND diff_110280_107400# GND efet w=720 l=5400
+ ad=0 pd=0 as=0 ps=0 
M2651 diff_111720_106680# GND GND GND efet w=480 l=5040
+ ad=0 pd=0 as=0 ps=0 
M2652 GND GND diff_117480_108840# GND efet w=660 l=7020
+ ad=0 pd=0 as=0 ps=0 
M2653 diff_118080_91560# GND GND GND efet w=600 l=5400
+ ad=0 pd=0 as=0 ps=0 
M2654 diff_128040_60120# diff_126240_106680# GND GND efet w=1140 l=960
+ ad=1.476e+07 pd=61920 as=0 ps=0 
M2655 GND GND diff_128040_60120# GND efet w=1080 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2656 GND GND GND GND efet w=540 l=5280
+ ad=0 pd=0 as=0 ps=0 
M2657 diff_126240_106680# GND diff_126240_106680# GND efet w=300 l=7260
+ ad=0 pd=0 as=0 ps=0 
M2658 GND GND diff_99120_25800# GND efet w=1620 l=1140
+ ad=0 pd=0 as=1.43136e+07 ps=57600 
M2659 diff_104880_119520# GND GND GND efet w=1080 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2660 diff_99120_118920# GND GND GND efet w=1020 l=1380
+ ad=0 pd=0 as=0 ps=0 
M2661 GND GND GND GND efet w=1800 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2662 diff_99120_118920# GND diff_99120_118920# GND efet w=240 l=5280
+ ad=0 pd=0 as=0 ps=0 
M2663 GND GND GND GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M2664 diff_104880_119520# GND GND GND efet w=1080 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2665 GND GND diff_98880_123960# GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M2666 GND GND diff_104880_119520# GND efet w=1140 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2667 GND GND diff_99120_118920# GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M2668 GND GND GND GND efet w=1440 l=1440
+ ad=0 pd=0 as=0 ps=0 
M2669 diff_172560_117720# GND diff_172560_117720# GND efet w=480 l=3720
+ ad=3.9744e+06 pd=14160 as=0 ps=0 
M2670 GND diff_183360_117720# GND GND efet w=2700 l=2100
+ ad=0 pd=0 as=0 ps=0 
M2671 diff_172560_117720# GND GND GND efet w=2100 l=1380
+ ad=0 pd=0 as=0 ps=0 
M2672 GND GND diff_177960_117720# GND efet w=660 l=3180
+ ad=0 pd=0 as=3.816e+06 ps=13440 
M2673 GND diff_165480_110160# GND GND efet w=4860 l=1500
+ ad=0 pd=0 as=0 ps=0 
M2674 GND GND diff_134400_26040# GND efet w=4500 l=1020
+ ad=0 pd=0 as=1.8576e+07 ps=68160 
M2675 diff_134400_26040# diff_219720_138000# diff_134400_26040# GND efet w=5400 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2676 diff_219720_138000# GND GND GND efet w=720 l=1320
+ ad=374400 pd=2880 as=0 ps=0 
M2677 GND GND diff_213360_134760# GND efet w=1080 l=2760
+ ad=0 pd=0 as=1.008e+07 ps=24240 
M2678 GND diff_165480_110160# diff_66000_145440# GND efet w=5400 l=1080
+ ad=0 pd=0 as=1.96704e+07 ps=53520 
M2679 GND diff_188760_119280# diff_89400_129240# GND efet w=3120 l=1200
+ ad=0 pd=0 as=1.71936e+07 ps=54000 
M2680 diff_66000_145440# diff_187800_118320# GND GND efet w=5820 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2681 diff_134400_26040# diff_219720_138000# GND GND efet w=1080 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2682 diff_213360_134760# diff_134400_26040# GND GND efet w=2280 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2683 diff_213360_134760# GND GND GND efet w=4020 l=1500
+ ad=0 pd=0 as=0 ps=0 
M2684 GND diff_187800_118320# diff_89400_129240# GND efet w=4380 l=2100
+ ad=0 pd=0 as=0 ps=0 
M2685 diff_66000_145440# diff_188760_119280# GND GND efet w=2400 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2686 GND GND diff_183360_117720# GND efet w=600 l=3360
+ ad=0 pd=0 as=4.2624e+06 ps=15840 
M2687 diff_177960_117720# GND GND GND efet w=1800 l=1620
+ ad=0 pd=0 as=0 ps=0 
M2688 GND diff_174480_111480# GND GND efet w=4680 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2689 GND diff_179880_112560# GND GND efet w=4620 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2690 GND GND diff_165480_110160# GND efet w=1260 l=1020
+ ad=0 pd=0 as=1.08864e+07 ps=38400 
M2691 diff_183360_117720# GND GND GND efet w=1740 l=1680
+ ad=0 pd=0 as=0 ps=0 
M2692 GND GND diff_188760_119280# GND efet w=780 l=2940
+ ad=0 pd=0 as=3.2832e+06 ps=12240 
M2693 diff_188760_119280# diff_187800_118320# GND GND efet w=2880 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2694 GND diff_185280_114120# GND GND efet w=4740 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2695 GND diff_192360_116040# diff_187800_118320# GND efet w=5340 l=1020
+ ad=0 pd=0 as=3.2832e+06 ps=18960 
M2696 GND GND GND GND efet w=720 l=960
+ ad=0 pd=0 as=0 ps=0 
M2697 diff_218280_127680# GND GND GND efet w=720 l=1440
+ ad=374400 pd=3600 as=0 ps=0 
M2698 GND diff_218280_127680# GND GND efet w=5700 l=600
+ ad=0 pd=0 as=0 ps=0 
M2699 GND diff_218280_127680# GND GND efet w=840 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2700 GND GND GND GND efet w=840 l=960
+ ad=0 pd=0 as=0 ps=0 
M2701 GND GND GND GND efet w=4080 l=3300
+ ad=0 pd=0 as=0 ps=0 
M2702 GND GND GND GND efet w=3480 l=1920
+ ad=0 pd=0 as=0 ps=0 
M2703 GND GND GND GND efet w=20760 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2704 GND GND GND GND efet w=18840 l=960
+ ad=0 pd=0 as=0 ps=0 
M2705 GND GND GND GND efet w=6000 l=3120
+ ad=0 pd=0 as=0 ps=0 
M2706 GND GND GND GND efet w=4800 l=1860
+ ad=0 pd=0 as=0 ps=0 
M2707 GND diff_188880_226560# diff_192360_116040# GND efet w=840 l=1080
+ ad=0 pd=0 as=446400 ps=3360 
M2708 GND GND GND GND efet w=3900 l=1380
+ ad=0 pd=0 as=0 ps=0 
M2709 GND GND GND GND efet w=1620 l=3480
+ ad=0 pd=0 as=0 ps=0 
M2710 diff_165480_110160# GND GND GND efet w=900 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2711 diff_98880_123960# GND diff_98880_123960# GND efet w=300 l=6180
+ ad=0 pd=0 as=0 ps=0 
M2712 GND GND GND GND efet w=960 l=2520
+ ad=0 pd=0 as=0 ps=0 
M2713 GND GND GND GND efet w=1020 l=4080
+ ad=0 pd=0 as=0 ps=0 
M2714 diff_187800_118320# GND GND GND efet w=780 l=4260
+ ad=0 pd=0 as=0 ps=0 
M2715 GND diff_188880_226560# diff_185280_114120# GND efet w=900 l=1140
+ ad=0 pd=0 as=374400 ps=3360 
M2716 GND GND GND GND efet w=101580 l=2100
+ ad=0 pd=0 as=0 ps=0 
M2717 GND diff_165480_110160# diff_165480_110160# GND efet w=3240 l=1560
+ ad=0 pd=0 as=0 ps=0 
M2718 GND GND diff_165480_110160# GND efet w=600 l=5760
+ ad=0 pd=0 as=0 ps=0 
M2719 diff_165480_110160# GND GND GND efet w=3060 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2720 GND diff_188880_226560# diff_179880_112560# GND efet w=900 l=1140
+ ad=0 pd=0 as=388800 ps=3360 
M2721 GND GND GND GND efet w=54420 l=900
+ ad=0 pd=0 as=0 ps=0 
M2722 diff_165480_110160# diff_173520_107280# diff_165480_110160# GND efet w=3120 l=3960
+ ad=0 pd=0 as=0 ps=0 
M2723 GND diff_188880_226560# diff_174480_111480# GND efet w=840 l=960
+ ad=0 pd=0 as=475200 ps=3360 
M2724 GND diff_173520_107280# diff_165480_110160# GND efet w=720 l=1680
+ ad=0 pd=0 as=0 ps=0 
M2725 GND GND GND GND efet w=3840 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2726 GND GND GND GND efet w=3300 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2727 GND GND diff_173520_107280# GND efet w=600 l=960
+ ad=0 pd=0 as=360000 ps=2400 
M2728 GND GND GND GND efet w=660 l=3000
+ ad=0 pd=0 as=0 ps=0 
M2729 GND GND GND GND efet w=960 l=1740
+ ad=0 pd=0 as=0 ps=0 
M2730 GND GND GND GND efet w=4440 l=840
+ ad=0 pd=0 as=0 ps=0 
M2731 GND GND diff_174240_97200# GND efet w=960 l=3120
+ ad=0 pd=0 as=4.7808e+06 ps=13680 
M2732 GND diff_108000_115920# diff_165720_88920# GND efet w=960 l=1020
+ ad=0 pd=0 as=2.5056e+06 ps=7200 
M2733 diff_182640_101160# GND GND GND efet w=600 l=1680
+ ad=1.02816e+07 pd=36480 as=0 ps=0 
M2734 GND diff_178920_94920# diff_193560_103560# GND efet w=4740 l=1260
+ ad=0 pd=0 as=2.4336e+06 ps=9840 
M2735 GND diff_178920_94920# diff_182640_101160# GND efet w=3540 l=900
+ ad=0 pd=0 as=0 ps=0 
M2736 GND GND diff_165720_88920# GND efet w=1080 l=7200
+ ad=0 pd=0 as=0 ps=0 
M2737 diff_165720_88920# GND GND GND efet w=1020 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2738 GND GND diff_133440_86160# GND efet w=1200 l=960
+ ad=0 pd=0 as=7.8192e+06 ps=27840 
M2739 GND diff_99120_118920# diff_131760_92520# GND efet w=960 l=900
+ ad=0 pd=0 as=6.7824e+06 ps=33120 
M2740 GND GND diff_171960_95040# GND efet w=720 l=2820
+ ad=0 pd=0 as=2.4912e+06 ps=7920 
M2741 GND GND diff_182640_101160# GND efet w=1740 l=1560
+ ad=0 pd=0 as=0 ps=0 
M2742 diff_55200_81120# diff_118080_91560# diff_118080_91560# GND efet w=840 l=1320
+ ad=4.70736e+07 pd=154560 as=0 ps=0 
M2743 diff_86760_94560# GND GND GND efet w=480 l=960
+ ad=403200 pd=2640 as=0 ps=0 
M2744 diff_92160_93720# GND diff_92160_93720# GND efet w=240 l=1560
+ ad=403200 pd=2640 as=0 ps=0 
M2745 diff_106320_90480# GND diff_102480_94560# GND efet w=1320 l=840
+ ad=1.07568e+07 pd=38640 as=2.52e+06 ps=8880 
M2746 diff_102480_94560# GND GND GND efet w=780 l=1440
+ ad=0 pd=0 as=0 ps=0 
M2747 diff_133440_86160# diff_142920_94680# diff_133440_86160# GND efet w=4980 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2748 diff_106320_90480# GND diff_104520_92040# GND efet w=660 l=1020
+ ad=0 pd=0 as=2.0376e+07 ps=66240 
M2749 diff_132720_93000# diff_131760_92520# diff_104520_92040# GND efet w=1200 l=960
+ ad=4.8816e+06 pd=18720 as=0 ps=0 
M2750 diff_104520_92040# GND GND GND efet w=840 l=2880
+ ad=0 pd=0 as=0 ps=0 
M2751 diff_104520_92040# GND GND GND efet w=3120 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2752 diff_118080_91560# diff_110280_107400# diff_106320_90480# GND efet w=1200 l=960
+ ad=0 pd=0 as=0 ps=0 
M2753 GND diff_97440_92520# diff_55200_81120# GND efet w=4740 l=840
+ ad=0 pd=0 as=0 ps=0 
M2754 GND GND diff_133440_86160# GND efet w=1140 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2755 diff_131760_92520# diff_147840_90120# diff_131760_92520# GND efet w=6600 l=1680
+ ad=0 pd=0 as=0 ps=0 
M2756 diff_119880_90240# diff_118920_89640# diff_106320_90480# GND efet w=840 l=1080
+ ad=1.01952e+07 pd=26400 as=0 ps=0 
M2757 GND diff_106320_90480# GND GND efet w=4920 l=960
+ ad=0 pd=0 as=0 ps=0 
M2758 GND GND GND GND efet w=840 l=2760
+ ad=0 pd=0 as=0 ps=0 
M2759 diff_90240_74760# diff_118080_91560# diff_106320_90480# GND efet w=600 l=960
+ ad=6.22656e+07 pd=174240 as=0 ps=0 
M2760 diff_133440_86160# diff_142920_94680# GND GND efet w=540 l=4020
+ ad=0 pd=0 as=0 ps=0 
M2761 GND GND diff_131760_92520# GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M2762 GND diff_104880_119520# diff_131640_42480# GND efet w=1200 l=960
+ ad=0 pd=0 as=9.9936e+06 ps=42240 
M2763 GND GND diff_131640_42480# GND efet w=1260 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2764 GND GND diff_118920_89640# GND efet w=1140 l=900
+ ad=0 pd=0 as=3.672e+06 ps=9120 
M2765 diff_98880_123960# diff_98880_123960# GND GND efet w=960 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2766 diff_174240_97200# GND GND GND efet w=1860 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2767 GND GND diff_193560_103560# GND efet w=3600 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2768 GND diff_174240_97200# diff_171960_95040# GND efet w=2400 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2769 GND diff_176280_101040# diff_174240_97200# GND efet w=2040 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2770 diff_182640_101160# diff_134400_26040# diff_176280_101040# GND efet w=840 l=960
+ ad=0 pd=0 as=1.4112e+06 ps=7680 
M2771 diff_111960_24480# diff_171960_95040# GND GND efet w=3420 l=1200
+ ad=3.22704e+07 pd=78960 as=0 ps=0 
M2772 diff_174240_97200# GND GND GND efet w=1920 l=960
+ ad=0 pd=0 as=0 ps=0 
M2773 GND diff_174240_97200# diff_111960_24480# GND efet w=3780 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2774 GND diff_159360_93840# diff_118920_89640# GND efet w=1080 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2775 GND diff_159360_93840# diff_98880_123960# GND efet w=1200 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2776 GND GND diff_98880_123960# GND efet w=480 l=5760
+ ad=0 pd=0 as=0 ps=0 
M2777 GND diff_147840_90120# diff_131760_92520# GND efet w=480 l=4800
+ ad=0 pd=0 as=0 ps=0 
M2778 diff_118920_89640# GND GND GND efet w=720 l=6600
+ ad=0 pd=0 as=0 ps=0 
M2779 diff_147840_90120# GND GND GND efet w=600 l=960
+ ad=878400 pd=5280 as=0 ps=0 
M2780 diff_142920_94680# GND GND GND efet w=660 l=840
+ ad=417600 pd=3120 as=0 ps=0 
M2781 diff_178920_94920# GND diff_185640_97320# GND efet w=900 l=1080
+ ad=0 pd=0 as=576000 ps=3360 
M2782 GND GND diff_194040_99480# GND efet w=3720 l=1320
+ ad=0 pd=0 as=2.952e+06 ps=10800 
M2783 diff_194040_99480# GND GND GND efet w=4080 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2784 GND diff_185640_97320# GND GND efet w=4920 l=780
+ ad=0 pd=0 as=0 ps=0 
M2785 GND diff_178920_94920# diff_178200_92400# GND efet w=10440 l=1080
+ ad=0 pd=0 as=6.5952e+06 ps=22560 
M2786 GND GND GND GND efet w=4620 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2787 diff_178200_92400# diff_134400_26040# GND GND efet w=7980 l=900
+ ad=0 pd=0 as=0 ps=0 
M2788 GND GND GND GND efet w=1260 l=2280
+ ad=0 pd=0 as=0 ps=0 
M2789 GND GND diff_188040_90240# GND efet w=3120 l=1320
+ ad=0 pd=0 as=2.808e+06 ps=12480 
M2790 GND GND diff_132720_93000# GND efet w=840 l=840
+ ad=0 pd=0 as=0 ps=0 
M2791 diff_132720_93000# diff_165720_88920# GND GND efet w=780 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2792 GND diff_96720_85440# diff_55200_81120# GND efet w=4440 l=840
+ ad=0 pd=0 as=0 ps=0 
M2793 diff_55200_81120# GND GND GND efet w=540 l=2400
+ ad=0 pd=0 as=0 ps=0 
M2794 GND diff_99120_25800# diff_96720_85440# GND efet w=720 l=840
+ ad=0 pd=0 as=3.2112e+06 ps=12960 
M2795 diff_132720_93000# diff_133440_86160# GND GND efet w=1320 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2796 GND GND diff_175680_35880# GND efet w=1080 l=960
+ ad=0 pd=0 as=1.02096e+07 ps=37440 
M2797 diff_175680_35880# GND GND GND efet w=1500 l=780
+ ad=0 pd=0 as=0 ps=0 
M2798 diff_188040_90240# GND GND GND efet w=780 l=3180
+ ad=0 pd=0 as=0 ps=0 
M2799 GND diff_188040_90240# GND GND efet w=5460 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2800 GND GND GND GND efet w=1140 l=960
+ ad=0 pd=0 as=0 ps=0 
M2801 diff_152520_82440# diff_132720_93000# diff_150960_82320# GND efet w=4920 l=960
+ ad=3.7296e+06 pd=14880 as=2.4768e+06 ps=10320 
M2802 GND diff_132720_93000# diff_153120_82680# GND efet w=5100 l=900
+ ad=0 pd=0 as=1.86192e+07 ps=57360 
M2803 GND diff_144480_78240# diff_90240_74760# GND efet w=5040 l=960
+ ad=0 pd=0 as=0 ps=0 
M2804 GND GND GND GND efet w=600 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2805 GND diff_96000_83640# GND GND efet w=4860 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2806 diff_106800_81960# diff_99120_25800# diff_96000_83640# GND efet w=660 l=1020
+ ad=2.2104e+07 pd=60720 as=2.7072e+06 ps=10560 
M2807 GND GND GND GND efet w=540 l=2700
+ ad=0 pd=0 as=0 ps=0 
M2808 GND diff_128040_60120# diff_106800_81960# GND efet w=1200 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2809 diff_90240_74760# diff_143280_82080# GND GND efet w=1080 l=840
+ ad=0 pd=0 as=0 ps=0 
M2810 diff_150960_82320# GND GND GND efet w=3660 l=900
+ ad=0 pd=0 as=0 ps=0 
M2811 GND diff_55200_81120# diff_56400_79440# GND efet w=1200 l=1440
+ ad=0 pd=0 as=3.8448e+06 ps=15600 
M2812 GND diff_24120_80040# GND GND efet w=2400 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2813 GND GND diff_28560_76560# GND efet w=540 l=960
+ ad=0 pd=0 as=460800 ps=2880 
M2814 diff_41040_77520# GND GND GND efet w=720 l=1080
+ ad=446400 pd=2880 as=0 ps=0 
M2815 GND GND GND GND efet w=6420 l=900
+ ad=0 pd=0 as=0 ps=0 
M2816 GND diff_28560_76560# GND GND efet w=480 l=2280
+ ad=0 pd=0 as=0 ps=0 
M2817 diff_24120_80040# GND diff_30240_71280# GND efet w=1320 l=840
+ ad=1.0368e+06 pd=5280 as=4.9392e+06 ps=17760 
M2818 diff_30240_71280# diff_28080_71160# GND GND efet w=2280 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2819 diff_28080_71160# GND diff_11280_215400# GND efet w=1200 l=960
+ ad=1.08e+06 pd=4800 as=1.05523e+08 ps=304560 
M2820 GND GND diff_30240_71280# GND efet w=720 l=3360
+ ad=0 pd=0 as=0 ps=0 
M2821 diff_20640_113640# diff_11280_215400# GND GND efet w=1920 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2822 GND GND diff_62400_80640# GND efet w=1080 l=960
+ ad=0 pd=0 as=1.7856e+06 ps=6240 
M2823 diff_70320_79920# diff_56400_79440# GND GND efet w=2340 l=960
+ ad=1.44e+06 pd=6000 as=0 ps=0 
M2824 GND GND diff_70320_79920# GND efet w=2400 l=960
+ ad=0 pd=0 as=0 ps=0 
M2825 GND GND GND GND efet w=900 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2826 GND GND GND GND efet w=1440 l=960
+ ad=0 pd=0 as=0 ps=0 
M2827 diff_106800_81960# GND GND GND efet w=840 l=3120
+ ad=0 pd=0 as=0 ps=0 
M2828 diff_56400_79440# GND diff_56400_73800# GND efet w=2340 l=840
+ ad=0 pd=0 as=8.5536e+06 ps=30240 
M2829 GND diff_27960_63360# diff_11280_215400# GND efet w=3180 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2830 diff_11280_215400# diff_24120_68040# GND GND efet w=3240 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2831 diff_27960_63360# diff_28680_63960# diff_27960_63360# GND efet w=5640 l=540
+ ad=8.0496e+06 pd=28800 as=0 ps=0 
M2832 diff_27960_63360# diff_24120_68040# GND GND efet w=2880 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2833 GND GND diff_28680_63960# GND efet w=480 l=1080
+ ad=0 pd=0 as=489600 ps=3120 
M2834 GND diff_28680_63960# diff_27960_63360# GND efet w=600 l=2160
+ ad=0 pd=0 as=0 ps=0 
M2835 GND GND diff_44280_73320# GND efet w=720 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2836 GND GND GND GND efet w=660 l=3780
+ ad=0 pd=0 as=0 ps=0 
M2837 GND GND GND GND efet w=600 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2838 GND GND diff_56400_73800# GND efet w=2760 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2839 diff_56400_73800# GND GND GND efet w=3120 l=960
+ ad=0 pd=0 as=0 ps=0 
M2840 diff_56400_79440# GND GND GND efet w=300 l=4380
+ ad=0 pd=0 as=0 ps=0 
M2841 GND GND GND GND efet w=480 l=2820
+ ad=0 pd=0 as=0 ps=0 
M2842 diff_62400_80640# GND GND GND efet w=480 l=5880
+ ad=0 pd=0 as=0 ps=0 
M2843 GND GND GND GND efet w=540 l=3900
+ ad=0 pd=0 as=0 ps=0 
M2844 GND GND GND GND efet w=720 l=4200
+ ad=0 pd=0 as=0 ps=0 
M2845 GND GND GND GND efet w=420 l=3780
+ ad=0 pd=0 as=0 ps=0 
M2846 GND GND diff_59400_45960# GND efet w=660 l=4260
+ ad=0 pd=0 as=1.49328e+07 ps=42960 
M2847 GND GND GND GND efet w=300 l=4260
+ ad=0 pd=0 as=0 ps=0 
M2848 GND GND GND GND efet w=2220 l=1620
+ ad=0 pd=0 as=0 ps=0 
M2849 GND GND diff_76560_120480# GND efet w=1800 l=960
+ ad=0 pd=0 as=1.38096e+07 ps=37920 
M2850 diff_55200_81120# diff_110280_107400# GND GND efet w=600 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2851 GND GND diff_106800_81960# GND efet w=4200 l=1860
+ ad=0 pd=0 as=0 ps=0 
M2852 GND GND GND GND efet w=1080 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2853 diff_104520_77760# GND GND GND efet w=780 l=3060
+ ad=1.99728e+07 pd=60480 as=0 ps=0 
M2854 GND diff_90000_47280# GND GND efet w=3600 l=900
+ ad=0 pd=0 as=0 ps=0 
M2855 diff_76560_120480# GND GND GND efet w=720 l=3720
+ ad=0 pd=0 as=0 ps=0 
M2856 GND diff_90240_74760# diff_72120_132600# GND efet w=3540 l=900
+ ad=0 pd=0 as=1.1448e+07 ps=37200 
M2857 GND GND diff_104520_77760# GND efet w=600 l=960
+ ad=0 pd=0 as=0 ps=0 
M2858 diff_90240_74760# diff_98880_123960# GND GND efet w=840 l=960
+ ad=0 pd=0 as=0 ps=0 
M2859 GND diff_144480_78240# diff_143280_82080# GND efet w=1020 l=1140
+ ad=0 pd=0 as=1.7856e+06 ps=6720 
M2860 diff_144480_78240# diff_153120_82680# diff_152520_82440# GND efet w=5040 l=1020
+ ad=6.336e+06 pd=23520 as=0 ps=0 
M2861 GND GND GND GND efet w=4980 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2862 diff_153120_82680# diff_153120_82680# GND GND efet w=3840 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2863 GND diff_106800_81960# diff_104520_77760# GND efet w=3000 l=960
+ ad=0 pd=0 as=0 ps=0 
M2864 diff_143280_82080# GND GND GND efet w=480 l=4920
+ ad=0 pd=0 as=0 ps=0 
M2865 diff_153120_82680# GND diff_159360_78360# GND efet w=5700 l=1440
+ ad=0 pd=0 as=4.8672e+06 ps=17040 
M2866 diff_159360_78360# diff_153120_82680# GND GND efet w=4620 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2867 diff_177840_83640# diff_182880_82560# GND GND efet w=1860 l=1020
+ ad=5.8608e+06 pd=18720 as=0 ps=0 
M2868 GND GND GND GND efet w=7740 l=900
+ ad=0 pd=0 as=0 ps=0 
M2869 diff_177840_83640# diff_175680_35880# diff_153120_82680# GND efet w=1140 l=900
+ ad=0 pd=0 as=0 ps=0 
M2870 GND diff_177480_79320# diff_177840_83640# GND efet w=1200 l=960
+ ad=0 pd=0 as=0 ps=0 
M2871 GND GND diff_159360_78360# GND efet w=480 l=5520
+ ad=0 pd=0 as=0 ps=0 
M2872 diff_90240_71400# diff_118080_91560# GND GND efet w=840 l=960
+ ad=5.66928e+07 pd=158160 as=0 ps=0 
M2873 diff_144480_78240# GND GND GND efet w=600 l=4440
+ ad=0 pd=0 as=0 ps=0 
M2874 diff_148800_77640# diff_147720_75720# diff_144480_78240# GND efet w=3000 l=1080
+ ad=5.8608e+06 pd=18960 as=0 ps=0 
M2875 GND GND diff_148800_77640# GND efet w=2940 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2876 diff_148800_77640# diff_132720_93000# GND GND efet w=3600 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2877 GND diff_153120_82680# diff_148800_77640# GND efet w=2940 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2878 diff_165240_79680# diff_159360_78360# GND GND efet w=960 l=960
+ ad=1.4256e+06 pd=7680 as=0 ps=0 
M2879 GND GND diff_165240_79680# GND efet w=600 l=5220
+ ad=0 pd=0 as=0 ps=0 
M2880 GND diff_87360_101640# diff_90240_74760# GND efet w=3360 l=960
+ ad=0 pd=0 as=0 ps=0 
M2881 GND diff_131640_42480# diff_104520_77760# GND efet w=1200 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2882 diff_182880_82560# GND GND GND efet w=360 l=3960
+ ad=1.4832e+06 pd=8640 as=0 ps=0 
M2883 GND diff_177480_79320# diff_182880_82560# GND efet w=1260 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2884 diff_177480_79320# GND diff_153120_82680# GND efet w=1260 l=1020
+ ad=1.37376e+07 pd=47520 as=0 ps=0 
M2885 diff_177480_79320# diff_182880_82560# GND GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M2886 GND diff_177480_79320# diff_177480_79320# GND efet w=1560 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2887 GND GND diff_188280_75600# GND efet w=600 l=960
+ ad=0 pd=0 as=2.52e+06 ps=9360 
M2888 diff_147720_75720# diff_165240_79680# GND GND efet w=1680 l=840
+ ad=9.5616e+06 pd=36000 as=0 ps=0 
M2889 GND diff_191520_73200# diff_188280_75600# GND efet w=1020 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2890 GND diff_188280_75600# diff_177480_79320# GND efet w=3480 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2891 diff_177480_79320# diff_179760_74400# diff_177480_79320# GND efet w=4260 l=1620
+ ad=0 pd=0 as=0 ps=0 
M2892 diff_177480_79320# diff_179760_74400# GND GND efet w=480 l=3960
+ ad=0 pd=0 as=0 ps=0 
M2893 GND diff_159360_78360# diff_147720_75720# GND efet w=1200 l=960
+ ad=0 pd=0 as=0 ps=0 
M2894 GND diff_144000_67920# diff_90240_71400# GND efet w=5220 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2895 GND diff_133080_73080# diff_128040_60120# GND efet w=480 l=3780
+ ad=0 pd=0 as=0 ps=0 
M2896 diff_128040_60120# diff_133080_73080# diff_128040_60120# GND efet w=6540 l=420
+ ad=0 pd=0 as=0 ps=0 
M2897 diff_72120_132600# GND GND GND efet w=720 l=3840
+ ad=0 pd=0 as=0 ps=0 
M2898 GND GND GND GND efet w=720 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2899 GND GND GND GND efet w=2940 l=840
+ ad=0 pd=0 as=0 ps=0 
M2900 diff_44280_73320# diff_44280_73320# GND GND efet w=1740 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2901 GND GND GND GND efet w=3420 l=1380
+ ad=0 pd=0 as=0 ps=0 
M2902 GND diff_44280_73320# diff_49440_63480# GND efet w=1020 l=1020
+ ad=0 pd=0 as=2.9952e+06 ps=12720 
M2903 GND GND GND GND efet w=1920 l=960
+ ad=0 pd=0 as=0 ps=0 
M2904 GND GND GND GND efet w=2940 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2905 GND diff_49440_63480# GND GND efet w=4200 l=840
+ ad=0 pd=0 as=0 ps=0 
M2906 diff_59400_45960# GND GND GND efet w=1200 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2907 GND GND GND GND efet w=1200 l=960
+ ad=0 pd=0 as=0 ps=0 
M2908 GND GND GND GND efet w=1320 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2909 GND GND GND GND efet w=1500 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2910 GND GND diff_59280_61920# GND efet w=480 l=4920
+ ad=0 pd=0 as=5.3136e+06 ps=20640 
M2911 GND diff_90240_71400# diff_72120_132600# GND efet w=3300 l=900
+ ad=0 pd=0 as=0 ps=0 
M2912 diff_90240_71400# diff_87360_101640# GND GND efet w=3300 l=960
+ ad=0 pd=0 as=0 ps=0 
M2913 GND GND diff_133080_73080# GND efet w=480 l=960
+ ad=0 pd=0 as=288000 ps=2160 
M2914 diff_90240_71400# diff_142320_69960# GND GND efet w=1320 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2915 GND GND diff_168720_72960# GND efet w=660 l=1020
+ ad=0 pd=0 as=633600 ps=4320 
M2916 GND diff_90000_47280# GND GND efet w=3300 l=960
+ ad=0 pd=0 as=0 ps=0 
M2917 diff_131160_70440# diff_128040_60120# diff_104520_69840# GND efet w=1200 l=1080
+ ad=1.35792e+07 pd=40560 as=1.77552e+07 ps=58800 
M2918 diff_152400_72000# diff_147720_75720# diff_149760_73320# GND efet w=4740 l=900
+ ad=4.0608e+06 pd=14400 as=3.2832e+06 ps=13200 
M2919 diff_149760_73320# diff_131160_70440# GND GND efet w=4800 l=960
+ ad=0 pd=0 as=0 ps=0 
M2920 diff_142320_69960# diff_153120_70680# diff_152400_72000# GND efet w=4980 l=960
+ ad=6.6528e+06 pd=21360 as=0 ps=0 
M2921 GND GND diff_76560_120480# GND efet w=1920 l=840
+ ad=0 pd=0 as=0 ps=0 
M2922 diff_104520_69840# GND GND GND efet w=900 l=2940
+ ad=0 pd=0 as=0 ps=0 
M2923 diff_104520_69840# GND diff_107760_66840# GND efet w=720 l=960
+ ad=0 pd=0 as=8.5248e+06 ps=33600 
M2924 diff_104520_69840# GND GND GND efet w=2700 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2925 diff_90240_74760# diff_110280_107400# diff_107760_66840# GND efet w=720 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2926 GND diff_142320_69960# diff_144000_67920# GND efet w=1020 l=900
+ ad=0 pd=0 as=2.0736e+06 ps=12000 
M2927 diff_147720_75720# diff_147720_75720# diff_160920_66360# GND efet w=4680 l=1200
+ ad=0 pd=0 as=9.864e+06 ps=30960 
M2928 diff_147720_75720# diff_131160_70440# GND GND efet w=5460 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2929 diff_160920_66360# diff_153120_70680# GND GND efet w=4020 l=900
+ ad=0 pd=0 as=0 ps=0 
M2930 GND diff_59280_61920# GND GND efet w=1440 l=960
+ ad=0 pd=0 as=0 ps=0 
M2931 diff_59280_61920# GND GND GND efet w=900 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2932 GND GND diff_57120_59640# GND efet w=540 l=5700
+ ad=0 pd=0 as=4.1472e+06 ps=18000 
M2933 diff_30240_59280# diff_28080_59280# GND GND efet w=2280 l=960
+ ad=4.7232e+06 pd=17280 as=0 ps=0 
M2934 diff_28080_59280# GND diff_21360_57480# GND efet w=1140 l=1020
+ ad=1.0224e+06 pd=4560 as=0 ps=0 
M2935 diff_24120_68040# GND diff_30240_59280# GND efet w=1200 l=960
+ ad=1.0368e+06 pd=5040 as=0 ps=0 
M2936 diff_30240_59280# GND diff_30240_59280# GND efet w=300 l=3480
+ ad=0 pd=0 as=0 ps=0 
M2937 GND diff_43680_56040# GND GND efet w=4080 l=960
+ ad=0 pd=0 as=0 ps=0 
M2938 diff_59280_61920# diff_44280_73320# diff_49440_63480# GND efet w=1020 l=840
+ ad=0 pd=0 as=0 ps=0 
M2939 diff_159360_66360# diff_153120_70680# diff_147720_75720# GND efet w=4740 l=1140
+ ad=1.04688e+07 pd=40560 as=0 ps=0 
M2940 diff_160920_66360# diff_131160_70440# diff_159360_66360# GND efet w=5580 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2941 diff_159360_66360# diff_168720_72960# diff_159360_66360# GND efet w=4140 l=1920
+ ad=0 pd=0 as=0 ps=0 
M2942 diff_179760_74400# GND GND GND efet w=720 l=960
+ ad=1.3104e+06 pd=5520 as=0 ps=0 
M2943 GND GND diff_191520_73200# GND efet w=1800 l=1320
+ ad=0 pd=0 as=3.9168e+06 ps=11040 
M2944 diff_191520_73200# GND GND GND efet w=900 l=2940
+ ad=0 pd=0 as=0 ps=0 
M2945 GND diff_131160_70440# diff_148680_65520# GND efet w=2880 l=1200
+ ad=0 pd=0 as=6.6096e+06 ps=19440 
M2946 GND diff_107760_66840# GND GND efet w=4920 l=960
+ ad=0 pd=0 as=0 ps=0 
M2947 diff_90240_71400# diff_98880_123960# diff_107760_66840# GND efet w=720 l=960
+ ad=0 pd=0 as=0 ps=0 
M2948 diff_144000_67920# GND GND GND efet w=600 l=4140
+ ad=0 pd=0 as=0 ps=0 
M2949 GND GND GND GND efet w=840 l=2760
+ ad=0 pd=0 as=0 ps=0 
M2950 diff_87000_54000# diff_118080_91560# diff_107760_66840# GND efet w=660 l=1140
+ ad=6.21792e+07 pd=171600 as=0 ps=0 
M2951 GND GND GND GND efet w=600 l=2760
+ ad=0 pd=0 as=0 ps=0 
M2952 GND GND GND GND efet w=4560 l=1200
+ ad=0 pd=0 as=0 ps=0 
M2953 GND diff_99120_25800# GND GND efet w=720 l=960
+ ad=0 pd=0 as=0 ps=0 
M2954 GND GND diff_131160_70440# GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M2955 diff_142320_69960# GND GND GND efet w=420 l=5700
+ ad=0 pd=0 as=0 ps=0 
M2956 diff_148680_65520# GND diff_142320_69960# GND efet w=2940 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2957 diff_148680_65520# diff_147720_75720# GND GND efet w=3600 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2958 GND diff_153120_70680# diff_148680_65520# GND efet w=3000 l=840
+ ad=0 pd=0 as=0 ps=0 
M2959 diff_131160_70440# diff_131640_42480# GND GND efet w=1320 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2960 diff_59400_45960# GND GND GND efet w=1500 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2961 GND GND GND GND efet w=960 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2962 GND GND GND GND efet w=1560 l=960
+ ad=0 pd=0 as=0 ps=0 
M2963 diff_20640_113640# diff_21360_57480# GND GND efet w=1920 l=1080
+ ad=0 pd=0 as=0 ps=0 
M2964 GND diff_49200_59400# diff_43680_56040# GND efet w=3240 l=960
+ ad=0 pd=0 as=7.2576e+06 ps=26160 
M2965 GND GND GND GND efet w=2640 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2966 GND diff_144360_54120# diff_87000_54000# GND efet w=5040 l=840
+ ad=0 pd=0 as=0 ps=0 
M2967 GND diff_168720_72960# diff_159360_66360# GND efet w=480 l=4260
+ ad=0 pd=0 as=0 ps=0 
M2968 diff_177360_65880# diff_175680_35880# diff_153120_70680# GND efet w=1200 l=960
+ ad=1.89792e+07 pd=63360 as=7.632e+06 ps=24480 
M2969 diff_177360_65880# diff_182160_70080# GND GND efet w=1680 l=960
+ ad=0 pd=0 as=0 ps=0 
M2970 diff_199440_72600# GND GND GND efet w=4740 l=1020
+ ad=7.7472e+06 pd=19680 as=0 ps=0 
M2971 GND GND GND GND efet w=2460 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2972 GND GND diff_199440_72600# GND efet w=900 l=3360
+ ad=0 pd=0 as=0 ps=0 
M2973 GND GND GND GND efet w=600 l=1320
+ ad=0 pd=0 as=0 ps=0 
M2974 GND GND GND GND efet w=600 l=1260
+ ad=0 pd=0 as=0 ps=0 
M2975 GND GND GND GND efet w=4500 l=2160
+ ad=0 pd=0 as=0 ps=0 
M2976 GND GND GND GND efet w=840 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2977 GND GND GND GND efet w=1020 l=1500
+ ad=0 pd=0 as=0 ps=0 
M2978 GND diff_177360_65880# diff_177360_65880# GND efet w=660 l=1500
+ ad=0 pd=0 as=0 ps=0 
M2979 GND diff_134400_26040# diff_199440_72600# GND efet w=2280 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2980 diff_182160_70080# GND GND GND efet w=420 l=4020
+ ad=1.7568e+06 pd=10080 as=0 ps=0 
M2981 diff_165120_67680# diff_159360_66360# GND GND efet w=1080 l=840
+ ad=1.4544e+06 pd=7920 as=0 ps=0 
M2982 GND GND diff_165120_67680# GND efet w=600 l=5220
+ ad=0 pd=0 as=0 ps=0 
M2983 GND diff_177360_65880# diff_182160_70080# GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M2984 GND GND GND GND efet w=1800 l=5580
+ ad=0 pd=0 as=0 ps=0 
M2985 GND GND diff_188160_64200# GND efet w=660 l=840
+ ad=0 pd=0 as=2.1888e+06 ps=7920 
M2986 diff_177360_65880# diff_182160_70080# GND GND efet w=1200 l=960
+ ad=0 pd=0 as=0 ps=0 
M2987 diff_177360_65880# GND diff_153120_70680# GND efet w=1500 l=1020
+ ad=0 pd=0 as=0 ps=0 
M2988 GND diff_177360_65880# diff_177360_65880# GND efet w=1200 l=1440
+ ad=0 pd=0 as=0 ps=0 
M2989 GND GND GND GND efet w=20820 l=1980
+ ad=0 pd=0 as=0 ps=0 
M2990 GND diff_191520_73200# diff_188160_64200# GND efet w=1020 l=1140
+ ad=0 pd=0 as=0 ps=0 
M2991 GND diff_165120_67680# GND GND efet w=1680 l=840
+ ad=0 pd=0 as=0 ps=0 
M2992 GND GND GND GND efet w=18780 l=960
+ ad=0 pd=0 as=0 ps=0 
M2993 GND diff_188160_64200# diff_177360_65880# GND efet w=3420 l=1500
+ ad=0 pd=0 as=0 ps=0 
M2994 GND diff_159360_66360# GND GND efet w=1200 l=840
+ ad=0 pd=0 as=0 ps=0 
M2995 diff_177360_65880# diff_179760_61200# diff_177360_65880# GND efet w=4140 l=1680
+ ad=0 pd=0 as=0 ps=0 
M2996 diff_177360_65880# diff_179760_61200# GND GND efet w=480 l=3600
+ ad=0 pd=0 as=0 ps=0 
M2997 GND diff_96120_61680# GND GND efet w=4680 l=960
+ ad=0 pd=0 as=0 ps=0 
M2998 diff_106800_59760# diff_99120_25800# diff_96120_61680# GND efet w=600 l=1080
+ ad=1.99728e+07 pd=55440 as=2.7504e+06 ps=10560 
M2999 GND GND GND GND efet w=720 l=2400
+ ad=0 pd=0 as=0 ps=0 
M3000 GND diff_27960_54240# diff_21360_57480# GND efet w=3420 l=900
+ ad=0 pd=0 as=0 ps=0 
M3001 diff_21360_57480# diff_24240_55920# GND GND efet w=3120 l=960
+ ad=0 pd=0 as=0 ps=0 
M3002 GND GND diff_43680_56040# GND efet w=1560 l=1320
+ ad=0 pd=0 as=0 ps=0 
M3003 diff_43680_56040# GND GND GND efet w=600 l=4080
+ ad=0 pd=0 as=0 ps=0 
M3004 diff_57120_59640# diff_44280_73320# diff_49200_59400# GND efet w=1020 l=1260
+ ad=0 pd=0 as=1.6848e+06 ps=10320 
M3005 GND diff_57120_59640# GND GND efet w=1440 l=840
+ ad=0 pd=0 as=0 ps=0 
M3006 GND GND diff_59400_45960# GND efet w=2040 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3007 GND GND GND GND efet w=900 l=1260
+ ad=0 pd=0 as=0 ps=0 
M3008 diff_57120_59640# GND GND GND efet w=1200 l=840
+ ad=0 pd=0 as=0 ps=0 
M3009 GND diff_128040_60120# diff_106800_59760# GND efet w=1260 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3010 diff_87000_54000# diff_143280_58080# GND GND efet w=1140 l=1260
+ ad=0 pd=0 as=0 ps=0 
M3011 diff_106800_59760# GND GND GND efet w=840 l=3420
+ ad=0 pd=0 as=0 ps=0 
M3012 GND GND GND GND efet w=1200 l=1200
+ ad=0 pd=0 as=0 ps=0 
M3013 GND GND GND GND efet w=2700 l=1140
+ ad=0 pd=0 as=0 ps=0 
M3014 GND diff_43680_56040# GND GND efet w=1920 l=960
+ ad=0 pd=0 as=0 ps=0 
M3015 GND GND GND GND efet w=600 l=4320
+ ad=0 pd=0 as=0 ps=0 
M3016 diff_27960_54240# diff_28680_52080# diff_27960_54240# GND efet w=5760 l=480
+ ad=7.128e+06 pd=28080 as=0 ps=0 
M3017 diff_27960_54240# diff_24240_55920# GND GND efet w=2700 l=1260
+ ad=0 pd=0 as=0 ps=0 
M3018 GND GND diff_28680_52080# GND efet w=540 l=1140
+ ad=0 pd=0 as=432000 ps=3360 
M3019 GND diff_28680_52080# diff_27960_54240# GND efet w=480 l=2040
+ ad=0 pd=0 as=0 ps=0 
M3020 GND diff_44280_73320# diff_49200_59400# GND efet w=840 l=960
+ ad=0 pd=0 as=0 ps=0 
M3021 GND GND diff_58920_54000# GND efet w=540 l=6060
+ ad=0 pd=0 as=2.7216e+06 ps=13680 
M3022 diff_58920_54000# diff_44280_73320# GND GND efet w=840 l=840
+ ad=0 pd=0 as=0 ps=0 
M3023 GND diff_58920_54000# GND GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M3024 diff_58920_54000# GND GND GND efet w=1260 l=900
+ ad=0 pd=0 as=0 ps=0 
M3025 GND GND diff_76560_120480# GND efet w=1920 l=960
+ ad=0 pd=0 as=0 ps=0 
M3026 diff_90240_71400# diff_110280_107400# GND GND efet w=600 l=1200
+ ad=0 pd=0 as=0 ps=0 
M3027 GND GND diff_106800_59760# GND efet w=4500 l=1800
+ ad=0 pd=0 as=0 ps=0 
M3028 diff_104520_55560# GND GND GND efet w=1020 l=3060
+ ad=2.00016e+07 pd=63600 as=0 ps=0 
M3029 GND diff_87000_54000# diff_72120_132600# GND efet w=3540 l=900
+ ad=0 pd=0 as=0 ps=0 
M3030 GND diff_90000_47280# GND GND efet w=3240 l=1140
+ ad=0 pd=0 as=0 ps=0 
M3031 diff_87000_54000# diff_98880_123960# GND GND efet w=660 l=960
+ ad=0 pd=0 as=0 ps=0 
M3032 GND GND diff_104520_55560# GND efet w=660 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3033 GND diff_106800_59760# diff_104520_55560# GND efet w=3000 l=960
+ ad=0 pd=0 as=0 ps=0 
M3034 diff_152400_58560# GND diff_149640_61440# GND efet w=4920 l=960
+ ad=4.4064e+06 pd=14880 as=3.528e+06 ps=13440 
M3035 diff_149640_61440# GND GND GND efet w=5040 l=840
+ ad=0 pd=0 as=0 ps=0 
M3036 diff_144360_54120# diff_148680_53520# diff_152400_58560# GND efet w=5400 l=900
+ ad=1.116e+07 pd=34800 as=0 ps=0 
M3037 GND GND GND GND efet w=5220 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3038 GND diff_144360_54120# diff_143280_58080# GND efet w=840 l=1020
+ ad=0 pd=0 as=1.5984e+06 ps=6480 
M3039 GND GND GND GND efet w=1260 l=900
+ ad=0 pd=0 as=0 ps=0 
M3040 diff_87000_49080# diff_118080_91560# GND GND efet w=780 l=1020
+ ad=5.14368e+07 pd=140640 as=0 ps=0 
M3041 diff_148680_53520# diff_148680_53520# GND GND efet w=4200 l=1080
+ ad=2.59776e+07 pd=81840 as=0 ps=0 
M3042 diff_148680_53520# GND diff_159360_54360# GND efet w=5640 l=1200
+ ad=0 pd=0 as=6.3936e+06 ps=20160 
M3043 diff_159360_54360# diff_148680_53520# GND GND efet w=4680 l=960
+ ad=0 pd=0 as=0 ps=0 
M3044 diff_143280_58080# GND GND GND efet w=480 l=5700
+ ad=0 pd=0 as=0 ps=0 
M3045 GND diff_87360_101640# diff_87000_54000# GND efet w=3540 l=960
+ ad=0 pd=0 as=0 ps=0 
M3046 GND diff_131640_42480# diff_104520_55560# GND efet w=1200 l=960
+ ad=0 pd=0 as=0 ps=0 
M3047 diff_144360_54120# GND GND GND efet w=600 l=4920
+ ad=0 pd=0 as=0 ps=0 
M3048 GND GND GND GND efet w=3360 l=1080
+ ad=0 pd=0 as=0 ps=0 
M3049 diff_30240_47160# diff_28080_47280# GND GND efet w=2280 l=960
+ ad=4.536e+06 pd=17280 as=0 ps=0 
M3050 diff_24240_55920# GND diff_30240_47160# GND efet w=1140 l=1020
+ ad=892800 pd=4800 as=0 ps=0 
M3051 diff_28080_47280# GND diff_21360_45480# GND efet w=1320 l=960
+ ad=892800 pd=4560 as=7.42752e+07 ps=188640 
M3052 GND GND GND GND efet w=3360 l=960
+ ad=0 pd=0 as=0 ps=0 
M3053 GND GND diff_59400_45960# GND efet w=1560 l=960
+ ad=0 pd=0 as=0 ps=0 
M3054 GND GND GND GND efet w=1620 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3055 GND GND GND GND efet w=1320 l=1200
+ ad=0 pd=0 as=0 ps=0 
M3056 GND GND GND GND efet w=2760 l=1080
+ ad=0 pd=0 as=0 ps=0 
M3057 diff_148680_53520# diff_144360_54120# diff_144360_54120# GND efet w=2460 l=1440
+ ad=0 pd=0 as=0 ps=0 
M3058 GND GND diff_148680_53520# GND efet w=3000 l=840
+ ad=0 pd=0 as=0 ps=0 
M3059 diff_148680_53520# GND GND GND efet w=3180 l=1380
+ ad=0 pd=0 as=0 ps=0 
M3060 GND diff_148680_53520# diff_148680_53520# GND efet w=3000 l=1440
+ ad=0 pd=0 as=0 ps=0 
M3061 diff_131640_42480# diff_133800_49440# diff_131640_42480# GND efet w=6720 l=360
+ ad=0 pd=0 as=0 ps=0 
M3062 GND GND diff_148680_53520# GND efet w=4680 l=1320
+ ad=0 pd=0 as=0 ps=0 
M3063 GND GND GND GND efet w=5700 l=3180
+ ad=0 pd=0 as=0 ps=0 
M3064 GND diff_191520_73200# GND GND efet w=1620 l=1440
+ ad=0 pd=0 as=0 ps=0 
M3065 GND GND GND GND efet w=4980 l=2100
+ ad=0 pd=0 as=0 ps=0 
M3066 diff_179760_61200# GND GND GND efet w=780 l=1020
+ ad=1.368e+06 pd=5280 as=0 ps=0 
M3067 GND GND diff_159360_54360# GND efet w=480 l=4800
+ ad=0 pd=0 as=0 ps=0 
M3068 diff_177480_52680# diff_182160_57120# GND GND efet w=1860 l=960
+ ad=1.73952e+07 pd=58560 as=0 ps=0 
M3069 diff_177480_52680# diff_175680_35880# diff_148680_53520# GND efet w=1320 l=900
+ ad=0 pd=0 as=0 ps=0 
M3070 GND diff_177480_52680# diff_177480_52680# GND efet w=720 l=1560
+ ad=0 pd=0 as=0 ps=0 
M3071 GND GND GND GND efet w=97500 l=2640
+ ad=0 pd=0 as=0 ps=0 
M3072 GND GND GND GND efet w=720 l=960
+ ad=0 pd=0 as=0 ps=0 
M3073 diff_197400_55440# diff_111960_24480# GND GND efet w=2160 l=1080
+ ad=5.7456e+06 pd=18240 as=0 ps=0 
M3074 diff_165120_55680# diff_159360_54360# GND GND efet w=1080 l=900
+ ad=1.3824e+06 pd=7680 as=0 ps=0 
M3075 GND GND diff_165120_55680# GND efet w=480 l=5280
+ ad=0 pd=0 as=0 ps=0 
M3076 diff_144360_54120# diff_165120_55680# GND GND efet w=1680 l=960
+ ad=0 pd=0 as=0 ps=0 
M3077 GND diff_159360_54360# diff_144360_54120# GND efet w=1260 l=900
+ ad=0 pd=0 as=0 ps=0 
M3078 GND GND diff_168960_46920# GND efet w=480 l=960
+ ad=0 pd=0 as=302400 ps=2400 
M3079 diff_182160_57120# GND GND GND efet w=420 l=3900
+ ad=1.584e+06 pd=9600 as=0 ps=0 
M3080 GND diff_177480_52680# diff_182160_57120# GND efet w=1140 l=1260
+ ad=0 pd=0 as=0 ps=0 
M3081 diff_177480_52680# diff_182160_57120# GND GND efet w=1320 l=1140
+ ad=0 pd=0 as=0 ps=0 
M3082 GND diff_177480_52680# diff_177480_52680# GND efet w=1140 l=1620
+ ad=0 pd=0 as=0 ps=0 
M3083 diff_177480_52680# GND diff_148680_53520# GND efet w=1260 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3084 GND GND GND GND efet w=49620 l=4500
+ ad=0 pd=0 as=0 ps=0 
M3085 GND GND diff_197400_55440# GND efet w=960 l=4320
+ ad=0 pd=0 as=0 ps=0 
M3086 diff_197400_55440# GND GND GND efet w=840 l=1440
+ ad=0 pd=0 as=0 ps=0 
M3087 diff_177480_52680# diff_180240_49440# GND GND efet w=720 l=4440
+ ad=0 pd=0 as=0 ps=0 
M3088 GND GND GND GND efet w=300 l=5340
+ ad=0 pd=0 as=0 ps=0 
M3089 GND diff_133800_49440# diff_131640_42480# GND efet w=540 l=3780
+ ad=0 pd=0 as=0 ps=0 
M3090 GND GND diff_30240_47160# GND efet w=600 l=3180
+ ad=0 pd=0 as=0 ps=0 
M3091 diff_20640_113640# diff_21360_45480# GND GND efet w=1860 l=960
+ ad=0 pd=0 as=0 ps=0 
M3092 GND GND GND GND efet w=720 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3093 GND GND GND GND efet w=600 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3094 GND diff_27960_42600# diff_21360_45480# GND efet w=3240 l=1080
+ ad=0 pd=0 as=0 ps=0 
M3095 GND GND GND GND efet w=1860 l=1200
+ ad=0 pd=0 as=0 ps=0 
M3096 GND GND GND GND efet w=1920 l=960
+ ad=0 pd=0 as=0 ps=0 
M3097 diff_21360_45480# diff_24240_43920# GND GND efet w=3180 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3098 diff_27960_42600# diff_28680_39960# diff_27960_42600# GND efet w=5640 l=480
+ ad=7.2576e+06 pd=28560 as=0 ps=0 
M3099 diff_27960_42600# diff_24240_43920# GND GND efet w=2280 l=960
+ ad=0 pd=0 as=0 ps=0 
M3100 GND GND diff_28680_39960# GND efet w=480 l=1020
+ ad=0 pd=0 as=504000 ps=3120 
M3101 GND diff_44280_73320# GND GND efet w=780 l=1140
+ ad=0 pd=0 as=0 ps=0 
M3102 GND GND diff_59400_45960# GND efet w=1140 l=1560
+ ad=0 pd=0 as=0 ps=0 
M3103 GND GND GND GND efet w=1260 l=900
+ ad=0 pd=0 as=0 ps=0 
M3104 GND GND GND GND efet w=960 l=840
+ ad=0 pd=0 as=0 ps=0 
M3105 GND diff_87000_49080# diff_72120_132600# GND efet w=3420 l=900
+ ad=0 pd=0 as=0 ps=0 
M3106 GND GND GND GND efet w=1440 l=840
+ ad=0 pd=0 as=0 ps=0 
M3107 GND GND GND GND efet w=1380 l=1500
+ ad=0 pd=0 as=0 ps=0 
M3108 GND GND GND GND efet w=2760 l=840
+ ad=0 pd=0 as=0 ps=0 
M3109 GND diff_28680_39960# diff_27960_42600# GND efet w=480 l=2160
+ ad=0 pd=0 as=0 ps=0 
M3110 diff_87000_49080# diff_87360_101640# GND GND efet w=3360 l=960
+ ad=0 pd=0 as=0 ps=0 
M3111 GND GND diff_133800_49440# GND efet w=480 l=840
+ ad=0 pd=0 as=230400 ps=1920 
M3112 diff_87000_49080# diff_142200_46080# GND GND efet w=1620 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3113 GND diff_90000_47280# GND GND efet w=3360 l=960
+ ad=0 pd=0 as=0 ps=0 
M3114 diff_131160_47160# diff_128040_60120# diff_104520_47640# GND efet w=1320 l=1140
+ ad=3.40848e+07 pd=131520 as=1.83024e+07 ps=60240 
M3115 GND GND GND GND efet w=5160 l=1320
+ ad=0 pd=0 as=0 ps=0 
M3116 GND diff_59400_45960# GND GND efet w=6000 l=960
+ ad=0 pd=0 as=0 ps=0 
M3117 GND GND GND GND efet w=5100 l=1380
+ ad=0 pd=0 as=0 ps=0 
M3118 GND GND GND GND efet w=6180 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3119 GND GND GND GND efet w=4500 l=1380
+ ad=0 pd=0 as=0 ps=0 
M3120 GND GND GND GND efet w=480 l=5520
+ ad=0 pd=0 as=0 ps=0 
M3121 GND diff_53880_36240# GND GND efet w=6360 l=600
+ ad=0 pd=0 as=0 ps=0 
M3122 GND GND GND GND efet w=2220 l=2580
+ ad=0 pd=0 as=0 ps=0 
M3123 diff_24240_43920# GND diff_30240_35160# GND efet w=1140 l=840
+ ad=950400 pd=5040 as=4.2624e+06 ps=17280 
M3124 diff_30240_35160# diff_28200_35160# GND GND efet w=2400 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3125 GND GND diff_30240_35160# GND efet w=420 l=3480
+ ad=0 pd=0 as=0 ps=0 
M3126 diff_28200_35160# GND diff_20640_113640# GND efet w=1080 l=960
+ ad=792000 pd=4080 as=0 ps=0 
M3127 GND GND GND GND efet w=3660 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3128 GND GND diff_53880_36240# GND efet w=360 l=1320
+ ad=0 pd=0 as=446400 ps=3360 
M3129 GND diff_53880_36240# GND GND efet w=840 l=2040
+ ad=0 pd=0 as=0 ps=0 
M3130 GND GND GND GND efet w=480 l=5520
+ ad=0 pd=0 as=0 ps=0 
M3131 GND GND diff_20640_113640# GND efet w=360 l=3240
+ ad=0 pd=0 as=0 ps=0 
M3132 GND diff_53880_29280# GND GND efet w=6360 l=840
+ ad=0 pd=0 as=0 ps=0 
M3133 GND GND GND GND efet w=2940 l=1740
+ ad=0 pd=0 as=0 ps=0 
M3134 GND GND GND GND efet w=9540 l=3180
+ ad=0 pd=0 as=0 ps=0 
M3135 GND GND GND GND efet w=3960 l=1560
+ ad=0 pd=0 as=0 ps=0 
M3136 GND GND GND GND efet w=3600 l=840
+ ad=0 pd=0 as=0 ps=0 
M3137 GND GND GND GND efet w=4560 l=1440
+ ad=0 pd=0 as=0 ps=0 
M3138 GND GND GND GND efet w=4920 l=960
+ ad=0 pd=0 as=0 ps=0 
M3139 GND GND GND GND efet w=4620 l=1320
+ ad=0 pd=0 as=0 ps=0 
M3140 GND GND GND GND efet w=4920 l=960
+ ad=0 pd=0 as=0 ps=0 
M3141 GND GND GND GND efet w=5040 l=840
+ ad=0 pd=0 as=0 ps=0 
M3142 GND GND diff_76560_120480# GND efet w=1920 l=960
+ ad=0 pd=0 as=0 ps=0 
M3143 diff_104520_47640# GND GND GND efet w=900 l=2940
+ ad=0 pd=0 as=0 ps=0 
M3144 GND diff_95880_45240# GND GND efet w=4440 l=1080
+ ad=0 pd=0 as=0 ps=0 
M3145 GND GND GND GND efet w=720 l=2880
+ ad=0 pd=0 as=0 ps=0 
M3146 GND GND GND GND efet w=4980 l=900
+ ad=0 pd=0 as=0 ps=0 
M3147 GND GND diff_53880_29280# GND efet w=660 l=1020
+ ad=0 pd=0 as=460800 ps=3360 
M3148 GND GND GND GND efet w=11580 l=1140
+ ad=0 pd=0 as=0 ps=0 
M3149 GND GND GND GND efet w=420 l=1980
+ ad=0 pd=0 as=0 ps=0 
M3150 GND GND GND GND efet w=540 l=1860
+ ad=0 pd=0 as=0 ps=0 
M3151 GND GND GND GND efet w=3360 l=1080
+ ad=0 pd=0 as=0 ps=0 
M3152 GND diff_53880_29280# GND GND efet w=840 l=2040
+ ad=0 pd=0 as=0 ps=0 
M3153 GND GND GND GND efet w=360 l=5280
+ ad=0 pd=0 as=0 ps=0 
M3154 GND diff_59400_45960# GND GND efet w=5100 l=900
+ ad=0 pd=0 as=0 ps=0 
M3155 diff_63960_26160# GND GND GND efet w=540 l=5640
+ ad=2.78496e+07 pd=79440 as=0 ps=0 
M3156 GND diff_56400_22080# GND GND efet w=6540 l=540
+ ad=0 pd=0 as=0 ps=0 
M3157 GND GND GND GND efet w=19080 l=3960
+ ad=0 pd=0 as=0 ps=0 
M3158 GND GND GND GND efet w=19020 l=3780
+ ad=0 pd=0 as=0 ps=0 
M3159 GND GND GND GND efet w=3120 l=1560
+ ad=0 pd=0 as=0 ps=0 
M3160 GND GND GND GND efet w=4920 l=960
+ ad=0 pd=0 as=0 ps=0 
M3161 GND GND GND GND efet w=6180 l=540
+ ad=0 pd=0 as=0 ps=0 
M3162 GND GND GND GND efet w=660 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3163 GND GND GND GND efet w=3540 l=1260
+ ad=0 pd=0 as=0 ps=0 
M3164 GND GND GND GND efet w=4980 l=1500
+ ad=0 pd=0 as=0 ps=0 
M3165 GND GND GND GND efet w=4980 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3166 GND GND GND GND efet w=4020 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3167 GND GND GND GND efet w=3720 l=1560
+ ad=0 pd=0 as=0 ps=0 
M3168 GND GND GND GND efet w=4440 l=1440
+ ad=0 pd=0 as=0 ps=0 
M3169 diff_56400_22080# GND diff_56400_22080# GND efet w=360 l=1320
+ ad=388800 pd=2640 as=0 ps=0 
M3170 GND diff_56400_22080# GND GND efet w=900 l=1980
+ ad=0 pd=0 as=0 ps=0 
M3171 GND GND GND GND efet w=780 l=1860
+ ad=0 pd=0 as=0 ps=0 
M3172 GND diff_59400_45960# diff_63960_26160# GND efet w=5160 l=1140
+ ad=0 pd=0 as=0 ps=0 
M3173 GND GND diff_63960_26160# GND efet w=5280 l=1320
+ ad=0 pd=0 as=0 ps=0 
M3174 GND GND diff_63960_26160# GND efet w=4980 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3175 GND GND GND GND efet w=3840 l=1320
+ ad=0 pd=0 as=0 ps=0 
M3176 GND GND diff_63960_26160# GND efet w=4260 l=1320
+ ad=0 pd=0 as=0 ps=0 
M3177 diff_104520_47640# GND diff_107760_44520# GND efet w=720 l=960
+ ad=0 pd=0 as=8.7264e+06 ps=32880 
M3178 diff_104520_47640# GND GND GND efet w=2820 l=1140
+ ad=0 pd=0 as=0 ps=0 
M3179 diff_87000_54000# diff_110280_107400# diff_107760_44520# GND efet w=720 l=960
+ ad=0 pd=0 as=0 ps=0 
M3180 GND diff_143880_43920# diff_87000_49080# GND efet w=5460 l=900
+ ad=0 pd=0 as=0 ps=0 
M3181 GND GND diff_177480_52680# GND efet w=3000 l=1560
+ ad=0 pd=0 as=0 ps=0 
M3182 diff_149640_49320# diff_131160_47160# GND GND efet w=4980 l=900
+ ad=3.5424e+06 pd=12960 as=0 ps=0 
M3183 GND diff_142200_46080# diff_143880_43920# GND efet w=1140 l=840
+ ad=0 pd=0 as=2.1744e+06 ps=10800 
M3184 diff_152400_46440# diff_144360_54120# diff_149640_49320# GND efet w=4680 l=960
+ ad=4.4784e+06 pd=15120 as=0 ps=0 
M3185 diff_142200_46080# diff_131160_47160# diff_152400_46440# GND efet w=5400 l=840
+ ad=6.912e+06 pd=23280 as=0 ps=0 
M3186 diff_131160_47160# diff_131160_47160# GND GND efet w=6120 l=1800
+ ad=0 pd=0 as=0 ps=0 
M3187 GND diff_131160_47160# diff_160800_42360# GND efet w=5100 l=2340
+ ad=0 pd=0 as=1.02384e+07 ps=30720 
M3188 GND diff_107760_44520# GND GND efet w=4860 l=1140
+ ad=0 pd=0 as=0 ps=0 
M3189 diff_87000_49080# diff_98880_123960# diff_107760_44520# GND efet w=780 l=900
+ ad=0 pd=0 as=0 ps=0 
M3190 GND GND GND GND efet w=780 l=2940
+ ad=0 pd=0 as=0 ps=0 
M3191 diff_87000_49080# diff_110280_107400# diff_118080_91560# GND efet w=1260 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3192 GND diff_99120_25800# diff_95880_45240# GND efet w=600 l=1080
+ ad=0 pd=0 as=2.6928e+06 ps=10560 
M3193 diff_118080_91560# diff_118080_91560# diff_107760_44520# GND efet w=1080 l=1140
+ ad=0 pd=0 as=0 ps=0 
M3194 diff_131160_47160# diff_131160_47160# diff_131160_47160# GND efet w=4620 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3195 GND diff_131160_47160# diff_131160_47160# GND efet w=2520 l=1440
+ ad=0 pd=0 as=0 ps=0 
M3196 diff_143880_43920# GND GND GND efet w=480 l=4800
+ ad=0 pd=0 as=0 ps=0 
M3197 GND GND diff_131160_47160# GND efet w=1140 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3198 diff_131160_47160# diff_119880_90240# diff_142200_46080# GND efet w=3120 l=840
+ ad=0 pd=0 as=0 ps=0 
M3199 diff_142200_46080# GND GND GND efet w=600 l=5400
+ ad=0 pd=0 as=0 ps=0 
M3200 diff_131160_47160# diff_131640_42480# GND GND efet w=1320 l=900
+ ad=0 pd=0 as=0 ps=0 
M3201 diff_160800_42360# diff_131160_47160# diff_131160_47160# GND efet w=5400 l=1440
+ ad=0 pd=0 as=0 ps=0 
M3202 diff_131160_47160# diff_144360_54120# GND GND efet w=3600 l=840
+ ad=0 pd=0 as=0 ps=0 
M3203 GND diff_131160_47160# diff_131160_47160# GND efet w=2940 l=1140
+ ad=0 pd=0 as=0 ps=0 
M3204 diff_131160_47160# diff_144360_54120# diff_160800_42360# GND efet w=4800 l=840
+ ad=0 pd=0 as=0 ps=0 
M3205 diff_177480_52680# diff_180240_49440# diff_177480_52680# GND efet w=3840 l=1740
+ ad=0 pd=0 as=0 ps=0 
M3206 diff_131160_47160# diff_168960_46920# diff_131160_47160# GND efet w=4740 l=2820
+ ad=0 pd=0 as=0 ps=0 
M3207 diff_180240_49440# GND GND GND efet w=1020 l=1080
+ ad=820800 pd=6000 as=0 ps=0 
M3208 GND GND GND GND efet w=3480 l=1740
+ ad=0 pd=0 as=0 ps=0 
M3209 GND diff_197400_55440# GND GND efet w=3300 l=1260
+ ad=0 pd=0 as=0 ps=0 
M3210 GND diff_168960_46920# diff_131160_47160# GND efet w=420 l=4320
+ ad=0 pd=0 as=0 ps=0 
M3211 GND GND GND GND efet w=840 l=3240
+ ad=0 pd=0 as=0 ps=0 
M3212 diff_177480_41640# diff_182040_45240# GND GND efet w=1740 l=1080
+ ad=1.91808e+07 pd=64080 as=0 ps=0 
M3213 GND GND GND GND efet w=5520 l=1380
+ ad=0 pd=0 as=0 ps=0 
M3214 diff_177480_41640# GND diff_131160_47160# GND efet w=1200 l=960
+ ad=0 pd=0 as=0 ps=0 
M3215 GND diff_111960_24480# GND GND efet w=3720 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3216 GND diff_177480_41640# diff_177480_41640# GND efet w=720 l=1440
+ ad=0 pd=0 as=0 ps=0 
M3217 diff_165360_43680# diff_131160_47160# GND GND efet w=1020 l=1020
+ ad=1.0656e+06 pd=6960 as=0 ps=0 
M3218 GND GND diff_165360_43680# GND efet w=480 l=5280
+ ad=0 pd=0 as=0 ps=0 
M3219 diff_119880_90240# diff_165360_43680# GND GND efet w=1560 l=960
+ ad=0 pd=0 as=0 ps=0 
M3220 diff_182040_45240# GND GND GND efet w=540 l=3780
+ ad=1.7568e+06 pd=9840 as=0 ps=0 
M3221 GND diff_177480_41640# diff_182040_45240# GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M3222 GND GND diff_190680_39840# GND efet w=780 l=720
+ ad=0 pd=0 as=2.1168e+06 ps=7680 
M3223 diff_177480_41640# diff_175680_35880# diff_131160_47160# GND efet w=1260 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3224 diff_177480_41640# diff_182040_45240# GND GND efet w=1140 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3225 GND diff_131160_47160# diff_119880_90240# GND efet w=1080 l=960
+ ad=0 pd=0 as=0 ps=0 
M3226 GND GND diff_182160_40080# GND efet w=540 l=780
+ ad=0 pd=0 as=288000 ps=2160 
M3227 GND diff_177480_41640# diff_177480_41640# GND efet w=1320 l=1320
+ ad=0 pd=0 as=0 ps=0 
M3228 GND diff_191520_73200# diff_190680_39840# GND efet w=1200 l=1200
+ ad=0 pd=0 as=0 ps=0 
M3229 diff_177480_41640# diff_182160_40080# diff_177480_41640# GND efet w=5640 l=480
+ ad=0 pd=0 as=0 ps=0 
M3230 GND diff_190680_39840# diff_177480_41640# GND efet w=3180 l=1140
+ ad=0 pd=0 as=0 ps=0 
M3231 GND GND GND GND efet w=9600 l=1080
+ ad=0 pd=0 as=0 ps=0 
M3232 diff_99120_25800# diff_99000_21120# diff_99120_25800# GND efet w=4740 l=1440
+ ad=0 pd=0 as=0 ps=0 
M3233 GND GND diff_63960_26160# GND efet w=4980 l=1140
+ ad=0 pd=0 as=0 ps=0 
M3234 GND GND diff_172440_35400# GND efet w=600 l=780
+ ad=0 pd=0 as=360000 ps=2880 
M3235 diff_177480_41640# diff_182160_40080# GND GND efet w=480 l=3360
+ ad=0 pd=0 as=0 ps=0 
M3236 diff_175680_35880# diff_172440_35400# diff_175680_35880# GND efet w=5520 l=480
+ ad=0 pd=0 as=0 ps=0 
M3237 diff_113400_27480# GND GND GND efet w=5940 l=1020
+ ad=1.20528e+07 pd=32640 as=0 ps=0 
M3238 GND diff_113400_27480# GND GND efet w=4080 l=960
+ ad=0 pd=0 as=0 ps=0 
M3239 GND diff_113400_27480# diff_117240_28320# GND efet w=1140 l=960
+ ad=0 pd=0 as=5.4432e+06 ps=18960 
M3240 GND GND GND GND efet w=9480 l=1200
+ ad=0 pd=0 as=0 ps=0 
M3241 diff_99120_25800# diff_99000_21120# GND GND efet w=600 l=4320
+ ad=0 pd=0 as=0 ps=0 
M3242 GND GND diff_99000_21120# GND efet w=720 l=1080
+ ad=0 pd=0 as=936000 ps=4560 
M3243 diff_113400_27480# diff_111960_24480# GND GND efet w=4260 l=1140
+ ad=0 pd=0 as=0 ps=0 
M3244 GND diff_111960_24480# diff_117240_28320# GND efet w=2100 l=960
+ ad=0 pd=0 as=0 ps=0 
M3245 GND diff_117240_28320# GND GND efet w=3180 l=1080
+ ad=0 pd=0 as=0 ps=0 
M3246 diff_113400_27480# GND GND GND efet w=840 l=3060
+ ad=0 pd=0 as=0 ps=0 
M3247 diff_117240_28320# GND GND GND efet w=480 l=4200
+ ad=0 pd=0 as=0 ps=0 
M3248 GND GND diff_135360_28440# GND efet w=4740 l=1020
+ ad=0 pd=0 as=5.9184e+06 ps=18000 
M3249 diff_135360_28440# GND GND GND efet w=1080 l=3240
+ ad=0 pd=0 as=0 ps=0 
M3250 diff_135360_28440# diff_134400_26040# diff_129000_14040# GND efet w=2280 l=960
+ ad=0 pd=0 as=2.232e+06 ps=7680 
M3251 GND diff_129000_14040# GND GND efet w=8220 l=900
+ ad=0 pd=0 as=0 ps=0 
M3252 GND GND GND GND efet w=53400 l=2640
+ ad=0 pd=0 as=0 ps=0 
M3253 GND GND GND GND efet w=4140 l=1620
+ ad=0 pd=0 as=0 ps=0 
M3254 GND GND GND GND efet w=10740 l=1980
+ ad=0 pd=0 as=0 ps=0 
M3255 GND GND GND GND efet w=10560 l=2160
+ ad=0 pd=0 as=0 ps=0 
M3256 GND GND GND GND efet w=600 l=1920
+ ad=0 pd=0 as=0 ps=0 
M3257 GND GND GND GND efet w=540 l=1980
+ ad=0 pd=0 as=0 ps=0 
M3258 GND GND GND GND efet w=3600 l=960
+ ad=0 pd=0 as=0 ps=0 
M3259 GND GND GND GND efet w=19080 l=3600
+ ad=0 pd=0 as=0 ps=0 
M3260 GND GND GND GND efet w=17940 l=4260
+ ad=0 pd=0 as=0 ps=0 
M3261 GND GND GND GND efet w=100200 l=1200
+ ad=0 pd=0 as=0 ps=0 
M3262 GND GND GND GND efet w=20520 l=960
+ ad=0 pd=0 as=0 ps=0 
M3263 GND GND GND GND efet w=780 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3264 GND GND GND GND efet w=900 l=1140
+ ad=0 pd=0 as=0 ps=0 
M3265 GND GND GND GND efet w=5400 l=1560
+ ad=0 pd=0 as=0 ps=0 
M3266 GND GND GND GND efet w=6780 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3267 GND GND GND GND efet w=18960 l=960
+ ad=0 pd=0 as=0 ps=0 
M3268 GND diff_136080_6840# GND GND efet w=840 l=960
+ ad=0 pd=0 as=0 ps=0 
M3269 GND diff_136080_6840# GND GND efet w=4800 l=2880
+ ad=0 pd=0 as=0 ps=0 
M3270 GND GND diff_136080_6840# GND efet w=840 l=1080
+ ad=0 pd=0 as=331200 ps=2880 
M3271 GND GND GND GND efet w=5520 l=1080
+ ad=0 pd=0 as=0 ps=0 
M3272 diff_175680_35880# diff_172440_35400# GND GND efet w=540 l=2760
+ ad=0 pd=0 as=0 ps=0 
M3273 GND GND GND GND efet w=8220 l=1260
+ ad=0 pd=0 as=0 ps=0 
M3274 GND GND GND GND efet w=3720 l=1320
+ ad=0 pd=0 as=0 ps=0 
M3275 diff_173520_28320# GND GND GND efet w=1380 l=900
+ ad=5.04e+06 pd=16080 as=0 ps=0 
M3276 GND diff_111960_24480# diff_173520_28320# GND efet w=2220 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3277 GND diff_111960_24480# GND GND efet w=3660 l=1140
+ ad=0 pd=0 as=0 ps=0 
M3278 GND GND diff_173520_28320# GND efet w=540 l=4620
+ ad=0 pd=0 as=0 ps=0 
M3279 GND diff_173520_28320# GND GND efet w=3240 l=960
+ ad=0 pd=0 as=0 ps=0 
M3280 GND GND GND GND efet w=540 l=3120
+ ad=0 pd=0 as=0 ps=0 
M3281 GND GND diff_191280_27720# GND efet w=4200 l=900
+ ad=0 pd=0 as=6.3792e+06 ps=18720 
M3282 diff_191280_27720# diff_134400_26040# GND GND efet w=2280 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3283 diff_191280_27720# GND GND GND efet w=900 l=3060
+ ad=0 pd=0 as=0 ps=0 
M3284 GND diff_111960_24480# GND GND efet w=4080 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3285 GND diff_202320_11520# GND GND efet w=3300 l=1020
+ ad=0 pd=0 as=0 ps=0 
M3286 GND GND GND GND efet w=2400 l=1200
+ ad=0 pd=0 as=0 ps=0 
M3287 GND GND GND GND efet w=54300 l=3060
+ ad=0 pd=0 as=0 ps=0 
M3288 GND GND GND GND efet w=2760 l=960
+ ad=0 pd=0 as=0 ps=0 
M3289 GND GND GND GND efet w=6120 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3290 GND GND GND GND efet w=20160 l=2760
+ ad=0 pd=0 as=0 ps=0 
M3291 GND GND GND GND efet w=600 l=960
+ ad=0 pd=0 as=0 ps=0 
M3292 GND GND GND GND efet w=780 l=1140
+ ad=0 pd=0 as=0 ps=0 
M3293 GND GND GND GND efet w=99600 l=1680
+ ad=0 pd=0 as=0 ps=0 
M3294 GND GND GND GND efet w=5040 l=1800
+ ad=0 pd=0 as=0 ps=0 
M3295 GND GND diff_202320_11520# GND efet w=780 l=4080
+ ad=0 pd=0 as=5.0976e+06 ps=18240 
M3296 GND GND diff_111960_24480# GND efet w=720 l=3000
+ ad=0 pd=0 as=0 ps=0 
M3297 GND diff_111960_24480# diff_111960_24480# GND efet w=4140 l=1740
+ ad=0 pd=0 as=0 ps=0 
M3298 GND GND GND GND efet w=6240 l=1080
+ ad=0 pd=0 as=0 ps=0 
M3299 GND GND GND GND efet w=18000 l=1920
+ ad=0 pd=0 as=0 ps=0 
M3300 GND GND GND GND efet w=840 l=1200
+ ad=0 pd=0 as=0 ps=0 
M3301 GND GND GND GND efet w=2940 l=4860
+ ad=0 pd=0 as=0 ps=0 
M3302 GND GND GND GND efet w=600 l=1140
+ ad=0 pd=0 as=0 ps=0 
M3303 GND diff_111960_24480# diff_202320_11520# GND efet w=1920 l=1320
+ ad=0 pd=0 as=0 ps=0 
M3304 diff_202320_11520# diff_111960_24480# GND GND efet w=1980 l=960
+ ad=0 pd=0 as=0 ps=0 
M3305 GND GND diff_111960_24480# GND efet w=7140 l=1260
+ ad=0 pd=0 as=0 ps=0 
M3306 GND GND GND GND efet w=9180 l=2220
+ ad=0 pd=0 as=0 ps=0 
M3307 GND GND GND GND efet w=2520 l=900
+ ad=0 pd=0 as=0 ps=0 
C0 metal_210600_287760# gnd! 23.1fF ;**FLOATING
C1 metal_209040_287400# gnd! 50.5fF ;**FLOATING
C2 metal_210000_293400# gnd! 19.9fF ;**FLOATING
C3 metal_207840_293640# gnd! 3.0fF ;**FLOATING
C4 metal_217320_295440# gnd! 5.2fF ;**FLOATING
C5 metal_221040_295200# gnd! 17.8fF ;**FLOATING
C6 metal_210000_295560# gnd! 42.7fF ;**FLOATING
C7 metal_221040_300120# gnd! 12.2fF ;**FLOATING
C8 metal_217320_298560# gnd! 9.4fF ;**FLOATING
C9 metal_8760_295200# gnd! 21.5fF ;**FLOATING
C10 metal_8760_299880# gnd! 20.6fF ;**FLOATING
C11 metal_207840_312240# gnd! 134.1fF ;**FLOATING
C12 metal_166920_313920# gnd! 151.8fF ;**FLOATING
C13 metal_107520_317040# gnd! 37.6fF ;**FLOATING
C14 metal_98520_313440# gnd! 38.1fF ;**FLOATING
C15 metal_92640_317040# gnd! 38.0fF ;**FLOATING
C16 metal_103440_313560# gnd! 38.0fF ;**FLOATING
C17 diff_191280_27720# gnd! 82.5fF
C18 diff_173520_28320# gnd! 104.2fF
C19 diff_202320_11520# gnd! 212.4fF
C20 diff_136080_6840# gnd! 85.9fF
C21 diff_129000_14040# gnd! 119.8fF
C22 diff_135360_28440# gnd! 77.1fF
C23 diff_117240_28320# gnd! 128.6fF
C24 diff_113400_27480# gnd! 197.8fF
C25 diff_172440_35400# gnd! 94.9fF
C26 diff_99000_21120# gnd! 105.5fF
C27 diff_182160_40080# gnd! 86.9fF
C28 diff_190680_39840# gnd! 60.1fF
C29 diff_165360_43680# gnd! 39.9fF
C30 diff_177480_41640# gnd! 335.3fF
C31 diff_182040_45240# gnd! 64.8fF
C32 diff_160800_42360# gnd! 150.7fF
C33 diff_152400_46440# gnd! 59.8fF
C34 diff_149640_49320# gnd! 48.3fF
C35 diff_56400_22080# gnd! 88.7fF
C36 diff_63960_26160# gnd! 444.0fF
C37 diff_95880_45240# gnd! 86.7fF
C38 diff_53880_29280# gnd! 91.2fF
C39 diff_30240_35160# gnd! 59.8fF
C40 diff_28200_35160# gnd! 33.9fF
C41 diff_53880_36240# gnd! 90.9fF
C42 diff_107760_44520# gnd! 164.9fF
C43 diff_131160_47160# gnd! 1041.0fF
C44 diff_142200_46080# gnd! 171.8fF
C45 diff_104520_47640# gnd! 243.3fF
C46 diff_28680_39960# gnd! 86.5fF
C47 diff_24240_43920# gnd! 85.9fF
C48 diff_27960_42600# gnd! 142.0fF
C49 diff_180240_49440# gnd! 95.6fF
C50 diff_168960_46920# gnd! 90.2fF
C51 diff_165120_55680# gnd! 43.2fF
C52 diff_197400_55440# gnd! 125.2fF
C53 diff_177480_52680# gnd! 315.8fF
C54 diff_182160_57120# gnd! 65.3fF
C55 diff_159360_54360# gnd! 176.4fF
C56 diff_143880_43920# gnd! 68.2fF
C57 diff_133800_49440# gnd! 88.5fF
C58 diff_30240_47160# gnd! 60.6fF
C59 diff_28080_47280# gnd! 34.7fF
C60 diff_87000_49080# gnd! 771.8fF
C61 diff_148680_53520# gnd! 563.6fF
C62 diff_152400_58560# gnd! 58.7fF
C63 diff_149640_61440# gnd! 48.7fF
C64 diff_104520_55560# gnd! 263.5fF
C65 diff_58920_54000# gnd! 131.4fF
C66 diff_28680_52080# gnd! 84.2fF
C67 diff_24240_55920# gnd! 85.4fF
C68 diff_27960_54240# gnd! 142.6fF
C69 diff_106800_59760# gnd! 296.2fF
C70 diff_143280_58080# gnd! 48.1fF
C71 diff_96120_61680# gnd! 72.1fF
C72 diff_179760_61200# gnd! 102.8fF
C73 diff_188160_64200# gnd! 65.0fF
C74 diff_165120_67680# gnd! 41.6fF
C75 diff_199440_72600# gnd! 96.8fF
C76 diff_177360_65880# gnd! 357.4fF
C77 diff_57120_59640# gnd! 150.3fF
C78 diff_49200_59400# gnd! 120.9fF
C79 diff_144360_54120# gnd! 408.9fF
C80 diff_87000_54000# gnd! 922.6fF
C81 diff_148680_65520# gnd! 98.7fF
C82 diff_182160_70080# gnd! 64.6fF
C83 diff_168720_72960# gnd! 99.4fF
C84 diff_43680_56040# gnd! 158.4fF
C85 diff_30240_59280# gnd! 62.6fF
C86 diff_160920_66360# gnd! 146.7fF
C87 diff_107760_66840# gnd! 165.7fF
C88 diff_153120_70680# gnd! 298.7fF
C89 diff_152400_72000# gnd! 54.9fF
C90 diff_149760_73320# gnd! 45.9fF
C91 diff_159360_66360# gnd! 233.5fF
C92 diff_131160_70440# gnd! 393.7fF
C93 diff_104520_69840# gnd! 236.1fF
C94 diff_142320_69960# gnd! 170.2fF
C95 diff_59280_61920# gnd! 159.3fF
C96 diff_28080_59280# gnd! 33.8fF
C97 diff_49440_63480# gnd! 100.5fF
C98 diff_133080_73080# gnd! 86.5fF
C99 diff_144000_67920# gnd! 69.5fF
C100 diff_179760_74400# gnd! 101.4fF
C101 diff_191520_73200# gnd! 232.0fF
C102 diff_188280_75600# gnd! 71.0fF
C103 diff_165240_79680# gnd! 41.2fF
C104 diff_159360_78360# gnd! 167.4fF
C105 diff_104520_77760# gnd! 260.1fF
C106 diff_90240_71400# gnd! 854.3fF
C107 diff_147720_75720# gnd! 351.7fF
C108 diff_148800_77640# gnd! 90.5fF
C109 diff_177480_79320# gnd! 245.3fF
C110 diff_177840_83640# gnd! 93.6fF
C111 diff_182880_82560# gnd! 60.2fF
C112 diff_153120_82680# gnd! 448.6fF
C113 diff_59400_45960# gnd! 403.0fF
C114 diff_28680_63960# gnd! 88.6fF
C115 diff_24120_68040# gnd! 87.0fF
C116 diff_27960_63360# gnd! 153.4fF
C117 diff_56400_73800# gnd! 115.4fF
C118 diff_70320_79920# gnd! 20.4fF
C119 diff_30240_71280# gnd! 65.2fF
C120 diff_28080_71160# gnd! 35.8fF
C121 diff_96000_83640# gnd! 72.9fF
C122 diff_106800_81960# gnd! 322.6fF
C123 diff_144480_78240# gnd! 159.2fF
C124 diff_152520_82440# gnd! 52.1fF
C125 diff_143280_82080# gnd! 47.1fF
C126 diff_150960_82320# gnd! 35.0fF
C127 diff_96720_85440# gnd! 78.2fF
C128 diff_175680_35880# gnd! 338.5fF
C129 diff_188040_90240# gnd! 78.5fF
C130 diff_178200_92400# gnd! 88.3fF
C131 diff_185640_97320# gnd! 41.1fF
C132 diff_194040_99480# gnd! 40.1fF
C133 diff_111960_24480# gnd! 1602.1fF
C134 diff_171960_95040# gnd! 60.1fF
C135 diff_176280_101040# gnd! 45.8fF
C136 diff_90240_74760# gnd! 912.3fF
C137 diff_119880_90240# gnd! 369.9fF
C138 diff_147840_90120# gnd! 120.3fF
C139 diff_132720_93000# gnd! 335.4fF
C140 diff_104520_92040# gnd! 269.8fF
C141 diff_118920_89640# gnd! 247.2fF
C142 diff_142920_94680# gnd! 98.3fF
C143 diff_106320_90480# gnd! 215.8fF
C144 diff_102480_94560# gnd! 34.0fF
C145 diff_131640_42480# gnd! 452.3fF
C146 diff_133440_86160# gnd! 188.7fF
C147 diff_193560_103560# gnd! 34.1fF
C148 diff_131760_92520# gnd! 192.2fF
C149 diff_165720_88920# gnd! 94.2fF
C150 diff_182640_101160# gnd! 137.4fF
C151 diff_174240_97200# gnd! 137.8fF
C152 diff_173520_107280# gnd! 92.4fF
C153 diff_218280_127680# gnd! 80.3fF
C154 diff_192360_116040# gnd! 46.1fF
C155 diff_185280_114120# gnd! 112.1fF
C156 diff_179880_112560# gnd! 131.3fF
C157 diff_213360_134760# gnd! 124.2fF
C158 diff_187800_118320# gnd! 178.1fF
C159 diff_188760_119280# gnd! 192.9fF
C160 diff_219720_138000# gnd! 84.2fF
C161 diff_134400_26040# gnd! 995.3fF
C162 diff_174480_111480# gnd! 157.8fF
C163 diff_128040_60120# gnd! 438.1fF
C164 diff_99120_25800# gnd! 440.3fF
C165 diff_126240_106680# gnd! 39.4fF
C166 diff_118080_91560# gnd! 660.1fF
C167 diff_117480_108840# gnd! 72.6fF
C168 diff_92160_93720# gnd! 106.1fF
C169 diff_86760_94560# gnd! 95.6fF
C170 diff_110280_107400# gnd! 426.8fF
C171 diff_97440_92520# gnd! 177.1fF
C172 diff_111720_106680# gnd! 59.9fF
C173 diff_131760_114840# gnd! 100.0fF
C174 diff_87360_101640# gnd! 541.7fF
C175 diff_90000_47280# gnd! 660.9fF
C176 diff_94440_111840# gnd! 70.4fF
C177 diff_108000_115920# gnd! 284.3fF
C178 diff_91800_105960# gnd! 194.4fF
C179 diff_28560_76560# gnd! 88.7fF
C180 diff_41040_77520# gnd! 76.0fF
C181 diff_24120_80040# gnd! 87.2fF
C182 diff_56400_79440# gnd! 121.0fF
C183 diff_62400_80640# gnd! 73.9fF
C184 diff_66480_87720# gnd! 31.7fF
C185 diff_62160_91320# gnd! 70.6fF
C186 diff_59040_94320# gnd! 124.1fF
C187 diff_48240_86520# gnd! 34.6fF
C188 diff_30240_84720# gnd! 62.7fF
C189 diff_28080_84600# gnd! 34.8fF
C190 diff_45240_90120# gnd! 60.6fF
C191 diff_47760_87000# gnd! 57.5fF
C192 diff_58680_100920# gnd! 88.4fF
C193 diff_28560_89520# gnd! 85.7fF
C194 diff_24120_93360# gnd! 87.2fF
C195 diff_27840_93120# gnd! 151.6fF
C196 diff_46680_91560# gnd! 175.1fF
C197 diff_94440_117120# gnd! 158.3fF
C198 diff_104880_119520# gnd! 421.6fF
C199 diff_99120_118920# gnd! 325.7fF
C200 diff_87480_109680# gnd! 123.6fF
C201 diff_60000_105000# gnd! 23.1fF
C202 diff_58440_105000# gnd! 22.7fF
C203 diff_58800_94080# gnd! 242.7fF
C204 diff_55200_105000# gnd! 20.4fF
C205 diff_60720_104520# gnd! 119.8fF
C206 diff_49560_105120# gnd! 48.1fF
C207 diff_30240_96720# gnd! 62.5fF
C208 diff_27960_96720# gnd! 37.0fF
C209 diff_51120_105120# gnd! 45.8fF
C210 diff_54240_108720# gnd! 142.3fF
C211 diff_98880_123960# gnd! 963.4fF
C212 diff_44280_73320# gnd! 886.7fF
C213 diff_84120_123480# gnd! 51.5fF
C214 diff_86760_128040# gnd! 49.4fF
C215 diff_28560_101520# gnd! 83.6fF
C216 diff_24120_105360# gnd! 86.1fF
C217 diff_65160_119400# gnd! 36.1fF
C218 diff_54720_116400# gnd! 95.2fF
C219 diff_63480_120120# gnd! 24.7fF
C220 diff_30240_108840# gnd! 63.8fF
C221 diff_27960_108600# gnd! 36.0fF
C222 diff_28560_113400# gnd! 81.1fF
C223 diff_24000_117480# gnd! 83.9fF
C224 diff_27840_112800# gnd! 157.3fF
C225 diff_65040_121200# gnd! 128.7fF
C226 diff_52200_120960# gnd! 19.4fF
C227 diff_45720_111480# gnd! 430.5fF
C228 diff_43560_89160# gnd! 299.5fF
C229 diff_56040_120960# gnd! 49.8fF
C230 diff_60720_122640# gnd! 73.3fF
C231 diff_84000_131040# gnd! 44.6fF
C232 diff_67080_124440# gnd! 35.7fF
C233 diff_70080_125040# gnd! 45.2fF
C234 diff_71040_129240# gnd! 31.2fF
C235 diff_28560_123960# gnd! 84.8fF
C236 diff_46320_121200# gnd! 54.0fF
C237 diff_41160_121200# gnd! 274.2fF
C238 diff_64680_127080# gnd! 98.7fF
C239 diff_74160_129960# gnd! 113.6fF
C240 diff_102000_133320# gnd! 448.6fF
C241 diff_55200_81120# gnd! 972.3fF
C242 diff_177960_117720# gnd! 230.2fF
C243 diff_84120_135360# gnd! 50.7fF
C244 diff_89400_137160# gnd! 541.2fF
C245 diff_76560_120480# gnd! 575.5fF
C246 diff_172560_117720# gnd! 235.2fF
C247 diff_183360_117720# gnd! 250.2fF
C248 diff_168960_143880# gnd! 30.7fF
C249 diff_77400_140520# gnd! 99.4fF
C250 diff_72120_132600# gnd! 594.2fF
C251 diff_75840_138120# gnd! 90.9fF
C252 diff_70560_140880# gnd! 200.9fF
C253 diff_27840_125040# gnd! 154.4fF
C254 diff_42960_134880# gnd! 298.9fF
C255 diff_66000_140160# gnd! 76.9fF
C256 diff_52440_136080# gnd! 35.1fF
C257 diff_27480_130800# gnd! 93.6fF
C258 diff_26040_133800# gnd! 57.9fF
C259 diff_30720_135000# gnd! 81.2fF
C260 diff_30000_135120# gnd! 151.9fF
C261 diff_53040_136920# gnd! 40.1fF
C262 diff_56400_140040# gnd! 79.6fF
C263 diff_60720_140760# gnd! 120.1fF
C264 diff_183600_148680# gnd! 18.4fF
C265 diff_180360_148200# gnd! 46.1fF
C266 diff_178560_149760# gnd! 55.4fF
C267 diff_159360_93840# gnd! 300.8fF
C268 diff_70080_105840# gnd! 724.7fF
C269 diff_165480_110160# gnd! 574.2fF
C270 diff_189960_159840# gnd! 58.2fF
C271 diff_178200_162000# gnd! 213.2fF
C272 diff_115920_125040# gnd! 271.6fF
C273 diff_106440_110160# gnd! 222.4fF
C274 diff_61320_141480# gnd! 24.6fF
C275 diff_55800_140760# gnd! 39.9fF
C276 diff_68400_139200# gnd! 60.3fF
C277 diff_55320_141960# gnd! 24.7fF
C278 diff_61320_143040# gnd! 25.8fF
C279 diff_41160_139680# gnd! 169.0fF
C280 diff_57000_124920# gnd! 193.1fF
C281 diff_74760_145920# gnd! 25.7fF
C282 diff_84840_148440# gnd! 57.3fF
C283 diff_55080_128160# gnd! 644.0fF
C284 diff_43560_137160# gnd! 53.3fF
C285 diff_66000_145440# gnd! 1005.0fF
C286 diff_49800_158880# gnd! 15.6fF
C287 diff_43800_159360# gnd! 60.6fF
C288 diff_168480_155400# gnd! 305.3fF
C289 diff_178200_154800# gnd! 276.6fF
C290 diff_208440_168000# gnd! 70.6fF
C291 diff_202560_165000# gnd! 114.6fF
C292 diff_197160_165000# gnd! 142.8fF
C293 diff_191760_165240# gnd! 162.7fF
C294 diff_209760_180360# gnd! 112.9fF
C295 diff_182160_172680# gnd! 199.2fF
C296 diff_182760_168000# gnd! 226.8fF
C297 diff_51360_158880# gnd! 141.8fF
C298 diff_173280_163200# gnd! 351.9fF
C299 diff_52680_161880# gnd! 33.2fF
C300 diff_52080_163800# gnd! 61.1fF
C301 diff_56040_162240# gnd! 123.7fF
C302 diff_58200_162360# gnd! 141.6fF
C303 diff_95160_164880# gnd! 202.3fF
C304 diff_207360_185520# gnd! 63.1fF
C305 diff_203520_184560# gnd! 16.6fF
C306 diff_207360_187080# gnd! 24.2fF
C307 diff_207360_188640# gnd! 27.5fF
C308 diff_195360_185760# gnd! 22.9fF
C309 diff_196920_186240# gnd! 87.0fF
C310 diff_65520_142080# gnd! 271.0fF
C311 diff_69720_171360# gnd! 894.8fF
C312 diff_47160_165840# gnd! 119.6fF
C313 diff_97800_109440# gnd! 452.4fF
C314 diff_206520_194880# gnd! 21.4fF
C315 diff_178920_94920# gnd! 805.8fF
C316 diff_201120_185760# gnd! 85.8fF
C317 diff_205680_196560# gnd! 26.8fF
C318 diff_205680_198000# gnd! 65.2fF
C319 diff_193320_187440# gnd! 96.4fF
C320 diff_180360_194040# gnd! 40.9fF
C321 diff_183600_181920# gnd! 216.0fF
C322 diff_179760_181440# gnd! 227.8fF
C323 diff_180120_190560# gnd! 152.5fF
C324 diff_176040_194040# gnd! 57.9fF
C325 diff_170880_192840# gnd! 18.1fF
C326 diff_169320_193320# gnd! 43.1fF
C327 diff_163800_185160# gnd! 18.1fF
C328 diff_159960_184200# gnd! 26.6fF
C329 diff_89160_121200# gnd! 470.4fF
C330 diff_165360_185160# gnd! 60.0fF
C331 diff_163800_191040# gnd! 18.1fF
C332 diff_159960_191040# gnd! 18.9fF
C333 diff_141720_184920# gnd! 152.6fF
C334 diff_82080_164400# gnd! 270.9fF
C335 diff_145200_181200# gnd! 57.6fF
C336 diff_148680_185160# gnd! 90.7fF
C337 diff_143400_186720# gnd! 70.1fF
C338 diff_153120_191040# gnd! 66.2fF
C339 diff_158400_186360# gnd! 62.6fF
C340 diff_174480_194280# gnd! 48.8fF
C341 diff_149880_184080# gnd! 167.8fF
C342 diff_153120_192360# gnd! 21.4fF
C343 diff_143400_188160# gnd! 58.2fF
C344 diff_135600_194640# gnd! 33.9fF
C345 diff_130080_189840# gnd! 35.1fF
C346 diff_89400_129240# gnd! 1261.1fF
C347 diff_128520_190200# gnd! 70.2fF
C348 diff_135600_195960# gnd! 121.5fF
C349 diff_198960_207240# gnd! 57.2fF
C350 diff_191520_202680# gnd! 103.8fF
C351 diff_181440_206520# gnd! 102.9fF
C352 diff_182160_210000# gnd! 100.7fF
C353 diff_180360_195360# gnd! 200.7fF
C354 diff_192240_207600# gnd! 318.6fF
C355 diff_200880_213960# gnd! 23.3fF
C356 diff_156600_191160# gnd! 159.7fF
C357 diff_123480_192240# gnd! 18.1fF
C358 diff_84720_181920# gnd! 20.4fF
C359 diff_118320_192240# gnd! 15.5fF
C360 diff_121680_193680# gnd! 21.5fF
C361 diff_120240_185760# gnd! 304.8fF
C362 diff_137400_197640# gnd! 87.6fF
C363 diff_141240_199080# gnd! 73.5fF
C364 diff_170760_206520# gnd! 97.0fF
C365 diff_162960_208080# gnd! 181.5fF
C366 diff_167280_200280# gnd! 120.0fF
C367 diff_174480_199320# gnd! 141.5fF
C368 diff_196440_216960# gnd! 37.2fF
C369 diff_188760_215400# gnd! 172.3fF
C370 diff_182880_214080# gnd! 25.6fF
C371 diff_182160_213240# gnd! 45.4fF
C372 diff_183120_215520# gnd! 178.4fF
C373 diff_188280_216360# gnd! 88.5fF
C374 diff_176640_214080# gnd! 23.2fF
C375 diff_119880_192240# gnd! 90.6fF
C376 diff_115200_193800# gnd! 64.4fF
C377 diff_110640_192240# gnd! 21.5fF
C378 diff_109080_192240# gnd! 21.4fF
C379 diff_90600_186120# gnd! 15.6fF
C380 diff_84720_183480# gnd! 141.8fF
C381 diff_83040_186840# gnd! 70.6fF
C382 diff_71760_186600# gnd! 15.6fF
C383 diff_71640_183960# gnd! 80.2fF
C384 diff_105120_200040# gnd! 20.9fF
C385 diff_84720_180000# gnd! 252.0fF
C386 diff_106680_199920# gnd! 27.4fF
C387 diff_158520_214320# gnd! 23.4fF
C388 diff_152280_214200# gnd! 23.3fF
C389 diff_175200_217320# gnd! 53.2fF
C390 diff_172080_217080# gnd! 36.4fF
C391 diff_109680_203520# gnd! 216.0fF
C392 diff_89040_188280# gnd! 644.9fF
C393 diff_124200_197520# gnd! 77.6fF
C394 diff_116040_208080# gnd! 21.8fF
C395 diff_115080_208680# gnd! 42.3fF
C396 diff_102600_202200# gnd! 89.1fF
C397 diff_112200_208080# gnd! 21.9fF
C398 diff_157920_213240# gnd! 48.3fF
C399 diff_134640_214200# gnd! 23.3fF
C400 diff_164520_215520# gnd! 274.1fF
C401 diff_158880_215640# gnd! 329.8fF
C402 diff_148200_217200# gnd! 36.1fF
C403 diff_133320_215640# gnd! 210.8fF
C404 diff_134040_213360# gnd! 46.8fF
C405 diff_134880_217080# gnd! 329.4fF
C406 diff_110640_210960# gnd! 35.8fF
C407 diff_117120_215640# gnd! 49.0fF
C408 diff_90840_198360# gnd! 120.9fF
C409 diff_72240_189360# gnd! 252.5fF
C410 diff_44040_172320# gnd! 119.4fF
C411 diff_49320_172200# gnd! 80.8fF
C412 diff_56280_181320# gnd! 23.3fF
C413 diff_50880_179400# gnd! 157.8fF
C414 diff_52440_182520# gnd! 27.4fF
C415 diff_47160_181560# gnd! 24.1fF
C416 diff_45600_181560# gnd! 24.6fF
C417 diff_44520_147840# gnd! 424.5fF
C418 diff_73200_192960# gnd! 60.0fF
C419 diff_74040_202080# gnd! 32.5fF
C420 diff_64920_198240# gnd! 113.0fF
C421 diff_66840_200160# gnd! 44.1fF
C422 diff_75120_202800# gnd! 129.5fF
C423 diff_77400_204960# gnd! 68.1fF
C424 diff_95880_204840# gnd! 107.8fF
C425 diff_92760_202560# gnd! 60.5fF
C426 diff_86640_208320# gnd! 77.8fF
C427 diff_70800_207960# gnd! 42.3fF
C428 diff_70800_206280# gnd! 221.4fF
C429 diff_52440_194280# gnd! 21.4fF
C430 diff_49320_194400# gnd! 20.4fF
C431 diff_45480_194400# gnd! 21.2fF
C432 diff_43800_194280# gnd! 24.2fF
C433 diff_51480_191880# gnd! 622.9fF
C434 diff_53040_193920# gnd! 260.0fF
C435 diff_44520_186120# gnd! 674.9fF
C436 diff_50880_194400# gnd! 65.4fF
C437 diff_49320_199200# gnd! 21.4fF
C438 diff_47040_199200# gnd! 40.9fF
C439 diff_64080_204360# gnd! 53.8fF
C440 diff_45720_176880# gnd! 174.5fF
C441 diff_80640_207120# gnd! 85.8fF
C442 diff_56520_205560# gnd! 95.5fF
C443 diff_57000_209520# gnd! 248.8fF
C444 diff_99360_215760# gnd! 180.5fF
C445 diff_164040_216360# gnd! 93.0fF
C446 diff_140640_215520# gnd! 276.9fF
C447 diff_140160_216480# gnd! 89.5fF
C448 diff_138120_220200# gnd! 498.3fF
C449 diff_188880_226560# gnd! 658.6fF
C450 diff_170640_228120# gnd! 118.8fF
C451 diff_161040_229440# gnd! 120.9fF
C452 diff_156120_226800# gnd! 119.8fF
C453 diff_151680_228720# gnd! 120.0fF
C454 diff_146760_226200# gnd! 119.3fF
C455 diff_133560_222480# gnd! 344.8fF
C456 diff_116040_220560# gnd! 21.6fF
C457 diff_87600_213720# gnd! 116.0fF
C458 diff_112200_220320# gnd! 22.6fF
C459 diff_82680_213840# gnd! 115.2fF
C460 diff_78120_219240# gnd! 116.5fF
C461 diff_73200_214320# gnd! 120.1fF
C462 diff_83400_222240# gnd! 143.3fF
C463 diff_115080_221040# gnd! 44.5fF
C464 diff_110640_223320# gnd! 36.8fF
C465 diff_74880_222120# gnd! 139.7fF
C466 diff_16920_200160# gnd! 77.0fF
C467 diff_21960_203880# gnd! 30.8fF
C468 diff_19080_201840# gnd! 52.9fF
C469 diff_20640_113640# gnd! 4117.4fF
C470 diff_30480_212760# gnd! 170.8fF
C471 diff_35040_214560# gnd! 123.4fF
C472 diff_110160_224880# gnd! 456.4fF
C473 diff_117120_227880# gnd! 49.0fF
C474 diff_99360_217440# gnd! 180.6fF
C475 diff_110040_208680# gnd! 309.5fF
C476 diff_110040_229200# gnd! 143.2fF
C477 diff_142320_226920# gnd! 119.4fF
C478 diff_137400_226080# gnd! 121.7fF
C479 diff_143160_236160# gnd! 257.8fF
C480 diff_38760_219600# gnd! 115.5fF
C481 diff_20760_213720# gnd! 86.2fF
C482 diff_23400_208080# gnd! 150.0fF
C483 diff_22800_212640# gnd! 101.2fF
C484 diff_58200_222720# gnd! 35.9fF
C485 diff_65760_223560# gnd! 36.7fF
C486 diff_62040_223560# gnd! 35.6fF
C487 diff_116040_234240# gnd! 22.3fF
C488 diff_164160_221520# gnd! 266.8fF
C489 diff_115080_234840# gnd! 43.5fF
C490 diff_112200_234120# gnd! 22.7fF
C491 diff_83160_218280# gnd! 179.7fF
C492 diff_110640_237120# gnd! 36.1fF
C493 diff_148080_240000# gnd! 250.8fF
C494 diff_138120_242040# gnd! 283.8fF
C495 diff_183360_241080# gnd! 198.4fF
C496 diff_69480_207240# gnd! 355.3fF
C497 diff_34560_231000# gnd! 88.1fF
C498 diff_63960_210840# gnd! 503.5fF
C499 diff_77640_236160# gnd! 191.6fF
C500 diff_72840_236280# gnd! 197.5fF
C501 diff_77640_238440# gnd! 85.4fF
C502 diff_71760_233040# gnd! 105.9fF
C503 diff_41520_198840# gnd! 341.4fF
C504 diff_117120_241680# gnd! 48.7fF
C505 diff_94080_215520# gnd! 234.8fF
C506 diff_128520_243360# gnd! 91.6fF
C507 diff_165720_226080# gnd! 357.5fF
C508 diff_176640_255840# gnd! 96.9fF
C509 diff_128520_245400# gnd! 93.0fF
C510 diff_161160_232920# gnd! 227.6fF
C511 diff_156720_230520# gnd! 229.8fF
C512 diff_116040_246960# gnd! 22.3fF
C513 diff_112200_247080# gnd! 22.0fF
C514 diff_115080_246600# gnd! 49.8fF
C515 diff_110640_249960# gnd! 41.4fF
C516 diff_93960_243360# gnd! 17.2fF
C517 diff_86400_243000# gnd! 17.6fF
C518 diff_82680_243840# gnd! 18.7fF
C519 diff_92160_246000# gnd! 27.2fF
C520 diff_87000_243000# gnd! 27.0fF
C521 diff_75120_243120# gnd! 16.9fF
C522 diff_39480_231000# gnd! 45.1fF
C523 diff_32040_231840# gnd! 100.2fF
C524 diff_40560_232800# gnd! 47.5fF
C525 diff_44400_224400# gnd! 279.2fF
C526 diff_21360_45480# gnd! 2310.6fF
C527 diff_21360_57480# gnd! 2453.1fF
C528 diff_35040_230160# gnd! 80.2fF
C529 diff_39480_236280# gnd! 37.8fF
C530 diff_11280_215400# gnd! 2539.5fF
C531 diff_81000_246000# gnd! 26.1fF
C532 diff_75840_243000# gnd! 26.0fF
C533 diff_93960_249000# gnd! 16.4fF
C534 diff_92160_247440# gnd! 27.1fF
C535 diff_105120_208440# gnd! 439.0fF
C536 diff_139680_251040# gnd! 836.3fF
C537 diff_147480_249360# gnd! 94.7fF
C538 diff_141600_255960# gnd! 95.4fF
C539 diff_117120_254520# gnd! 49.8fF
C540 diff_94080_217680# gnd! 262.1fF
C541 diff_134880_253320# gnd! 108.1fF
C542 diff_133560_235080# gnd! 2628.3fF
C543 diff_179520_261120# gnd! 14.5fF
C544 diff_172080_260640# gnd! 16.3fF
C545 diff_168360_261840# gnd! 15.7fF
C546 diff_177840_263520# gnd! 30.7fF
C547 diff_172680_260520# gnd! 28.2fF
C548 diff_160800_260640# gnd! 18.1fF
C549 diff_157200_261120# gnd! 18.0fF
C550 diff_166680_263640# gnd! 27.7fF
C551 diff_161520_260520# gnd! 26.4fF
C552 diff_179520_266520# gnd! 16.7fF
C553 diff_177840_265080# gnd! 28.2fF
C554 diff_179520_270000# gnd! 14.4fF
C555 diff_171960_268200# gnd! 15.8fF
C556 diff_168360_266520# gnd! 16.6fF
C557 diff_149640_260640# gnd! 18.4fF
C558 diff_146040_261120# gnd! 17.9fF
C559 diff_110040_234240# gnd! 329.1fF
C560 diff_109800_255840# gnd! 149.4fF
C561 diff_155520_263640# gnd! 26.3fF
C562 diff_150360_260520# gnd! 25.8fF
C563 diff_172560_268320# gnd! 27.9fF
C564 diff_166680_265080# gnd! 26.9fF
C565 diff_161520_265080# gnd! 27.0fF
C566 diff_160800_268080# gnd! 16.2fF
C567 diff_157200_266640# gnd! 16.8fF
C568 diff_138480_260760# gnd! 16.4fF
C569 diff_144240_263640# gnd! 26.6fF
C570 diff_139080_260640# gnd! 26.8fF
C571 diff_155520_265080# gnd! 26.4fF
C572 diff_171960_269520# gnd! 16.3fF
C573 diff_168360_270000# gnd! 16.3fF
C574 diff_177840_272520# gnd! 28.3fF
C575 diff_172680_269400# gnd! 26.9fF
C576 diff_160800_269520# gnd! 18.0fF
C577 diff_157200_270000# gnd! 17.3fF
C578 diff_149640_268200# gnd! 16.9fF
C579 diff_146040_266640# gnd! 16.8fF
C580 diff_150240_268320# gnd! 28.8fF
C581 diff_166680_272520# gnd! 26.8fF
C582 diff_161400_269520# gnd! 26.4fF
C583 diff_179520_275400# gnd! 14.9fF
C584 diff_177840_273960# gnd! 28.2fF
C585 diff_179520_278760# gnd! 13.9fF
C586 diff_171960_276960# gnd! 17.8fF
C587 diff_168360_275520# gnd! 15.8fF
C588 diff_172680_273960# gnd! 25.3fF
C589 diff_144240_265200# gnd! 25.4fF
C590 diff_149640_269640# gnd! 17.8fF
C591 diff_146040_270000# gnd! 16.7fF
C592 diff_138480_268200# gnd! 16.4fF
C593 diff_93960_252240# gnd! 16.8fF
C594 diff_86400_250320# gnd! 16.5fF
C595 diff_82800_249000# gnd! 16.4fF
C596 diff_87000_250680# gnd! 27.7fF
C597 diff_81000_247440# gnd! 26.6fF
C598 diff_75120_250560# gnd! 17.0fF
C599 diff_40440_238080# gnd! 52.5fF
C600 diff_54240_245520# gnd! 288.2fF
C601 diff_75840_250680# gnd! 26.6fF
C602 diff_82680_252360# gnd! 17.9fF
C603 diff_86400_251880# gnd! 17.7fF
C604 diff_92160_254880# gnd! 27.0fF
C605 diff_87000_251880# gnd! 26.3fF
C606 diff_75120_251880# gnd! 17.9fF
C607 diff_81000_254880# gnd! 25.9fF
C608 diff_93960_257880# gnd! 17.3fF
C609 diff_75840_251880# gnd! 26.4fF
C610 diff_92160_256320# gnd! 26.6fF
C611 diff_139080_268320# gnd! 27.8fF
C612 diff_155520_272520# gnd! 26.4fF
C613 diff_150360_269400# gnd! 26.8fF
C614 diff_166680_273960# gnd! 26.7fF
C615 diff_160800_276960# gnd! 16.7fF
C616 diff_157200_275520# gnd! 16.4fF
C617 diff_161400_277200# gnd! 26.1fF
C618 diff_138480_269640# gnd! 16.5fF
C619 diff_144240_272520# gnd! 26.8fF
C620 diff_139080_269520# gnd! 26.8fF
C621 diff_155400_274320# gnd! 26.2fF
C622 diff_171960_278400# gnd! 17.5fF
C623 diff_168360_278880# gnd! 14.8fF
C624 diff_177840_281280# gnd! 30.6fF
C625 diff_172680_278280# gnd! 26.4fF
C626 diff_179520_284280# gnd! 14.2fF
C627 diff_160800_278400# gnd! 17.7fF
C628 diff_157200_278880# gnd! 16.1fF
C629 diff_149640_276960# gnd! 16.4fF
C630 diff_146040_275520# gnd! 16.7fF
C631 diff_150240_277080# gnd! 25.8fF
C632 diff_144240_273960# gnd! 27.7fF
C633 diff_166560_281400# gnd! 27.4fF
C634 diff_161400_278280# gnd! 25.3fF
C635 diff_177840_282840# gnd! 28.8fF
C636 diff_149640_278400# gnd! 17.3fF
C637 diff_138480_276960# gnd! 16.4fF
C638 diff_139080_277080# gnd! 25.9fF
C639 diff_145920_280320# gnd! 16.8fF
C640 diff_155400_281400# gnd! 27.2fF
C641 diff_150240_278280# gnd! 25.6fF
C642 diff_171960_285840# gnd! 17.2fF
C643 diff_179520_287640# gnd! 13.7fF
C644 diff_172680_282840# gnd! 25.3fF
C645 diff_168360_284280# gnd! 14.9fF
C646 diff_166560_282840# gnd! 27.8fF
C647 diff_171960_287280# gnd! 17.3fF
C648 diff_168360_287640# gnd! 13.9fF
C649 diff_160800_285840# gnd! 17.4fF
C650 diff_138360_278640# gnd! 16.7fF
C651 diff_144240_281400# gnd! 26.6fF
C652 diff_139080_278280# gnd! 26.4fF
C653 diff_157080_284280# gnd! 17.6fF
C654 diff_161400_286080# gnd! 25.2fF
C655 diff_155400_282840# gnd! 26.8fF
C656 diff_172680_287040# gnd! 27.6fF
C657 diff_174360_263520# gnd! 226.3fF
C658 diff_149520_286080# gnd! 17.4fF
C659 diff_145920_284400# gnd! 17.8fF
C660 diff_150240_286080# gnd! 26.4fF
C661 diff_160800_287280# gnd! 16.7fF
C662 diff_157200_287760# gnd! 14.5fF
C663 diff_166560_290280# gnd! 29.2fF
C664 diff_161400_287160# gnd! 25.6fF
C665 diff_179520_293160# gnd! 13.7fF
C666 diff_177840_291720# gnd! 28.4fF
C667 diff_172440_294840# gnd! 28.9fF
C668 diff_171960_294720# gnd! 14.3fF
C669 diff_168360_293160# gnd! 14.4fF
C670 diff_179280_254400# gnd! 239.8fF
C671 diff_144240_282840# gnd! 26.2fF
C672 diff_149520_287400# gnd! 16.7fF
C673 diff_145920_287880# gnd! 17.1fF
C674 diff_138360_286080# gnd! 16.6fF
C675 diff_109920_264000# gnd! 263.4fF
C676 diff_86400_259200# gnd! 18.2fF
C677 diff_82680_258240# gnd! 18.9fF
C678 diff_87000_259560# gnd! 26.0fF
C679 diff_81000_256320# gnd! 25.9fF
C680 diff_93960_261240# gnd! 16.6fF
C681 diff_86400_260760# gnd! 18.7fF
C682 diff_75120_259560# gnd! 16.5fF
C683 diff_75840_259440# gnd! 26.8fF
C684 diff_82680_261240# gnd! 19.8fF
C685 diff_92160_263760# gnd! 27.5fF
C686 diff_87000_260760# gnd! 26.5fF
C687 diff_75120_260760# gnd! 18.0fF
C688 diff_81000_263760# gnd! 24.5fF
C689 diff_75840_260760# gnd! 26.2fF
C690 diff_93960_266640# gnd! 17.6fF
C691 diff_92160_265200# gnd! 27.1fF
C692 diff_93960_270120# gnd! 17.7fF
C693 diff_86280_268320# gnd! 18.3fF
C694 diff_82680_266760# gnd! 18.8fF
C695 diff_87000_268440# gnd! 26.8fF
C696 diff_81000_265200# gnd! 24.7fF
C697 diff_86400_269640# gnd! 19.4fF
C698 diff_82800_269880# gnd! 17.9fF
C699 diff_75840_268440# gnd! 27.1fF
C700 diff_75120_268440# gnd! 16.5fF
C701 diff_92160_272640# gnd! 26.7fF
C702 diff_87000_269640# gnd! 25.2fF
C703 diff_75120_269640# gnd! 17.5fF
C704 diff_81000_272640# gnd! 26.2fF
C705 diff_75840_269640# gnd! 27.4fF
C706 diff_93960_275640# gnd! 17.4fF
C707 diff_92160_274080# gnd! 26.4fF
C708 diff_138960_286080# gnd! 27.0fF
C709 diff_155400_290280# gnd! 27.9fF
C710 diff_150240_287160# gnd! 26.1fF
C711 diff_138360_287280# gnd! 17.9fF
C712 diff_144240_290280# gnd! 27.5fF
C713 diff_138960_287280# gnd! 26.4fF
C714 diff_153840_254520# gnd! 216.0fF
C715 diff_151440_254520# gnd! 216.4fF
C716 diff_142200_254520# gnd! 215.5fF
C717 diff_139680_254520# gnd! 217.5fF
C718 diff_166560_291720# gnd! 29.6fF
C719 diff_167640_254400# gnd! 229.8fF
C720 diff_160800_294960# gnd! 14.5fF
C721 diff_157200_293280# gnd! 13.7fF
C722 diff_161280_294840# gnd! 27.8fF
C723 diff_155400_291720# gnd! 29.1fF
C724 diff_149640_294720# gnd! 16.8fF
C725 diff_146040_293280# gnd! 14.3fF
C726 diff_150240_291840# gnd! 26.8fF
C727 diff_144240_291720# gnd! 28.7fF
C728 diff_138480_294720# gnd! 14.8fF
C729 diff_93960_279120# gnd! 18.2fF
C730 diff_86400_276960# gnd! 18.3fF
C731 diff_82800_275640# gnd! 16.8fF
C732 diff_87000_277320# gnd! 26.4fF
C733 diff_81000_274080# gnd! 26.9fF
C734 diff_117960_280920# gnd! 343.9fF
C735 diff_86400_278520# gnd! 19.3fF
C736 diff_82680_279240# gnd! 17.9fF
C737 diff_75840_277320# gnd! 28.0fF
C738 diff_75240_277200# gnd! 15.8fF
C739 diff_92280_281520# gnd! 26.5fF
C740 diff_87000_278520# gnd! 25.3fF
C741 diff_75120_278520# gnd! 17.7fF
C742 diff_81000_281520# gnd! 26.0fF
C743 diff_75840_278520# gnd! 27.6fF
C744 diff_93960_284400# gnd! 18.2fF
C745 diff_92280_282960# gnd! 25.7fF
C746 diff_93960_288000# gnd! 17.6fF
C747 diff_86400_286080# gnd! 18.9fF
C748 diff_82800_284400# gnd! 18.3fF
C749 diff_87120_286080# gnd! 26.1fF
C750 diff_117840_290880# gnd! 359.5fF
C751 diff_123240_258000# gnd! 503.7fF
C752 diff_117960_263280# gnd! 8796.1fF
C753 diff_171480_208680# gnd! 566.0fF
C754 diff_81000_282960# gnd! 26.0fF
C755 diff_86400_287400# gnd! 19.3fF
C756 diff_82800_287520# gnd! 18.6fF
C757 diff_75240_286080# gnd! 16.0fF
C758 diff_75840_286320# gnd! 28.7fF
C759 diff_92280_290400# gnd! 27.0fF
C760 diff_87000_287520# gnd! 26.0fF
C761 diff_75120_287520# gnd! 17.4fF
C762 diff_81000_290400# gnd! 26.3fF
C763 diff_75840_287400# gnd! 28.2fF
C764 diff_78120_238200# gnd! 302.8fF
C765 diff_75720_237120# gnd! 300.4fF
C766 diff_93960_293280# gnd! 17.9fF
C767 diff_86760_205920# gnd! 619.5fF
C768 diff_92280_291840# gnd! 24.1fF
C769 diff_86400_294960# gnd! 14.9fF
C770 diff_82800_293280# gnd! 17.4fF
C771 diff_87000_295200# gnd! 29.0fF
C772 diff_81000_291840# gnd! 24.7fF
C773 diff_85440_237000# gnd! 300.7fF
C774 diff_28320_238920# gnd! 135.9fF
C775 diff_42000_244200# gnd! 347.3fF
C776 diff_36120_243120# gnd! 103.7fF
C777 diff_40680_247920# gnd! 85.8fF
C778 diff_26760_254160# gnd! 149.6fF
C779 diff_24720_254040# gnd! 130.4fF
C780 diff_24240_254880# gnd! 209.0fF
C781 diff_54240_263880# gnd! 282.9fF
C782 diff_54240_272160# gnd! 281.8fF
C783 diff_60240_235200# gnd! 328.7fF
C784 diff_29760_255720# gnd! 12.7fF
C785 diff_26760_255720# gnd! 16.6fF
C786 diff_24720_255720# gnd! 9.8fF
C787 diff_40680_263760# gnd! 83.9fF
C788 diff_42000_267240# gnd! 343.1fF
C789 diff_31320_260160# gnd! 191.6fF
C790 diff_36600_265200# gnd! 98.3fF
C791 diff_42000_270960# gnd! 348.2fF
C792 diff_29880_257280# gnd! 175.1fF
C793 diff_40800_274440# gnd! 86.2fF
C794 diff_4200_259560# gnd! 803.4fF
C795 diff_26760_257280# gnd! 115.3fF
C796 diff_24720_257280# gnd! 135.8fF
C797 diff_27240_279000# gnd! 194.9fF
C798 diff_27600_280080# gnd! 100.8fF
C799 diff_40800_290280# gnd! 91.2fF
C800 diff_64920_237000# gnd! 356.8fF
C801 diff_52080_238440# gnd! 397.9fF
C802 diff_50160_238320# gnd! 2180.7fF
C803 diff_42000_294000# gnd! 358.2fF
C804 diff_75240_295200# gnd! 16.5fF
C805 diff_75840_295200# gnd! 29.1fF
C806 diff_73440_237000# gnd! 306.9fF
C807 diff_51960_227760# gnd! 1443.7fF
C808 diff_51480_235440# gnd! 4651.0fF
C809 diff_28560_293760# gnd! 196.9fF
C810 diff_36720_291840# gnd! 95.9fF
C811 diff_26520_220920# gnd! 846.6fF
C812 test gnd! 1619.7fF
C813 reset gnd! 1652.9fF
